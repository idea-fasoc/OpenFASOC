* NGSPICE file created from diff_pair_sample_1362.ext - technology: sky130A

.subckt diff_pair_sample_1362 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=4.173 ps=22.18 w=10.7 l=0.74
X1 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=4.173 ps=22.18 w=10.7 l=0.74
X2 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=0.74
X3 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=0.74
X4 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=0.74
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=0 ps=0 w=10.7 l=0.74
X6 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=4.173 ps=22.18 w=10.7 l=0.74
X7 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.173 pd=22.18 as=4.173 ps=22.18 w=10.7 l=0.74
R0 VP.n0 VP.t0 601.612
R1 VP.n0 VP.t1 562.859
R2 VP VP.n0 0.0516364
R3 VTAIL.n226 VTAIL.n174 289.615
R4 VTAIL.n52 VTAIL.n0 289.615
R5 VTAIL.n168 VTAIL.n116 289.615
R6 VTAIL.n110 VTAIL.n58 289.615
R7 VTAIL.n193 VTAIL.n192 185
R8 VTAIL.n190 VTAIL.n189 185
R9 VTAIL.n199 VTAIL.n198 185
R10 VTAIL.n201 VTAIL.n200 185
R11 VTAIL.n186 VTAIL.n185 185
R12 VTAIL.n207 VTAIL.n206 185
R13 VTAIL.n210 VTAIL.n209 185
R14 VTAIL.n208 VTAIL.n182 185
R15 VTAIL.n215 VTAIL.n181 185
R16 VTAIL.n217 VTAIL.n216 185
R17 VTAIL.n219 VTAIL.n218 185
R18 VTAIL.n178 VTAIL.n177 185
R19 VTAIL.n225 VTAIL.n224 185
R20 VTAIL.n227 VTAIL.n226 185
R21 VTAIL.n19 VTAIL.n18 185
R22 VTAIL.n16 VTAIL.n15 185
R23 VTAIL.n25 VTAIL.n24 185
R24 VTAIL.n27 VTAIL.n26 185
R25 VTAIL.n12 VTAIL.n11 185
R26 VTAIL.n33 VTAIL.n32 185
R27 VTAIL.n36 VTAIL.n35 185
R28 VTAIL.n34 VTAIL.n8 185
R29 VTAIL.n41 VTAIL.n7 185
R30 VTAIL.n43 VTAIL.n42 185
R31 VTAIL.n45 VTAIL.n44 185
R32 VTAIL.n4 VTAIL.n3 185
R33 VTAIL.n51 VTAIL.n50 185
R34 VTAIL.n53 VTAIL.n52 185
R35 VTAIL.n169 VTAIL.n168 185
R36 VTAIL.n167 VTAIL.n166 185
R37 VTAIL.n120 VTAIL.n119 185
R38 VTAIL.n161 VTAIL.n160 185
R39 VTAIL.n159 VTAIL.n158 185
R40 VTAIL.n157 VTAIL.n123 185
R41 VTAIL.n127 VTAIL.n124 185
R42 VTAIL.n152 VTAIL.n151 185
R43 VTAIL.n150 VTAIL.n149 185
R44 VTAIL.n129 VTAIL.n128 185
R45 VTAIL.n144 VTAIL.n143 185
R46 VTAIL.n142 VTAIL.n141 185
R47 VTAIL.n133 VTAIL.n132 185
R48 VTAIL.n136 VTAIL.n135 185
R49 VTAIL.n111 VTAIL.n110 185
R50 VTAIL.n109 VTAIL.n108 185
R51 VTAIL.n62 VTAIL.n61 185
R52 VTAIL.n103 VTAIL.n102 185
R53 VTAIL.n101 VTAIL.n100 185
R54 VTAIL.n99 VTAIL.n65 185
R55 VTAIL.n69 VTAIL.n66 185
R56 VTAIL.n94 VTAIL.n93 185
R57 VTAIL.n92 VTAIL.n91 185
R58 VTAIL.n71 VTAIL.n70 185
R59 VTAIL.n86 VTAIL.n85 185
R60 VTAIL.n84 VTAIL.n83 185
R61 VTAIL.n75 VTAIL.n74 185
R62 VTAIL.n78 VTAIL.n77 185
R63 VTAIL.t1 VTAIL.n191 149.524
R64 VTAIL.t3 VTAIL.n17 149.524
R65 VTAIL.t2 VTAIL.n134 149.524
R66 VTAIL.t0 VTAIL.n76 149.524
R67 VTAIL.n192 VTAIL.n189 104.615
R68 VTAIL.n199 VTAIL.n189 104.615
R69 VTAIL.n200 VTAIL.n199 104.615
R70 VTAIL.n200 VTAIL.n185 104.615
R71 VTAIL.n207 VTAIL.n185 104.615
R72 VTAIL.n209 VTAIL.n207 104.615
R73 VTAIL.n209 VTAIL.n208 104.615
R74 VTAIL.n208 VTAIL.n181 104.615
R75 VTAIL.n217 VTAIL.n181 104.615
R76 VTAIL.n218 VTAIL.n217 104.615
R77 VTAIL.n218 VTAIL.n177 104.615
R78 VTAIL.n225 VTAIL.n177 104.615
R79 VTAIL.n226 VTAIL.n225 104.615
R80 VTAIL.n18 VTAIL.n15 104.615
R81 VTAIL.n25 VTAIL.n15 104.615
R82 VTAIL.n26 VTAIL.n25 104.615
R83 VTAIL.n26 VTAIL.n11 104.615
R84 VTAIL.n33 VTAIL.n11 104.615
R85 VTAIL.n35 VTAIL.n33 104.615
R86 VTAIL.n35 VTAIL.n34 104.615
R87 VTAIL.n34 VTAIL.n7 104.615
R88 VTAIL.n43 VTAIL.n7 104.615
R89 VTAIL.n44 VTAIL.n43 104.615
R90 VTAIL.n44 VTAIL.n3 104.615
R91 VTAIL.n51 VTAIL.n3 104.615
R92 VTAIL.n52 VTAIL.n51 104.615
R93 VTAIL.n168 VTAIL.n167 104.615
R94 VTAIL.n167 VTAIL.n119 104.615
R95 VTAIL.n160 VTAIL.n119 104.615
R96 VTAIL.n160 VTAIL.n159 104.615
R97 VTAIL.n159 VTAIL.n123 104.615
R98 VTAIL.n127 VTAIL.n123 104.615
R99 VTAIL.n151 VTAIL.n127 104.615
R100 VTAIL.n151 VTAIL.n150 104.615
R101 VTAIL.n150 VTAIL.n128 104.615
R102 VTAIL.n143 VTAIL.n128 104.615
R103 VTAIL.n143 VTAIL.n142 104.615
R104 VTAIL.n142 VTAIL.n132 104.615
R105 VTAIL.n135 VTAIL.n132 104.615
R106 VTAIL.n110 VTAIL.n109 104.615
R107 VTAIL.n109 VTAIL.n61 104.615
R108 VTAIL.n102 VTAIL.n61 104.615
R109 VTAIL.n102 VTAIL.n101 104.615
R110 VTAIL.n101 VTAIL.n65 104.615
R111 VTAIL.n69 VTAIL.n65 104.615
R112 VTAIL.n93 VTAIL.n69 104.615
R113 VTAIL.n93 VTAIL.n92 104.615
R114 VTAIL.n92 VTAIL.n70 104.615
R115 VTAIL.n85 VTAIL.n70 104.615
R116 VTAIL.n85 VTAIL.n84 104.615
R117 VTAIL.n84 VTAIL.n74 104.615
R118 VTAIL.n77 VTAIL.n74 104.615
R119 VTAIL.n192 VTAIL.t1 52.3082
R120 VTAIL.n18 VTAIL.t3 52.3082
R121 VTAIL.n135 VTAIL.t2 52.3082
R122 VTAIL.n77 VTAIL.t0 52.3082
R123 VTAIL.n231 VTAIL.n230 32.5732
R124 VTAIL.n57 VTAIL.n56 32.5732
R125 VTAIL.n173 VTAIL.n172 32.5732
R126 VTAIL.n115 VTAIL.n114 32.5732
R127 VTAIL.n115 VTAIL.n57 23.4531
R128 VTAIL.n231 VTAIL.n173 22.5307
R129 VTAIL.n216 VTAIL.n215 13.1884
R130 VTAIL.n42 VTAIL.n41 13.1884
R131 VTAIL.n158 VTAIL.n157 13.1884
R132 VTAIL.n100 VTAIL.n99 13.1884
R133 VTAIL.n214 VTAIL.n182 12.8005
R134 VTAIL.n219 VTAIL.n180 12.8005
R135 VTAIL.n40 VTAIL.n8 12.8005
R136 VTAIL.n45 VTAIL.n6 12.8005
R137 VTAIL.n161 VTAIL.n122 12.8005
R138 VTAIL.n156 VTAIL.n124 12.8005
R139 VTAIL.n103 VTAIL.n64 12.8005
R140 VTAIL.n98 VTAIL.n66 12.8005
R141 VTAIL.n211 VTAIL.n210 12.0247
R142 VTAIL.n220 VTAIL.n178 12.0247
R143 VTAIL.n37 VTAIL.n36 12.0247
R144 VTAIL.n46 VTAIL.n4 12.0247
R145 VTAIL.n162 VTAIL.n120 12.0247
R146 VTAIL.n153 VTAIL.n152 12.0247
R147 VTAIL.n104 VTAIL.n62 12.0247
R148 VTAIL.n95 VTAIL.n94 12.0247
R149 VTAIL.n206 VTAIL.n184 11.249
R150 VTAIL.n224 VTAIL.n223 11.249
R151 VTAIL.n32 VTAIL.n10 11.249
R152 VTAIL.n50 VTAIL.n49 11.249
R153 VTAIL.n166 VTAIL.n165 11.249
R154 VTAIL.n149 VTAIL.n126 11.249
R155 VTAIL.n108 VTAIL.n107 11.249
R156 VTAIL.n91 VTAIL.n68 11.249
R157 VTAIL.n205 VTAIL.n186 10.4732
R158 VTAIL.n227 VTAIL.n176 10.4732
R159 VTAIL.n31 VTAIL.n12 10.4732
R160 VTAIL.n53 VTAIL.n2 10.4732
R161 VTAIL.n169 VTAIL.n118 10.4732
R162 VTAIL.n148 VTAIL.n129 10.4732
R163 VTAIL.n111 VTAIL.n60 10.4732
R164 VTAIL.n90 VTAIL.n71 10.4732
R165 VTAIL.n193 VTAIL.n191 10.2747
R166 VTAIL.n19 VTAIL.n17 10.2747
R167 VTAIL.n136 VTAIL.n134 10.2747
R168 VTAIL.n78 VTAIL.n76 10.2747
R169 VTAIL.n202 VTAIL.n201 9.69747
R170 VTAIL.n228 VTAIL.n174 9.69747
R171 VTAIL.n28 VTAIL.n27 9.69747
R172 VTAIL.n54 VTAIL.n0 9.69747
R173 VTAIL.n170 VTAIL.n116 9.69747
R174 VTAIL.n145 VTAIL.n144 9.69747
R175 VTAIL.n112 VTAIL.n58 9.69747
R176 VTAIL.n87 VTAIL.n86 9.69747
R177 VTAIL.n230 VTAIL.n229 9.45567
R178 VTAIL.n56 VTAIL.n55 9.45567
R179 VTAIL.n172 VTAIL.n171 9.45567
R180 VTAIL.n114 VTAIL.n113 9.45567
R181 VTAIL.n229 VTAIL.n228 9.3005
R182 VTAIL.n176 VTAIL.n175 9.3005
R183 VTAIL.n223 VTAIL.n222 9.3005
R184 VTAIL.n221 VTAIL.n220 9.3005
R185 VTAIL.n180 VTAIL.n179 9.3005
R186 VTAIL.n195 VTAIL.n194 9.3005
R187 VTAIL.n197 VTAIL.n196 9.3005
R188 VTAIL.n188 VTAIL.n187 9.3005
R189 VTAIL.n203 VTAIL.n202 9.3005
R190 VTAIL.n205 VTAIL.n204 9.3005
R191 VTAIL.n184 VTAIL.n183 9.3005
R192 VTAIL.n212 VTAIL.n211 9.3005
R193 VTAIL.n214 VTAIL.n213 9.3005
R194 VTAIL.n55 VTAIL.n54 9.3005
R195 VTAIL.n2 VTAIL.n1 9.3005
R196 VTAIL.n49 VTAIL.n48 9.3005
R197 VTAIL.n47 VTAIL.n46 9.3005
R198 VTAIL.n6 VTAIL.n5 9.3005
R199 VTAIL.n21 VTAIL.n20 9.3005
R200 VTAIL.n23 VTAIL.n22 9.3005
R201 VTAIL.n14 VTAIL.n13 9.3005
R202 VTAIL.n29 VTAIL.n28 9.3005
R203 VTAIL.n31 VTAIL.n30 9.3005
R204 VTAIL.n10 VTAIL.n9 9.3005
R205 VTAIL.n38 VTAIL.n37 9.3005
R206 VTAIL.n40 VTAIL.n39 9.3005
R207 VTAIL.n138 VTAIL.n137 9.3005
R208 VTAIL.n140 VTAIL.n139 9.3005
R209 VTAIL.n131 VTAIL.n130 9.3005
R210 VTAIL.n146 VTAIL.n145 9.3005
R211 VTAIL.n148 VTAIL.n147 9.3005
R212 VTAIL.n126 VTAIL.n125 9.3005
R213 VTAIL.n154 VTAIL.n153 9.3005
R214 VTAIL.n156 VTAIL.n155 9.3005
R215 VTAIL.n171 VTAIL.n170 9.3005
R216 VTAIL.n118 VTAIL.n117 9.3005
R217 VTAIL.n165 VTAIL.n164 9.3005
R218 VTAIL.n163 VTAIL.n162 9.3005
R219 VTAIL.n122 VTAIL.n121 9.3005
R220 VTAIL.n80 VTAIL.n79 9.3005
R221 VTAIL.n82 VTAIL.n81 9.3005
R222 VTAIL.n73 VTAIL.n72 9.3005
R223 VTAIL.n88 VTAIL.n87 9.3005
R224 VTAIL.n90 VTAIL.n89 9.3005
R225 VTAIL.n68 VTAIL.n67 9.3005
R226 VTAIL.n96 VTAIL.n95 9.3005
R227 VTAIL.n98 VTAIL.n97 9.3005
R228 VTAIL.n113 VTAIL.n112 9.3005
R229 VTAIL.n60 VTAIL.n59 9.3005
R230 VTAIL.n107 VTAIL.n106 9.3005
R231 VTAIL.n105 VTAIL.n104 9.3005
R232 VTAIL.n64 VTAIL.n63 9.3005
R233 VTAIL.n198 VTAIL.n188 8.92171
R234 VTAIL.n24 VTAIL.n14 8.92171
R235 VTAIL.n141 VTAIL.n131 8.92171
R236 VTAIL.n83 VTAIL.n73 8.92171
R237 VTAIL.n197 VTAIL.n190 8.14595
R238 VTAIL.n23 VTAIL.n16 8.14595
R239 VTAIL.n140 VTAIL.n133 8.14595
R240 VTAIL.n82 VTAIL.n75 8.14595
R241 VTAIL.n194 VTAIL.n193 7.3702
R242 VTAIL.n20 VTAIL.n19 7.3702
R243 VTAIL.n137 VTAIL.n136 7.3702
R244 VTAIL.n79 VTAIL.n78 7.3702
R245 VTAIL.n194 VTAIL.n190 5.81868
R246 VTAIL.n20 VTAIL.n16 5.81868
R247 VTAIL.n137 VTAIL.n133 5.81868
R248 VTAIL.n79 VTAIL.n75 5.81868
R249 VTAIL.n198 VTAIL.n197 5.04292
R250 VTAIL.n24 VTAIL.n23 5.04292
R251 VTAIL.n141 VTAIL.n140 5.04292
R252 VTAIL.n83 VTAIL.n82 5.04292
R253 VTAIL.n201 VTAIL.n188 4.26717
R254 VTAIL.n230 VTAIL.n174 4.26717
R255 VTAIL.n27 VTAIL.n14 4.26717
R256 VTAIL.n56 VTAIL.n0 4.26717
R257 VTAIL.n172 VTAIL.n116 4.26717
R258 VTAIL.n144 VTAIL.n131 4.26717
R259 VTAIL.n114 VTAIL.n58 4.26717
R260 VTAIL.n86 VTAIL.n73 4.26717
R261 VTAIL.n202 VTAIL.n186 3.49141
R262 VTAIL.n228 VTAIL.n227 3.49141
R263 VTAIL.n28 VTAIL.n12 3.49141
R264 VTAIL.n54 VTAIL.n53 3.49141
R265 VTAIL.n170 VTAIL.n169 3.49141
R266 VTAIL.n145 VTAIL.n129 3.49141
R267 VTAIL.n112 VTAIL.n111 3.49141
R268 VTAIL.n87 VTAIL.n71 3.49141
R269 VTAIL.n195 VTAIL.n191 2.84303
R270 VTAIL.n21 VTAIL.n17 2.84303
R271 VTAIL.n138 VTAIL.n134 2.84303
R272 VTAIL.n80 VTAIL.n76 2.84303
R273 VTAIL.n206 VTAIL.n205 2.71565
R274 VTAIL.n224 VTAIL.n176 2.71565
R275 VTAIL.n32 VTAIL.n31 2.71565
R276 VTAIL.n50 VTAIL.n2 2.71565
R277 VTAIL.n166 VTAIL.n118 2.71565
R278 VTAIL.n149 VTAIL.n148 2.71565
R279 VTAIL.n108 VTAIL.n60 2.71565
R280 VTAIL.n91 VTAIL.n90 2.71565
R281 VTAIL.n210 VTAIL.n184 1.93989
R282 VTAIL.n223 VTAIL.n178 1.93989
R283 VTAIL.n36 VTAIL.n10 1.93989
R284 VTAIL.n49 VTAIL.n4 1.93989
R285 VTAIL.n165 VTAIL.n120 1.93989
R286 VTAIL.n152 VTAIL.n126 1.93989
R287 VTAIL.n107 VTAIL.n62 1.93989
R288 VTAIL.n94 VTAIL.n68 1.93989
R289 VTAIL.n211 VTAIL.n182 1.16414
R290 VTAIL.n220 VTAIL.n219 1.16414
R291 VTAIL.n37 VTAIL.n8 1.16414
R292 VTAIL.n46 VTAIL.n45 1.16414
R293 VTAIL.n162 VTAIL.n161 1.16414
R294 VTAIL.n153 VTAIL.n124 1.16414
R295 VTAIL.n104 VTAIL.n103 1.16414
R296 VTAIL.n95 VTAIL.n66 1.16414
R297 VTAIL.n173 VTAIL.n115 0.931535
R298 VTAIL VTAIL.n57 0.759121
R299 VTAIL.n215 VTAIL.n214 0.388379
R300 VTAIL.n216 VTAIL.n180 0.388379
R301 VTAIL.n41 VTAIL.n40 0.388379
R302 VTAIL.n42 VTAIL.n6 0.388379
R303 VTAIL.n158 VTAIL.n122 0.388379
R304 VTAIL.n157 VTAIL.n156 0.388379
R305 VTAIL.n100 VTAIL.n64 0.388379
R306 VTAIL.n99 VTAIL.n98 0.388379
R307 VTAIL VTAIL.n231 0.172914
R308 VTAIL.n196 VTAIL.n195 0.155672
R309 VTAIL.n196 VTAIL.n187 0.155672
R310 VTAIL.n203 VTAIL.n187 0.155672
R311 VTAIL.n204 VTAIL.n203 0.155672
R312 VTAIL.n204 VTAIL.n183 0.155672
R313 VTAIL.n212 VTAIL.n183 0.155672
R314 VTAIL.n213 VTAIL.n212 0.155672
R315 VTAIL.n213 VTAIL.n179 0.155672
R316 VTAIL.n221 VTAIL.n179 0.155672
R317 VTAIL.n222 VTAIL.n221 0.155672
R318 VTAIL.n222 VTAIL.n175 0.155672
R319 VTAIL.n229 VTAIL.n175 0.155672
R320 VTAIL.n22 VTAIL.n21 0.155672
R321 VTAIL.n22 VTAIL.n13 0.155672
R322 VTAIL.n29 VTAIL.n13 0.155672
R323 VTAIL.n30 VTAIL.n29 0.155672
R324 VTAIL.n30 VTAIL.n9 0.155672
R325 VTAIL.n38 VTAIL.n9 0.155672
R326 VTAIL.n39 VTAIL.n38 0.155672
R327 VTAIL.n39 VTAIL.n5 0.155672
R328 VTAIL.n47 VTAIL.n5 0.155672
R329 VTAIL.n48 VTAIL.n47 0.155672
R330 VTAIL.n48 VTAIL.n1 0.155672
R331 VTAIL.n55 VTAIL.n1 0.155672
R332 VTAIL.n171 VTAIL.n117 0.155672
R333 VTAIL.n164 VTAIL.n117 0.155672
R334 VTAIL.n164 VTAIL.n163 0.155672
R335 VTAIL.n163 VTAIL.n121 0.155672
R336 VTAIL.n155 VTAIL.n121 0.155672
R337 VTAIL.n155 VTAIL.n154 0.155672
R338 VTAIL.n154 VTAIL.n125 0.155672
R339 VTAIL.n147 VTAIL.n125 0.155672
R340 VTAIL.n147 VTAIL.n146 0.155672
R341 VTAIL.n146 VTAIL.n130 0.155672
R342 VTAIL.n139 VTAIL.n130 0.155672
R343 VTAIL.n139 VTAIL.n138 0.155672
R344 VTAIL.n113 VTAIL.n59 0.155672
R345 VTAIL.n106 VTAIL.n59 0.155672
R346 VTAIL.n106 VTAIL.n105 0.155672
R347 VTAIL.n105 VTAIL.n63 0.155672
R348 VTAIL.n97 VTAIL.n63 0.155672
R349 VTAIL.n97 VTAIL.n96 0.155672
R350 VTAIL.n96 VTAIL.n67 0.155672
R351 VTAIL.n89 VTAIL.n67 0.155672
R352 VTAIL.n89 VTAIL.n88 0.155672
R353 VTAIL.n88 VTAIL.n72 0.155672
R354 VTAIL.n81 VTAIL.n72 0.155672
R355 VTAIL.n81 VTAIL.n80 0.155672
R356 VDD1.n52 VDD1.n0 289.615
R357 VDD1.n109 VDD1.n57 289.615
R358 VDD1.n53 VDD1.n52 185
R359 VDD1.n51 VDD1.n50 185
R360 VDD1.n4 VDD1.n3 185
R361 VDD1.n45 VDD1.n44 185
R362 VDD1.n43 VDD1.n42 185
R363 VDD1.n41 VDD1.n7 185
R364 VDD1.n11 VDD1.n8 185
R365 VDD1.n36 VDD1.n35 185
R366 VDD1.n34 VDD1.n33 185
R367 VDD1.n13 VDD1.n12 185
R368 VDD1.n28 VDD1.n27 185
R369 VDD1.n26 VDD1.n25 185
R370 VDD1.n17 VDD1.n16 185
R371 VDD1.n20 VDD1.n19 185
R372 VDD1.n76 VDD1.n75 185
R373 VDD1.n73 VDD1.n72 185
R374 VDD1.n82 VDD1.n81 185
R375 VDD1.n84 VDD1.n83 185
R376 VDD1.n69 VDD1.n68 185
R377 VDD1.n90 VDD1.n89 185
R378 VDD1.n93 VDD1.n92 185
R379 VDD1.n91 VDD1.n65 185
R380 VDD1.n98 VDD1.n64 185
R381 VDD1.n100 VDD1.n99 185
R382 VDD1.n102 VDD1.n101 185
R383 VDD1.n61 VDD1.n60 185
R384 VDD1.n108 VDD1.n107 185
R385 VDD1.n110 VDD1.n109 185
R386 VDD1.t1 VDD1.n18 149.524
R387 VDD1.t0 VDD1.n74 149.524
R388 VDD1.n52 VDD1.n51 104.615
R389 VDD1.n51 VDD1.n3 104.615
R390 VDD1.n44 VDD1.n3 104.615
R391 VDD1.n44 VDD1.n43 104.615
R392 VDD1.n43 VDD1.n7 104.615
R393 VDD1.n11 VDD1.n7 104.615
R394 VDD1.n35 VDD1.n11 104.615
R395 VDD1.n35 VDD1.n34 104.615
R396 VDD1.n34 VDD1.n12 104.615
R397 VDD1.n27 VDD1.n12 104.615
R398 VDD1.n27 VDD1.n26 104.615
R399 VDD1.n26 VDD1.n16 104.615
R400 VDD1.n19 VDD1.n16 104.615
R401 VDD1.n75 VDD1.n72 104.615
R402 VDD1.n82 VDD1.n72 104.615
R403 VDD1.n83 VDD1.n82 104.615
R404 VDD1.n83 VDD1.n68 104.615
R405 VDD1.n90 VDD1.n68 104.615
R406 VDD1.n92 VDD1.n90 104.615
R407 VDD1.n92 VDD1.n91 104.615
R408 VDD1.n91 VDD1.n64 104.615
R409 VDD1.n100 VDD1.n64 104.615
R410 VDD1.n101 VDD1.n100 104.615
R411 VDD1.n101 VDD1.n60 104.615
R412 VDD1.n108 VDD1.n60 104.615
R413 VDD1.n109 VDD1.n108 104.615
R414 VDD1 VDD1.n113 84.7531
R415 VDD1.n19 VDD1.t1 52.3082
R416 VDD1.n75 VDD1.t0 52.3082
R417 VDD1 VDD1.n56 49.5408
R418 VDD1.n42 VDD1.n41 13.1884
R419 VDD1.n99 VDD1.n98 13.1884
R420 VDD1.n45 VDD1.n6 12.8005
R421 VDD1.n40 VDD1.n8 12.8005
R422 VDD1.n97 VDD1.n65 12.8005
R423 VDD1.n102 VDD1.n63 12.8005
R424 VDD1.n46 VDD1.n4 12.0247
R425 VDD1.n37 VDD1.n36 12.0247
R426 VDD1.n94 VDD1.n93 12.0247
R427 VDD1.n103 VDD1.n61 12.0247
R428 VDD1.n50 VDD1.n49 11.249
R429 VDD1.n33 VDD1.n10 11.249
R430 VDD1.n89 VDD1.n67 11.249
R431 VDD1.n107 VDD1.n106 11.249
R432 VDD1.n53 VDD1.n2 10.4732
R433 VDD1.n32 VDD1.n13 10.4732
R434 VDD1.n88 VDD1.n69 10.4732
R435 VDD1.n110 VDD1.n59 10.4732
R436 VDD1.n20 VDD1.n18 10.2747
R437 VDD1.n76 VDD1.n74 10.2747
R438 VDD1.n54 VDD1.n0 9.69747
R439 VDD1.n29 VDD1.n28 9.69747
R440 VDD1.n85 VDD1.n84 9.69747
R441 VDD1.n111 VDD1.n57 9.69747
R442 VDD1.n56 VDD1.n55 9.45567
R443 VDD1.n113 VDD1.n112 9.45567
R444 VDD1.n22 VDD1.n21 9.3005
R445 VDD1.n24 VDD1.n23 9.3005
R446 VDD1.n15 VDD1.n14 9.3005
R447 VDD1.n30 VDD1.n29 9.3005
R448 VDD1.n32 VDD1.n31 9.3005
R449 VDD1.n10 VDD1.n9 9.3005
R450 VDD1.n38 VDD1.n37 9.3005
R451 VDD1.n40 VDD1.n39 9.3005
R452 VDD1.n55 VDD1.n54 9.3005
R453 VDD1.n2 VDD1.n1 9.3005
R454 VDD1.n49 VDD1.n48 9.3005
R455 VDD1.n47 VDD1.n46 9.3005
R456 VDD1.n6 VDD1.n5 9.3005
R457 VDD1.n112 VDD1.n111 9.3005
R458 VDD1.n59 VDD1.n58 9.3005
R459 VDD1.n106 VDD1.n105 9.3005
R460 VDD1.n104 VDD1.n103 9.3005
R461 VDD1.n63 VDD1.n62 9.3005
R462 VDD1.n78 VDD1.n77 9.3005
R463 VDD1.n80 VDD1.n79 9.3005
R464 VDD1.n71 VDD1.n70 9.3005
R465 VDD1.n86 VDD1.n85 9.3005
R466 VDD1.n88 VDD1.n87 9.3005
R467 VDD1.n67 VDD1.n66 9.3005
R468 VDD1.n95 VDD1.n94 9.3005
R469 VDD1.n97 VDD1.n96 9.3005
R470 VDD1.n25 VDD1.n15 8.92171
R471 VDD1.n81 VDD1.n71 8.92171
R472 VDD1.n24 VDD1.n17 8.14595
R473 VDD1.n80 VDD1.n73 8.14595
R474 VDD1.n21 VDD1.n20 7.3702
R475 VDD1.n77 VDD1.n76 7.3702
R476 VDD1.n21 VDD1.n17 5.81868
R477 VDD1.n77 VDD1.n73 5.81868
R478 VDD1.n25 VDD1.n24 5.04292
R479 VDD1.n81 VDD1.n80 5.04292
R480 VDD1.n56 VDD1.n0 4.26717
R481 VDD1.n28 VDD1.n15 4.26717
R482 VDD1.n84 VDD1.n71 4.26717
R483 VDD1.n113 VDD1.n57 4.26717
R484 VDD1.n54 VDD1.n53 3.49141
R485 VDD1.n29 VDD1.n13 3.49141
R486 VDD1.n85 VDD1.n69 3.49141
R487 VDD1.n111 VDD1.n110 3.49141
R488 VDD1.n22 VDD1.n18 2.84303
R489 VDD1.n78 VDD1.n74 2.84303
R490 VDD1.n50 VDD1.n2 2.71565
R491 VDD1.n33 VDD1.n32 2.71565
R492 VDD1.n89 VDD1.n88 2.71565
R493 VDD1.n107 VDD1.n59 2.71565
R494 VDD1.n49 VDD1.n4 1.93989
R495 VDD1.n36 VDD1.n10 1.93989
R496 VDD1.n93 VDD1.n67 1.93989
R497 VDD1.n106 VDD1.n61 1.93989
R498 VDD1.n46 VDD1.n45 1.16414
R499 VDD1.n37 VDD1.n8 1.16414
R500 VDD1.n94 VDD1.n65 1.16414
R501 VDD1.n103 VDD1.n102 1.16414
R502 VDD1.n42 VDD1.n6 0.388379
R503 VDD1.n41 VDD1.n40 0.388379
R504 VDD1.n98 VDD1.n97 0.388379
R505 VDD1.n99 VDD1.n63 0.388379
R506 VDD1.n55 VDD1.n1 0.155672
R507 VDD1.n48 VDD1.n1 0.155672
R508 VDD1.n48 VDD1.n47 0.155672
R509 VDD1.n47 VDD1.n5 0.155672
R510 VDD1.n39 VDD1.n5 0.155672
R511 VDD1.n39 VDD1.n38 0.155672
R512 VDD1.n38 VDD1.n9 0.155672
R513 VDD1.n31 VDD1.n9 0.155672
R514 VDD1.n31 VDD1.n30 0.155672
R515 VDD1.n30 VDD1.n14 0.155672
R516 VDD1.n23 VDD1.n14 0.155672
R517 VDD1.n23 VDD1.n22 0.155672
R518 VDD1.n79 VDD1.n78 0.155672
R519 VDD1.n79 VDD1.n70 0.155672
R520 VDD1.n86 VDD1.n70 0.155672
R521 VDD1.n87 VDD1.n86 0.155672
R522 VDD1.n87 VDD1.n66 0.155672
R523 VDD1.n95 VDD1.n66 0.155672
R524 VDD1.n96 VDD1.n95 0.155672
R525 VDD1.n96 VDD1.n62 0.155672
R526 VDD1.n104 VDD1.n62 0.155672
R527 VDD1.n105 VDD1.n104 0.155672
R528 VDD1.n105 VDD1.n58 0.155672
R529 VDD1.n112 VDD1.n58 0.155672
R530 B.n385 B.n384 585
R531 B.n385 B.n30 585
R532 B.n388 B.n387 585
R533 B.n389 B.n77 585
R534 B.n391 B.n390 585
R535 B.n393 B.n76 585
R536 B.n396 B.n395 585
R537 B.n397 B.n75 585
R538 B.n399 B.n398 585
R539 B.n401 B.n74 585
R540 B.n404 B.n403 585
R541 B.n405 B.n73 585
R542 B.n407 B.n406 585
R543 B.n409 B.n72 585
R544 B.n412 B.n411 585
R545 B.n413 B.n71 585
R546 B.n415 B.n414 585
R547 B.n417 B.n70 585
R548 B.n420 B.n419 585
R549 B.n421 B.n69 585
R550 B.n423 B.n422 585
R551 B.n425 B.n68 585
R552 B.n428 B.n427 585
R553 B.n429 B.n67 585
R554 B.n431 B.n430 585
R555 B.n433 B.n66 585
R556 B.n436 B.n435 585
R557 B.n437 B.n65 585
R558 B.n439 B.n438 585
R559 B.n441 B.n64 585
R560 B.n444 B.n443 585
R561 B.n445 B.n63 585
R562 B.n447 B.n446 585
R563 B.n449 B.n62 585
R564 B.n452 B.n451 585
R565 B.n453 B.n61 585
R566 B.n455 B.n454 585
R567 B.n457 B.n60 585
R568 B.n460 B.n459 585
R569 B.n462 B.n57 585
R570 B.n464 B.n463 585
R571 B.n466 B.n56 585
R572 B.n469 B.n468 585
R573 B.n470 B.n55 585
R574 B.n472 B.n471 585
R575 B.n474 B.n54 585
R576 B.n476 B.n475 585
R577 B.n478 B.n477 585
R578 B.n481 B.n480 585
R579 B.n482 B.n49 585
R580 B.n484 B.n483 585
R581 B.n486 B.n48 585
R582 B.n489 B.n488 585
R583 B.n490 B.n47 585
R584 B.n492 B.n491 585
R585 B.n494 B.n46 585
R586 B.n497 B.n496 585
R587 B.n498 B.n45 585
R588 B.n500 B.n499 585
R589 B.n502 B.n44 585
R590 B.n505 B.n504 585
R591 B.n506 B.n43 585
R592 B.n508 B.n507 585
R593 B.n510 B.n42 585
R594 B.n513 B.n512 585
R595 B.n514 B.n41 585
R596 B.n516 B.n515 585
R597 B.n518 B.n40 585
R598 B.n521 B.n520 585
R599 B.n522 B.n39 585
R600 B.n524 B.n523 585
R601 B.n526 B.n38 585
R602 B.n529 B.n528 585
R603 B.n530 B.n37 585
R604 B.n532 B.n531 585
R605 B.n534 B.n36 585
R606 B.n537 B.n536 585
R607 B.n538 B.n35 585
R608 B.n540 B.n539 585
R609 B.n542 B.n34 585
R610 B.n545 B.n544 585
R611 B.n546 B.n33 585
R612 B.n548 B.n547 585
R613 B.n550 B.n32 585
R614 B.n553 B.n552 585
R615 B.n554 B.n31 585
R616 B.n383 B.n29 585
R617 B.n557 B.n29 585
R618 B.n382 B.n28 585
R619 B.n558 B.n28 585
R620 B.n381 B.n27 585
R621 B.n559 B.n27 585
R622 B.n380 B.n379 585
R623 B.n379 B.n23 585
R624 B.n378 B.n22 585
R625 B.n565 B.n22 585
R626 B.n377 B.n21 585
R627 B.n566 B.n21 585
R628 B.n376 B.n20 585
R629 B.n567 B.n20 585
R630 B.n375 B.n374 585
R631 B.n374 B.n16 585
R632 B.n373 B.n15 585
R633 B.n573 B.n15 585
R634 B.n372 B.n14 585
R635 B.n574 B.n14 585
R636 B.n371 B.n13 585
R637 B.n575 B.n13 585
R638 B.n370 B.n369 585
R639 B.n369 B.n12 585
R640 B.n368 B.n367 585
R641 B.n368 B.n8 585
R642 B.n366 B.n7 585
R643 B.n582 B.n7 585
R644 B.n365 B.n6 585
R645 B.n583 B.n6 585
R646 B.n364 B.n5 585
R647 B.n584 B.n5 585
R648 B.n363 B.n362 585
R649 B.n362 B.n4 585
R650 B.n361 B.n78 585
R651 B.n361 B.n360 585
R652 B.n350 B.n79 585
R653 B.n353 B.n79 585
R654 B.n352 B.n351 585
R655 B.n354 B.n352 585
R656 B.n349 B.n84 585
R657 B.n84 B.n83 585
R658 B.n348 B.n347 585
R659 B.n347 B.n346 585
R660 B.n86 B.n85 585
R661 B.n87 B.n86 585
R662 B.n339 B.n338 585
R663 B.n340 B.n339 585
R664 B.n337 B.n92 585
R665 B.n92 B.n91 585
R666 B.n336 B.n335 585
R667 B.n335 B.n334 585
R668 B.n94 B.n93 585
R669 B.n95 B.n94 585
R670 B.n327 B.n326 585
R671 B.n328 B.n327 585
R672 B.n325 B.n100 585
R673 B.n100 B.n99 585
R674 B.n324 B.n323 585
R675 B.n323 B.n322 585
R676 B.n319 B.n104 585
R677 B.n318 B.n317 585
R678 B.n315 B.n105 585
R679 B.n315 B.n103 585
R680 B.n314 B.n313 585
R681 B.n312 B.n311 585
R682 B.n310 B.n107 585
R683 B.n308 B.n307 585
R684 B.n306 B.n108 585
R685 B.n305 B.n304 585
R686 B.n302 B.n109 585
R687 B.n300 B.n299 585
R688 B.n298 B.n110 585
R689 B.n297 B.n296 585
R690 B.n294 B.n111 585
R691 B.n292 B.n291 585
R692 B.n290 B.n112 585
R693 B.n289 B.n288 585
R694 B.n286 B.n113 585
R695 B.n284 B.n283 585
R696 B.n282 B.n114 585
R697 B.n281 B.n280 585
R698 B.n278 B.n115 585
R699 B.n276 B.n275 585
R700 B.n274 B.n116 585
R701 B.n273 B.n272 585
R702 B.n270 B.n117 585
R703 B.n268 B.n267 585
R704 B.n266 B.n118 585
R705 B.n265 B.n264 585
R706 B.n262 B.n119 585
R707 B.n260 B.n259 585
R708 B.n258 B.n120 585
R709 B.n257 B.n256 585
R710 B.n254 B.n121 585
R711 B.n252 B.n251 585
R712 B.n250 B.n122 585
R713 B.n249 B.n248 585
R714 B.n246 B.n123 585
R715 B.n244 B.n243 585
R716 B.n242 B.n124 585
R717 B.n241 B.n240 585
R718 B.n238 B.n128 585
R719 B.n236 B.n235 585
R720 B.n234 B.n129 585
R721 B.n233 B.n232 585
R722 B.n230 B.n130 585
R723 B.n228 B.n227 585
R724 B.n225 B.n131 585
R725 B.n224 B.n223 585
R726 B.n221 B.n134 585
R727 B.n219 B.n218 585
R728 B.n217 B.n135 585
R729 B.n216 B.n215 585
R730 B.n213 B.n136 585
R731 B.n211 B.n210 585
R732 B.n209 B.n137 585
R733 B.n208 B.n207 585
R734 B.n205 B.n138 585
R735 B.n203 B.n202 585
R736 B.n201 B.n139 585
R737 B.n200 B.n199 585
R738 B.n197 B.n140 585
R739 B.n195 B.n194 585
R740 B.n193 B.n141 585
R741 B.n192 B.n191 585
R742 B.n189 B.n142 585
R743 B.n187 B.n186 585
R744 B.n185 B.n143 585
R745 B.n184 B.n183 585
R746 B.n181 B.n144 585
R747 B.n179 B.n178 585
R748 B.n177 B.n145 585
R749 B.n176 B.n175 585
R750 B.n173 B.n146 585
R751 B.n171 B.n170 585
R752 B.n169 B.n147 585
R753 B.n168 B.n167 585
R754 B.n165 B.n148 585
R755 B.n163 B.n162 585
R756 B.n161 B.n149 585
R757 B.n160 B.n159 585
R758 B.n157 B.n150 585
R759 B.n155 B.n154 585
R760 B.n153 B.n152 585
R761 B.n102 B.n101 585
R762 B.n321 B.n320 585
R763 B.n322 B.n321 585
R764 B.n98 B.n97 585
R765 B.n99 B.n98 585
R766 B.n330 B.n329 585
R767 B.n329 B.n328 585
R768 B.n331 B.n96 585
R769 B.n96 B.n95 585
R770 B.n333 B.n332 585
R771 B.n334 B.n333 585
R772 B.n90 B.n89 585
R773 B.n91 B.n90 585
R774 B.n342 B.n341 585
R775 B.n341 B.n340 585
R776 B.n343 B.n88 585
R777 B.n88 B.n87 585
R778 B.n345 B.n344 585
R779 B.n346 B.n345 585
R780 B.n82 B.n81 585
R781 B.n83 B.n82 585
R782 B.n356 B.n355 585
R783 B.n355 B.n354 585
R784 B.n357 B.n80 585
R785 B.n353 B.n80 585
R786 B.n359 B.n358 585
R787 B.n360 B.n359 585
R788 B.n3 B.n0 585
R789 B.n4 B.n3 585
R790 B.n581 B.n1 585
R791 B.n582 B.n581 585
R792 B.n580 B.n579 585
R793 B.n580 B.n8 585
R794 B.n578 B.n9 585
R795 B.n12 B.n9 585
R796 B.n577 B.n576 585
R797 B.n576 B.n575 585
R798 B.n11 B.n10 585
R799 B.n574 B.n11 585
R800 B.n572 B.n571 585
R801 B.n573 B.n572 585
R802 B.n570 B.n17 585
R803 B.n17 B.n16 585
R804 B.n569 B.n568 585
R805 B.n568 B.n567 585
R806 B.n19 B.n18 585
R807 B.n566 B.n19 585
R808 B.n564 B.n563 585
R809 B.n565 B.n564 585
R810 B.n562 B.n24 585
R811 B.n24 B.n23 585
R812 B.n561 B.n560 585
R813 B.n560 B.n559 585
R814 B.n26 B.n25 585
R815 B.n558 B.n26 585
R816 B.n556 B.n555 585
R817 B.n557 B.n556 585
R818 B.n585 B.n584 585
R819 B.n583 B.n2 585
R820 B.n50 B.t2 550.972
R821 B.n58 B.t13 550.972
R822 B.n132 B.t10 550.972
R823 B.n125 B.t6 550.972
R824 B.n556 B.n31 506.916
R825 B.n385 B.n29 506.916
R826 B.n323 B.n102 506.916
R827 B.n321 B.n104 506.916
R828 B.n58 B.t14 280.498
R829 B.n132 B.t12 280.498
R830 B.n50 B.t4 280.498
R831 B.n125 B.t9 280.498
R832 B.n59 B.t15 259.748
R833 B.n133 B.t11 259.748
R834 B.n51 B.t5 259.748
R835 B.n126 B.t8 259.748
R836 B.n386 B.n30 256.663
R837 B.n392 B.n30 256.663
R838 B.n394 B.n30 256.663
R839 B.n400 B.n30 256.663
R840 B.n402 B.n30 256.663
R841 B.n408 B.n30 256.663
R842 B.n410 B.n30 256.663
R843 B.n416 B.n30 256.663
R844 B.n418 B.n30 256.663
R845 B.n424 B.n30 256.663
R846 B.n426 B.n30 256.663
R847 B.n432 B.n30 256.663
R848 B.n434 B.n30 256.663
R849 B.n440 B.n30 256.663
R850 B.n442 B.n30 256.663
R851 B.n448 B.n30 256.663
R852 B.n450 B.n30 256.663
R853 B.n456 B.n30 256.663
R854 B.n458 B.n30 256.663
R855 B.n465 B.n30 256.663
R856 B.n467 B.n30 256.663
R857 B.n473 B.n30 256.663
R858 B.n53 B.n30 256.663
R859 B.n479 B.n30 256.663
R860 B.n485 B.n30 256.663
R861 B.n487 B.n30 256.663
R862 B.n493 B.n30 256.663
R863 B.n495 B.n30 256.663
R864 B.n501 B.n30 256.663
R865 B.n503 B.n30 256.663
R866 B.n509 B.n30 256.663
R867 B.n511 B.n30 256.663
R868 B.n517 B.n30 256.663
R869 B.n519 B.n30 256.663
R870 B.n525 B.n30 256.663
R871 B.n527 B.n30 256.663
R872 B.n533 B.n30 256.663
R873 B.n535 B.n30 256.663
R874 B.n541 B.n30 256.663
R875 B.n543 B.n30 256.663
R876 B.n549 B.n30 256.663
R877 B.n551 B.n30 256.663
R878 B.n316 B.n103 256.663
R879 B.n106 B.n103 256.663
R880 B.n309 B.n103 256.663
R881 B.n303 B.n103 256.663
R882 B.n301 B.n103 256.663
R883 B.n295 B.n103 256.663
R884 B.n293 B.n103 256.663
R885 B.n287 B.n103 256.663
R886 B.n285 B.n103 256.663
R887 B.n279 B.n103 256.663
R888 B.n277 B.n103 256.663
R889 B.n271 B.n103 256.663
R890 B.n269 B.n103 256.663
R891 B.n263 B.n103 256.663
R892 B.n261 B.n103 256.663
R893 B.n255 B.n103 256.663
R894 B.n253 B.n103 256.663
R895 B.n247 B.n103 256.663
R896 B.n245 B.n103 256.663
R897 B.n239 B.n103 256.663
R898 B.n237 B.n103 256.663
R899 B.n231 B.n103 256.663
R900 B.n229 B.n103 256.663
R901 B.n222 B.n103 256.663
R902 B.n220 B.n103 256.663
R903 B.n214 B.n103 256.663
R904 B.n212 B.n103 256.663
R905 B.n206 B.n103 256.663
R906 B.n204 B.n103 256.663
R907 B.n198 B.n103 256.663
R908 B.n196 B.n103 256.663
R909 B.n190 B.n103 256.663
R910 B.n188 B.n103 256.663
R911 B.n182 B.n103 256.663
R912 B.n180 B.n103 256.663
R913 B.n174 B.n103 256.663
R914 B.n172 B.n103 256.663
R915 B.n166 B.n103 256.663
R916 B.n164 B.n103 256.663
R917 B.n158 B.n103 256.663
R918 B.n156 B.n103 256.663
R919 B.n151 B.n103 256.663
R920 B.n587 B.n586 256.663
R921 B.n552 B.n550 163.367
R922 B.n548 B.n33 163.367
R923 B.n544 B.n542 163.367
R924 B.n540 B.n35 163.367
R925 B.n536 B.n534 163.367
R926 B.n532 B.n37 163.367
R927 B.n528 B.n526 163.367
R928 B.n524 B.n39 163.367
R929 B.n520 B.n518 163.367
R930 B.n516 B.n41 163.367
R931 B.n512 B.n510 163.367
R932 B.n508 B.n43 163.367
R933 B.n504 B.n502 163.367
R934 B.n500 B.n45 163.367
R935 B.n496 B.n494 163.367
R936 B.n492 B.n47 163.367
R937 B.n488 B.n486 163.367
R938 B.n484 B.n49 163.367
R939 B.n480 B.n478 163.367
R940 B.n475 B.n474 163.367
R941 B.n472 B.n55 163.367
R942 B.n468 B.n466 163.367
R943 B.n464 B.n57 163.367
R944 B.n459 B.n457 163.367
R945 B.n455 B.n61 163.367
R946 B.n451 B.n449 163.367
R947 B.n447 B.n63 163.367
R948 B.n443 B.n441 163.367
R949 B.n439 B.n65 163.367
R950 B.n435 B.n433 163.367
R951 B.n431 B.n67 163.367
R952 B.n427 B.n425 163.367
R953 B.n423 B.n69 163.367
R954 B.n419 B.n417 163.367
R955 B.n415 B.n71 163.367
R956 B.n411 B.n409 163.367
R957 B.n407 B.n73 163.367
R958 B.n403 B.n401 163.367
R959 B.n399 B.n75 163.367
R960 B.n395 B.n393 163.367
R961 B.n391 B.n77 163.367
R962 B.n387 B.n385 163.367
R963 B.n323 B.n100 163.367
R964 B.n327 B.n100 163.367
R965 B.n327 B.n94 163.367
R966 B.n335 B.n94 163.367
R967 B.n335 B.n92 163.367
R968 B.n339 B.n92 163.367
R969 B.n339 B.n86 163.367
R970 B.n347 B.n86 163.367
R971 B.n347 B.n84 163.367
R972 B.n352 B.n84 163.367
R973 B.n352 B.n79 163.367
R974 B.n361 B.n79 163.367
R975 B.n362 B.n361 163.367
R976 B.n362 B.n5 163.367
R977 B.n6 B.n5 163.367
R978 B.n7 B.n6 163.367
R979 B.n368 B.n7 163.367
R980 B.n369 B.n368 163.367
R981 B.n369 B.n13 163.367
R982 B.n14 B.n13 163.367
R983 B.n15 B.n14 163.367
R984 B.n374 B.n15 163.367
R985 B.n374 B.n20 163.367
R986 B.n21 B.n20 163.367
R987 B.n22 B.n21 163.367
R988 B.n379 B.n22 163.367
R989 B.n379 B.n27 163.367
R990 B.n28 B.n27 163.367
R991 B.n29 B.n28 163.367
R992 B.n317 B.n315 163.367
R993 B.n315 B.n314 163.367
R994 B.n311 B.n310 163.367
R995 B.n308 B.n108 163.367
R996 B.n304 B.n302 163.367
R997 B.n300 B.n110 163.367
R998 B.n296 B.n294 163.367
R999 B.n292 B.n112 163.367
R1000 B.n288 B.n286 163.367
R1001 B.n284 B.n114 163.367
R1002 B.n280 B.n278 163.367
R1003 B.n276 B.n116 163.367
R1004 B.n272 B.n270 163.367
R1005 B.n268 B.n118 163.367
R1006 B.n264 B.n262 163.367
R1007 B.n260 B.n120 163.367
R1008 B.n256 B.n254 163.367
R1009 B.n252 B.n122 163.367
R1010 B.n248 B.n246 163.367
R1011 B.n244 B.n124 163.367
R1012 B.n240 B.n238 163.367
R1013 B.n236 B.n129 163.367
R1014 B.n232 B.n230 163.367
R1015 B.n228 B.n131 163.367
R1016 B.n223 B.n221 163.367
R1017 B.n219 B.n135 163.367
R1018 B.n215 B.n213 163.367
R1019 B.n211 B.n137 163.367
R1020 B.n207 B.n205 163.367
R1021 B.n203 B.n139 163.367
R1022 B.n199 B.n197 163.367
R1023 B.n195 B.n141 163.367
R1024 B.n191 B.n189 163.367
R1025 B.n187 B.n143 163.367
R1026 B.n183 B.n181 163.367
R1027 B.n179 B.n145 163.367
R1028 B.n175 B.n173 163.367
R1029 B.n171 B.n147 163.367
R1030 B.n167 B.n165 163.367
R1031 B.n163 B.n149 163.367
R1032 B.n159 B.n157 163.367
R1033 B.n155 B.n152 163.367
R1034 B.n321 B.n98 163.367
R1035 B.n329 B.n98 163.367
R1036 B.n329 B.n96 163.367
R1037 B.n333 B.n96 163.367
R1038 B.n333 B.n90 163.367
R1039 B.n341 B.n90 163.367
R1040 B.n341 B.n88 163.367
R1041 B.n345 B.n88 163.367
R1042 B.n345 B.n82 163.367
R1043 B.n355 B.n82 163.367
R1044 B.n355 B.n80 163.367
R1045 B.n359 B.n80 163.367
R1046 B.n359 B.n3 163.367
R1047 B.n585 B.n3 163.367
R1048 B.n581 B.n2 163.367
R1049 B.n581 B.n580 163.367
R1050 B.n580 B.n9 163.367
R1051 B.n576 B.n9 163.367
R1052 B.n576 B.n11 163.367
R1053 B.n572 B.n11 163.367
R1054 B.n572 B.n17 163.367
R1055 B.n568 B.n17 163.367
R1056 B.n568 B.n19 163.367
R1057 B.n564 B.n19 163.367
R1058 B.n564 B.n24 163.367
R1059 B.n560 B.n24 163.367
R1060 B.n560 B.n26 163.367
R1061 B.n556 B.n26 163.367
R1062 B.n322 B.n103 80.4631
R1063 B.n557 B.n30 80.4631
R1064 B.n551 B.n31 71.676
R1065 B.n550 B.n549 71.676
R1066 B.n543 B.n33 71.676
R1067 B.n542 B.n541 71.676
R1068 B.n535 B.n35 71.676
R1069 B.n534 B.n533 71.676
R1070 B.n527 B.n37 71.676
R1071 B.n526 B.n525 71.676
R1072 B.n519 B.n39 71.676
R1073 B.n518 B.n517 71.676
R1074 B.n511 B.n41 71.676
R1075 B.n510 B.n509 71.676
R1076 B.n503 B.n43 71.676
R1077 B.n502 B.n501 71.676
R1078 B.n495 B.n45 71.676
R1079 B.n494 B.n493 71.676
R1080 B.n487 B.n47 71.676
R1081 B.n486 B.n485 71.676
R1082 B.n479 B.n49 71.676
R1083 B.n478 B.n53 71.676
R1084 B.n474 B.n473 71.676
R1085 B.n467 B.n55 71.676
R1086 B.n466 B.n465 71.676
R1087 B.n458 B.n57 71.676
R1088 B.n457 B.n456 71.676
R1089 B.n450 B.n61 71.676
R1090 B.n449 B.n448 71.676
R1091 B.n442 B.n63 71.676
R1092 B.n441 B.n440 71.676
R1093 B.n434 B.n65 71.676
R1094 B.n433 B.n432 71.676
R1095 B.n426 B.n67 71.676
R1096 B.n425 B.n424 71.676
R1097 B.n418 B.n69 71.676
R1098 B.n417 B.n416 71.676
R1099 B.n410 B.n71 71.676
R1100 B.n409 B.n408 71.676
R1101 B.n402 B.n73 71.676
R1102 B.n401 B.n400 71.676
R1103 B.n394 B.n75 71.676
R1104 B.n393 B.n392 71.676
R1105 B.n386 B.n77 71.676
R1106 B.n387 B.n386 71.676
R1107 B.n392 B.n391 71.676
R1108 B.n395 B.n394 71.676
R1109 B.n400 B.n399 71.676
R1110 B.n403 B.n402 71.676
R1111 B.n408 B.n407 71.676
R1112 B.n411 B.n410 71.676
R1113 B.n416 B.n415 71.676
R1114 B.n419 B.n418 71.676
R1115 B.n424 B.n423 71.676
R1116 B.n427 B.n426 71.676
R1117 B.n432 B.n431 71.676
R1118 B.n435 B.n434 71.676
R1119 B.n440 B.n439 71.676
R1120 B.n443 B.n442 71.676
R1121 B.n448 B.n447 71.676
R1122 B.n451 B.n450 71.676
R1123 B.n456 B.n455 71.676
R1124 B.n459 B.n458 71.676
R1125 B.n465 B.n464 71.676
R1126 B.n468 B.n467 71.676
R1127 B.n473 B.n472 71.676
R1128 B.n475 B.n53 71.676
R1129 B.n480 B.n479 71.676
R1130 B.n485 B.n484 71.676
R1131 B.n488 B.n487 71.676
R1132 B.n493 B.n492 71.676
R1133 B.n496 B.n495 71.676
R1134 B.n501 B.n500 71.676
R1135 B.n504 B.n503 71.676
R1136 B.n509 B.n508 71.676
R1137 B.n512 B.n511 71.676
R1138 B.n517 B.n516 71.676
R1139 B.n520 B.n519 71.676
R1140 B.n525 B.n524 71.676
R1141 B.n528 B.n527 71.676
R1142 B.n533 B.n532 71.676
R1143 B.n536 B.n535 71.676
R1144 B.n541 B.n540 71.676
R1145 B.n544 B.n543 71.676
R1146 B.n549 B.n548 71.676
R1147 B.n552 B.n551 71.676
R1148 B.n316 B.n104 71.676
R1149 B.n314 B.n106 71.676
R1150 B.n310 B.n309 71.676
R1151 B.n303 B.n108 71.676
R1152 B.n302 B.n301 71.676
R1153 B.n295 B.n110 71.676
R1154 B.n294 B.n293 71.676
R1155 B.n287 B.n112 71.676
R1156 B.n286 B.n285 71.676
R1157 B.n279 B.n114 71.676
R1158 B.n278 B.n277 71.676
R1159 B.n271 B.n116 71.676
R1160 B.n270 B.n269 71.676
R1161 B.n263 B.n118 71.676
R1162 B.n262 B.n261 71.676
R1163 B.n255 B.n120 71.676
R1164 B.n254 B.n253 71.676
R1165 B.n247 B.n122 71.676
R1166 B.n246 B.n245 71.676
R1167 B.n239 B.n124 71.676
R1168 B.n238 B.n237 71.676
R1169 B.n231 B.n129 71.676
R1170 B.n230 B.n229 71.676
R1171 B.n222 B.n131 71.676
R1172 B.n221 B.n220 71.676
R1173 B.n214 B.n135 71.676
R1174 B.n213 B.n212 71.676
R1175 B.n206 B.n137 71.676
R1176 B.n205 B.n204 71.676
R1177 B.n198 B.n139 71.676
R1178 B.n197 B.n196 71.676
R1179 B.n190 B.n141 71.676
R1180 B.n189 B.n188 71.676
R1181 B.n182 B.n143 71.676
R1182 B.n181 B.n180 71.676
R1183 B.n174 B.n145 71.676
R1184 B.n173 B.n172 71.676
R1185 B.n166 B.n147 71.676
R1186 B.n165 B.n164 71.676
R1187 B.n158 B.n149 71.676
R1188 B.n157 B.n156 71.676
R1189 B.n152 B.n151 71.676
R1190 B.n317 B.n316 71.676
R1191 B.n311 B.n106 71.676
R1192 B.n309 B.n308 71.676
R1193 B.n304 B.n303 71.676
R1194 B.n301 B.n300 71.676
R1195 B.n296 B.n295 71.676
R1196 B.n293 B.n292 71.676
R1197 B.n288 B.n287 71.676
R1198 B.n285 B.n284 71.676
R1199 B.n280 B.n279 71.676
R1200 B.n277 B.n276 71.676
R1201 B.n272 B.n271 71.676
R1202 B.n269 B.n268 71.676
R1203 B.n264 B.n263 71.676
R1204 B.n261 B.n260 71.676
R1205 B.n256 B.n255 71.676
R1206 B.n253 B.n252 71.676
R1207 B.n248 B.n247 71.676
R1208 B.n245 B.n244 71.676
R1209 B.n240 B.n239 71.676
R1210 B.n237 B.n236 71.676
R1211 B.n232 B.n231 71.676
R1212 B.n229 B.n228 71.676
R1213 B.n223 B.n222 71.676
R1214 B.n220 B.n219 71.676
R1215 B.n215 B.n214 71.676
R1216 B.n212 B.n211 71.676
R1217 B.n207 B.n206 71.676
R1218 B.n204 B.n203 71.676
R1219 B.n199 B.n198 71.676
R1220 B.n196 B.n195 71.676
R1221 B.n191 B.n190 71.676
R1222 B.n188 B.n187 71.676
R1223 B.n183 B.n182 71.676
R1224 B.n180 B.n179 71.676
R1225 B.n175 B.n174 71.676
R1226 B.n172 B.n171 71.676
R1227 B.n167 B.n166 71.676
R1228 B.n164 B.n163 71.676
R1229 B.n159 B.n158 71.676
R1230 B.n156 B.n155 71.676
R1231 B.n151 B.n102 71.676
R1232 B.n586 B.n585 71.676
R1233 B.n586 B.n2 71.676
R1234 B.n52 B.n51 59.5399
R1235 B.n461 B.n59 59.5399
R1236 B.n226 B.n133 59.5399
R1237 B.n127 B.n126 59.5399
R1238 B.n322 B.n99 46.7651
R1239 B.n328 B.n99 46.7651
R1240 B.n328 B.n95 46.7651
R1241 B.n334 B.n95 46.7651
R1242 B.n340 B.n91 46.7651
R1243 B.n340 B.n87 46.7651
R1244 B.n346 B.n87 46.7651
R1245 B.n346 B.n83 46.7651
R1246 B.n354 B.n83 46.7651
R1247 B.n354 B.n353 46.7651
R1248 B.n360 B.n4 46.7651
R1249 B.n584 B.n4 46.7651
R1250 B.n584 B.n583 46.7651
R1251 B.n583 B.n582 46.7651
R1252 B.n582 B.n8 46.7651
R1253 B.n575 B.n12 46.7651
R1254 B.n575 B.n574 46.7651
R1255 B.n574 B.n573 46.7651
R1256 B.n573 B.n16 46.7651
R1257 B.n567 B.n16 46.7651
R1258 B.n567 B.n566 46.7651
R1259 B.n565 B.n23 46.7651
R1260 B.n559 B.n23 46.7651
R1261 B.n559 B.n558 46.7651
R1262 B.n558 B.n557 46.7651
R1263 B.n334 B.t7 45.3897
R1264 B.t3 B.n565 45.3897
R1265 B.n320 B.n319 32.9371
R1266 B.n324 B.n101 32.9371
R1267 B.n384 B.n383 32.9371
R1268 B.n555 B.n554 32.9371
R1269 B.n360 B.t0 31.6354
R1270 B.t1 B.n8 31.6354
R1271 B.n51 B.n50 20.752
R1272 B.n59 B.n58 20.752
R1273 B.n133 B.n132 20.752
R1274 B.n126 B.n125 20.752
R1275 B B.n587 18.0485
R1276 B.n353 B.t0 15.1302
R1277 B.n12 B.t1 15.1302
R1278 B.n320 B.n97 10.6151
R1279 B.n330 B.n97 10.6151
R1280 B.n331 B.n330 10.6151
R1281 B.n332 B.n331 10.6151
R1282 B.n332 B.n89 10.6151
R1283 B.n342 B.n89 10.6151
R1284 B.n343 B.n342 10.6151
R1285 B.n344 B.n343 10.6151
R1286 B.n344 B.n81 10.6151
R1287 B.n356 B.n81 10.6151
R1288 B.n357 B.n356 10.6151
R1289 B.n358 B.n357 10.6151
R1290 B.n358 B.n0 10.6151
R1291 B.n319 B.n318 10.6151
R1292 B.n318 B.n105 10.6151
R1293 B.n313 B.n105 10.6151
R1294 B.n313 B.n312 10.6151
R1295 B.n312 B.n107 10.6151
R1296 B.n307 B.n107 10.6151
R1297 B.n307 B.n306 10.6151
R1298 B.n306 B.n305 10.6151
R1299 B.n305 B.n109 10.6151
R1300 B.n299 B.n109 10.6151
R1301 B.n299 B.n298 10.6151
R1302 B.n298 B.n297 10.6151
R1303 B.n297 B.n111 10.6151
R1304 B.n291 B.n111 10.6151
R1305 B.n291 B.n290 10.6151
R1306 B.n290 B.n289 10.6151
R1307 B.n289 B.n113 10.6151
R1308 B.n283 B.n113 10.6151
R1309 B.n283 B.n282 10.6151
R1310 B.n282 B.n281 10.6151
R1311 B.n281 B.n115 10.6151
R1312 B.n275 B.n115 10.6151
R1313 B.n275 B.n274 10.6151
R1314 B.n274 B.n273 10.6151
R1315 B.n273 B.n117 10.6151
R1316 B.n267 B.n117 10.6151
R1317 B.n267 B.n266 10.6151
R1318 B.n266 B.n265 10.6151
R1319 B.n265 B.n119 10.6151
R1320 B.n259 B.n119 10.6151
R1321 B.n259 B.n258 10.6151
R1322 B.n258 B.n257 10.6151
R1323 B.n257 B.n121 10.6151
R1324 B.n251 B.n121 10.6151
R1325 B.n251 B.n250 10.6151
R1326 B.n250 B.n249 10.6151
R1327 B.n249 B.n123 10.6151
R1328 B.n243 B.n242 10.6151
R1329 B.n242 B.n241 10.6151
R1330 B.n241 B.n128 10.6151
R1331 B.n235 B.n128 10.6151
R1332 B.n235 B.n234 10.6151
R1333 B.n234 B.n233 10.6151
R1334 B.n233 B.n130 10.6151
R1335 B.n227 B.n130 10.6151
R1336 B.n225 B.n224 10.6151
R1337 B.n224 B.n134 10.6151
R1338 B.n218 B.n134 10.6151
R1339 B.n218 B.n217 10.6151
R1340 B.n217 B.n216 10.6151
R1341 B.n216 B.n136 10.6151
R1342 B.n210 B.n136 10.6151
R1343 B.n210 B.n209 10.6151
R1344 B.n209 B.n208 10.6151
R1345 B.n208 B.n138 10.6151
R1346 B.n202 B.n138 10.6151
R1347 B.n202 B.n201 10.6151
R1348 B.n201 B.n200 10.6151
R1349 B.n200 B.n140 10.6151
R1350 B.n194 B.n140 10.6151
R1351 B.n194 B.n193 10.6151
R1352 B.n193 B.n192 10.6151
R1353 B.n192 B.n142 10.6151
R1354 B.n186 B.n142 10.6151
R1355 B.n186 B.n185 10.6151
R1356 B.n185 B.n184 10.6151
R1357 B.n184 B.n144 10.6151
R1358 B.n178 B.n144 10.6151
R1359 B.n178 B.n177 10.6151
R1360 B.n177 B.n176 10.6151
R1361 B.n176 B.n146 10.6151
R1362 B.n170 B.n146 10.6151
R1363 B.n170 B.n169 10.6151
R1364 B.n169 B.n168 10.6151
R1365 B.n168 B.n148 10.6151
R1366 B.n162 B.n148 10.6151
R1367 B.n162 B.n161 10.6151
R1368 B.n161 B.n160 10.6151
R1369 B.n160 B.n150 10.6151
R1370 B.n154 B.n150 10.6151
R1371 B.n154 B.n153 10.6151
R1372 B.n153 B.n101 10.6151
R1373 B.n325 B.n324 10.6151
R1374 B.n326 B.n325 10.6151
R1375 B.n326 B.n93 10.6151
R1376 B.n336 B.n93 10.6151
R1377 B.n337 B.n336 10.6151
R1378 B.n338 B.n337 10.6151
R1379 B.n338 B.n85 10.6151
R1380 B.n348 B.n85 10.6151
R1381 B.n349 B.n348 10.6151
R1382 B.n351 B.n349 10.6151
R1383 B.n351 B.n350 10.6151
R1384 B.n350 B.n78 10.6151
R1385 B.n363 B.n78 10.6151
R1386 B.n364 B.n363 10.6151
R1387 B.n365 B.n364 10.6151
R1388 B.n366 B.n365 10.6151
R1389 B.n367 B.n366 10.6151
R1390 B.n370 B.n367 10.6151
R1391 B.n371 B.n370 10.6151
R1392 B.n372 B.n371 10.6151
R1393 B.n373 B.n372 10.6151
R1394 B.n375 B.n373 10.6151
R1395 B.n376 B.n375 10.6151
R1396 B.n377 B.n376 10.6151
R1397 B.n378 B.n377 10.6151
R1398 B.n380 B.n378 10.6151
R1399 B.n381 B.n380 10.6151
R1400 B.n382 B.n381 10.6151
R1401 B.n383 B.n382 10.6151
R1402 B.n579 B.n1 10.6151
R1403 B.n579 B.n578 10.6151
R1404 B.n578 B.n577 10.6151
R1405 B.n577 B.n10 10.6151
R1406 B.n571 B.n10 10.6151
R1407 B.n571 B.n570 10.6151
R1408 B.n570 B.n569 10.6151
R1409 B.n569 B.n18 10.6151
R1410 B.n563 B.n18 10.6151
R1411 B.n563 B.n562 10.6151
R1412 B.n562 B.n561 10.6151
R1413 B.n561 B.n25 10.6151
R1414 B.n555 B.n25 10.6151
R1415 B.n554 B.n553 10.6151
R1416 B.n553 B.n32 10.6151
R1417 B.n547 B.n32 10.6151
R1418 B.n547 B.n546 10.6151
R1419 B.n546 B.n545 10.6151
R1420 B.n545 B.n34 10.6151
R1421 B.n539 B.n34 10.6151
R1422 B.n539 B.n538 10.6151
R1423 B.n538 B.n537 10.6151
R1424 B.n537 B.n36 10.6151
R1425 B.n531 B.n36 10.6151
R1426 B.n531 B.n530 10.6151
R1427 B.n530 B.n529 10.6151
R1428 B.n529 B.n38 10.6151
R1429 B.n523 B.n38 10.6151
R1430 B.n523 B.n522 10.6151
R1431 B.n522 B.n521 10.6151
R1432 B.n521 B.n40 10.6151
R1433 B.n515 B.n40 10.6151
R1434 B.n515 B.n514 10.6151
R1435 B.n514 B.n513 10.6151
R1436 B.n513 B.n42 10.6151
R1437 B.n507 B.n42 10.6151
R1438 B.n507 B.n506 10.6151
R1439 B.n506 B.n505 10.6151
R1440 B.n505 B.n44 10.6151
R1441 B.n499 B.n44 10.6151
R1442 B.n499 B.n498 10.6151
R1443 B.n498 B.n497 10.6151
R1444 B.n497 B.n46 10.6151
R1445 B.n491 B.n46 10.6151
R1446 B.n491 B.n490 10.6151
R1447 B.n490 B.n489 10.6151
R1448 B.n489 B.n48 10.6151
R1449 B.n483 B.n48 10.6151
R1450 B.n483 B.n482 10.6151
R1451 B.n482 B.n481 10.6151
R1452 B.n477 B.n476 10.6151
R1453 B.n476 B.n54 10.6151
R1454 B.n471 B.n54 10.6151
R1455 B.n471 B.n470 10.6151
R1456 B.n470 B.n469 10.6151
R1457 B.n469 B.n56 10.6151
R1458 B.n463 B.n56 10.6151
R1459 B.n463 B.n462 10.6151
R1460 B.n460 B.n60 10.6151
R1461 B.n454 B.n60 10.6151
R1462 B.n454 B.n453 10.6151
R1463 B.n453 B.n452 10.6151
R1464 B.n452 B.n62 10.6151
R1465 B.n446 B.n62 10.6151
R1466 B.n446 B.n445 10.6151
R1467 B.n445 B.n444 10.6151
R1468 B.n444 B.n64 10.6151
R1469 B.n438 B.n64 10.6151
R1470 B.n438 B.n437 10.6151
R1471 B.n437 B.n436 10.6151
R1472 B.n436 B.n66 10.6151
R1473 B.n430 B.n66 10.6151
R1474 B.n430 B.n429 10.6151
R1475 B.n429 B.n428 10.6151
R1476 B.n428 B.n68 10.6151
R1477 B.n422 B.n68 10.6151
R1478 B.n422 B.n421 10.6151
R1479 B.n421 B.n420 10.6151
R1480 B.n420 B.n70 10.6151
R1481 B.n414 B.n70 10.6151
R1482 B.n414 B.n413 10.6151
R1483 B.n413 B.n412 10.6151
R1484 B.n412 B.n72 10.6151
R1485 B.n406 B.n72 10.6151
R1486 B.n406 B.n405 10.6151
R1487 B.n405 B.n404 10.6151
R1488 B.n404 B.n74 10.6151
R1489 B.n398 B.n74 10.6151
R1490 B.n398 B.n397 10.6151
R1491 B.n397 B.n396 10.6151
R1492 B.n396 B.n76 10.6151
R1493 B.n390 B.n76 10.6151
R1494 B.n390 B.n389 10.6151
R1495 B.n389 B.n388 10.6151
R1496 B.n388 B.n384 10.6151
R1497 B.n587 B.n0 8.11757
R1498 B.n587 B.n1 8.11757
R1499 B.n243 B.n127 7.18099
R1500 B.n227 B.n226 7.18099
R1501 B.n477 B.n52 7.18099
R1502 B.n462 B.n461 7.18099
R1503 B.n127 B.n123 3.43465
R1504 B.n226 B.n225 3.43465
R1505 B.n481 B.n52 3.43465
R1506 B.n461 B.n460 3.43465
R1507 B.t7 B.n91 1.37593
R1508 B.n566 B.t3 1.37593
R1509 VN VN.t0 601.994
R1510 VN VN.t1 562.909
R1511 VDD2.n109 VDD2.n57 289.615
R1512 VDD2.n52 VDD2.n0 289.615
R1513 VDD2.n110 VDD2.n109 185
R1514 VDD2.n108 VDD2.n107 185
R1515 VDD2.n61 VDD2.n60 185
R1516 VDD2.n102 VDD2.n101 185
R1517 VDD2.n100 VDD2.n99 185
R1518 VDD2.n98 VDD2.n64 185
R1519 VDD2.n68 VDD2.n65 185
R1520 VDD2.n93 VDD2.n92 185
R1521 VDD2.n91 VDD2.n90 185
R1522 VDD2.n70 VDD2.n69 185
R1523 VDD2.n85 VDD2.n84 185
R1524 VDD2.n83 VDD2.n82 185
R1525 VDD2.n74 VDD2.n73 185
R1526 VDD2.n77 VDD2.n76 185
R1527 VDD2.n19 VDD2.n18 185
R1528 VDD2.n16 VDD2.n15 185
R1529 VDD2.n25 VDD2.n24 185
R1530 VDD2.n27 VDD2.n26 185
R1531 VDD2.n12 VDD2.n11 185
R1532 VDD2.n33 VDD2.n32 185
R1533 VDD2.n36 VDD2.n35 185
R1534 VDD2.n34 VDD2.n8 185
R1535 VDD2.n41 VDD2.n7 185
R1536 VDD2.n43 VDD2.n42 185
R1537 VDD2.n45 VDD2.n44 185
R1538 VDD2.n4 VDD2.n3 185
R1539 VDD2.n51 VDD2.n50 185
R1540 VDD2.n53 VDD2.n52 185
R1541 VDD2.t1 VDD2.n75 149.524
R1542 VDD2.t0 VDD2.n17 149.524
R1543 VDD2.n109 VDD2.n108 104.615
R1544 VDD2.n108 VDD2.n60 104.615
R1545 VDD2.n101 VDD2.n60 104.615
R1546 VDD2.n101 VDD2.n100 104.615
R1547 VDD2.n100 VDD2.n64 104.615
R1548 VDD2.n68 VDD2.n64 104.615
R1549 VDD2.n92 VDD2.n68 104.615
R1550 VDD2.n92 VDD2.n91 104.615
R1551 VDD2.n91 VDD2.n69 104.615
R1552 VDD2.n84 VDD2.n69 104.615
R1553 VDD2.n84 VDD2.n83 104.615
R1554 VDD2.n83 VDD2.n73 104.615
R1555 VDD2.n76 VDD2.n73 104.615
R1556 VDD2.n18 VDD2.n15 104.615
R1557 VDD2.n25 VDD2.n15 104.615
R1558 VDD2.n26 VDD2.n25 104.615
R1559 VDD2.n26 VDD2.n11 104.615
R1560 VDD2.n33 VDD2.n11 104.615
R1561 VDD2.n35 VDD2.n33 104.615
R1562 VDD2.n35 VDD2.n34 104.615
R1563 VDD2.n34 VDD2.n7 104.615
R1564 VDD2.n43 VDD2.n7 104.615
R1565 VDD2.n44 VDD2.n43 104.615
R1566 VDD2.n44 VDD2.n3 104.615
R1567 VDD2.n51 VDD2.n3 104.615
R1568 VDD2.n52 VDD2.n51 104.615
R1569 VDD2.n114 VDD2.n56 83.9977
R1570 VDD2.n76 VDD2.t1 52.3082
R1571 VDD2.n18 VDD2.t0 52.3082
R1572 VDD2.n114 VDD2.n113 49.252
R1573 VDD2.n99 VDD2.n98 13.1884
R1574 VDD2.n42 VDD2.n41 13.1884
R1575 VDD2.n102 VDD2.n63 12.8005
R1576 VDD2.n97 VDD2.n65 12.8005
R1577 VDD2.n40 VDD2.n8 12.8005
R1578 VDD2.n45 VDD2.n6 12.8005
R1579 VDD2.n103 VDD2.n61 12.0247
R1580 VDD2.n94 VDD2.n93 12.0247
R1581 VDD2.n37 VDD2.n36 12.0247
R1582 VDD2.n46 VDD2.n4 12.0247
R1583 VDD2.n107 VDD2.n106 11.249
R1584 VDD2.n90 VDD2.n67 11.249
R1585 VDD2.n32 VDD2.n10 11.249
R1586 VDD2.n50 VDD2.n49 11.249
R1587 VDD2.n110 VDD2.n59 10.4732
R1588 VDD2.n89 VDD2.n70 10.4732
R1589 VDD2.n31 VDD2.n12 10.4732
R1590 VDD2.n53 VDD2.n2 10.4732
R1591 VDD2.n77 VDD2.n75 10.2747
R1592 VDD2.n19 VDD2.n17 10.2747
R1593 VDD2.n111 VDD2.n57 9.69747
R1594 VDD2.n86 VDD2.n85 9.69747
R1595 VDD2.n28 VDD2.n27 9.69747
R1596 VDD2.n54 VDD2.n0 9.69747
R1597 VDD2.n113 VDD2.n112 9.45567
R1598 VDD2.n56 VDD2.n55 9.45567
R1599 VDD2.n79 VDD2.n78 9.3005
R1600 VDD2.n81 VDD2.n80 9.3005
R1601 VDD2.n72 VDD2.n71 9.3005
R1602 VDD2.n87 VDD2.n86 9.3005
R1603 VDD2.n89 VDD2.n88 9.3005
R1604 VDD2.n67 VDD2.n66 9.3005
R1605 VDD2.n95 VDD2.n94 9.3005
R1606 VDD2.n97 VDD2.n96 9.3005
R1607 VDD2.n112 VDD2.n111 9.3005
R1608 VDD2.n59 VDD2.n58 9.3005
R1609 VDD2.n106 VDD2.n105 9.3005
R1610 VDD2.n104 VDD2.n103 9.3005
R1611 VDD2.n63 VDD2.n62 9.3005
R1612 VDD2.n55 VDD2.n54 9.3005
R1613 VDD2.n2 VDD2.n1 9.3005
R1614 VDD2.n49 VDD2.n48 9.3005
R1615 VDD2.n47 VDD2.n46 9.3005
R1616 VDD2.n6 VDD2.n5 9.3005
R1617 VDD2.n21 VDD2.n20 9.3005
R1618 VDD2.n23 VDD2.n22 9.3005
R1619 VDD2.n14 VDD2.n13 9.3005
R1620 VDD2.n29 VDD2.n28 9.3005
R1621 VDD2.n31 VDD2.n30 9.3005
R1622 VDD2.n10 VDD2.n9 9.3005
R1623 VDD2.n38 VDD2.n37 9.3005
R1624 VDD2.n40 VDD2.n39 9.3005
R1625 VDD2.n82 VDD2.n72 8.92171
R1626 VDD2.n24 VDD2.n14 8.92171
R1627 VDD2.n81 VDD2.n74 8.14595
R1628 VDD2.n23 VDD2.n16 8.14595
R1629 VDD2.n78 VDD2.n77 7.3702
R1630 VDD2.n20 VDD2.n19 7.3702
R1631 VDD2.n78 VDD2.n74 5.81868
R1632 VDD2.n20 VDD2.n16 5.81868
R1633 VDD2.n82 VDD2.n81 5.04292
R1634 VDD2.n24 VDD2.n23 5.04292
R1635 VDD2.n113 VDD2.n57 4.26717
R1636 VDD2.n85 VDD2.n72 4.26717
R1637 VDD2.n27 VDD2.n14 4.26717
R1638 VDD2.n56 VDD2.n0 4.26717
R1639 VDD2.n111 VDD2.n110 3.49141
R1640 VDD2.n86 VDD2.n70 3.49141
R1641 VDD2.n28 VDD2.n12 3.49141
R1642 VDD2.n54 VDD2.n53 3.49141
R1643 VDD2.n79 VDD2.n75 2.84303
R1644 VDD2.n21 VDD2.n17 2.84303
R1645 VDD2.n107 VDD2.n59 2.71565
R1646 VDD2.n90 VDD2.n89 2.71565
R1647 VDD2.n32 VDD2.n31 2.71565
R1648 VDD2.n50 VDD2.n2 2.71565
R1649 VDD2.n106 VDD2.n61 1.93989
R1650 VDD2.n93 VDD2.n67 1.93989
R1651 VDD2.n36 VDD2.n10 1.93989
R1652 VDD2.n49 VDD2.n4 1.93989
R1653 VDD2.n103 VDD2.n102 1.16414
R1654 VDD2.n94 VDD2.n65 1.16414
R1655 VDD2.n37 VDD2.n8 1.16414
R1656 VDD2.n46 VDD2.n45 1.16414
R1657 VDD2.n99 VDD2.n63 0.388379
R1658 VDD2.n98 VDD2.n97 0.388379
R1659 VDD2.n41 VDD2.n40 0.388379
R1660 VDD2.n42 VDD2.n6 0.388379
R1661 VDD2 VDD2.n114 0.289293
R1662 VDD2.n112 VDD2.n58 0.155672
R1663 VDD2.n105 VDD2.n58 0.155672
R1664 VDD2.n105 VDD2.n104 0.155672
R1665 VDD2.n104 VDD2.n62 0.155672
R1666 VDD2.n96 VDD2.n62 0.155672
R1667 VDD2.n96 VDD2.n95 0.155672
R1668 VDD2.n95 VDD2.n66 0.155672
R1669 VDD2.n88 VDD2.n66 0.155672
R1670 VDD2.n88 VDD2.n87 0.155672
R1671 VDD2.n87 VDD2.n71 0.155672
R1672 VDD2.n80 VDD2.n71 0.155672
R1673 VDD2.n80 VDD2.n79 0.155672
R1674 VDD2.n22 VDD2.n21 0.155672
R1675 VDD2.n22 VDD2.n13 0.155672
R1676 VDD2.n29 VDD2.n13 0.155672
R1677 VDD2.n30 VDD2.n29 0.155672
R1678 VDD2.n30 VDD2.n9 0.155672
R1679 VDD2.n38 VDD2.n9 0.155672
R1680 VDD2.n39 VDD2.n38 0.155672
R1681 VDD2.n39 VDD2.n5 0.155672
R1682 VDD2.n47 VDD2.n5 0.155672
R1683 VDD2.n48 VDD2.n47 0.155672
R1684 VDD2.n48 VDD2.n1 0.155672
R1685 VDD2.n55 VDD2.n1 0.155672
C0 VTAIL VN 1.38804f
C1 VTAIL VDD1 5.1207f
C2 VP VN 4.337f
C3 VDD2 VTAIL 5.15568f
C4 VP VDD1 1.93408f
C5 VDD1 VN 0.14894f
C6 VDD2 VP 0.256798f
C7 VDD2 VN 1.83006f
C8 VDD2 VDD1 0.465632f
C9 VTAIL VP 1.40258f
C10 VDD2 B 3.523321f
C11 VDD1 B 5.23227f
C12 VTAIL B 5.903802f
C13 VN B 6.71103f
C14 VP B 3.986009f
C15 VDD2.n0 B 0.021233f
C16 VDD2.n1 B 0.015554f
C17 VDD2.n2 B 0.008358f
C18 VDD2.n3 B 0.019755f
C19 VDD2.n4 B 0.00885f
C20 VDD2.n5 B 0.015554f
C21 VDD2.n6 B 0.008358f
C22 VDD2.n7 B 0.019755f
C23 VDD2.n8 B 0.00885f
C24 VDD2.n9 B 0.015554f
C25 VDD2.n10 B 0.008358f
C26 VDD2.n11 B 0.019755f
C27 VDD2.n12 B 0.00885f
C28 VDD2.n13 B 0.015554f
C29 VDD2.n14 B 0.008358f
C30 VDD2.n15 B 0.019755f
C31 VDD2.n16 B 0.00885f
C32 VDD2.n17 B 0.104381f
C33 VDD2.t0 B 0.033257f
C34 VDD2.n18 B 0.014817f
C35 VDD2.n19 B 0.013966f
C36 VDD2.n20 B 0.008358f
C37 VDD2.n21 B 0.694735f
C38 VDD2.n22 B 0.015554f
C39 VDD2.n23 B 0.008358f
C40 VDD2.n24 B 0.00885f
C41 VDD2.n25 B 0.019755f
C42 VDD2.n26 B 0.019755f
C43 VDD2.n27 B 0.00885f
C44 VDD2.n28 B 0.008358f
C45 VDD2.n29 B 0.015554f
C46 VDD2.n30 B 0.015554f
C47 VDD2.n31 B 0.008358f
C48 VDD2.n32 B 0.00885f
C49 VDD2.n33 B 0.019755f
C50 VDD2.n34 B 0.019755f
C51 VDD2.n35 B 0.019755f
C52 VDD2.n36 B 0.00885f
C53 VDD2.n37 B 0.008358f
C54 VDD2.n38 B 0.015554f
C55 VDD2.n39 B 0.015554f
C56 VDD2.n40 B 0.008358f
C57 VDD2.n41 B 0.008604f
C58 VDD2.n42 B 0.008604f
C59 VDD2.n43 B 0.019755f
C60 VDD2.n44 B 0.019755f
C61 VDD2.n45 B 0.00885f
C62 VDD2.n46 B 0.008358f
C63 VDD2.n47 B 0.015554f
C64 VDD2.n48 B 0.015554f
C65 VDD2.n49 B 0.008358f
C66 VDD2.n50 B 0.00885f
C67 VDD2.n51 B 0.019755f
C68 VDD2.n52 B 0.041654f
C69 VDD2.n53 B 0.00885f
C70 VDD2.n54 B 0.008358f
C71 VDD2.n55 B 0.036377f
C72 VDD2.n56 B 0.355f
C73 VDD2.n57 B 0.021233f
C74 VDD2.n58 B 0.015554f
C75 VDD2.n59 B 0.008358f
C76 VDD2.n60 B 0.019755f
C77 VDD2.n61 B 0.00885f
C78 VDD2.n62 B 0.015554f
C79 VDD2.n63 B 0.008358f
C80 VDD2.n64 B 0.019755f
C81 VDD2.n65 B 0.00885f
C82 VDD2.n66 B 0.015554f
C83 VDD2.n67 B 0.008358f
C84 VDD2.n68 B 0.019755f
C85 VDD2.n69 B 0.019755f
C86 VDD2.n70 B 0.00885f
C87 VDD2.n71 B 0.015554f
C88 VDD2.n72 B 0.008358f
C89 VDD2.n73 B 0.019755f
C90 VDD2.n74 B 0.00885f
C91 VDD2.n75 B 0.104381f
C92 VDD2.t1 B 0.033257f
C93 VDD2.n76 B 0.014817f
C94 VDD2.n77 B 0.013966f
C95 VDD2.n78 B 0.008358f
C96 VDD2.n79 B 0.694735f
C97 VDD2.n80 B 0.015554f
C98 VDD2.n81 B 0.008358f
C99 VDD2.n82 B 0.00885f
C100 VDD2.n83 B 0.019755f
C101 VDD2.n84 B 0.019755f
C102 VDD2.n85 B 0.00885f
C103 VDD2.n86 B 0.008358f
C104 VDD2.n87 B 0.015554f
C105 VDD2.n88 B 0.015554f
C106 VDD2.n89 B 0.008358f
C107 VDD2.n90 B 0.00885f
C108 VDD2.n91 B 0.019755f
C109 VDD2.n92 B 0.019755f
C110 VDD2.n93 B 0.00885f
C111 VDD2.n94 B 0.008358f
C112 VDD2.n95 B 0.015554f
C113 VDD2.n96 B 0.015554f
C114 VDD2.n97 B 0.008358f
C115 VDD2.n98 B 0.008604f
C116 VDD2.n99 B 0.008604f
C117 VDD2.n100 B 0.019755f
C118 VDD2.n101 B 0.019755f
C119 VDD2.n102 B 0.00885f
C120 VDD2.n103 B 0.008358f
C121 VDD2.n104 B 0.015554f
C122 VDD2.n105 B 0.015554f
C123 VDD2.n106 B 0.008358f
C124 VDD2.n107 B 0.00885f
C125 VDD2.n108 B 0.019755f
C126 VDD2.n109 B 0.041654f
C127 VDD2.n110 B 0.00885f
C128 VDD2.n111 B 0.008358f
C129 VDD2.n112 B 0.036377f
C130 VDD2.n113 B 0.033942f
C131 VDD2.n114 B 1.58946f
C132 VN.t1 B 0.786535f
C133 VN.t0 B 0.87411f
C134 VDD1.n0 B 0.020597f
C135 VDD1.n1 B 0.015088f
C136 VDD1.n2 B 0.008108f
C137 VDD1.n3 B 0.019164f
C138 VDD1.n4 B 0.008585f
C139 VDD1.n5 B 0.015088f
C140 VDD1.n6 B 0.008108f
C141 VDD1.n7 B 0.019164f
C142 VDD1.n8 B 0.008585f
C143 VDD1.n9 B 0.015088f
C144 VDD1.n10 B 0.008108f
C145 VDD1.n11 B 0.019164f
C146 VDD1.n12 B 0.019164f
C147 VDD1.n13 B 0.008585f
C148 VDD1.n14 B 0.015088f
C149 VDD1.n15 B 0.008108f
C150 VDD1.n16 B 0.019164f
C151 VDD1.n17 B 0.008585f
C152 VDD1.n18 B 0.101255f
C153 VDD1.t1 B 0.032261f
C154 VDD1.n19 B 0.014373f
C155 VDD1.n20 B 0.013547f
C156 VDD1.n21 B 0.008108f
C157 VDD1.n22 B 0.67393f
C158 VDD1.n23 B 0.015088f
C159 VDD1.n24 B 0.008108f
C160 VDD1.n25 B 0.008585f
C161 VDD1.n26 B 0.019164f
C162 VDD1.n27 B 0.019164f
C163 VDD1.n28 B 0.008585f
C164 VDD1.n29 B 0.008108f
C165 VDD1.n30 B 0.015088f
C166 VDD1.n31 B 0.015088f
C167 VDD1.n32 B 0.008108f
C168 VDD1.n33 B 0.008585f
C169 VDD1.n34 B 0.019164f
C170 VDD1.n35 B 0.019164f
C171 VDD1.n36 B 0.008585f
C172 VDD1.n37 B 0.008108f
C173 VDD1.n38 B 0.015088f
C174 VDD1.n39 B 0.015088f
C175 VDD1.n40 B 0.008108f
C176 VDD1.n41 B 0.008346f
C177 VDD1.n42 B 0.008346f
C178 VDD1.n43 B 0.019164f
C179 VDD1.n44 B 0.019164f
C180 VDD1.n45 B 0.008585f
C181 VDD1.n46 B 0.008108f
C182 VDD1.n47 B 0.015088f
C183 VDD1.n48 B 0.015088f
C184 VDD1.n49 B 0.008108f
C185 VDD1.n50 B 0.008585f
C186 VDD1.n51 B 0.019164f
C187 VDD1.n52 B 0.040406f
C188 VDD1.n53 B 0.008585f
C189 VDD1.n54 B 0.008108f
C190 VDD1.n55 B 0.035288f
C191 VDD1.n56 B 0.033178f
C192 VDD1.n57 B 0.020597f
C193 VDD1.n58 B 0.015088f
C194 VDD1.n59 B 0.008108f
C195 VDD1.n60 B 0.019164f
C196 VDD1.n61 B 0.008585f
C197 VDD1.n62 B 0.015088f
C198 VDD1.n63 B 0.008108f
C199 VDD1.n64 B 0.019164f
C200 VDD1.n65 B 0.008585f
C201 VDD1.n66 B 0.015088f
C202 VDD1.n67 B 0.008108f
C203 VDD1.n68 B 0.019164f
C204 VDD1.n69 B 0.008585f
C205 VDD1.n70 B 0.015088f
C206 VDD1.n71 B 0.008108f
C207 VDD1.n72 B 0.019164f
C208 VDD1.n73 B 0.008585f
C209 VDD1.n74 B 0.101255f
C210 VDD1.t0 B 0.032261f
C211 VDD1.n75 B 0.014373f
C212 VDD1.n76 B 0.013547f
C213 VDD1.n77 B 0.008108f
C214 VDD1.n78 B 0.67393f
C215 VDD1.n79 B 0.015088f
C216 VDD1.n80 B 0.008108f
C217 VDD1.n81 B 0.008585f
C218 VDD1.n82 B 0.019164f
C219 VDD1.n83 B 0.019164f
C220 VDD1.n84 B 0.008585f
C221 VDD1.n85 B 0.008108f
C222 VDD1.n86 B 0.015088f
C223 VDD1.n87 B 0.015088f
C224 VDD1.n88 B 0.008108f
C225 VDD1.n89 B 0.008585f
C226 VDD1.n90 B 0.019164f
C227 VDD1.n91 B 0.019164f
C228 VDD1.n92 B 0.019164f
C229 VDD1.n93 B 0.008585f
C230 VDD1.n94 B 0.008108f
C231 VDD1.n95 B 0.015088f
C232 VDD1.n96 B 0.015088f
C233 VDD1.n97 B 0.008108f
C234 VDD1.n98 B 0.008346f
C235 VDD1.n99 B 0.008346f
C236 VDD1.n100 B 0.019164f
C237 VDD1.n101 B 0.019164f
C238 VDD1.n102 B 0.008585f
C239 VDD1.n103 B 0.008108f
C240 VDD1.n104 B 0.015088f
C241 VDD1.n105 B 0.015088f
C242 VDD1.n106 B 0.008108f
C243 VDD1.n107 B 0.008585f
C244 VDD1.n108 B 0.019164f
C245 VDD1.n109 B 0.040406f
C246 VDD1.n110 B 0.008585f
C247 VDD1.n111 B 0.008108f
C248 VDD1.n112 B 0.035288f
C249 VDD1.n113 B 0.364142f
C250 VTAIL.n0 B 0.022603f
C251 VTAIL.n1 B 0.016557f
C252 VTAIL.n2 B 0.008897f
C253 VTAIL.n3 B 0.02103f
C254 VTAIL.n4 B 0.009421f
C255 VTAIL.n5 B 0.016557f
C256 VTAIL.n6 B 0.008897f
C257 VTAIL.n7 B 0.02103f
C258 VTAIL.n8 B 0.009421f
C259 VTAIL.n9 B 0.016557f
C260 VTAIL.n10 B 0.008897f
C261 VTAIL.n11 B 0.02103f
C262 VTAIL.n12 B 0.009421f
C263 VTAIL.n13 B 0.016557f
C264 VTAIL.n14 B 0.008897f
C265 VTAIL.n15 B 0.02103f
C266 VTAIL.n16 B 0.009421f
C267 VTAIL.n17 B 0.111113f
C268 VTAIL.t3 B 0.035402f
C269 VTAIL.n18 B 0.015772f
C270 VTAIL.n19 B 0.014866f
C271 VTAIL.n20 B 0.008897f
C272 VTAIL.n21 B 0.739547f
C273 VTAIL.n22 B 0.016557f
C274 VTAIL.n23 B 0.008897f
C275 VTAIL.n24 B 0.009421f
C276 VTAIL.n25 B 0.02103f
C277 VTAIL.n26 B 0.02103f
C278 VTAIL.n27 B 0.009421f
C279 VTAIL.n28 B 0.008897f
C280 VTAIL.n29 B 0.016557f
C281 VTAIL.n30 B 0.016557f
C282 VTAIL.n31 B 0.008897f
C283 VTAIL.n32 B 0.009421f
C284 VTAIL.n33 B 0.02103f
C285 VTAIL.n34 B 0.02103f
C286 VTAIL.n35 B 0.02103f
C287 VTAIL.n36 B 0.009421f
C288 VTAIL.n37 B 0.008897f
C289 VTAIL.n38 B 0.016557f
C290 VTAIL.n39 B 0.016557f
C291 VTAIL.n40 B 0.008897f
C292 VTAIL.n41 B 0.009159f
C293 VTAIL.n42 B 0.009159f
C294 VTAIL.n43 B 0.02103f
C295 VTAIL.n44 B 0.02103f
C296 VTAIL.n45 B 0.009421f
C297 VTAIL.n46 B 0.008897f
C298 VTAIL.n47 B 0.016557f
C299 VTAIL.n48 B 0.016557f
C300 VTAIL.n49 B 0.008897f
C301 VTAIL.n50 B 0.009421f
C302 VTAIL.n51 B 0.02103f
C303 VTAIL.n52 B 0.04434f
C304 VTAIL.n53 B 0.009421f
C305 VTAIL.n54 B 0.008897f
C306 VTAIL.n55 B 0.038724f
C307 VTAIL.n56 B 0.024702f
C308 VTAIL.n57 B 0.871244f
C309 VTAIL.n58 B 0.022603f
C310 VTAIL.n59 B 0.016557f
C311 VTAIL.n60 B 0.008897f
C312 VTAIL.n61 B 0.02103f
C313 VTAIL.n62 B 0.009421f
C314 VTAIL.n63 B 0.016557f
C315 VTAIL.n64 B 0.008897f
C316 VTAIL.n65 B 0.02103f
C317 VTAIL.n66 B 0.009421f
C318 VTAIL.n67 B 0.016557f
C319 VTAIL.n68 B 0.008897f
C320 VTAIL.n69 B 0.02103f
C321 VTAIL.n70 B 0.02103f
C322 VTAIL.n71 B 0.009421f
C323 VTAIL.n72 B 0.016557f
C324 VTAIL.n73 B 0.008897f
C325 VTAIL.n74 B 0.02103f
C326 VTAIL.n75 B 0.009421f
C327 VTAIL.n76 B 0.111113f
C328 VTAIL.t0 B 0.035402f
C329 VTAIL.n77 B 0.015772f
C330 VTAIL.n78 B 0.014866f
C331 VTAIL.n79 B 0.008897f
C332 VTAIL.n80 B 0.739547f
C333 VTAIL.n81 B 0.016557f
C334 VTAIL.n82 B 0.008897f
C335 VTAIL.n83 B 0.009421f
C336 VTAIL.n84 B 0.02103f
C337 VTAIL.n85 B 0.02103f
C338 VTAIL.n86 B 0.009421f
C339 VTAIL.n87 B 0.008897f
C340 VTAIL.n88 B 0.016557f
C341 VTAIL.n89 B 0.016557f
C342 VTAIL.n90 B 0.008897f
C343 VTAIL.n91 B 0.009421f
C344 VTAIL.n92 B 0.02103f
C345 VTAIL.n93 B 0.02103f
C346 VTAIL.n94 B 0.009421f
C347 VTAIL.n95 B 0.008897f
C348 VTAIL.n96 B 0.016557f
C349 VTAIL.n97 B 0.016557f
C350 VTAIL.n98 B 0.008897f
C351 VTAIL.n99 B 0.009159f
C352 VTAIL.n100 B 0.009159f
C353 VTAIL.n101 B 0.02103f
C354 VTAIL.n102 B 0.02103f
C355 VTAIL.n103 B 0.009421f
C356 VTAIL.n104 B 0.008897f
C357 VTAIL.n105 B 0.016557f
C358 VTAIL.n106 B 0.016557f
C359 VTAIL.n107 B 0.008897f
C360 VTAIL.n108 B 0.009421f
C361 VTAIL.n109 B 0.02103f
C362 VTAIL.n110 B 0.04434f
C363 VTAIL.n111 B 0.009421f
C364 VTAIL.n112 B 0.008897f
C365 VTAIL.n113 B 0.038724f
C366 VTAIL.n114 B 0.024702f
C367 VTAIL.n115 B 0.880443f
C368 VTAIL.n116 B 0.022603f
C369 VTAIL.n117 B 0.016557f
C370 VTAIL.n118 B 0.008897f
C371 VTAIL.n119 B 0.02103f
C372 VTAIL.n120 B 0.009421f
C373 VTAIL.n121 B 0.016557f
C374 VTAIL.n122 B 0.008897f
C375 VTAIL.n123 B 0.02103f
C376 VTAIL.n124 B 0.009421f
C377 VTAIL.n125 B 0.016557f
C378 VTAIL.n126 B 0.008897f
C379 VTAIL.n127 B 0.02103f
C380 VTAIL.n128 B 0.02103f
C381 VTAIL.n129 B 0.009421f
C382 VTAIL.n130 B 0.016557f
C383 VTAIL.n131 B 0.008897f
C384 VTAIL.n132 B 0.02103f
C385 VTAIL.n133 B 0.009421f
C386 VTAIL.n134 B 0.111113f
C387 VTAIL.t2 B 0.035402f
C388 VTAIL.n135 B 0.015772f
C389 VTAIL.n136 B 0.014866f
C390 VTAIL.n137 B 0.008897f
C391 VTAIL.n138 B 0.739547f
C392 VTAIL.n139 B 0.016557f
C393 VTAIL.n140 B 0.008897f
C394 VTAIL.n141 B 0.009421f
C395 VTAIL.n142 B 0.02103f
C396 VTAIL.n143 B 0.02103f
C397 VTAIL.n144 B 0.009421f
C398 VTAIL.n145 B 0.008897f
C399 VTAIL.n146 B 0.016557f
C400 VTAIL.n147 B 0.016557f
C401 VTAIL.n148 B 0.008897f
C402 VTAIL.n149 B 0.009421f
C403 VTAIL.n150 B 0.02103f
C404 VTAIL.n151 B 0.02103f
C405 VTAIL.n152 B 0.009421f
C406 VTAIL.n153 B 0.008897f
C407 VTAIL.n154 B 0.016557f
C408 VTAIL.n155 B 0.016557f
C409 VTAIL.n156 B 0.008897f
C410 VTAIL.n157 B 0.009159f
C411 VTAIL.n158 B 0.009159f
C412 VTAIL.n159 B 0.02103f
C413 VTAIL.n160 B 0.02103f
C414 VTAIL.n161 B 0.009421f
C415 VTAIL.n162 B 0.008897f
C416 VTAIL.n163 B 0.016557f
C417 VTAIL.n164 B 0.016557f
C418 VTAIL.n165 B 0.008897f
C419 VTAIL.n166 B 0.009421f
C420 VTAIL.n167 B 0.02103f
C421 VTAIL.n168 B 0.04434f
C422 VTAIL.n169 B 0.009421f
C423 VTAIL.n170 B 0.008897f
C424 VTAIL.n171 B 0.038724f
C425 VTAIL.n172 B 0.024702f
C426 VTAIL.n173 B 0.831231f
C427 VTAIL.n174 B 0.022603f
C428 VTAIL.n175 B 0.016557f
C429 VTAIL.n176 B 0.008897f
C430 VTAIL.n177 B 0.02103f
C431 VTAIL.n178 B 0.009421f
C432 VTAIL.n179 B 0.016557f
C433 VTAIL.n180 B 0.008897f
C434 VTAIL.n181 B 0.02103f
C435 VTAIL.n182 B 0.009421f
C436 VTAIL.n183 B 0.016557f
C437 VTAIL.n184 B 0.008897f
C438 VTAIL.n185 B 0.02103f
C439 VTAIL.n186 B 0.009421f
C440 VTAIL.n187 B 0.016557f
C441 VTAIL.n188 B 0.008897f
C442 VTAIL.n189 B 0.02103f
C443 VTAIL.n190 B 0.009421f
C444 VTAIL.n191 B 0.111113f
C445 VTAIL.t1 B 0.035402f
C446 VTAIL.n192 B 0.015772f
C447 VTAIL.n193 B 0.014866f
C448 VTAIL.n194 B 0.008897f
C449 VTAIL.n195 B 0.739547f
C450 VTAIL.n196 B 0.016557f
C451 VTAIL.n197 B 0.008897f
C452 VTAIL.n198 B 0.009421f
C453 VTAIL.n199 B 0.02103f
C454 VTAIL.n200 B 0.02103f
C455 VTAIL.n201 B 0.009421f
C456 VTAIL.n202 B 0.008897f
C457 VTAIL.n203 B 0.016557f
C458 VTAIL.n204 B 0.016557f
C459 VTAIL.n205 B 0.008897f
C460 VTAIL.n206 B 0.009421f
C461 VTAIL.n207 B 0.02103f
C462 VTAIL.n208 B 0.02103f
C463 VTAIL.n209 B 0.02103f
C464 VTAIL.n210 B 0.009421f
C465 VTAIL.n211 B 0.008897f
C466 VTAIL.n212 B 0.016557f
C467 VTAIL.n213 B 0.016557f
C468 VTAIL.n214 B 0.008897f
C469 VTAIL.n215 B 0.009159f
C470 VTAIL.n216 B 0.009159f
C471 VTAIL.n217 B 0.02103f
C472 VTAIL.n218 B 0.02103f
C473 VTAIL.n219 B 0.009421f
C474 VTAIL.n220 B 0.008897f
C475 VTAIL.n221 B 0.016557f
C476 VTAIL.n222 B 0.016557f
C477 VTAIL.n223 B 0.008897f
C478 VTAIL.n224 B 0.009421f
C479 VTAIL.n225 B 0.02103f
C480 VTAIL.n226 B 0.04434f
C481 VTAIL.n227 B 0.009421f
C482 VTAIL.n228 B 0.008897f
C483 VTAIL.n229 B 0.038724f
C484 VTAIL.n230 B 0.024702f
C485 VTAIL.n231 B 0.790757f
C486 VP.t0 B 0.880973f
C487 VP.t1 B 0.79462f
C488 VP.n0 B 2.61265f
.ends

