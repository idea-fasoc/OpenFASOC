* NGSPICE file created from diff_pair_sample_1736.ext - technology: sky130A

.subckt diff_pair_sample_1736 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=5.2182 ps=27.54 w=13.38 l=0.67
X1 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=0 ps=0 w=13.38 l=0.67
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=0 ps=0 w=13.38 l=0.67
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=5.2182 ps=27.54 w=13.38 l=0.67
X4 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=5.2182 ps=27.54 w=13.38 l=0.67
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=0 ps=0 w=13.38 l=0.67
X6 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=5.2182 ps=27.54 w=13.38 l=0.67
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.2182 pd=27.54 as=0 ps=0 w=13.38 l=0.67
R0 VN VN.t0 742.912
R1 VN VN.t1 701.982
R2 VTAIL.n282 VTAIL.n216 214.453
R3 VTAIL.n66 VTAIL.n0 214.453
R4 VTAIL.n210 VTAIL.n144 214.453
R5 VTAIL.n138 VTAIL.n72 214.453
R6 VTAIL.n241 VTAIL.n240 185
R7 VTAIL.n243 VTAIL.n242 185
R8 VTAIL.n236 VTAIL.n235 185
R9 VTAIL.n249 VTAIL.n248 185
R10 VTAIL.n251 VTAIL.n250 185
R11 VTAIL.n232 VTAIL.n231 185
R12 VTAIL.n257 VTAIL.n256 185
R13 VTAIL.n259 VTAIL.n258 185
R14 VTAIL.n228 VTAIL.n227 185
R15 VTAIL.n265 VTAIL.n264 185
R16 VTAIL.n267 VTAIL.n266 185
R17 VTAIL.n224 VTAIL.n223 185
R18 VTAIL.n273 VTAIL.n272 185
R19 VTAIL.n275 VTAIL.n274 185
R20 VTAIL.n220 VTAIL.n219 185
R21 VTAIL.n281 VTAIL.n280 185
R22 VTAIL.n283 VTAIL.n282 185
R23 VTAIL.n25 VTAIL.n24 185
R24 VTAIL.n27 VTAIL.n26 185
R25 VTAIL.n20 VTAIL.n19 185
R26 VTAIL.n33 VTAIL.n32 185
R27 VTAIL.n35 VTAIL.n34 185
R28 VTAIL.n16 VTAIL.n15 185
R29 VTAIL.n41 VTAIL.n40 185
R30 VTAIL.n43 VTAIL.n42 185
R31 VTAIL.n12 VTAIL.n11 185
R32 VTAIL.n49 VTAIL.n48 185
R33 VTAIL.n51 VTAIL.n50 185
R34 VTAIL.n8 VTAIL.n7 185
R35 VTAIL.n57 VTAIL.n56 185
R36 VTAIL.n59 VTAIL.n58 185
R37 VTAIL.n4 VTAIL.n3 185
R38 VTAIL.n65 VTAIL.n64 185
R39 VTAIL.n67 VTAIL.n66 185
R40 VTAIL.n211 VTAIL.n210 185
R41 VTAIL.n209 VTAIL.n208 185
R42 VTAIL.n148 VTAIL.n147 185
R43 VTAIL.n203 VTAIL.n202 185
R44 VTAIL.n201 VTAIL.n200 185
R45 VTAIL.n152 VTAIL.n151 185
R46 VTAIL.n195 VTAIL.n194 185
R47 VTAIL.n193 VTAIL.n192 185
R48 VTAIL.n156 VTAIL.n155 185
R49 VTAIL.n187 VTAIL.n186 185
R50 VTAIL.n185 VTAIL.n184 185
R51 VTAIL.n160 VTAIL.n159 185
R52 VTAIL.n179 VTAIL.n178 185
R53 VTAIL.n177 VTAIL.n176 185
R54 VTAIL.n164 VTAIL.n163 185
R55 VTAIL.n171 VTAIL.n170 185
R56 VTAIL.n169 VTAIL.n168 185
R57 VTAIL.n139 VTAIL.n138 185
R58 VTAIL.n137 VTAIL.n136 185
R59 VTAIL.n76 VTAIL.n75 185
R60 VTAIL.n131 VTAIL.n130 185
R61 VTAIL.n129 VTAIL.n128 185
R62 VTAIL.n80 VTAIL.n79 185
R63 VTAIL.n123 VTAIL.n122 185
R64 VTAIL.n121 VTAIL.n120 185
R65 VTAIL.n84 VTAIL.n83 185
R66 VTAIL.n115 VTAIL.n114 185
R67 VTAIL.n113 VTAIL.n112 185
R68 VTAIL.n88 VTAIL.n87 185
R69 VTAIL.n107 VTAIL.n106 185
R70 VTAIL.n105 VTAIL.n104 185
R71 VTAIL.n92 VTAIL.n91 185
R72 VTAIL.n99 VTAIL.n98 185
R73 VTAIL.n97 VTAIL.n96 185
R74 VTAIL.n239 VTAIL.t3 147.659
R75 VTAIL.n23 VTAIL.t0 147.659
R76 VTAIL.n167 VTAIL.t1 147.659
R77 VTAIL.n95 VTAIL.t2 147.659
R78 VTAIL.n242 VTAIL.n241 104.615
R79 VTAIL.n242 VTAIL.n235 104.615
R80 VTAIL.n249 VTAIL.n235 104.615
R81 VTAIL.n250 VTAIL.n249 104.615
R82 VTAIL.n250 VTAIL.n231 104.615
R83 VTAIL.n257 VTAIL.n231 104.615
R84 VTAIL.n258 VTAIL.n257 104.615
R85 VTAIL.n258 VTAIL.n227 104.615
R86 VTAIL.n265 VTAIL.n227 104.615
R87 VTAIL.n266 VTAIL.n265 104.615
R88 VTAIL.n266 VTAIL.n223 104.615
R89 VTAIL.n273 VTAIL.n223 104.615
R90 VTAIL.n274 VTAIL.n273 104.615
R91 VTAIL.n274 VTAIL.n219 104.615
R92 VTAIL.n281 VTAIL.n219 104.615
R93 VTAIL.n282 VTAIL.n281 104.615
R94 VTAIL.n26 VTAIL.n25 104.615
R95 VTAIL.n26 VTAIL.n19 104.615
R96 VTAIL.n33 VTAIL.n19 104.615
R97 VTAIL.n34 VTAIL.n33 104.615
R98 VTAIL.n34 VTAIL.n15 104.615
R99 VTAIL.n41 VTAIL.n15 104.615
R100 VTAIL.n42 VTAIL.n41 104.615
R101 VTAIL.n42 VTAIL.n11 104.615
R102 VTAIL.n49 VTAIL.n11 104.615
R103 VTAIL.n50 VTAIL.n49 104.615
R104 VTAIL.n50 VTAIL.n7 104.615
R105 VTAIL.n57 VTAIL.n7 104.615
R106 VTAIL.n58 VTAIL.n57 104.615
R107 VTAIL.n58 VTAIL.n3 104.615
R108 VTAIL.n65 VTAIL.n3 104.615
R109 VTAIL.n66 VTAIL.n65 104.615
R110 VTAIL.n210 VTAIL.n209 104.615
R111 VTAIL.n209 VTAIL.n147 104.615
R112 VTAIL.n202 VTAIL.n147 104.615
R113 VTAIL.n202 VTAIL.n201 104.615
R114 VTAIL.n201 VTAIL.n151 104.615
R115 VTAIL.n194 VTAIL.n151 104.615
R116 VTAIL.n194 VTAIL.n193 104.615
R117 VTAIL.n193 VTAIL.n155 104.615
R118 VTAIL.n186 VTAIL.n155 104.615
R119 VTAIL.n186 VTAIL.n185 104.615
R120 VTAIL.n185 VTAIL.n159 104.615
R121 VTAIL.n178 VTAIL.n159 104.615
R122 VTAIL.n178 VTAIL.n177 104.615
R123 VTAIL.n177 VTAIL.n163 104.615
R124 VTAIL.n170 VTAIL.n163 104.615
R125 VTAIL.n170 VTAIL.n169 104.615
R126 VTAIL.n138 VTAIL.n137 104.615
R127 VTAIL.n137 VTAIL.n75 104.615
R128 VTAIL.n130 VTAIL.n75 104.615
R129 VTAIL.n130 VTAIL.n129 104.615
R130 VTAIL.n129 VTAIL.n79 104.615
R131 VTAIL.n122 VTAIL.n79 104.615
R132 VTAIL.n122 VTAIL.n121 104.615
R133 VTAIL.n121 VTAIL.n83 104.615
R134 VTAIL.n114 VTAIL.n83 104.615
R135 VTAIL.n114 VTAIL.n113 104.615
R136 VTAIL.n113 VTAIL.n87 104.615
R137 VTAIL.n106 VTAIL.n87 104.615
R138 VTAIL.n106 VTAIL.n105 104.615
R139 VTAIL.n105 VTAIL.n91 104.615
R140 VTAIL.n98 VTAIL.n91 104.615
R141 VTAIL.n98 VTAIL.n97 104.615
R142 VTAIL.n241 VTAIL.t3 52.3082
R143 VTAIL.n25 VTAIL.t0 52.3082
R144 VTAIL.n169 VTAIL.t1 52.3082
R145 VTAIL.n97 VTAIL.t2 52.3082
R146 VTAIL.n287 VTAIL.n286 35.6763
R147 VTAIL.n71 VTAIL.n70 35.6763
R148 VTAIL.n215 VTAIL.n214 35.6763
R149 VTAIL.n143 VTAIL.n142 35.6763
R150 VTAIL.n143 VTAIL.n71 25.6427
R151 VTAIL.n287 VTAIL.n215 24.7807
R152 VTAIL.n240 VTAIL.n239 15.6677
R153 VTAIL.n24 VTAIL.n23 15.6677
R154 VTAIL.n168 VTAIL.n167 15.6677
R155 VTAIL.n96 VTAIL.n95 15.6677
R156 VTAIL.n243 VTAIL.n238 12.8005
R157 VTAIL.n284 VTAIL.n283 12.8005
R158 VTAIL.n27 VTAIL.n22 12.8005
R159 VTAIL.n68 VTAIL.n67 12.8005
R160 VTAIL.n212 VTAIL.n211 12.8005
R161 VTAIL.n171 VTAIL.n166 12.8005
R162 VTAIL.n140 VTAIL.n139 12.8005
R163 VTAIL.n99 VTAIL.n94 12.8005
R164 VTAIL.n244 VTAIL.n236 12.0247
R165 VTAIL.n280 VTAIL.n218 12.0247
R166 VTAIL.n28 VTAIL.n20 12.0247
R167 VTAIL.n64 VTAIL.n2 12.0247
R168 VTAIL.n208 VTAIL.n146 12.0247
R169 VTAIL.n172 VTAIL.n164 12.0247
R170 VTAIL.n136 VTAIL.n74 12.0247
R171 VTAIL.n100 VTAIL.n92 12.0247
R172 VTAIL.n248 VTAIL.n247 11.249
R173 VTAIL.n279 VTAIL.n220 11.249
R174 VTAIL.n32 VTAIL.n31 11.249
R175 VTAIL.n63 VTAIL.n4 11.249
R176 VTAIL.n207 VTAIL.n148 11.249
R177 VTAIL.n176 VTAIL.n175 11.249
R178 VTAIL.n135 VTAIL.n76 11.249
R179 VTAIL.n104 VTAIL.n103 11.249
R180 VTAIL.n251 VTAIL.n234 10.4732
R181 VTAIL.n276 VTAIL.n275 10.4732
R182 VTAIL.n35 VTAIL.n18 10.4732
R183 VTAIL.n60 VTAIL.n59 10.4732
R184 VTAIL.n204 VTAIL.n203 10.4732
R185 VTAIL.n179 VTAIL.n162 10.4732
R186 VTAIL.n132 VTAIL.n131 10.4732
R187 VTAIL.n107 VTAIL.n90 10.4732
R188 VTAIL.n252 VTAIL.n232 9.69747
R189 VTAIL.n272 VTAIL.n222 9.69747
R190 VTAIL.n36 VTAIL.n16 9.69747
R191 VTAIL.n56 VTAIL.n6 9.69747
R192 VTAIL.n200 VTAIL.n150 9.69747
R193 VTAIL.n180 VTAIL.n160 9.69747
R194 VTAIL.n128 VTAIL.n78 9.69747
R195 VTAIL.n108 VTAIL.n88 9.69747
R196 VTAIL.n286 VTAIL.n285 9.45567
R197 VTAIL.n70 VTAIL.n69 9.45567
R198 VTAIL.n214 VTAIL.n213 9.45567
R199 VTAIL.n142 VTAIL.n141 9.45567
R200 VTAIL.n261 VTAIL.n260 9.3005
R201 VTAIL.n230 VTAIL.n229 9.3005
R202 VTAIL.n255 VTAIL.n254 9.3005
R203 VTAIL.n253 VTAIL.n252 9.3005
R204 VTAIL.n234 VTAIL.n233 9.3005
R205 VTAIL.n247 VTAIL.n246 9.3005
R206 VTAIL.n245 VTAIL.n244 9.3005
R207 VTAIL.n238 VTAIL.n237 9.3005
R208 VTAIL.n263 VTAIL.n262 9.3005
R209 VTAIL.n226 VTAIL.n225 9.3005
R210 VTAIL.n269 VTAIL.n268 9.3005
R211 VTAIL.n271 VTAIL.n270 9.3005
R212 VTAIL.n222 VTAIL.n221 9.3005
R213 VTAIL.n277 VTAIL.n276 9.3005
R214 VTAIL.n279 VTAIL.n278 9.3005
R215 VTAIL.n218 VTAIL.n217 9.3005
R216 VTAIL.n285 VTAIL.n284 9.3005
R217 VTAIL.n45 VTAIL.n44 9.3005
R218 VTAIL.n14 VTAIL.n13 9.3005
R219 VTAIL.n39 VTAIL.n38 9.3005
R220 VTAIL.n37 VTAIL.n36 9.3005
R221 VTAIL.n18 VTAIL.n17 9.3005
R222 VTAIL.n31 VTAIL.n30 9.3005
R223 VTAIL.n29 VTAIL.n28 9.3005
R224 VTAIL.n22 VTAIL.n21 9.3005
R225 VTAIL.n47 VTAIL.n46 9.3005
R226 VTAIL.n10 VTAIL.n9 9.3005
R227 VTAIL.n53 VTAIL.n52 9.3005
R228 VTAIL.n55 VTAIL.n54 9.3005
R229 VTAIL.n6 VTAIL.n5 9.3005
R230 VTAIL.n61 VTAIL.n60 9.3005
R231 VTAIL.n63 VTAIL.n62 9.3005
R232 VTAIL.n2 VTAIL.n1 9.3005
R233 VTAIL.n69 VTAIL.n68 9.3005
R234 VTAIL.n154 VTAIL.n153 9.3005
R235 VTAIL.n197 VTAIL.n196 9.3005
R236 VTAIL.n199 VTAIL.n198 9.3005
R237 VTAIL.n150 VTAIL.n149 9.3005
R238 VTAIL.n205 VTAIL.n204 9.3005
R239 VTAIL.n207 VTAIL.n206 9.3005
R240 VTAIL.n146 VTAIL.n145 9.3005
R241 VTAIL.n213 VTAIL.n212 9.3005
R242 VTAIL.n191 VTAIL.n190 9.3005
R243 VTAIL.n189 VTAIL.n188 9.3005
R244 VTAIL.n158 VTAIL.n157 9.3005
R245 VTAIL.n183 VTAIL.n182 9.3005
R246 VTAIL.n181 VTAIL.n180 9.3005
R247 VTAIL.n162 VTAIL.n161 9.3005
R248 VTAIL.n175 VTAIL.n174 9.3005
R249 VTAIL.n173 VTAIL.n172 9.3005
R250 VTAIL.n166 VTAIL.n165 9.3005
R251 VTAIL.n82 VTAIL.n81 9.3005
R252 VTAIL.n125 VTAIL.n124 9.3005
R253 VTAIL.n127 VTAIL.n126 9.3005
R254 VTAIL.n78 VTAIL.n77 9.3005
R255 VTAIL.n133 VTAIL.n132 9.3005
R256 VTAIL.n135 VTAIL.n134 9.3005
R257 VTAIL.n74 VTAIL.n73 9.3005
R258 VTAIL.n141 VTAIL.n140 9.3005
R259 VTAIL.n119 VTAIL.n118 9.3005
R260 VTAIL.n117 VTAIL.n116 9.3005
R261 VTAIL.n86 VTAIL.n85 9.3005
R262 VTAIL.n111 VTAIL.n110 9.3005
R263 VTAIL.n109 VTAIL.n108 9.3005
R264 VTAIL.n90 VTAIL.n89 9.3005
R265 VTAIL.n103 VTAIL.n102 9.3005
R266 VTAIL.n101 VTAIL.n100 9.3005
R267 VTAIL.n94 VTAIL.n93 9.3005
R268 VTAIL.n256 VTAIL.n255 8.92171
R269 VTAIL.n271 VTAIL.n224 8.92171
R270 VTAIL.n40 VTAIL.n39 8.92171
R271 VTAIL.n55 VTAIL.n8 8.92171
R272 VTAIL.n199 VTAIL.n152 8.92171
R273 VTAIL.n184 VTAIL.n183 8.92171
R274 VTAIL.n127 VTAIL.n80 8.92171
R275 VTAIL.n112 VTAIL.n111 8.92171
R276 VTAIL.n286 VTAIL.n216 8.2187
R277 VTAIL.n70 VTAIL.n0 8.2187
R278 VTAIL.n214 VTAIL.n144 8.2187
R279 VTAIL.n142 VTAIL.n72 8.2187
R280 VTAIL.n259 VTAIL.n230 8.14595
R281 VTAIL.n268 VTAIL.n267 8.14595
R282 VTAIL.n43 VTAIL.n14 8.14595
R283 VTAIL.n52 VTAIL.n51 8.14595
R284 VTAIL.n196 VTAIL.n195 8.14595
R285 VTAIL.n187 VTAIL.n158 8.14595
R286 VTAIL.n124 VTAIL.n123 8.14595
R287 VTAIL.n115 VTAIL.n86 8.14595
R288 VTAIL.n260 VTAIL.n228 7.3702
R289 VTAIL.n264 VTAIL.n226 7.3702
R290 VTAIL.n44 VTAIL.n12 7.3702
R291 VTAIL.n48 VTAIL.n10 7.3702
R292 VTAIL.n192 VTAIL.n154 7.3702
R293 VTAIL.n188 VTAIL.n156 7.3702
R294 VTAIL.n120 VTAIL.n82 7.3702
R295 VTAIL.n116 VTAIL.n84 7.3702
R296 VTAIL.n263 VTAIL.n228 6.59444
R297 VTAIL.n264 VTAIL.n263 6.59444
R298 VTAIL.n47 VTAIL.n12 6.59444
R299 VTAIL.n48 VTAIL.n47 6.59444
R300 VTAIL.n192 VTAIL.n191 6.59444
R301 VTAIL.n191 VTAIL.n156 6.59444
R302 VTAIL.n120 VTAIL.n119 6.59444
R303 VTAIL.n119 VTAIL.n84 6.59444
R304 VTAIL.n260 VTAIL.n259 5.81868
R305 VTAIL.n267 VTAIL.n226 5.81868
R306 VTAIL.n44 VTAIL.n43 5.81868
R307 VTAIL.n51 VTAIL.n10 5.81868
R308 VTAIL.n195 VTAIL.n154 5.81868
R309 VTAIL.n188 VTAIL.n187 5.81868
R310 VTAIL.n123 VTAIL.n82 5.81868
R311 VTAIL.n116 VTAIL.n115 5.81868
R312 VTAIL.n284 VTAIL.n216 5.3904
R313 VTAIL.n68 VTAIL.n0 5.3904
R314 VTAIL.n212 VTAIL.n144 5.3904
R315 VTAIL.n140 VTAIL.n72 5.3904
R316 VTAIL.n256 VTAIL.n230 5.04292
R317 VTAIL.n268 VTAIL.n224 5.04292
R318 VTAIL.n40 VTAIL.n14 5.04292
R319 VTAIL.n52 VTAIL.n8 5.04292
R320 VTAIL.n196 VTAIL.n152 5.04292
R321 VTAIL.n184 VTAIL.n158 5.04292
R322 VTAIL.n124 VTAIL.n80 5.04292
R323 VTAIL.n112 VTAIL.n86 5.04292
R324 VTAIL.n239 VTAIL.n237 4.38563
R325 VTAIL.n23 VTAIL.n21 4.38563
R326 VTAIL.n167 VTAIL.n165 4.38563
R327 VTAIL.n95 VTAIL.n93 4.38563
R328 VTAIL.n255 VTAIL.n232 4.26717
R329 VTAIL.n272 VTAIL.n271 4.26717
R330 VTAIL.n39 VTAIL.n16 4.26717
R331 VTAIL.n56 VTAIL.n55 4.26717
R332 VTAIL.n200 VTAIL.n199 4.26717
R333 VTAIL.n183 VTAIL.n160 4.26717
R334 VTAIL.n128 VTAIL.n127 4.26717
R335 VTAIL.n111 VTAIL.n88 4.26717
R336 VTAIL.n252 VTAIL.n251 3.49141
R337 VTAIL.n275 VTAIL.n222 3.49141
R338 VTAIL.n36 VTAIL.n35 3.49141
R339 VTAIL.n59 VTAIL.n6 3.49141
R340 VTAIL.n203 VTAIL.n150 3.49141
R341 VTAIL.n180 VTAIL.n179 3.49141
R342 VTAIL.n131 VTAIL.n78 3.49141
R343 VTAIL.n108 VTAIL.n107 3.49141
R344 VTAIL.n248 VTAIL.n234 2.71565
R345 VTAIL.n276 VTAIL.n220 2.71565
R346 VTAIL.n32 VTAIL.n18 2.71565
R347 VTAIL.n60 VTAIL.n4 2.71565
R348 VTAIL.n204 VTAIL.n148 2.71565
R349 VTAIL.n176 VTAIL.n162 2.71565
R350 VTAIL.n132 VTAIL.n76 2.71565
R351 VTAIL.n104 VTAIL.n90 2.71565
R352 VTAIL.n247 VTAIL.n236 1.93989
R353 VTAIL.n280 VTAIL.n279 1.93989
R354 VTAIL.n31 VTAIL.n20 1.93989
R355 VTAIL.n64 VTAIL.n63 1.93989
R356 VTAIL.n208 VTAIL.n207 1.93989
R357 VTAIL.n175 VTAIL.n164 1.93989
R358 VTAIL.n136 VTAIL.n135 1.93989
R359 VTAIL.n103 VTAIL.n92 1.93989
R360 VTAIL.n244 VTAIL.n243 1.16414
R361 VTAIL.n283 VTAIL.n218 1.16414
R362 VTAIL.n28 VTAIL.n27 1.16414
R363 VTAIL.n67 VTAIL.n2 1.16414
R364 VTAIL.n211 VTAIL.n146 1.16414
R365 VTAIL.n172 VTAIL.n171 1.16414
R366 VTAIL.n139 VTAIL.n74 1.16414
R367 VTAIL.n100 VTAIL.n99 1.16414
R368 VTAIL.n215 VTAIL.n143 0.901362
R369 VTAIL VTAIL.n71 0.744035
R370 VTAIL.n240 VTAIL.n238 0.388379
R371 VTAIL.n24 VTAIL.n22 0.388379
R372 VTAIL.n168 VTAIL.n166 0.388379
R373 VTAIL.n96 VTAIL.n94 0.388379
R374 VTAIL VTAIL.n287 0.157828
R375 VTAIL.n245 VTAIL.n237 0.155672
R376 VTAIL.n246 VTAIL.n245 0.155672
R377 VTAIL.n246 VTAIL.n233 0.155672
R378 VTAIL.n253 VTAIL.n233 0.155672
R379 VTAIL.n254 VTAIL.n253 0.155672
R380 VTAIL.n254 VTAIL.n229 0.155672
R381 VTAIL.n261 VTAIL.n229 0.155672
R382 VTAIL.n262 VTAIL.n261 0.155672
R383 VTAIL.n262 VTAIL.n225 0.155672
R384 VTAIL.n269 VTAIL.n225 0.155672
R385 VTAIL.n270 VTAIL.n269 0.155672
R386 VTAIL.n270 VTAIL.n221 0.155672
R387 VTAIL.n277 VTAIL.n221 0.155672
R388 VTAIL.n278 VTAIL.n277 0.155672
R389 VTAIL.n278 VTAIL.n217 0.155672
R390 VTAIL.n285 VTAIL.n217 0.155672
R391 VTAIL.n29 VTAIL.n21 0.155672
R392 VTAIL.n30 VTAIL.n29 0.155672
R393 VTAIL.n30 VTAIL.n17 0.155672
R394 VTAIL.n37 VTAIL.n17 0.155672
R395 VTAIL.n38 VTAIL.n37 0.155672
R396 VTAIL.n38 VTAIL.n13 0.155672
R397 VTAIL.n45 VTAIL.n13 0.155672
R398 VTAIL.n46 VTAIL.n45 0.155672
R399 VTAIL.n46 VTAIL.n9 0.155672
R400 VTAIL.n53 VTAIL.n9 0.155672
R401 VTAIL.n54 VTAIL.n53 0.155672
R402 VTAIL.n54 VTAIL.n5 0.155672
R403 VTAIL.n61 VTAIL.n5 0.155672
R404 VTAIL.n62 VTAIL.n61 0.155672
R405 VTAIL.n62 VTAIL.n1 0.155672
R406 VTAIL.n69 VTAIL.n1 0.155672
R407 VTAIL.n213 VTAIL.n145 0.155672
R408 VTAIL.n206 VTAIL.n145 0.155672
R409 VTAIL.n206 VTAIL.n205 0.155672
R410 VTAIL.n205 VTAIL.n149 0.155672
R411 VTAIL.n198 VTAIL.n149 0.155672
R412 VTAIL.n198 VTAIL.n197 0.155672
R413 VTAIL.n197 VTAIL.n153 0.155672
R414 VTAIL.n190 VTAIL.n153 0.155672
R415 VTAIL.n190 VTAIL.n189 0.155672
R416 VTAIL.n189 VTAIL.n157 0.155672
R417 VTAIL.n182 VTAIL.n157 0.155672
R418 VTAIL.n182 VTAIL.n181 0.155672
R419 VTAIL.n181 VTAIL.n161 0.155672
R420 VTAIL.n174 VTAIL.n161 0.155672
R421 VTAIL.n174 VTAIL.n173 0.155672
R422 VTAIL.n173 VTAIL.n165 0.155672
R423 VTAIL.n141 VTAIL.n73 0.155672
R424 VTAIL.n134 VTAIL.n73 0.155672
R425 VTAIL.n134 VTAIL.n133 0.155672
R426 VTAIL.n133 VTAIL.n77 0.155672
R427 VTAIL.n126 VTAIL.n77 0.155672
R428 VTAIL.n126 VTAIL.n125 0.155672
R429 VTAIL.n125 VTAIL.n81 0.155672
R430 VTAIL.n118 VTAIL.n81 0.155672
R431 VTAIL.n118 VTAIL.n117 0.155672
R432 VTAIL.n117 VTAIL.n85 0.155672
R433 VTAIL.n110 VTAIL.n85 0.155672
R434 VTAIL.n110 VTAIL.n109 0.155672
R435 VTAIL.n109 VTAIL.n89 0.155672
R436 VTAIL.n102 VTAIL.n89 0.155672
R437 VTAIL.n102 VTAIL.n101 0.155672
R438 VTAIL.n101 VTAIL.n93 0.155672
R439 VDD2.n137 VDD2.n71 214.453
R440 VDD2.n66 VDD2.n0 214.453
R441 VDD2.n138 VDD2.n137 185
R442 VDD2.n136 VDD2.n135 185
R443 VDD2.n75 VDD2.n74 185
R444 VDD2.n130 VDD2.n129 185
R445 VDD2.n128 VDD2.n127 185
R446 VDD2.n79 VDD2.n78 185
R447 VDD2.n122 VDD2.n121 185
R448 VDD2.n120 VDD2.n119 185
R449 VDD2.n83 VDD2.n82 185
R450 VDD2.n114 VDD2.n113 185
R451 VDD2.n112 VDD2.n111 185
R452 VDD2.n87 VDD2.n86 185
R453 VDD2.n106 VDD2.n105 185
R454 VDD2.n104 VDD2.n103 185
R455 VDD2.n91 VDD2.n90 185
R456 VDD2.n98 VDD2.n97 185
R457 VDD2.n96 VDD2.n95 185
R458 VDD2.n25 VDD2.n24 185
R459 VDD2.n27 VDD2.n26 185
R460 VDD2.n20 VDD2.n19 185
R461 VDD2.n33 VDD2.n32 185
R462 VDD2.n35 VDD2.n34 185
R463 VDD2.n16 VDD2.n15 185
R464 VDD2.n41 VDD2.n40 185
R465 VDD2.n43 VDD2.n42 185
R466 VDD2.n12 VDD2.n11 185
R467 VDD2.n49 VDD2.n48 185
R468 VDD2.n51 VDD2.n50 185
R469 VDD2.n8 VDD2.n7 185
R470 VDD2.n57 VDD2.n56 185
R471 VDD2.n59 VDD2.n58 185
R472 VDD2.n4 VDD2.n3 185
R473 VDD2.n65 VDD2.n64 185
R474 VDD2.n67 VDD2.n66 185
R475 VDD2.n23 VDD2.t0 147.659
R476 VDD2.n94 VDD2.t1 147.659
R477 VDD2.n137 VDD2.n136 104.615
R478 VDD2.n136 VDD2.n74 104.615
R479 VDD2.n129 VDD2.n74 104.615
R480 VDD2.n129 VDD2.n128 104.615
R481 VDD2.n128 VDD2.n78 104.615
R482 VDD2.n121 VDD2.n78 104.615
R483 VDD2.n121 VDD2.n120 104.615
R484 VDD2.n120 VDD2.n82 104.615
R485 VDD2.n113 VDD2.n82 104.615
R486 VDD2.n113 VDD2.n112 104.615
R487 VDD2.n112 VDD2.n86 104.615
R488 VDD2.n105 VDD2.n86 104.615
R489 VDD2.n105 VDD2.n104 104.615
R490 VDD2.n104 VDD2.n90 104.615
R491 VDD2.n97 VDD2.n90 104.615
R492 VDD2.n97 VDD2.n96 104.615
R493 VDD2.n26 VDD2.n25 104.615
R494 VDD2.n26 VDD2.n19 104.615
R495 VDD2.n33 VDD2.n19 104.615
R496 VDD2.n34 VDD2.n33 104.615
R497 VDD2.n34 VDD2.n15 104.615
R498 VDD2.n41 VDD2.n15 104.615
R499 VDD2.n42 VDD2.n41 104.615
R500 VDD2.n42 VDD2.n11 104.615
R501 VDD2.n49 VDD2.n11 104.615
R502 VDD2.n50 VDD2.n49 104.615
R503 VDD2.n50 VDD2.n7 104.615
R504 VDD2.n57 VDD2.n7 104.615
R505 VDD2.n58 VDD2.n57 104.615
R506 VDD2.n58 VDD2.n3 104.615
R507 VDD2.n65 VDD2.n3 104.615
R508 VDD2.n66 VDD2.n65 104.615
R509 VDD2.n142 VDD2.n70 89.2904
R510 VDD2.n142 VDD2.n141 52.355
R511 VDD2.n96 VDD2.t1 52.3082
R512 VDD2.n25 VDD2.t0 52.3082
R513 VDD2.n95 VDD2.n94 15.6677
R514 VDD2.n24 VDD2.n23 15.6677
R515 VDD2.n139 VDD2.n138 12.8005
R516 VDD2.n98 VDD2.n93 12.8005
R517 VDD2.n27 VDD2.n22 12.8005
R518 VDD2.n68 VDD2.n67 12.8005
R519 VDD2.n135 VDD2.n73 12.0247
R520 VDD2.n99 VDD2.n91 12.0247
R521 VDD2.n28 VDD2.n20 12.0247
R522 VDD2.n64 VDD2.n2 12.0247
R523 VDD2.n134 VDD2.n75 11.249
R524 VDD2.n103 VDD2.n102 11.249
R525 VDD2.n32 VDD2.n31 11.249
R526 VDD2.n63 VDD2.n4 11.249
R527 VDD2.n131 VDD2.n130 10.4732
R528 VDD2.n106 VDD2.n89 10.4732
R529 VDD2.n35 VDD2.n18 10.4732
R530 VDD2.n60 VDD2.n59 10.4732
R531 VDD2.n127 VDD2.n77 9.69747
R532 VDD2.n107 VDD2.n87 9.69747
R533 VDD2.n36 VDD2.n16 9.69747
R534 VDD2.n56 VDD2.n6 9.69747
R535 VDD2.n141 VDD2.n140 9.45567
R536 VDD2.n70 VDD2.n69 9.45567
R537 VDD2.n81 VDD2.n80 9.3005
R538 VDD2.n124 VDD2.n123 9.3005
R539 VDD2.n126 VDD2.n125 9.3005
R540 VDD2.n77 VDD2.n76 9.3005
R541 VDD2.n132 VDD2.n131 9.3005
R542 VDD2.n134 VDD2.n133 9.3005
R543 VDD2.n73 VDD2.n72 9.3005
R544 VDD2.n140 VDD2.n139 9.3005
R545 VDD2.n118 VDD2.n117 9.3005
R546 VDD2.n116 VDD2.n115 9.3005
R547 VDD2.n85 VDD2.n84 9.3005
R548 VDD2.n110 VDD2.n109 9.3005
R549 VDD2.n108 VDD2.n107 9.3005
R550 VDD2.n89 VDD2.n88 9.3005
R551 VDD2.n102 VDD2.n101 9.3005
R552 VDD2.n100 VDD2.n99 9.3005
R553 VDD2.n93 VDD2.n92 9.3005
R554 VDD2.n45 VDD2.n44 9.3005
R555 VDD2.n14 VDD2.n13 9.3005
R556 VDD2.n39 VDD2.n38 9.3005
R557 VDD2.n37 VDD2.n36 9.3005
R558 VDD2.n18 VDD2.n17 9.3005
R559 VDD2.n31 VDD2.n30 9.3005
R560 VDD2.n29 VDD2.n28 9.3005
R561 VDD2.n22 VDD2.n21 9.3005
R562 VDD2.n47 VDD2.n46 9.3005
R563 VDD2.n10 VDD2.n9 9.3005
R564 VDD2.n53 VDD2.n52 9.3005
R565 VDD2.n55 VDD2.n54 9.3005
R566 VDD2.n6 VDD2.n5 9.3005
R567 VDD2.n61 VDD2.n60 9.3005
R568 VDD2.n63 VDD2.n62 9.3005
R569 VDD2.n2 VDD2.n1 9.3005
R570 VDD2.n69 VDD2.n68 9.3005
R571 VDD2.n126 VDD2.n79 8.92171
R572 VDD2.n111 VDD2.n110 8.92171
R573 VDD2.n40 VDD2.n39 8.92171
R574 VDD2.n55 VDD2.n8 8.92171
R575 VDD2.n141 VDD2.n71 8.2187
R576 VDD2.n70 VDD2.n0 8.2187
R577 VDD2.n123 VDD2.n122 8.14595
R578 VDD2.n114 VDD2.n85 8.14595
R579 VDD2.n43 VDD2.n14 8.14595
R580 VDD2.n52 VDD2.n51 8.14595
R581 VDD2.n119 VDD2.n81 7.3702
R582 VDD2.n115 VDD2.n83 7.3702
R583 VDD2.n44 VDD2.n12 7.3702
R584 VDD2.n48 VDD2.n10 7.3702
R585 VDD2.n119 VDD2.n118 6.59444
R586 VDD2.n118 VDD2.n83 6.59444
R587 VDD2.n47 VDD2.n12 6.59444
R588 VDD2.n48 VDD2.n47 6.59444
R589 VDD2.n122 VDD2.n81 5.81868
R590 VDD2.n115 VDD2.n114 5.81868
R591 VDD2.n44 VDD2.n43 5.81868
R592 VDD2.n51 VDD2.n10 5.81868
R593 VDD2.n139 VDD2.n71 5.3904
R594 VDD2.n68 VDD2.n0 5.3904
R595 VDD2.n123 VDD2.n79 5.04292
R596 VDD2.n111 VDD2.n85 5.04292
R597 VDD2.n40 VDD2.n14 5.04292
R598 VDD2.n52 VDD2.n8 5.04292
R599 VDD2.n23 VDD2.n21 4.38563
R600 VDD2.n94 VDD2.n92 4.38563
R601 VDD2.n127 VDD2.n126 4.26717
R602 VDD2.n110 VDD2.n87 4.26717
R603 VDD2.n39 VDD2.n16 4.26717
R604 VDD2.n56 VDD2.n55 4.26717
R605 VDD2.n130 VDD2.n77 3.49141
R606 VDD2.n107 VDD2.n106 3.49141
R607 VDD2.n36 VDD2.n35 3.49141
R608 VDD2.n59 VDD2.n6 3.49141
R609 VDD2.n131 VDD2.n75 2.71565
R610 VDD2.n103 VDD2.n89 2.71565
R611 VDD2.n32 VDD2.n18 2.71565
R612 VDD2.n60 VDD2.n4 2.71565
R613 VDD2.n135 VDD2.n134 1.93989
R614 VDD2.n102 VDD2.n91 1.93989
R615 VDD2.n31 VDD2.n20 1.93989
R616 VDD2.n64 VDD2.n63 1.93989
R617 VDD2.n138 VDD2.n73 1.16414
R618 VDD2.n99 VDD2.n98 1.16414
R619 VDD2.n28 VDD2.n27 1.16414
R620 VDD2.n67 VDD2.n2 1.16414
R621 VDD2.n95 VDD2.n93 0.388379
R622 VDD2.n24 VDD2.n22 0.388379
R623 VDD2 VDD2.n142 0.274207
R624 VDD2.n140 VDD2.n72 0.155672
R625 VDD2.n133 VDD2.n72 0.155672
R626 VDD2.n133 VDD2.n132 0.155672
R627 VDD2.n132 VDD2.n76 0.155672
R628 VDD2.n125 VDD2.n76 0.155672
R629 VDD2.n125 VDD2.n124 0.155672
R630 VDD2.n124 VDD2.n80 0.155672
R631 VDD2.n117 VDD2.n80 0.155672
R632 VDD2.n117 VDD2.n116 0.155672
R633 VDD2.n116 VDD2.n84 0.155672
R634 VDD2.n109 VDD2.n84 0.155672
R635 VDD2.n109 VDD2.n108 0.155672
R636 VDD2.n108 VDD2.n88 0.155672
R637 VDD2.n101 VDD2.n88 0.155672
R638 VDD2.n101 VDD2.n100 0.155672
R639 VDD2.n100 VDD2.n92 0.155672
R640 VDD2.n29 VDD2.n21 0.155672
R641 VDD2.n30 VDD2.n29 0.155672
R642 VDD2.n30 VDD2.n17 0.155672
R643 VDD2.n37 VDD2.n17 0.155672
R644 VDD2.n38 VDD2.n37 0.155672
R645 VDD2.n38 VDD2.n13 0.155672
R646 VDD2.n45 VDD2.n13 0.155672
R647 VDD2.n46 VDD2.n45 0.155672
R648 VDD2.n46 VDD2.n9 0.155672
R649 VDD2.n53 VDD2.n9 0.155672
R650 VDD2.n54 VDD2.n53 0.155672
R651 VDD2.n54 VDD2.n5 0.155672
R652 VDD2.n61 VDD2.n5 0.155672
R653 VDD2.n62 VDD2.n61 0.155672
R654 VDD2.n62 VDD2.n1 0.155672
R655 VDD2.n69 VDD2.n1 0.155672
R656 B.n144 B.t13 684.631
R657 B.n137 B.t2 684.631
R658 B.n53 B.t10 684.631
R659 B.n61 B.t6 684.631
R660 B.n430 B.n429 585
R661 B.n430 B.n29 585
R662 B.n433 B.n432 585
R663 B.n434 B.n84 585
R664 B.n436 B.n435 585
R665 B.n438 B.n83 585
R666 B.n441 B.n440 585
R667 B.n442 B.n82 585
R668 B.n444 B.n443 585
R669 B.n446 B.n81 585
R670 B.n449 B.n448 585
R671 B.n450 B.n80 585
R672 B.n452 B.n451 585
R673 B.n454 B.n79 585
R674 B.n457 B.n456 585
R675 B.n458 B.n78 585
R676 B.n460 B.n459 585
R677 B.n462 B.n77 585
R678 B.n465 B.n464 585
R679 B.n466 B.n76 585
R680 B.n468 B.n467 585
R681 B.n470 B.n75 585
R682 B.n473 B.n472 585
R683 B.n474 B.n74 585
R684 B.n476 B.n475 585
R685 B.n478 B.n73 585
R686 B.n481 B.n480 585
R687 B.n482 B.n72 585
R688 B.n484 B.n483 585
R689 B.n486 B.n71 585
R690 B.n489 B.n488 585
R691 B.n490 B.n70 585
R692 B.n492 B.n491 585
R693 B.n494 B.n69 585
R694 B.n497 B.n496 585
R695 B.n498 B.n68 585
R696 B.n500 B.n499 585
R697 B.n502 B.n67 585
R698 B.n505 B.n504 585
R699 B.n506 B.n66 585
R700 B.n508 B.n507 585
R701 B.n510 B.n65 585
R702 B.n513 B.n512 585
R703 B.n514 B.n64 585
R704 B.n516 B.n515 585
R705 B.n518 B.n63 585
R706 B.n521 B.n520 585
R707 B.n523 B.n60 585
R708 B.n525 B.n524 585
R709 B.n527 B.n59 585
R710 B.n530 B.n529 585
R711 B.n531 B.n58 585
R712 B.n533 B.n532 585
R713 B.n535 B.n57 585
R714 B.n537 B.n536 585
R715 B.n539 B.n538 585
R716 B.n542 B.n541 585
R717 B.n543 B.n52 585
R718 B.n545 B.n544 585
R719 B.n547 B.n51 585
R720 B.n550 B.n549 585
R721 B.n551 B.n50 585
R722 B.n553 B.n552 585
R723 B.n555 B.n49 585
R724 B.n558 B.n557 585
R725 B.n559 B.n48 585
R726 B.n561 B.n560 585
R727 B.n563 B.n47 585
R728 B.n566 B.n565 585
R729 B.n567 B.n46 585
R730 B.n569 B.n568 585
R731 B.n571 B.n45 585
R732 B.n574 B.n573 585
R733 B.n575 B.n44 585
R734 B.n577 B.n576 585
R735 B.n579 B.n43 585
R736 B.n582 B.n581 585
R737 B.n583 B.n42 585
R738 B.n585 B.n584 585
R739 B.n587 B.n41 585
R740 B.n590 B.n589 585
R741 B.n591 B.n40 585
R742 B.n593 B.n592 585
R743 B.n595 B.n39 585
R744 B.n598 B.n597 585
R745 B.n599 B.n38 585
R746 B.n601 B.n600 585
R747 B.n603 B.n37 585
R748 B.n606 B.n605 585
R749 B.n607 B.n36 585
R750 B.n609 B.n608 585
R751 B.n611 B.n35 585
R752 B.n614 B.n613 585
R753 B.n615 B.n34 585
R754 B.n617 B.n616 585
R755 B.n619 B.n33 585
R756 B.n622 B.n621 585
R757 B.n623 B.n32 585
R758 B.n625 B.n624 585
R759 B.n627 B.n31 585
R760 B.n630 B.n629 585
R761 B.n631 B.n30 585
R762 B.n428 B.n28 585
R763 B.n634 B.n28 585
R764 B.n427 B.n27 585
R765 B.n635 B.n27 585
R766 B.n426 B.n26 585
R767 B.n636 B.n26 585
R768 B.n425 B.n424 585
R769 B.n424 B.n22 585
R770 B.n423 B.n21 585
R771 B.n642 B.n21 585
R772 B.n422 B.n20 585
R773 B.n643 B.n20 585
R774 B.n421 B.n19 585
R775 B.n644 B.n19 585
R776 B.n420 B.n419 585
R777 B.n419 B.n15 585
R778 B.n418 B.n14 585
R779 B.n650 B.n14 585
R780 B.n417 B.n13 585
R781 B.n651 B.n13 585
R782 B.n416 B.n12 585
R783 B.n652 B.n12 585
R784 B.n415 B.n414 585
R785 B.n414 B.n8 585
R786 B.n413 B.n7 585
R787 B.n658 B.n7 585
R788 B.n412 B.n6 585
R789 B.n659 B.n6 585
R790 B.n411 B.n5 585
R791 B.n660 B.n5 585
R792 B.n410 B.n409 585
R793 B.n409 B.n4 585
R794 B.n408 B.n85 585
R795 B.n408 B.n407 585
R796 B.n398 B.n86 585
R797 B.n87 B.n86 585
R798 B.n400 B.n399 585
R799 B.n401 B.n400 585
R800 B.n397 B.n92 585
R801 B.n92 B.n91 585
R802 B.n396 B.n395 585
R803 B.n395 B.n394 585
R804 B.n94 B.n93 585
R805 B.n95 B.n94 585
R806 B.n387 B.n386 585
R807 B.n388 B.n387 585
R808 B.n385 B.n100 585
R809 B.n100 B.n99 585
R810 B.n384 B.n383 585
R811 B.n383 B.n382 585
R812 B.n102 B.n101 585
R813 B.n103 B.n102 585
R814 B.n375 B.n374 585
R815 B.n376 B.n375 585
R816 B.n373 B.n108 585
R817 B.n108 B.n107 585
R818 B.n372 B.n371 585
R819 B.n371 B.n370 585
R820 B.n367 B.n112 585
R821 B.n366 B.n365 585
R822 B.n363 B.n113 585
R823 B.n363 B.n111 585
R824 B.n362 B.n361 585
R825 B.n360 B.n359 585
R826 B.n358 B.n115 585
R827 B.n356 B.n355 585
R828 B.n354 B.n116 585
R829 B.n353 B.n352 585
R830 B.n350 B.n117 585
R831 B.n348 B.n347 585
R832 B.n346 B.n118 585
R833 B.n345 B.n344 585
R834 B.n342 B.n119 585
R835 B.n340 B.n339 585
R836 B.n338 B.n120 585
R837 B.n337 B.n336 585
R838 B.n334 B.n121 585
R839 B.n332 B.n331 585
R840 B.n330 B.n122 585
R841 B.n329 B.n328 585
R842 B.n326 B.n123 585
R843 B.n324 B.n323 585
R844 B.n322 B.n124 585
R845 B.n321 B.n320 585
R846 B.n318 B.n125 585
R847 B.n316 B.n315 585
R848 B.n314 B.n126 585
R849 B.n313 B.n312 585
R850 B.n310 B.n127 585
R851 B.n308 B.n307 585
R852 B.n306 B.n128 585
R853 B.n305 B.n304 585
R854 B.n302 B.n129 585
R855 B.n300 B.n299 585
R856 B.n298 B.n130 585
R857 B.n297 B.n296 585
R858 B.n294 B.n131 585
R859 B.n292 B.n291 585
R860 B.n290 B.n132 585
R861 B.n289 B.n288 585
R862 B.n286 B.n133 585
R863 B.n284 B.n283 585
R864 B.n282 B.n134 585
R865 B.n281 B.n280 585
R866 B.n278 B.n135 585
R867 B.n276 B.n275 585
R868 B.n274 B.n136 585
R869 B.n273 B.n272 585
R870 B.n270 B.n140 585
R871 B.n268 B.n267 585
R872 B.n266 B.n141 585
R873 B.n265 B.n264 585
R874 B.n262 B.n142 585
R875 B.n260 B.n259 585
R876 B.n257 B.n143 585
R877 B.n256 B.n255 585
R878 B.n253 B.n146 585
R879 B.n251 B.n250 585
R880 B.n249 B.n147 585
R881 B.n248 B.n247 585
R882 B.n245 B.n148 585
R883 B.n243 B.n242 585
R884 B.n241 B.n149 585
R885 B.n240 B.n239 585
R886 B.n237 B.n150 585
R887 B.n235 B.n234 585
R888 B.n233 B.n151 585
R889 B.n232 B.n231 585
R890 B.n229 B.n152 585
R891 B.n227 B.n226 585
R892 B.n225 B.n153 585
R893 B.n224 B.n223 585
R894 B.n221 B.n154 585
R895 B.n219 B.n218 585
R896 B.n217 B.n155 585
R897 B.n216 B.n215 585
R898 B.n213 B.n156 585
R899 B.n211 B.n210 585
R900 B.n209 B.n157 585
R901 B.n208 B.n207 585
R902 B.n205 B.n158 585
R903 B.n203 B.n202 585
R904 B.n201 B.n159 585
R905 B.n200 B.n199 585
R906 B.n197 B.n160 585
R907 B.n195 B.n194 585
R908 B.n193 B.n161 585
R909 B.n192 B.n191 585
R910 B.n189 B.n162 585
R911 B.n187 B.n186 585
R912 B.n185 B.n163 585
R913 B.n184 B.n183 585
R914 B.n181 B.n164 585
R915 B.n179 B.n178 585
R916 B.n177 B.n165 585
R917 B.n176 B.n175 585
R918 B.n173 B.n166 585
R919 B.n171 B.n170 585
R920 B.n169 B.n168 585
R921 B.n110 B.n109 585
R922 B.n369 B.n368 585
R923 B.n370 B.n369 585
R924 B.n106 B.n105 585
R925 B.n107 B.n106 585
R926 B.n378 B.n377 585
R927 B.n377 B.n376 585
R928 B.n379 B.n104 585
R929 B.n104 B.n103 585
R930 B.n381 B.n380 585
R931 B.n382 B.n381 585
R932 B.n98 B.n97 585
R933 B.n99 B.n98 585
R934 B.n390 B.n389 585
R935 B.n389 B.n388 585
R936 B.n391 B.n96 585
R937 B.n96 B.n95 585
R938 B.n393 B.n392 585
R939 B.n394 B.n393 585
R940 B.n90 B.n89 585
R941 B.n91 B.n90 585
R942 B.n403 B.n402 585
R943 B.n402 B.n401 585
R944 B.n404 B.n88 585
R945 B.n88 B.n87 585
R946 B.n406 B.n405 585
R947 B.n407 B.n406 585
R948 B.n2 B.n0 585
R949 B.n4 B.n2 585
R950 B.n3 B.n1 585
R951 B.n659 B.n3 585
R952 B.n657 B.n656 585
R953 B.n658 B.n657 585
R954 B.n655 B.n9 585
R955 B.n9 B.n8 585
R956 B.n654 B.n653 585
R957 B.n653 B.n652 585
R958 B.n11 B.n10 585
R959 B.n651 B.n11 585
R960 B.n649 B.n648 585
R961 B.n650 B.n649 585
R962 B.n647 B.n16 585
R963 B.n16 B.n15 585
R964 B.n646 B.n645 585
R965 B.n645 B.n644 585
R966 B.n18 B.n17 585
R967 B.n643 B.n18 585
R968 B.n641 B.n640 585
R969 B.n642 B.n641 585
R970 B.n639 B.n23 585
R971 B.n23 B.n22 585
R972 B.n638 B.n637 585
R973 B.n637 B.n636 585
R974 B.n25 B.n24 585
R975 B.n635 B.n25 585
R976 B.n633 B.n632 585
R977 B.n634 B.n633 585
R978 B.n662 B.n661 585
R979 B.n661 B.n660 585
R980 B.n369 B.n112 502.111
R981 B.n633 B.n30 502.111
R982 B.n371 B.n110 502.111
R983 B.n430 B.n28 502.111
R984 B.n144 B.t15 325.214
R985 B.n61 B.t8 325.214
R986 B.n137 B.t5 325.214
R987 B.n53 B.t11 325.214
R988 B.n145 B.t14 305.82
R989 B.n62 B.t9 305.82
R990 B.n138 B.t4 305.82
R991 B.n54 B.t12 305.82
R992 B.n431 B.n29 256.663
R993 B.n437 B.n29 256.663
R994 B.n439 B.n29 256.663
R995 B.n445 B.n29 256.663
R996 B.n447 B.n29 256.663
R997 B.n453 B.n29 256.663
R998 B.n455 B.n29 256.663
R999 B.n461 B.n29 256.663
R1000 B.n463 B.n29 256.663
R1001 B.n469 B.n29 256.663
R1002 B.n471 B.n29 256.663
R1003 B.n477 B.n29 256.663
R1004 B.n479 B.n29 256.663
R1005 B.n485 B.n29 256.663
R1006 B.n487 B.n29 256.663
R1007 B.n493 B.n29 256.663
R1008 B.n495 B.n29 256.663
R1009 B.n501 B.n29 256.663
R1010 B.n503 B.n29 256.663
R1011 B.n509 B.n29 256.663
R1012 B.n511 B.n29 256.663
R1013 B.n517 B.n29 256.663
R1014 B.n519 B.n29 256.663
R1015 B.n526 B.n29 256.663
R1016 B.n528 B.n29 256.663
R1017 B.n534 B.n29 256.663
R1018 B.n56 B.n29 256.663
R1019 B.n540 B.n29 256.663
R1020 B.n546 B.n29 256.663
R1021 B.n548 B.n29 256.663
R1022 B.n554 B.n29 256.663
R1023 B.n556 B.n29 256.663
R1024 B.n562 B.n29 256.663
R1025 B.n564 B.n29 256.663
R1026 B.n570 B.n29 256.663
R1027 B.n572 B.n29 256.663
R1028 B.n578 B.n29 256.663
R1029 B.n580 B.n29 256.663
R1030 B.n586 B.n29 256.663
R1031 B.n588 B.n29 256.663
R1032 B.n594 B.n29 256.663
R1033 B.n596 B.n29 256.663
R1034 B.n602 B.n29 256.663
R1035 B.n604 B.n29 256.663
R1036 B.n610 B.n29 256.663
R1037 B.n612 B.n29 256.663
R1038 B.n618 B.n29 256.663
R1039 B.n620 B.n29 256.663
R1040 B.n626 B.n29 256.663
R1041 B.n628 B.n29 256.663
R1042 B.n364 B.n111 256.663
R1043 B.n114 B.n111 256.663
R1044 B.n357 B.n111 256.663
R1045 B.n351 B.n111 256.663
R1046 B.n349 B.n111 256.663
R1047 B.n343 B.n111 256.663
R1048 B.n341 B.n111 256.663
R1049 B.n335 B.n111 256.663
R1050 B.n333 B.n111 256.663
R1051 B.n327 B.n111 256.663
R1052 B.n325 B.n111 256.663
R1053 B.n319 B.n111 256.663
R1054 B.n317 B.n111 256.663
R1055 B.n311 B.n111 256.663
R1056 B.n309 B.n111 256.663
R1057 B.n303 B.n111 256.663
R1058 B.n301 B.n111 256.663
R1059 B.n295 B.n111 256.663
R1060 B.n293 B.n111 256.663
R1061 B.n287 B.n111 256.663
R1062 B.n285 B.n111 256.663
R1063 B.n279 B.n111 256.663
R1064 B.n277 B.n111 256.663
R1065 B.n271 B.n111 256.663
R1066 B.n269 B.n111 256.663
R1067 B.n263 B.n111 256.663
R1068 B.n261 B.n111 256.663
R1069 B.n254 B.n111 256.663
R1070 B.n252 B.n111 256.663
R1071 B.n246 B.n111 256.663
R1072 B.n244 B.n111 256.663
R1073 B.n238 B.n111 256.663
R1074 B.n236 B.n111 256.663
R1075 B.n230 B.n111 256.663
R1076 B.n228 B.n111 256.663
R1077 B.n222 B.n111 256.663
R1078 B.n220 B.n111 256.663
R1079 B.n214 B.n111 256.663
R1080 B.n212 B.n111 256.663
R1081 B.n206 B.n111 256.663
R1082 B.n204 B.n111 256.663
R1083 B.n198 B.n111 256.663
R1084 B.n196 B.n111 256.663
R1085 B.n190 B.n111 256.663
R1086 B.n188 B.n111 256.663
R1087 B.n182 B.n111 256.663
R1088 B.n180 B.n111 256.663
R1089 B.n174 B.n111 256.663
R1090 B.n172 B.n111 256.663
R1091 B.n167 B.n111 256.663
R1092 B.n369 B.n106 163.367
R1093 B.n377 B.n106 163.367
R1094 B.n377 B.n104 163.367
R1095 B.n381 B.n104 163.367
R1096 B.n381 B.n98 163.367
R1097 B.n389 B.n98 163.367
R1098 B.n389 B.n96 163.367
R1099 B.n393 B.n96 163.367
R1100 B.n393 B.n90 163.367
R1101 B.n402 B.n90 163.367
R1102 B.n402 B.n88 163.367
R1103 B.n406 B.n88 163.367
R1104 B.n406 B.n2 163.367
R1105 B.n661 B.n2 163.367
R1106 B.n661 B.n3 163.367
R1107 B.n657 B.n3 163.367
R1108 B.n657 B.n9 163.367
R1109 B.n653 B.n9 163.367
R1110 B.n653 B.n11 163.367
R1111 B.n649 B.n11 163.367
R1112 B.n649 B.n16 163.367
R1113 B.n645 B.n16 163.367
R1114 B.n645 B.n18 163.367
R1115 B.n641 B.n18 163.367
R1116 B.n641 B.n23 163.367
R1117 B.n637 B.n23 163.367
R1118 B.n637 B.n25 163.367
R1119 B.n633 B.n25 163.367
R1120 B.n365 B.n363 163.367
R1121 B.n363 B.n362 163.367
R1122 B.n359 B.n358 163.367
R1123 B.n356 B.n116 163.367
R1124 B.n352 B.n350 163.367
R1125 B.n348 B.n118 163.367
R1126 B.n344 B.n342 163.367
R1127 B.n340 B.n120 163.367
R1128 B.n336 B.n334 163.367
R1129 B.n332 B.n122 163.367
R1130 B.n328 B.n326 163.367
R1131 B.n324 B.n124 163.367
R1132 B.n320 B.n318 163.367
R1133 B.n316 B.n126 163.367
R1134 B.n312 B.n310 163.367
R1135 B.n308 B.n128 163.367
R1136 B.n304 B.n302 163.367
R1137 B.n300 B.n130 163.367
R1138 B.n296 B.n294 163.367
R1139 B.n292 B.n132 163.367
R1140 B.n288 B.n286 163.367
R1141 B.n284 B.n134 163.367
R1142 B.n280 B.n278 163.367
R1143 B.n276 B.n136 163.367
R1144 B.n272 B.n270 163.367
R1145 B.n268 B.n141 163.367
R1146 B.n264 B.n262 163.367
R1147 B.n260 B.n143 163.367
R1148 B.n255 B.n253 163.367
R1149 B.n251 B.n147 163.367
R1150 B.n247 B.n245 163.367
R1151 B.n243 B.n149 163.367
R1152 B.n239 B.n237 163.367
R1153 B.n235 B.n151 163.367
R1154 B.n231 B.n229 163.367
R1155 B.n227 B.n153 163.367
R1156 B.n223 B.n221 163.367
R1157 B.n219 B.n155 163.367
R1158 B.n215 B.n213 163.367
R1159 B.n211 B.n157 163.367
R1160 B.n207 B.n205 163.367
R1161 B.n203 B.n159 163.367
R1162 B.n199 B.n197 163.367
R1163 B.n195 B.n161 163.367
R1164 B.n191 B.n189 163.367
R1165 B.n187 B.n163 163.367
R1166 B.n183 B.n181 163.367
R1167 B.n179 B.n165 163.367
R1168 B.n175 B.n173 163.367
R1169 B.n171 B.n168 163.367
R1170 B.n371 B.n108 163.367
R1171 B.n375 B.n108 163.367
R1172 B.n375 B.n102 163.367
R1173 B.n383 B.n102 163.367
R1174 B.n383 B.n100 163.367
R1175 B.n387 B.n100 163.367
R1176 B.n387 B.n94 163.367
R1177 B.n395 B.n94 163.367
R1178 B.n395 B.n92 163.367
R1179 B.n400 B.n92 163.367
R1180 B.n400 B.n86 163.367
R1181 B.n408 B.n86 163.367
R1182 B.n409 B.n408 163.367
R1183 B.n409 B.n5 163.367
R1184 B.n6 B.n5 163.367
R1185 B.n7 B.n6 163.367
R1186 B.n414 B.n7 163.367
R1187 B.n414 B.n12 163.367
R1188 B.n13 B.n12 163.367
R1189 B.n14 B.n13 163.367
R1190 B.n419 B.n14 163.367
R1191 B.n419 B.n19 163.367
R1192 B.n20 B.n19 163.367
R1193 B.n21 B.n20 163.367
R1194 B.n424 B.n21 163.367
R1195 B.n424 B.n26 163.367
R1196 B.n27 B.n26 163.367
R1197 B.n28 B.n27 163.367
R1198 B.n629 B.n627 163.367
R1199 B.n625 B.n32 163.367
R1200 B.n621 B.n619 163.367
R1201 B.n617 B.n34 163.367
R1202 B.n613 B.n611 163.367
R1203 B.n609 B.n36 163.367
R1204 B.n605 B.n603 163.367
R1205 B.n601 B.n38 163.367
R1206 B.n597 B.n595 163.367
R1207 B.n593 B.n40 163.367
R1208 B.n589 B.n587 163.367
R1209 B.n585 B.n42 163.367
R1210 B.n581 B.n579 163.367
R1211 B.n577 B.n44 163.367
R1212 B.n573 B.n571 163.367
R1213 B.n569 B.n46 163.367
R1214 B.n565 B.n563 163.367
R1215 B.n561 B.n48 163.367
R1216 B.n557 B.n555 163.367
R1217 B.n553 B.n50 163.367
R1218 B.n549 B.n547 163.367
R1219 B.n545 B.n52 163.367
R1220 B.n541 B.n539 163.367
R1221 B.n536 B.n535 163.367
R1222 B.n533 B.n58 163.367
R1223 B.n529 B.n527 163.367
R1224 B.n525 B.n60 163.367
R1225 B.n520 B.n518 163.367
R1226 B.n516 B.n64 163.367
R1227 B.n512 B.n510 163.367
R1228 B.n508 B.n66 163.367
R1229 B.n504 B.n502 163.367
R1230 B.n500 B.n68 163.367
R1231 B.n496 B.n494 163.367
R1232 B.n492 B.n70 163.367
R1233 B.n488 B.n486 163.367
R1234 B.n484 B.n72 163.367
R1235 B.n480 B.n478 163.367
R1236 B.n476 B.n74 163.367
R1237 B.n472 B.n470 163.367
R1238 B.n468 B.n76 163.367
R1239 B.n464 B.n462 163.367
R1240 B.n460 B.n78 163.367
R1241 B.n456 B.n454 163.367
R1242 B.n452 B.n80 163.367
R1243 B.n448 B.n446 163.367
R1244 B.n444 B.n82 163.367
R1245 B.n440 B.n438 163.367
R1246 B.n436 B.n84 163.367
R1247 B.n432 B.n430 163.367
R1248 B.n370 B.n111 72.4503
R1249 B.n634 B.n29 72.4503
R1250 B.n364 B.n112 71.676
R1251 B.n362 B.n114 71.676
R1252 B.n358 B.n357 71.676
R1253 B.n351 B.n116 71.676
R1254 B.n350 B.n349 71.676
R1255 B.n343 B.n118 71.676
R1256 B.n342 B.n341 71.676
R1257 B.n335 B.n120 71.676
R1258 B.n334 B.n333 71.676
R1259 B.n327 B.n122 71.676
R1260 B.n326 B.n325 71.676
R1261 B.n319 B.n124 71.676
R1262 B.n318 B.n317 71.676
R1263 B.n311 B.n126 71.676
R1264 B.n310 B.n309 71.676
R1265 B.n303 B.n128 71.676
R1266 B.n302 B.n301 71.676
R1267 B.n295 B.n130 71.676
R1268 B.n294 B.n293 71.676
R1269 B.n287 B.n132 71.676
R1270 B.n286 B.n285 71.676
R1271 B.n279 B.n134 71.676
R1272 B.n278 B.n277 71.676
R1273 B.n271 B.n136 71.676
R1274 B.n270 B.n269 71.676
R1275 B.n263 B.n141 71.676
R1276 B.n262 B.n261 71.676
R1277 B.n254 B.n143 71.676
R1278 B.n253 B.n252 71.676
R1279 B.n246 B.n147 71.676
R1280 B.n245 B.n244 71.676
R1281 B.n238 B.n149 71.676
R1282 B.n237 B.n236 71.676
R1283 B.n230 B.n151 71.676
R1284 B.n229 B.n228 71.676
R1285 B.n222 B.n153 71.676
R1286 B.n221 B.n220 71.676
R1287 B.n214 B.n155 71.676
R1288 B.n213 B.n212 71.676
R1289 B.n206 B.n157 71.676
R1290 B.n205 B.n204 71.676
R1291 B.n198 B.n159 71.676
R1292 B.n197 B.n196 71.676
R1293 B.n190 B.n161 71.676
R1294 B.n189 B.n188 71.676
R1295 B.n182 B.n163 71.676
R1296 B.n181 B.n180 71.676
R1297 B.n174 B.n165 71.676
R1298 B.n173 B.n172 71.676
R1299 B.n168 B.n167 71.676
R1300 B.n628 B.n30 71.676
R1301 B.n627 B.n626 71.676
R1302 B.n620 B.n32 71.676
R1303 B.n619 B.n618 71.676
R1304 B.n612 B.n34 71.676
R1305 B.n611 B.n610 71.676
R1306 B.n604 B.n36 71.676
R1307 B.n603 B.n602 71.676
R1308 B.n596 B.n38 71.676
R1309 B.n595 B.n594 71.676
R1310 B.n588 B.n40 71.676
R1311 B.n587 B.n586 71.676
R1312 B.n580 B.n42 71.676
R1313 B.n579 B.n578 71.676
R1314 B.n572 B.n44 71.676
R1315 B.n571 B.n570 71.676
R1316 B.n564 B.n46 71.676
R1317 B.n563 B.n562 71.676
R1318 B.n556 B.n48 71.676
R1319 B.n555 B.n554 71.676
R1320 B.n548 B.n50 71.676
R1321 B.n547 B.n546 71.676
R1322 B.n540 B.n52 71.676
R1323 B.n539 B.n56 71.676
R1324 B.n535 B.n534 71.676
R1325 B.n528 B.n58 71.676
R1326 B.n527 B.n526 71.676
R1327 B.n519 B.n60 71.676
R1328 B.n518 B.n517 71.676
R1329 B.n511 B.n64 71.676
R1330 B.n510 B.n509 71.676
R1331 B.n503 B.n66 71.676
R1332 B.n502 B.n501 71.676
R1333 B.n495 B.n68 71.676
R1334 B.n494 B.n493 71.676
R1335 B.n487 B.n70 71.676
R1336 B.n486 B.n485 71.676
R1337 B.n479 B.n72 71.676
R1338 B.n478 B.n477 71.676
R1339 B.n471 B.n74 71.676
R1340 B.n470 B.n469 71.676
R1341 B.n463 B.n76 71.676
R1342 B.n462 B.n461 71.676
R1343 B.n455 B.n78 71.676
R1344 B.n454 B.n453 71.676
R1345 B.n447 B.n80 71.676
R1346 B.n446 B.n445 71.676
R1347 B.n439 B.n82 71.676
R1348 B.n438 B.n437 71.676
R1349 B.n431 B.n84 71.676
R1350 B.n432 B.n431 71.676
R1351 B.n437 B.n436 71.676
R1352 B.n440 B.n439 71.676
R1353 B.n445 B.n444 71.676
R1354 B.n448 B.n447 71.676
R1355 B.n453 B.n452 71.676
R1356 B.n456 B.n455 71.676
R1357 B.n461 B.n460 71.676
R1358 B.n464 B.n463 71.676
R1359 B.n469 B.n468 71.676
R1360 B.n472 B.n471 71.676
R1361 B.n477 B.n476 71.676
R1362 B.n480 B.n479 71.676
R1363 B.n485 B.n484 71.676
R1364 B.n488 B.n487 71.676
R1365 B.n493 B.n492 71.676
R1366 B.n496 B.n495 71.676
R1367 B.n501 B.n500 71.676
R1368 B.n504 B.n503 71.676
R1369 B.n509 B.n508 71.676
R1370 B.n512 B.n511 71.676
R1371 B.n517 B.n516 71.676
R1372 B.n520 B.n519 71.676
R1373 B.n526 B.n525 71.676
R1374 B.n529 B.n528 71.676
R1375 B.n534 B.n533 71.676
R1376 B.n536 B.n56 71.676
R1377 B.n541 B.n540 71.676
R1378 B.n546 B.n545 71.676
R1379 B.n549 B.n548 71.676
R1380 B.n554 B.n553 71.676
R1381 B.n557 B.n556 71.676
R1382 B.n562 B.n561 71.676
R1383 B.n565 B.n564 71.676
R1384 B.n570 B.n569 71.676
R1385 B.n573 B.n572 71.676
R1386 B.n578 B.n577 71.676
R1387 B.n581 B.n580 71.676
R1388 B.n586 B.n585 71.676
R1389 B.n589 B.n588 71.676
R1390 B.n594 B.n593 71.676
R1391 B.n597 B.n596 71.676
R1392 B.n602 B.n601 71.676
R1393 B.n605 B.n604 71.676
R1394 B.n610 B.n609 71.676
R1395 B.n613 B.n612 71.676
R1396 B.n618 B.n617 71.676
R1397 B.n621 B.n620 71.676
R1398 B.n626 B.n625 71.676
R1399 B.n629 B.n628 71.676
R1400 B.n365 B.n364 71.676
R1401 B.n359 B.n114 71.676
R1402 B.n357 B.n356 71.676
R1403 B.n352 B.n351 71.676
R1404 B.n349 B.n348 71.676
R1405 B.n344 B.n343 71.676
R1406 B.n341 B.n340 71.676
R1407 B.n336 B.n335 71.676
R1408 B.n333 B.n332 71.676
R1409 B.n328 B.n327 71.676
R1410 B.n325 B.n324 71.676
R1411 B.n320 B.n319 71.676
R1412 B.n317 B.n316 71.676
R1413 B.n312 B.n311 71.676
R1414 B.n309 B.n308 71.676
R1415 B.n304 B.n303 71.676
R1416 B.n301 B.n300 71.676
R1417 B.n296 B.n295 71.676
R1418 B.n293 B.n292 71.676
R1419 B.n288 B.n287 71.676
R1420 B.n285 B.n284 71.676
R1421 B.n280 B.n279 71.676
R1422 B.n277 B.n276 71.676
R1423 B.n272 B.n271 71.676
R1424 B.n269 B.n268 71.676
R1425 B.n264 B.n263 71.676
R1426 B.n261 B.n260 71.676
R1427 B.n255 B.n254 71.676
R1428 B.n252 B.n251 71.676
R1429 B.n247 B.n246 71.676
R1430 B.n244 B.n243 71.676
R1431 B.n239 B.n238 71.676
R1432 B.n236 B.n235 71.676
R1433 B.n231 B.n230 71.676
R1434 B.n228 B.n227 71.676
R1435 B.n223 B.n222 71.676
R1436 B.n220 B.n219 71.676
R1437 B.n215 B.n214 71.676
R1438 B.n212 B.n211 71.676
R1439 B.n207 B.n206 71.676
R1440 B.n204 B.n203 71.676
R1441 B.n199 B.n198 71.676
R1442 B.n196 B.n195 71.676
R1443 B.n191 B.n190 71.676
R1444 B.n188 B.n187 71.676
R1445 B.n183 B.n182 71.676
R1446 B.n180 B.n179 71.676
R1447 B.n175 B.n174 71.676
R1448 B.n172 B.n171 71.676
R1449 B.n167 B.n110 71.676
R1450 B.n258 B.n145 59.5399
R1451 B.n139 B.n138 59.5399
R1452 B.n55 B.n54 59.5399
R1453 B.n522 B.n62 59.5399
R1454 B.n370 B.n107 40.054
R1455 B.n376 B.n107 40.054
R1456 B.n376 B.n103 40.054
R1457 B.n382 B.n103 40.054
R1458 B.n388 B.n99 40.054
R1459 B.n388 B.n95 40.054
R1460 B.n394 B.n95 40.054
R1461 B.n394 B.n91 40.054
R1462 B.n401 B.n91 40.054
R1463 B.n407 B.n87 40.054
R1464 B.n407 B.n4 40.054
R1465 B.n660 B.n4 40.054
R1466 B.n660 B.n659 40.054
R1467 B.n659 B.n658 40.054
R1468 B.n658 B.n8 40.054
R1469 B.n652 B.n651 40.054
R1470 B.n651 B.n650 40.054
R1471 B.n650 B.n15 40.054
R1472 B.n644 B.n15 40.054
R1473 B.n644 B.n643 40.054
R1474 B.n642 B.n22 40.054
R1475 B.n636 B.n22 40.054
R1476 B.n636 B.n635 40.054
R1477 B.n635 B.n634 40.054
R1478 B.n401 B.t0 37.1089
R1479 B.n652 B.t1 37.1089
R1480 B.n632 B.n631 32.6249
R1481 B.n429 B.n428 32.6249
R1482 B.n372 B.n109 32.6249
R1483 B.n368 B.n367 32.6249
R1484 B.n382 B.t3 31.2187
R1485 B.t7 B.n642 31.2187
R1486 B.n145 B.n144 19.3944
R1487 B.n138 B.n137 19.3944
R1488 B.n54 B.n53 19.3944
R1489 B.n62 B.n61 19.3944
R1490 B B.n662 18.0485
R1491 B.n631 B.n630 10.6151
R1492 B.n630 B.n31 10.6151
R1493 B.n624 B.n31 10.6151
R1494 B.n624 B.n623 10.6151
R1495 B.n623 B.n622 10.6151
R1496 B.n622 B.n33 10.6151
R1497 B.n616 B.n33 10.6151
R1498 B.n616 B.n615 10.6151
R1499 B.n615 B.n614 10.6151
R1500 B.n614 B.n35 10.6151
R1501 B.n608 B.n35 10.6151
R1502 B.n608 B.n607 10.6151
R1503 B.n607 B.n606 10.6151
R1504 B.n606 B.n37 10.6151
R1505 B.n600 B.n37 10.6151
R1506 B.n600 B.n599 10.6151
R1507 B.n599 B.n598 10.6151
R1508 B.n598 B.n39 10.6151
R1509 B.n592 B.n39 10.6151
R1510 B.n592 B.n591 10.6151
R1511 B.n591 B.n590 10.6151
R1512 B.n590 B.n41 10.6151
R1513 B.n584 B.n41 10.6151
R1514 B.n584 B.n583 10.6151
R1515 B.n583 B.n582 10.6151
R1516 B.n582 B.n43 10.6151
R1517 B.n576 B.n43 10.6151
R1518 B.n576 B.n575 10.6151
R1519 B.n575 B.n574 10.6151
R1520 B.n574 B.n45 10.6151
R1521 B.n568 B.n45 10.6151
R1522 B.n568 B.n567 10.6151
R1523 B.n567 B.n566 10.6151
R1524 B.n566 B.n47 10.6151
R1525 B.n560 B.n47 10.6151
R1526 B.n560 B.n559 10.6151
R1527 B.n559 B.n558 10.6151
R1528 B.n558 B.n49 10.6151
R1529 B.n552 B.n49 10.6151
R1530 B.n552 B.n551 10.6151
R1531 B.n551 B.n550 10.6151
R1532 B.n550 B.n51 10.6151
R1533 B.n544 B.n51 10.6151
R1534 B.n544 B.n543 10.6151
R1535 B.n543 B.n542 10.6151
R1536 B.n538 B.n537 10.6151
R1537 B.n537 B.n57 10.6151
R1538 B.n532 B.n57 10.6151
R1539 B.n532 B.n531 10.6151
R1540 B.n531 B.n530 10.6151
R1541 B.n530 B.n59 10.6151
R1542 B.n524 B.n59 10.6151
R1543 B.n524 B.n523 10.6151
R1544 B.n521 B.n63 10.6151
R1545 B.n515 B.n63 10.6151
R1546 B.n515 B.n514 10.6151
R1547 B.n514 B.n513 10.6151
R1548 B.n513 B.n65 10.6151
R1549 B.n507 B.n65 10.6151
R1550 B.n507 B.n506 10.6151
R1551 B.n506 B.n505 10.6151
R1552 B.n505 B.n67 10.6151
R1553 B.n499 B.n67 10.6151
R1554 B.n499 B.n498 10.6151
R1555 B.n498 B.n497 10.6151
R1556 B.n497 B.n69 10.6151
R1557 B.n491 B.n69 10.6151
R1558 B.n491 B.n490 10.6151
R1559 B.n490 B.n489 10.6151
R1560 B.n489 B.n71 10.6151
R1561 B.n483 B.n71 10.6151
R1562 B.n483 B.n482 10.6151
R1563 B.n482 B.n481 10.6151
R1564 B.n481 B.n73 10.6151
R1565 B.n475 B.n73 10.6151
R1566 B.n475 B.n474 10.6151
R1567 B.n474 B.n473 10.6151
R1568 B.n473 B.n75 10.6151
R1569 B.n467 B.n75 10.6151
R1570 B.n467 B.n466 10.6151
R1571 B.n466 B.n465 10.6151
R1572 B.n465 B.n77 10.6151
R1573 B.n459 B.n77 10.6151
R1574 B.n459 B.n458 10.6151
R1575 B.n458 B.n457 10.6151
R1576 B.n457 B.n79 10.6151
R1577 B.n451 B.n79 10.6151
R1578 B.n451 B.n450 10.6151
R1579 B.n450 B.n449 10.6151
R1580 B.n449 B.n81 10.6151
R1581 B.n443 B.n81 10.6151
R1582 B.n443 B.n442 10.6151
R1583 B.n442 B.n441 10.6151
R1584 B.n441 B.n83 10.6151
R1585 B.n435 B.n83 10.6151
R1586 B.n435 B.n434 10.6151
R1587 B.n434 B.n433 10.6151
R1588 B.n433 B.n429 10.6151
R1589 B.n373 B.n372 10.6151
R1590 B.n374 B.n373 10.6151
R1591 B.n374 B.n101 10.6151
R1592 B.n384 B.n101 10.6151
R1593 B.n385 B.n384 10.6151
R1594 B.n386 B.n385 10.6151
R1595 B.n386 B.n93 10.6151
R1596 B.n396 B.n93 10.6151
R1597 B.n397 B.n396 10.6151
R1598 B.n399 B.n397 10.6151
R1599 B.n399 B.n398 10.6151
R1600 B.n398 B.n85 10.6151
R1601 B.n410 B.n85 10.6151
R1602 B.n411 B.n410 10.6151
R1603 B.n412 B.n411 10.6151
R1604 B.n413 B.n412 10.6151
R1605 B.n415 B.n413 10.6151
R1606 B.n416 B.n415 10.6151
R1607 B.n417 B.n416 10.6151
R1608 B.n418 B.n417 10.6151
R1609 B.n420 B.n418 10.6151
R1610 B.n421 B.n420 10.6151
R1611 B.n422 B.n421 10.6151
R1612 B.n423 B.n422 10.6151
R1613 B.n425 B.n423 10.6151
R1614 B.n426 B.n425 10.6151
R1615 B.n427 B.n426 10.6151
R1616 B.n428 B.n427 10.6151
R1617 B.n367 B.n366 10.6151
R1618 B.n366 B.n113 10.6151
R1619 B.n361 B.n113 10.6151
R1620 B.n361 B.n360 10.6151
R1621 B.n360 B.n115 10.6151
R1622 B.n355 B.n115 10.6151
R1623 B.n355 B.n354 10.6151
R1624 B.n354 B.n353 10.6151
R1625 B.n353 B.n117 10.6151
R1626 B.n347 B.n117 10.6151
R1627 B.n347 B.n346 10.6151
R1628 B.n346 B.n345 10.6151
R1629 B.n345 B.n119 10.6151
R1630 B.n339 B.n119 10.6151
R1631 B.n339 B.n338 10.6151
R1632 B.n338 B.n337 10.6151
R1633 B.n337 B.n121 10.6151
R1634 B.n331 B.n121 10.6151
R1635 B.n331 B.n330 10.6151
R1636 B.n330 B.n329 10.6151
R1637 B.n329 B.n123 10.6151
R1638 B.n323 B.n123 10.6151
R1639 B.n323 B.n322 10.6151
R1640 B.n322 B.n321 10.6151
R1641 B.n321 B.n125 10.6151
R1642 B.n315 B.n125 10.6151
R1643 B.n315 B.n314 10.6151
R1644 B.n314 B.n313 10.6151
R1645 B.n313 B.n127 10.6151
R1646 B.n307 B.n127 10.6151
R1647 B.n307 B.n306 10.6151
R1648 B.n306 B.n305 10.6151
R1649 B.n305 B.n129 10.6151
R1650 B.n299 B.n129 10.6151
R1651 B.n299 B.n298 10.6151
R1652 B.n298 B.n297 10.6151
R1653 B.n297 B.n131 10.6151
R1654 B.n291 B.n131 10.6151
R1655 B.n291 B.n290 10.6151
R1656 B.n290 B.n289 10.6151
R1657 B.n289 B.n133 10.6151
R1658 B.n283 B.n133 10.6151
R1659 B.n283 B.n282 10.6151
R1660 B.n282 B.n281 10.6151
R1661 B.n281 B.n135 10.6151
R1662 B.n275 B.n274 10.6151
R1663 B.n274 B.n273 10.6151
R1664 B.n273 B.n140 10.6151
R1665 B.n267 B.n140 10.6151
R1666 B.n267 B.n266 10.6151
R1667 B.n266 B.n265 10.6151
R1668 B.n265 B.n142 10.6151
R1669 B.n259 B.n142 10.6151
R1670 B.n257 B.n256 10.6151
R1671 B.n256 B.n146 10.6151
R1672 B.n250 B.n146 10.6151
R1673 B.n250 B.n249 10.6151
R1674 B.n249 B.n248 10.6151
R1675 B.n248 B.n148 10.6151
R1676 B.n242 B.n148 10.6151
R1677 B.n242 B.n241 10.6151
R1678 B.n241 B.n240 10.6151
R1679 B.n240 B.n150 10.6151
R1680 B.n234 B.n150 10.6151
R1681 B.n234 B.n233 10.6151
R1682 B.n233 B.n232 10.6151
R1683 B.n232 B.n152 10.6151
R1684 B.n226 B.n152 10.6151
R1685 B.n226 B.n225 10.6151
R1686 B.n225 B.n224 10.6151
R1687 B.n224 B.n154 10.6151
R1688 B.n218 B.n154 10.6151
R1689 B.n218 B.n217 10.6151
R1690 B.n217 B.n216 10.6151
R1691 B.n216 B.n156 10.6151
R1692 B.n210 B.n156 10.6151
R1693 B.n210 B.n209 10.6151
R1694 B.n209 B.n208 10.6151
R1695 B.n208 B.n158 10.6151
R1696 B.n202 B.n158 10.6151
R1697 B.n202 B.n201 10.6151
R1698 B.n201 B.n200 10.6151
R1699 B.n200 B.n160 10.6151
R1700 B.n194 B.n160 10.6151
R1701 B.n194 B.n193 10.6151
R1702 B.n193 B.n192 10.6151
R1703 B.n192 B.n162 10.6151
R1704 B.n186 B.n162 10.6151
R1705 B.n186 B.n185 10.6151
R1706 B.n185 B.n184 10.6151
R1707 B.n184 B.n164 10.6151
R1708 B.n178 B.n164 10.6151
R1709 B.n178 B.n177 10.6151
R1710 B.n177 B.n176 10.6151
R1711 B.n176 B.n166 10.6151
R1712 B.n170 B.n166 10.6151
R1713 B.n170 B.n169 10.6151
R1714 B.n169 B.n109 10.6151
R1715 B.n368 B.n105 10.6151
R1716 B.n378 B.n105 10.6151
R1717 B.n379 B.n378 10.6151
R1718 B.n380 B.n379 10.6151
R1719 B.n380 B.n97 10.6151
R1720 B.n390 B.n97 10.6151
R1721 B.n391 B.n390 10.6151
R1722 B.n392 B.n391 10.6151
R1723 B.n392 B.n89 10.6151
R1724 B.n403 B.n89 10.6151
R1725 B.n404 B.n403 10.6151
R1726 B.n405 B.n404 10.6151
R1727 B.n405 B.n0 10.6151
R1728 B.n656 B.n1 10.6151
R1729 B.n656 B.n655 10.6151
R1730 B.n655 B.n654 10.6151
R1731 B.n654 B.n10 10.6151
R1732 B.n648 B.n10 10.6151
R1733 B.n648 B.n647 10.6151
R1734 B.n647 B.n646 10.6151
R1735 B.n646 B.n17 10.6151
R1736 B.n640 B.n17 10.6151
R1737 B.n640 B.n639 10.6151
R1738 B.n639 B.n638 10.6151
R1739 B.n638 B.n24 10.6151
R1740 B.n632 B.n24 10.6151
R1741 B.t3 B.n99 8.83584
R1742 B.n643 B.t7 8.83584
R1743 B.n538 B.n55 7.18099
R1744 B.n523 B.n522 7.18099
R1745 B.n275 B.n139 7.18099
R1746 B.n259 B.n258 7.18099
R1747 B.n542 B.n55 3.43465
R1748 B.n522 B.n521 3.43465
R1749 B.n139 B.n135 3.43465
R1750 B.n258 B.n257 3.43465
R1751 B.t0 B.n87 2.94561
R1752 B.t1 B.n8 2.94561
R1753 B.n662 B.n0 2.81026
R1754 B.n662 B.n1 2.81026
R1755 VP.n0 VP.t0 742.53
R1756 VP.n0 VP.t1 701.932
R1757 VP VP.n0 0.0516364
R1758 VDD1.n66 VDD1.n0 214.453
R1759 VDD1.n137 VDD1.n71 214.453
R1760 VDD1.n67 VDD1.n66 185
R1761 VDD1.n65 VDD1.n64 185
R1762 VDD1.n4 VDD1.n3 185
R1763 VDD1.n59 VDD1.n58 185
R1764 VDD1.n57 VDD1.n56 185
R1765 VDD1.n8 VDD1.n7 185
R1766 VDD1.n51 VDD1.n50 185
R1767 VDD1.n49 VDD1.n48 185
R1768 VDD1.n12 VDD1.n11 185
R1769 VDD1.n43 VDD1.n42 185
R1770 VDD1.n41 VDD1.n40 185
R1771 VDD1.n16 VDD1.n15 185
R1772 VDD1.n35 VDD1.n34 185
R1773 VDD1.n33 VDD1.n32 185
R1774 VDD1.n20 VDD1.n19 185
R1775 VDD1.n27 VDD1.n26 185
R1776 VDD1.n25 VDD1.n24 185
R1777 VDD1.n96 VDD1.n95 185
R1778 VDD1.n98 VDD1.n97 185
R1779 VDD1.n91 VDD1.n90 185
R1780 VDD1.n104 VDD1.n103 185
R1781 VDD1.n106 VDD1.n105 185
R1782 VDD1.n87 VDD1.n86 185
R1783 VDD1.n112 VDD1.n111 185
R1784 VDD1.n114 VDD1.n113 185
R1785 VDD1.n83 VDD1.n82 185
R1786 VDD1.n120 VDD1.n119 185
R1787 VDD1.n122 VDD1.n121 185
R1788 VDD1.n79 VDD1.n78 185
R1789 VDD1.n128 VDD1.n127 185
R1790 VDD1.n130 VDD1.n129 185
R1791 VDD1.n75 VDD1.n74 185
R1792 VDD1.n136 VDD1.n135 185
R1793 VDD1.n138 VDD1.n137 185
R1794 VDD1.n94 VDD1.t0 147.659
R1795 VDD1.n23 VDD1.t1 147.659
R1796 VDD1.n66 VDD1.n65 104.615
R1797 VDD1.n65 VDD1.n3 104.615
R1798 VDD1.n58 VDD1.n3 104.615
R1799 VDD1.n58 VDD1.n57 104.615
R1800 VDD1.n57 VDD1.n7 104.615
R1801 VDD1.n50 VDD1.n7 104.615
R1802 VDD1.n50 VDD1.n49 104.615
R1803 VDD1.n49 VDD1.n11 104.615
R1804 VDD1.n42 VDD1.n11 104.615
R1805 VDD1.n42 VDD1.n41 104.615
R1806 VDD1.n41 VDD1.n15 104.615
R1807 VDD1.n34 VDD1.n15 104.615
R1808 VDD1.n34 VDD1.n33 104.615
R1809 VDD1.n33 VDD1.n19 104.615
R1810 VDD1.n26 VDD1.n19 104.615
R1811 VDD1.n26 VDD1.n25 104.615
R1812 VDD1.n97 VDD1.n96 104.615
R1813 VDD1.n97 VDD1.n90 104.615
R1814 VDD1.n104 VDD1.n90 104.615
R1815 VDD1.n105 VDD1.n104 104.615
R1816 VDD1.n105 VDD1.n86 104.615
R1817 VDD1.n112 VDD1.n86 104.615
R1818 VDD1.n113 VDD1.n112 104.615
R1819 VDD1.n113 VDD1.n82 104.615
R1820 VDD1.n120 VDD1.n82 104.615
R1821 VDD1.n121 VDD1.n120 104.615
R1822 VDD1.n121 VDD1.n78 104.615
R1823 VDD1.n128 VDD1.n78 104.615
R1824 VDD1.n129 VDD1.n128 104.615
R1825 VDD1.n129 VDD1.n74 104.615
R1826 VDD1.n136 VDD1.n74 104.615
R1827 VDD1.n137 VDD1.n136 104.615
R1828 VDD1 VDD1.n141 90.0307
R1829 VDD1 VDD1.n70 52.6288
R1830 VDD1.n25 VDD1.t1 52.3082
R1831 VDD1.n96 VDD1.t0 52.3082
R1832 VDD1.n24 VDD1.n23 15.6677
R1833 VDD1.n95 VDD1.n94 15.6677
R1834 VDD1.n68 VDD1.n67 12.8005
R1835 VDD1.n27 VDD1.n22 12.8005
R1836 VDD1.n98 VDD1.n93 12.8005
R1837 VDD1.n139 VDD1.n138 12.8005
R1838 VDD1.n64 VDD1.n2 12.0247
R1839 VDD1.n28 VDD1.n20 12.0247
R1840 VDD1.n99 VDD1.n91 12.0247
R1841 VDD1.n135 VDD1.n73 12.0247
R1842 VDD1.n63 VDD1.n4 11.249
R1843 VDD1.n32 VDD1.n31 11.249
R1844 VDD1.n103 VDD1.n102 11.249
R1845 VDD1.n134 VDD1.n75 11.249
R1846 VDD1.n60 VDD1.n59 10.4732
R1847 VDD1.n35 VDD1.n18 10.4732
R1848 VDD1.n106 VDD1.n89 10.4732
R1849 VDD1.n131 VDD1.n130 10.4732
R1850 VDD1.n56 VDD1.n6 9.69747
R1851 VDD1.n36 VDD1.n16 9.69747
R1852 VDD1.n107 VDD1.n87 9.69747
R1853 VDD1.n127 VDD1.n77 9.69747
R1854 VDD1.n70 VDD1.n69 9.45567
R1855 VDD1.n141 VDD1.n140 9.45567
R1856 VDD1.n10 VDD1.n9 9.3005
R1857 VDD1.n53 VDD1.n52 9.3005
R1858 VDD1.n55 VDD1.n54 9.3005
R1859 VDD1.n6 VDD1.n5 9.3005
R1860 VDD1.n61 VDD1.n60 9.3005
R1861 VDD1.n63 VDD1.n62 9.3005
R1862 VDD1.n2 VDD1.n1 9.3005
R1863 VDD1.n69 VDD1.n68 9.3005
R1864 VDD1.n47 VDD1.n46 9.3005
R1865 VDD1.n45 VDD1.n44 9.3005
R1866 VDD1.n14 VDD1.n13 9.3005
R1867 VDD1.n39 VDD1.n38 9.3005
R1868 VDD1.n37 VDD1.n36 9.3005
R1869 VDD1.n18 VDD1.n17 9.3005
R1870 VDD1.n31 VDD1.n30 9.3005
R1871 VDD1.n29 VDD1.n28 9.3005
R1872 VDD1.n22 VDD1.n21 9.3005
R1873 VDD1.n116 VDD1.n115 9.3005
R1874 VDD1.n85 VDD1.n84 9.3005
R1875 VDD1.n110 VDD1.n109 9.3005
R1876 VDD1.n108 VDD1.n107 9.3005
R1877 VDD1.n89 VDD1.n88 9.3005
R1878 VDD1.n102 VDD1.n101 9.3005
R1879 VDD1.n100 VDD1.n99 9.3005
R1880 VDD1.n93 VDD1.n92 9.3005
R1881 VDD1.n118 VDD1.n117 9.3005
R1882 VDD1.n81 VDD1.n80 9.3005
R1883 VDD1.n124 VDD1.n123 9.3005
R1884 VDD1.n126 VDD1.n125 9.3005
R1885 VDD1.n77 VDD1.n76 9.3005
R1886 VDD1.n132 VDD1.n131 9.3005
R1887 VDD1.n134 VDD1.n133 9.3005
R1888 VDD1.n73 VDD1.n72 9.3005
R1889 VDD1.n140 VDD1.n139 9.3005
R1890 VDD1.n55 VDD1.n8 8.92171
R1891 VDD1.n40 VDD1.n39 8.92171
R1892 VDD1.n111 VDD1.n110 8.92171
R1893 VDD1.n126 VDD1.n79 8.92171
R1894 VDD1.n70 VDD1.n0 8.2187
R1895 VDD1.n141 VDD1.n71 8.2187
R1896 VDD1.n52 VDD1.n51 8.14595
R1897 VDD1.n43 VDD1.n14 8.14595
R1898 VDD1.n114 VDD1.n85 8.14595
R1899 VDD1.n123 VDD1.n122 8.14595
R1900 VDD1.n48 VDD1.n10 7.3702
R1901 VDD1.n44 VDD1.n12 7.3702
R1902 VDD1.n115 VDD1.n83 7.3702
R1903 VDD1.n119 VDD1.n81 7.3702
R1904 VDD1.n48 VDD1.n47 6.59444
R1905 VDD1.n47 VDD1.n12 6.59444
R1906 VDD1.n118 VDD1.n83 6.59444
R1907 VDD1.n119 VDD1.n118 6.59444
R1908 VDD1.n51 VDD1.n10 5.81868
R1909 VDD1.n44 VDD1.n43 5.81868
R1910 VDD1.n115 VDD1.n114 5.81868
R1911 VDD1.n122 VDD1.n81 5.81868
R1912 VDD1.n68 VDD1.n0 5.3904
R1913 VDD1.n139 VDD1.n71 5.3904
R1914 VDD1.n52 VDD1.n8 5.04292
R1915 VDD1.n40 VDD1.n14 5.04292
R1916 VDD1.n111 VDD1.n85 5.04292
R1917 VDD1.n123 VDD1.n79 5.04292
R1918 VDD1.n94 VDD1.n92 4.38563
R1919 VDD1.n23 VDD1.n21 4.38563
R1920 VDD1.n56 VDD1.n55 4.26717
R1921 VDD1.n39 VDD1.n16 4.26717
R1922 VDD1.n110 VDD1.n87 4.26717
R1923 VDD1.n127 VDD1.n126 4.26717
R1924 VDD1.n59 VDD1.n6 3.49141
R1925 VDD1.n36 VDD1.n35 3.49141
R1926 VDD1.n107 VDD1.n106 3.49141
R1927 VDD1.n130 VDD1.n77 3.49141
R1928 VDD1.n60 VDD1.n4 2.71565
R1929 VDD1.n32 VDD1.n18 2.71565
R1930 VDD1.n103 VDD1.n89 2.71565
R1931 VDD1.n131 VDD1.n75 2.71565
R1932 VDD1.n64 VDD1.n63 1.93989
R1933 VDD1.n31 VDD1.n20 1.93989
R1934 VDD1.n102 VDD1.n91 1.93989
R1935 VDD1.n135 VDD1.n134 1.93989
R1936 VDD1.n67 VDD1.n2 1.16414
R1937 VDD1.n28 VDD1.n27 1.16414
R1938 VDD1.n99 VDD1.n98 1.16414
R1939 VDD1.n138 VDD1.n73 1.16414
R1940 VDD1.n24 VDD1.n22 0.388379
R1941 VDD1.n95 VDD1.n93 0.388379
R1942 VDD1.n69 VDD1.n1 0.155672
R1943 VDD1.n62 VDD1.n1 0.155672
R1944 VDD1.n62 VDD1.n61 0.155672
R1945 VDD1.n61 VDD1.n5 0.155672
R1946 VDD1.n54 VDD1.n5 0.155672
R1947 VDD1.n54 VDD1.n53 0.155672
R1948 VDD1.n53 VDD1.n9 0.155672
R1949 VDD1.n46 VDD1.n9 0.155672
R1950 VDD1.n46 VDD1.n45 0.155672
R1951 VDD1.n45 VDD1.n13 0.155672
R1952 VDD1.n38 VDD1.n13 0.155672
R1953 VDD1.n38 VDD1.n37 0.155672
R1954 VDD1.n37 VDD1.n17 0.155672
R1955 VDD1.n30 VDD1.n17 0.155672
R1956 VDD1.n30 VDD1.n29 0.155672
R1957 VDD1.n29 VDD1.n21 0.155672
R1958 VDD1.n100 VDD1.n92 0.155672
R1959 VDD1.n101 VDD1.n100 0.155672
R1960 VDD1.n101 VDD1.n88 0.155672
R1961 VDD1.n108 VDD1.n88 0.155672
R1962 VDD1.n109 VDD1.n108 0.155672
R1963 VDD1.n109 VDD1.n84 0.155672
R1964 VDD1.n116 VDD1.n84 0.155672
R1965 VDD1.n117 VDD1.n116 0.155672
R1966 VDD1.n117 VDD1.n80 0.155672
R1967 VDD1.n124 VDD1.n80 0.155672
R1968 VDD1.n125 VDD1.n124 0.155672
R1969 VDD1.n125 VDD1.n76 0.155672
R1970 VDD1.n132 VDD1.n76 0.155672
R1971 VDD1.n133 VDD1.n132 0.155672
R1972 VDD1.n133 VDD1.n72 0.155672
R1973 VDD1.n140 VDD1.n72 0.155672
C0 VDD1 VN 0.148242f
C1 VDD2 VN 2.15237f
C2 VP VTAIL 1.59336f
C3 VDD1 VTAIL 6.22402f
C4 VDD2 VTAIL 6.25676f
C5 VP VDD1 2.25288f
C6 VP VDD2 0.253632f
C7 VDD1 VDD2 0.459664f
C8 VN VTAIL 1.57869f
C9 VP VN 4.80584f
C10 VDD2 B 3.994073f
C11 VDD1 B 6.57274f
C12 VTAIL B 6.893832f
C13 VN B 8.473651f
C14 VP B 4.086743f
C15 VDD1.n0 B 0.029155f
C16 VDD1.n1 B 0.021046f
C17 VDD1.n2 B 0.011309f
C18 VDD1.n3 B 0.026731f
C19 VDD1.n4 B 0.011974f
C20 VDD1.n5 B 0.021046f
C21 VDD1.n6 B 0.011309f
C22 VDD1.n7 B 0.026731f
C23 VDD1.n8 B 0.011974f
C24 VDD1.n9 B 0.021046f
C25 VDD1.n10 B 0.011309f
C26 VDD1.n11 B 0.026731f
C27 VDD1.n12 B 0.011974f
C28 VDD1.n13 B 0.021046f
C29 VDD1.n14 B 0.011309f
C30 VDD1.n15 B 0.026731f
C31 VDD1.n16 B 0.011974f
C32 VDD1.n17 B 0.021046f
C33 VDD1.n18 B 0.011309f
C34 VDD1.n19 B 0.026731f
C35 VDD1.n20 B 0.011974f
C36 VDD1.n21 B 1.21302f
C37 VDD1.n22 B 0.011309f
C38 VDD1.t1 B 0.043959f
C39 VDD1.n23 B 0.128717f
C40 VDD1.n24 B 0.015791f
C41 VDD1.n25 B 0.020048f
C42 VDD1.n26 B 0.026731f
C43 VDD1.n27 B 0.011974f
C44 VDD1.n28 B 0.011309f
C45 VDD1.n29 B 0.021046f
C46 VDD1.n30 B 0.021046f
C47 VDD1.n31 B 0.011309f
C48 VDD1.n32 B 0.011974f
C49 VDD1.n33 B 0.026731f
C50 VDD1.n34 B 0.026731f
C51 VDD1.n35 B 0.011974f
C52 VDD1.n36 B 0.011309f
C53 VDD1.n37 B 0.021046f
C54 VDD1.n38 B 0.021046f
C55 VDD1.n39 B 0.011309f
C56 VDD1.n40 B 0.011974f
C57 VDD1.n41 B 0.026731f
C58 VDD1.n42 B 0.026731f
C59 VDD1.n43 B 0.011974f
C60 VDD1.n44 B 0.011309f
C61 VDD1.n45 B 0.021046f
C62 VDD1.n46 B 0.021046f
C63 VDD1.n47 B 0.011309f
C64 VDD1.n48 B 0.011974f
C65 VDD1.n49 B 0.026731f
C66 VDD1.n50 B 0.026731f
C67 VDD1.n51 B 0.011974f
C68 VDD1.n52 B 0.011309f
C69 VDD1.n53 B 0.021046f
C70 VDD1.n54 B 0.021046f
C71 VDD1.n55 B 0.011309f
C72 VDD1.n56 B 0.011974f
C73 VDD1.n57 B 0.026731f
C74 VDD1.n58 B 0.026731f
C75 VDD1.n59 B 0.011974f
C76 VDD1.n60 B 0.011309f
C77 VDD1.n61 B 0.021046f
C78 VDD1.n62 B 0.021046f
C79 VDD1.n63 B 0.011309f
C80 VDD1.n64 B 0.011974f
C81 VDD1.n65 B 0.026731f
C82 VDD1.n66 B 0.055083f
C83 VDD1.n67 B 0.011974f
C84 VDD1.n68 B 0.022113f
C85 VDD1.n69 B 0.053822f
C86 VDD1.n70 B 0.072202f
C87 VDD1.n71 B 0.029155f
C88 VDD1.n72 B 0.021046f
C89 VDD1.n73 B 0.011309f
C90 VDD1.n74 B 0.026731f
C91 VDD1.n75 B 0.011974f
C92 VDD1.n76 B 0.021046f
C93 VDD1.n77 B 0.011309f
C94 VDD1.n78 B 0.026731f
C95 VDD1.n79 B 0.011974f
C96 VDD1.n80 B 0.021046f
C97 VDD1.n81 B 0.011309f
C98 VDD1.n82 B 0.026731f
C99 VDD1.n83 B 0.011974f
C100 VDD1.n84 B 0.021046f
C101 VDD1.n85 B 0.011309f
C102 VDD1.n86 B 0.026731f
C103 VDD1.n87 B 0.011974f
C104 VDD1.n88 B 0.021046f
C105 VDD1.n89 B 0.011309f
C106 VDD1.n90 B 0.026731f
C107 VDD1.n91 B 0.011974f
C108 VDD1.n92 B 1.21302f
C109 VDD1.n93 B 0.011309f
C110 VDD1.t0 B 0.043959f
C111 VDD1.n94 B 0.128717f
C112 VDD1.n95 B 0.015791f
C113 VDD1.n96 B 0.020048f
C114 VDD1.n97 B 0.026731f
C115 VDD1.n98 B 0.011974f
C116 VDD1.n99 B 0.011309f
C117 VDD1.n100 B 0.021046f
C118 VDD1.n101 B 0.021046f
C119 VDD1.n102 B 0.011309f
C120 VDD1.n103 B 0.011974f
C121 VDD1.n104 B 0.026731f
C122 VDD1.n105 B 0.026731f
C123 VDD1.n106 B 0.011974f
C124 VDD1.n107 B 0.011309f
C125 VDD1.n108 B 0.021046f
C126 VDD1.n109 B 0.021046f
C127 VDD1.n110 B 0.011309f
C128 VDD1.n111 B 0.011974f
C129 VDD1.n112 B 0.026731f
C130 VDD1.n113 B 0.026731f
C131 VDD1.n114 B 0.011974f
C132 VDD1.n115 B 0.011309f
C133 VDD1.n116 B 0.021046f
C134 VDD1.n117 B 0.021046f
C135 VDD1.n118 B 0.011309f
C136 VDD1.n119 B 0.011974f
C137 VDD1.n120 B 0.026731f
C138 VDD1.n121 B 0.026731f
C139 VDD1.n122 B 0.011974f
C140 VDD1.n123 B 0.011309f
C141 VDD1.n124 B 0.021046f
C142 VDD1.n125 B 0.021046f
C143 VDD1.n126 B 0.011309f
C144 VDD1.n127 B 0.011974f
C145 VDD1.n128 B 0.026731f
C146 VDD1.n129 B 0.026731f
C147 VDD1.n130 B 0.011974f
C148 VDD1.n131 B 0.011309f
C149 VDD1.n132 B 0.021046f
C150 VDD1.n133 B 0.021046f
C151 VDD1.n134 B 0.011309f
C152 VDD1.n135 B 0.011974f
C153 VDD1.n136 B 0.026731f
C154 VDD1.n137 B 0.055083f
C155 VDD1.n138 B 0.011974f
C156 VDD1.n139 B 0.022113f
C157 VDD1.n140 B 0.053822f
C158 VDD1.n141 B 0.588825f
C159 VP.t0 B 1.43811f
C160 VP.t1 B 1.31719f
C161 VP.n0 B 4.32906f
C162 VDD2.n0 B 0.029424f
C163 VDD2.n1 B 0.02124f
C164 VDD2.n2 B 0.011413f
C165 VDD2.n3 B 0.026977f
C166 VDD2.n4 B 0.012085f
C167 VDD2.n5 B 0.02124f
C168 VDD2.n6 B 0.011413f
C169 VDD2.n7 B 0.026977f
C170 VDD2.n8 B 0.012085f
C171 VDD2.n9 B 0.02124f
C172 VDD2.n10 B 0.011413f
C173 VDD2.n11 B 0.026977f
C174 VDD2.n12 B 0.012085f
C175 VDD2.n13 B 0.02124f
C176 VDD2.n14 B 0.011413f
C177 VDD2.n15 B 0.026977f
C178 VDD2.n16 B 0.012085f
C179 VDD2.n17 B 0.02124f
C180 VDD2.n18 B 0.011413f
C181 VDD2.n19 B 0.026977f
C182 VDD2.n20 B 0.012085f
C183 VDD2.n21 B 1.22421f
C184 VDD2.n22 B 0.011413f
C185 VDD2.t0 B 0.044364f
C186 VDD2.n23 B 0.129905f
C187 VDD2.n24 B 0.015936f
C188 VDD2.n25 B 0.020233f
C189 VDD2.n26 B 0.026977f
C190 VDD2.n27 B 0.012085f
C191 VDD2.n28 B 0.011413f
C192 VDD2.n29 B 0.02124f
C193 VDD2.n30 B 0.02124f
C194 VDD2.n31 B 0.011413f
C195 VDD2.n32 B 0.012085f
C196 VDD2.n33 B 0.026977f
C197 VDD2.n34 B 0.026977f
C198 VDD2.n35 B 0.012085f
C199 VDD2.n36 B 0.011413f
C200 VDD2.n37 B 0.02124f
C201 VDD2.n38 B 0.02124f
C202 VDD2.n39 B 0.011413f
C203 VDD2.n40 B 0.012085f
C204 VDD2.n41 B 0.026977f
C205 VDD2.n42 B 0.026977f
C206 VDD2.n43 B 0.012085f
C207 VDD2.n44 B 0.011413f
C208 VDD2.n45 B 0.02124f
C209 VDD2.n46 B 0.02124f
C210 VDD2.n47 B 0.011413f
C211 VDD2.n48 B 0.012085f
C212 VDD2.n49 B 0.026977f
C213 VDD2.n50 B 0.026977f
C214 VDD2.n51 B 0.012085f
C215 VDD2.n52 B 0.011413f
C216 VDD2.n53 B 0.02124f
C217 VDD2.n54 B 0.02124f
C218 VDD2.n55 B 0.011413f
C219 VDD2.n56 B 0.012085f
C220 VDD2.n57 B 0.026977f
C221 VDD2.n58 B 0.026977f
C222 VDD2.n59 B 0.012085f
C223 VDD2.n60 B 0.011413f
C224 VDD2.n61 B 0.02124f
C225 VDD2.n62 B 0.02124f
C226 VDD2.n63 B 0.011413f
C227 VDD2.n64 B 0.012085f
C228 VDD2.n65 B 0.026977f
C229 VDD2.n66 B 0.055591f
C230 VDD2.n67 B 0.012085f
C231 VDD2.n68 B 0.022317f
C232 VDD2.n69 B 0.054318f
C233 VDD2.n70 B 0.566413f
C234 VDD2.n71 B 0.029424f
C235 VDD2.n72 B 0.02124f
C236 VDD2.n73 B 0.011413f
C237 VDD2.n74 B 0.026977f
C238 VDD2.n75 B 0.012085f
C239 VDD2.n76 B 0.02124f
C240 VDD2.n77 B 0.011413f
C241 VDD2.n78 B 0.026977f
C242 VDD2.n79 B 0.012085f
C243 VDD2.n80 B 0.02124f
C244 VDD2.n81 B 0.011413f
C245 VDD2.n82 B 0.026977f
C246 VDD2.n83 B 0.012085f
C247 VDD2.n84 B 0.02124f
C248 VDD2.n85 B 0.011413f
C249 VDD2.n86 B 0.026977f
C250 VDD2.n87 B 0.012085f
C251 VDD2.n88 B 0.02124f
C252 VDD2.n89 B 0.011413f
C253 VDD2.n90 B 0.026977f
C254 VDD2.n91 B 0.012085f
C255 VDD2.n92 B 1.22421f
C256 VDD2.n93 B 0.011413f
C257 VDD2.t1 B 0.044364f
C258 VDD2.n94 B 0.129905f
C259 VDD2.n95 B 0.015936f
C260 VDD2.n96 B 0.020233f
C261 VDD2.n97 B 0.026977f
C262 VDD2.n98 B 0.012085f
C263 VDD2.n99 B 0.011413f
C264 VDD2.n100 B 0.02124f
C265 VDD2.n101 B 0.02124f
C266 VDD2.n102 B 0.011413f
C267 VDD2.n103 B 0.012085f
C268 VDD2.n104 B 0.026977f
C269 VDD2.n105 B 0.026977f
C270 VDD2.n106 B 0.012085f
C271 VDD2.n107 B 0.011413f
C272 VDD2.n108 B 0.02124f
C273 VDD2.n109 B 0.02124f
C274 VDD2.n110 B 0.011413f
C275 VDD2.n111 B 0.012085f
C276 VDD2.n112 B 0.026977f
C277 VDD2.n113 B 0.026977f
C278 VDD2.n114 B 0.012085f
C279 VDD2.n115 B 0.011413f
C280 VDD2.n116 B 0.02124f
C281 VDD2.n117 B 0.02124f
C282 VDD2.n118 B 0.011413f
C283 VDD2.n119 B 0.012085f
C284 VDD2.n120 B 0.026977f
C285 VDD2.n121 B 0.026977f
C286 VDD2.n122 B 0.012085f
C287 VDD2.n123 B 0.011413f
C288 VDD2.n124 B 0.02124f
C289 VDD2.n125 B 0.02124f
C290 VDD2.n126 B 0.011413f
C291 VDD2.n127 B 0.012085f
C292 VDD2.n128 B 0.026977f
C293 VDD2.n129 B 0.026977f
C294 VDD2.n130 B 0.012085f
C295 VDD2.n131 B 0.011413f
C296 VDD2.n132 B 0.02124f
C297 VDD2.n133 B 0.02124f
C298 VDD2.n134 B 0.011413f
C299 VDD2.n135 B 0.012085f
C300 VDD2.n136 B 0.026977f
C301 VDD2.n137 B 0.055591f
C302 VDD2.n138 B 0.012085f
C303 VDD2.n139 B 0.022317f
C304 VDD2.n140 B 0.054318f
C305 VDD2.n141 B 0.072543f
C306 VDD2.n142 B 2.42115f
C307 VTAIL.n0 B 0.022966f
C308 VTAIL.n1 B 0.016578f
C309 VTAIL.n2 B 0.008908f
C310 VTAIL.n3 B 0.021056f
C311 VTAIL.n4 B 0.009432f
C312 VTAIL.n5 B 0.016578f
C313 VTAIL.n6 B 0.008908f
C314 VTAIL.n7 B 0.021056f
C315 VTAIL.n8 B 0.009432f
C316 VTAIL.n9 B 0.016578f
C317 VTAIL.n10 B 0.008908f
C318 VTAIL.n11 B 0.021056f
C319 VTAIL.n12 B 0.009432f
C320 VTAIL.n13 B 0.016578f
C321 VTAIL.n14 B 0.008908f
C322 VTAIL.n15 B 0.021056f
C323 VTAIL.n16 B 0.009432f
C324 VTAIL.n17 B 0.016578f
C325 VTAIL.n18 B 0.008908f
C326 VTAIL.n19 B 0.021056f
C327 VTAIL.n20 B 0.009432f
C328 VTAIL.n21 B 0.955502f
C329 VTAIL.n22 B 0.008908f
C330 VTAIL.t0 B 0.034626f
C331 VTAIL.n23 B 0.101391f
C332 VTAIL.n24 B 0.012438f
C333 VTAIL.n25 B 0.015792f
C334 VTAIL.n26 B 0.021056f
C335 VTAIL.n27 B 0.009432f
C336 VTAIL.n28 B 0.008908f
C337 VTAIL.n29 B 0.016578f
C338 VTAIL.n30 B 0.016578f
C339 VTAIL.n31 B 0.008908f
C340 VTAIL.n32 B 0.009432f
C341 VTAIL.n33 B 0.021056f
C342 VTAIL.n34 B 0.021056f
C343 VTAIL.n35 B 0.009432f
C344 VTAIL.n36 B 0.008908f
C345 VTAIL.n37 B 0.016578f
C346 VTAIL.n38 B 0.016578f
C347 VTAIL.n39 B 0.008908f
C348 VTAIL.n40 B 0.009432f
C349 VTAIL.n41 B 0.021056f
C350 VTAIL.n42 B 0.021056f
C351 VTAIL.n43 B 0.009432f
C352 VTAIL.n44 B 0.008908f
C353 VTAIL.n45 B 0.016578f
C354 VTAIL.n46 B 0.016578f
C355 VTAIL.n47 B 0.008908f
C356 VTAIL.n48 B 0.009432f
C357 VTAIL.n49 B 0.021056f
C358 VTAIL.n50 B 0.021056f
C359 VTAIL.n51 B 0.009432f
C360 VTAIL.n52 B 0.008908f
C361 VTAIL.n53 B 0.016578f
C362 VTAIL.n54 B 0.016578f
C363 VTAIL.n55 B 0.008908f
C364 VTAIL.n56 B 0.009432f
C365 VTAIL.n57 B 0.021056f
C366 VTAIL.n58 B 0.021056f
C367 VTAIL.n59 B 0.009432f
C368 VTAIL.n60 B 0.008908f
C369 VTAIL.n61 B 0.016578f
C370 VTAIL.n62 B 0.016578f
C371 VTAIL.n63 B 0.008908f
C372 VTAIL.n64 B 0.009432f
C373 VTAIL.n65 B 0.021056f
C374 VTAIL.n66 B 0.043389f
C375 VTAIL.n67 B 0.009432f
C376 VTAIL.n68 B 0.017419f
C377 VTAIL.n69 B 0.042396f
C378 VTAIL.n70 B 0.045201f
C379 VTAIL.n71 B 0.990543f
C380 VTAIL.n72 B 0.022966f
C381 VTAIL.n73 B 0.016578f
C382 VTAIL.n74 B 0.008908f
C383 VTAIL.n75 B 0.021056f
C384 VTAIL.n76 B 0.009432f
C385 VTAIL.n77 B 0.016578f
C386 VTAIL.n78 B 0.008908f
C387 VTAIL.n79 B 0.021056f
C388 VTAIL.n80 B 0.009432f
C389 VTAIL.n81 B 0.016578f
C390 VTAIL.n82 B 0.008908f
C391 VTAIL.n83 B 0.021056f
C392 VTAIL.n84 B 0.009432f
C393 VTAIL.n85 B 0.016578f
C394 VTAIL.n86 B 0.008908f
C395 VTAIL.n87 B 0.021056f
C396 VTAIL.n88 B 0.009432f
C397 VTAIL.n89 B 0.016578f
C398 VTAIL.n90 B 0.008908f
C399 VTAIL.n91 B 0.021056f
C400 VTAIL.n92 B 0.009432f
C401 VTAIL.n93 B 0.955502f
C402 VTAIL.n94 B 0.008908f
C403 VTAIL.t2 B 0.034626f
C404 VTAIL.n95 B 0.101391f
C405 VTAIL.n96 B 0.012438f
C406 VTAIL.n97 B 0.015792f
C407 VTAIL.n98 B 0.021056f
C408 VTAIL.n99 B 0.009432f
C409 VTAIL.n100 B 0.008908f
C410 VTAIL.n101 B 0.016578f
C411 VTAIL.n102 B 0.016578f
C412 VTAIL.n103 B 0.008908f
C413 VTAIL.n104 B 0.009432f
C414 VTAIL.n105 B 0.021056f
C415 VTAIL.n106 B 0.021056f
C416 VTAIL.n107 B 0.009432f
C417 VTAIL.n108 B 0.008908f
C418 VTAIL.n109 B 0.016578f
C419 VTAIL.n110 B 0.016578f
C420 VTAIL.n111 B 0.008908f
C421 VTAIL.n112 B 0.009432f
C422 VTAIL.n113 B 0.021056f
C423 VTAIL.n114 B 0.021056f
C424 VTAIL.n115 B 0.009432f
C425 VTAIL.n116 B 0.008908f
C426 VTAIL.n117 B 0.016578f
C427 VTAIL.n118 B 0.016578f
C428 VTAIL.n119 B 0.008908f
C429 VTAIL.n120 B 0.009432f
C430 VTAIL.n121 B 0.021056f
C431 VTAIL.n122 B 0.021056f
C432 VTAIL.n123 B 0.009432f
C433 VTAIL.n124 B 0.008908f
C434 VTAIL.n125 B 0.016578f
C435 VTAIL.n126 B 0.016578f
C436 VTAIL.n127 B 0.008908f
C437 VTAIL.n128 B 0.009432f
C438 VTAIL.n129 B 0.021056f
C439 VTAIL.n130 B 0.021056f
C440 VTAIL.n131 B 0.009432f
C441 VTAIL.n132 B 0.008908f
C442 VTAIL.n133 B 0.016578f
C443 VTAIL.n134 B 0.016578f
C444 VTAIL.n135 B 0.008908f
C445 VTAIL.n136 B 0.009432f
C446 VTAIL.n137 B 0.021056f
C447 VTAIL.n138 B 0.043389f
C448 VTAIL.n139 B 0.009432f
C449 VTAIL.n140 B 0.017419f
C450 VTAIL.n141 B 0.042396f
C451 VTAIL.n142 B 0.045201f
C452 VTAIL.n143 B 0.998947f
C453 VTAIL.n144 B 0.022966f
C454 VTAIL.n145 B 0.016578f
C455 VTAIL.n146 B 0.008908f
C456 VTAIL.n147 B 0.021056f
C457 VTAIL.n148 B 0.009432f
C458 VTAIL.n149 B 0.016578f
C459 VTAIL.n150 B 0.008908f
C460 VTAIL.n151 B 0.021056f
C461 VTAIL.n152 B 0.009432f
C462 VTAIL.n153 B 0.016578f
C463 VTAIL.n154 B 0.008908f
C464 VTAIL.n155 B 0.021056f
C465 VTAIL.n156 B 0.009432f
C466 VTAIL.n157 B 0.016578f
C467 VTAIL.n158 B 0.008908f
C468 VTAIL.n159 B 0.021056f
C469 VTAIL.n160 B 0.009432f
C470 VTAIL.n161 B 0.016578f
C471 VTAIL.n162 B 0.008908f
C472 VTAIL.n163 B 0.021056f
C473 VTAIL.n164 B 0.009432f
C474 VTAIL.n165 B 0.955502f
C475 VTAIL.n166 B 0.008908f
C476 VTAIL.t1 B 0.034626f
C477 VTAIL.n167 B 0.101391f
C478 VTAIL.n168 B 0.012438f
C479 VTAIL.n169 B 0.015792f
C480 VTAIL.n170 B 0.021056f
C481 VTAIL.n171 B 0.009432f
C482 VTAIL.n172 B 0.008908f
C483 VTAIL.n173 B 0.016578f
C484 VTAIL.n174 B 0.016578f
C485 VTAIL.n175 B 0.008908f
C486 VTAIL.n176 B 0.009432f
C487 VTAIL.n177 B 0.021056f
C488 VTAIL.n178 B 0.021056f
C489 VTAIL.n179 B 0.009432f
C490 VTAIL.n180 B 0.008908f
C491 VTAIL.n181 B 0.016578f
C492 VTAIL.n182 B 0.016578f
C493 VTAIL.n183 B 0.008908f
C494 VTAIL.n184 B 0.009432f
C495 VTAIL.n185 B 0.021056f
C496 VTAIL.n186 B 0.021056f
C497 VTAIL.n187 B 0.009432f
C498 VTAIL.n188 B 0.008908f
C499 VTAIL.n189 B 0.016578f
C500 VTAIL.n190 B 0.016578f
C501 VTAIL.n191 B 0.008908f
C502 VTAIL.n192 B 0.009432f
C503 VTAIL.n193 B 0.021056f
C504 VTAIL.n194 B 0.021056f
C505 VTAIL.n195 B 0.009432f
C506 VTAIL.n196 B 0.008908f
C507 VTAIL.n197 B 0.016578f
C508 VTAIL.n198 B 0.016578f
C509 VTAIL.n199 B 0.008908f
C510 VTAIL.n200 B 0.009432f
C511 VTAIL.n201 B 0.021056f
C512 VTAIL.n202 B 0.021056f
C513 VTAIL.n203 B 0.009432f
C514 VTAIL.n204 B 0.008908f
C515 VTAIL.n205 B 0.016578f
C516 VTAIL.n206 B 0.016578f
C517 VTAIL.n207 B 0.008908f
C518 VTAIL.n208 B 0.009432f
C519 VTAIL.n209 B 0.021056f
C520 VTAIL.n210 B 0.043389f
C521 VTAIL.n211 B 0.009432f
C522 VTAIL.n212 B 0.017419f
C523 VTAIL.n213 B 0.042396f
C524 VTAIL.n214 B 0.045201f
C525 VTAIL.n215 B 0.952897f
C526 VTAIL.n216 B 0.022966f
C527 VTAIL.n217 B 0.016578f
C528 VTAIL.n218 B 0.008908f
C529 VTAIL.n219 B 0.021056f
C530 VTAIL.n220 B 0.009432f
C531 VTAIL.n221 B 0.016578f
C532 VTAIL.n222 B 0.008908f
C533 VTAIL.n223 B 0.021056f
C534 VTAIL.n224 B 0.009432f
C535 VTAIL.n225 B 0.016578f
C536 VTAIL.n226 B 0.008908f
C537 VTAIL.n227 B 0.021056f
C538 VTAIL.n228 B 0.009432f
C539 VTAIL.n229 B 0.016578f
C540 VTAIL.n230 B 0.008908f
C541 VTAIL.n231 B 0.021056f
C542 VTAIL.n232 B 0.009432f
C543 VTAIL.n233 B 0.016578f
C544 VTAIL.n234 B 0.008908f
C545 VTAIL.n235 B 0.021056f
C546 VTAIL.n236 B 0.009432f
C547 VTAIL.n237 B 0.955502f
C548 VTAIL.n238 B 0.008908f
C549 VTAIL.t3 B 0.034626f
C550 VTAIL.n239 B 0.101391f
C551 VTAIL.n240 B 0.012438f
C552 VTAIL.n241 B 0.015792f
C553 VTAIL.n242 B 0.021056f
C554 VTAIL.n243 B 0.009432f
C555 VTAIL.n244 B 0.008908f
C556 VTAIL.n245 B 0.016578f
C557 VTAIL.n246 B 0.016578f
C558 VTAIL.n247 B 0.008908f
C559 VTAIL.n248 B 0.009432f
C560 VTAIL.n249 B 0.021056f
C561 VTAIL.n250 B 0.021056f
C562 VTAIL.n251 B 0.009432f
C563 VTAIL.n252 B 0.008908f
C564 VTAIL.n253 B 0.016578f
C565 VTAIL.n254 B 0.016578f
C566 VTAIL.n255 B 0.008908f
C567 VTAIL.n256 B 0.009432f
C568 VTAIL.n257 B 0.021056f
C569 VTAIL.n258 B 0.021056f
C570 VTAIL.n259 B 0.009432f
C571 VTAIL.n260 B 0.008908f
C572 VTAIL.n261 B 0.016578f
C573 VTAIL.n262 B 0.016578f
C574 VTAIL.n263 B 0.008908f
C575 VTAIL.n264 B 0.009432f
C576 VTAIL.n265 B 0.021056f
C577 VTAIL.n266 B 0.021056f
C578 VTAIL.n267 B 0.009432f
C579 VTAIL.n268 B 0.008908f
C580 VTAIL.n269 B 0.016578f
C581 VTAIL.n270 B 0.016578f
C582 VTAIL.n271 B 0.008908f
C583 VTAIL.n272 B 0.009432f
C584 VTAIL.n273 B 0.021056f
C585 VTAIL.n274 B 0.021056f
C586 VTAIL.n275 B 0.009432f
C587 VTAIL.n276 B 0.008908f
C588 VTAIL.n277 B 0.016578f
C589 VTAIL.n278 B 0.016578f
C590 VTAIL.n279 B 0.008908f
C591 VTAIL.n280 B 0.009432f
C592 VTAIL.n281 B 0.021056f
C593 VTAIL.n282 B 0.043389f
C594 VTAIL.n283 B 0.009432f
C595 VTAIL.n284 B 0.017419f
C596 VTAIL.n285 B 0.042396f
C597 VTAIL.n286 B 0.045201f
C598 VTAIL.n287 B 0.913179f
C599 VN.t1 B 1.28659f
C600 VN.t0 B 1.4074f
.ends

