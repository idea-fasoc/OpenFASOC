* NGSPICE file created from diff_pair_sample_0795.ext - technology: sky130A

.subckt diff_pair_sample_0795 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
X1 VTAIL.t12 VP.t1 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
X2 VTAIL.t6 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=1.68
X3 VDD1.t5 VP.t2 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=1.68
X4 B.t20 B.t18 B.t19 B.t15 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=1.68
X5 VTAIL.t13 VP.t3 VDD1.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=1.68
X6 VDD1.t3 VP.t4 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=1.68
X7 VTAIL.t10 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
X8 VDD1.t1 VP.t6 VTAIL.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
X9 VDD2.t6 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=1.68
X10 VTAIL.t1 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
X11 VDD2.t4 VN.t3 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=6.4155 ps=33.68 w=16.45 l=1.68
X12 VTAIL.t4 VN.t4 VDD2.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
X13 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=1.68
X14 VTAIL.t11 VP.t7 VDD1.t0 B.t21 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=1.68
X15 VDD2.t2 VN.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
X16 VTAIL.t15 VN.t6 VDD2.t1 B.t21 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=2.71425 ps=16.78 w=16.45 l=1.68
X17 B.t13 B.t11 B.t12 B.t8 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=1.68
X18 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=6.4155 pd=33.68 as=0 ps=0 w=16.45 l=1.68
X19 VDD2.t0 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.71425 pd=16.78 as=2.71425 ps=16.78 w=16.45 l=1.68
R0 VP.n12 VP.t7 263.481
R1 VP.n31 VP.t3 235.98
R2 VP.n38 VP.t6 235.98
R3 VP.n46 VP.t5 235.98
R4 VP.n53 VP.t4 235.98
R5 VP.n28 VP.t2 235.98
R6 VP.n21 VP.t1 235.98
R7 VP.n13 VP.t0 235.98
R8 VP.n31 VP.n30 185.034
R9 VP.n54 VP.n53 185.034
R10 VP.n29 VP.n28 185.034
R11 VP.n14 VP.n11 161.3
R12 VP.n16 VP.n15 161.3
R13 VP.n17 VP.n10 161.3
R14 VP.n19 VP.n18 161.3
R15 VP.n20 VP.n9 161.3
R16 VP.n23 VP.n22 161.3
R17 VP.n24 VP.n8 161.3
R18 VP.n26 VP.n25 161.3
R19 VP.n27 VP.n7 161.3
R20 VP.n52 VP.n0 161.3
R21 VP.n51 VP.n50 161.3
R22 VP.n49 VP.n1 161.3
R23 VP.n48 VP.n47 161.3
R24 VP.n45 VP.n2 161.3
R25 VP.n44 VP.n43 161.3
R26 VP.n42 VP.n3 161.3
R27 VP.n41 VP.n40 161.3
R28 VP.n39 VP.n4 161.3
R29 VP.n37 VP.n36 161.3
R30 VP.n35 VP.n5 161.3
R31 VP.n34 VP.n33 161.3
R32 VP.n32 VP.n6 161.3
R33 VP.n13 VP.n12 68.7155
R34 VP.n30 VP.n29 49.7884
R35 VP.n33 VP.n5 41.4647
R36 VP.n51 VP.n1 41.4647
R37 VP.n26 VP.n8 41.4647
R38 VP.n40 VP.n3 40.4934
R39 VP.n44 VP.n3 40.4934
R40 VP.n19 VP.n10 40.4934
R41 VP.n15 VP.n10 40.4934
R42 VP.n37 VP.n5 39.5221
R43 VP.n47 VP.n1 39.5221
R44 VP.n22 VP.n8 39.5221
R45 VP.n33 VP.n32 24.4675
R46 VP.n40 VP.n39 24.4675
R47 VP.n45 VP.n44 24.4675
R48 VP.n52 VP.n51 24.4675
R49 VP.n27 VP.n26 24.4675
R50 VP.n20 VP.n19 24.4675
R51 VP.n15 VP.n14 24.4675
R52 VP.n38 VP.n37 24.2228
R53 VP.n47 VP.n46 24.2228
R54 VP.n22 VP.n21 24.2228
R55 VP.n12 VP.n11 18.9997
R56 VP.n32 VP.n31 0.73451
R57 VP.n53 VP.n52 0.73451
R58 VP.n28 VP.n27 0.73451
R59 VP.n39 VP.n38 0.24517
R60 VP.n46 VP.n45 0.24517
R61 VP.n21 VP.n20 0.24517
R62 VP.n14 VP.n13 0.24517
R63 VP.n16 VP.n11 0.189894
R64 VP.n17 VP.n16 0.189894
R65 VP.n18 VP.n17 0.189894
R66 VP.n18 VP.n9 0.189894
R67 VP.n23 VP.n9 0.189894
R68 VP.n24 VP.n23 0.189894
R69 VP.n25 VP.n24 0.189894
R70 VP.n25 VP.n7 0.189894
R71 VP.n29 VP.n7 0.189894
R72 VP.n30 VP.n6 0.189894
R73 VP.n34 VP.n6 0.189894
R74 VP.n35 VP.n34 0.189894
R75 VP.n36 VP.n35 0.189894
R76 VP.n36 VP.n4 0.189894
R77 VP.n41 VP.n4 0.189894
R78 VP.n42 VP.n41 0.189894
R79 VP.n43 VP.n42 0.189894
R80 VP.n43 VP.n2 0.189894
R81 VP.n48 VP.n2 0.189894
R82 VP.n49 VP.n48 0.189894
R83 VP.n50 VP.n49 0.189894
R84 VP.n50 VP.n0 0.189894
R85 VP.n54 VP.n0 0.189894
R86 VP VP.n54 0.0516364
R87 VTAIL.n11 VTAIL.t11 45.4684
R88 VTAIL.n10 VTAIL.t0 45.4684
R89 VTAIL.n7 VTAIL.t6 45.4684
R90 VTAIL.n14 VTAIL.t7 45.4682
R91 VTAIL.n15 VTAIL.t3 45.4682
R92 VTAIL.n2 VTAIL.t15 45.4682
R93 VTAIL.n3 VTAIL.t14 45.4682
R94 VTAIL.n6 VTAIL.t13 45.4682
R95 VTAIL.n13 VTAIL.n12 44.2648
R96 VTAIL.n9 VTAIL.n8 44.2648
R97 VTAIL.n1 VTAIL.n0 44.2646
R98 VTAIL.n5 VTAIL.n4 44.2646
R99 VTAIL.n15 VTAIL.n14 28.2807
R100 VTAIL.n7 VTAIL.n6 28.2807
R101 VTAIL.n9 VTAIL.n7 1.73326
R102 VTAIL.n10 VTAIL.n9 1.73326
R103 VTAIL.n13 VTAIL.n11 1.73326
R104 VTAIL.n14 VTAIL.n13 1.73326
R105 VTAIL.n6 VTAIL.n5 1.73326
R106 VTAIL.n5 VTAIL.n3 1.73326
R107 VTAIL.n2 VTAIL.n1 1.73326
R108 VTAIL VTAIL.n15 1.67507
R109 VTAIL.n0 VTAIL.t2 1.20415
R110 VTAIL.n0 VTAIL.t1 1.20415
R111 VTAIL.n4 VTAIL.t8 1.20415
R112 VTAIL.n4 VTAIL.t10 1.20415
R113 VTAIL.n12 VTAIL.t9 1.20415
R114 VTAIL.n12 VTAIL.t12 1.20415
R115 VTAIL.n8 VTAIL.t5 1.20415
R116 VTAIL.n8 VTAIL.t4 1.20415
R117 VTAIL.n11 VTAIL.n10 0.470328
R118 VTAIL.n3 VTAIL.n2 0.470328
R119 VTAIL VTAIL.n1 0.0586897
R120 VDD1 VDD1.n0 61.8681
R121 VDD1.n3 VDD1.n2 61.7544
R122 VDD1.n3 VDD1.n1 61.7544
R123 VDD1.n5 VDD1.n4 60.9434
R124 VDD1.n5 VDD1.n3 46.2768
R125 VDD1.n4 VDD1.t6 1.20415
R126 VDD1.n4 VDD1.t5 1.20415
R127 VDD1.n0 VDD1.t0 1.20415
R128 VDD1.n0 VDD1.t7 1.20415
R129 VDD1.n2 VDD1.t2 1.20415
R130 VDD1.n2 VDD1.t3 1.20415
R131 VDD1.n1 VDD1.t4 1.20415
R132 VDD1.n1 VDD1.t1 1.20415
R133 VDD1 VDD1.n5 0.80869
R134 B.n908 B.n907 585
R135 B.n909 B.n908 585
R136 B.n371 B.n130 585
R137 B.n370 B.n369 585
R138 B.n368 B.n367 585
R139 B.n366 B.n365 585
R140 B.n364 B.n363 585
R141 B.n362 B.n361 585
R142 B.n360 B.n359 585
R143 B.n358 B.n357 585
R144 B.n356 B.n355 585
R145 B.n354 B.n353 585
R146 B.n352 B.n351 585
R147 B.n350 B.n349 585
R148 B.n348 B.n347 585
R149 B.n346 B.n345 585
R150 B.n344 B.n343 585
R151 B.n342 B.n341 585
R152 B.n340 B.n339 585
R153 B.n338 B.n337 585
R154 B.n336 B.n335 585
R155 B.n334 B.n333 585
R156 B.n332 B.n331 585
R157 B.n330 B.n329 585
R158 B.n328 B.n327 585
R159 B.n326 B.n325 585
R160 B.n324 B.n323 585
R161 B.n322 B.n321 585
R162 B.n320 B.n319 585
R163 B.n318 B.n317 585
R164 B.n316 B.n315 585
R165 B.n314 B.n313 585
R166 B.n312 B.n311 585
R167 B.n310 B.n309 585
R168 B.n308 B.n307 585
R169 B.n306 B.n305 585
R170 B.n304 B.n303 585
R171 B.n302 B.n301 585
R172 B.n300 B.n299 585
R173 B.n298 B.n297 585
R174 B.n296 B.n295 585
R175 B.n294 B.n293 585
R176 B.n292 B.n291 585
R177 B.n290 B.n289 585
R178 B.n288 B.n287 585
R179 B.n286 B.n285 585
R180 B.n284 B.n283 585
R181 B.n282 B.n281 585
R182 B.n280 B.n279 585
R183 B.n278 B.n277 585
R184 B.n276 B.n275 585
R185 B.n274 B.n273 585
R186 B.n272 B.n271 585
R187 B.n270 B.n269 585
R188 B.n268 B.n267 585
R189 B.n266 B.n265 585
R190 B.n264 B.n263 585
R191 B.n262 B.n261 585
R192 B.n260 B.n259 585
R193 B.n258 B.n257 585
R194 B.n256 B.n255 585
R195 B.n254 B.n253 585
R196 B.n252 B.n251 585
R197 B.n250 B.n249 585
R198 B.n248 B.n247 585
R199 B.n245 B.n244 585
R200 B.n243 B.n242 585
R201 B.n241 B.n240 585
R202 B.n239 B.n238 585
R203 B.n237 B.n236 585
R204 B.n235 B.n234 585
R205 B.n233 B.n232 585
R206 B.n231 B.n230 585
R207 B.n229 B.n228 585
R208 B.n227 B.n226 585
R209 B.n225 B.n224 585
R210 B.n223 B.n222 585
R211 B.n221 B.n220 585
R212 B.n219 B.n218 585
R213 B.n217 B.n216 585
R214 B.n215 B.n214 585
R215 B.n213 B.n212 585
R216 B.n211 B.n210 585
R217 B.n209 B.n208 585
R218 B.n207 B.n206 585
R219 B.n205 B.n204 585
R220 B.n203 B.n202 585
R221 B.n201 B.n200 585
R222 B.n199 B.n198 585
R223 B.n197 B.n196 585
R224 B.n195 B.n194 585
R225 B.n193 B.n192 585
R226 B.n191 B.n190 585
R227 B.n189 B.n188 585
R228 B.n187 B.n186 585
R229 B.n185 B.n184 585
R230 B.n183 B.n182 585
R231 B.n181 B.n180 585
R232 B.n179 B.n178 585
R233 B.n177 B.n176 585
R234 B.n175 B.n174 585
R235 B.n173 B.n172 585
R236 B.n171 B.n170 585
R237 B.n169 B.n168 585
R238 B.n167 B.n166 585
R239 B.n165 B.n164 585
R240 B.n163 B.n162 585
R241 B.n161 B.n160 585
R242 B.n159 B.n158 585
R243 B.n157 B.n156 585
R244 B.n155 B.n154 585
R245 B.n153 B.n152 585
R246 B.n151 B.n150 585
R247 B.n149 B.n148 585
R248 B.n147 B.n146 585
R249 B.n145 B.n144 585
R250 B.n143 B.n142 585
R251 B.n141 B.n140 585
R252 B.n139 B.n138 585
R253 B.n137 B.n136 585
R254 B.n906 B.n70 585
R255 B.n910 B.n70 585
R256 B.n905 B.n69 585
R257 B.n911 B.n69 585
R258 B.n904 B.n903 585
R259 B.n903 B.n65 585
R260 B.n902 B.n64 585
R261 B.n917 B.n64 585
R262 B.n901 B.n63 585
R263 B.n918 B.n63 585
R264 B.n900 B.n62 585
R265 B.n919 B.n62 585
R266 B.n899 B.n898 585
R267 B.n898 B.n61 585
R268 B.n897 B.n57 585
R269 B.n925 B.n57 585
R270 B.n896 B.n56 585
R271 B.n926 B.n56 585
R272 B.n895 B.n55 585
R273 B.n927 B.n55 585
R274 B.n894 B.n893 585
R275 B.n893 B.n51 585
R276 B.n892 B.n50 585
R277 B.n933 B.n50 585
R278 B.n891 B.n49 585
R279 B.n934 B.n49 585
R280 B.n890 B.n48 585
R281 B.n935 B.n48 585
R282 B.n889 B.n888 585
R283 B.n888 B.n44 585
R284 B.n887 B.n43 585
R285 B.n941 B.n43 585
R286 B.n886 B.n42 585
R287 B.n942 B.n42 585
R288 B.n885 B.n41 585
R289 B.n943 B.n41 585
R290 B.n884 B.n883 585
R291 B.n883 B.n37 585
R292 B.n882 B.n36 585
R293 B.n949 B.n36 585
R294 B.n881 B.n35 585
R295 B.n950 B.n35 585
R296 B.n880 B.n34 585
R297 B.n951 B.n34 585
R298 B.n879 B.n878 585
R299 B.n878 B.n30 585
R300 B.n877 B.n29 585
R301 B.n957 B.n29 585
R302 B.n876 B.n28 585
R303 B.n958 B.n28 585
R304 B.n875 B.n27 585
R305 B.n959 B.n27 585
R306 B.n874 B.n873 585
R307 B.n873 B.n23 585
R308 B.n872 B.n22 585
R309 B.n965 B.n22 585
R310 B.n871 B.n21 585
R311 B.n966 B.n21 585
R312 B.n870 B.n20 585
R313 B.n967 B.n20 585
R314 B.n869 B.n868 585
R315 B.n868 B.n16 585
R316 B.n867 B.n15 585
R317 B.n973 B.n15 585
R318 B.n866 B.n14 585
R319 B.n974 B.n14 585
R320 B.n865 B.n13 585
R321 B.n975 B.n13 585
R322 B.n864 B.n863 585
R323 B.n863 B.n12 585
R324 B.n862 B.n861 585
R325 B.n862 B.n8 585
R326 B.n860 B.n7 585
R327 B.n982 B.n7 585
R328 B.n859 B.n6 585
R329 B.n983 B.n6 585
R330 B.n858 B.n5 585
R331 B.n984 B.n5 585
R332 B.n857 B.n856 585
R333 B.n856 B.n4 585
R334 B.n855 B.n372 585
R335 B.n855 B.n854 585
R336 B.n845 B.n373 585
R337 B.n374 B.n373 585
R338 B.n847 B.n846 585
R339 B.n848 B.n847 585
R340 B.n844 B.n378 585
R341 B.n382 B.n378 585
R342 B.n843 B.n842 585
R343 B.n842 B.n841 585
R344 B.n380 B.n379 585
R345 B.n381 B.n380 585
R346 B.n834 B.n833 585
R347 B.n835 B.n834 585
R348 B.n832 B.n387 585
R349 B.n387 B.n386 585
R350 B.n831 B.n830 585
R351 B.n830 B.n829 585
R352 B.n389 B.n388 585
R353 B.n390 B.n389 585
R354 B.n822 B.n821 585
R355 B.n823 B.n822 585
R356 B.n820 B.n395 585
R357 B.n395 B.n394 585
R358 B.n819 B.n818 585
R359 B.n818 B.n817 585
R360 B.n397 B.n396 585
R361 B.n398 B.n397 585
R362 B.n810 B.n809 585
R363 B.n811 B.n810 585
R364 B.n808 B.n403 585
R365 B.n403 B.n402 585
R366 B.n807 B.n806 585
R367 B.n806 B.n805 585
R368 B.n405 B.n404 585
R369 B.n406 B.n405 585
R370 B.n798 B.n797 585
R371 B.n799 B.n798 585
R372 B.n796 B.n411 585
R373 B.n411 B.n410 585
R374 B.n795 B.n794 585
R375 B.n794 B.n793 585
R376 B.n413 B.n412 585
R377 B.n414 B.n413 585
R378 B.n786 B.n785 585
R379 B.n787 B.n786 585
R380 B.n784 B.n419 585
R381 B.n419 B.n418 585
R382 B.n783 B.n782 585
R383 B.n782 B.n781 585
R384 B.n421 B.n420 585
R385 B.n422 B.n421 585
R386 B.n774 B.n773 585
R387 B.n775 B.n774 585
R388 B.n772 B.n427 585
R389 B.n427 B.n426 585
R390 B.n771 B.n770 585
R391 B.n770 B.n769 585
R392 B.n429 B.n428 585
R393 B.n762 B.n429 585
R394 B.n761 B.n760 585
R395 B.n763 B.n761 585
R396 B.n759 B.n434 585
R397 B.n434 B.n433 585
R398 B.n758 B.n757 585
R399 B.n757 B.n756 585
R400 B.n436 B.n435 585
R401 B.n437 B.n436 585
R402 B.n749 B.n748 585
R403 B.n750 B.n749 585
R404 B.n747 B.n442 585
R405 B.n442 B.n441 585
R406 B.n741 B.n740 585
R407 B.n739 B.n503 585
R408 B.n738 B.n502 585
R409 B.n743 B.n502 585
R410 B.n737 B.n736 585
R411 B.n735 B.n734 585
R412 B.n733 B.n732 585
R413 B.n731 B.n730 585
R414 B.n729 B.n728 585
R415 B.n727 B.n726 585
R416 B.n725 B.n724 585
R417 B.n723 B.n722 585
R418 B.n721 B.n720 585
R419 B.n719 B.n718 585
R420 B.n717 B.n716 585
R421 B.n715 B.n714 585
R422 B.n713 B.n712 585
R423 B.n711 B.n710 585
R424 B.n709 B.n708 585
R425 B.n707 B.n706 585
R426 B.n705 B.n704 585
R427 B.n703 B.n702 585
R428 B.n701 B.n700 585
R429 B.n699 B.n698 585
R430 B.n697 B.n696 585
R431 B.n695 B.n694 585
R432 B.n693 B.n692 585
R433 B.n691 B.n690 585
R434 B.n689 B.n688 585
R435 B.n687 B.n686 585
R436 B.n685 B.n684 585
R437 B.n683 B.n682 585
R438 B.n681 B.n680 585
R439 B.n679 B.n678 585
R440 B.n677 B.n676 585
R441 B.n675 B.n674 585
R442 B.n673 B.n672 585
R443 B.n671 B.n670 585
R444 B.n669 B.n668 585
R445 B.n667 B.n666 585
R446 B.n665 B.n664 585
R447 B.n663 B.n662 585
R448 B.n661 B.n660 585
R449 B.n659 B.n658 585
R450 B.n657 B.n656 585
R451 B.n655 B.n654 585
R452 B.n653 B.n652 585
R453 B.n651 B.n650 585
R454 B.n649 B.n648 585
R455 B.n647 B.n646 585
R456 B.n645 B.n644 585
R457 B.n643 B.n642 585
R458 B.n641 B.n640 585
R459 B.n639 B.n638 585
R460 B.n637 B.n636 585
R461 B.n635 B.n634 585
R462 B.n633 B.n632 585
R463 B.n631 B.n630 585
R464 B.n629 B.n628 585
R465 B.n627 B.n626 585
R466 B.n625 B.n624 585
R467 B.n623 B.n622 585
R468 B.n621 B.n620 585
R469 B.n619 B.n618 585
R470 B.n617 B.n616 585
R471 B.n614 B.n613 585
R472 B.n612 B.n611 585
R473 B.n610 B.n609 585
R474 B.n608 B.n607 585
R475 B.n606 B.n605 585
R476 B.n604 B.n603 585
R477 B.n602 B.n601 585
R478 B.n600 B.n599 585
R479 B.n598 B.n597 585
R480 B.n596 B.n595 585
R481 B.n594 B.n593 585
R482 B.n592 B.n591 585
R483 B.n590 B.n589 585
R484 B.n588 B.n587 585
R485 B.n586 B.n585 585
R486 B.n584 B.n583 585
R487 B.n582 B.n581 585
R488 B.n580 B.n579 585
R489 B.n578 B.n577 585
R490 B.n576 B.n575 585
R491 B.n574 B.n573 585
R492 B.n572 B.n571 585
R493 B.n570 B.n569 585
R494 B.n568 B.n567 585
R495 B.n566 B.n565 585
R496 B.n564 B.n563 585
R497 B.n562 B.n561 585
R498 B.n560 B.n559 585
R499 B.n558 B.n557 585
R500 B.n556 B.n555 585
R501 B.n554 B.n553 585
R502 B.n552 B.n551 585
R503 B.n550 B.n549 585
R504 B.n548 B.n547 585
R505 B.n546 B.n545 585
R506 B.n544 B.n543 585
R507 B.n542 B.n541 585
R508 B.n540 B.n539 585
R509 B.n538 B.n537 585
R510 B.n536 B.n535 585
R511 B.n534 B.n533 585
R512 B.n532 B.n531 585
R513 B.n530 B.n529 585
R514 B.n528 B.n527 585
R515 B.n526 B.n525 585
R516 B.n524 B.n523 585
R517 B.n522 B.n521 585
R518 B.n520 B.n519 585
R519 B.n518 B.n517 585
R520 B.n516 B.n515 585
R521 B.n514 B.n513 585
R522 B.n512 B.n511 585
R523 B.n510 B.n509 585
R524 B.n444 B.n443 585
R525 B.n746 B.n745 585
R526 B.n440 B.n439 585
R527 B.n441 B.n440 585
R528 B.n752 B.n751 585
R529 B.n751 B.n750 585
R530 B.n753 B.n438 585
R531 B.n438 B.n437 585
R532 B.n755 B.n754 585
R533 B.n756 B.n755 585
R534 B.n432 B.n431 585
R535 B.n433 B.n432 585
R536 B.n765 B.n764 585
R537 B.n764 B.n763 585
R538 B.n766 B.n430 585
R539 B.n762 B.n430 585
R540 B.n768 B.n767 585
R541 B.n769 B.n768 585
R542 B.n425 B.n424 585
R543 B.n426 B.n425 585
R544 B.n777 B.n776 585
R545 B.n776 B.n775 585
R546 B.n778 B.n423 585
R547 B.n423 B.n422 585
R548 B.n780 B.n779 585
R549 B.n781 B.n780 585
R550 B.n417 B.n416 585
R551 B.n418 B.n417 585
R552 B.n789 B.n788 585
R553 B.n788 B.n787 585
R554 B.n790 B.n415 585
R555 B.n415 B.n414 585
R556 B.n792 B.n791 585
R557 B.n793 B.n792 585
R558 B.n409 B.n408 585
R559 B.n410 B.n409 585
R560 B.n801 B.n800 585
R561 B.n800 B.n799 585
R562 B.n802 B.n407 585
R563 B.n407 B.n406 585
R564 B.n804 B.n803 585
R565 B.n805 B.n804 585
R566 B.n401 B.n400 585
R567 B.n402 B.n401 585
R568 B.n813 B.n812 585
R569 B.n812 B.n811 585
R570 B.n814 B.n399 585
R571 B.n399 B.n398 585
R572 B.n816 B.n815 585
R573 B.n817 B.n816 585
R574 B.n393 B.n392 585
R575 B.n394 B.n393 585
R576 B.n825 B.n824 585
R577 B.n824 B.n823 585
R578 B.n826 B.n391 585
R579 B.n391 B.n390 585
R580 B.n828 B.n827 585
R581 B.n829 B.n828 585
R582 B.n385 B.n384 585
R583 B.n386 B.n385 585
R584 B.n837 B.n836 585
R585 B.n836 B.n835 585
R586 B.n838 B.n383 585
R587 B.n383 B.n381 585
R588 B.n840 B.n839 585
R589 B.n841 B.n840 585
R590 B.n377 B.n376 585
R591 B.n382 B.n377 585
R592 B.n850 B.n849 585
R593 B.n849 B.n848 585
R594 B.n851 B.n375 585
R595 B.n375 B.n374 585
R596 B.n853 B.n852 585
R597 B.n854 B.n853 585
R598 B.n3 B.n0 585
R599 B.n4 B.n3 585
R600 B.n981 B.n1 585
R601 B.n982 B.n981 585
R602 B.n980 B.n979 585
R603 B.n980 B.n8 585
R604 B.n978 B.n9 585
R605 B.n12 B.n9 585
R606 B.n977 B.n976 585
R607 B.n976 B.n975 585
R608 B.n11 B.n10 585
R609 B.n974 B.n11 585
R610 B.n972 B.n971 585
R611 B.n973 B.n972 585
R612 B.n970 B.n17 585
R613 B.n17 B.n16 585
R614 B.n969 B.n968 585
R615 B.n968 B.n967 585
R616 B.n19 B.n18 585
R617 B.n966 B.n19 585
R618 B.n964 B.n963 585
R619 B.n965 B.n964 585
R620 B.n962 B.n24 585
R621 B.n24 B.n23 585
R622 B.n961 B.n960 585
R623 B.n960 B.n959 585
R624 B.n26 B.n25 585
R625 B.n958 B.n26 585
R626 B.n956 B.n955 585
R627 B.n957 B.n956 585
R628 B.n954 B.n31 585
R629 B.n31 B.n30 585
R630 B.n953 B.n952 585
R631 B.n952 B.n951 585
R632 B.n33 B.n32 585
R633 B.n950 B.n33 585
R634 B.n948 B.n947 585
R635 B.n949 B.n948 585
R636 B.n946 B.n38 585
R637 B.n38 B.n37 585
R638 B.n945 B.n944 585
R639 B.n944 B.n943 585
R640 B.n40 B.n39 585
R641 B.n942 B.n40 585
R642 B.n940 B.n939 585
R643 B.n941 B.n940 585
R644 B.n938 B.n45 585
R645 B.n45 B.n44 585
R646 B.n937 B.n936 585
R647 B.n936 B.n935 585
R648 B.n47 B.n46 585
R649 B.n934 B.n47 585
R650 B.n932 B.n931 585
R651 B.n933 B.n932 585
R652 B.n930 B.n52 585
R653 B.n52 B.n51 585
R654 B.n929 B.n928 585
R655 B.n928 B.n927 585
R656 B.n54 B.n53 585
R657 B.n926 B.n54 585
R658 B.n924 B.n923 585
R659 B.n925 B.n924 585
R660 B.n922 B.n58 585
R661 B.n61 B.n58 585
R662 B.n921 B.n920 585
R663 B.n920 B.n919 585
R664 B.n60 B.n59 585
R665 B.n918 B.n60 585
R666 B.n916 B.n915 585
R667 B.n917 B.n916 585
R668 B.n914 B.n66 585
R669 B.n66 B.n65 585
R670 B.n913 B.n912 585
R671 B.n912 B.n911 585
R672 B.n68 B.n67 585
R673 B.n910 B.n68 585
R674 B.n985 B.n984 585
R675 B.n983 B.n2 585
R676 B.n136 B.n68 526.135
R677 B.n908 B.n70 526.135
R678 B.n745 B.n442 526.135
R679 B.n741 B.n440 526.135
R680 B.n134 B.t11 442.031
R681 B.n131 B.t7 442.031
R682 B.n507 B.t18 442.031
R683 B.n504 B.t14 442.031
R684 B.n909 B.n129 256.663
R685 B.n909 B.n128 256.663
R686 B.n909 B.n127 256.663
R687 B.n909 B.n126 256.663
R688 B.n909 B.n125 256.663
R689 B.n909 B.n124 256.663
R690 B.n909 B.n123 256.663
R691 B.n909 B.n122 256.663
R692 B.n909 B.n121 256.663
R693 B.n909 B.n120 256.663
R694 B.n909 B.n119 256.663
R695 B.n909 B.n118 256.663
R696 B.n909 B.n117 256.663
R697 B.n909 B.n116 256.663
R698 B.n909 B.n115 256.663
R699 B.n909 B.n114 256.663
R700 B.n909 B.n113 256.663
R701 B.n909 B.n112 256.663
R702 B.n909 B.n111 256.663
R703 B.n909 B.n110 256.663
R704 B.n909 B.n109 256.663
R705 B.n909 B.n108 256.663
R706 B.n909 B.n107 256.663
R707 B.n909 B.n106 256.663
R708 B.n909 B.n105 256.663
R709 B.n909 B.n104 256.663
R710 B.n909 B.n103 256.663
R711 B.n909 B.n102 256.663
R712 B.n909 B.n101 256.663
R713 B.n909 B.n100 256.663
R714 B.n909 B.n99 256.663
R715 B.n909 B.n98 256.663
R716 B.n909 B.n97 256.663
R717 B.n909 B.n96 256.663
R718 B.n909 B.n95 256.663
R719 B.n909 B.n94 256.663
R720 B.n909 B.n93 256.663
R721 B.n909 B.n92 256.663
R722 B.n909 B.n91 256.663
R723 B.n909 B.n90 256.663
R724 B.n909 B.n89 256.663
R725 B.n909 B.n88 256.663
R726 B.n909 B.n87 256.663
R727 B.n909 B.n86 256.663
R728 B.n909 B.n85 256.663
R729 B.n909 B.n84 256.663
R730 B.n909 B.n83 256.663
R731 B.n909 B.n82 256.663
R732 B.n909 B.n81 256.663
R733 B.n909 B.n80 256.663
R734 B.n909 B.n79 256.663
R735 B.n909 B.n78 256.663
R736 B.n909 B.n77 256.663
R737 B.n909 B.n76 256.663
R738 B.n909 B.n75 256.663
R739 B.n909 B.n74 256.663
R740 B.n909 B.n73 256.663
R741 B.n909 B.n72 256.663
R742 B.n909 B.n71 256.663
R743 B.n743 B.n742 256.663
R744 B.n743 B.n445 256.663
R745 B.n743 B.n446 256.663
R746 B.n743 B.n447 256.663
R747 B.n743 B.n448 256.663
R748 B.n743 B.n449 256.663
R749 B.n743 B.n450 256.663
R750 B.n743 B.n451 256.663
R751 B.n743 B.n452 256.663
R752 B.n743 B.n453 256.663
R753 B.n743 B.n454 256.663
R754 B.n743 B.n455 256.663
R755 B.n743 B.n456 256.663
R756 B.n743 B.n457 256.663
R757 B.n743 B.n458 256.663
R758 B.n743 B.n459 256.663
R759 B.n743 B.n460 256.663
R760 B.n743 B.n461 256.663
R761 B.n743 B.n462 256.663
R762 B.n743 B.n463 256.663
R763 B.n743 B.n464 256.663
R764 B.n743 B.n465 256.663
R765 B.n743 B.n466 256.663
R766 B.n743 B.n467 256.663
R767 B.n743 B.n468 256.663
R768 B.n743 B.n469 256.663
R769 B.n743 B.n470 256.663
R770 B.n743 B.n471 256.663
R771 B.n743 B.n472 256.663
R772 B.n743 B.n473 256.663
R773 B.n743 B.n474 256.663
R774 B.n743 B.n475 256.663
R775 B.n743 B.n476 256.663
R776 B.n743 B.n477 256.663
R777 B.n743 B.n478 256.663
R778 B.n743 B.n479 256.663
R779 B.n743 B.n480 256.663
R780 B.n743 B.n481 256.663
R781 B.n743 B.n482 256.663
R782 B.n743 B.n483 256.663
R783 B.n743 B.n484 256.663
R784 B.n743 B.n485 256.663
R785 B.n743 B.n486 256.663
R786 B.n743 B.n487 256.663
R787 B.n743 B.n488 256.663
R788 B.n743 B.n489 256.663
R789 B.n743 B.n490 256.663
R790 B.n743 B.n491 256.663
R791 B.n743 B.n492 256.663
R792 B.n743 B.n493 256.663
R793 B.n743 B.n494 256.663
R794 B.n743 B.n495 256.663
R795 B.n743 B.n496 256.663
R796 B.n743 B.n497 256.663
R797 B.n743 B.n498 256.663
R798 B.n743 B.n499 256.663
R799 B.n743 B.n500 256.663
R800 B.n743 B.n501 256.663
R801 B.n744 B.n743 256.663
R802 B.n987 B.n986 256.663
R803 B.n140 B.n139 163.367
R804 B.n144 B.n143 163.367
R805 B.n148 B.n147 163.367
R806 B.n152 B.n151 163.367
R807 B.n156 B.n155 163.367
R808 B.n160 B.n159 163.367
R809 B.n164 B.n163 163.367
R810 B.n168 B.n167 163.367
R811 B.n172 B.n171 163.367
R812 B.n176 B.n175 163.367
R813 B.n180 B.n179 163.367
R814 B.n184 B.n183 163.367
R815 B.n188 B.n187 163.367
R816 B.n192 B.n191 163.367
R817 B.n196 B.n195 163.367
R818 B.n200 B.n199 163.367
R819 B.n204 B.n203 163.367
R820 B.n208 B.n207 163.367
R821 B.n212 B.n211 163.367
R822 B.n216 B.n215 163.367
R823 B.n220 B.n219 163.367
R824 B.n224 B.n223 163.367
R825 B.n228 B.n227 163.367
R826 B.n232 B.n231 163.367
R827 B.n236 B.n235 163.367
R828 B.n240 B.n239 163.367
R829 B.n244 B.n243 163.367
R830 B.n249 B.n248 163.367
R831 B.n253 B.n252 163.367
R832 B.n257 B.n256 163.367
R833 B.n261 B.n260 163.367
R834 B.n265 B.n264 163.367
R835 B.n269 B.n268 163.367
R836 B.n273 B.n272 163.367
R837 B.n277 B.n276 163.367
R838 B.n281 B.n280 163.367
R839 B.n285 B.n284 163.367
R840 B.n289 B.n288 163.367
R841 B.n293 B.n292 163.367
R842 B.n297 B.n296 163.367
R843 B.n301 B.n300 163.367
R844 B.n305 B.n304 163.367
R845 B.n309 B.n308 163.367
R846 B.n313 B.n312 163.367
R847 B.n317 B.n316 163.367
R848 B.n321 B.n320 163.367
R849 B.n325 B.n324 163.367
R850 B.n329 B.n328 163.367
R851 B.n333 B.n332 163.367
R852 B.n337 B.n336 163.367
R853 B.n341 B.n340 163.367
R854 B.n345 B.n344 163.367
R855 B.n349 B.n348 163.367
R856 B.n353 B.n352 163.367
R857 B.n357 B.n356 163.367
R858 B.n361 B.n360 163.367
R859 B.n365 B.n364 163.367
R860 B.n369 B.n368 163.367
R861 B.n908 B.n130 163.367
R862 B.n749 B.n442 163.367
R863 B.n749 B.n436 163.367
R864 B.n757 B.n436 163.367
R865 B.n757 B.n434 163.367
R866 B.n761 B.n434 163.367
R867 B.n761 B.n429 163.367
R868 B.n770 B.n429 163.367
R869 B.n770 B.n427 163.367
R870 B.n774 B.n427 163.367
R871 B.n774 B.n421 163.367
R872 B.n782 B.n421 163.367
R873 B.n782 B.n419 163.367
R874 B.n786 B.n419 163.367
R875 B.n786 B.n413 163.367
R876 B.n794 B.n413 163.367
R877 B.n794 B.n411 163.367
R878 B.n798 B.n411 163.367
R879 B.n798 B.n405 163.367
R880 B.n806 B.n405 163.367
R881 B.n806 B.n403 163.367
R882 B.n810 B.n403 163.367
R883 B.n810 B.n397 163.367
R884 B.n818 B.n397 163.367
R885 B.n818 B.n395 163.367
R886 B.n822 B.n395 163.367
R887 B.n822 B.n389 163.367
R888 B.n830 B.n389 163.367
R889 B.n830 B.n387 163.367
R890 B.n834 B.n387 163.367
R891 B.n834 B.n380 163.367
R892 B.n842 B.n380 163.367
R893 B.n842 B.n378 163.367
R894 B.n847 B.n378 163.367
R895 B.n847 B.n373 163.367
R896 B.n855 B.n373 163.367
R897 B.n856 B.n855 163.367
R898 B.n856 B.n5 163.367
R899 B.n6 B.n5 163.367
R900 B.n7 B.n6 163.367
R901 B.n862 B.n7 163.367
R902 B.n863 B.n862 163.367
R903 B.n863 B.n13 163.367
R904 B.n14 B.n13 163.367
R905 B.n15 B.n14 163.367
R906 B.n868 B.n15 163.367
R907 B.n868 B.n20 163.367
R908 B.n21 B.n20 163.367
R909 B.n22 B.n21 163.367
R910 B.n873 B.n22 163.367
R911 B.n873 B.n27 163.367
R912 B.n28 B.n27 163.367
R913 B.n29 B.n28 163.367
R914 B.n878 B.n29 163.367
R915 B.n878 B.n34 163.367
R916 B.n35 B.n34 163.367
R917 B.n36 B.n35 163.367
R918 B.n883 B.n36 163.367
R919 B.n883 B.n41 163.367
R920 B.n42 B.n41 163.367
R921 B.n43 B.n42 163.367
R922 B.n888 B.n43 163.367
R923 B.n888 B.n48 163.367
R924 B.n49 B.n48 163.367
R925 B.n50 B.n49 163.367
R926 B.n893 B.n50 163.367
R927 B.n893 B.n55 163.367
R928 B.n56 B.n55 163.367
R929 B.n57 B.n56 163.367
R930 B.n898 B.n57 163.367
R931 B.n898 B.n62 163.367
R932 B.n63 B.n62 163.367
R933 B.n64 B.n63 163.367
R934 B.n903 B.n64 163.367
R935 B.n903 B.n69 163.367
R936 B.n70 B.n69 163.367
R937 B.n503 B.n502 163.367
R938 B.n736 B.n502 163.367
R939 B.n734 B.n733 163.367
R940 B.n730 B.n729 163.367
R941 B.n726 B.n725 163.367
R942 B.n722 B.n721 163.367
R943 B.n718 B.n717 163.367
R944 B.n714 B.n713 163.367
R945 B.n710 B.n709 163.367
R946 B.n706 B.n705 163.367
R947 B.n702 B.n701 163.367
R948 B.n698 B.n697 163.367
R949 B.n694 B.n693 163.367
R950 B.n690 B.n689 163.367
R951 B.n686 B.n685 163.367
R952 B.n682 B.n681 163.367
R953 B.n678 B.n677 163.367
R954 B.n674 B.n673 163.367
R955 B.n670 B.n669 163.367
R956 B.n666 B.n665 163.367
R957 B.n662 B.n661 163.367
R958 B.n658 B.n657 163.367
R959 B.n654 B.n653 163.367
R960 B.n650 B.n649 163.367
R961 B.n646 B.n645 163.367
R962 B.n642 B.n641 163.367
R963 B.n638 B.n637 163.367
R964 B.n634 B.n633 163.367
R965 B.n630 B.n629 163.367
R966 B.n626 B.n625 163.367
R967 B.n622 B.n621 163.367
R968 B.n618 B.n617 163.367
R969 B.n613 B.n612 163.367
R970 B.n609 B.n608 163.367
R971 B.n605 B.n604 163.367
R972 B.n601 B.n600 163.367
R973 B.n597 B.n596 163.367
R974 B.n593 B.n592 163.367
R975 B.n589 B.n588 163.367
R976 B.n585 B.n584 163.367
R977 B.n581 B.n580 163.367
R978 B.n577 B.n576 163.367
R979 B.n573 B.n572 163.367
R980 B.n569 B.n568 163.367
R981 B.n565 B.n564 163.367
R982 B.n561 B.n560 163.367
R983 B.n557 B.n556 163.367
R984 B.n553 B.n552 163.367
R985 B.n549 B.n548 163.367
R986 B.n545 B.n544 163.367
R987 B.n541 B.n540 163.367
R988 B.n537 B.n536 163.367
R989 B.n533 B.n532 163.367
R990 B.n529 B.n528 163.367
R991 B.n525 B.n524 163.367
R992 B.n521 B.n520 163.367
R993 B.n517 B.n516 163.367
R994 B.n513 B.n512 163.367
R995 B.n509 B.n444 163.367
R996 B.n751 B.n440 163.367
R997 B.n751 B.n438 163.367
R998 B.n755 B.n438 163.367
R999 B.n755 B.n432 163.367
R1000 B.n764 B.n432 163.367
R1001 B.n764 B.n430 163.367
R1002 B.n768 B.n430 163.367
R1003 B.n768 B.n425 163.367
R1004 B.n776 B.n425 163.367
R1005 B.n776 B.n423 163.367
R1006 B.n780 B.n423 163.367
R1007 B.n780 B.n417 163.367
R1008 B.n788 B.n417 163.367
R1009 B.n788 B.n415 163.367
R1010 B.n792 B.n415 163.367
R1011 B.n792 B.n409 163.367
R1012 B.n800 B.n409 163.367
R1013 B.n800 B.n407 163.367
R1014 B.n804 B.n407 163.367
R1015 B.n804 B.n401 163.367
R1016 B.n812 B.n401 163.367
R1017 B.n812 B.n399 163.367
R1018 B.n816 B.n399 163.367
R1019 B.n816 B.n393 163.367
R1020 B.n824 B.n393 163.367
R1021 B.n824 B.n391 163.367
R1022 B.n828 B.n391 163.367
R1023 B.n828 B.n385 163.367
R1024 B.n836 B.n385 163.367
R1025 B.n836 B.n383 163.367
R1026 B.n840 B.n383 163.367
R1027 B.n840 B.n377 163.367
R1028 B.n849 B.n377 163.367
R1029 B.n849 B.n375 163.367
R1030 B.n853 B.n375 163.367
R1031 B.n853 B.n3 163.367
R1032 B.n985 B.n3 163.367
R1033 B.n981 B.n2 163.367
R1034 B.n981 B.n980 163.367
R1035 B.n980 B.n9 163.367
R1036 B.n976 B.n9 163.367
R1037 B.n976 B.n11 163.367
R1038 B.n972 B.n11 163.367
R1039 B.n972 B.n17 163.367
R1040 B.n968 B.n17 163.367
R1041 B.n968 B.n19 163.367
R1042 B.n964 B.n19 163.367
R1043 B.n964 B.n24 163.367
R1044 B.n960 B.n24 163.367
R1045 B.n960 B.n26 163.367
R1046 B.n956 B.n26 163.367
R1047 B.n956 B.n31 163.367
R1048 B.n952 B.n31 163.367
R1049 B.n952 B.n33 163.367
R1050 B.n948 B.n33 163.367
R1051 B.n948 B.n38 163.367
R1052 B.n944 B.n38 163.367
R1053 B.n944 B.n40 163.367
R1054 B.n940 B.n40 163.367
R1055 B.n940 B.n45 163.367
R1056 B.n936 B.n45 163.367
R1057 B.n936 B.n47 163.367
R1058 B.n932 B.n47 163.367
R1059 B.n932 B.n52 163.367
R1060 B.n928 B.n52 163.367
R1061 B.n928 B.n54 163.367
R1062 B.n924 B.n54 163.367
R1063 B.n924 B.n58 163.367
R1064 B.n920 B.n58 163.367
R1065 B.n920 B.n60 163.367
R1066 B.n916 B.n60 163.367
R1067 B.n916 B.n66 163.367
R1068 B.n912 B.n66 163.367
R1069 B.n912 B.n68 163.367
R1070 B.n131 B.t9 108.853
R1071 B.n507 B.t20 108.853
R1072 B.n134 B.t12 108.832
R1073 B.n504 B.t17 108.832
R1074 B.n136 B.n71 71.676
R1075 B.n140 B.n72 71.676
R1076 B.n144 B.n73 71.676
R1077 B.n148 B.n74 71.676
R1078 B.n152 B.n75 71.676
R1079 B.n156 B.n76 71.676
R1080 B.n160 B.n77 71.676
R1081 B.n164 B.n78 71.676
R1082 B.n168 B.n79 71.676
R1083 B.n172 B.n80 71.676
R1084 B.n176 B.n81 71.676
R1085 B.n180 B.n82 71.676
R1086 B.n184 B.n83 71.676
R1087 B.n188 B.n84 71.676
R1088 B.n192 B.n85 71.676
R1089 B.n196 B.n86 71.676
R1090 B.n200 B.n87 71.676
R1091 B.n204 B.n88 71.676
R1092 B.n208 B.n89 71.676
R1093 B.n212 B.n90 71.676
R1094 B.n216 B.n91 71.676
R1095 B.n220 B.n92 71.676
R1096 B.n224 B.n93 71.676
R1097 B.n228 B.n94 71.676
R1098 B.n232 B.n95 71.676
R1099 B.n236 B.n96 71.676
R1100 B.n240 B.n97 71.676
R1101 B.n244 B.n98 71.676
R1102 B.n249 B.n99 71.676
R1103 B.n253 B.n100 71.676
R1104 B.n257 B.n101 71.676
R1105 B.n261 B.n102 71.676
R1106 B.n265 B.n103 71.676
R1107 B.n269 B.n104 71.676
R1108 B.n273 B.n105 71.676
R1109 B.n277 B.n106 71.676
R1110 B.n281 B.n107 71.676
R1111 B.n285 B.n108 71.676
R1112 B.n289 B.n109 71.676
R1113 B.n293 B.n110 71.676
R1114 B.n297 B.n111 71.676
R1115 B.n301 B.n112 71.676
R1116 B.n305 B.n113 71.676
R1117 B.n309 B.n114 71.676
R1118 B.n313 B.n115 71.676
R1119 B.n317 B.n116 71.676
R1120 B.n321 B.n117 71.676
R1121 B.n325 B.n118 71.676
R1122 B.n329 B.n119 71.676
R1123 B.n333 B.n120 71.676
R1124 B.n337 B.n121 71.676
R1125 B.n341 B.n122 71.676
R1126 B.n345 B.n123 71.676
R1127 B.n349 B.n124 71.676
R1128 B.n353 B.n125 71.676
R1129 B.n357 B.n126 71.676
R1130 B.n361 B.n127 71.676
R1131 B.n365 B.n128 71.676
R1132 B.n369 B.n129 71.676
R1133 B.n130 B.n129 71.676
R1134 B.n368 B.n128 71.676
R1135 B.n364 B.n127 71.676
R1136 B.n360 B.n126 71.676
R1137 B.n356 B.n125 71.676
R1138 B.n352 B.n124 71.676
R1139 B.n348 B.n123 71.676
R1140 B.n344 B.n122 71.676
R1141 B.n340 B.n121 71.676
R1142 B.n336 B.n120 71.676
R1143 B.n332 B.n119 71.676
R1144 B.n328 B.n118 71.676
R1145 B.n324 B.n117 71.676
R1146 B.n320 B.n116 71.676
R1147 B.n316 B.n115 71.676
R1148 B.n312 B.n114 71.676
R1149 B.n308 B.n113 71.676
R1150 B.n304 B.n112 71.676
R1151 B.n300 B.n111 71.676
R1152 B.n296 B.n110 71.676
R1153 B.n292 B.n109 71.676
R1154 B.n288 B.n108 71.676
R1155 B.n284 B.n107 71.676
R1156 B.n280 B.n106 71.676
R1157 B.n276 B.n105 71.676
R1158 B.n272 B.n104 71.676
R1159 B.n268 B.n103 71.676
R1160 B.n264 B.n102 71.676
R1161 B.n260 B.n101 71.676
R1162 B.n256 B.n100 71.676
R1163 B.n252 B.n99 71.676
R1164 B.n248 B.n98 71.676
R1165 B.n243 B.n97 71.676
R1166 B.n239 B.n96 71.676
R1167 B.n235 B.n95 71.676
R1168 B.n231 B.n94 71.676
R1169 B.n227 B.n93 71.676
R1170 B.n223 B.n92 71.676
R1171 B.n219 B.n91 71.676
R1172 B.n215 B.n90 71.676
R1173 B.n211 B.n89 71.676
R1174 B.n207 B.n88 71.676
R1175 B.n203 B.n87 71.676
R1176 B.n199 B.n86 71.676
R1177 B.n195 B.n85 71.676
R1178 B.n191 B.n84 71.676
R1179 B.n187 B.n83 71.676
R1180 B.n183 B.n82 71.676
R1181 B.n179 B.n81 71.676
R1182 B.n175 B.n80 71.676
R1183 B.n171 B.n79 71.676
R1184 B.n167 B.n78 71.676
R1185 B.n163 B.n77 71.676
R1186 B.n159 B.n76 71.676
R1187 B.n155 B.n75 71.676
R1188 B.n151 B.n74 71.676
R1189 B.n147 B.n73 71.676
R1190 B.n143 B.n72 71.676
R1191 B.n139 B.n71 71.676
R1192 B.n742 B.n741 71.676
R1193 B.n736 B.n445 71.676
R1194 B.n733 B.n446 71.676
R1195 B.n729 B.n447 71.676
R1196 B.n725 B.n448 71.676
R1197 B.n721 B.n449 71.676
R1198 B.n717 B.n450 71.676
R1199 B.n713 B.n451 71.676
R1200 B.n709 B.n452 71.676
R1201 B.n705 B.n453 71.676
R1202 B.n701 B.n454 71.676
R1203 B.n697 B.n455 71.676
R1204 B.n693 B.n456 71.676
R1205 B.n689 B.n457 71.676
R1206 B.n685 B.n458 71.676
R1207 B.n681 B.n459 71.676
R1208 B.n677 B.n460 71.676
R1209 B.n673 B.n461 71.676
R1210 B.n669 B.n462 71.676
R1211 B.n665 B.n463 71.676
R1212 B.n661 B.n464 71.676
R1213 B.n657 B.n465 71.676
R1214 B.n653 B.n466 71.676
R1215 B.n649 B.n467 71.676
R1216 B.n645 B.n468 71.676
R1217 B.n641 B.n469 71.676
R1218 B.n637 B.n470 71.676
R1219 B.n633 B.n471 71.676
R1220 B.n629 B.n472 71.676
R1221 B.n625 B.n473 71.676
R1222 B.n621 B.n474 71.676
R1223 B.n617 B.n475 71.676
R1224 B.n612 B.n476 71.676
R1225 B.n608 B.n477 71.676
R1226 B.n604 B.n478 71.676
R1227 B.n600 B.n479 71.676
R1228 B.n596 B.n480 71.676
R1229 B.n592 B.n481 71.676
R1230 B.n588 B.n482 71.676
R1231 B.n584 B.n483 71.676
R1232 B.n580 B.n484 71.676
R1233 B.n576 B.n485 71.676
R1234 B.n572 B.n486 71.676
R1235 B.n568 B.n487 71.676
R1236 B.n564 B.n488 71.676
R1237 B.n560 B.n489 71.676
R1238 B.n556 B.n490 71.676
R1239 B.n552 B.n491 71.676
R1240 B.n548 B.n492 71.676
R1241 B.n544 B.n493 71.676
R1242 B.n540 B.n494 71.676
R1243 B.n536 B.n495 71.676
R1244 B.n532 B.n496 71.676
R1245 B.n528 B.n497 71.676
R1246 B.n524 B.n498 71.676
R1247 B.n520 B.n499 71.676
R1248 B.n516 B.n500 71.676
R1249 B.n512 B.n501 71.676
R1250 B.n744 B.n444 71.676
R1251 B.n742 B.n503 71.676
R1252 B.n734 B.n445 71.676
R1253 B.n730 B.n446 71.676
R1254 B.n726 B.n447 71.676
R1255 B.n722 B.n448 71.676
R1256 B.n718 B.n449 71.676
R1257 B.n714 B.n450 71.676
R1258 B.n710 B.n451 71.676
R1259 B.n706 B.n452 71.676
R1260 B.n702 B.n453 71.676
R1261 B.n698 B.n454 71.676
R1262 B.n694 B.n455 71.676
R1263 B.n690 B.n456 71.676
R1264 B.n686 B.n457 71.676
R1265 B.n682 B.n458 71.676
R1266 B.n678 B.n459 71.676
R1267 B.n674 B.n460 71.676
R1268 B.n670 B.n461 71.676
R1269 B.n666 B.n462 71.676
R1270 B.n662 B.n463 71.676
R1271 B.n658 B.n464 71.676
R1272 B.n654 B.n465 71.676
R1273 B.n650 B.n466 71.676
R1274 B.n646 B.n467 71.676
R1275 B.n642 B.n468 71.676
R1276 B.n638 B.n469 71.676
R1277 B.n634 B.n470 71.676
R1278 B.n630 B.n471 71.676
R1279 B.n626 B.n472 71.676
R1280 B.n622 B.n473 71.676
R1281 B.n618 B.n474 71.676
R1282 B.n613 B.n475 71.676
R1283 B.n609 B.n476 71.676
R1284 B.n605 B.n477 71.676
R1285 B.n601 B.n478 71.676
R1286 B.n597 B.n479 71.676
R1287 B.n593 B.n480 71.676
R1288 B.n589 B.n481 71.676
R1289 B.n585 B.n482 71.676
R1290 B.n581 B.n483 71.676
R1291 B.n577 B.n484 71.676
R1292 B.n573 B.n485 71.676
R1293 B.n569 B.n486 71.676
R1294 B.n565 B.n487 71.676
R1295 B.n561 B.n488 71.676
R1296 B.n557 B.n489 71.676
R1297 B.n553 B.n490 71.676
R1298 B.n549 B.n491 71.676
R1299 B.n545 B.n492 71.676
R1300 B.n541 B.n493 71.676
R1301 B.n537 B.n494 71.676
R1302 B.n533 B.n495 71.676
R1303 B.n529 B.n496 71.676
R1304 B.n525 B.n497 71.676
R1305 B.n521 B.n498 71.676
R1306 B.n517 B.n499 71.676
R1307 B.n513 B.n500 71.676
R1308 B.n509 B.n501 71.676
R1309 B.n745 B.n744 71.676
R1310 B.n986 B.n985 71.676
R1311 B.n986 B.n2 71.676
R1312 B.n132 B.t10 69.8713
R1313 B.n508 B.t19 69.8713
R1314 B.n135 B.t13 69.8495
R1315 B.n505 B.t16 69.8495
R1316 B.n743 B.n441 68.3549
R1317 B.n910 B.n909 68.3549
R1318 B.n246 B.n135 59.5399
R1319 B.n133 B.n132 59.5399
R1320 B.n615 B.n508 59.5399
R1321 B.n506 B.n505 59.5399
R1322 B.n135 B.n134 38.9823
R1323 B.n132 B.n131 38.9823
R1324 B.n508 B.n507 38.9823
R1325 B.n505 B.n504 38.9823
R1326 B.n750 B.n441 34.4309
R1327 B.n750 B.n437 34.4309
R1328 B.n756 B.n437 34.4309
R1329 B.n756 B.n433 34.4309
R1330 B.n763 B.n433 34.4309
R1331 B.n763 B.n762 34.4309
R1332 B.n769 B.n426 34.4309
R1333 B.n775 B.n426 34.4309
R1334 B.n775 B.n422 34.4309
R1335 B.n781 B.n422 34.4309
R1336 B.n781 B.n418 34.4309
R1337 B.n787 B.n418 34.4309
R1338 B.n787 B.n414 34.4309
R1339 B.n793 B.n414 34.4309
R1340 B.n799 B.n410 34.4309
R1341 B.n799 B.n406 34.4309
R1342 B.n805 B.n406 34.4309
R1343 B.n805 B.n402 34.4309
R1344 B.n811 B.n402 34.4309
R1345 B.n817 B.n398 34.4309
R1346 B.n817 B.n394 34.4309
R1347 B.n823 B.n394 34.4309
R1348 B.n823 B.n390 34.4309
R1349 B.n829 B.n390 34.4309
R1350 B.n835 B.n386 34.4309
R1351 B.n835 B.n381 34.4309
R1352 B.n841 B.n381 34.4309
R1353 B.n841 B.n382 34.4309
R1354 B.n848 B.n374 34.4309
R1355 B.n854 B.n374 34.4309
R1356 B.n854 B.n4 34.4309
R1357 B.n984 B.n4 34.4309
R1358 B.n984 B.n983 34.4309
R1359 B.n983 B.n982 34.4309
R1360 B.n982 B.n8 34.4309
R1361 B.n12 B.n8 34.4309
R1362 B.n975 B.n12 34.4309
R1363 B.n974 B.n973 34.4309
R1364 B.n973 B.n16 34.4309
R1365 B.n967 B.n16 34.4309
R1366 B.n967 B.n966 34.4309
R1367 B.n965 B.n23 34.4309
R1368 B.n959 B.n23 34.4309
R1369 B.n959 B.n958 34.4309
R1370 B.n958 B.n957 34.4309
R1371 B.n957 B.n30 34.4309
R1372 B.n951 B.n950 34.4309
R1373 B.n950 B.n949 34.4309
R1374 B.n949 B.n37 34.4309
R1375 B.n943 B.n37 34.4309
R1376 B.n943 B.n942 34.4309
R1377 B.n941 B.n44 34.4309
R1378 B.n935 B.n44 34.4309
R1379 B.n935 B.n934 34.4309
R1380 B.n934 B.n933 34.4309
R1381 B.n933 B.n51 34.4309
R1382 B.n927 B.n51 34.4309
R1383 B.n927 B.n926 34.4309
R1384 B.n926 B.n925 34.4309
R1385 B.n919 B.n61 34.4309
R1386 B.n919 B.n918 34.4309
R1387 B.n918 B.n917 34.4309
R1388 B.n917 B.n65 34.4309
R1389 B.n911 B.n65 34.4309
R1390 B.n911 B.n910 34.4309
R1391 B.n740 B.n439 34.1859
R1392 B.n747 B.n746 34.1859
R1393 B.n907 B.n906 34.1859
R1394 B.n137 B.n67 34.1859
R1395 B.t4 B.n386 33.4182
R1396 B.n966 B.t2 33.4182
R1397 B.n382 B.t0 32.4056
R1398 B.t21 B.n974 32.4056
R1399 B.n769 B.t15 31.3929
R1400 B.n925 B.t8 31.3929
R1401 B.t5 B.n398 30.3802
R1402 B.t1 B.n30 30.3802
R1403 B.t6 B.n410 27.3423
R1404 B.n942 B.t3 27.3423
R1405 B B.n987 18.0485
R1406 B.n752 B.n439 10.6151
R1407 B.n753 B.n752 10.6151
R1408 B.n754 B.n753 10.6151
R1409 B.n754 B.n431 10.6151
R1410 B.n765 B.n431 10.6151
R1411 B.n766 B.n765 10.6151
R1412 B.n767 B.n766 10.6151
R1413 B.n767 B.n424 10.6151
R1414 B.n777 B.n424 10.6151
R1415 B.n778 B.n777 10.6151
R1416 B.n779 B.n778 10.6151
R1417 B.n779 B.n416 10.6151
R1418 B.n789 B.n416 10.6151
R1419 B.n790 B.n789 10.6151
R1420 B.n791 B.n790 10.6151
R1421 B.n791 B.n408 10.6151
R1422 B.n801 B.n408 10.6151
R1423 B.n802 B.n801 10.6151
R1424 B.n803 B.n802 10.6151
R1425 B.n803 B.n400 10.6151
R1426 B.n813 B.n400 10.6151
R1427 B.n814 B.n813 10.6151
R1428 B.n815 B.n814 10.6151
R1429 B.n815 B.n392 10.6151
R1430 B.n825 B.n392 10.6151
R1431 B.n826 B.n825 10.6151
R1432 B.n827 B.n826 10.6151
R1433 B.n827 B.n384 10.6151
R1434 B.n837 B.n384 10.6151
R1435 B.n838 B.n837 10.6151
R1436 B.n839 B.n838 10.6151
R1437 B.n839 B.n376 10.6151
R1438 B.n850 B.n376 10.6151
R1439 B.n851 B.n850 10.6151
R1440 B.n852 B.n851 10.6151
R1441 B.n852 B.n0 10.6151
R1442 B.n740 B.n739 10.6151
R1443 B.n739 B.n738 10.6151
R1444 B.n738 B.n737 10.6151
R1445 B.n737 B.n735 10.6151
R1446 B.n735 B.n732 10.6151
R1447 B.n732 B.n731 10.6151
R1448 B.n731 B.n728 10.6151
R1449 B.n728 B.n727 10.6151
R1450 B.n727 B.n724 10.6151
R1451 B.n724 B.n723 10.6151
R1452 B.n723 B.n720 10.6151
R1453 B.n720 B.n719 10.6151
R1454 B.n719 B.n716 10.6151
R1455 B.n716 B.n715 10.6151
R1456 B.n715 B.n712 10.6151
R1457 B.n712 B.n711 10.6151
R1458 B.n711 B.n708 10.6151
R1459 B.n708 B.n707 10.6151
R1460 B.n707 B.n704 10.6151
R1461 B.n704 B.n703 10.6151
R1462 B.n703 B.n700 10.6151
R1463 B.n700 B.n699 10.6151
R1464 B.n699 B.n696 10.6151
R1465 B.n696 B.n695 10.6151
R1466 B.n695 B.n692 10.6151
R1467 B.n692 B.n691 10.6151
R1468 B.n691 B.n688 10.6151
R1469 B.n688 B.n687 10.6151
R1470 B.n687 B.n684 10.6151
R1471 B.n684 B.n683 10.6151
R1472 B.n683 B.n680 10.6151
R1473 B.n680 B.n679 10.6151
R1474 B.n679 B.n676 10.6151
R1475 B.n676 B.n675 10.6151
R1476 B.n675 B.n672 10.6151
R1477 B.n672 B.n671 10.6151
R1478 B.n671 B.n668 10.6151
R1479 B.n668 B.n667 10.6151
R1480 B.n667 B.n664 10.6151
R1481 B.n664 B.n663 10.6151
R1482 B.n663 B.n660 10.6151
R1483 B.n660 B.n659 10.6151
R1484 B.n659 B.n656 10.6151
R1485 B.n656 B.n655 10.6151
R1486 B.n655 B.n652 10.6151
R1487 B.n652 B.n651 10.6151
R1488 B.n651 B.n648 10.6151
R1489 B.n648 B.n647 10.6151
R1490 B.n647 B.n644 10.6151
R1491 B.n644 B.n643 10.6151
R1492 B.n643 B.n640 10.6151
R1493 B.n640 B.n639 10.6151
R1494 B.n639 B.n636 10.6151
R1495 B.n636 B.n635 10.6151
R1496 B.n632 B.n631 10.6151
R1497 B.n631 B.n628 10.6151
R1498 B.n628 B.n627 10.6151
R1499 B.n627 B.n624 10.6151
R1500 B.n624 B.n623 10.6151
R1501 B.n623 B.n620 10.6151
R1502 B.n620 B.n619 10.6151
R1503 B.n619 B.n616 10.6151
R1504 B.n614 B.n611 10.6151
R1505 B.n611 B.n610 10.6151
R1506 B.n610 B.n607 10.6151
R1507 B.n607 B.n606 10.6151
R1508 B.n606 B.n603 10.6151
R1509 B.n603 B.n602 10.6151
R1510 B.n602 B.n599 10.6151
R1511 B.n599 B.n598 10.6151
R1512 B.n598 B.n595 10.6151
R1513 B.n595 B.n594 10.6151
R1514 B.n594 B.n591 10.6151
R1515 B.n591 B.n590 10.6151
R1516 B.n590 B.n587 10.6151
R1517 B.n587 B.n586 10.6151
R1518 B.n586 B.n583 10.6151
R1519 B.n583 B.n582 10.6151
R1520 B.n582 B.n579 10.6151
R1521 B.n579 B.n578 10.6151
R1522 B.n578 B.n575 10.6151
R1523 B.n575 B.n574 10.6151
R1524 B.n574 B.n571 10.6151
R1525 B.n571 B.n570 10.6151
R1526 B.n570 B.n567 10.6151
R1527 B.n567 B.n566 10.6151
R1528 B.n566 B.n563 10.6151
R1529 B.n563 B.n562 10.6151
R1530 B.n562 B.n559 10.6151
R1531 B.n559 B.n558 10.6151
R1532 B.n558 B.n555 10.6151
R1533 B.n555 B.n554 10.6151
R1534 B.n554 B.n551 10.6151
R1535 B.n551 B.n550 10.6151
R1536 B.n550 B.n547 10.6151
R1537 B.n547 B.n546 10.6151
R1538 B.n546 B.n543 10.6151
R1539 B.n543 B.n542 10.6151
R1540 B.n542 B.n539 10.6151
R1541 B.n539 B.n538 10.6151
R1542 B.n538 B.n535 10.6151
R1543 B.n535 B.n534 10.6151
R1544 B.n534 B.n531 10.6151
R1545 B.n531 B.n530 10.6151
R1546 B.n530 B.n527 10.6151
R1547 B.n527 B.n526 10.6151
R1548 B.n526 B.n523 10.6151
R1549 B.n523 B.n522 10.6151
R1550 B.n522 B.n519 10.6151
R1551 B.n519 B.n518 10.6151
R1552 B.n518 B.n515 10.6151
R1553 B.n515 B.n514 10.6151
R1554 B.n514 B.n511 10.6151
R1555 B.n511 B.n510 10.6151
R1556 B.n510 B.n443 10.6151
R1557 B.n746 B.n443 10.6151
R1558 B.n748 B.n747 10.6151
R1559 B.n748 B.n435 10.6151
R1560 B.n758 B.n435 10.6151
R1561 B.n759 B.n758 10.6151
R1562 B.n760 B.n759 10.6151
R1563 B.n760 B.n428 10.6151
R1564 B.n771 B.n428 10.6151
R1565 B.n772 B.n771 10.6151
R1566 B.n773 B.n772 10.6151
R1567 B.n773 B.n420 10.6151
R1568 B.n783 B.n420 10.6151
R1569 B.n784 B.n783 10.6151
R1570 B.n785 B.n784 10.6151
R1571 B.n785 B.n412 10.6151
R1572 B.n795 B.n412 10.6151
R1573 B.n796 B.n795 10.6151
R1574 B.n797 B.n796 10.6151
R1575 B.n797 B.n404 10.6151
R1576 B.n807 B.n404 10.6151
R1577 B.n808 B.n807 10.6151
R1578 B.n809 B.n808 10.6151
R1579 B.n809 B.n396 10.6151
R1580 B.n819 B.n396 10.6151
R1581 B.n820 B.n819 10.6151
R1582 B.n821 B.n820 10.6151
R1583 B.n821 B.n388 10.6151
R1584 B.n831 B.n388 10.6151
R1585 B.n832 B.n831 10.6151
R1586 B.n833 B.n832 10.6151
R1587 B.n833 B.n379 10.6151
R1588 B.n843 B.n379 10.6151
R1589 B.n844 B.n843 10.6151
R1590 B.n846 B.n844 10.6151
R1591 B.n846 B.n845 10.6151
R1592 B.n845 B.n372 10.6151
R1593 B.n857 B.n372 10.6151
R1594 B.n858 B.n857 10.6151
R1595 B.n859 B.n858 10.6151
R1596 B.n860 B.n859 10.6151
R1597 B.n861 B.n860 10.6151
R1598 B.n864 B.n861 10.6151
R1599 B.n865 B.n864 10.6151
R1600 B.n866 B.n865 10.6151
R1601 B.n867 B.n866 10.6151
R1602 B.n869 B.n867 10.6151
R1603 B.n870 B.n869 10.6151
R1604 B.n871 B.n870 10.6151
R1605 B.n872 B.n871 10.6151
R1606 B.n874 B.n872 10.6151
R1607 B.n875 B.n874 10.6151
R1608 B.n876 B.n875 10.6151
R1609 B.n877 B.n876 10.6151
R1610 B.n879 B.n877 10.6151
R1611 B.n880 B.n879 10.6151
R1612 B.n881 B.n880 10.6151
R1613 B.n882 B.n881 10.6151
R1614 B.n884 B.n882 10.6151
R1615 B.n885 B.n884 10.6151
R1616 B.n886 B.n885 10.6151
R1617 B.n887 B.n886 10.6151
R1618 B.n889 B.n887 10.6151
R1619 B.n890 B.n889 10.6151
R1620 B.n891 B.n890 10.6151
R1621 B.n892 B.n891 10.6151
R1622 B.n894 B.n892 10.6151
R1623 B.n895 B.n894 10.6151
R1624 B.n896 B.n895 10.6151
R1625 B.n897 B.n896 10.6151
R1626 B.n899 B.n897 10.6151
R1627 B.n900 B.n899 10.6151
R1628 B.n901 B.n900 10.6151
R1629 B.n902 B.n901 10.6151
R1630 B.n904 B.n902 10.6151
R1631 B.n905 B.n904 10.6151
R1632 B.n906 B.n905 10.6151
R1633 B.n979 B.n1 10.6151
R1634 B.n979 B.n978 10.6151
R1635 B.n978 B.n977 10.6151
R1636 B.n977 B.n10 10.6151
R1637 B.n971 B.n10 10.6151
R1638 B.n971 B.n970 10.6151
R1639 B.n970 B.n969 10.6151
R1640 B.n969 B.n18 10.6151
R1641 B.n963 B.n18 10.6151
R1642 B.n963 B.n962 10.6151
R1643 B.n962 B.n961 10.6151
R1644 B.n961 B.n25 10.6151
R1645 B.n955 B.n25 10.6151
R1646 B.n955 B.n954 10.6151
R1647 B.n954 B.n953 10.6151
R1648 B.n953 B.n32 10.6151
R1649 B.n947 B.n32 10.6151
R1650 B.n947 B.n946 10.6151
R1651 B.n946 B.n945 10.6151
R1652 B.n945 B.n39 10.6151
R1653 B.n939 B.n39 10.6151
R1654 B.n939 B.n938 10.6151
R1655 B.n938 B.n937 10.6151
R1656 B.n937 B.n46 10.6151
R1657 B.n931 B.n46 10.6151
R1658 B.n931 B.n930 10.6151
R1659 B.n930 B.n929 10.6151
R1660 B.n929 B.n53 10.6151
R1661 B.n923 B.n53 10.6151
R1662 B.n923 B.n922 10.6151
R1663 B.n922 B.n921 10.6151
R1664 B.n921 B.n59 10.6151
R1665 B.n915 B.n59 10.6151
R1666 B.n915 B.n914 10.6151
R1667 B.n914 B.n913 10.6151
R1668 B.n913 B.n67 10.6151
R1669 B.n138 B.n137 10.6151
R1670 B.n141 B.n138 10.6151
R1671 B.n142 B.n141 10.6151
R1672 B.n145 B.n142 10.6151
R1673 B.n146 B.n145 10.6151
R1674 B.n149 B.n146 10.6151
R1675 B.n150 B.n149 10.6151
R1676 B.n153 B.n150 10.6151
R1677 B.n154 B.n153 10.6151
R1678 B.n157 B.n154 10.6151
R1679 B.n158 B.n157 10.6151
R1680 B.n161 B.n158 10.6151
R1681 B.n162 B.n161 10.6151
R1682 B.n165 B.n162 10.6151
R1683 B.n166 B.n165 10.6151
R1684 B.n169 B.n166 10.6151
R1685 B.n170 B.n169 10.6151
R1686 B.n173 B.n170 10.6151
R1687 B.n174 B.n173 10.6151
R1688 B.n177 B.n174 10.6151
R1689 B.n178 B.n177 10.6151
R1690 B.n181 B.n178 10.6151
R1691 B.n182 B.n181 10.6151
R1692 B.n185 B.n182 10.6151
R1693 B.n186 B.n185 10.6151
R1694 B.n189 B.n186 10.6151
R1695 B.n190 B.n189 10.6151
R1696 B.n193 B.n190 10.6151
R1697 B.n194 B.n193 10.6151
R1698 B.n197 B.n194 10.6151
R1699 B.n198 B.n197 10.6151
R1700 B.n201 B.n198 10.6151
R1701 B.n202 B.n201 10.6151
R1702 B.n205 B.n202 10.6151
R1703 B.n206 B.n205 10.6151
R1704 B.n209 B.n206 10.6151
R1705 B.n210 B.n209 10.6151
R1706 B.n213 B.n210 10.6151
R1707 B.n214 B.n213 10.6151
R1708 B.n217 B.n214 10.6151
R1709 B.n218 B.n217 10.6151
R1710 B.n221 B.n218 10.6151
R1711 B.n222 B.n221 10.6151
R1712 B.n225 B.n222 10.6151
R1713 B.n226 B.n225 10.6151
R1714 B.n229 B.n226 10.6151
R1715 B.n230 B.n229 10.6151
R1716 B.n233 B.n230 10.6151
R1717 B.n234 B.n233 10.6151
R1718 B.n237 B.n234 10.6151
R1719 B.n238 B.n237 10.6151
R1720 B.n241 B.n238 10.6151
R1721 B.n242 B.n241 10.6151
R1722 B.n245 B.n242 10.6151
R1723 B.n250 B.n247 10.6151
R1724 B.n251 B.n250 10.6151
R1725 B.n254 B.n251 10.6151
R1726 B.n255 B.n254 10.6151
R1727 B.n258 B.n255 10.6151
R1728 B.n259 B.n258 10.6151
R1729 B.n262 B.n259 10.6151
R1730 B.n263 B.n262 10.6151
R1731 B.n267 B.n266 10.6151
R1732 B.n270 B.n267 10.6151
R1733 B.n271 B.n270 10.6151
R1734 B.n274 B.n271 10.6151
R1735 B.n275 B.n274 10.6151
R1736 B.n278 B.n275 10.6151
R1737 B.n279 B.n278 10.6151
R1738 B.n282 B.n279 10.6151
R1739 B.n283 B.n282 10.6151
R1740 B.n286 B.n283 10.6151
R1741 B.n287 B.n286 10.6151
R1742 B.n290 B.n287 10.6151
R1743 B.n291 B.n290 10.6151
R1744 B.n294 B.n291 10.6151
R1745 B.n295 B.n294 10.6151
R1746 B.n298 B.n295 10.6151
R1747 B.n299 B.n298 10.6151
R1748 B.n302 B.n299 10.6151
R1749 B.n303 B.n302 10.6151
R1750 B.n306 B.n303 10.6151
R1751 B.n307 B.n306 10.6151
R1752 B.n310 B.n307 10.6151
R1753 B.n311 B.n310 10.6151
R1754 B.n314 B.n311 10.6151
R1755 B.n315 B.n314 10.6151
R1756 B.n318 B.n315 10.6151
R1757 B.n319 B.n318 10.6151
R1758 B.n322 B.n319 10.6151
R1759 B.n323 B.n322 10.6151
R1760 B.n326 B.n323 10.6151
R1761 B.n327 B.n326 10.6151
R1762 B.n330 B.n327 10.6151
R1763 B.n331 B.n330 10.6151
R1764 B.n334 B.n331 10.6151
R1765 B.n335 B.n334 10.6151
R1766 B.n338 B.n335 10.6151
R1767 B.n339 B.n338 10.6151
R1768 B.n342 B.n339 10.6151
R1769 B.n343 B.n342 10.6151
R1770 B.n346 B.n343 10.6151
R1771 B.n347 B.n346 10.6151
R1772 B.n350 B.n347 10.6151
R1773 B.n351 B.n350 10.6151
R1774 B.n354 B.n351 10.6151
R1775 B.n355 B.n354 10.6151
R1776 B.n358 B.n355 10.6151
R1777 B.n359 B.n358 10.6151
R1778 B.n362 B.n359 10.6151
R1779 B.n363 B.n362 10.6151
R1780 B.n366 B.n363 10.6151
R1781 B.n367 B.n366 10.6151
R1782 B.n370 B.n367 10.6151
R1783 B.n371 B.n370 10.6151
R1784 B.n907 B.n371 10.6151
R1785 B.n987 B.n0 8.11757
R1786 B.n987 B.n1 8.11757
R1787 B.n793 B.t6 7.08911
R1788 B.t3 B.n941 7.08911
R1789 B.n632 B.n506 6.5566
R1790 B.n616 B.n615 6.5566
R1791 B.n247 B.n246 6.5566
R1792 B.n263 B.n133 6.5566
R1793 B.n635 B.n506 4.05904
R1794 B.n615 B.n614 4.05904
R1795 B.n246 B.n245 4.05904
R1796 B.n266 B.n133 4.05904
R1797 B.n811 B.t5 4.05113
R1798 B.n951 B.t1 4.05113
R1799 B.n762 B.t15 3.03847
R1800 B.n61 B.t8 3.03847
R1801 B.n848 B.t0 2.02582
R1802 B.n975 B.t21 2.02582
R1803 B.n829 B.t4 1.01316
R1804 B.t2 B.n965 1.01316
R1805 VN.n5 VN.t6 263.481
R1806 VN.n28 VN.t1 263.481
R1807 VN.n6 VN.t7 235.98
R1808 VN.n14 VN.t2 235.98
R1809 VN.n21 VN.t3 235.98
R1810 VN.n29 VN.t4 235.98
R1811 VN.n37 VN.t5 235.98
R1812 VN.n44 VN.t0 235.98
R1813 VN.n22 VN.n21 185.034
R1814 VN.n45 VN.n44 185.034
R1815 VN.n43 VN.n23 161.3
R1816 VN.n42 VN.n41 161.3
R1817 VN.n40 VN.n24 161.3
R1818 VN.n39 VN.n38 161.3
R1819 VN.n36 VN.n25 161.3
R1820 VN.n35 VN.n34 161.3
R1821 VN.n33 VN.n26 161.3
R1822 VN.n32 VN.n31 161.3
R1823 VN.n30 VN.n27 161.3
R1824 VN.n20 VN.n0 161.3
R1825 VN.n19 VN.n18 161.3
R1826 VN.n17 VN.n1 161.3
R1827 VN.n16 VN.n15 161.3
R1828 VN.n13 VN.n2 161.3
R1829 VN.n12 VN.n11 161.3
R1830 VN.n10 VN.n3 161.3
R1831 VN.n9 VN.n8 161.3
R1832 VN.n7 VN.n4 161.3
R1833 VN.n6 VN.n5 68.7155
R1834 VN.n29 VN.n28 68.7155
R1835 VN VN.n45 50.1691
R1836 VN.n19 VN.n1 41.4647
R1837 VN.n42 VN.n24 41.4647
R1838 VN.n8 VN.n3 40.4934
R1839 VN.n12 VN.n3 40.4934
R1840 VN.n31 VN.n26 40.4934
R1841 VN.n35 VN.n26 40.4934
R1842 VN.n15 VN.n1 39.5221
R1843 VN.n38 VN.n24 39.5221
R1844 VN.n8 VN.n7 24.4675
R1845 VN.n13 VN.n12 24.4675
R1846 VN.n20 VN.n19 24.4675
R1847 VN.n31 VN.n30 24.4675
R1848 VN.n36 VN.n35 24.4675
R1849 VN.n43 VN.n42 24.4675
R1850 VN.n15 VN.n14 24.2228
R1851 VN.n38 VN.n37 24.2228
R1852 VN.n28 VN.n27 18.9997
R1853 VN.n5 VN.n4 18.9997
R1854 VN.n21 VN.n20 0.73451
R1855 VN.n44 VN.n43 0.73451
R1856 VN.n7 VN.n6 0.24517
R1857 VN.n14 VN.n13 0.24517
R1858 VN.n30 VN.n29 0.24517
R1859 VN.n37 VN.n36 0.24517
R1860 VN.n45 VN.n23 0.189894
R1861 VN.n41 VN.n23 0.189894
R1862 VN.n41 VN.n40 0.189894
R1863 VN.n40 VN.n39 0.189894
R1864 VN.n39 VN.n25 0.189894
R1865 VN.n34 VN.n25 0.189894
R1866 VN.n34 VN.n33 0.189894
R1867 VN.n33 VN.n32 0.189894
R1868 VN.n32 VN.n27 0.189894
R1869 VN.n9 VN.n4 0.189894
R1870 VN.n10 VN.n9 0.189894
R1871 VN.n11 VN.n10 0.189894
R1872 VN.n11 VN.n2 0.189894
R1873 VN.n16 VN.n2 0.189894
R1874 VN.n17 VN.n16 0.189894
R1875 VN.n18 VN.n17 0.189894
R1876 VN.n18 VN.n0 0.189894
R1877 VN.n22 VN.n0 0.189894
R1878 VN VN.n22 0.0516364
R1879 VDD2.n2 VDD2.n1 61.7544
R1880 VDD2.n2 VDD2.n0 61.7544
R1881 VDD2 VDD2.n5 61.7516
R1882 VDD2.n4 VDD2.n3 60.9436
R1883 VDD2.n4 VDD2.n2 45.6937
R1884 VDD2.n5 VDD2.t3 1.20415
R1885 VDD2.n5 VDD2.t6 1.20415
R1886 VDD2.n3 VDD2.t7 1.20415
R1887 VDD2.n3 VDD2.t2 1.20415
R1888 VDD2.n1 VDD2.t5 1.20415
R1889 VDD2.n1 VDD2.t4 1.20415
R1890 VDD2.n0 VDD2.t1 1.20415
R1891 VDD2.n0 VDD2.t0 1.20415
R1892 VDD2 VDD2.n4 0.925069
C0 VP VTAIL 10.5071f
C1 VDD1 VDD2 1.29537f
C2 VN VDD1 0.149573f
C3 VP VDD1 10.8547f
C4 VTAIL VDD1 10.2078f
C5 VN VDD2 10.5839f
C6 VP VDD2 0.421282f
C7 VTAIL VDD2 10.2561f
C8 VN VP 7.36462f
C9 VN VTAIL 10.493f
C10 VDD2 B 4.805187f
C11 VDD1 B 5.141833f
C12 VTAIL B 12.390697f
C13 VN B 12.47026f
C14 VP B 10.780178f
C15 VDD2.t1 B 0.324f
C16 VDD2.t0 B 0.324f
C17 VDD2.n0 B 2.94632f
C18 VDD2.t5 B 0.324f
C19 VDD2.t4 B 0.324f
C20 VDD2.n1 B 2.94632f
C21 VDD2.n2 B 3.01334f
C22 VDD2.t7 B 0.324f
C23 VDD2.t2 B 0.324f
C24 VDD2.n3 B 2.9408f
C25 VDD2.n4 B 2.96163f
C26 VDD2.t3 B 0.324f
C27 VDD2.t6 B 0.324f
C28 VDD2.n5 B 2.94628f
C29 VN.n0 B 0.028369f
C30 VN.t3 B 2.15265f
C31 VN.n1 B 0.02297f
C32 VN.n2 B 0.028369f
C33 VN.t2 B 2.15265f
C34 VN.n3 B 0.022934f
C35 VN.n4 B 0.179147f
C36 VN.t7 B 2.15265f
C37 VN.t6 B 2.24413f
C38 VN.n5 B 0.840042f
C39 VN.n6 B 0.806254f
C40 VN.n7 B 0.027029f
C41 VN.n8 B 0.056384f
C42 VN.n9 B 0.028369f
C43 VN.n10 B 0.028369f
C44 VN.n11 B 0.028369f
C45 VN.n12 B 0.056384f
C46 VN.n13 B 0.027029f
C47 VN.n14 B 0.758494f
C48 VN.n15 B 0.056387f
C49 VN.n16 B 0.028369f
C50 VN.n17 B 0.028369f
C51 VN.n18 B 0.028369f
C52 VN.n19 B 0.056081f
C53 VN.n20 B 0.027551f
C54 VN.n21 B 0.813459f
C55 VN.n22 B 0.030072f
C56 VN.n23 B 0.028369f
C57 VN.t0 B 2.15265f
C58 VN.n24 B 0.02297f
C59 VN.n25 B 0.028369f
C60 VN.t5 B 2.15265f
C61 VN.n26 B 0.022934f
C62 VN.n27 B 0.179147f
C63 VN.t4 B 2.15265f
C64 VN.t1 B 2.24413f
C65 VN.n28 B 0.840042f
C66 VN.n29 B 0.806254f
C67 VN.n30 B 0.027029f
C68 VN.n31 B 0.056384f
C69 VN.n32 B 0.028369f
C70 VN.n33 B 0.028369f
C71 VN.n34 B 0.028369f
C72 VN.n35 B 0.056384f
C73 VN.n36 B 0.027029f
C74 VN.n37 B 0.758494f
C75 VN.n38 B 0.056387f
C76 VN.n39 B 0.028369f
C77 VN.n40 B 0.028369f
C78 VN.n41 B 0.028369f
C79 VN.n42 B 0.056081f
C80 VN.n43 B 0.027551f
C81 VN.n44 B 0.813459f
C82 VN.n45 B 1.55907f
C83 VDD1.t0 B 0.325666f
C84 VDD1.t7 B 0.325666f
C85 VDD1.n0 B 2.96236f
C86 VDD1.t4 B 0.325666f
C87 VDD1.t1 B 0.325666f
C88 VDD1.n1 B 2.96147f
C89 VDD1.t2 B 0.325666f
C90 VDD1.t3 B 0.325666f
C91 VDD1.n2 B 2.96147f
C92 VDD1.n3 B 3.08136f
C93 VDD1.t6 B 0.325666f
C94 VDD1.t5 B 0.325666f
C95 VDD1.n4 B 2.95591f
C96 VDD1.n5 B 3.00748f
C97 VTAIL.t2 B 0.240732f
C98 VTAIL.t1 B 0.240732f
C99 VTAIL.n0 B 2.1288f
C100 VTAIL.n1 B 0.290623f
C101 VTAIL.t15 B 2.71798f
C102 VTAIL.n2 B 0.382548f
C103 VTAIL.t14 B 2.71798f
C104 VTAIL.n3 B 0.382548f
C105 VTAIL.t8 B 0.240732f
C106 VTAIL.t10 B 0.240732f
C107 VTAIL.n4 B 2.1288f
C108 VTAIL.n5 B 0.390547f
C109 VTAIL.t13 B 2.71798f
C110 VTAIL.n6 B 1.55568f
C111 VTAIL.t6 B 2.71798f
C112 VTAIL.n7 B 1.55567f
C113 VTAIL.t5 B 0.240732f
C114 VTAIL.t4 B 0.240732f
C115 VTAIL.n8 B 2.1288f
C116 VTAIL.n9 B 0.390544f
C117 VTAIL.t0 B 2.71798f
C118 VTAIL.n10 B 0.382545f
C119 VTAIL.t11 B 2.71798f
C120 VTAIL.n11 B 0.382545f
C121 VTAIL.t9 B 0.240732f
C122 VTAIL.t12 B 0.240732f
C123 VTAIL.n12 B 2.1288f
C124 VTAIL.n13 B 0.390544f
C125 VTAIL.t7 B 2.71798f
C126 VTAIL.n14 B 1.55568f
C127 VTAIL.t3 B 2.71798f
C128 VTAIL.n15 B 1.5522f
C129 VP.n0 B 0.028708f
C130 VP.t4 B 2.17836f
C131 VP.n1 B 0.023245f
C132 VP.n2 B 0.028708f
C133 VP.t5 B 2.17836f
C134 VP.n3 B 0.023208f
C135 VP.n4 B 0.028708f
C136 VP.t6 B 2.17836f
C137 VP.n5 B 0.023245f
C138 VP.n6 B 0.028708f
C139 VP.t3 B 2.17836f
C140 VP.n7 B 0.028708f
C141 VP.t2 B 2.17836f
C142 VP.n8 B 0.023245f
C143 VP.n9 B 0.028708f
C144 VP.t1 B 2.17836f
C145 VP.n10 B 0.023208f
C146 VP.n11 B 0.181286f
C147 VP.t0 B 2.17836f
C148 VP.t7 B 2.27093f
C149 VP.n12 B 0.850074f
C150 VP.n13 B 0.815882f
C151 VP.n14 B 0.027352f
C152 VP.n15 B 0.057057f
C153 VP.n16 B 0.028708f
C154 VP.n17 B 0.028708f
C155 VP.n18 B 0.028708f
C156 VP.n19 B 0.057057f
C157 VP.n20 B 0.027352f
C158 VP.n21 B 0.767552f
C159 VP.n22 B 0.057061f
C160 VP.n23 B 0.028708f
C161 VP.n24 B 0.028708f
C162 VP.n25 B 0.028708f
C163 VP.n26 B 0.056751f
C164 VP.n27 B 0.02788f
C165 VP.n28 B 0.823173f
C166 VP.n29 B 1.55902f
C167 VP.n30 B 1.57975f
C168 VP.n31 B 0.823173f
C169 VP.n32 B 0.02788f
C170 VP.n33 B 0.056751f
C171 VP.n34 B 0.028708f
C172 VP.n35 B 0.028708f
C173 VP.n36 B 0.028708f
C174 VP.n37 B 0.057061f
C175 VP.n38 B 0.767552f
C176 VP.n39 B 0.027352f
C177 VP.n40 B 0.057057f
C178 VP.n41 B 0.028708f
C179 VP.n42 B 0.028708f
C180 VP.n43 B 0.028708f
C181 VP.n44 B 0.057057f
C182 VP.n45 B 0.027352f
C183 VP.n46 B 0.767552f
C184 VP.n47 B 0.057061f
C185 VP.n48 B 0.028708f
C186 VP.n49 B 0.028708f
C187 VP.n50 B 0.028708f
C188 VP.n51 B 0.056751f
C189 VP.n52 B 0.02788f
C190 VP.n53 B 0.823173f
C191 VP.n54 B 0.030432f
.ends

