* NGSPICE file created from diff_pair_sample_0905.ext - technology: sky130A

.subckt diff_pair_sample_0905 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=2.5212 ps=15.61 w=15.28 l=0.66
X1 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=0 ps=0 w=15.28 l=0.66
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=0 ps=0 w=15.28 l=0.66
X3 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=2.5212 ps=15.61 w=15.28 l=0.66
X4 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=0 ps=0 w=15.28 l=0.66
X5 VDD2.t2 VN.t1 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5212 pd=15.61 as=5.9592 ps=31.34 w=15.28 l=0.66
X6 VDD1.t2 VP.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5212 pd=15.61 as=5.9592 ps=31.34 w=15.28 l=0.66
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=0 ps=0 w=15.28 l=0.66
X8 VTAIL.t2 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=2.5212 ps=15.61 w=15.28 l=0.66
X9 VTAIL.t5 VP.t2 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.9592 pd=31.34 as=2.5212 ps=15.61 w=15.28 l=0.66
X10 VDD1.t3 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5212 pd=15.61 as=5.9592 ps=31.34 w=15.28 l=0.66
X11 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5212 pd=15.61 as=5.9592 ps=31.34 w=15.28 l=0.66
R0 VP.n1 VP.t2 638.467
R1 VP.n1 VP.t3 638.418
R2 VP.n3 VP.t0 617.471
R3 VP.n5 VP.t1 617.471
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 87.4045
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VDD1 VDD1.n1 99.6952
R14 VDD1 VDD1.n0 59.7812
R15 VDD1.n0 VDD1.t0 1.29631
R16 VDD1.n0 VDD1.t3 1.29631
R17 VDD1.n1 VDD1.t1 1.29631
R18 VDD1.n1 VDD1.t2 1.29631
R19 VTAIL.n6 VTAIL.t4 44.3401
R20 VTAIL.n5 VTAIL.t5 44.34
R21 VTAIL.n4 VTAIL.t3 44.34
R22 VTAIL.n3 VTAIL.t2 44.34
R23 VTAIL.n7 VTAIL.t1 44.3399
R24 VTAIL.n0 VTAIL.t0 44.3399
R25 VTAIL.n1 VTAIL.t6 44.3399
R26 VTAIL.n2 VTAIL.t7 44.3399
R27 VTAIL.n7 VTAIL.n6 26.3927
R28 VTAIL.n3 VTAIL.n2 26.3927
R29 VTAIL.n4 VTAIL.n3 0.853948
R30 VTAIL.n6 VTAIL.n5 0.853948
R31 VTAIL.n2 VTAIL.n1 0.853948
R32 VTAIL VTAIL.n0 0.485414
R33 VTAIL.n5 VTAIL.n4 0.470328
R34 VTAIL.n1 VTAIL.n0 0.470328
R35 VTAIL VTAIL.n7 0.369034
R36 B.n411 B.t4 761.438
R37 B.n408 B.t15 761.438
R38 B.n93 B.t12 761.438
R39 B.n91 B.t8 761.438
R40 B.n709 B.n708 585
R41 B.n317 B.n90 585
R42 B.n316 B.n315 585
R43 B.n314 B.n313 585
R44 B.n312 B.n311 585
R45 B.n310 B.n309 585
R46 B.n308 B.n307 585
R47 B.n306 B.n305 585
R48 B.n304 B.n303 585
R49 B.n302 B.n301 585
R50 B.n300 B.n299 585
R51 B.n298 B.n297 585
R52 B.n296 B.n295 585
R53 B.n294 B.n293 585
R54 B.n292 B.n291 585
R55 B.n290 B.n289 585
R56 B.n288 B.n287 585
R57 B.n286 B.n285 585
R58 B.n284 B.n283 585
R59 B.n282 B.n281 585
R60 B.n280 B.n279 585
R61 B.n278 B.n277 585
R62 B.n276 B.n275 585
R63 B.n274 B.n273 585
R64 B.n272 B.n271 585
R65 B.n270 B.n269 585
R66 B.n268 B.n267 585
R67 B.n266 B.n265 585
R68 B.n264 B.n263 585
R69 B.n262 B.n261 585
R70 B.n260 B.n259 585
R71 B.n258 B.n257 585
R72 B.n256 B.n255 585
R73 B.n254 B.n253 585
R74 B.n252 B.n251 585
R75 B.n250 B.n249 585
R76 B.n248 B.n247 585
R77 B.n246 B.n245 585
R78 B.n244 B.n243 585
R79 B.n242 B.n241 585
R80 B.n240 B.n239 585
R81 B.n238 B.n237 585
R82 B.n236 B.n235 585
R83 B.n234 B.n233 585
R84 B.n232 B.n231 585
R85 B.n230 B.n229 585
R86 B.n228 B.n227 585
R87 B.n226 B.n225 585
R88 B.n224 B.n223 585
R89 B.n222 B.n221 585
R90 B.n220 B.n219 585
R91 B.n217 B.n216 585
R92 B.n215 B.n214 585
R93 B.n213 B.n212 585
R94 B.n211 B.n210 585
R95 B.n209 B.n208 585
R96 B.n207 B.n206 585
R97 B.n205 B.n204 585
R98 B.n203 B.n202 585
R99 B.n201 B.n200 585
R100 B.n199 B.n198 585
R101 B.n196 B.n195 585
R102 B.n194 B.n193 585
R103 B.n192 B.n191 585
R104 B.n190 B.n189 585
R105 B.n188 B.n187 585
R106 B.n186 B.n185 585
R107 B.n184 B.n183 585
R108 B.n182 B.n181 585
R109 B.n180 B.n179 585
R110 B.n178 B.n177 585
R111 B.n176 B.n175 585
R112 B.n174 B.n173 585
R113 B.n172 B.n171 585
R114 B.n170 B.n169 585
R115 B.n168 B.n167 585
R116 B.n166 B.n165 585
R117 B.n164 B.n163 585
R118 B.n162 B.n161 585
R119 B.n160 B.n159 585
R120 B.n158 B.n157 585
R121 B.n156 B.n155 585
R122 B.n154 B.n153 585
R123 B.n152 B.n151 585
R124 B.n150 B.n149 585
R125 B.n148 B.n147 585
R126 B.n146 B.n145 585
R127 B.n144 B.n143 585
R128 B.n142 B.n141 585
R129 B.n140 B.n139 585
R130 B.n138 B.n137 585
R131 B.n136 B.n135 585
R132 B.n134 B.n133 585
R133 B.n132 B.n131 585
R134 B.n130 B.n129 585
R135 B.n128 B.n127 585
R136 B.n126 B.n125 585
R137 B.n124 B.n123 585
R138 B.n122 B.n121 585
R139 B.n120 B.n119 585
R140 B.n118 B.n117 585
R141 B.n116 B.n115 585
R142 B.n114 B.n113 585
R143 B.n112 B.n111 585
R144 B.n110 B.n109 585
R145 B.n108 B.n107 585
R146 B.n106 B.n105 585
R147 B.n104 B.n103 585
R148 B.n102 B.n101 585
R149 B.n100 B.n99 585
R150 B.n98 B.n97 585
R151 B.n96 B.n95 585
R152 B.n707 B.n34 585
R153 B.n712 B.n34 585
R154 B.n706 B.n33 585
R155 B.n713 B.n33 585
R156 B.n705 B.n704 585
R157 B.n704 B.n29 585
R158 B.n703 B.n28 585
R159 B.n719 B.n28 585
R160 B.n702 B.n27 585
R161 B.n720 B.n27 585
R162 B.n701 B.n26 585
R163 B.n721 B.n26 585
R164 B.n700 B.n699 585
R165 B.n699 B.n22 585
R166 B.n698 B.n21 585
R167 B.n727 B.n21 585
R168 B.n697 B.n20 585
R169 B.n728 B.n20 585
R170 B.n696 B.n19 585
R171 B.n729 B.n19 585
R172 B.n695 B.n694 585
R173 B.n694 B.n15 585
R174 B.n693 B.n14 585
R175 B.n735 B.n14 585
R176 B.n692 B.n13 585
R177 B.n736 B.n13 585
R178 B.n691 B.n12 585
R179 B.n737 B.n12 585
R180 B.n690 B.n689 585
R181 B.n689 B.n8 585
R182 B.n688 B.n7 585
R183 B.n743 B.n7 585
R184 B.n687 B.n6 585
R185 B.n744 B.n6 585
R186 B.n686 B.n5 585
R187 B.n745 B.n5 585
R188 B.n685 B.n684 585
R189 B.n684 B.n4 585
R190 B.n683 B.n318 585
R191 B.n683 B.n682 585
R192 B.n673 B.n319 585
R193 B.n320 B.n319 585
R194 B.n675 B.n674 585
R195 B.n676 B.n675 585
R196 B.n672 B.n325 585
R197 B.n325 B.n324 585
R198 B.n671 B.n670 585
R199 B.n670 B.n669 585
R200 B.n327 B.n326 585
R201 B.n328 B.n327 585
R202 B.n662 B.n661 585
R203 B.n663 B.n662 585
R204 B.n660 B.n333 585
R205 B.n333 B.n332 585
R206 B.n659 B.n658 585
R207 B.n658 B.n657 585
R208 B.n335 B.n334 585
R209 B.n336 B.n335 585
R210 B.n650 B.n649 585
R211 B.n651 B.n650 585
R212 B.n648 B.n340 585
R213 B.n344 B.n340 585
R214 B.n647 B.n646 585
R215 B.n646 B.n645 585
R216 B.n342 B.n341 585
R217 B.n343 B.n342 585
R218 B.n638 B.n637 585
R219 B.n639 B.n638 585
R220 B.n636 B.n349 585
R221 B.n349 B.n348 585
R222 B.n631 B.n630 585
R223 B.n629 B.n407 585
R224 B.n628 B.n406 585
R225 B.n633 B.n406 585
R226 B.n627 B.n626 585
R227 B.n625 B.n624 585
R228 B.n623 B.n622 585
R229 B.n621 B.n620 585
R230 B.n619 B.n618 585
R231 B.n617 B.n616 585
R232 B.n615 B.n614 585
R233 B.n613 B.n612 585
R234 B.n611 B.n610 585
R235 B.n609 B.n608 585
R236 B.n607 B.n606 585
R237 B.n605 B.n604 585
R238 B.n603 B.n602 585
R239 B.n601 B.n600 585
R240 B.n599 B.n598 585
R241 B.n597 B.n596 585
R242 B.n595 B.n594 585
R243 B.n593 B.n592 585
R244 B.n591 B.n590 585
R245 B.n589 B.n588 585
R246 B.n587 B.n586 585
R247 B.n585 B.n584 585
R248 B.n583 B.n582 585
R249 B.n581 B.n580 585
R250 B.n579 B.n578 585
R251 B.n577 B.n576 585
R252 B.n575 B.n574 585
R253 B.n573 B.n572 585
R254 B.n571 B.n570 585
R255 B.n569 B.n568 585
R256 B.n567 B.n566 585
R257 B.n565 B.n564 585
R258 B.n563 B.n562 585
R259 B.n561 B.n560 585
R260 B.n559 B.n558 585
R261 B.n557 B.n556 585
R262 B.n555 B.n554 585
R263 B.n553 B.n552 585
R264 B.n551 B.n550 585
R265 B.n549 B.n548 585
R266 B.n547 B.n546 585
R267 B.n545 B.n544 585
R268 B.n543 B.n542 585
R269 B.n541 B.n540 585
R270 B.n539 B.n538 585
R271 B.n537 B.n536 585
R272 B.n535 B.n534 585
R273 B.n533 B.n532 585
R274 B.n531 B.n530 585
R275 B.n529 B.n528 585
R276 B.n527 B.n526 585
R277 B.n525 B.n524 585
R278 B.n523 B.n522 585
R279 B.n521 B.n520 585
R280 B.n519 B.n518 585
R281 B.n517 B.n516 585
R282 B.n515 B.n514 585
R283 B.n513 B.n512 585
R284 B.n511 B.n510 585
R285 B.n509 B.n508 585
R286 B.n507 B.n506 585
R287 B.n505 B.n504 585
R288 B.n503 B.n502 585
R289 B.n501 B.n500 585
R290 B.n499 B.n498 585
R291 B.n497 B.n496 585
R292 B.n495 B.n494 585
R293 B.n493 B.n492 585
R294 B.n491 B.n490 585
R295 B.n489 B.n488 585
R296 B.n487 B.n486 585
R297 B.n485 B.n484 585
R298 B.n483 B.n482 585
R299 B.n481 B.n480 585
R300 B.n479 B.n478 585
R301 B.n477 B.n476 585
R302 B.n475 B.n474 585
R303 B.n473 B.n472 585
R304 B.n471 B.n470 585
R305 B.n469 B.n468 585
R306 B.n467 B.n466 585
R307 B.n465 B.n464 585
R308 B.n463 B.n462 585
R309 B.n461 B.n460 585
R310 B.n459 B.n458 585
R311 B.n457 B.n456 585
R312 B.n455 B.n454 585
R313 B.n453 B.n452 585
R314 B.n451 B.n450 585
R315 B.n449 B.n448 585
R316 B.n447 B.n446 585
R317 B.n445 B.n444 585
R318 B.n443 B.n442 585
R319 B.n441 B.n440 585
R320 B.n439 B.n438 585
R321 B.n437 B.n436 585
R322 B.n435 B.n434 585
R323 B.n433 B.n432 585
R324 B.n431 B.n430 585
R325 B.n429 B.n428 585
R326 B.n427 B.n426 585
R327 B.n425 B.n424 585
R328 B.n423 B.n422 585
R329 B.n421 B.n420 585
R330 B.n419 B.n418 585
R331 B.n417 B.n416 585
R332 B.n415 B.n414 585
R333 B.n351 B.n350 585
R334 B.n635 B.n634 585
R335 B.n634 B.n633 585
R336 B.n347 B.n346 585
R337 B.n348 B.n347 585
R338 B.n641 B.n640 585
R339 B.n640 B.n639 585
R340 B.n642 B.n345 585
R341 B.n345 B.n343 585
R342 B.n644 B.n643 585
R343 B.n645 B.n644 585
R344 B.n339 B.n338 585
R345 B.n344 B.n339 585
R346 B.n653 B.n652 585
R347 B.n652 B.n651 585
R348 B.n654 B.n337 585
R349 B.n337 B.n336 585
R350 B.n656 B.n655 585
R351 B.n657 B.n656 585
R352 B.n331 B.n330 585
R353 B.n332 B.n331 585
R354 B.n665 B.n664 585
R355 B.n664 B.n663 585
R356 B.n666 B.n329 585
R357 B.n329 B.n328 585
R358 B.n668 B.n667 585
R359 B.n669 B.n668 585
R360 B.n323 B.n322 585
R361 B.n324 B.n323 585
R362 B.n678 B.n677 585
R363 B.n677 B.n676 585
R364 B.n679 B.n321 585
R365 B.n321 B.n320 585
R366 B.n681 B.n680 585
R367 B.n682 B.n681 585
R368 B.n2 B.n0 585
R369 B.n4 B.n2 585
R370 B.n3 B.n1 585
R371 B.n744 B.n3 585
R372 B.n742 B.n741 585
R373 B.n743 B.n742 585
R374 B.n740 B.n9 585
R375 B.n9 B.n8 585
R376 B.n739 B.n738 585
R377 B.n738 B.n737 585
R378 B.n11 B.n10 585
R379 B.n736 B.n11 585
R380 B.n734 B.n733 585
R381 B.n735 B.n734 585
R382 B.n732 B.n16 585
R383 B.n16 B.n15 585
R384 B.n731 B.n730 585
R385 B.n730 B.n729 585
R386 B.n18 B.n17 585
R387 B.n728 B.n18 585
R388 B.n726 B.n725 585
R389 B.n727 B.n726 585
R390 B.n724 B.n23 585
R391 B.n23 B.n22 585
R392 B.n723 B.n722 585
R393 B.n722 B.n721 585
R394 B.n25 B.n24 585
R395 B.n720 B.n25 585
R396 B.n718 B.n717 585
R397 B.n719 B.n718 585
R398 B.n716 B.n30 585
R399 B.n30 B.n29 585
R400 B.n715 B.n714 585
R401 B.n714 B.n713 585
R402 B.n32 B.n31 585
R403 B.n712 B.n32 585
R404 B.n747 B.n746 585
R405 B.n746 B.n745 585
R406 B.n631 B.n347 482.89
R407 B.n95 B.n32 482.89
R408 B.n634 B.n349 482.89
R409 B.n709 B.n34 482.89
R410 B.n711 B.n710 256.663
R411 B.n711 B.n89 256.663
R412 B.n711 B.n88 256.663
R413 B.n711 B.n87 256.663
R414 B.n711 B.n86 256.663
R415 B.n711 B.n85 256.663
R416 B.n711 B.n84 256.663
R417 B.n711 B.n83 256.663
R418 B.n711 B.n82 256.663
R419 B.n711 B.n81 256.663
R420 B.n711 B.n80 256.663
R421 B.n711 B.n79 256.663
R422 B.n711 B.n78 256.663
R423 B.n711 B.n77 256.663
R424 B.n711 B.n76 256.663
R425 B.n711 B.n75 256.663
R426 B.n711 B.n74 256.663
R427 B.n711 B.n73 256.663
R428 B.n711 B.n72 256.663
R429 B.n711 B.n71 256.663
R430 B.n711 B.n70 256.663
R431 B.n711 B.n69 256.663
R432 B.n711 B.n68 256.663
R433 B.n711 B.n67 256.663
R434 B.n711 B.n66 256.663
R435 B.n711 B.n65 256.663
R436 B.n711 B.n64 256.663
R437 B.n711 B.n63 256.663
R438 B.n711 B.n62 256.663
R439 B.n711 B.n61 256.663
R440 B.n711 B.n60 256.663
R441 B.n711 B.n59 256.663
R442 B.n711 B.n58 256.663
R443 B.n711 B.n57 256.663
R444 B.n711 B.n56 256.663
R445 B.n711 B.n55 256.663
R446 B.n711 B.n54 256.663
R447 B.n711 B.n53 256.663
R448 B.n711 B.n52 256.663
R449 B.n711 B.n51 256.663
R450 B.n711 B.n50 256.663
R451 B.n711 B.n49 256.663
R452 B.n711 B.n48 256.663
R453 B.n711 B.n47 256.663
R454 B.n711 B.n46 256.663
R455 B.n711 B.n45 256.663
R456 B.n711 B.n44 256.663
R457 B.n711 B.n43 256.663
R458 B.n711 B.n42 256.663
R459 B.n711 B.n41 256.663
R460 B.n711 B.n40 256.663
R461 B.n711 B.n39 256.663
R462 B.n711 B.n38 256.663
R463 B.n711 B.n37 256.663
R464 B.n711 B.n36 256.663
R465 B.n711 B.n35 256.663
R466 B.n633 B.n632 256.663
R467 B.n633 B.n352 256.663
R468 B.n633 B.n353 256.663
R469 B.n633 B.n354 256.663
R470 B.n633 B.n355 256.663
R471 B.n633 B.n356 256.663
R472 B.n633 B.n357 256.663
R473 B.n633 B.n358 256.663
R474 B.n633 B.n359 256.663
R475 B.n633 B.n360 256.663
R476 B.n633 B.n361 256.663
R477 B.n633 B.n362 256.663
R478 B.n633 B.n363 256.663
R479 B.n633 B.n364 256.663
R480 B.n633 B.n365 256.663
R481 B.n633 B.n366 256.663
R482 B.n633 B.n367 256.663
R483 B.n633 B.n368 256.663
R484 B.n633 B.n369 256.663
R485 B.n633 B.n370 256.663
R486 B.n633 B.n371 256.663
R487 B.n633 B.n372 256.663
R488 B.n633 B.n373 256.663
R489 B.n633 B.n374 256.663
R490 B.n633 B.n375 256.663
R491 B.n633 B.n376 256.663
R492 B.n633 B.n377 256.663
R493 B.n633 B.n378 256.663
R494 B.n633 B.n379 256.663
R495 B.n633 B.n380 256.663
R496 B.n633 B.n381 256.663
R497 B.n633 B.n382 256.663
R498 B.n633 B.n383 256.663
R499 B.n633 B.n384 256.663
R500 B.n633 B.n385 256.663
R501 B.n633 B.n386 256.663
R502 B.n633 B.n387 256.663
R503 B.n633 B.n388 256.663
R504 B.n633 B.n389 256.663
R505 B.n633 B.n390 256.663
R506 B.n633 B.n391 256.663
R507 B.n633 B.n392 256.663
R508 B.n633 B.n393 256.663
R509 B.n633 B.n394 256.663
R510 B.n633 B.n395 256.663
R511 B.n633 B.n396 256.663
R512 B.n633 B.n397 256.663
R513 B.n633 B.n398 256.663
R514 B.n633 B.n399 256.663
R515 B.n633 B.n400 256.663
R516 B.n633 B.n401 256.663
R517 B.n633 B.n402 256.663
R518 B.n633 B.n403 256.663
R519 B.n633 B.n404 256.663
R520 B.n633 B.n405 256.663
R521 B.n640 B.n347 163.367
R522 B.n640 B.n345 163.367
R523 B.n644 B.n345 163.367
R524 B.n644 B.n339 163.367
R525 B.n652 B.n339 163.367
R526 B.n652 B.n337 163.367
R527 B.n656 B.n337 163.367
R528 B.n656 B.n331 163.367
R529 B.n664 B.n331 163.367
R530 B.n664 B.n329 163.367
R531 B.n668 B.n329 163.367
R532 B.n668 B.n323 163.367
R533 B.n677 B.n323 163.367
R534 B.n677 B.n321 163.367
R535 B.n681 B.n321 163.367
R536 B.n681 B.n2 163.367
R537 B.n746 B.n2 163.367
R538 B.n746 B.n3 163.367
R539 B.n742 B.n3 163.367
R540 B.n742 B.n9 163.367
R541 B.n738 B.n9 163.367
R542 B.n738 B.n11 163.367
R543 B.n734 B.n11 163.367
R544 B.n734 B.n16 163.367
R545 B.n730 B.n16 163.367
R546 B.n730 B.n18 163.367
R547 B.n726 B.n18 163.367
R548 B.n726 B.n23 163.367
R549 B.n722 B.n23 163.367
R550 B.n722 B.n25 163.367
R551 B.n718 B.n25 163.367
R552 B.n718 B.n30 163.367
R553 B.n714 B.n30 163.367
R554 B.n714 B.n32 163.367
R555 B.n407 B.n406 163.367
R556 B.n626 B.n406 163.367
R557 B.n624 B.n623 163.367
R558 B.n620 B.n619 163.367
R559 B.n616 B.n615 163.367
R560 B.n612 B.n611 163.367
R561 B.n608 B.n607 163.367
R562 B.n604 B.n603 163.367
R563 B.n600 B.n599 163.367
R564 B.n596 B.n595 163.367
R565 B.n592 B.n591 163.367
R566 B.n588 B.n587 163.367
R567 B.n584 B.n583 163.367
R568 B.n580 B.n579 163.367
R569 B.n576 B.n575 163.367
R570 B.n572 B.n571 163.367
R571 B.n568 B.n567 163.367
R572 B.n564 B.n563 163.367
R573 B.n560 B.n559 163.367
R574 B.n556 B.n555 163.367
R575 B.n552 B.n551 163.367
R576 B.n548 B.n547 163.367
R577 B.n544 B.n543 163.367
R578 B.n540 B.n539 163.367
R579 B.n536 B.n535 163.367
R580 B.n532 B.n531 163.367
R581 B.n528 B.n527 163.367
R582 B.n524 B.n523 163.367
R583 B.n520 B.n519 163.367
R584 B.n516 B.n515 163.367
R585 B.n512 B.n511 163.367
R586 B.n508 B.n507 163.367
R587 B.n504 B.n503 163.367
R588 B.n500 B.n499 163.367
R589 B.n496 B.n495 163.367
R590 B.n492 B.n491 163.367
R591 B.n488 B.n487 163.367
R592 B.n484 B.n483 163.367
R593 B.n480 B.n479 163.367
R594 B.n476 B.n475 163.367
R595 B.n472 B.n471 163.367
R596 B.n468 B.n467 163.367
R597 B.n464 B.n463 163.367
R598 B.n460 B.n459 163.367
R599 B.n456 B.n455 163.367
R600 B.n452 B.n451 163.367
R601 B.n448 B.n447 163.367
R602 B.n444 B.n443 163.367
R603 B.n440 B.n439 163.367
R604 B.n436 B.n435 163.367
R605 B.n432 B.n431 163.367
R606 B.n428 B.n427 163.367
R607 B.n424 B.n423 163.367
R608 B.n420 B.n419 163.367
R609 B.n416 B.n415 163.367
R610 B.n634 B.n351 163.367
R611 B.n638 B.n349 163.367
R612 B.n638 B.n342 163.367
R613 B.n646 B.n342 163.367
R614 B.n646 B.n340 163.367
R615 B.n650 B.n340 163.367
R616 B.n650 B.n335 163.367
R617 B.n658 B.n335 163.367
R618 B.n658 B.n333 163.367
R619 B.n662 B.n333 163.367
R620 B.n662 B.n327 163.367
R621 B.n670 B.n327 163.367
R622 B.n670 B.n325 163.367
R623 B.n675 B.n325 163.367
R624 B.n675 B.n319 163.367
R625 B.n683 B.n319 163.367
R626 B.n684 B.n683 163.367
R627 B.n684 B.n5 163.367
R628 B.n6 B.n5 163.367
R629 B.n7 B.n6 163.367
R630 B.n689 B.n7 163.367
R631 B.n689 B.n12 163.367
R632 B.n13 B.n12 163.367
R633 B.n14 B.n13 163.367
R634 B.n694 B.n14 163.367
R635 B.n694 B.n19 163.367
R636 B.n20 B.n19 163.367
R637 B.n21 B.n20 163.367
R638 B.n699 B.n21 163.367
R639 B.n699 B.n26 163.367
R640 B.n27 B.n26 163.367
R641 B.n28 B.n27 163.367
R642 B.n704 B.n28 163.367
R643 B.n704 B.n33 163.367
R644 B.n34 B.n33 163.367
R645 B.n99 B.n98 163.367
R646 B.n103 B.n102 163.367
R647 B.n107 B.n106 163.367
R648 B.n111 B.n110 163.367
R649 B.n115 B.n114 163.367
R650 B.n119 B.n118 163.367
R651 B.n123 B.n122 163.367
R652 B.n127 B.n126 163.367
R653 B.n131 B.n130 163.367
R654 B.n135 B.n134 163.367
R655 B.n139 B.n138 163.367
R656 B.n143 B.n142 163.367
R657 B.n147 B.n146 163.367
R658 B.n151 B.n150 163.367
R659 B.n155 B.n154 163.367
R660 B.n159 B.n158 163.367
R661 B.n163 B.n162 163.367
R662 B.n167 B.n166 163.367
R663 B.n171 B.n170 163.367
R664 B.n175 B.n174 163.367
R665 B.n179 B.n178 163.367
R666 B.n183 B.n182 163.367
R667 B.n187 B.n186 163.367
R668 B.n191 B.n190 163.367
R669 B.n195 B.n194 163.367
R670 B.n200 B.n199 163.367
R671 B.n204 B.n203 163.367
R672 B.n208 B.n207 163.367
R673 B.n212 B.n211 163.367
R674 B.n216 B.n215 163.367
R675 B.n221 B.n220 163.367
R676 B.n225 B.n224 163.367
R677 B.n229 B.n228 163.367
R678 B.n233 B.n232 163.367
R679 B.n237 B.n236 163.367
R680 B.n241 B.n240 163.367
R681 B.n245 B.n244 163.367
R682 B.n249 B.n248 163.367
R683 B.n253 B.n252 163.367
R684 B.n257 B.n256 163.367
R685 B.n261 B.n260 163.367
R686 B.n265 B.n264 163.367
R687 B.n269 B.n268 163.367
R688 B.n273 B.n272 163.367
R689 B.n277 B.n276 163.367
R690 B.n281 B.n280 163.367
R691 B.n285 B.n284 163.367
R692 B.n289 B.n288 163.367
R693 B.n293 B.n292 163.367
R694 B.n297 B.n296 163.367
R695 B.n301 B.n300 163.367
R696 B.n305 B.n304 163.367
R697 B.n309 B.n308 163.367
R698 B.n313 B.n312 163.367
R699 B.n315 B.n90 163.367
R700 B.n411 B.t7 92.8463
R701 B.n91 B.t10 92.8463
R702 B.n408 B.t17 92.8265
R703 B.n93 B.t13 92.8265
R704 B.n412 B.t6 73.6463
R705 B.n92 B.t11 73.6463
R706 B.n409 B.t16 73.6265
R707 B.n94 B.t14 73.6265
R708 B.n632 B.n631 71.676
R709 B.n626 B.n352 71.676
R710 B.n623 B.n353 71.676
R711 B.n619 B.n354 71.676
R712 B.n615 B.n355 71.676
R713 B.n611 B.n356 71.676
R714 B.n607 B.n357 71.676
R715 B.n603 B.n358 71.676
R716 B.n599 B.n359 71.676
R717 B.n595 B.n360 71.676
R718 B.n591 B.n361 71.676
R719 B.n587 B.n362 71.676
R720 B.n583 B.n363 71.676
R721 B.n579 B.n364 71.676
R722 B.n575 B.n365 71.676
R723 B.n571 B.n366 71.676
R724 B.n567 B.n367 71.676
R725 B.n563 B.n368 71.676
R726 B.n559 B.n369 71.676
R727 B.n555 B.n370 71.676
R728 B.n551 B.n371 71.676
R729 B.n547 B.n372 71.676
R730 B.n543 B.n373 71.676
R731 B.n539 B.n374 71.676
R732 B.n535 B.n375 71.676
R733 B.n531 B.n376 71.676
R734 B.n527 B.n377 71.676
R735 B.n523 B.n378 71.676
R736 B.n519 B.n379 71.676
R737 B.n515 B.n380 71.676
R738 B.n511 B.n381 71.676
R739 B.n507 B.n382 71.676
R740 B.n503 B.n383 71.676
R741 B.n499 B.n384 71.676
R742 B.n495 B.n385 71.676
R743 B.n491 B.n386 71.676
R744 B.n487 B.n387 71.676
R745 B.n483 B.n388 71.676
R746 B.n479 B.n389 71.676
R747 B.n475 B.n390 71.676
R748 B.n471 B.n391 71.676
R749 B.n467 B.n392 71.676
R750 B.n463 B.n393 71.676
R751 B.n459 B.n394 71.676
R752 B.n455 B.n395 71.676
R753 B.n451 B.n396 71.676
R754 B.n447 B.n397 71.676
R755 B.n443 B.n398 71.676
R756 B.n439 B.n399 71.676
R757 B.n435 B.n400 71.676
R758 B.n431 B.n401 71.676
R759 B.n427 B.n402 71.676
R760 B.n423 B.n403 71.676
R761 B.n419 B.n404 71.676
R762 B.n415 B.n405 71.676
R763 B.n95 B.n35 71.676
R764 B.n99 B.n36 71.676
R765 B.n103 B.n37 71.676
R766 B.n107 B.n38 71.676
R767 B.n111 B.n39 71.676
R768 B.n115 B.n40 71.676
R769 B.n119 B.n41 71.676
R770 B.n123 B.n42 71.676
R771 B.n127 B.n43 71.676
R772 B.n131 B.n44 71.676
R773 B.n135 B.n45 71.676
R774 B.n139 B.n46 71.676
R775 B.n143 B.n47 71.676
R776 B.n147 B.n48 71.676
R777 B.n151 B.n49 71.676
R778 B.n155 B.n50 71.676
R779 B.n159 B.n51 71.676
R780 B.n163 B.n52 71.676
R781 B.n167 B.n53 71.676
R782 B.n171 B.n54 71.676
R783 B.n175 B.n55 71.676
R784 B.n179 B.n56 71.676
R785 B.n183 B.n57 71.676
R786 B.n187 B.n58 71.676
R787 B.n191 B.n59 71.676
R788 B.n195 B.n60 71.676
R789 B.n200 B.n61 71.676
R790 B.n204 B.n62 71.676
R791 B.n208 B.n63 71.676
R792 B.n212 B.n64 71.676
R793 B.n216 B.n65 71.676
R794 B.n221 B.n66 71.676
R795 B.n225 B.n67 71.676
R796 B.n229 B.n68 71.676
R797 B.n233 B.n69 71.676
R798 B.n237 B.n70 71.676
R799 B.n241 B.n71 71.676
R800 B.n245 B.n72 71.676
R801 B.n249 B.n73 71.676
R802 B.n253 B.n74 71.676
R803 B.n257 B.n75 71.676
R804 B.n261 B.n76 71.676
R805 B.n265 B.n77 71.676
R806 B.n269 B.n78 71.676
R807 B.n273 B.n79 71.676
R808 B.n277 B.n80 71.676
R809 B.n281 B.n81 71.676
R810 B.n285 B.n82 71.676
R811 B.n289 B.n83 71.676
R812 B.n293 B.n84 71.676
R813 B.n297 B.n85 71.676
R814 B.n301 B.n86 71.676
R815 B.n305 B.n87 71.676
R816 B.n309 B.n88 71.676
R817 B.n313 B.n89 71.676
R818 B.n710 B.n90 71.676
R819 B.n710 B.n709 71.676
R820 B.n315 B.n89 71.676
R821 B.n312 B.n88 71.676
R822 B.n308 B.n87 71.676
R823 B.n304 B.n86 71.676
R824 B.n300 B.n85 71.676
R825 B.n296 B.n84 71.676
R826 B.n292 B.n83 71.676
R827 B.n288 B.n82 71.676
R828 B.n284 B.n81 71.676
R829 B.n280 B.n80 71.676
R830 B.n276 B.n79 71.676
R831 B.n272 B.n78 71.676
R832 B.n268 B.n77 71.676
R833 B.n264 B.n76 71.676
R834 B.n260 B.n75 71.676
R835 B.n256 B.n74 71.676
R836 B.n252 B.n73 71.676
R837 B.n248 B.n72 71.676
R838 B.n244 B.n71 71.676
R839 B.n240 B.n70 71.676
R840 B.n236 B.n69 71.676
R841 B.n232 B.n68 71.676
R842 B.n228 B.n67 71.676
R843 B.n224 B.n66 71.676
R844 B.n220 B.n65 71.676
R845 B.n215 B.n64 71.676
R846 B.n211 B.n63 71.676
R847 B.n207 B.n62 71.676
R848 B.n203 B.n61 71.676
R849 B.n199 B.n60 71.676
R850 B.n194 B.n59 71.676
R851 B.n190 B.n58 71.676
R852 B.n186 B.n57 71.676
R853 B.n182 B.n56 71.676
R854 B.n178 B.n55 71.676
R855 B.n174 B.n54 71.676
R856 B.n170 B.n53 71.676
R857 B.n166 B.n52 71.676
R858 B.n162 B.n51 71.676
R859 B.n158 B.n50 71.676
R860 B.n154 B.n49 71.676
R861 B.n150 B.n48 71.676
R862 B.n146 B.n47 71.676
R863 B.n142 B.n46 71.676
R864 B.n138 B.n45 71.676
R865 B.n134 B.n44 71.676
R866 B.n130 B.n43 71.676
R867 B.n126 B.n42 71.676
R868 B.n122 B.n41 71.676
R869 B.n118 B.n40 71.676
R870 B.n114 B.n39 71.676
R871 B.n110 B.n38 71.676
R872 B.n106 B.n37 71.676
R873 B.n102 B.n36 71.676
R874 B.n98 B.n35 71.676
R875 B.n632 B.n407 71.676
R876 B.n624 B.n352 71.676
R877 B.n620 B.n353 71.676
R878 B.n616 B.n354 71.676
R879 B.n612 B.n355 71.676
R880 B.n608 B.n356 71.676
R881 B.n604 B.n357 71.676
R882 B.n600 B.n358 71.676
R883 B.n596 B.n359 71.676
R884 B.n592 B.n360 71.676
R885 B.n588 B.n361 71.676
R886 B.n584 B.n362 71.676
R887 B.n580 B.n363 71.676
R888 B.n576 B.n364 71.676
R889 B.n572 B.n365 71.676
R890 B.n568 B.n366 71.676
R891 B.n564 B.n367 71.676
R892 B.n560 B.n368 71.676
R893 B.n556 B.n369 71.676
R894 B.n552 B.n370 71.676
R895 B.n548 B.n371 71.676
R896 B.n544 B.n372 71.676
R897 B.n540 B.n373 71.676
R898 B.n536 B.n374 71.676
R899 B.n532 B.n375 71.676
R900 B.n528 B.n376 71.676
R901 B.n524 B.n377 71.676
R902 B.n520 B.n378 71.676
R903 B.n516 B.n379 71.676
R904 B.n512 B.n380 71.676
R905 B.n508 B.n381 71.676
R906 B.n504 B.n382 71.676
R907 B.n500 B.n383 71.676
R908 B.n496 B.n384 71.676
R909 B.n492 B.n385 71.676
R910 B.n488 B.n386 71.676
R911 B.n484 B.n387 71.676
R912 B.n480 B.n388 71.676
R913 B.n476 B.n389 71.676
R914 B.n472 B.n390 71.676
R915 B.n468 B.n391 71.676
R916 B.n464 B.n392 71.676
R917 B.n460 B.n393 71.676
R918 B.n456 B.n394 71.676
R919 B.n452 B.n395 71.676
R920 B.n448 B.n396 71.676
R921 B.n444 B.n397 71.676
R922 B.n440 B.n398 71.676
R923 B.n436 B.n399 71.676
R924 B.n432 B.n400 71.676
R925 B.n428 B.n401 71.676
R926 B.n424 B.n402 71.676
R927 B.n420 B.n403 71.676
R928 B.n416 B.n404 71.676
R929 B.n405 B.n351 71.676
R930 B.n633 B.n348 60.4724
R931 B.n712 B.n711 60.4724
R932 B.n413 B.n412 59.5399
R933 B.n410 B.n409 59.5399
R934 B.n197 B.n94 59.5399
R935 B.n218 B.n92 59.5399
R936 B.n639 B.n348 36.3907
R937 B.n639 B.n343 36.3907
R938 B.n645 B.n343 36.3907
R939 B.n645 B.n344 36.3907
R940 B.n651 B.n336 36.3907
R941 B.n657 B.n336 36.3907
R942 B.n657 B.n332 36.3907
R943 B.n663 B.n332 36.3907
R944 B.n663 B.n328 36.3907
R945 B.n669 B.n328 36.3907
R946 B.n676 B.n324 36.3907
R947 B.n682 B.n320 36.3907
R948 B.n682 B.n4 36.3907
R949 B.n745 B.n4 36.3907
R950 B.n745 B.n744 36.3907
R951 B.n744 B.n743 36.3907
R952 B.n743 B.n8 36.3907
R953 B.n737 B.n736 36.3907
R954 B.n735 B.n15 36.3907
R955 B.n729 B.n15 36.3907
R956 B.n729 B.n728 36.3907
R957 B.n728 B.n727 36.3907
R958 B.n727 B.n22 36.3907
R959 B.n721 B.n22 36.3907
R960 B.n720 B.n719 36.3907
R961 B.n719 B.n29 36.3907
R962 B.n713 B.n29 36.3907
R963 B.n713 B.n712 36.3907
R964 B.t2 B.n324 35.3204
R965 B.n736 B.t1 35.3204
R966 B.n676 B.t3 34.2501
R967 B.n737 B.t0 34.2501
R968 B.n344 B.t5 33.1798
R969 B.t9 B.n720 33.1798
R970 B.n96 B.n31 31.3761
R971 B.n708 B.n707 31.3761
R972 B.n636 B.n635 31.3761
R973 B.n630 B.n346 31.3761
R974 B.n412 B.n411 19.2005
R975 B.n409 B.n408 19.2005
R976 B.n94 B.n93 19.2005
R977 B.n92 B.n91 19.2005
R978 B B.n747 18.0485
R979 B.n97 B.n96 10.6151
R980 B.n100 B.n97 10.6151
R981 B.n101 B.n100 10.6151
R982 B.n104 B.n101 10.6151
R983 B.n105 B.n104 10.6151
R984 B.n108 B.n105 10.6151
R985 B.n109 B.n108 10.6151
R986 B.n112 B.n109 10.6151
R987 B.n113 B.n112 10.6151
R988 B.n116 B.n113 10.6151
R989 B.n117 B.n116 10.6151
R990 B.n120 B.n117 10.6151
R991 B.n121 B.n120 10.6151
R992 B.n124 B.n121 10.6151
R993 B.n125 B.n124 10.6151
R994 B.n128 B.n125 10.6151
R995 B.n129 B.n128 10.6151
R996 B.n132 B.n129 10.6151
R997 B.n133 B.n132 10.6151
R998 B.n136 B.n133 10.6151
R999 B.n137 B.n136 10.6151
R1000 B.n140 B.n137 10.6151
R1001 B.n141 B.n140 10.6151
R1002 B.n144 B.n141 10.6151
R1003 B.n145 B.n144 10.6151
R1004 B.n148 B.n145 10.6151
R1005 B.n149 B.n148 10.6151
R1006 B.n152 B.n149 10.6151
R1007 B.n153 B.n152 10.6151
R1008 B.n156 B.n153 10.6151
R1009 B.n157 B.n156 10.6151
R1010 B.n160 B.n157 10.6151
R1011 B.n161 B.n160 10.6151
R1012 B.n164 B.n161 10.6151
R1013 B.n165 B.n164 10.6151
R1014 B.n168 B.n165 10.6151
R1015 B.n169 B.n168 10.6151
R1016 B.n172 B.n169 10.6151
R1017 B.n173 B.n172 10.6151
R1018 B.n176 B.n173 10.6151
R1019 B.n177 B.n176 10.6151
R1020 B.n180 B.n177 10.6151
R1021 B.n181 B.n180 10.6151
R1022 B.n184 B.n181 10.6151
R1023 B.n185 B.n184 10.6151
R1024 B.n188 B.n185 10.6151
R1025 B.n189 B.n188 10.6151
R1026 B.n192 B.n189 10.6151
R1027 B.n193 B.n192 10.6151
R1028 B.n196 B.n193 10.6151
R1029 B.n201 B.n198 10.6151
R1030 B.n202 B.n201 10.6151
R1031 B.n205 B.n202 10.6151
R1032 B.n206 B.n205 10.6151
R1033 B.n209 B.n206 10.6151
R1034 B.n210 B.n209 10.6151
R1035 B.n213 B.n210 10.6151
R1036 B.n214 B.n213 10.6151
R1037 B.n217 B.n214 10.6151
R1038 B.n222 B.n219 10.6151
R1039 B.n223 B.n222 10.6151
R1040 B.n226 B.n223 10.6151
R1041 B.n227 B.n226 10.6151
R1042 B.n230 B.n227 10.6151
R1043 B.n231 B.n230 10.6151
R1044 B.n234 B.n231 10.6151
R1045 B.n235 B.n234 10.6151
R1046 B.n238 B.n235 10.6151
R1047 B.n239 B.n238 10.6151
R1048 B.n242 B.n239 10.6151
R1049 B.n243 B.n242 10.6151
R1050 B.n246 B.n243 10.6151
R1051 B.n247 B.n246 10.6151
R1052 B.n250 B.n247 10.6151
R1053 B.n251 B.n250 10.6151
R1054 B.n254 B.n251 10.6151
R1055 B.n255 B.n254 10.6151
R1056 B.n258 B.n255 10.6151
R1057 B.n259 B.n258 10.6151
R1058 B.n262 B.n259 10.6151
R1059 B.n263 B.n262 10.6151
R1060 B.n266 B.n263 10.6151
R1061 B.n267 B.n266 10.6151
R1062 B.n270 B.n267 10.6151
R1063 B.n271 B.n270 10.6151
R1064 B.n274 B.n271 10.6151
R1065 B.n275 B.n274 10.6151
R1066 B.n278 B.n275 10.6151
R1067 B.n279 B.n278 10.6151
R1068 B.n282 B.n279 10.6151
R1069 B.n283 B.n282 10.6151
R1070 B.n286 B.n283 10.6151
R1071 B.n287 B.n286 10.6151
R1072 B.n290 B.n287 10.6151
R1073 B.n291 B.n290 10.6151
R1074 B.n294 B.n291 10.6151
R1075 B.n295 B.n294 10.6151
R1076 B.n298 B.n295 10.6151
R1077 B.n299 B.n298 10.6151
R1078 B.n302 B.n299 10.6151
R1079 B.n303 B.n302 10.6151
R1080 B.n306 B.n303 10.6151
R1081 B.n307 B.n306 10.6151
R1082 B.n310 B.n307 10.6151
R1083 B.n311 B.n310 10.6151
R1084 B.n314 B.n311 10.6151
R1085 B.n316 B.n314 10.6151
R1086 B.n317 B.n316 10.6151
R1087 B.n708 B.n317 10.6151
R1088 B.n637 B.n636 10.6151
R1089 B.n637 B.n341 10.6151
R1090 B.n647 B.n341 10.6151
R1091 B.n648 B.n647 10.6151
R1092 B.n649 B.n648 10.6151
R1093 B.n649 B.n334 10.6151
R1094 B.n659 B.n334 10.6151
R1095 B.n660 B.n659 10.6151
R1096 B.n661 B.n660 10.6151
R1097 B.n661 B.n326 10.6151
R1098 B.n671 B.n326 10.6151
R1099 B.n672 B.n671 10.6151
R1100 B.n674 B.n672 10.6151
R1101 B.n674 B.n673 10.6151
R1102 B.n673 B.n318 10.6151
R1103 B.n685 B.n318 10.6151
R1104 B.n686 B.n685 10.6151
R1105 B.n687 B.n686 10.6151
R1106 B.n688 B.n687 10.6151
R1107 B.n690 B.n688 10.6151
R1108 B.n691 B.n690 10.6151
R1109 B.n692 B.n691 10.6151
R1110 B.n693 B.n692 10.6151
R1111 B.n695 B.n693 10.6151
R1112 B.n696 B.n695 10.6151
R1113 B.n697 B.n696 10.6151
R1114 B.n698 B.n697 10.6151
R1115 B.n700 B.n698 10.6151
R1116 B.n701 B.n700 10.6151
R1117 B.n702 B.n701 10.6151
R1118 B.n703 B.n702 10.6151
R1119 B.n705 B.n703 10.6151
R1120 B.n706 B.n705 10.6151
R1121 B.n707 B.n706 10.6151
R1122 B.n630 B.n629 10.6151
R1123 B.n629 B.n628 10.6151
R1124 B.n628 B.n627 10.6151
R1125 B.n627 B.n625 10.6151
R1126 B.n625 B.n622 10.6151
R1127 B.n622 B.n621 10.6151
R1128 B.n621 B.n618 10.6151
R1129 B.n618 B.n617 10.6151
R1130 B.n617 B.n614 10.6151
R1131 B.n614 B.n613 10.6151
R1132 B.n613 B.n610 10.6151
R1133 B.n610 B.n609 10.6151
R1134 B.n609 B.n606 10.6151
R1135 B.n606 B.n605 10.6151
R1136 B.n605 B.n602 10.6151
R1137 B.n602 B.n601 10.6151
R1138 B.n601 B.n598 10.6151
R1139 B.n598 B.n597 10.6151
R1140 B.n597 B.n594 10.6151
R1141 B.n594 B.n593 10.6151
R1142 B.n593 B.n590 10.6151
R1143 B.n590 B.n589 10.6151
R1144 B.n589 B.n586 10.6151
R1145 B.n586 B.n585 10.6151
R1146 B.n585 B.n582 10.6151
R1147 B.n582 B.n581 10.6151
R1148 B.n581 B.n578 10.6151
R1149 B.n578 B.n577 10.6151
R1150 B.n577 B.n574 10.6151
R1151 B.n574 B.n573 10.6151
R1152 B.n573 B.n570 10.6151
R1153 B.n570 B.n569 10.6151
R1154 B.n569 B.n566 10.6151
R1155 B.n566 B.n565 10.6151
R1156 B.n565 B.n562 10.6151
R1157 B.n562 B.n561 10.6151
R1158 B.n561 B.n558 10.6151
R1159 B.n558 B.n557 10.6151
R1160 B.n557 B.n554 10.6151
R1161 B.n554 B.n553 10.6151
R1162 B.n553 B.n550 10.6151
R1163 B.n550 B.n549 10.6151
R1164 B.n549 B.n546 10.6151
R1165 B.n546 B.n545 10.6151
R1166 B.n545 B.n542 10.6151
R1167 B.n542 B.n541 10.6151
R1168 B.n541 B.n538 10.6151
R1169 B.n538 B.n537 10.6151
R1170 B.n537 B.n534 10.6151
R1171 B.n534 B.n533 10.6151
R1172 B.n530 B.n529 10.6151
R1173 B.n529 B.n526 10.6151
R1174 B.n526 B.n525 10.6151
R1175 B.n525 B.n522 10.6151
R1176 B.n522 B.n521 10.6151
R1177 B.n521 B.n518 10.6151
R1178 B.n518 B.n517 10.6151
R1179 B.n517 B.n514 10.6151
R1180 B.n514 B.n513 10.6151
R1181 B.n510 B.n509 10.6151
R1182 B.n509 B.n506 10.6151
R1183 B.n506 B.n505 10.6151
R1184 B.n505 B.n502 10.6151
R1185 B.n502 B.n501 10.6151
R1186 B.n501 B.n498 10.6151
R1187 B.n498 B.n497 10.6151
R1188 B.n497 B.n494 10.6151
R1189 B.n494 B.n493 10.6151
R1190 B.n493 B.n490 10.6151
R1191 B.n490 B.n489 10.6151
R1192 B.n489 B.n486 10.6151
R1193 B.n486 B.n485 10.6151
R1194 B.n485 B.n482 10.6151
R1195 B.n482 B.n481 10.6151
R1196 B.n481 B.n478 10.6151
R1197 B.n478 B.n477 10.6151
R1198 B.n477 B.n474 10.6151
R1199 B.n474 B.n473 10.6151
R1200 B.n473 B.n470 10.6151
R1201 B.n470 B.n469 10.6151
R1202 B.n469 B.n466 10.6151
R1203 B.n466 B.n465 10.6151
R1204 B.n465 B.n462 10.6151
R1205 B.n462 B.n461 10.6151
R1206 B.n461 B.n458 10.6151
R1207 B.n458 B.n457 10.6151
R1208 B.n457 B.n454 10.6151
R1209 B.n454 B.n453 10.6151
R1210 B.n453 B.n450 10.6151
R1211 B.n450 B.n449 10.6151
R1212 B.n449 B.n446 10.6151
R1213 B.n446 B.n445 10.6151
R1214 B.n445 B.n442 10.6151
R1215 B.n442 B.n441 10.6151
R1216 B.n441 B.n438 10.6151
R1217 B.n438 B.n437 10.6151
R1218 B.n437 B.n434 10.6151
R1219 B.n434 B.n433 10.6151
R1220 B.n433 B.n430 10.6151
R1221 B.n430 B.n429 10.6151
R1222 B.n429 B.n426 10.6151
R1223 B.n426 B.n425 10.6151
R1224 B.n425 B.n422 10.6151
R1225 B.n422 B.n421 10.6151
R1226 B.n421 B.n418 10.6151
R1227 B.n418 B.n417 10.6151
R1228 B.n417 B.n414 10.6151
R1229 B.n414 B.n350 10.6151
R1230 B.n635 B.n350 10.6151
R1231 B.n641 B.n346 10.6151
R1232 B.n642 B.n641 10.6151
R1233 B.n643 B.n642 10.6151
R1234 B.n643 B.n338 10.6151
R1235 B.n653 B.n338 10.6151
R1236 B.n654 B.n653 10.6151
R1237 B.n655 B.n654 10.6151
R1238 B.n655 B.n330 10.6151
R1239 B.n665 B.n330 10.6151
R1240 B.n666 B.n665 10.6151
R1241 B.n667 B.n666 10.6151
R1242 B.n667 B.n322 10.6151
R1243 B.n678 B.n322 10.6151
R1244 B.n679 B.n678 10.6151
R1245 B.n680 B.n679 10.6151
R1246 B.n680 B.n0 10.6151
R1247 B.n741 B.n1 10.6151
R1248 B.n741 B.n740 10.6151
R1249 B.n740 B.n739 10.6151
R1250 B.n739 B.n10 10.6151
R1251 B.n733 B.n10 10.6151
R1252 B.n733 B.n732 10.6151
R1253 B.n732 B.n731 10.6151
R1254 B.n731 B.n17 10.6151
R1255 B.n725 B.n17 10.6151
R1256 B.n725 B.n724 10.6151
R1257 B.n724 B.n723 10.6151
R1258 B.n723 B.n24 10.6151
R1259 B.n717 B.n24 10.6151
R1260 B.n717 B.n716 10.6151
R1261 B.n716 B.n715 10.6151
R1262 B.n715 B.n31 10.6151
R1263 B.n197 B.n196 9.36635
R1264 B.n219 B.n218 9.36635
R1265 B.n533 B.n410 9.36635
R1266 B.n510 B.n413 9.36635
R1267 B.n651 B.t5 3.2114
R1268 B.n721 B.t9 3.2114
R1269 B.n747 B.n0 2.81026
R1270 B.n747 B.n1 2.81026
R1271 B.t3 B.n320 2.1411
R1272 B.t0 B.n8 2.1411
R1273 B.n198 B.n197 1.24928
R1274 B.n218 B.n217 1.24928
R1275 B.n530 B.n410 1.24928
R1276 B.n513 B.n413 1.24928
R1277 B.n669 B.t2 1.0708
R1278 B.t1 B.n735 1.0708
R1279 VN.n0 VN.t0 638.467
R1280 VN.n1 VN.t1 638.467
R1281 VN.n0 VN.t3 638.418
R1282 VN.n1 VN.t2 638.418
R1283 VN VN.n1 87.7852
R1284 VN VN.n0 44.7132
R1285 VDD2.n2 VDD2.n0 99.1704
R1286 VDD2.n2 VDD2.n1 59.723
R1287 VDD2.n1 VDD2.t1 1.29631
R1288 VDD2.n1 VDD2.t2 1.29631
R1289 VDD2.n0 VDD2.t3 1.29631
R1290 VDD2.n0 VDD2.t0 1.29631
R1291 VDD2 VDD2.n2 0.0586897
C0 VTAIL VN 3.30287f
C1 VP VN 5.40142f
C2 VTAIL VDD2 8.47583f
C3 VP VDD2 0.270999f
C4 VN VDD1 0.147386f
C5 VP VTAIL 3.31697f
C6 VDD1 VDD2 0.557286f
C7 VTAIL VDD1 8.434629f
C8 VP VDD1 3.9666f
C9 VN VDD2 3.84323f
C10 VDD2 B 2.933042f
C11 VDD1 B 7.0432f
C12 VTAIL B 10.588008f
C13 VN B 8.578951f
C14 VP B 5.037591f
C15 VDD2.t3 B 0.344217f
C16 VDD2.t0 B 0.344217f
C17 VDD2.n0 B 3.85316f
C18 VDD2.t1 B 0.344217f
C19 VDD2.t2 B 0.344217f
C20 VDD2.n1 B 3.10482f
C21 VDD2.n2 B 3.88062f
C22 VN.t0 B 1.4489f
C23 VN.t3 B 1.44885f
C24 VN.n0 B 1.07007f
C25 VN.t1 B 1.4489f
C26 VN.t2 B 1.44885f
C27 VN.n1 B 2.17958f
C28 VTAIL.t0 B 2.1787f
C29 VTAIL.n0 B 0.277253f
C30 VTAIL.t6 B 2.1787f
C31 VTAIL.n1 B 0.29643f
C32 VTAIL.t7 B 2.1787f
C33 VTAIL.n2 B 1.22116f
C34 VTAIL.t2 B 2.17871f
C35 VTAIL.n3 B 1.22115f
C36 VTAIL.t3 B 2.17871f
C37 VTAIL.n4 B 0.296417f
C38 VTAIL.t5 B 2.17871f
C39 VTAIL.n5 B 0.296417f
C40 VTAIL.t4 B 2.17871f
C41 VTAIL.n6 B 1.22116f
C42 VTAIL.t1 B 2.1787f
C43 VTAIL.n7 B 1.19593f
C44 VDD1.t0 B 0.34407f
C45 VDD1.t3 B 0.34407f
C46 VDD1.n0 B 3.10382f
C47 VDD1.t1 B 0.34407f
C48 VDD1.t2 B 0.34407f
C49 VDD1.n1 B 3.88049f
C50 VP.n0 B 0.051024f
C51 VP.t3 B 1.48035f
C52 VP.t2 B 1.4804f
C53 VP.n1 B 2.20548f
C54 VP.n2 B 3.37343f
C55 VP.t0 B 1.46188f
C56 VP.n3 B 0.559116f
C57 VP.n4 B 0.011578f
C58 VP.t1 B 1.46188f
C59 VP.n5 B 0.559116f
C60 VP.n6 B 0.039542f
.ends

