* NGSPICE file created from diff_pair_sample_0064.ext - technology: sky130A

.subckt diff_pair_sample_0064 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t18 VN.t0 VDD2.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X1 VDD2.t4 VN.t1 VTAIL.t17 B.t22 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.5265 ps=3.48 w=1.35 l=2.44
X2 VTAIL.t16 VN.t2 VDD2.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X3 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0 ps=0 w=1.35 l=2.44
X4 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.5265 ps=3.48 w=1.35 l=2.44
X5 VDD2.t5 VN.t3 VTAIL.t15 B.t5 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X6 VTAIL.t14 VN.t4 VDD2.t2 B.t23 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X7 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0 ps=0 w=1.35 l=2.44
X8 VDD1.t8 VP.t1 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0.22275 ps=1.68 w=1.35 l=2.44
X9 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0 ps=0 w=1.35 l=2.44
X10 VTAIL.t2 VP.t2 VDD1.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X11 VTAIL.t13 VN.t5 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X12 VTAIL.t1 VP.t3 VDD1.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X13 VDD2.t7 VN.t6 VTAIL.t12 B.t3 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.5265 ps=3.48 w=1.35 l=2.44
X14 VDD2.t6 VN.t7 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0.22275 ps=1.68 w=1.35 l=2.44
X15 VDD1.t5 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X16 VTAIL.t7 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X17 VDD2.t0 VN.t8 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0.22275 ps=1.68 w=1.35 l=2.44
X18 VTAIL.t19 VP.t6 VDD1.t3 B.t23 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X19 VDD2.t9 VN.t9 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
X20 VDD1.t2 VP.t7 VTAIL.t8 B.t22 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.5265 ps=3.48 w=1.35 l=2.44
X21 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0 ps=0 w=1.35 l=2.44
X22 VDD1.t1 VP.t8 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=0.5265 pd=3.48 as=0.22275 ps=1.68 w=1.35 l=2.44
X23 VDD1.t0 VP.t9 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=0.22275 pd=1.68 as=0.22275 ps=1.68 w=1.35 l=2.44
R0 VN.n77 VN.n40 161.3
R1 VN.n76 VN.n75 161.3
R2 VN.n74 VN.n41 161.3
R3 VN.n73 VN.n72 161.3
R4 VN.n71 VN.n42 161.3
R5 VN.n69 VN.n68 161.3
R6 VN.n67 VN.n43 161.3
R7 VN.n66 VN.n65 161.3
R8 VN.n64 VN.n44 161.3
R9 VN.n63 VN.n62 161.3
R10 VN.n61 VN.n45 161.3
R11 VN.n60 VN.n59 161.3
R12 VN.n58 VN.n46 161.3
R13 VN.n57 VN.n56 161.3
R14 VN.n55 VN.n48 161.3
R15 VN.n54 VN.n53 161.3
R16 VN.n52 VN.n49 161.3
R17 VN.n37 VN.n0 161.3
R18 VN.n36 VN.n35 161.3
R19 VN.n34 VN.n1 161.3
R20 VN.n33 VN.n32 161.3
R21 VN.n31 VN.n2 161.3
R22 VN.n29 VN.n28 161.3
R23 VN.n27 VN.n3 161.3
R24 VN.n26 VN.n25 161.3
R25 VN.n24 VN.n4 161.3
R26 VN.n23 VN.n22 161.3
R27 VN.n21 VN.n5 161.3
R28 VN.n20 VN.n19 161.3
R29 VN.n17 VN.n6 161.3
R30 VN.n16 VN.n15 161.3
R31 VN.n14 VN.n7 161.3
R32 VN.n13 VN.n12 161.3
R33 VN.n11 VN.n8 161.3
R34 VN.n39 VN.n38 96.5656
R35 VN.n79 VN.n78 96.5656
R36 VN.n10 VN.n9 71.4859
R37 VN.n51 VN.n50 71.4859
R38 VN.n16 VN.n7 53.6055
R39 VN.n25 VN.n24 53.6055
R40 VN.n57 VN.n48 53.6055
R41 VN.n65 VN.n64 53.6055
R42 VN.n32 VN.n1 49.7204
R43 VN.n72 VN.n41 49.7204
R44 VN.n9 VN.t7 45.4455
R45 VN.n50 VN.t6 45.4455
R46 VN VN.n79 44.5019
R47 VN.n36 VN.n1 31.2664
R48 VN.n76 VN.n41 31.2664
R49 VN.n17 VN.n16 27.3813
R50 VN.n24 VN.n23 27.3813
R51 VN.n58 VN.n57 27.3813
R52 VN.n64 VN.n63 27.3813
R53 VN.n12 VN.n11 24.4675
R54 VN.n12 VN.n7 24.4675
R55 VN.n19 VN.n17 24.4675
R56 VN.n23 VN.n5 24.4675
R57 VN.n25 VN.n3 24.4675
R58 VN.n29 VN.n3 24.4675
R59 VN.n32 VN.n31 24.4675
R60 VN.n37 VN.n36 24.4675
R61 VN.n53 VN.n48 24.4675
R62 VN.n53 VN.n52 24.4675
R63 VN.n63 VN.n45 24.4675
R64 VN.n59 VN.n58 24.4675
R65 VN.n72 VN.n71 24.4675
R66 VN.n69 VN.n43 24.4675
R67 VN.n65 VN.n43 24.4675
R68 VN.n77 VN.n76 24.4675
R69 VN.n31 VN.n30 23.4888
R70 VN.n71 VN.n70 23.4888
R71 VN.n38 VN.n37 14.1914
R72 VN.n78 VN.n77 14.1914
R73 VN.n10 VN.t4 13.3345
R74 VN.n18 VN.t3 13.3345
R75 VN.n30 VN.t2 13.3345
R76 VN.n38 VN.t1 13.3345
R77 VN.n51 VN.t5 13.3345
R78 VN.n47 VN.t9 13.3345
R79 VN.n70 VN.t0 13.3345
R80 VN.n78 VN.t8 13.3345
R81 VN.n19 VN.n18 12.234
R82 VN.n18 VN.n5 12.234
R83 VN.n47 VN.n45 12.234
R84 VN.n59 VN.n47 12.234
R85 VN.n50 VN.n49 9.60581
R86 VN.n9 VN.n8 9.60581
R87 VN.n11 VN.n10 0.97918
R88 VN.n30 VN.n29 0.97918
R89 VN.n52 VN.n51 0.97918
R90 VN.n70 VN.n69 0.97918
R91 VN.n79 VN.n40 0.278367
R92 VN.n39 VN.n0 0.278367
R93 VN.n75 VN.n40 0.189894
R94 VN.n75 VN.n74 0.189894
R95 VN.n74 VN.n73 0.189894
R96 VN.n73 VN.n42 0.189894
R97 VN.n68 VN.n42 0.189894
R98 VN.n68 VN.n67 0.189894
R99 VN.n67 VN.n66 0.189894
R100 VN.n66 VN.n44 0.189894
R101 VN.n62 VN.n44 0.189894
R102 VN.n62 VN.n61 0.189894
R103 VN.n61 VN.n60 0.189894
R104 VN.n60 VN.n46 0.189894
R105 VN.n56 VN.n46 0.189894
R106 VN.n56 VN.n55 0.189894
R107 VN.n55 VN.n54 0.189894
R108 VN.n54 VN.n49 0.189894
R109 VN.n13 VN.n8 0.189894
R110 VN.n14 VN.n13 0.189894
R111 VN.n15 VN.n14 0.189894
R112 VN.n15 VN.n6 0.189894
R113 VN.n20 VN.n6 0.189894
R114 VN.n21 VN.n20 0.189894
R115 VN.n22 VN.n21 0.189894
R116 VN.n22 VN.n4 0.189894
R117 VN.n26 VN.n4 0.189894
R118 VN.n27 VN.n26 0.189894
R119 VN.n28 VN.n27 0.189894
R120 VN.n28 VN.n2 0.189894
R121 VN.n33 VN.n2 0.189894
R122 VN.n34 VN.n33 0.189894
R123 VN.n35 VN.n34 0.189894
R124 VN.n35 VN.n0 0.189894
R125 VN VN.n39 0.153454
R126 VDD2.n1 VDD2.t6 176.333
R127 VDD2.n4 VDD2.t0 173.945
R128 VDD2.n3 VDD2.n2 149.523
R129 VDD2 VDD2.n7 149.519
R130 VDD2.n1 VDD2.n0 147.786
R131 VDD2.n6 VDD2.n5 147.786
R132 VDD2.n4 VDD2.n3 36.2218
R133 VDD2.n7 VDD2.t1 14.6672
R134 VDD2.n7 VDD2.t7 14.6672
R135 VDD2.n5 VDD2.t3 14.6672
R136 VDD2.n5 VDD2.t9 14.6672
R137 VDD2.n2 VDD2.t8 14.6672
R138 VDD2.n2 VDD2.t4 14.6672
R139 VDD2.n0 VDD2.t2 14.6672
R140 VDD2.n0 VDD2.t5 14.6672
R141 VDD2.n6 VDD2.n4 2.38843
R142 VDD2 VDD2.n6 0.655672
R143 VDD2.n3 VDD2.n1 0.542137
R144 VTAIL.n17 VTAIL.t17 157.266
R145 VTAIL.n2 VTAIL.t3 157.266
R146 VTAIL.n16 VTAIL.t8 157.266
R147 VTAIL.n11 VTAIL.t12 157.266
R148 VTAIL.n19 VTAIL.n18 131.107
R149 VTAIL.n1 VTAIL.n0 131.107
R150 VTAIL.n4 VTAIL.n3 131.107
R151 VTAIL.n6 VTAIL.n5 131.107
R152 VTAIL.n15 VTAIL.n14 131.107
R153 VTAIL.n13 VTAIL.n12 131.107
R154 VTAIL.n10 VTAIL.n9 131.107
R155 VTAIL.n8 VTAIL.n7 131.107
R156 VTAIL.n8 VTAIL.n6 18.3065
R157 VTAIL.n17 VTAIL.n16 15.9186
R158 VTAIL.n18 VTAIL.t15 14.6672
R159 VTAIL.n18 VTAIL.t16 14.6672
R160 VTAIL.n0 VTAIL.t11 14.6672
R161 VTAIL.n0 VTAIL.t14 14.6672
R162 VTAIL.n3 VTAIL.t0 14.6672
R163 VTAIL.n3 VTAIL.t2 14.6672
R164 VTAIL.n5 VTAIL.t4 14.6672
R165 VTAIL.n5 VTAIL.t7 14.6672
R166 VTAIL.n14 VTAIL.t5 14.6672
R167 VTAIL.n14 VTAIL.t1 14.6672
R168 VTAIL.n12 VTAIL.t6 14.6672
R169 VTAIL.n12 VTAIL.t19 14.6672
R170 VTAIL.n9 VTAIL.t9 14.6672
R171 VTAIL.n9 VTAIL.t13 14.6672
R172 VTAIL.n7 VTAIL.t10 14.6672
R173 VTAIL.n7 VTAIL.t18 14.6672
R174 VTAIL.n10 VTAIL.n8 2.38843
R175 VTAIL.n11 VTAIL.n10 2.38843
R176 VTAIL.n15 VTAIL.n13 2.38843
R177 VTAIL.n16 VTAIL.n15 2.38843
R178 VTAIL.n6 VTAIL.n4 2.38843
R179 VTAIL.n4 VTAIL.n2 2.38843
R180 VTAIL.n19 VTAIL.n17 2.38843
R181 VTAIL VTAIL.n1 1.84964
R182 VTAIL.n13 VTAIL.n11 1.66429
R183 VTAIL.n2 VTAIL.n1 1.66429
R184 VTAIL VTAIL.n19 0.539293
R185 B.n619 B.n618 585
R186 B.n182 B.n119 585
R187 B.n181 B.n180 585
R188 B.n179 B.n178 585
R189 B.n177 B.n176 585
R190 B.n175 B.n174 585
R191 B.n173 B.n172 585
R192 B.n171 B.n170 585
R193 B.n169 B.n168 585
R194 B.n167 B.n166 585
R195 B.n165 B.n164 585
R196 B.n163 B.n162 585
R197 B.n161 B.n160 585
R198 B.n159 B.n158 585
R199 B.n157 B.n156 585
R200 B.n155 B.n154 585
R201 B.n153 B.n152 585
R202 B.n151 B.n150 585
R203 B.n149 B.n148 585
R204 B.n147 B.n146 585
R205 B.n145 B.n144 585
R206 B.n143 B.n142 585
R207 B.n141 B.n140 585
R208 B.n139 B.n138 585
R209 B.n137 B.n136 585
R210 B.n135 B.n134 585
R211 B.n133 B.n132 585
R212 B.n131 B.n130 585
R213 B.n129 B.n128 585
R214 B.n127 B.n126 585
R215 B.n617 B.n104 585
R216 B.n622 B.n104 585
R217 B.n616 B.n103 585
R218 B.n623 B.n103 585
R219 B.n615 B.n614 585
R220 B.n614 B.n99 585
R221 B.n613 B.n98 585
R222 B.n629 B.n98 585
R223 B.n612 B.n97 585
R224 B.n630 B.n97 585
R225 B.n611 B.n96 585
R226 B.n631 B.n96 585
R227 B.n610 B.n609 585
R228 B.n609 B.n92 585
R229 B.n608 B.n91 585
R230 B.n637 B.n91 585
R231 B.n607 B.n90 585
R232 B.n638 B.n90 585
R233 B.n606 B.n89 585
R234 B.n639 B.n89 585
R235 B.n605 B.n604 585
R236 B.n604 B.n85 585
R237 B.n603 B.n84 585
R238 B.n645 B.n84 585
R239 B.n602 B.n83 585
R240 B.n646 B.n83 585
R241 B.n601 B.n82 585
R242 B.n647 B.n82 585
R243 B.n600 B.n599 585
R244 B.n599 B.n78 585
R245 B.n598 B.n77 585
R246 B.n653 B.n77 585
R247 B.n597 B.n76 585
R248 B.n654 B.n76 585
R249 B.n596 B.n75 585
R250 B.n655 B.n75 585
R251 B.n595 B.n594 585
R252 B.n594 B.n74 585
R253 B.n593 B.n70 585
R254 B.n661 B.n70 585
R255 B.n592 B.n69 585
R256 B.n662 B.n69 585
R257 B.n591 B.n68 585
R258 B.n663 B.n68 585
R259 B.n590 B.n589 585
R260 B.n589 B.n64 585
R261 B.n588 B.n63 585
R262 B.n669 B.n63 585
R263 B.n587 B.n62 585
R264 B.n670 B.n62 585
R265 B.n586 B.n61 585
R266 B.n671 B.n61 585
R267 B.n585 B.n584 585
R268 B.n584 B.n60 585
R269 B.n583 B.n56 585
R270 B.n677 B.n56 585
R271 B.n582 B.n55 585
R272 B.n678 B.n55 585
R273 B.n581 B.n54 585
R274 B.n679 B.n54 585
R275 B.n580 B.n579 585
R276 B.n579 B.n50 585
R277 B.n578 B.n49 585
R278 B.n685 B.n49 585
R279 B.n577 B.n48 585
R280 B.n686 B.n48 585
R281 B.n576 B.n47 585
R282 B.n687 B.n47 585
R283 B.n575 B.n574 585
R284 B.n574 B.n43 585
R285 B.n573 B.n42 585
R286 B.n693 B.n42 585
R287 B.n572 B.n41 585
R288 B.n694 B.n41 585
R289 B.n571 B.n40 585
R290 B.n695 B.n40 585
R291 B.n570 B.n569 585
R292 B.n569 B.n36 585
R293 B.n568 B.n35 585
R294 B.n701 B.n35 585
R295 B.n567 B.n34 585
R296 B.n702 B.n34 585
R297 B.n566 B.n33 585
R298 B.n703 B.n33 585
R299 B.n565 B.n564 585
R300 B.n564 B.n29 585
R301 B.n563 B.n28 585
R302 B.n709 B.n28 585
R303 B.n562 B.n27 585
R304 B.n710 B.n27 585
R305 B.n561 B.n26 585
R306 B.n711 B.n26 585
R307 B.n560 B.n559 585
R308 B.n559 B.n22 585
R309 B.n558 B.n21 585
R310 B.n717 B.n21 585
R311 B.n557 B.n20 585
R312 B.n718 B.n20 585
R313 B.n556 B.n19 585
R314 B.n719 B.n19 585
R315 B.n555 B.n554 585
R316 B.n554 B.n15 585
R317 B.n553 B.n14 585
R318 B.n725 B.n14 585
R319 B.n552 B.n13 585
R320 B.n726 B.n13 585
R321 B.n551 B.n12 585
R322 B.n727 B.n12 585
R323 B.n550 B.n549 585
R324 B.n549 B.n8 585
R325 B.n548 B.n7 585
R326 B.n733 B.n7 585
R327 B.n547 B.n6 585
R328 B.n734 B.n6 585
R329 B.n546 B.n5 585
R330 B.n735 B.n5 585
R331 B.n545 B.n544 585
R332 B.n544 B.n4 585
R333 B.n543 B.n183 585
R334 B.n543 B.n542 585
R335 B.n533 B.n184 585
R336 B.n185 B.n184 585
R337 B.n535 B.n534 585
R338 B.n536 B.n535 585
R339 B.n532 B.n190 585
R340 B.n190 B.n189 585
R341 B.n531 B.n530 585
R342 B.n530 B.n529 585
R343 B.n192 B.n191 585
R344 B.n193 B.n192 585
R345 B.n522 B.n521 585
R346 B.n523 B.n522 585
R347 B.n520 B.n198 585
R348 B.n198 B.n197 585
R349 B.n519 B.n518 585
R350 B.n518 B.n517 585
R351 B.n200 B.n199 585
R352 B.n201 B.n200 585
R353 B.n510 B.n509 585
R354 B.n511 B.n510 585
R355 B.n508 B.n206 585
R356 B.n206 B.n205 585
R357 B.n507 B.n506 585
R358 B.n506 B.n505 585
R359 B.n208 B.n207 585
R360 B.n209 B.n208 585
R361 B.n498 B.n497 585
R362 B.n499 B.n498 585
R363 B.n496 B.n214 585
R364 B.n214 B.n213 585
R365 B.n495 B.n494 585
R366 B.n494 B.n493 585
R367 B.n216 B.n215 585
R368 B.n217 B.n216 585
R369 B.n486 B.n485 585
R370 B.n487 B.n486 585
R371 B.n484 B.n222 585
R372 B.n222 B.n221 585
R373 B.n483 B.n482 585
R374 B.n482 B.n481 585
R375 B.n224 B.n223 585
R376 B.n225 B.n224 585
R377 B.n474 B.n473 585
R378 B.n475 B.n474 585
R379 B.n472 B.n230 585
R380 B.n230 B.n229 585
R381 B.n471 B.n470 585
R382 B.n470 B.n469 585
R383 B.n232 B.n231 585
R384 B.n233 B.n232 585
R385 B.n462 B.n461 585
R386 B.n463 B.n462 585
R387 B.n460 B.n238 585
R388 B.n238 B.n237 585
R389 B.n459 B.n458 585
R390 B.n458 B.n457 585
R391 B.n240 B.n239 585
R392 B.n450 B.n240 585
R393 B.n449 B.n448 585
R394 B.n451 B.n449 585
R395 B.n447 B.n245 585
R396 B.n245 B.n244 585
R397 B.n446 B.n445 585
R398 B.n445 B.n444 585
R399 B.n247 B.n246 585
R400 B.n248 B.n247 585
R401 B.n437 B.n436 585
R402 B.n438 B.n437 585
R403 B.n435 B.n253 585
R404 B.n253 B.n252 585
R405 B.n434 B.n433 585
R406 B.n433 B.n432 585
R407 B.n255 B.n254 585
R408 B.n425 B.n255 585
R409 B.n424 B.n423 585
R410 B.n426 B.n424 585
R411 B.n422 B.n260 585
R412 B.n260 B.n259 585
R413 B.n421 B.n420 585
R414 B.n420 B.n419 585
R415 B.n262 B.n261 585
R416 B.n263 B.n262 585
R417 B.n412 B.n411 585
R418 B.n413 B.n412 585
R419 B.n410 B.n268 585
R420 B.n268 B.n267 585
R421 B.n409 B.n408 585
R422 B.n408 B.n407 585
R423 B.n270 B.n269 585
R424 B.n271 B.n270 585
R425 B.n400 B.n399 585
R426 B.n401 B.n400 585
R427 B.n398 B.n276 585
R428 B.n276 B.n275 585
R429 B.n397 B.n396 585
R430 B.n396 B.n395 585
R431 B.n278 B.n277 585
R432 B.n279 B.n278 585
R433 B.n388 B.n387 585
R434 B.n389 B.n388 585
R435 B.n386 B.n284 585
R436 B.n284 B.n283 585
R437 B.n385 B.n384 585
R438 B.n384 B.n383 585
R439 B.n286 B.n285 585
R440 B.n287 B.n286 585
R441 B.n376 B.n375 585
R442 B.n377 B.n376 585
R443 B.n374 B.n292 585
R444 B.n292 B.n291 585
R445 B.n369 B.n368 585
R446 B.n367 B.n309 585
R447 B.n366 B.n308 585
R448 B.n371 B.n308 585
R449 B.n365 B.n364 585
R450 B.n363 B.n362 585
R451 B.n361 B.n360 585
R452 B.n359 B.n358 585
R453 B.n357 B.n356 585
R454 B.n355 B.n354 585
R455 B.n353 B.n352 585
R456 B.n350 B.n349 585
R457 B.n348 B.n347 585
R458 B.n346 B.n345 585
R459 B.n344 B.n343 585
R460 B.n342 B.n341 585
R461 B.n340 B.n339 585
R462 B.n338 B.n337 585
R463 B.n336 B.n335 585
R464 B.n334 B.n333 585
R465 B.n332 B.n331 585
R466 B.n329 B.n328 585
R467 B.n327 B.n326 585
R468 B.n325 B.n324 585
R469 B.n323 B.n322 585
R470 B.n321 B.n320 585
R471 B.n319 B.n318 585
R472 B.n317 B.n316 585
R473 B.n315 B.n314 585
R474 B.n294 B.n293 585
R475 B.n373 B.n372 585
R476 B.n372 B.n371 585
R477 B.n290 B.n289 585
R478 B.n291 B.n290 585
R479 B.n379 B.n378 585
R480 B.n378 B.n377 585
R481 B.n380 B.n288 585
R482 B.n288 B.n287 585
R483 B.n382 B.n381 585
R484 B.n383 B.n382 585
R485 B.n282 B.n281 585
R486 B.n283 B.n282 585
R487 B.n391 B.n390 585
R488 B.n390 B.n389 585
R489 B.n392 B.n280 585
R490 B.n280 B.n279 585
R491 B.n394 B.n393 585
R492 B.n395 B.n394 585
R493 B.n274 B.n273 585
R494 B.n275 B.n274 585
R495 B.n403 B.n402 585
R496 B.n402 B.n401 585
R497 B.n404 B.n272 585
R498 B.n272 B.n271 585
R499 B.n406 B.n405 585
R500 B.n407 B.n406 585
R501 B.n266 B.n265 585
R502 B.n267 B.n266 585
R503 B.n415 B.n414 585
R504 B.n414 B.n413 585
R505 B.n416 B.n264 585
R506 B.n264 B.n263 585
R507 B.n418 B.n417 585
R508 B.n419 B.n418 585
R509 B.n258 B.n257 585
R510 B.n259 B.n258 585
R511 B.n428 B.n427 585
R512 B.n427 B.n426 585
R513 B.n429 B.n256 585
R514 B.n425 B.n256 585
R515 B.n431 B.n430 585
R516 B.n432 B.n431 585
R517 B.n251 B.n250 585
R518 B.n252 B.n251 585
R519 B.n440 B.n439 585
R520 B.n439 B.n438 585
R521 B.n441 B.n249 585
R522 B.n249 B.n248 585
R523 B.n443 B.n442 585
R524 B.n444 B.n443 585
R525 B.n243 B.n242 585
R526 B.n244 B.n243 585
R527 B.n453 B.n452 585
R528 B.n452 B.n451 585
R529 B.n454 B.n241 585
R530 B.n450 B.n241 585
R531 B.n456 B.n455 585
R532 B.n457 B.n456 585
R533 B.n236 B.n235 585
R534 B.n237 B.n236 585
R535 B.n465 B.n464 585
R536 B.n464 B.n463 585
R537 B.n466 B.n234 585
R538 B.n234 B.n233 585
R539 B.n468 B.n467 585
R540 B.n469 B.n468 585
R541 B.n228 B.n227 585
R542 B.n229 B.n228 585
R543 B.n477 B.n476 585
R544 B.n476 B.n475 585
R545 B.n478 B.n226 585
R546 B.n226 B.n225 585
R547 B.n480 B.n479 585
R548 B.n481 B.n480 585
R549 B.n220 B.n219 585
R550 B.n221 B.n220 585
R551 B.n489 B.n488 585
R552 B.n488 B.n487 585
R553 B.n490 B.n218 585
R554 B.n218 B.n217 585
R555 B.n492 B.n491 585
R556 B.n493 B.n492 585
R557 B.n212 B.n211 585
R558 B.n213 B.n212 585
R559 B.n501 B.n500 585
R560 B.n500 B.n499 585
R561 B.n502 B.n210 585
R562 B.n210 B.n209 585
R563 B.n504 B.n503 585
R564 B.n505 B.n504 585
R565 B.n204 B.n203 585
R566 B.n205 B.n204 585
R567 B.n513 B.n512 585
R568 B.n512 B.n511 585
R569 B.n514 B.n202 585
R570 B.n202 B.n201 585
R571 B.n516 B.n515 585
R572 B.n517 B.n516 585
R573 B.n196 B.n195 585
R574 B.n197 B.n196 585
R575 B.n525 B.n524 585
R576 B.n524 B.n523 585
R577 B.n526 B.n194 585
R578 B.n194 B.n193 585
R579 B.n528 B.n527 585
R580 B.n529 B.n528 585
R581 B.n188 B.n187 585
R582 B.n189 B.n188 585
R583 B.n538 B.n537 585
R584 B.n537 B.n536 585
R585 B.n539 B.n186 585
R586 B.n186 B.n185 585
R587 B.n541 B.n540 585
R588 B.n542 B.n541 585
R589 B.n2 B.n0 585
R590 B.n4 B.n2 585
R591 B.n3 B.n1 585
R592 B.n734 B.n3 585
R593 B.n732 B.n731 585
R594 B.n733 B.n732 585
R595 B.n730 B.n9 585
R596 B.n9 B.n8 585
R597 B.n729 B.n728 585
R598 B.n728 B.n727 585
R599 B.n11 B.n10 585
R600 B.n726 B.n11 585
R601 B.n724 B.n723 585
R602 B.n725 B.n724 585
R603 B.n722 B.n16 585
R604 B.n16 B.n15 585
R605 B.n721 B.n720 585
R606 B.n720 B.n719 585
R607 B.n18 B.n17 585
R608 B.n718 B.n18 585
R609 B.n716 B.n715 585
R610 B.n717 B.n716 585
R611 B.n714 B.n23 585
R612 B.n23 B.n22 585
R613 B.n713 B.n712 585
R614 B.n712 B.n711 585
R615 B.n25 B.n24 585
R616 B.n710 B.n25 585
R617 B.n708 B.n707 585
R618 B.n709 B.n708 585
R619 B.n706 B.n30 585
R620 B.n30 B.n29 585
R621 B.n705 B.n704 585
R622 B.n704 B.n703 585
R623 B.n32 B.n31 585
R624 B.n702 B.n32 585
R625 B.n700 B.n699 585
R626 B.n701 B.n700 585
R627 B.n698 B.n37 585
R628 B.n37 B.n36 585
R629 B.n697 B.n696 585
R630 B.n696 B.n695 585
R631 B.n39 B.n38 585
R632 B.n694 B.n39 585
R633 B.n692 B.n691 585
R634 B.n693 B.n692 585
R635 B.n690 B.n44 585
R636 B.n44 B.n43 585
R637 B.n689 B.n688 585
R638 B.n688 B.n687 585
R639 B.n46 B.n45 585
R640 B.n686 B.n46 585
R641 B.n684 B.n683 585
R642 B.n685 B.n684 585
R643 B.n682 B.n51 585
R644 B.n51 B.n50 585
R645 B.n681 B.n680 585
R646 B.n680 B.n679 585
R647 B.n53 B.n52 585
R648 B.n678 B.n53 585
R649 B.n676 B.n675 585
R650 B.n677 B.n676 585
R651 B.n674 B.n57 585
R652 B.n60 B.n57 585
R653 B.n673 B.n672 585
R654 B.n672 B.n671 585
R655 B.n59 B.n58 585
R656 B.n670 B.n59 585
R657 B.n668 B.n667 585
R658 B.n669 B.n668 585
R659 B.n666 B.n65 585
R660 B.n65 B.n64 585
R661 B.n665 B.n664 585
R662 B.n664 B.n663 585
R663 B.n67 B.n66 585
R664 B.n662 B.n67 585
R665 B.n660 B.n659 585
R666 B.n661 B.n660 585
R667 B.n658 B.n71 585
R668 B.n74 B.n71 585
R669 B.n657 B.n656 585
R670 B.n656 B.n655 585
R671 B.n73 B.n72 585
R672 B.n654 B.n73 585
R673 B.n652 B.n651 585
R674 B.n653 B.n652 585
R675 B.n650 B.n79 585
R676 B.n79 B.n78 585
R677 B.n649 B.n648 585
R678 B.n648 B.n647 585
R679 B.n81 B.n80 585
R680 B.n646 B.n81 585
R681 B.n644 B.n643 585
R682 B.n645 B.n644 585
R683 B.n642 B.n86 585
R684 B.n86 B.n85 585
R685 B.n641 B.n640 585
R686 B.n640 B.n639 585
R687 B.n88 B.n87 585
R688 B.n638 B.n88 585
R689 B.n636 B.n635 585
R690 B.n637 B.n636 585
R691 B.n634 B.n93 585
R692 B.n93 B.n92 585
R693 B.n633 B.n632 585
R694 B.n632 B.n631 585
R695 B.n95 B.n94 585
R696 B.n630 B.n95 585
R697 B.n628 B.n627 585
R698 B.n629 B.n628 585
R699 B.n626 B.n100 585
R700 B.n100 B.n99 585
R701 B.n625 B.n624 585
R702 B.n624 B.n623 585
R703 B.n102 B.n101 585
R704 B.n622 B.n102 585
R705 B.n737 B.n736 585
R706 B.n736 B.n735 585
R707 B.n369 B.n290 511.721
R708 B.n126 B.n102 511.721
R709 B.n372 B.n292 511.721
R710 B.n619 B.n104 511.721
R711 B.n621 B.n620 256.663
R712 B.n621 B.n118 256.663
R713 B.n621 B.n117 256.663
R714 B.n621 B.n116 256.663
R715 B.n621 B.n115 256.663
R716 B.n621 B.n114 256.663
R717 B.n621 B.n113 256.663
R718 B.n621 B.n112 256.663
R719 B.n621 B.n111 256.663
R720 B.n621 B.n110 256.663
R721 B.n621 B.n109 256.663
R722 B.n621 B.n108 256.663
R723 B.n621 B.n107 256.663
R724 B.n621 B.n106 256.663
R725 B.n621 B.n105 256.663
R726 B.n371 B.n370 256.663
R727 B.n371 B.n295 256.663
R728 B.n371 B.n296 256.663
R729 B.n371 B.n297 256.663
R730 B.n371 B.n298 256.663
R731 B.n371 B.n299 256.663
R732 B.n371 B.n300 256.663
R733 B.n371 B.n301 256.663
R734 B.n371 B.n302 256.663
R735 B.n371 B.n303 256.663
R736 B.n371 B.n304 256.663
R737 B.n371 B.n305 256.663
R738 B.n371 B.n306 256.663
R739 B.n371 B.n307 256.663
R740 B.n312 B.t12 208.524
R741 B.n310 B.t19 208.524
R742 B.n123 B.t16 208.524
R743 B.n120 B.t8 208.524
R744 B.n312 B.t15 204.869
R745 B.n310 B.t21 204.869
R746 B.n123 B.t17 204.869
R747 B.n120 B.t10 204.869
R748 B.n371 B.n291 204.226
R749 B.n622 B.n621 204.226
R750 B.n378 B.n290 163.367
R751 B.n378 B.n288 163.367
R752 B.n382 B.n288 163.367
R753 B.n382 B.n282 163.367
R754 B.n390 B.n282 163.367
R755 B.n390 B.n280 163.367
R756 B.n394 B.n280 163.367
R757 B.n394 B.n274 163.367
R758 B.n402 B.n274 163.367
R759 B.n402 B.n272 163.367
R760 B.n406 B.n272 163.367
R761 B.n406 B.n266 163.367
R762 B.n414 B.n266 163.367
R763 B.n414 B.n264 163.367
R764 B.n418 B.n264 163.367
R765 B.n418 B.n258 163.367
R766 B.n427 B.n258 163.367
R767 B.n427 B.n256 163.367
R768 B.n431 B.n256 163.367
R769 B.n431 B.n251 163.367
R770 B.n439 B.n251 163.367
R771 B.n439 B.n249 163.367
R772 B.n443 B.n249 163.367
R773 B.n443 B.n243 163.367
R774 B.n452 B.n243 163.367
R775 B.n452 B.n241 163.367
R776 B.n456 B.n241 163.367
R777 B.n456 B.n236 163.367
R778 B.n464 B.n236 163.367
R779 B.n464 B.n234 163.367
R780 B.n468 B.n234 163.367
R781 B.n468 B.n228 163.367
R782 B.n476 B.n228 163.367
R783 B.n476 B.n226 163.367
R784 B.n480 B.n226 163.367
R785 B.n480 B.n220 163.367
R786 B.n488 B.n220 163.367
R787 B.n488 B.n218 163.367
R788 B.n492 B.n218 163.367
R789 B.n492 B.n212 163.367
R790 B.n500 B.n212 163.367
R791 B.n500 B.n210 163.367
R792 B.n504 B.n210 163.367
R793 B.n504 B.n204 163.367
R794 B.n512 B.n204 163.367
R795 B.n512 B.n202 163.367
R796 B.n516 B.n202 163.367
R797 B.n516 B.n196 163.367
R798 B.n524 B.n196 163.367
R799 B.n524 B.n194 163.367
R800 B.n528 B.n194 163.367
R801 B.n528 B.n188 163.367
R802 B.n537 B.n188 163.367
R803 B.n537 B.n186 163.367
R804 B.n541 B.n186 163.367
R805 B.n541 B.n2 163.367
R806 B.n736 B.n2 163.367
R807 B.n736 B.n3 163.367
R808 B.n732 B.n3 163.367
R809 B.n732 B.n9 163.367
R810 B.n728 B.n9 163.367
R811 B.n728 B.n11 163.367
R812 B.n724 B.n11 163.367
R813 B.n724 B.n16 163.367
R814 B.n720 B.n16 163.367
R815 B.n720 B.n18 163.367
R816 B.n716 B.n18 163.367
R817 B.n716 B.n23 163.367
R818 B.n712 B.n23 163.367
R819 B.n712 B.n25 163.367
R820 B.n708 B.n25 163.367
R821 B.n708 B.n30 163.367
R822 B.n704 B.n30 163.367
R823 B.n704 B.n32 163.367
R824 B.n700 B.n32 163.367
R825 B.n700 B.n37 163.367
R826 B.n696 B.n37 163.367
R827 B.n696 B.n39 163.367
R828 B.n692 B.n39 163.367
R829 B.n692 B.n44 163.367
R830 B.n688 B.n44 163.367
R831 B.n688 B.n46 163.367
R832 B.n684 B.n46 163.367
R833 B.n684 B.n51 163.367
R834 B.n680 B.n51 163.367
R835 B.n680 B.n53 163.367
R836 B.n676 B.n53 163.367
R837 B.n676 B.n57 163.367
R838 B.n672 B.n57 163.367
R839 B.n672 B.n59 163.367
R840 B.n668 B.n59 163.367
R841 B.n668 B.n65 163.367
R842 B.n664 B.n65 163.367
R843 B.n664 B.n67 163.367
R844 B.n660 B.n67 163.367
R845 B.n660 B.n71 163.367
R846 B.n656 B.n71 163.367
R847 B.n656 B.n73 163.367
R848 B.n652 B.n73 163.367
R849 B.n652 B.n79 163.367
R850 B.n648 B.n79 163.367
R851 B.n648 B.n81 163.367
R852 B.n644 B.n81 163.367
R853 B.n644 B.n86 163.367
R854 B.n640 B.n86 163.367
R855 B.n640 B.n88 163.367
R856 B.n636 B.n88 163.367
R857 B.n636 B.n93 163.367
R858 B.n632 B.n93 163.367
R859 B.n632 B.n95 163.367
R860 B.n628 B.n95 163.367
R861 B.n628 B.n100 163.367
R862 B.n624 B.n100 163.367
R863 B.n624 B.n102 163.367
R864 B.n309 B.n308 163.367
R865 B.n364 B.n308 163.367
R866 B.n362 B.n361 163.367
R867 B.n358 B.n357 163.367
R868 B.n354 B.n353 163.367
R869 B.n349 B.n348 163.367
R870 B.n345 B.n344 163.367
R871 B.n341 B.n340 163.367
R872 B.n337 B.n336 163.367
R873 B.n333 B.n332 163.367
R874 B.n328 B.n327 163.367
R875 B.n324 B.n323 163.367
R876 B.n320 B.n319 163.367
R877 B.n316 B.n315 163.367
R878 B.n372 B.n294 163.367
R879 B.n376 B.n292 163.367
R880 B.n376 B.n286 163.367
R881 B.n384 B.n286 163.367
R882 B.n384 B.n284 163.367
R883 B.n388 B.n284 163.367
R884 B.n388 B.n278 163.367
R885 B.n396 B.n278 163.367
R886 B.n396 B.n276 163.367
R887 B.n400 B.n276 163.367
R888 B.n400 B.n270 163.367
R889 B.n408 B.n270 163.367
R890 B.n408 B.n268 163.367
R891 B.n412 B.n268 163.367
R892 B.n412 B.n262 163.367
R893 B.n420 B.n262 163.367
R894 B.n420 B.n260 163.367
R895 B.n424 B.n260 163.367
R896 B.n424 B.n255 163.367
R897 B.n433 B.n255 163.367
R898 B.n433 B.n253 163.367
R899 B.n437 B.n253 163.367
R900 B.n437 B.n247 163.367
R901 B.n445 B.n247 163.367
R902 B.n445 B.n245 163.367
R903 B.n449 B.n245 163.367
R904 B.n449 B.n240 163.367
R905 B.n458 B.n240 163.367
R906 B.n458 B.n238 163.367
R907 B.n462 B.n238 163.367
R908 B.n462 B.n232 163.367
R909 B.n470 B.n232 163.367
R910 B.n470 B.n230 163.367
R911 B.n474 B.n230 163.367
R912 B.n474 B.n224 163.367
R913 B.n482 B.n224 163.367
R914 B.n482 B.n222 163.367
R915 B.n486 B.n222 163.367
R916 B.n486 B.n216 163.367
R917 B.n494 B.n216 163.367
R918 B.n494 B.n214 163.367
R919 B.n498 B.n214 163.367
R920 B.n498 B.n208 163.367
R921 B.n506 B.n208 163.367
R922 B.n506 B.n206 163.367
R923 B.n510 B.n206 163.367
R924 B.n510 B.n200 163.367
R925 B.n518 B.n200 163.367
R926 B.n518 B.n198 163.367
R927 B.n522 B.n198 163.367
R928 B.n522 B.n192 163.367
R929 B.n530 B.n192 163.367
R930 B.n530 B.n190 163.367
R931 B.n535 B.n190 163.367
R932 B.n535 B.n184 163.367
R933 B.n543 B.n184 163.367
R934 B.n544 B.n543 163.367
R935 B.n544 B.n5 163.367
R936 B.n6 B.n5 163.367
R937 B.n7 B.n6 163.367
R938 B.n549 B.n7 163.367
R939 B.n549 B.n12 163.367
R940 B.n13 B.n12 163.367
R941 B.n14 B.n13 163.367
R942 B.n554 B.n14 163.367
R943 B.n554 B.n19 163.367
R944 B.n20 B.n19 163.367
R945 B.n21 B.n20 163.367
R946 B.n559 B.n21 163.367
R947 B.n559 B.n26 163.367
R948 B.n27 B.n26 163.367
R949 B.n28 B.n27 163.367
R950 B.n564 B.n28 163.367
R951 B.n564 B.n33 163.367
R952 B.n34 B.n33 163.367
R953 B.n35 B.n34 163.367
R954 B.n569 B.n35 163.367
R955 B.n569 B.n40 163.367
R956 B.n41 B.n40 163.367
R957 B.n42 B.n41 163.367
R958 B.n574 B.n42 163.367
R959 B.n574 B.n47 163.367
R960 B.n48 B.n47 163.367
R961 B.n49 B.n48 163.367
R962 B.n579 B.n49 163.367
R963 B.n579 B.n54 163.367
R964 B.n55 B.n54 163.367
R965 B.n56 B.n55 163.367
R966 B.n584 B.n56 163.367
R967 B.n584 B.n61 163.367
R968 B.n62 B.n61 163.367
R969 B.n63 B.n62 163.367
R970 B.n589 B.n63 163.367
R971 B.n589 B.n68 163.367
R972 B.n69 B.n68 163.367
R973 B.n70 B.n69 163.367
R974 B.n594 B.n70 163.367
R975 B.n594 B.n75 163.367
R976 B.n76 B.n75 163.367
R977 B.n77 B.n76 163.367
R978 B.n599 B.n77 163.367
R979 B.n599 B.n82 163.367
R980 B.n83 B.n82 163.367
R981 B.n84 B.n83 163.367
R982 B.n604 B.n84 163.367
R983 B.n604 B.n89 163.367
R984 B.n90 B.n89 163.367
R985 B.n91 B.n90 163.367
R986 B.n609 B.n91 163.367
R987 B.n609 B.n96 163.367
R988 B.n97 B.n96 163.367
R989 B.n98 B.n97 163.367
R990 B.n614 B.n98 163.367
R991 B.n614 B.n103 163.367
R992 B.n104 B.n103 163.367
R993 B.n130 B.n129 163.367
R994 B.n134 B.n133 163.367
R995 B.n138 B.n137 163.367
R996 B.n142 B.n141 163.367
R997 B.n146 B.n145 163.367
R998 B.n150 B.n149 163.367
R999 B.n154 B.n153 163.367
R1000 B.n158 B.n157 163.367
R1001 B.n162 B.n161 163.367
R1002 B.n166 B.n165 163.367
R1003 B.n170 B.n169 163.367
R1004 B.n174 B.n173 163.367
R1005 B.n178 B.n177 163.367
R1006 B.n180 B.n119 163.367
R1007 B.n313 B.t14 151.149
R1008 B.n311 B.t20 151.149
R1009 B.n124 B.t18 151.149
R1010 B.n121 B.t11 151.149
R1011 B.n377 B.n291 112.906
R1012 B.n377 B.n287 112.906
R1013 B.n383 B.n287 112.906
R1014 B.n383 B.n283 112.906
R1015 B.n389 B.n283 112.906
R1016 B.n389 B.n279 112.906
R1017 B.n395 B.n279 112.906
R1018 B.n401 B.n275 112.906
R1019 B.n401 B.n271 112.906
R1020 B.n407 B.n271 112.906
R1021 B.n407 B.n267 112.906
R1022 B.n413 B.n267 112.906
R1023 B.n413 B.n263 112.906
R1024 B.n419 B.n263 112.906
R1025 B.n419 B.n259 112.906
R1026 B.n426 B.n259 112.906
R1027 B.n426 B.n425 112.906
R1028 B.n432 B.n252 112.906
R1029 B.n438 B.n252 112.906
R1030 B.n438 B.n248 112.906
R1031 B.n444 B.n248 112.906
R1032 B.n444 B.n244 112.906
R1033 B.n451 B.n244 112.906
R1034 B.n451 B.n450 112.906
R1035 B.n457 B.n237 112.906
R1036 B.n463 B.n237 112.906
R1037 B.n463 B.n233 112.906
R1038 B.n469 B.n233 112.906
R1039 B.n469 B.n229 112.906
R1040 B.n475 B.n229 112.906
R1041 B.n475 B.n225 112.906
R1042 B.n481 B.n225 112.906
R1043 B.n487 B.n221 112.906
R1044 B.n487 B.n217 112.906
R1045 B.n493 B.n217 112.906
R1046 B.n493 B.n213 112.906
R1047 B.n499 B.n213 112.906
R1048 B.n499 B.n209 112.906
R1049 B.n505 B.n209 112.906
R1050 B.n511 B.n205 112.906
R1051 B.n511 B.n201 112.906
R1052 B.n517 B.n201 112.906
R1053 B.n517 B.n197 112.906
R1054 B.n523 B.n197 112.906
R1055 B.n523 B.n193 112.906
R1056 B.n529 B.n193 112.906
R1057 B.n536 B.n189 112.906
R1058 B.n536 B.n185 112.906
R1059 B.n542 B.n185 112.906
R1060 B.n542 B.n4 112.906
R1061 B.n735 B.n4 112.906
R1062 B.n735 B.n734 112.906
R1063 B.n734 B.n733 112.906
R1064 B.n733 B.n8 112.906
R1065 B.n727 B.n8 112.906
R1066 B.n727 B.n726 112.906
R1067 B.n725 B.n15 112.906
R1068 B.n719 B.n15 112.906
R1069 B.n719 B.n718 112.906
R1070 B.n718 B.n717 112.906
R1071 B.n717 B.n22 112.906
R1072 B.n711 B.n22 112.906
R1073 B.n711 B.n710 112.906
R1074 B.n709 B.n29 112.906
R1075 B.n703 B.n29 112.906
R1076 B.n703 B.n702 112.906
R1077 B.n702 B.n701 112.906
R1078 B.n701 B.n36 112.906
R1079 B.n695 B.n36 112.906
R1080 B.n695 B.n694 112.906
R1081 B.n693 B.n43 112.906
R1082 B.n687 B.n43 112.906
R1083 B.n687 B.n686 112.906
R1084 B.n686 B.n685 112.906
R1085 B.n685 B.n50 112.906
R1086 B.n679 B.n50 112.906
R1087 B.n679 B.n678 112.906
R1088 B.n678 B.n677 112.906
R1089 B.n671 B.n60 112.906
R1090 B.n671 B.n670 112.906
R1091 B.n670 B.n669 112.906
R1092 B.n669 B.n64 112.906
R1093 B.n663 B.n64 112.906
R1094 B.n663 B.n662 112.906
R1095 B.n662 B.n661 112.906
R1096 B.n655 B.n74 112.906
R1097 B.n655 B.n654 112.906
R1098 B.n654 B.n653 112.906
R1099 B.n653 B.n78 112.906
R1100 B.n647 B.n78 112.906
R1101 B.n647 B.n646 112.906
R1102 B.n646 B.n645 112.906
R1103 B.n645 B.n85 112.906
R1104 B.n639 B.n85 112.906
R1105 B.n639 B.n638 112.906
R1106 B.n637 B.n92 112.906
R1107 B.n631 B.n92 112.906
R1108 B.n631 B.n630 112.906
R1109 B.n630 B.n629 112.906
R1110 B.n629 B.n99 112.906
R1111 B.n623 B.n99 112.906
R1112 B.n623 B.n622 112.906
R1113 B.t0 B.n221 109.585
R1114 B.n694 B.t5 109.585
R1115 B.n450 B.t7 99.6231
R1116 B.n60 B.t1 99.6231
R1117 B.t2 B.n205 92.9816
R1118 B.n710 B.t23 92.9816
R1119 B.n425 B.t4 83.0194
R1120 B.n74 B.t22 83.0194
R1121 B.t3 B.n189 76.3779
R1122 B.n726 B.t6 76.3779
R1123 B.n370 B.n369 71.676
R1124 B.n364 B.n295 71.676
R1125 B.n361 B.n296 71.676
R1126 B.n357 B.n297 71.676
R1127 B.n353 B.n298 71.676
R1128 B.n348 B.n299 71.676
R1129 B.n344 B.n300 71.676
R1130 B.n340 B.n301 71.676
R1131 B.n336 B.n302 71.676
R1132 B.n332 B.n303 71.676
R1133 B.n327 B.n304 71.676
R1134 B.n323 B.n305 71.676
R1135 B.n319 B.n306 71.676
R1136 B.n315 B.n307 71.676
R1137 B.n126 B.n105 71.676
R1138 B.n130 B.n106 71.676
R1139 B.n134 B.n107 71.676
R1140 B.n138 B.n108 71.676
R1141 B.n142 B.n109 71.676
R1142 B.n146 B.n110 71.676
R1143 B.n150 B.n111 71.676
R1144 B.n154 B.n112 71.676
R1145 B.n158 B.n113 71.676
R1146 B.n162 B.n114 71.676
R1147 B.n166 B.n115 71.676
R1148 B.n170 B.n116 71.676
R1149 B.n174 B.n117 71.676
R1150 B.n178 B.n118 71.676
R1151 B.n620 B.n119 71.676
R1152 B.n620 B.n619 71.676
R1153 B.n180 B.n118 71.676
R1154 B.n177 B.n117 71.676
R1155 B.n173 B.n116 71.676
R1156 B.n169 B.n115 71.676
R1157 B.n165 B.n114 71.676
R1158 B.n161 B.n113 71.676
R1159 B.n157 B.n112 71.676
R1160 B.n153 B.n111 71.676
R1161 B.n149 B.n110 71.676
R1162 B.n145 B.n109 71.676
R1163 B.n141 B.n108 71.676
R1164 B.n137 B.n107 71.676
R1165 B.n133 B.n106 71.676
R1166 B.n129 B.n105 71.676
R1167 B.n370 B.n309 71.676
R1168 B.n362 B.n295 71.676
R1169 B.n358 B.n296 71.676
R1170 B.n354 B.n297 71.676
R1171 B.n349 B.n298 71.676
R1172 B.n345 B.n299 71.676
R1173 B.n341 B.n300 71.676
R1174 B.n337 B.n301 71.676
R1175 B.n333 B.n302 71.676
R1176 B.n328 B.n303 71.676
R1177 B.n324 B.n304 71.676
R1178 B.n320 B.n305 71.676
R1179 B.n316 B.n306 71.676
R1180 B.n307 B.n294 71.676
R1181 B.t13 B.n275 69.7364
R1182 B.n638 B.t9 69.7364
R1183 B.n330 B.n313 59.5399
R1184 B.n351 B.n311 59.5399
R1185 B.n125 B.n124 59.5399
R1186 B.n122 B.n121 59.5399
R1187 B.n313 B.n312 53.7217
R1188 B.n311 B.n310 53.7217
R1189 B.n124 B.n123 53.7217
R1190 B.n121 B.n120 53.7217
R1191 B.n395 B.t13 43.1703
R1192 B.t9 B.n637 43.1703
R1193 B.n529 B.t3 36.5288
R1194 B.t6 B.n725 36.5288
R1195 B.n127 B.n101 33.2493
R1196 B.n618 B.n617 33.2493
R1197 B.n374 B.n373 33.2493
R1198 B.n368 B.n289 33.2493
R1199 B.n432 B.t4 29.8873
R1200 B.n661 B.t22 29.8873
R1201 B.n505 B.t2 19.925
R1202 B.t23 B.n709 19.925
R1203 B B.n737 18.0485
R1204 B.n457 B.t7 13.2835
R1205 B.n677 B.t1 13.2835
R1206 B.n128 B.n127 10.6151
R1207 B.n131 B.n128 10.6151
R1208 B.n132 B.n131 10.6151
R1209 B.n135 B.n132 10.6151
R1210 B.n136 B.n135 10.6151
R1211 B.n139 B.n136 10.6151
R1212 B.n140 B.n139 10.6151
R1213 B.n143 B.n140 10.6151
R1214 B.n144 B.n143 10.6151
R1215 B.n148 B.n147 10.6151
R1216 B.n151 B.n148 10.6151
R1217 B.n152 B.n151 10.6151
R1218 B.n155 B.n152 10.6151
R1219 B.n156 B.n155 10.6151
R1220 B.n159 B.n156 10.6151
R1221 B.n160 B.n159 10.6151
R1222 B.n163 B.n160 10.6151
R1223 B.n164 B.n163 10.6151
R1224 B.n168 B.n167 10.6151
R1225 B.n171 B.n168 10.6151
R1226 B.n172 B.n171 10.6151
R1227 B.n175 B.n172 10.6151
R1228 B.n176 B.n175 10.6151
R1229 B.n179 B.n176 10.6151
R1230 B.n181 B.n179 10.6151
R1231 B.n182 B.n181 10.6151
R1232 B.n618 B.n182 10.6151
R1233 B.n375 B.n374 10.6151
R1234 B.n375 B.n285 10.6151
R1235 B.n385 B.n285 10.6151
R1236 B.n386 B.n385 10.6151
R1237 B.n387 B.n386 10.6151
R1238 B.n387 B.n277 10.6151
R1239 B.n397 B.n277 10.6151
R1240 B.n398 B.n397 10.6151
R1241 B.n399 B.n398 10.6151
R1242 B.n399 B.n269 10.6151
R1243 B.n409 B.n269 10.6151
R1244 B.n410 B.n409 10.6151
R1245 B.n411 B.n410 10.6151
R1246 B.n411 B.n261 10.6151
R1247 B.n421 B.n261 10.6151
R1248 B.n422 B.n421 10.6151
R1249 B.n423 B.n422 10.6151
R1250 B.n423 B.n254 10.6151
R1251 B.n434 B.n254 10.6151
R1252 B.n435 B.n434 10.6151
R1253 B.n436 B.n435 10.6151
R1254 B.n436 B.n246 10.6151
R1255 B.n446 B.n246 10.6151
R1256 B.n447 B.n446 10.6151
R1257 B.n448 B.n447 10.6151
R1258 B.n448 B.n239 10.6151
R1259 B.n459 B.n239 10.6151
R1260 B.n460 B.n459 10.6151
R1261 B.n461 B.n460 10.6151
R1262 B.n461 B.n231 10.6151
R1263 B.n471 B.n231 10.6151
R1264 B.n472 B.n471 10.6151
R1265 B.n473 B.n472 10.6151
R1266 B.n473 B.n223 10.6151
R1267 B.n483 B.n223 10.6151
R1268 B.n484 B.n483 10.6151
R1269 B.n485 B.n484 10.6151
R1270 B.n485 B.n215 10.6151
R1271 B.n495 B.n215 10.6151
R1272 B.n496 B.n495 10.6151
R1273 B.n497 B.n496 10.6151
R1274 B.n497 B.n207 10.6151
R1275 B.n507 B.n207 10.6151
R1276 B.n508 B.n507 10.6151
R1277 B.n509 B.n508 10.6151
R1278 B.n509 B.n199 10.6151
R1279 B.n519 B.n199 10.6151
R1280 B.n520 B.n519 10.6151
R1281 B.n521 B.n520 10.6151
R1282 B.n521 B.n191 10.6151
R1283 B.n531 B.n191 10.6151
R1284 B.n532 B.n531 10.6151
R1285 B.n534 B.n532 10.6151
R1286 B.n534 B.n533 10.6151
R1287 B.n533 B.n183 10.6151
R1288 B.n545 B.n183 10.6151
R1289 B.n546 B.n545 10.6151
R1290 B.n547 B.n546 10.6151
R1291 B.n548 B.n547 10.6151
R1292 B.n550 B.n548 10.6151
R1293 B.n551 B.n550 10.6151
R1294 B.n552 B.n551 10.6151
R1295 B.n553 B.n552 10.6151
R1296 B.n555 B.n553 10.6151
R1297 B.n556 B.n555 10.6151
R1298 B.n557 B.n556 10.6151
R1299 B.n558 B.n557 10.6151
R1300 B.n560 B.n558 10.6151
R1301 B.n561 B.n560 10.6151
R1302 B.n562 B.n561 10.6151
R1303 B.n563 B.n562 10.6151
R1304 B.n565 B.n563 10.6151
R1305 B.n566 B.n565 10.6151
R1306 B.n567 B.n566 10.6151
R1307 B.n568 B.n567 10.6151
R1308 B.n570 B.n568 10.6151
R1309 B.n571 B.n570 10.6151
R1310 B.n572 B.n571 10.6151
R1311 B.n573 B.n572 10.6151
R1312 B.n575 B.n573 10.6151
R1313 B.n576 B.n575 10.6151
R1314 B.n577 B.n576 10.6151
R1315 B.n578 B.n577 10.6151
R1316 B.n580 B.n578 10.6151
R1317 B.n581 B.n580 10.6151
R1318 B.n582 B.n581 10.6151
R1319 B.n583 B.n582 10.6151
R1320 B.n585 B.n583 10.6151
R1321 B.n586 B.n585 10.6151
R1322 B.n587 B.n586 10.6151
R1323 B.n588 B.n587 10.6151
R1324 B.n590 B.n588 10.6151
R1325 B.n591 B.n590 10.6151
R1326 B.n592 B.n591 10.6151
R1327 B.n593 B.n592 10.6151
R1328 B.n595 B.n593 10.6151
R1329 B.n596 B.n595 10.6151
R1330 B.n597 B.n596 10.6151
R1331 B.n598 B.n597 10.6151
R1332 B.n600 B.n598 10.6151
R1333 B.n601 B.n600 10.6151
R1334 B.n602 B.n601 10.6151
R1335 B.n603 B.n602 10.6151
R1336 B.n605 B.n603 10.6151
R1337 B.n606 B.n605 10.6151
R1338 B.n607 B.n606 10.6151
R1339 B.n608 B.n607 10.6151
R1340 B.n610 B.n608 10.6151
R1341 B.n611 B.n610 10.6151
R1342 B.n612 B.n611 10.6151
R1343 B.n613 B.n612 10.6151
R1344 B.n615 B.n613 10.6151
R1345 B.n616 B.n615 10.6151
R1346 B.n617 B.n616 10.6151
R1347 B.n368 B.n367 10.6151
R1348 B.n367 B.n366 10.6151
R1349 B.n366 B.n365 10.6151
R1350 B.n365 B.n363 10.6151
R1351 B.n363 B.n360 10.6151
R1352 B.n360 B.n359 10.6151
R1353 B.n359 B.n356 10.6151
R1354 B.n356 B.n355 10.6151
R1355 B.n355 B.n352 10.6151
R1356 B.n350 B.n347 10.6151
R1357 B.n347 B.n346 10.6151
R1358 B.n346 B.n343 10.6151
R1359 B.n343 B.n342 10.6151
R1360 B.n342 B.n339 10.6151
R1361 B.n339 B.n338 10.6151
R1362 B.n338 B.n335 10.6151
R1363 B.n335 B.n334 10.6151
R1364 B.n334 B.n331 10.6151
R1365 B.n329 B.n326 10.6151
R1366 B.n326 B.n325 10.6151
R1367 B.n325 B.n322 10.6151
R1368 B.n322 B.n321 10.6151
R1369 B.n321 B.n318 10.6151
R1370 B.n318 B.n317 10.6151
R1371 B.n317 B.n314 10.6151
R1372 B.n314 B.n293 10.6151
R1373 B.n373 B.n293 10.6151
R1374 B.n379 B.n289 10.6151
R1375 B.n380 B.n379 10.6151
R1376 B.n381 B.n380 10.6151
R1377 B.n381 B.n281 10.6151
R1378 B.n391 B.n281 10.6151
R1379 B.n392 B.n391 10.6151
R1380 B.n393 B.n392 10.6151
R1381 B.n393 B.n273 10.6151
R1382 B.n403 B.n273 10.6151
R1383 B.n404 B.n403 10.6151
R1384 B.n405 B.n404 10.6151
R1385 B.n405 B.n265 10.6151
R1386 B.n415 B.n265 10.6151
R1387 B.n416 B.n415 10.6151
R1388 B.n417 B.n416 10.6151
R1389 B.n417 B.n257 10.6151
R1390 B.n428 B.n257 10.6151
R1391 B.n429 B.n428 10.6151
R1392 B.n430 B.n429 10.6151
R1393 B.n430 B.n250 10.6151
R1394 B.n440 B.n250 10.6151
R1395 B.n441 B.n440 10.6151
R1396 B.n442 B.n441 10.6151
R1397 B.n442 B.n242 10.6151
R1398 B.n453 B.n242 10.6151
R1399 B.n454 B.n453 10.6151
R1400 B.n455 B.n454 10.6151
R1401 B.n455 B.n235 10.6151
R1402 B.n465 B.n235 10.6151
R1403 B.n466 B.n465 10.6151
R1404 B.n467 B.n466 10.6151
R1405 B.n467 B.n227 10.6151
R1406 B.n477 B.n227 10.6151
R1407 B.n478 B.n477 10.6151
R1408 B.n479 B.n478 10.6151
R1409 B.n479 B.n219 10.6151
R1410 B.n489 B.n219 10.6151
R1411 B.n490 B.n489 10.6151
R1412 B.n491 B.n490 10.6151
R1413 B.n491 B.n211 10.6151
R1414 B.n501 B.n211 10.6151
R1415 B.n502 B.n501 10.6151
R1416 B.n503 B.n502 10.6151
R1417 B.n503 B.n203 10.6151
R1418 B.n513 B.n203 10.6151
R1419 B.n514 B.n513 10.6151
R1420 B.n515 B.n514 10.6151
R1421 B.n515 B.n195 10.6151
R1422 B.n525 B.n195 10.6151
R1423 B.n526 B.n525 10.6151
R1424 B.n527 B.n526 10.6151
R1425 B.n527 B.n187 10.6151
R1426 B.n538 B.n187 10.6151
R1427 B.n539 B.n538 10.6151
R1428 B.n540 B.n539 10.6151
R1429 B.n540 B.n0 10.6151
R1430 B.n731 B.n1 10.6151
R1431 B.n731 B.n730 10.6151
R1432 B.n730 B.n729 10.6151
R1433 B.n729 B.n10 10.6151
R1434 B.n723 B.n10 10.6151
R1435 B.n723 B.n722 10.6151
R1436 B.n722 B.n721 10.6151
R1437 B.n721 B.n17 10.6151
R1438 B.n715 B.n17 10.6151
R1439 B.n715 B.n714 10.6151
R1440 B.n714 B.n713 10.6151
R1441 B.n713 B.n24 10.6151
R1442 B.n707 B.n24 10.6151
R1443 B.n707 B.n706 10.6151
R1444 B.n706 B.n705 10.6151
R1445 B.n705 B.n31 10.6151
R1446 B.n699 B.n31 10.6151
R1447 B.n699 B.n698 10.6151
R1448 B.n698 B.n697 10.6151
R1449 B.n697 B.n38 10.6151
R1450 B.n691 B.n38 10.6151
R1451 B.n691 B.n690 10.6151
R1452 B.n690 B.n689 10.6151
R1453 B.n689 B.n45 10.6151
R1454 B.n683 B.n45 10.6151
R1455 B.n683 B.n682 10.6151
R1456 B.n682 B.n681 10.6151
R1457 B.n681 B.n52 10.6151
R1458 B.n675 B.n52 10.6151
R1459 B.n675 B.n674 10.6151
R1460 B.n674 B.n673 10.6151
R1461 B.n673 B.n58 10.6151
R1462 B.n667 B.n58 10.6151
R1463 B.n667 B.n666 10.6151
R1464 B.n666 B.n665 10.6151
R1465 B.n665 B.n66 10.6151
R1466 B.n659 B.n66 10.6151
R1467 B.n659 B.n658 10.6151
R1468 B.n658 B.n657 10.6151
R1469 B.n657 B.n72 10.6151
R1470 B.n651 B.n72 10.6151
R1471 B.n651 B.n650 10.6151
R1472 B.n650 B.n649 10.6151
R1473 B.n649 B.n80 10.6151
R1474 B.n643 B.n80 10.6151
R1475 B.n643 B.n642 10.6151
R1476 B.n642 B.n641 10.6151
R1477 B.n641 B.n87 10.6151
R1478 B.n635 B.n87 10.6151
R1479 B.n635 B.n634 10.6151
R1480 B.n634 B.n633 10.6151
R1481 B.n633 B.n94 10.6151
R1482 B.n627 B.n94 10.6151
R1483 B.n627 B.n626 10.6151
R1484 B.n626 B.n625 10.6151
R1485 B.n625 B.n101 10.6151
R1486 B.n144 B.n125 9.36635
R1487 B.n167 B.n122 9.36635
R1488 B.n352 B.n351 9.36635
R1489 B.n330 B.n329 9.36635
R1490 B.n481 B.t0 3.32125
R1491 B.t5 B.n693 3.32125
R1492 B.n737 B.n0 2.81026
R1493 B.n737 B.n1 2.81026
R1494 B.n147 B.n125 1.24928
R1495 B.n164 B.n122 1.24928
R1496 B.n351 B.n350 1.24928
R1497 B.n331 B.n330 1.24928
R1498 VP.n23 VP.n20 161.3
R1499 VP.n25 VP.n24 161.3
R1500 VP.n26 VP.n19 161.3
R1501 VP.n28 VP.n27 161.3
R1502 VP.n29 VP.n18 161.3
R1503 VP.n32 VP.n31 161.3
R1504 VP.n33 VP.n17 161.3
R1505 VP.n35 VP.n34 161.3
R1506 VP.n36 VP.n16 161.3
R1507 VP.n38 VP.n37 161.3
R1508 VP.n39 VP.n15 161.3
R1509 VP.n41 VP.n40 161.3
R1510 VP.n43 VP.n14 161.3
R1511 VP.n45 VP.n44 161.3
R1512 VP.n46 VP.n13 161.3
R1513 VP.n48 VP.n47 161.3
R1514 VP.n49 VP.n12 161.3
R1515 VP.n88 VP.n0 161.3
R1516 VP.n87 VP.n86 161.3
R1517 VP.n85 VP.n1 161.3
R1518 VP.n84 VP.n83 161.3
R1519 VP.n82 VP.n2 161.3
R1520 VP.n80 VP.n79 161.3
R1521 VP.n78 VP.n3 161.3
R1522 VP.n77 VP.n76 161.3
R1523 VP.n75 VP.n4 161.3
R1524 VP.n74 VP.n73 161.3
R1525 VP.n72 VP.n5 161.3
R1526 VP.n71 VP.n70 161.3
R1527 VP.n68 VP.n6 161.3
R1528 VP.n67 VP.n66 161.3
R1529 VP.n65 VP.n7 161.3
R1530 VP.n64 VP.n63 161.3
R1531 VP.n62 VP.n8 161.3
R1532 VP.n60 VP.n59 161.3
R1533 VP.n58 VP.n9 161.3
R1534 VP.n57 VP.n56 161.3
R1535 VP.n55 VP.n10 161.3
R1536 VP.n54 VP.n53 161.3
R1537 VP.n52 VP.n11 96.5656
R1538 VP.n90 VP.n89 96.5656
R1539 VP.n51 VP.n50 96.5656
R1540 VP.n22 VP.n21 71.4859
R1541 VP.n67 VP.n7 53.6055
R1542 VP.n76 VP.n75 53.6055
R1543 VP.n37 VP.n36 53.6055
R1544 VP.n28 VP.n19 53.6055
R1545 VP.n56 VP.n9 49.7204
R1546 VP.n83 VP.n1 49.7204
R1547 VP.n44 VP.n13 49.7204
R1548 VP.n21 VP.t8 45.4455
R1549 VP.n52 VP.n51 44.2231
R1550 VP.n56 VP.n55 31.2664
R1551 VP.n87 VP.n1 31.2664
R1552 VP.n48 VP.n13 31.2664
R1553 VP.n68 VP.n67 27.3813
R1554 VP.n75 VP.n74 27.3813
R1555 VP.n36 VP.n35 27.3813
R1556 VP.n29 VP.n28 27.3813
R1557 VP.n55 VP.n54 24.4675
R1558 VP.n60 VP.n9 24.4675
R1559 VP.n63 VP.n62 24.4675
R1560 VP.n63 VP.n7 24.4675
R1561 VP.n70 VP.n68 24.4675
R1562 VP.n74 VP.n5 24.4675
R1563 VP.n76 VP.n3 24.4675
R1564 VP.n80 VP.n3 24.4675
R1565 VP.n83 VP.n82 24.4675
R1566 VP.n88 VP.n87 24.4675
R1567 VP.n49 VP.n48 24.4675
R1568 VP.n37 VP.n15 24.4675
R1569 VP.n41 VP.n15 24.4675
R1570 VP.n44 VP.n43 24.4675
R1571 VP.n31 VP.n29 24.4675
R1572 VP.n35 VP.n17 24.4675
R1573 VP.n24 VP.n23 24.4675
R1574 VP.n24 VP.n19 24.4675
R1575 VP.n61 VP.n60 23.4888
R1576 VP.n82 VP.n81 23.4888
R1577 VP.n43 VP.n42 23.4888
R1578 VP.n54 VP.n11 14.1914
R1579 VP.n89 VP.n88 14.1914
R1580 VP.n50 VP.n49 14.1914
R1581 VP.n11 VP.t1 13.3345
R1582 VP.n61 VP.t5 13.3345
R1583 VP.n69 VP.t4 13.3345
R1584 VP.n81 VP.t2 13.3345
R1585 VP.n89 VP.t0 13.3345
R1586 VP.n50 VP.t7 13.3345
R1587 VP.n42 VP.t3 13.3345
R1588 VP.n30 VP.t9 13.3345
R1589 VP.n22 VP.t6 13.3345
R1590 VP.n70 VP.n69 12.234
R1591 VP.n69 VP.n5 12.234
R1592 VP.n31 VP.n30 12.234
R1593 VP.n30 VP.n17 12.234
R1594 VP.n21 VP.n20 9.60581
R1595 VP.n62 VP.n61 0.97918
R1596 VP.n81 VP.n80 0.97918
R1597 VP.n42 VP.n41 0.97918
R1598 VP.n23 VP.n22 0.97918
R1599 VP.n51 VP.n12 0.278367
R1600 VP.n53 VP.n52 0.278367
R1601 VP.n90 VP.n0 0.278367
R1602 VP.n25 VP.n20 0.189894
R1603 VP.n26 VP.n25 0.189894
R1604 VP.n27 VP.n26 0.189894
R1605 VP.n27 VP.n18 0.189894
R1606 VP.n32 VP.n18 0.189894
R1607 VP.n33 VP.n32 0.189894
R1608 VP.n34 VP.n33 0.189894
R1609 VP.n34 VP.n16 0.189894
R1610 VP.n38 VP.n16 0.189894
R1611 VP.n39 VP.n38 0.189894
R1612 VP.n40 VP.n39 0.189894
R1613 VP.n40 VP.n14 0.189894
R1614 VP.n45 VP.n14 0.189894
R1615 VP.n46 VP.n45 0.189894
R1616 VP.n47 VP.n46 0.189894
R1617 VP.n47 VP.n12 0.189894
R1618 VP.n53 VP.n10 0.189894
R1619 VP.n57 VP.n10 0.189894
R1620 VP.n58 VP.n57 0.189894
R1621 VP.n59 VP.n58 0.189894
R1622 VP.n59 VP.n8 0.189894
R1623 VP.n64 VP.n8 0.189894
R1624 VP.n65 VP.n64 0.189894
R1625 VP.n66 VP.n65 0.189894
R1626 VP.n66 VP.n6 0.189894
R1627 VP.n71 VP.n6 0.189894
R1628 VP.n72 VP.n71 0.189894
R1629 VP.n73 VP.n72 0.189894
R1630 VP.n73 VP.n4 0.189894
R1631 VP.n77 VP.n4 0.189894
R1632 VP.n78 VP.n77 0.189894
R1633 VP.n79 VP.n78 0.189894
R1634 VP.n79 VP.n2 0.189894
R1635 VP.n84 VP.n2 0.189894
R1636 VP.n85 VP.n84 0.189894
R1637 VP.n86 VP.n85 0.189894
R1638 VP.n86 VP.n0 0.189894
R1639 VP VP.n90 0.153454
R1640 VDD1.n3 VDD1.t8 176.333
R1641 VDD1.n1 VDD1.t1 176.333
R1642 VDD1.n5 VDD1.n4 149.523
R1643 VDD1.n7 VDD1.n6 147.786
R1644 VDD1.n3 VDD1.n2 147.786
R1645 VDD1.n1 VDD1.n0 147.786
R1646 VDD1.n7 VDD1.n5 37.9987
R1647 VDD1.n6 VDD1.t6 14.6672
R1648 VDD1.n6 VDD1.t2 14.6672
R1649 VDD1.n0 VDD1.t3 14.6672
R1650 VDD1.n0 VDD1.t0 14.6672
R1651 VDD1.n4 VDD1.t7 14.6672
R1652 VDD1.n4 VDD1.t9 14.6672
R1653 VDD1.n2 VDD1.t4 14.6672
R1654 VDD1.n2 VDD1.t5 14.6672
R1655 VDD1 VDD1.n7 1.73326
R1656 VDD1 VDD1.n1 0.655672
R1657 VDD1.n5 VDD1.n3 0.542137
C0 VN VTAIL 3.05865f
C1 VTAIL VDD1 5.29794f
C2 VP VDD2 0.571408f
C3 VP VN 6.19752f
C4 VDD2 VN 1.64493f
C5 VP VDD1 2.05185f
C6 VP VTAIL 3.07278f
C7 VDD2 VDD1 2.06871f
C8 VDD2 VTAIL 5.35026f
C9 VN VDD1 0.160404f
C10 VDD2 B 5.144701f
C11 VDD1 B 5.142118f
C12 VTAIL B 3.337582f
C13 VN B 16.34097f
C14 VP B 14.898612f
C15 VDD1.t1 B 0.232004f
C16 VDD1.t3 B 0.03371f
C17 VDD1.t0 B 0.03371f
C18 VDD1.n0 B 0.169215f
C19 VDD1.n1 B 1.05876f
C20 VDD1.t8 B 0.232004f
C21 VDD1.t4 B 0.03371f
C22 VDD1.t5 B 0.03371f
C23 VDD1.n2 B 0.169216f
C24 VDD1.n3 B 1.04855f
C25 VDD1.t7 B 0.03371f
C26 VDD1.t9 B 0.03371f
C27 VDD1.n4 B 0.176934f
C28 VDD1.n5 B 2.88414f
C29 VDD1.t6 B 0.03371f
C30 VDD1.t2 B 0.03371f
C31 VDD1.n6 B 0.169216f
C32 VDD1.n7 B 2.84714f
C33 VP.n0 B 0.044839f
C34 VP.t0 B 0.236436f
C35 VP.n1 B 0.031653f
C36 VP.n2 B 0.03401f
C37 VP.t2 B 0.236436f
C38 VP.n3 B 0.063386f
C39 VP.n4 B 0.03401f
C40 VP.n5 B 0.047739f
C41 VP.n6 B 0.03401f
C42 VP.n7 B 0.059984f
C43 VP.n8 B 0.03401f
C44 VP.t5 B 0.236436f
C45 VP.n9 B 0.06275f
C46 VP.n10 B 0.03401f
C47 VP.t1 B 0.236436f
C48 VP.n11 B 0.2508f
C49 VP.n12 B 0.044839f
C50 VP.t7 B 0.236436f
C51 VP.n13 B 0.031653f
C52 VP.n14 B 0.03401f
C53 VP.t3 B 0.236436f
C54 VP.n15 B 0.063386f
C55 VP.n16 B 0.03401f
C56 VP.n17 B 0.047739f
C57 VP.n18 B 0.03401f
C58 VP.n19 B 0.059984f
C59 VP.n20 B 0.297678f
C60 VP.t6 B 0.236436f
C61 VP.t8 B 0.471083f
C62 VP.n21 B 0.221107f
C63 VP.n22 B 0.217674f
C64 VP.n23 B 0.033344f
C65 VP.n24 B 0.063386f
C66 VP.n25 B 0.03401f
C67 VP.n26 B 0.03401f
C68 VP.n27 B 0.03401f
C69 VP.n28 B 0.036388f
C70 VP.n29 B 0.066316f
C71 VP.t9 B 0.236436f
C72 VP.n30 B 0.135946f
C73 VP.n31 B 0.047739f
C74 VP.n32 B 0.03401f
C75 VP.n33 B 0.03401f
C76 VP.n34 B 0.03401f
C77 VP.n35 B 0.066316f
C78 VP.n36 B 0.036388f
C79 VP.n37 B 0.059984f
C80 VP.n38 B 0.03401f
C81 VP.n39 B 0.03401f
C82 VP.n40 B 0.03401f
C83 VP.n41 B 0.033344f
C84 VP.n42 B 0.135946f
C85 VP.n43 B 0.062134f
C86 VP.n44 B 0.06275f
C87 VP.n45 B 0.03401f
C88 VP.n46 B 0.03401f
C89 VP.n47 B 0.03401f
C90 VP.n48 B 0.068285f
C91 VP.n49 B 0.050242f
C92 VP.n50 B 0.2508f
C93 VP.n51 B 1.56584f
C94 VP.n52 B 1.59348f
C95 VP.n53 B 0.044839f
C96 VP.n54 B 0.050242f
C97 VP.n55 B 0.068285f
C98 VP.n56 B 0.031653f
C99 VP.n57 B 0.03401f
C100 VP.n58 B 0.03401f
C101 VP.n59 B 0.03401f
C102 VP.n60 B 0.062134f
C103 VP.n61 B 0.135946f
C104 VP.n62 B 0.033344f
C105 VP.n63 B 0.063386f
C106 VP.n64 B 0.03401f
C107 VP.n65 B 0.03401f
C108 VP.n66 B 0.03401f
C109 VP.n67 B 0.036388f
C110 VP.n68 B 0.066316f
C111 VP.t4 B 0.236436f
C112 VP.n69 B 0.135946f
C113 VP.n70 B 0.047739f
C114 VP.n71 B 0.03401f
C115 VP.n72 B 0.03401f
C116 VP.n73 B 0.03401f
C117 VP.n74 B 0.066316f
C118 VP.n75 B 0.036388f
C119 VP.n76 B 0.059984f
C120 VP.n77 B 0.03401f
C121 VP.n78 B 0.03401f
C122 VP.n79 B 0.03401f
C123 VP.n80 B 0.033344f
C124 VP.n81 B 0.135946f
C125 VP.n82 B 0.062134f
C126 VP.n83 B 0.06275f
C127 VP.n84 B 0.03401f
C128 VP.n85 B 0.03401f
C129 VP.n86 B 0.03401f
C130 VP.n87 B 0.068285f
C131 VP.n88 B 0.050242f
C132 VP.n89 B 0.2508f
C133 VP.n90 B 0.049895f
C134 VTAIL.t11 B 0.042442f
C135 VTAIL.t14 B 0.042442f
C136 VTAIL.n0 B 0.176857f
C137 VTAIL.n1 B 0.724465f
C138 VTAIL.t3 B 0.248152f
C139 VTAIL.n2 B 0.837989f
C140 VTAIL.t0 B 0.042442f
C141 VTAIL.t2 B 0.042442f
C142 VTAIL.n3 B 0.176857f
C143 VTAIL.n4 B 0.886362f
C144 VTAIL.t4 B 0.042442f
C145 VTAIL.t7 B 0.042442f
C146 VTAIL.n5 B 0.176857f
C147 VTAIL.n6 B 1.88207f
C148 VTAIL.t10 B 0.042442f
C149 VTAIL.t18 B 0.042442f
C150 VTAIL.n7 B 0.176856f
C151 VTAIL.n8 B 1.88208f
C152 VTAIL.t9 B 0.042442f
C153 VTAIL.t13 B 0.042442f
C154 VTAIL.n9 B 0.176856f
C155 VTAIL.n10 B 0.886363f
C156 VTAIL.t12 B 0.248152f
C157 VTAIL.n11 B 0.837989f
C158 VTAIL.t6 B 0.042442f
C159 VTAIL.t19 B 0.042442f
C160 VTAIL.n12 B 0.176856f
C161 VTAIL.n13 B 0.793535f
C162 VTAIL.t5 B 0.042442f
C163 VTAIL.t1 B 0.042442f
C164 VTAIL.n14 B 0.176856f
C165 VTAIL.n15 B 0.886363f
C166 VTAIL.t8 B 0.248152f
C167 VTAIL.n16 B 1.62042f
C168 VTAIL.t17 B 0.248152f
C169 VTAIL.n17 B 1.62042f
C170 VTAIL.t15 B 0.042442f
C171 VTAIL.t16 B 0.042442f
C172 VTAIL.n18 B 0.176857f
C173 VTAIL.n19 B 0.649319f
C174 VDD2.t6 B 0.185439f
C175 VDD2.t2 B 0.026944f
C176 VDD2.t5 B 0.026944f
C177 VDD2.n0 B 0.135253f
C178 VDD2.n1 B 0.838102f
C179 VDD2.t8 B 0.026944f
C180 VDD2.t4 B 0.026944f
C181 VDD2.n2 B 0.141422f
C182 VDD2.n3 B 2.19314f
C183 VDD2.t0 B 0.179767f
C184 VDD2.n4 B 2.1825f
C185 VDD2.t3 B 0.026944f
C186 VDD2.t9 B 0.026944f
C187 VDD2.n5 B 0.135253f
C188 VDD2.n6 B 0.433055f
C189 VDD2.t1 B 0.026944f
C190 VDD2.t7 B 0.026944f
C191 VDD2.n7 B 0.141406f
C192 VN.n0 B 0.036426f
C193 VN.t1 B 0.192076f
C194 VN.n1 B 0.025715f
C195 VN.n2 B 0.027629f
C196 VN.t2 B 0.192076f
C197 VN.n3 B 0.051493f
C198 VN.n4 B 0.027629f
C199 VN.n5 B 0.038782f
C200 VN.n6 B 0.027629f
C201 VN.n7 B 0.04873f
C202 VN.n8 B 0.241828f
C203 VN.t4 B 0.192076f
C204 VN.t7 B 0.382699f
C205 VN.n9 B 0.179624f
C206 VN.n10 B 0.176834f
C207 VN.n11 B 0.027088f
C208 VN.n12 B 0.051493f
C209 VN.n13 B 0.027629f
C210 VN.n14 B 0.027629f
C211 VN.n15 B 0.027629f
C212 VN.n16 B 0.029561f
C213 VN.n17 B 0.053874f
C214 VN.t3 B 0.192076f
C215 VN.n18 B 0.11044f
C216 VN.n19 B 0.038782f
C217 VN.n20 B 0.027629f
C218 VN.n21 B 0.027629f
C219 VN.n22 B 0.027629f
C220 VN.n23 B 0.053874f
C221 VN.n24 B 0.029561f
C222 VN.n25 B 0.04873f
C223 VN.n26 B 0.027629f
C224 VN.n27 B 0.027629f
C225 VN.n28 B 0.027629f
C226 VN.n29 B 0.027088f
C227 VN.n30 B 0.11044f
C228 VN.n31 B 0.050477f
C229 VN.n32 B 0.050977f
C230 VN.n33 B 0.027629f
C231 VN.n34 B 0.027629f
C232 VN.n35 B 0.027629f
C233 VN.n36 B 0.055474f
C234 VN.n37 B 0.040816f
C235 VN.n38 B 0.203745f
C236 VN.n39 B 0.040534f
C237 VN.n40 B 0.036426f
C238 VN.t8 B 0.192076f
C239 VN.n41 B 0.025715f
C240 VN.n42 B 0.027629f
C241 VN.t0 B 0.192076f
C242 VN.n43 B 0.051493f
C243 VN.n44 B 0.027629f
C244 VN.n45 B 0.038782f
C245 VN.n46 B 0.027629f
C246 VN.t9 B 0.192076f
C247 VN.n47 B 0.11044f
C248 VN.n48 B 0.04873f
C249 VN.n49 B 0.241828f
C250 VN.t5 B 0.192076f
C251 VN.t6 B 0.382699f
C252 VN.n50 B 0.179624f
C253 VN.n51 B 0.176834f
C254 VN.n52 B 0.027088f
C255 VN.n53 B 0.051493f
C256 VN.n54 B 0.027629f
C257 VN.n55 B 0.027629f
C258 VN.n56 B 0.027629f
C259 VN.n57 B 0.029561f
C260 VN.n58 B 0.053874f
C261 VN.n59 B 0.038782f
C262 VN.n60 B 0.027629f
C263 VN.n61 B 0.027629f
C264 VN.n62 B 0.027629f
C265 VN.n63 B 0.053874f
C266 VN.n64 B 0.029561f
C267 VN.n65 B 0.04873f
C268 VN.n66 B 0.027629f
C269 VN.n67 B 0.027629f
C270 VN.n68 B 0.027629f
C271 VN.n69 B 0.027088f
C272 VN.n70 B 0.11044f
C273 VN.n71 B 0.050477f
C274 VN.n72 B 0.050977f
C275 VN.n73 B 0.027629f
C276 VN.n74 B 0.027629f
C277 VN.n75 B 0.027629f
C278 VN.n76 B 0.055474f
C279 VN.n77 B 0.040816f
C280 VN.n78 B 0.203745f
C281 VN.n79 B 1.28721f
.ends

