* NGSPICE file created from diff_pair_sample_0792.ext - technology: sky130A

.subckt diff_pair_sample_0792 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t3 VN.t0 VTAIL.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=3.56
X1 VDD1.t3 VP.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=3.56
X2 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=3.56
X3 VTAIL.t6 VP.t1 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=3.56
X4 VTAIL.t2 VN.t1 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=3.56
X5 VTAIL.t4 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=3.56
X6 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=3.56
X7 VDD2.t1 VN.t2 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=3.56
X8 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=3.56
X9 VTAIL.t3 VN.t3 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=1.749 ps=10.93 w=10.6 l=3.56
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.134 pd=21.98 as=0 ps=0 w=10.6 l=3.56
X11 VDD1.t0 VP.t3 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=1.749 pd=10.93 as=4.134 ps=21.98 w=10.6 l=3.56
R0 VN.n1 VN.t2 106.547
R1 VN.n0 VN.t3 106.547
R2 VN.n0 VN.t0 105.311
R3 VN.n1 VN.t1 105.311
R4 VN VN.n1 50.5597
R5 VN VN.n0 2.1317
R6 VTAIL.n458 VTAIL.n406 289.615
R7 VTAIL.n52 VTAIL.n0 289.615
R8 VTAIL.n110 VTAIL.n58 289.615
R9 VTAIL.n168 VTAIL.n116 289.615
R10 VTAIL.n400 VTAIL.n348 289.615
R11 VTAIL.n342 VTAIL.n290 289.615
R12 VTAIL.n284 VTAIL.n232 289.615
R13 VTAIL.n226 VTAIL.n174 289.615
R14 VTAIL.n425 VTAIL.n424 185
R15 VTAIL.n422 VTAIL.n421 185
R16 VTAIL.n431 VTAIL.n430 185
R17 VTAIL.n433 VTAIL.n432 185
R18 VTAIL.n418 VTAIL.n417 185
R19 VTAIL.n439 VTAIL.n438 185
R20 VTAIL.n442 VTAIL.n441 185
R21 VTAIL.n440 VTAIL.n414 185
R22 VTAIL.n447 VTAIL.n413 185
R23 VTAIL.n449 VTAIL.n448 185
R24 VTAIL.n451 VTAIL.n450 185
R25 VTAIL.n410 VTAIL.n409 185
R26 VTAIL.n457 VTAIL.n456 185
R27 VTAIL.n459 VTAIL.n458 185
R28 VTAIL.n19 VTAIL.n18 185
R29 VTAIL.n16 VTAIL.n15 185
R30 VTAIL.n25 VTAIL.n24 185
R31 VTAIL.n27 VTAIL.n26 185
R32 VTAIL.n12 VTAIL.n11 185
R33 VTAIL.n33 VTAIL.n32 185
R34 VTAIL.n36 VTAIL.n35 185
R35 VTAIL.n34 VTAIL.n8 185
R36 VTAIL.n41 VTAIL.n7 185
R37 VTAIL.n43 VTAIL.n42 185
R38 VTAIL.n45 VTAIL.n44 185
R39 VTAIL.n4 VTAIL.n3 185
R40 VTAIL.n51 VTAIL.n50 185
R41 VTAIL.n53 VTAIL.n52 185
R42 VTAIL.n77 VTAIL.n76 185
R43 VTAIL.n74 VTAIL.n73 185
R44 VTAIL.n83 VTAIL.n82 185
R45 VTAIL.n85 VTAIL.n84 185
R46 VTAIL.n70 VTAIL.n69 185
R47 VTAIL.n91 VTAIL.n90 185
R48 VTAIL.n94 VTAIL.n93 185
R49 VTAIL.n92 VTAIL.n66 185
R50 VTAIL.n99 VTAIL.n65 185
R51 VTAIL.n101 VTAIL.n100 185
R52 VTAIL.n103 VTAIL.n102 185
R53 VTAIL.n62 VTAIL.n61 185
R54 VTAIL.n109 VTAIL.n108 185
R55 VTAIL.n111 VTAIL.n110 185
R56 VTAIL.n135 VTAIL.n134 185
R57 VTAIL.n132 VTAIL.n131 185
R58 VTAIL.n141 VTAIL.n140 185
R59 VTAIL.n143 VTAIL.n142 185
R60 VTAIL.n128 VTAIL.n127 185
R61 VTAIL.n149 VTAIL.n148 185
R62 VTAIL.n152 VTAIL.n151 185
R63 VTAIL.n150 VTAIL.n124 185
R64 VTAIL.n157 VTAIL.n123 185
R65 VTAIL.n159 VTAIL.n158 185
R66 VTAIL.n161 VTAIL.n160 185
R67 VTAIL.n120 VTAIL.n119 185
R68 VTAIL.n167 VTAIL.n166 185
R69 VTAIL.n169 VTAIL.n168 185
R70 VTAIL.n401 VTAIL.n400 185
R71 VTAIL.n399 VTAIL.n398 185
R72 VTAIL.n352 VTAIL.n351 185
R73 VTAIL.n393 VTAIL.n392 185
R74 VTAIL.n391 VTAIL.n390 185
R75 VTAIL.n389 VTAIL.n355 185
R76 VTAIL.n359 VTAIL.n356 185
R77 VTAIL.n384 VTAIL.n383 185
R78 VTAIL.n382 VTAIL.n381 185
R79 VTAIL.n361 VTAIL.n360 185
R80 VTAIL.n376 VTAIL.n375 185
R81 VTAIL.n374 VTAIL.n373 185
R82 VTAIL.n365 VTAIL.n364 185
R83 VTAIL.n368 VTAIL.n367 185
R84 VTAIL.n343 VTAIL.n342 185
R85 VTAIL.n341 VTAIL.n340 185
R86 VTAIL.n294 VTAIL.n293 185
R87 VTAIL.n335 VTAIL.n334 185
R88 VTAIL.n333 VTAIL.n332 185
R89 VTAIL.n331 VTAIL.n297 185
R90 VTAIL.n301 VTAIL.n298 185
R91 VTAIL.n326 VTAIL.n325 185
R92 VTAIL.n324 VTAIL.n323 185
R93 VTAIL.n303 VTAIL.n302 185
R94 VTAIL.n318 VTAIL.n317 185
R95 VTAIL.n316 VTAIL.n315 185
R96 VTAIL.n307 VTAIL.n306 185
R97 VTAIL.n310 VTAIL.n309 185
R98 VTAIL.n285 VTAIL.n284 185
R99 VTAIL.n283 VTAIL.n282 185
R100 VTAIL.n236 VTAIL.n235 185
R101 VTAIL.n277 VTAIL.n276 185
R102 VTAIL.n275 VTAIL.n274 185
R103 VTAIL.n273 VTAIL.n239 185
R104 VTAIL.n243 VTAIL.n240 185
R105 VTAIL.n268 VTAIL.n267 185
R106 VTAIL.n266 VTAIL.n265 185
R107 VTAIL.n245 VTAIL.n244 185
R108 VTAIL.n260 VTAIL.n259 185
R109 VTAIL.n258 VTAIL.n257 185
R110 VTAIL.n249 VTAIL.n248 185
R111 VTAIL.n252 VTAIL.n251 185
R112 VTAIL.n227 VTAIL.n226 185
R113 VTAIL.n225 VTAIL.n224 185
R114 VTAIL.n178 VTAIL.n177 185
R115 VTAIL.n219 VTAIL.n218 185
R116 VTAIL.n217 VTAIL.n216 185
R117 VTAIL.n215 VTAIL.n181 185
R118 VTAIL.n185 VTAIL.n182 185
R119 VTAIL.n210 VTAIL.n209 185
R120 VTAIL.n208 VTAIL.n207 185
R121 VTAIL.n187 VTAIL.n186 185
R122 VTAIL.n202 VTAIL.n201 185
R123 VTAIL.n200 VTAIL.n199 185
R124 VTAIL.n191 VTAIL.n190 185
R125 VTAIL.n194 VTAIL.n193 185
R126 VTAIL.t1 VTAIL.n423 149.524
R127 VTAIL.t3 VTAIL.n17 149.524
R128 VTAIL.t5 VTAIL.n75 149.524
R129 VTAIL.t6 VTAIL.n133 149.524
R130 VTAIL.t7 VTAIL.n366 149.524
R131 VTAIL.t4 VTAIL.n308 149.524
R132 VTAIL.t0 VTAIL.n250 149.524
R133 VTAIL.t2 VTAIL.n192 149.524
R134 VTAIL.n424 VTAIL.n421 104.615
R135 VTAIL.n431 VTAIL.n421 104.615
R136 VTAIL.n432 VTAIL.n431 104.615
R137 VTAIL.n432 VTAIL.n417 104.615
R138 VTAIL.n439 VTAIL.n417 104.615
R139 VTAIL.n441 VTAIL.n439 104.615
R140 VTAIL.n441 VTAIL.n440 104.615
R141 VTAIL.n440 VTAIL.n413 104.615
R142 VTAIL.n449 VTAIL.n413 104.615
R143 VTAIL.n450 VTAIL.n449 104.615
R144 VTAIL.n450 VTAIL.n409 104.615
R145 VTAIL.n457 VTAIL.n409 104.615
R146 VTAIL.n458 VTAIL.n457 104.615
R147 VTAIL.n18 VTAIL.n15 104.615
R148 VTAIL.n25 VTAIL.n15 104.615
R149 VTAIL.n26 VTAIL.n25 104.615
R150 VTAIL.n26 VTAIL.n11 104.615
R151 VTAIL.n33 VTAIL.n11 104.615
R152 VTAIL.n35 VTAIL.n33 104.615
R153 VTAIL.n35 VTAIL.n34 104.615
R154 VTAIL.n34 VTAIL.n7 104.615
R155 VTAIL.n43 VTAIL.n7 104.615
R156 VTAIL.n44 VTAIL.n43 104.615
R157 VTAIL.n44 VTAIL.n3 104.615
R158 VTAIL.n51 VTAIL.n3 104.615
R159 VTAIL.n52 VTAIL.n51 104.615
R160 VTAIL.n76 VTAIL.n73 104.615
R161 VTAIL.n83 VTAIL.n73 104.615
R162 VTAIL.n84 VTAIL.n83 104.615
R163 VTAIL.n84 VTAIL.n69 104.615
R164 VTAIL.n91 VTAIL.n69 104.615
R165 VTAIL.n93 VTAIL.n91 104.615
R166 VTAIL.n93 VTAIL.n92 104.615
R167 VTAIL.n92 VTAIL.n65 104.615
R168 VTAIL.n101 VTAIL.n65 104.615
R169 VTAIL.n102 VTAIL.n101 104.615
R170 VTAIL.n102 VTAIL.n61 104.615
R171 VTAIL.n109 VTAIL.n61 104.615
R172 VTAIL.n110 VTAIL.n109 104.615
R173 VTAIL.n134 VTAIL.n131 104.615
R174 VTAIL.n141 VTAIL.n131 104.615
R175 VTAIL.n142 VTAIL.n141 104.615
R176 VTAIL.n142 VTAIL.n127 104.615
R177 VTAIL.n149 VTAIL.n127 104.615
R178 VTAIL.n151 VTAIL.n149 104.615
R179 VTAIL.n151 VTAIL.n150 104.615
R180 VTAIL.n150 VTAIL.n123 104.615
R181 VTAIL.n159 VTAIL.n123 104.615
R182 VTAIL.n160 VTAIL.n159 104.615
R183 VTAIL.n160 VTAIL.n119 104.615
R184 VTAIL.n167 VTAIL.n119 104.615
R185 VTAIL.n168 VTAIL.n167 104.615
R186 VTAIL.n400 VTAIL.n399 104.615
R187 VTAIL.n399 VTAIL.n351 104.615
R188 VTAIL.n392 VTAIL.n351 104.615
R189 VTAIL.n392 VTAIL.n391 104.615
R190 VTAIL.n391 VTAIL.n355 104.615
R191 VTAIL.n359 VTAIL.n355 104.615
R192 VTAIL.n383 VTAIL.n359 104.615
R193 VTAIL.n383 VTAIL.n382 104.615
R194 VTAIL.n382 VTAIL.n360 104.615
R195 VTAIL.n375 VTAIL.n360 104.615
R196 VTAIL.n375 VTAIL.n374 104.615
R197 VTAIL.n374 VTAIL.n364 104.615
R198 VTAIL.n367 VTAIL.n364 104.615
R199 VTAIL.n342 VTAIL.n341 104.615
R200 VTAIL.n341 VTAIL.n293 104.615
R201 VTAIL.n334 VTAIL.n293 104.615
R202 VTAIL.n334 VTAIL.n333 104.615
R203 VTAIL.n333 VTAIL.n297 104.615
R204 VTAIL.n301 VTAIL.n297 104.615
R205 VTAIL.n325 VTAIL.n301 104.615
R206 VTAIL.n325 VTAIL.n324 104.615
R207 VTAIL.n324 VTAIL.n302 104.615
R208 VTAIL.n317 VTAIL.n302 104.615
R209 VTAIL.n317 VTAIL.n316 104.615
R210 VTAIL.n316 VTAIL.n306 104.615
R211 VTAIL.n309 VTAIL.n306 104.615
R212 VTAIL.n284 VTAIL.n283 104.615
R213 VTAIL.n283 VTAIL.n235 104.615
R214 VTAIL.n276 VTAIL.n235 104.615
R215 VTAIL.n276 VTAIL.n275 104.615
R216 VTAIL.n275 VTAIL.n239 104.615
R217 VTAIL.n243 VTAIL.n239 104.615
R218 VTAIL.n267 VTAIL.n243 104.615
R219 VTAIL.n267 VTAIL.n266 104.615
R220 VTAIL.n266 VTAIL.n244 104.615
R221 VTAIL.n259 VTAIL.n244 104.615
R222 VTAIL.n259 VTAIL.n258 104.615
R223 VTAIL.n258 VTAIL.n248 104.615
R224 VTAIL.n251 VTAIL.n248 104.615
R225 VTAIL.n226 VTAIL.n225 104.615
R226 VTAIL.n225 VTAIL.n177 104.615
R227 VTAIL.n218 VTAIL.n177 104.615
R228 VTAIL.n218 VTAIL.n217 104.615
R229 VTAIL.n217 VTAIL.n181 104.615
R230 VTAIL.n185 VTAIL.n181 104.615
R231 VTAIL.n209 VTAIL.n185 104.615
R232 VTAIL.n209 VTAIL.n208 104.615
R233 VTAIL.n208 VTAIL.n186 104.615
R234 VTAIL.n201 VTAIL.n186 104.615
R235 VTAIL.n201 VTAIL.n200 104.615
R236 VTAIL.n200 VTAIL.n190 104.615
R237 VTAIL.n193 VTAIL.n190 104.615
R238 VTAIL.n424 VTAIL.t1 52.3082
R239 VTAIL.n18 VTAIL.t3 52.3082
R240 VTAIL.n76 VTAIL.t5 52.3082
R241 VTAIL.n134 VTAIL.t6 52.3082
R242 VTAIL.n367 VTAIL.t7 52.3082
R243 VTAIL.n309 VTAIL.t4 52.3082
R244 VTAIL.n251 VTAIL.t0 52.3082
R245 VTAIL.n193 VTAIL.t2 52.3082
R246 VTAIL.n463 VTAIL.n462 30.6338
R247 VTAIL.n57 VTAIL.n56 30.6338
R248 VTAIL.n115 VTAIL.n114 30.6338
R249 VTAIL.n173 VTAIL.n172 30.6338
R250 VTAIL.n405 VTAIL.n404 30.6338
R251 VTAIL.n347 VTAIL.n346 30.6338
R252 VTAIL.n289 VTAIL.n288 30.6338
R253 VTAIL.n231 VTAIL.n230 30.6338
R254 VTAIL.n463 VTAIL.n405 24.8583
R255 VTAIL.n231 VTAIL.n173 24.8583
R256 VTAIL.n448 VTAIL.n447 13.1884
R257 VTAIL.n42 VTAIL.n41 13.1884
R258 VTAIL.n100 VTAIL.n99 13.1884
R259 VTAIL.n158 VTAIL.n157 13.1884
R260 VTAIL.n390 VTAIL.n389 13.1884
R261 VTAIL.n332 VTAIL.n331 13.1884
R262 VTAIL.n274 VTAIL.n273 13.1884
R263 VTAIL.n216 VTAIL.n215 13.1884
R264 VTAIL.n446 VTAIL.n414 12.8005
R265 VTAIL.n451 VTAIL.n412 12.8005
R266 VTAIL.n40 VTAIL.n8 12.8005
R267 VTAIL.n45 VTAIL.n6 12.8005
R268 VTAIL.n98 VTAIL.n66 12.8005
R269 VTAIL.n103 VTAIL.n64 12.8005
R270 VTAIL.n156 VTAIL.n124 12.8005
R271 VTAIL.n161 VTAIL.n122 12.8005
R272 VTAIL.n393 VTAIL.n354 12.8005
R273 VTAIL.n388 VTAIL.n356 12.8005
R274 VTAIL.n335 VTAIL.n296 12.8005
R275 VTAIL.n330 VTAIL.n298 12.8005
R276 VTAIL.n277 VTAIL.n238 12.8005
R277 VTAIL.n272 VTAIL.n240 12.8005
R278 VTAIL.n219 VTAIL.n180 12.8005
R279 VTAIL.n214 VTAIL.n182 12.8005
R280 VTAIL.n443 VTAIL.n442 12.0247
R281 VTAIL.n452 VTAIL.n410 12.0247
R282 VTAIL.n37 VTAIL.n36 12.0247
R283 VTAIL.n46 VTAIL.n4 12.0247
R284 VTAIL.n95 VTAIL.n94 12.0247
R285 VTAIL.n104 VTAIL.n62 12.0247
R286 VTAIL.n153 VTAIL.n152 12.0247
R287 VTAIL.n162 VTAIL.n120 12.0247
R288 VTAIL.n394 VTAIL.n352 12.0247
R289 VTAIL.n385 VTAIL.n384 12.0247
R290 VTAIL.n336 VTAIL.n294 12.0247
R291 VTAIL.n327 VTAIL.n326 12.0247
R292 VTAIL.n278 VTAIL.n236 12.0247
R293 VTAIL.n269 VTAIL.n268 12.0247
R294 VTAIL.n220 VTAIL.n178 12.0247
R295 VTAIL.n211 VTAIL.n210 12.0247
R296 VTAIL.n438 VTAIL.n416 11.249
R297 VTAIL.n456 VTAIL.n455 11.249
R298 VTAIL.n32 VTAIL.n10 11.249
R299 VTAIL.n50 VTAIL.n49 11.249
R300 VTAIL.n90 VTAIL.n68 11.249
R301 VTAIL.n108 VTAIL.n107 11.249
R302 VTAIL.n148 VTAIL.n126 11.249
R303 VTAIL.n166 VTAIL.n165 11.249
R304 VTAIL.n398 VTAIL.n397 11.249
R305 VTAIL.n381 VTAIL.n358 11.249
R306 VTAIL.n340 VTAIL.n339 11.249
R307 VTAIL.n323 VTAIL.n300 11.249
R308 VTAIL.n282 VTAIL.n281 11.249
R309 VTAIL.n265 VTAIL.n242 11.249
R310 VTAIL.n224 VTAIL.n223 11.249
R311 VTAIL.n207 VTAIL.n184 11.249
R312 VTAIL.n437 VTAIL.n418 10.4732
R313 VTAIL.n459 VTAIL.n408 10.4732
R314 VTAIL.n31 VTAIL.n12 10.4732
R315 VTAIL.n53 VTAIL.n2 10.4732
R316 VTAIL.n89 VTAIL.n70 10.4732
R317 VTAIL.n111 VTAIL.n60 10.4732
R318 VTAIL.n147 VTAIL.n128 10.4732
R319 VTAIL.n169 VTAIL.n118 10.4732
R320 VTAIL.n401 VTAIL.n350 10.4732
R321 VTAIL.n380 VTAIL.n361 10.4732
R322 VTAIL.n343 VTAIL.n292 10.4732
R323 VTAIL.n322 VTAIL.n303 10.4732
R324 VTAIL.n285 VTAIL.n234 10.4732
R325 VTAIL.n264 VTAIL.n245 10.4732
R326 VTAIL.n227 VTAIL.n176 10.4732
R327 VTAIL.n206 VTAIL.n187 10.4732
R328 VTAIL.n425 VTAIL.n423 10.2747
R329 VTAIL.n19 VTAIL.n17 10.2747
R330 VTAIL.n77 VTAIL.n75 10.2747
R331 VTAIL.n135 VTAIL.n133 10.2747
R332 VTAIL.n368 VTAIL.n366 10.2747
R333 VTAIL.n310 VTAIL.n308 10.2747
R334 VTAIL.n252 VTAIL.n250 10.2747
R335 VTAIL.n194 VTAIL.n192 10.2747
R336 VTAIL.n434 VTAIL.n433 9.69747
R337 VTAIL.n460 VTAIL.n406 9.69747
R338 VTAIL.n28 VTAIL.n27 9.69747
R339 VTAIL.n54 VTAIL.n0 9.69747
R340 VTAIL.n86 VTAIL.n85 9.69747
R341 VTAIL.n112 VTAIL.n58 9.69747
R342 VTAIL.n144 VTAIL.n143 9.69747
R343 VTAIL.n170 VTAIL.n116 9.69747
R344 VTAIL.n402 VTAIL.n348 9.69747
R345 VTAIL.n377 VTAIL.n376 9.69747
R346 VTAIL.n344 VTAIL.n290 9.69747
R347 VTAIL.n319 VTAIL.n318 9.69747
R348 VTAIL.n286 VTAIL.n232 9.69747
R349 VTAIL.n261 VTAIL.n260 9.69747
R350 VTAIL.n228 VTAIL.n174 9.69747
R351 VTAIL.n203 VTAIL.n202 9.69747
R352 VTAIL.n462 VTAIL.n461 9.45567
R353 VTAIL.n56 VTAIL.n55 9.45567
R354 VTAIL.n114 VTAIL.n113 9.45567
R355 VTAIL.n172 VTAIL.n171 9.45567
R356 VTAIL.n404 VTAIL.n403 9.45567
R357 VTAIL.n346 VTAIL.n345 9.45567
R358 VTAIL.n288 VTAIL.n287 9.45567
R359 VTAIL.n230 VTAIL.n229 9.45567
R360 VTAIL.n461 VTAIL.n460 9.3005
R361 VTAIL.n408 VTAIL.n407 9.3005
R362 VTAIL.n455 VTAIL.n454 9.3005
R363 VTAIL.n453 VTAIL.n452 9.3005
R364 VTAIL.n412 VTAIL.n411 9.3005
R365 VTAIL.n427 VTAIL.n426 9.3005
R366 VTAIL.n429 VTAIL.n428 9.3005
R367 VTAIL.n420 VTAIL.n419 9.3005
R368 VTAIL.n435 VTAIL.n434 9.3005
R369 VTAIL.n437 VTAIL.n436 9.3005
R370 VTAIL.n416 VTAIL.n415 9.3005
R371 VTAIL.n444 VTAIL.n443 9.3005
R372 VTAIL.n446 VTAIL.n445 9.3005
R373 VTAIL.n55 VTAIL.n54 9.3005
R374 VTAIL.n2 VTAIL.n1 9.3005
R375 VTAIL.n49 VTAIL.n48 9.3005
R376 VTAIL.n47 VTAIL.n46 9.3005
R377 VTAIL.n6 VTAIL.n5 9.3005
R378 VTAIL.n21 VTAIL.n20 9.3005
R379 VTAIL.n23 VTAIL.n22 9.3005
R380 VTAIL.n14 VTAIL.n13 9.3005
R381 VTAIL.n29 VTAIL.n28 9.3005
R382 VTAIL.n31 VTAIL.n30 9.3005
R383 VTAIL.n10 VTAIL.n9 9.3005
R384 VTAIL.n38 VTAIL.n37 9.3005
R385 VTAIL.n40 VTAIL.n39 9.3005
R386 VTAIL.n113 VTAIL.n112 9.3005
R387 VTAIL.n60 VTAIL.n59 9.3005
R388 VTAIL.n107 VTAIL.n106 9.3005
R389 VTAIL.n105 VTAIL.n104 9.3005
R390 VTAIL.n64 VTAIL.n63 9.3005
R391 VTAIL.n79 VTAIL.n78 9.3005
R392 VTAIL.n81 VTAIL.n80 9.3005
R393 VTAIL.n72 VTAIL.n71 9.3005
R394 VTAIL.n87 VTAIL.n86 9.3005
R395 VTAIL.n89 VTAIL.n88 9.3005
R396 VTAIL.n68 VTAIL.n67 9.3005
R397 VTAIL.n96 VTAIL.n95 9.3005
R398 VTAIL.n98 VTAIL.n97 9.3005
R399 VTAIL.n171 VTAIL.n170 9.3005
R400 VTAIL.n118 VTAIL.n117 9.3005
R401 VTAIL.n165 VTAIL.n164 9.3005
R402 VTAIL.n163 VTAIL.n162 9.3005
R403 VTAIL.n122 VTAIL.n121 9.3005
R404 VTAIL.n137 VTAIL.n136 9.3005
R405 VTAIL.n139 VTAIL.n138 9.3005
R406 VTAIL.n130 VTAIL.n129 9.3005
R407 VTAIL.n145 VTAIL.n144 9.3005
R408 VTAIL.n147 VTAIL.n146 9.3005
R409 VTAIL.n126 VTAIL.n125 9.3005
R410 VTAIL.n154 VTAIL.n153 9.3005
R411 VTAIL.n156 VTAIL.n155 9.3005
R412 VTAIL.n370 VTAIL.n369 9.3005
R413 VTAIL.n372 VTAIL.n371 9.3005
R414 VTAIL.n363 VTAIL.n362 9.3005
R415 VTAIL.n378 VTAIL.n377 9.3005
R416 VTAIL.n380 VTAIL.n379 9.3005
R417 VTAIL.n358 VTAIL.n357 9.3005
R418 VTAIL.n386 VTAIL.n385 9.3005
R419 VTAIL.n388 VTAIL.n387 9.3005
R420 VTAIL.n403 VTAIL.n402 9.3005
R421 VTAIL.n350 VTAIL.n349 9.3005
R422 VTAIL.n397 VTAIL.n396 9.3005
R423 VTAIL.n395 VTAIL.n394 9.3005
R424 VTAIL.n354 VTAIL.n353 9.3005
R425 VTAIL.n312 VTAIL.n311 9.3005
R426 VTAIL.n314 VTAIL.n313 9.3005
R427 VTAIL.n305 VTAIL.n304 9.3005
R428 VTAIL.n320 VTAIL.n319 9.3005
R429 VTAIL.n322 VTAIL.n321 9.3005
R430 VTAIL.n300 VTAIL.n299 9.3005
R431 VTAIL.n328 VTAIL.n327 9.3005
R432 VTAIL.n330 VTAIL.n329 9.3005
R433 VTAIL.n345 VTAIL.n344 9.3005
R434 VTAIL.n292 VTAIL.n291 9.3005
R435 VTAIL.n339 VTAIL.n338 9.3005
R436 VTAIL.n337 VTAIL.n336 9.3005
R437 VTAIL.n296 VTAIL.n295 9.3005
R438 VTAIL.n254 VTAIL.n253 9.3005
R439 VTAIL.n256 VTAIL.n255 9.3005
R440 VTAIL.n247 VTAIL.n246 9.3005
R441 VTAIL.n262 VTAIL.n261 9.3005
R442 VTAIL.n264 VTAIL.n263 9.3005
R443 VTAIL.n242 VTAIL.n241 9.3005
R444 VTAIL.n270 VTAIL.n269 9.3005
R445 VTAIL.n272 VTAIL.n271 9.3005
R446 VTAIL.n287 VTAIL.n286 9.3005
R447 VTAIL.n234 VTAIL.n233 9.3005
R448 VTAIL.n281 VTAIL.n280 9.3005
R449 VTAIL.n279 VTAIL.n278 9.3005
R450 VTAIL.n238 VTAIL.n237 9.3005
R451 VTAIL.n196 VTAIL.n195 9.3005
R452 VTAIL.n198 VTAIL.n197 9.3005
R453 VTAIL.n189 VTAIL.n188 9.3005
R454 VTAIL.n204 VTAIL.n203 9.3005
R455 VTAIL.n206 VTAIL.n205 9.3005
R456 VTAIL.n184 VTAIL.n183 9.3005
R457 VTAIL.n212 VTAIL.n211 9.3005
R458 VTAIL.n214 VTAIL.n213 9.3005
R459 VTAIL.n229 VTAIL.n228 9.3005
R460 VTAIL.n176 VTAIL.n175 9.3005
R461 VTAIL.n223 VTAIL.n222 9.3005
R462 VTAIL.n221 VTAIL.n220 9.3005
R463 VTAIL.n180 VTAIL.n179 9.3005
R464 VTAIL.n430 VTAIL.n420 8.92171
R465 VTAIL.n24 VTAIL.n14 8.92171
R466 VTAIL.n82 VTAIL.n72 8.92171
R467 VTAIL.n140 VTAIL.n130 8.92171
R468 VTAIL.n373 VTAIL.n363 8.92171
R469 VTAIL.n315 VTAIL.n305 8.92171
R470 VTAIL.n257 VTAIL.n247 8.92171
R471 VTAIL.n199 VTAIL.n189 8.92171
R472 VTAIL.n429 VTAIL.n422 8.14595
R473 VTAIL.n23 VTAIL.n16 8.14595
R474 VTAIL.n81 VTAIL.n74 8.14595
R475 VTAIL.n139 VTAIL.n132 8.14595
R476 VTAIL.n372 VTAIL.n365 8.14595
R477 VTAIL.n314 VTAIL.n307 8.14595
R478 VTAIL.n256 VTAIL.n249 8.14595
R479 VTAIL.n198 VTAIL.n191 8.14595
R480 VTAIL.n426 VTAIL.n425 7.3702
R481 VTAIL.n20 VTAIL.n19 7.3702
R482 VTAIL.n78 VTAIL.n77 7.3702
R483 VTAIL.n136 VTAIL.n135 7.3702
R484 VTAIL.n369 VTAIL.n368 7.3702
R485 VTAIL.n311 VTAIL.n310 7.3702
R486 VTAIL.n253 VTAIL.n252 7.3702
R487 VTAIL.n195 VTAIL.n194 7.3702
R488 VTAIL.n426 VTAIL.n422 5.81868
R489 VTAIL.n20 VTAIL.n16 5.81868
R490 VTAIL.n78 VTAIL.n74 5.81868
R491 VTAIL.n136 VTAIL.n132 5.81868
R492 VTAIL.n369 VTAIL.n365 5.81868
R493 VTAIL.n311 VTAIL.n307 5.81868
R494 VTAIL.n253 VTAIL.n249 5.81868
R495 VTAIL.n195 VTAIL.n191 5.81868
R496 VTAIL.n430 VTAIL.n429 5.04292
R497 VTAIL.n24 VTAIL.n23 5.04292
R498 VTAIL.n82 VTAIL.n81 5.04292
R499 VTAIL.n140 VTAIL.n139 5.04292
R500 VTAIL.n373 VTAIL.n372 5.04292
R501 VTAIL.n315 VTAIL.n314 5.04292
R502 VTAIL.n257 VTAIL.n256 5.04292
R503 VTAIL.n199 VTAIL.n198 5.04292
R504 VTAIL.n433 VTAIL.n420 4.26717
R505 VTAIL.n462 VTAIL.n406 4.26717
R506 VTAIL.n27 VTAIL.n14 4.26717
R507 VTAIL.n56 VTAIL.n0 4.26717
R508 VTAIL.n85 VTAIL.n72 4.26717
R509 VTAIL.n114 VTAIL.n58 4.26717
R510 VTAIL.n143 VTAIL.n130 4.26717
R511 VTAIL.n172 VTAIL.n116 4.26717
R512 VTAIL.n404 VTAIL.n348 4.26717
R513 VTAIL.n376 VTAIL.n363 4.26717
R514 VTAIL.n346 VTAIL.n290 4.26717
R515 VTAIL.n318 VTAIL.n305 4.26717
R516 VTAIL.n288 VTAIL.n232 4.26717
R517 VTAIL.n260 VTAIL.n247 4.26717
R518 VTAIL.n230 VTAIL.n174 4.26717
R519 VTAIL.n202 VTAIL.n189 4.26717
R520 VTAIL.n434 VTAIL.n418 3.49141
R521 VTAIL.n460 VTAIL.n459 3.49141
R522 VTAIL.n28 VTAIL.n12 3.49141
R523 VTAIL.n54 VTAIL.n53 3.49141
R524 VTAIL.n86 VTAIL.n70 3.49141
R525 VTAIL.n112 VTAIL.n111 3.49141
R526 VTAIL.n144 VTAIL.n128 3.49141
R527 VTAIL.n170 VTAIL.n169 3.49141
R528 VTAIL.n402 VTAIL.n401 3.49141
R529 VTAIL.n377 VTAIL.n361 3.49141
R530 VTAIL.n344 VTAIL.n343 3.49141
R531 VTAIL.n319 VTAIL.n303 3.49141
R532 VTAIL.n286 VTAIL.n285 3.49141
R533 VTAIL.n261 VTAIL.n245 3.49141
R534 VTAIL.n228 VTAIL.n227 3.49141
R535 VTAIL.n203 VTAIL.n187 3.49141
R536 VTAIL.n289 VTAIL.n231 3.35395
R537 VTAIL.n405 VTAIL.n347 3.35395
R538 VTAIL.n173 VTAIL.n115 3.35395
R539 VTAIL.n427 VTAIL.n423 2.84303
R540 VTAIL.n21 VTAIL.n17 2.84303
R541 VTAIL.n79 VTAIL.n75 2.84303
R542 VTAIL.n137 VTAIL.n133 2.84303
R543 VTAIL.n370 VTAIL.n366 2.84303
R544 VTAIL.n312 VTAIL.n308 2.84303
R545 VTAIL.n254 VTAIL.n250 2.84303
R546 VTAIL.n196 VTAIL.n192 2.84303
R547 VTAIL.n438 VTAIL.n437 2.71565
R548 VTAIL.n456 VTAIL.n408 2.71565
R549 VTAIL.n32 VTAIL.n31 2.71565
R550 VTAIL.n50 VTAIL.n2 2.71565
R551 VTAIL.n90 VTAIL.n89 2.71565
R552 VTAIL.n108 VTAIL.n60 2.71565
R553 VTAIL.n148 VTAIL.n147 2.71565
R554 VTAIL.n166 VTAIL.n118 2.71565
R555 VTAIL.n398 VTAIL.n350 2.71565
R556 VTAIL.n381 VTAIL.n380 2.71565
R557 VTAIL.n340 VTAIL.n292 2.71565
R558 VTAIL.n323 VTAIL.n322 2.71565
R559 VTAIL.n282 VTAIL.n234 2.71565
R560 VTAIL.n265 VTAIL.n264 2.71565
R561 VTAIL.n224 VTAIL.n176 2.71565
R562 VTAIL.n207 VTAIL.n206 2.71565
R563 VTAIL.n442 VTAIL.n416 1.93989
R564 VTAIL.n455 VTAIL.n410 1.93989
R565 VTAIL.n36 VTAIL.n10 1.93989
R566 VTAIL.n49 VTAIL.n4 1.93989
R567 VTAIL.n94 VTAIL.n68 1.93989
R568 VTAIL.n107 VTAIL.n62 1.93989
R569 VTAIL.n152 VTAIL.n126 1.93989
R570 VTAIL.n165 VTAIL.n120 1.93989
R571 VTAIL.n397 VTAIL.n352 1.93989
R572 VTAIL.n384 VTAIL.n358 1.93989
R573 VTAIL.n339 VTAIL.n294 1.93989
R574 VTAIL.n326 VTAIL.n300 1.93989
R575 VTAIL.n281 VTAIL.n236 1.93989
R576 VTAIL.n268 VTAIL.n242 1.93989
R577 VTAIL.n223 VTAIL.n178 1.93989
R578 VTAIL.n210 VTAIL.n184 1.93989
R579 VTAIL VTAIL.n57 1.73541
R580 VTAIL VTAIL.n463 1.61903
R581 VTAIL.n443 VTAIL.n414 1.16414
R582 VTAIL.n452 VTAIL.n451 1.16414
R583 VTAIL.n37 VTAIL.n8 1.16414
R584 VTAIL.n46 VTAIL.n45 1.16414
R585 VTAIL.n95 VTAIL.n66 1.16414
R586 VTAIL.n104 VTAIL.n103 1.16414
R587 VTAIL.n153 VTAIL.n124 1.16414
R588 VTAIL.n162 VTAIL.n161 1.16414
R589 VTAIL.n394 VTAIL.n393 1.16414
R590 VTAIL.n385 VTAIL.n356 1.16414
R591 VTAIL.n336 VTAIL.n335 1.16414
R592 VTAIL.n327 VTAIL.n298 1.16414
R593 VTAIL.n278 VTAIL.n277 1.16414
R594 VTAIL.n269 VTAIL.n240 1.16414
R595 VTAIL.n220 VTAIL.n219 1.16414
R596 VTAIL.n211 VTAIL.n182 1.16414
R597 VTAIL.n347 VTAIL.n289 0.470328
R598 VTAIL.n115 VTAIL.n57 0.470328
R599 VTAIL.n447 VTAIL.n446 0.388379
R600 VTAIL.n448 VTAIL.n412 0.388379
R601 VTAIL.n41 VTAIL.n40 0.388379
R602 VTAIL.n42 VTAIL.n6 0.388379
R603 VTAIL.n99 VTAIL.n98 0.388379
R604 VTAIL.n100 VTAIL.n64 0.388379
R605 VTAIL.n157 VTAIL.n156 0.388379
R606 VTAIL.n158 VTAIL.n122 0.388379
R607 VTAIL.n390 VTAIL.n354 0.388379
R608 VTAIL.n389 VTAIL.n388 0.388379
R609 VTAIL.n332 VTAIL.n296 0.388379
R610 VTAIL.n331 VTAIL.n330 0.388379
R611 VTAIL.n274 VTAIL.n238 0.388379
R612 VTAIL.n273 VTAIL.n272 0.388379
R613 VTAIL.n216 VTAIL.n180 0.388379
R614 VTAIL.n215 VTAIL.n214 0.388379
R615 VTAIL.n428 VTAIL.n427 0.155672
R616 VTAIL.n428 VTAIL.n419 0.155672
R617 VTAIL.n435 VTAIL.n419 0.155672
R618 VTAIL.n436 VTAIL.n435 0.155672
R619 VTAIL.n436 VTAIL.n415 0.155672
R620 VTAIL.n444 VTAIL.n415 0.155672
R621 VTAIL.n445 VTAIL.n444 0.155672
R622 VTAIL.n445 VTAIL.n411 0.155672
R623 VTAIL.n453 VTAIL.n411 0.155672
R624 VTAIL.n454 VTAIL.n453 0.155672
R625 VTAIL.n454 VTAIL.n407 0.155672
R626 VTAIL.n461 VTAIL.n407 0.155672
R627 VTAIL.n22 VTAIL.n21 0.155672
R628 VTAIL.n22 VTAIL.n13 0.155672
R629 VTAIL.n29 VTAIL.n13 0.155672
R630 VTAIL.n30 VTAIL.n29 0.155672
R631 VTAIL.n30 VTAIL.n9 0.155672
R632 VTAIL.n38 VTAIL.n9 0.155672
R633 VTAIL.n39 VTAIL.n38 0.155672
R634 VTAIL.n39 VTAIL.n5 0.155672
R635 VTAIL.n47 VTAIL.n5 0.155672
R636 VTAIL.n48 VTAIL.n47 0.155672
R637 VTAIL.n48 VTAIL.n1 0.155672
R638 VTAIL.n55 VTAIL.n1 0.155672
R639 VTAIL.n80 VTAIL.n79 0.155672
R640 VTAIL.n80 VTAIL.n71 0.155672
R641 VTAIL.n87 VTAIL.n71 0.155672
R642 VTAIL.n88 VTAIL.n87 0.155672
R643 VTAIL.n88 VTAIL.n67 0.155672
R644 VTAIL.n96 VTAIL.n67 0.155672
R645 VTAIL.n97 VTAIL.n96 0.155672
R646 VTAIL.n97 VTAIL.n63 0.155672
R647 VTAIL.n105 VTAIL.n63 0.155672
R648 VTAIL.n106 VTAIL.n105 0.155672
R649 VTAIL.n106 VTAIL.n59 0.155672
R650 VTAIL.n113 VTAIL.n59 0.155672
R651 VTAIL.n138 VTAIL.n137 0.155672
R652 VTAIL.n138 VTAIL.n129 0.155672
R653 VTAIL.n145 VTAIL.n129 0.155672
R654 VTAIL.n146 VTAIL.n145 0.155672
R655 VTAIL.n146 VTAIL.n125 0.155672
R656 VTAIL.n154 VTAIL.n125 0.155672
R657 VTAIL.n155 VTAIL.n154 0.155672
R658 VTAIL.n155 VTAIL.n121 0.155672
R659 VTAIL.n163 VTAIL.n121 0.155672
R660 VTAIL.n164 VTAIL.n163 0.155672
R661 VTAIL.n164 VTAIL.n117 0.155672
R662 VTAIL.n171 VTAIL.n117 0.155672
R663 VTAIL.n403 VTAIL.n349 0.155672
R664 VTAIL.n396 VTAIL.n349 0.155672
R665 VTAIL.n396 VTAIL.n395 0.155672
R666 VTAIL.n395 VTAIL.n353 0.155672
R667 VTAIL.n387 VTAIL.n353 0.155672
R668 VTAIL.n387 VTAIL.n386 0.155672
R669 VTAIL.n386 VTAIL.n357 0.155672
R670 VTAIL.n379 VTAIL.n357 0.155672
R671 VTAIL.n379 VTAIL.n378 0.155672
R672 VTAIL.n378 VTAIL.n362 0.155672
R673 VTAIL.n371 VTAIL.n362 0.155672
R674 VTAIL.n371 VTAIL.n370 0.155672
R675 VTAIL.n345 VTAIL.n291 0.155672
R676 VTAIL.n338 VTAIL.n291 0.155672
R677 VTAIL.n338 VTAIL.n337 0.155672
R678 VTAIL.n337 VTAIL.n295 0.155672
R679 VTAIL.n329 VTAIL.n295 0.155672
R680 VTAIL.n329 VTAIL.n328 0.155672
R681 VTAIL.n328 VTAIL.n299 0.155672
R682 VTAIL.n321 VTAIL.n299 0.155672
R683 VTAIL.n321 VTAIL.n320 0.155672
R684 VTAIL.n320 VTAIL.n304 0.155672
R685 VTAIL.n313 VTAIL.n304 0.155672
R686 VTAIL.n313 VTAIL.n312 0.155672
R687 VTAIL.n287 VTAIL.n233 0.155672
R688 VTAIL.n280 VTAIL.n233 0.155672
R689 VTAIL.n280 VTAIL.n279 0.155672
R690 VTAIL.n279 VTAIL.n237 0.155672
R691 VTAIL.n271 VTAIL.n237 0.155672
R692 VTAIL.n271 VTAIL.n270 0.155672
R693 VTAIL.n270 VTAIL.n241 0.155672
R694 VTAIL.n263 VTAIL.n241 0.155672
R695 VTAIL.n263 VTAIL.n262 0.155672
R696 VTAIL.n262 VTAIL.n246 0.155672
R697 VTAIL.n255 VTAIL.n246 0.155672
R698 VTAIL.n255 VTAIL.n254 0.155672
R699 VTAIL.n229 VTAIL.n175 0.155672
R700 VTAIL.n222 VTAIL.n175 0.155672
R701 VTAIL.n222 VTAIL.n221 0.155672
R702 VTAIL.n221 VTAIL.n179 0.155672
R703 VTAIL.n213 VTAIL.n179 0.155672
R704 VTAIL.n213 VTAIL.n212 0.155672
R705 VTAIL.n212 VTAIL.n183 0.155672
R706 VTAIL.n205 VTAIL.n183 0.155672
R707 VTAIL.n205 VTAIL.n204 0.155672
R708 VTAIL.n204 VTAIL.n188 0.155672
R709 VTAIL.n197 VTAIL.n188 0.155672
R710 VTAIL.n197 VTAIL.n196 0.155672
R711 VDD2.n2 VDD2.n0 103.701
R712 VDD2.n2 VDD2.n1 60.7886
R713 VDD2.n1 VDD2.t2 1.86842
R714 VDD2.n1 VDD2.t1 1.86842
R715 VDD2.n0 VDD2.t0 1.86842
R716 VDD2.n0 VDD2.t3 1.86842
R717 VDD2 VDD2.n2 0.0586897
R718 B.n609 B.n608 585
R719 B.n609 B.n79 585
R720 B.n612 B.n611 585
R721 B.n613 B.n126 585
R722 B.n615 B.n614 585
R723 B.n617 B.n125 585
R724 B.n620 B.n619 585
R725 B.n621 B.n124 585
R726 B.n623 B.n622 585
R727 B.n625 B.n123 585
R728 B.n628 B.n627 585
R729 B.n629 B.n122 585
R730 B.n631 B.n630 585
R731 B.n633 B.n121 585
R732 B.n636 B.n635 585
R733 B.n637 B.n120 585
R734 B.n639 B.n638 585
R735 B.n641 B.n119 585
R736 B.n644 B.n643 585
R737 B.n645 B.n118 585
R738 B.n647 B.n646 585
R739 B.n649 B.n117 585
R740 B.n652 B.n651 585
R741 B.n653 B.n116 585
R742 B.n655 B.n654 585
R743 B.n657 B.n115 585
R744 B.n660 B.n659 585
R745 B.n661 B.n114 585
R746 B.n663 B.n662 585
R747 B.n665 B.n113 585
R748 B.n668 B.n667 585
R749 B.n669 B.n112 585
R750 B.n671 B.n670 585
R751 B.n673 B.n111 585
R752 B.n676 B.n675 585
R753 B.n677 B.n110 585
R754 B.n679 B.n678 585
R755 B.n681 B.n109 585
R756 B.n684 B.n683 585
R757 B.n686 B.n106 585
R758 B.n688 B.n687 585
R759 B.n690 B.n105 585
R760 B.n693 B.n692 585
R761 B.n694 B.n104 585
R762 B.n696 B.n695 585
R763 B.n698 B.n103 585
R764 B.n700 B.n699 585
R765 B.n702 B.n701 585
R766 B.n705 B.n704 585
R767 B.n706 B.n98 585
R768 B.n708 B.n707 585
R769 B.n710 B.n97 585
R770 B.n713 B.n712 585
R771 B.n714 B.n96 585
R772 B.n716 B.n715 585
R773 B.n718 B.n95 585
R774 B.n721 B.n720 585
R775 B.n722 B.n94 585
R776 B.n724 B.n723 585
R777 B.n726 B.n93 585
R778 B.n729 B.n728 585
R779 B.n730 B.n92 585
R780 B.n732 B.n731 585
R781 B.n734 B.n91 585
R782 B.n737 B.n736 585
R783 B.n738 B.n90 585
R784 B.n740 B.n739 585
R785 B.n742 B.n89 585
R786 B.n745 B.n744 585
R787 B.n746 B.n88 585
R788 B.n748 B.n747 585
R789 B.n750 B.n87 585
R790 B.n753 B.n752 585
R791 B.n754 B.n86 585
R792 B.n756 B.n755 585
R793 B.n758 B.n85 585
R794 B.n761 B.n760 585
R795 B.n762 B.n84 585
R796 B.n764 B.n763 585
R797 B.n766 B.n83 585
R798 B.n769 B.n768 585
R799 B.n770 B.n82 585
R800 B.n772 B.n771 585
R801 B.n774 B.n81 585
R802 B.n777 B.n776 585
R803 B.n778 B.n80 585
R804 B.n607 B.n78 585
R805 B.n781 B.n78 585
R806 B.n606 B.n77 585
R807 B.n782 B.n77 585
R808 B.n605 B.n76 585
R809 B.n783 B.n76 585
R810 B.n604 B.n603 585
R811 B.n603 B.n72 585
R812 B.n602 B.n71 585
R813 B.n789 B.n71 585
R814 B.n601 B.n70 585
R815 B.n790 B.n70 585
R816 B.n600 B.n69 585
R817 B.n791 B.n69 585
R818 B.n599 B.n598 585
R819 B.n598 B.n65 585
R820 B.n597 B.n64 585
R821 B.n797 B.n64 585
R822 B.n596 B.n63 585
R823 B.n798 B.n63 585
R824 B.n595 B.n62 585
R825 B.n799 B.n62 585
R826 B.n594 B.n593 585
R827 B.n593 B.n58 585
R828 B.n592 B.n57 585
R829 B.n805 B.n57 585
R830 B.n591 B.n56 585
R831 B.n806 B.n56 585
R832 B.n590 B.n55 585
R833 B.n807 B.n55 585
R834 B.n589 B.n588 585
R835 B.n588 B.n51 585
R836 B.n587 B.n50 585
R837 B.n813 B.n50 585
R838 B.n586 B.n49 585
R839 B.n814 B.n49 585
R840 B.n585 B.n48 585
R841 B.n815 B.n48 585
R842 B.n584 B.n583 585
R843 B.n583 B.n44 585
R844 B.n582 B.n43 585
R845 B.n821 B.n43 585
R846 B.n581 B.n42 585
R847 B.n822 B.n42 585
R848 B.n580 B.n41 585
R849 B.n823 B.n41 585
R850 B.n579 B.n578 585
R851 B.n578 B.n40 585
R852 B.n577 B.n36 585
R853 B.n829 B.n36 585
R854 B.n576 B.n35 585
R855 B.n830 B.n35 585
R856 B.n575 B.n34 585
R857 B.n831 B.n34 585
R858 B.n574 B.n573 585
R859 B.n573 B.n30 585
R860 B.n572 B.n29 585
R861 B.n837 B.n29 585
R862 B.n571 B.n28 585
R863 B.n838 B.n28 585
R864 B.n570 B.n27 585
R865 B.n839 B.n27 585
R866 B.n569 B.n568 585
R867 B.n568 B.n23 585
R868 B.n567 B.n22 585
R869 B.n845 B.n22 585
R870 B.n566 B.n21 585
R871 B.n846 B.n21 585
R872 B.n565 B.n20 585
R873 B.n847 B.n20 585
R874 B.n564 B.n563 585
R875 B.n563 B.n19 585
R876 B.n562 B.n15 585
R877 B.n853 B.n15 585
R878 B.n561 B.n14 585
R879 B.n854 B.n14 585
R880 B.n560 B.n13 585
R881 B.n855 B.n13 585
R882 B.n559 B.n558 585
R883 B.n558 B.n12 585
R884 B.n557 B.n556 585
R885 B.n557 B.n8 585
R886 B.n555 B.n7 585
R887 B.n862 B.n7 585
R888 B.n554 B.n6 585
R889 B.n863 B.n6 585
R890 B.n553 B.n5 585
R891 B.n864 B.n5 585
R892 B.n552 B.n551 585
R893 B.n551 B.n4 585
R894 B.n550 B.n127 585
R895 B.n550 B.n549 585
R896 B.n540 B.n128 585
R897 B.n129 B.n128 585
R898 B.n542 B.n541 585
R899 B.n543 B.n542 585
R900 B.n539 B.n134 585
R901 B.n134 B.n133 585
R902 B.n538 B.n537 585
R903 B.n537 B.n536 585
R904 B.n136 B.n135 585
R905 B.n529 B.n136 585
R906 B.n528 B.n527 585
R907 B.n530 B.n528 585
R908 B.n526 B.n141 585
R909 B.n141 B.n140 585
R910 B.n525 B.n524 585
R911 B.n524 B.n523 585
R912 B.n143 B.n142 585
R913 B.n144 B.n143 585
R914 B.n516 B.n515 585
R915 B.n517 B.n516 585
R916 B.n514 B.n149 585
R917 B.n149 B.n148 585
R918 B.n513 B.n512 585
R919 B.n512 B.n511 585
R920 B.n151 B.n150 585
R921 B.n152 B.n151 585
R922 B.n504 B.n503 585
R923 B.n505 B.n504 585
R924 B.n502 B.n157 585
R925 B.n157 B.n156 585
R926 B.n501 B.n500 585
R927 B.n500 B.n499 585
R928 B.n159 B.n158 585
R929 B.n492 B.n159 585
R930 B.n491 B.n490 585
R931 B.n493 B.n491 585
R932 B.n489 B.n164 585
R933 B.n164 B.n163 585
R934 B.n488 B.n487 585
R935 B.n487 B.n486 585
R936 B.n166 B.n165 585
R937 B.n167 B.n166 585
R938 B.n479 B.n478 585
R939 B.n480 B.n479 585
R940 B.n477 B.n172 585
R941 B.n172 B.n171 585
R942 B.n476 B.n475 585
R943 B.n475 B.n474 585
R944 B.n174 B.n173 585
R945 B.n175 B.n174 585
R946 B.n467 B.n466 585
R947 B.n468 B.n467 585
R948 B.n465 B.n180 585
R949 B.n180 B.n179 585
R950 B.n464 B.n463 585
R951 B.n463 B.n462 585
R952 B.n182 B.n181 585
R953 B.n183 B.n182 585
R954 B.n455 B.n454 585
R955 B.n456 B.n455 585
R956 B.n453 B.n187 585
R957 B.n191 B.n187 585
R958 B.n452 B.n451 585
R959 B.n451 B.n450 585
R960 B.n189 B.n188 585
R961 B.n190 B.n189 585
R962 B.n443 B.n442 585
R963 B.n444 B.n443 585
R964 B.n441 B.n196 585
R965 B.n196 B.n195 585
R966 B.n440 B.n439 585
R967 B.n439 B.n438 585
R968 B.n198 B.n197 585
R969 B.n199 B.n198 585
R970 B.n431 B.n430 585
R971 B.n432 B.n431 585
R972 B.n429 B.n204 585
R973 B.n204 B.n203 585
R974 B.n428 B.n427 585
R975 B.n427 B.n426 585
R976 B.n423 B.n208 585
R977 B.n422 B.n421 585
R978 B.n419 B.n209 585
R979 B.n419 B.n207 585
R980 B.n418 B.n417 585
R981 B.n416 B.n415 585
R982 B.n414 B.n211 585
R983 B.n412 B.n411 585
R984 B.n410 B.n212 585
R985 B.n409 B.n408 585
R986 B.n406 B.n213 585
R987 B.n404 B.n403 585
R988 B.n402 B.n214 585
R989 B.n401 B.n400 585
R990 B.n398 B.n215 585
R991 B.n396 B.n395 585
R992 B.n394 B.n216 585
R993 B.n393 B.n392 585
R994 B.n390 B.n217 585
R995 B.n388 B.n387 585
R996 B.n386 B.n218 585
R997 B.n385 B.n384 585
R998 B.n382 B.n219 585
R999 B.n380 B.n379 585
R1000 B.n378 B.n220 585
R1001 B.n377 B.n376 585
R1002 B.n374 B.n221 585
R1003 B.n372 B.n371 585
R1004 B.n370 B.n222 585
R1005 B.n369 B.n368 585
R1006 B.n366 B.n223 585
R1007 B.n364 B.n363 585
R1008 B.n362 B.n224 585
R1009 B.n361 B.n360 585
R1010 B.n358 B.n225 585
R1011 B.n356 B.n355 585
R1012 B.n354 B.n226 585
R1013 B.n353 B.n352 585
R1014 B.n350 B.n227 585
R1015 B.n348 B.n347 585
R1016 B.n346 B.n228 585
R1017 B.n345 B.n344 585
R1018 B.n342 B.n232 585
R1019 B.n340 B.n339 585
R1020 B.n338 B.n233 585
R1021 B.n337 B.n336 585
R1022 B.n334 B.n234 585
R1023 B.n332 B.n331 585
R1024 B.n329 B.n235 585
R1025 B.n328 B.n327 585
R1026 B.n325 B.n238 585
R1027 B.n323 B.n322 585
R1028 B.n321 B.n239 585
R1029 B.n320 B.n319 585
R1030 B.n317 B.n240 585
R1031 B.n315 B.n314 585
R1032 B.n313 B.n241 585
R1033 B.n312 B.n311 585
R1034 B.n309 B.n242 585
R1035 B.n307 B.n306 585
R1036 B.n305 B.n243 585
R1037 B.n304 B.n303 585
R1038 B.n301 B.n244 585
R1039 B.n299 B.n298 585
R1040 B.n297 B.n245 585
R1041 B.n296 B.n295 585
R1042 B.n293 B.n246 585
R1043 B.n291 B.n290 585
R1044 B.n289 B.n247 585
R1045 B.n288 B.n287 585
R1046 B.n285 B.n248 585
R1047 B.n283 B.n282 585
R1048 B.n281 B.n249 585
R1049 B.n280 B.n279 585
R1050 B.n277 B.n250 585
R1051 B.n275 B.n274 585
R1052 B.n273 B.n251 585
R1053 B.n272 B.n271 585
R1054 B.n269 B.n252 585
R1055 B.n267 B.n266 585
R1056 B.n265 B.n253 585
R1057 B.n264 B.n263 585
R1058 B.n261 B.n254 585
R1059 B.n259 B.n258 585
R1060 B.n257 B.n256 585
R1061 B.n206 B.n205 585
R1062 B.n425 B.n424 585
R1063 B.n426 B.n425 585
R1064 B.n202 B.n201 585
R1065 B.n203 B.n202 585
R1066 B.n434 B.n433 585
R1067 B.n433 B.n432 585
R1068 B.n435 B.n200 585
R1069 B.n200 B.n199 585
R1070 B.n437 B.n436 585
R1071 B.n438 B.n437 585
R1072 B.n194 B.n193 585
R1073 B.n195 B.n194 585
R1074 B.n446 B.n445 585
R1075 B.n445 B.n444 585
R1076 B.n447 B.n192 585
R1077 B.n192 B.n190 585
R1078 B.n449 B.n448 585
R1079 B.n450 B.n449 585
R1080 B.n186 B.n185 585
R1081 B.n191 B.n186 585
R1082 B.n458 B.n457 585
R1083 B.n457 B.n456 585
R1084 B.n459 B.n184 585
R1085 B.n184 B.n183 585
R1086 B.n461 B.n460 585
R1087 B.n462 B.n461 585
R1088 B.n178 B.n177 585
R1089 B.n179 B.n178 585
R1090 B.n470 B.n469 585
R1091 B.n469 B.n468 585
R1092 B.n471 B.n176 585
R1093 B.n176 B.n175 585
R1094 B.n473 B.n472 585
R1095 B.n474 B.n473 585
R1096 B.n170 B.n169 585
R1097 B.n171 B.n170 585
R1098 B.n482 B.n481 585
R1099 B.n481 B.n480 585
R1100 B.n483 B.n168 585
R1101 B.n168 B.n167 585
R1102 B.n485 B.n484 585
R1103 B.n486 B.n485 585
R1104 B.n162 B.n161 585
R1105 B.n163 B.n162 585
R1106 B.n495 B.n494 585
R1107 B.n494 B.n493 585
R1108 B.n496 B.n160 585
R1109 B.n492 B.n160 585
R1110 B.n498 B.n497 585
R1111 B.n499 B.n498 585
R1112 B.n155 B.n154 585
R1113 B.n156 B.n155 585
R1114 B.n507 B.n506 585
R1115 B.n506 B.n505 585
R1116 B.n508 B.n153 585
R1117 B.n153 B.n152 585
R1118 B.n510 B.n509 585
R1119 B.n511 B.n510 585
R1120 B.n147 B.n146 585
R1121 B.n148 B.n147 585
R1122 B.n519 B.n518 585
R1123 B.n518 B.n517 585
R1124 B.n520 B.n145 585
R1125 B.n145 B.n144 585
R1126 B.n522 B.n521 585
R1127 B.n523 B.n522 585
R1128 B.n139 B.n138 585
R1129 B.n140 B.n139 585
R1130 B.n532 B.n531 585
R1131 B.n531 B.n530 585
R1132 B.n533 B.n137 585
R1133 B.n529 B.n137 585
R1134 B.n535 B.n534 585
R1135 B.n536 B.n535 585
R1136 B.n132 B.n131 585
R1137 B.n133 B.n132 585
R1138 B.n545 B.n544 585
R1139 B.n544 B.n543 585
R1140 B.n546 B.n130 585
R1141 B.n130 B.n129 585
R1142 B.n548 B.n547 585
R1143 B.n549 B.n548 585
R1144 B.n3 B.n0 585
R1145 B.n4 B.n3 585
R1146 B.n861 B.n1 585
R1147 B.n862 B.n861 585
R1148 B.n860 B.n859 585
R1149 B.n860 B.n8 585
R1150 B.n858 B.n9 585
R1151 B.n12 B.n9 585
R1152 B.n857 B.n856 585
R1153 B.n856 B.n855 585
R1154 B.n11 B.n10 585
R1155 B.n854 B.n11 585
R1156 B.n852 B.n851 585
R1157 B.n853 B.n852 585
R1158 B.n850 B.n16 585
R1159 B.n19 B.n16 585
R1160 B.n849 B.n848 585
R1161 B.n848 B.n847 585
R1162 B.n18 B.n17 585
R1163 B.n846 B.n18 585
R1164 B.n844 B.n843 585
R1165 B.n845 B.n844 585
R1166 B.n842 B.n24 585
R1167 B.n24 B.n23 585
R1168 B.n841 B.n840 585
R1169 B.n840 B.n839 585
R1170 B.n26 B.n25 585
R1171 B.n838 B.n26 585
R1172 B.n836 B.n835 585
R1173 B.n837 B.n836 585
R1174 B.n834 B.n31 585
R1175 B.n31 B.n30 585
R1176 B.n833 B.n832 585
R1177 B.n832 B.n831 585
R1178 B.n33 B.n32 585
R1179 B.n830 B.n33 585
R1180 B.n828 B.n827 585
R1181 B.n829 B.n828 585
R1182 B.n826 B.n37 585
R1183 B.n40 B.n37 585
R1184 B.n825 B.n824 585
R1185 B.n824 B.n823 585
R1186 B.n39 B.n38 585
R1187 B.n822 B.n39 585
R1188 B.n820 B.n819 585
R1189 B.n821 B.n820 585
R1190 B.n818 B.n45 585
R1191 B.n45 B.n44 585
R1192 B.n817 B.n816 585
R1193 B.n816 B.n815 585
R1194 B.n47 B.n46 585
R1195 B.n814 B.n47 585
R1196 B.n812 B.n811 585
R1197 B.n813 B.n812 585
R1198 B.n810 B.n52 585
R1199 B.n52 B.n51 585
R1200 B.n809 B.n808 585
R1201 B.n808 B.n807 585
R1202 B.n54 B.n53 585
R1203 B.n806 B.n54 585
R1204 B.n804 B.n803 585
R1205 B.n805 B.n804 585
R1206 B.n802 B.n59 585
R1207 B.n59 B.n58 585
R1208 B.n801 B.n800 585
R1209 B.n800 B.n799 585
R1210 B.n61 B.n60 585
R1211 B.n798 B.n61 585
R1212 B.n796 B.n795 585
R1213 B.n797 B.n796 585
R1214 B.n794 B.n66 585
R1215 B.n66 B.n65 585
R1216 B.n793 B.n792 585
R1217 B.n792 B.n791 585
R1218 B.n68 B.n67 585
R1219 B.n790 B.n68 585
R1220 B.n788 B.n787 585
R1221 B.n789 B.n788 585
R1222 B.n786 B.n73 585
R1223 B.n73 B.n72 585
R1224 B.n785 B.n784 585
R1225 B.n784 B.n783 585
R1226 B.n75 B.n74 585
R1227 B.n782 B.n75 585
R1228 B.n780 B.n779 585
R1229 B.n781 B.n780 585
R1230 B.n865 B.n864 585
R1231 B.n863 B.n2 585
R1232 B.n780 B.n80 454.062
R1233 B.n609 B.n78 454.062
R1234 B.n427 B.n206 454.062
R1235 B.n425 B.n208 454.062
R1236 B.n107 B.t13 333.25
R1237 B.n236 B.t10 333.25
R1238 B.n99 B.t16 333.25
R1239 B.n229 B.t7 333.25
R1240 B.n99 B.t15 280.906
R1241 B.n107 B.t11 280.906
R1242 B.n236 B.t8 280.906
R1243 B.n229 B.t4 280.906
R1244 B.n108 B.t14 257.808
R1245 B.n237 B.t9 257.808
R1246 B.n100 B.t17 257.808
R1247 B.n230 B.t6 257.808
R1248 B.n610 B.n79 256.663
R1249 B.n616 B.n79 256.663
R1250 B.n618 B.n79 256.663
R1251 B.n624 B.n79 256.663
R1252 B.n626 B.n79 256.663
R1253 B.n632 B.n79 256.663
R1254 B.n634 B.n79 256.663
R1255 B.n640 B.n79 256.663
R1256 B.n642 B.n79 256.663
R1257 B.n648 B.n79 256.663
R1258 B.n650 B.n79 256.663
R1259 B.n656 B.n79 256.663
R1260 B.n658 B.n79 256.663
R1261 B.n664 B.n79 256.663
R1262 B.n666 B.n79 256.663
R1263 B.n672 B.n79 256.663
R1264 B.n674 B.n79 256.663
R1265 B.n680 B.n79 256.663
R1266 B.n682 B.n79 256.663
R1267 B.n689 B.n79 256.663
R1268 B.n691 B.n79 256.663
R1269 B.n697 B.n79 256.663
R1270 B.n102 B.n79 256.663
R1271 B.n703 B.n79 256.663
R1272 B.n709 B.n79 256.663
R1273 B.n711 B.n79 256.663
R1274 B.n717 B.n79 256.663
R1275 B.n719 B.n79 256.663
R1276 B.n725 B.n79 256.663
R1277 B.n727 B.n79 256.663
R1278 B.n733 B.n79 256.663
R1279 B.n735 B.n79 256.663
R1280 B.n741 B.n79 256.663
R1281 B.n743 B.n79 256.663
R1282 B.n749 B.n79 256.663
R1283 B.n751 B.n79 256.663
R1284 B.n757 B.n79 256.663
R1285 B.n759 B.n79 256.663
R1286 B.n765 B.n79 256.663
R1287 B.n767 B.n79 256.663
R1288 B.n773 B.n79 256.663
R1289 B.n775 B.n79 256.663
R1290 B.n420 B.n207 256.663
R1291 B.n210 B.n207 256.663
R1292 B.n413 B.n207 256.663
R1293 B.n407 B.n207 256.663
R1294 B.n405 B.n207 256.663
R1295 B.n399 B.n207 256.663
R1296 B.n397 B.n207 256.663
R1297 B.n391 B.n207 256.663
R1298 B.n389 B.n207 256.663
R1299 B.n383 B.n207 256.663
R1300 B.n381 B.n207 256.663
R1301 B.n375 B.n207 256.663
R1302 B.n373 B.n207 256.663
R1303 B.n367 B.n207 256.663
R1304 B.n365 B.n207 256.663
R1305 B.n359 B.n207 256.663
R1306 B.n357 B.n207 256.663
R1307 B.n351 B.n207 256.663
R1308 B.n349 B.n207 256.663
R1309 B.n343 B.n207 256.663
R1310 B.n341 B.n207 256.663
R1311 B.n335 B.n207 256.663
R1312 B.n333 B.n207 256.663
R1313 B.n326 B.n207 256.663
R1314 B.n324 B.n207 256.663
R1315 B.n318 B.n207 256.663
R1316 B.n316 B.n207 256.663
R1317 B.n310 B.n207 256.663
R1318 B.n308 B.n207 256.663
R1319 B.n302 B.n207 256.663
R1320 B.n300 B.n207 256.663
R1321 B.n294 B.n207 256.663
R1322 B.n292 B.n207 256.663
R1323 B.n286 B.n207 256.663
R1324 B.n284 B.n207 256.663
R1325 B.n278 B.n207 256.663
R1326 B.n276 B.n207 256.663
R1327 B.n270 B.n207 256.663
R1328 B.n268 B.n207 256.663
R1329 B.n262 B.n207 256.663
R1330 B.n260 B.n207 256.663
R1331 B.n255 B.n207 256.663
R1332 B.n867 B.n866 256.663
R1333 B.n776 B.n774 163.367
R1334 B.n772 B.n82 163.367
R1335 B.n768 B.n766 163.367
R1336 B.n764 B.n84 163.367
R1337 B.n760 B.n758 163.367
R1338 B.n756 B.n86 163.367
R1339 B.n752 B.n750 163.367
R1340 B.n748 B.n88 163.367
R1341 B.n744 B.n742 163.367
R1342 B.n740 B.n90 163.367
R1343 B.n736 B.n734 163.367
R1344 B.n732 B.n92 163.367
R1345 B.n728 B.n726 163.367
R1346 B.n724 B.n94 163.367
R1347 B.n720 B.n718 163.367
R1348 B.n716 B.n96 163.367
R1349 B.n712 B.n710 163.367
R1350 B.n708 B.n98 163.367
R1351 B.n704 B.n702 163.367
R1352 B.n699 B.n698 163.367
R1353 B.n696 B.n104 163.367
R1354 B.n692 B.n690 163.367
R1355 B.n688 B.n106 163.367
R1356 B.n683 B.n681 163.367
R1357 B.n679 B.n110 163.367
R1358 B.n675 B.n673 163.367
R1359 B.n671 B.n112 163.367
R1360 B.n667 B.n665 163.367
R1361 B.n663 B.n114 163.367
R1362 B.n659 B.n657 163.367
R1363 B.n655 B.n116 163.367
R1364 B.n651 B.n649 163.367
R1365 B.n647 B.n118 163.367
R1366 B.n643 B.n641 163.367
R1367 B.n639 B.n120 163.367
R1368 B.n635 B.n633 163.367
R1369 B.n631 B.n122 163.367
R1370 B.n627 B.n625 163.367
R1371 B.n623 B.n124 163.367
R1372 B.n619 B.n617 163.367
R1373 B.n615 B.n126 163.367
R1374 B.n611 B.n609 163.367
R1375 B.n427 B.n204 163.367
R1376 B.n431 B.n204 163.367
R1377 B.n431 B.n198 163.367
R1378 B.n439 B.n198 163.367
R1379 B.n439 B.n196 163.367
R1380 B.n443 B.n196 163.367
R1381 B.n443 B.n189 163.367
R1382 B.n451 B.n189 163.367
R1383 B.n451 B.n187 163.367
R1384 B.n455 B.n187 163.367
R1385 B.n455 B.n182 163.367
R1386 B.n463 B.n182 163.367
R1387 B.n463 B.n180 163.367
R1388 B.n467 B.n180 163.367
R1389 B.n467 B.n174 163.367
R1390 B.n475 B.n174 163.367
R1391 B.n475 B.n172 163.367
R1392 B.n479 B.n172 163.367
R1393 B.n479 B.n166 163.367
R1394 B.n487 B.n166 163.367
R1395 B.n487 B.n164 163.367
R1396 B.n491 B.n164 163.367
R1397 B.n491 B.n159 163.367
R1398 B.n500 B.n159 163.367
R1399 B.n500 B.n157 163.367
R1400 B.n504 B.n157 163.367
R1401 B.n504 B.n151 163.367
R1402 B.n512 B.n151 163.367
R1403 B.n512 B.n149 163.367
R1404 B.n516 B.n149 163.367
R1405 B.n516 B.n143 163.367
R1406 B.n524 B.n143 163.367
R1407 B.n524 B.n141 163.367
R1408 B.n528 B.n141 163.367
R1409 B.n528 B.n136 163.367
R1410 B.n537 B.n136 163.367
R1411 B.n537 B.n134 163.367
R1412 B.n542 B.n134 163.367
R1413 B.n542 B.n128 163.367
R1414 B.n550 B.n128 163.367
R1415 B.n551 B.n550 163.367
R1416 B.n551 B.n5 163.367
R1417 B.n6 B.n5 163.367
R1418 B.n7 B.n6 163.367
R1419 B.n557 B.n7 163.367
R1420 B.n558 B.n557 163.367
R1421 B.n558 B.n13 163.367
R1422 B.n14 B.n13 163.367
R1423 B.n15 B.n14 163.367
R1424 B.n563 B.n15 163.367
R1425 B.n563 B.n20 163.367
R1426 B.n21 B.n20 163.367
R1427 B.n22 B.n21 163.367
R1428 B.n568 B.n22 163.367
R1429 B.n568 B.n27 163.367
R1430 B.n28 B.n27 163.367
R1431 B.n29 B.n28 163.367
R1432 B.n573 B.n29 163.367
R1433 B.n573 B.n34 163.367
R1434 B.n35 B.n34 163.367
R1435 B.n36 B.n35 163.367
R1436 B.n578 B.n36 163.367
R1437 B.n578 B.n41 163.367
R1438 B.n42 B.n41 163.367
R1439 B.n43 B.n42 163.367
R1440 B.n583 B.n43 163.367
R1441 B.n583 B.n48 163.367
R1442 B.n49 B.n48 163.367
R1443 B.n50 B.n49 163.367
R1444 B.n588 B.n50 163.367
R1445 B.n588 B.n55 163.367
R1446 B.n56 B.n55 163.367
R1447 B.n57 B.n56 163.367
R1448 B.n593 B.n57 163.367
R1449 B.n593 B.n62 163.367
R1450 B.n63 B.n62 163.367
R1451 B.n64 B.n63 163.367
R1452 B.n598 B.n64 163.367
R1453 B.n598 B.n69 163.367
R1454 B.n70 B.n69 163.367
R1455 B.n71 B.n70 163.367
R1456 B.n603 B.n71 163.367
R1457 B.n603 B.n76 163.367
R1458 B.n77 B.n76 163.367
R1459 B.n78 B.n77 163.367
R1460 B.n421 B.n419 163.367
R1461 B.n419 B.n418 163.367
R1462 B.n415 B.n414 163.367
R1463 B.n412 B.n212 163.367
R1464 B.n408 B.n406 163.367
R1465 B.n404 B.n214 163.367
R1466 B.n400 B.n398 163.367
R1467 B.n396 B.n216 163.367
R1468 B.n392 B.n390 163.367
R1469 B.n388 B.n218 163.367
R1470 B.n384 B.n382 163.367
R1471 B.n380 B.n220 163.367
R1472 B.n376 B.n374 163.367
R1473 B.n372 B.n222 163.367
R1474 B.n368 B.n366 163.367
R1475 B.n364 B.n224 163.367
R1476 B.n360 B.n358 163.367
R1477 B.n356 B.n226 163.367
R1478 B.n352 B.n350 163.367
R1479 B.n348 B.n228 163.367
R1480 B.n344 B.n342 163.367
R1481 B.n340 B.n233 163.367
R1482 B.n336 B.n334 163.367
R1483 B.n332 B.n235 163.367
R1484 B.n327 B.n325 163.367
R1485 B.n323 B.n239 163.367
R1486 B.n319 B.n317 163.367
R1487 B.n315 B.n241 163.367
R1488 B.n311 B.n309 163.367
R1489 B.n307 B.n243 163.367
R1490 B.n303 B.n301 163.367
R1491 B.n299 B.n245 163.367
R1492 B.n295 B.n293 163.367
R1493 B.n291 B.n247 163.367
R1494 B.n287 B.n285 163.367
R1495 B.n283 B.n249 163.367
R1496 B.n279 B.n277 163.367
R1497 B.n275 B.n251 163.367
R1498 B.n271 B.n269 163.367
R1499 B.n267 B.n253 163.367
R1500 B.n263 B.n261 163.367
R1501 B.n259 B.n256 163.367
R1502 B.n425 B.n202 163.367
R1503 B.n433 B.n202 163.367
R1504 B.n433 B.n200 163.367
R1505 B.n437 B.n200 163.367
R1506 B.n437 B.n194 163.367
R1507 B.n445 B.n194 163.367
R1508 B.n445 B.n192 163.367
R1509 B.n449 B.n192 163.367
R1510 B.n449 B.n186 163.367
R1511 B.n457 B.n186 163.367
R1512 B.n457 B.n184 163.367
R1513 B.n461 B.n184 163.367
R1514 B.n461 B.n178 163.367
R1515 B.n469 B.n178 163.367
R1516 B.n469 B.n176 163.367
R1517 B.n473 B.n176 163.367
R1518 B.n473 B.n170 163.367
R1519 B.n481 B.n170 163.367
R1520 B.n481 B.n168 163.367
R1521 B.n485 B.n168 163.367
R1522 B.n485 B.n162 163.367
R1523 B.n494 B.n162 163.367
R1524 B.n494 B.n160 163.367
R1525 B.n498 B.n160 163.367
R1526 B.n498 B.n155 163.367
R1527 B.n506 B.n155 163.367
R1528 B.n506 B.n153 163.367
R1529 B.n510 B.n153 163.367
R1530 B.n510 B.n147 163.367
R1531 B.n518 B.n147 163.367
R1532 B.n518 B.n145 163.367
R1533 B.n522 B.n145 163.367
R1534 B.n522 B.n139 163.367
R1535 B.n531 B.n139 163.367
R1536 B.n531 B.n137 163.367
R1537 B.n535 B.n137 163.367
R1538 B.n535 B.n132 163.367
R1539 B.n544 B.n132 163.367
R1540 B.n544 B.n130 163.367
R1541 B.n548 B.n130 163.367
R1542 B.n548 B.n3 163.367
R1543 B.n865 B.n3 163.367
R1544 B.n861 B.n2 163.367
R1545 B.n861 B.n860 163.367
R1546 B.n860 B.n9 163.367
R1547 B.n856 B.n9 163.367
R1548 B.n856 B.n11 163.367
R1549 B.n852 B.n11 163.367
R1550 B.n852 B.n16 163.367
R1551 B.n848 B.n16 163.367
R1552 B.n848 B.n18 163.367
R1553 B.n844 B.n18 163.367
R1554 B.n844 B.n24 163.367
R1555 B.n840 B.n24 163.367
R1556 B.n840 B.n26 163.367
R1557 B.n836 B.n26 163.367
R1558 B.n836 B.n31 163.367
R1559 B.n832 B.n31 163.367
R1560 B.n832 B.n33 163.367
R1561 B.n828 B.n33 163.367
R1562 B.n828 B.n37 163.367
R1563 B.n824 B.n37 163.367
R1564 B.n824 B.n39 163.367
R1565 B.n820 B.n39 163.367
R1566 B.n820 B.n45 163.367
R1567 B.n816 B.n45 163.367
R1568 B.n816 B.n47 163.367
R1569 B.n812 B.n47 163.367
R1570 B.n812 B.n52 163.367
R1571 B.n808 B.n52 163.367
R1572 B.n808 B.n54 163.367
R1573 B.n804 B.n54 163.367
R1574 B.n804 B.n59 163.367
R1575 B.n800 B.n59 163.367
R1576 B.n800 B.n61 163.367
R1577 B.n796 B.n61 163.367
R1578 B.n796 B.n66 163.367
R1579 B.n792 B.n66 163.367
R1580 B.n792 B.n68 163.367
R1581 B.n788 B.n68 163.367
R1582 B.n788 B.n73 163.367
R1583 B.n784 B.n73 163.367
R1584 B.n784 B.n75 163.367
R1585 B.n780 B.n75 163.367
R1586 B.n426 B.n207 82.4572
R1587 B.n781 B.n79 82.4572
R1588 B.n100 B.n99 75.4429
R1589 B.n108 B.n107 75.4429
R1590 B.n237 B.n236 75.4429
R1591 B.n230 B.n229 75.4429
R1592 B.n775 B.n80 71.676
R1593 B.n774 B.n773 71.676
R1594 B.n767 B.n82 71.676
R1595 B.n766 B.n765 71.676
R1596 B.n759 B.n84 71.676
R1597 B.n758 B.n757 71.676
R1598 B.n751 B.n86 71.676
R1599 B.n750 B.n749 71.676
R1600 B.n743 B.n88 71.676
R1601 B.n742 B.n741 71.676
R1602 B.n735 B.n90 71.676
R1603 B.n734 B.n733 71.676
R1604 B.n727 B.n92 71.676
R1605 B.n726 B.n725 71.676
R1606 B.n719 B.n94 71.676
R1607 B.n718 B.n717 71.676
R1608 B.n711 B.n96 71.676
R1609 B.n710 B.n709 71.676
R1610 B.n703 B.n98 71.676
R1611 B.n702 B.n102 71.676
R1612 B.n698 B.n697 71.676
R1613 B.n691 B.n104 71.676
R1614 B.n690 B.n689 71.676
R1615 B.n682 B.n106 71.676
R1616 B.n681 B.n680 71.676
R1617 B.n674 B.n110 71.676
R1618 B.n673 B.n672 71.676
R1619 B.n666 B.n112 71.676
R1620 B.n665 B.n664 71.676
R1621 B.n658 B.n114 71.676
R1622 B.n657 B.n656 71.676
R1623 B.n650 B.n116 71.676
R1624 B.n649 B.n648 71.676
R1625 B.n642 B.n118 71.676
R1626 B.n641 B.n640 71.676
R1627 B.n634 B.n120 71.676
R1628 B.n633 B.n632 71.676
R1629 B.n626 B.n122 71.676
R1630 B.n625 B.n624 71.676
R1631 B.n618 B.n124 71.676
R1632 B.n617 B.n616 71.676
R1633 B.n610 B.n126 71.676
R1634 B.n611 B.n610 71.676
R1635 B.n616 B.n615 71.676
R1636 B.n619 B.n618 71.676
R1637 B.n624 B.n623 71.676
R1638 B.n627 B.n626 71.676
R1639 B.n632 B.n631 71.676
R1640 B.n635 B.n634 71.676
R1641 B.n640 B.n639 71.676
R1642 B.n643 B.n642 71.676
R1643 B.n648 B.n647 71.676
R1644 B.n651 B.n650 71.676
R1645 B.n656 B.n655 71.676
R1646 B.n659 B.n658 71.676
R1647 B.n664 B.n663 71.676
R1648 B.n667 B.n666 71.676
R1649 B.n672 B.n671 71.676
R1650 B.n675 B.n674 71.676
R1651 B.n680 B.n679 71.676
R1652 B.n683 B.n682 71.676
R1653 B.n689 B.n688 71.676
R1654 B.n692 B.n691 71.676
R1655 B.n697 B.n696 71.676
R1656 B.n699 B.n102 71.676
R1657 B.n704 B.n703 71.676
R1658 B.n709 B.n708 71.676
R1659 B.n712 B.n711 71.676
R1660 B.n717 B.n716 71.676
R1661 B.n720 B.n719 71.676
R1662 B.n725 B.n724 71.676
R1663 B.n728 B.n727 71.676
R1664 B.n733 B.n732 71.676
R1665 B.n736 B.n735 71.676
R1666 B.n741 B.n740 71.676
R1667 B.n744 B.n743 71.676
R1668 B.n749 B.n748 71.676
R1669 B.n752 B.n751 71.676
R1670 B.n757 B.n756 71.676
R1671 B.n760 B.n759 71.676
R1672 B.n765 B.n764 71.676
R1673 B.n768 B.n767 71.676
R1674 B.n773 B.n772 71.676
R1675 B.n776 B.n775 71.676
R1676 B.n420 B.n208 71.676
R1677 B.n418 B.n210 71.676
R1678 B.n414 B.n413 71.676
R1679 B.n407 B.n212 71.676
R1680 B.n406 B.n405 71.676
R1681 B.n399 B.n214 71.676
R1682 B.n398 B.n397 71.676
R1683 B.n391 B.n216 71.676
R1684 B.n390 B.n389 71.676
R1685 B.n383 B.n218 71.676
R1686 B.n382 B.n381 71.676
R1687 B.n375 B.n220 71.676
R1688 B.n374 B.n373 71.676
R1689 B.n367 B.n222 71.676
R1690 B.n366 B.n365 71.676
R1691 B.n359 B.n224 71.676
R1692 B.n358 B.n357 71.676
R1693 B.n351 B.n226 71.676
R1694 B.n350 B.n349 71.676
R1695 B.n343 B.n228 71.676
R1696 B.n342 B.n341 71.676
R1697 B.n335 B.n233 71.676
R1698 B.n334 B.n333 71.676
R1699 B.n326 B.n235 71.676
R1700 B.n325 B.n324 71.676
R1701 B.n318 B.n239 71.676
R1702 B.n317 B.n316 71.676
R1703 B.n310 B.n241 71.676
R1704 B.n309 B.n308 71.676
R1705 B.n302 B.n243 71.676
R1706 B.n301 B.n300 71.676
R1707 B.n294 B.n245 71.676
R1708 B.n293 B.n292 71.676
R1709 B.n286 B.n247 71.676
R1710 B.n285 B.n284 71.676
R1711 B.n278 B.n249 71.676
R1712 B.n277 B.n276 71.676
R1713 B.n270 B.n251 71.676
R1714 B.n269 B.n268 71.676
R1715 B.n262 B.n253 71.676
R1716 B.n261 B.n260 71.676
R1717 B.n256 B.n255 71.676
R1718 B.n421 B.n420 71.676
R1719 B.n415 B.n210 71.676
R1720 B.n413 B.n412 71.676
R1721 B.n408 B.n407 71.676
R1722 B.n405 B.n404 71.676
R1723 B.n400 B.n399 71.676
R1724 B.n397 B.n396 71.676
R1725 B.n392 B.n391 71.676
R1726 B.n389 B.n388 71.676
R1727 B.n384 B.n383 71.676
R1728 B.n381 B.n380 71.676
R1729 B.n376 B.n375 71.676
R1730 B.n373 B.n372 71.676
R1731 B.n368 B.n367 71.676
R1732 B.n365 B.n364 71.676
R1733 B.n360 B.n359 71.676
R1734 B.n357 B.n356 71.676
R1735 B.n352 B.n351 71.676
R1736 B.n349 B.n348 71.676
R1737 B.n344 B.n343 71.676
R1738 B.n341 B.n340 71.676
R1739 B.n336 B.n335 71.676
R1740 B.n333 B.n332 71.676
R1741 B.n327 B.n326 71.676
R1742 B.n324 B.n323 71.676
R1743 B.n319 B.n318 71.676
R1744 B.n316 B.n315 71.676
R1745 B.n311 B.n310 71.676
R1746 B.n308 B.n307 71.676
R1747 B.n303 B.n302 71.676
R1748 B.n300 B.n299 71.676
R1749 B.n295 B.n294 71.676
R1750 B.n292 B.n291 71.676
R1751 B.n287 B.n286 71.676
R1752 B.n284 B.n283 71.676
R1753 B.n279 B.n278 71.676
R1754 B.n276 B.n275 71.676
R1755 B.n271 B.n270 71.676
R1756 B.n268 B.n267 71.676
R1757 B.n263 B.n262 71.676
R1758 B.n260 B.n259 71.676
R1759 B.n255 B.n206 71.676
R1760 B.n866 B.n865 71.676
R1761 B.n866 B.n2 71.676
R1762 B.n101 B.n100 59.5399
R1763 B.n685 B.n108 59.5399
R1764 B.n330 B.n237 59.5399
R1765 B.n231 B.n230 59.5399
R1766 B.n426 B.n203 47.1186
R1767 B.n432 B.n203 47.1186
R1768 B.n432 B.n199 47.1186
R1769 B.n438 B.n199 47.1186
R1770 B.n438 B.n195 47.1186
R1771 B.n444 B.n195 47.1186
R1772 B.n444 B.n190 47.1186
R1773 B.n450 B.n190 47.1186
R1774 B.n450 B.n191 47.1186
R1775 B.n456 B.n183 47.1186
R1776 B.n462 B.n183 47.1186
R1777 B.n462 B.n179 47.1186
R1778 B.n468 B.n179 47.1186
R1779 B.n468 B.n175 47.1186
R1780 B.n474 B.n175 47.1186
R1781 B.n474 B.n171 47.1186
R1782 B.n480 B.n171 47.1186
R1783 B.n480 B.n167 47.1186
R1784 B.n486 B.n167 47.1186
R1785 B.n486 B.n163 47.1186
R1786 B.n493 B.n163 47.1186
R1787 B.n493 B.n492 47.1186
R1788 B.n499 B.n156 47.1186
R1789 B.n505 B.n156 47.1186
R1790 B.n505 B.n152 47.1186
R1791 B.n511 B.n152 47.1186
R1792 B.n511 B.n148 47.1186
R1793 B.n517 B.n148 47.1186
R1794 B.n517 B.n144 47.1186
R1795 B.n523 B.n144 47.1186
R1796 B.n523 B.n140 47.1186
R1797 B.n530 B.n140 47.1186
R1798 B.n530 B.n529 47.1186
R1799 B.n536 B.n133 47.1186
R1800 B.n543 B.n133 47.1186
R1801 B.n543 B.n129 47.1186
R1802 B.n549 B.n129 47.1186
R1803 B.n549 B.n4 47.1186
R1804 B.n864 B.n4 47.1186
R1805 B.n864 B.n863 47.1186
R1806 B.n863 B.n862 47.1186
R1807 B.n862 B.n8 47.1186
R1808 B.n12 B.n8 47.1186
R1809 B.n855 B.n12 47.1186
R1810 B.n855 B.n854 47.1186
R1811 B.n854 B.n853 47.1186
R1812 B.n847 B.n19 47.1186
R1813 B.n847 B.n846 47.1186
R1814 B.n846 B.n845 47.1186
R1815 B.n845 B.n23 47.1186
R1816 B.n839 B.n23 47.1186
R1817 B.n839 B.n838 47.1186
R1818 B.n838 B.n837 47.1186
R1819 B.n837 B.n30 47.1186
R1820 B.n831 B.n30 47.1186
R1821 B.n831 B.n830 47.1186
R1822 B.n830 B.n829 47.1186
R1823 B.n823 B.n40 47.1186
R1824 B.n823 B.n822 47.1186
R1825 B.n822 B.n821 47.1186
R1826 B.n821 B.n44 47.1186
R1827 B.n815 B.n44 47.1186
R1828 B.n815 B.n814 47.1186
R1829 B.n814 B.n813 47.1186
R1830 B.n813 B.n51 47.1186
R1831 B.n807 B.n51 47.1186
R1832 B.n807 B.n806 47.1186
R1833 B.n806 B.n805 47.1186
R1834 B.n805 B.n58 47.1186
R1835 B.n799 B.n58 47.1186
R1836 B.n798 B.n797 47.1186
R1837 B.n797 B.n65 47.1186
R1838 B.n791 B.n65 47.1186
R1839 B.n791 B.n790 47.1186
R1840 B.n790 B.n789 47.1186
R1841 B.n789 B.n72 47.1186
R1842 B.n783 B.n72 47.1186
R1843 B.n783 B.n782 47.1186
R1844 B.n782 B.n781 47.1186
R1845 B.n456 B.t5 42.9611
R1846 B.n799 B.t12 42.9611
R1847 B.n536 B.t1 38.8037
R1848 B.n853 B.t0 38.8037
R1849 B.n492 B.t2 34.6462
R1850 B.n40 B.t3 34.6462
R1851 B.n608 B.n607 29.5029
R1852 B.n424 B.n423 29.5029
R1853 B.n428 B.n205 29.5029
R1854 B.n779 B.n778 29.5029
R1855 B B.n867 18.0485
R1856 B.n499 B.t2 12.4729
R1857 B.n829 B.t3 12.4729
R1858 B.n424 B.n201 10.6151
R1859 B.n434 B.n201 10.6151
R1860 B.n435 B.n434 10.6151
R1861 B.n436 B.n435 10.6151
R1862 B.n436 B.n193 10.6151
R1863 B.n446 B.n193 10.6151
R1864 B.n447 B.n446 10.6151
R1865 B.n448 B.n447 10.6151
R1866 B.n448 B.n185 10.6151
R1867 B.n458 B.n185 10.6151
R1868 B.n459 B.n458 10.6151
R1869 B.n460 B.n459 10.6151
R1870 B.n460 B.n177 10.6151
R1871 B.n470 B.n177 10.6151
R1872 B.n471 B.n470 10.6151
R1873 B.n472 B.n471 10.6151
R1874 B.n472 B.n169 10.6151
R1875 B.n482 B.n169 10.6151
R1876 B.n483 B.n482 10.6151
R1877 B.n484 B.n483 10.6151
R1878 B.n484 B.n161 10.6151
R1879 B.n495 B.n161 10.6151
R1880 B.n496 B.n495 10.6151
R1881 B.n497 B.n496 10.6151
R1882 B.n497 B.n154 10.6151
R1883 B.n507 B.n154 10.6151
R1884 B.n508 B.n507 10.6151
R1885 B.n509 B.n508 10.6151
R1886 B.n509 B.n146 10.6151
R1887 B.n519 B.n146 10.6151
R1888 B.n520 B.n519 10.6151
R1889 B.n521 B.n520 10.6151
R1890 B.n521 B.n138 10.6151
R1891 B.n532 B.n138 10.6151
R1892 B.n533 B.n532 10.6151
R1893 B.n534 B.n533 10.6151
R1894 B.n534 B.n131 10.6151
R1895 B.n545 B.n131 10.6151
R1896 B.n546 B.n545 10.6151
R1897 B.n547 B.n546 10.6151
R1898 B.n547 B.n0 10.6151
R1899 B.n423 B.n422 10.6151
R1900 B.n422 B.n209 10.6151
R1901 B.n417 B.n209 10.6151
R1902 B.n417 B.n416 10.6151
R1903 B.n416 B.n211 10.6151
R1904 B.n411 B.n211 10.6151
R1905 B.n411 B.n410 10.6151
R1906 B.n410 B.n409 10.6151
R1907 B.n409 B.n213 10.6151
R1908 B.n403 B.n213 10.6151
R1909 B.n403 B.n402 10.6151
R1910 B.n402 B.n401 10.6151
R1911 B.n401 B.n215 10.6151
R1912 B.n395 B.n215 10.6151
R1913 B.n395 B.n394 10.6151
R1914 B.n394 B.n393 10.6151
R1915 B.n393 B.n217 10.6151
R1916 B.n387 B.n217 10.6151
R1917 B.n387 B.n386 10.6151
R1918 B.n386 B.n385 10.6151
R1919 B.n385 B.n219 10.6151
R1920 B.n379 B.n219 10.6151
R1921 B.n379 B.n378 10.6151
R1922 B.n378 B.n377 10.6151
R1923 B.n377 B.n221 10.6151
R1924 B.n371 B.n221 10.6151
R1925 B.n371 B.n370 10.6151
R1926 B.n370 B.n369 10.6151
R1927 B.n369 B.n223 10.6151
R1928 B.n363 B.n223 10.6151
R1929 B.n363 B.n362 10.6151
R1930 B.n362 B.n361 10.6151
R1931 B.n361 B.n225 10.6151
R1932 B.n355 B.n225 10.6151
R1933 B.n355 B.n354 10.6151
R1934 B.n354 B.n353 10.6151
R1935 B.n353 B.n227 10.6151
R1936 B.n347 B.n346 10.6151
R1937 B.n346 B.n345 10.6151
R1938 B.n345 B.n232 10.6151
R1939 B.n339 B.n232 10.6151
R1940 B.n339 B.n338 10.6151
R1941 B.n338 B.n337 10.6151
R1942 B.n337 B.n234 10.6151
R1943 B.n331 B.n234 10.6151
R1944 B.n329 B.n328 10.6151
R1945 B.n328 B.n238 10.6151
R1946 B.n322 B.n238 10.6151
R1947 B.n322 B.n321 10.6151
R1948 B.n321 B.n320 10.6151
R1949 B.n320 B.n240 10.6151
R1950 B.n314 B.n240 10.6151
R1951 B.n314 B.n313 10.6151
R1952 B.n313 B.n312 10.6151
R1953 B.n312 B.n242 10.6151
R1954 B.n306 B.n242 10.6151
R1955 B.n306 B.n305 10.6151
R1956 B.n305 B.n304 10.6151
R1957 B.n304 B.n244 10.6151
R1958 B.n298 B.n244 10.6151
R1959 B.n298 B.n297 10.6151
R1960 B.n297 B.n296 10.6151
R1961 B.n296 B.n246 10.6151
R1962 B.n290 B.n246 10.6151
R1963 B.n290 B.n289 10.6151
R1964 B.n289 B.n288 10.6151
R1965 B.n288 B.n248 10.6151
R1966 B.n282 B.n248 10.6151
R1967 B.n282 B.n281 10.6151
R1968 B.n281 B.n280 10.6151
R1969 B.n280 B.n250 10.6151
R1970 B.n274 B.n250 10.6151
R1971 B.n274 B.n273 10.6151
R1972 B.n273 B.n272 10.6151
R1973 B.n272 B.n252 10.6151
R1974 B.n266 B.n252 10.6151
R1975 B.n266 B.n265 10.6151
R1976 B.n265 B.n264 10.6151
R1977 B.n264 B.n254 10.6151
R1978 B.n258 B.n254 10.6151
R1979 B.n258 B.n257 10.6151
R1980 B.n257 B.n205 10.6151
R1981 B.n429 B.n428 10.6151
R1982 B.n430 B.n429 10.6151
R1983 B.n430 B.n197 10.6151
R1984 B.n440 B.n197 10.6151
R1985 B.n441 B.n440 10.6151
R1986 B.n442 B.n441 10.6151
R1987 B.n442 B.n188 10.6151
R1988 B.n452 B.n188 10.6151
R1989 B.n453 B.n452 10.6151
R1990 B.n454 B.n453 10.6151
R1991 B.n454 B.n181 10.6151
R1992 B.n464 B.n181 10.6151
R1993 B.n465 B.n464 10.6151
R1994 B.n466 B.n465 10.6151
R1995 B.n466 B.n173 10.6151
R1996 B.n476 B.n173 10.6151
R1997 B.n477 B.n476 10.6151
R1998 B.n478 B.n477 10.6151
R1999 B.n478 B.n165 10.6151
R2000 B.n488 B.n165 10.6151
R2001 B.n489 B.n488 10.6151
R2002 B.n490 B.n489 10.6151
R2003 B.n490 B.n158 10.6151
R2004 B.n501 B.n158 10.6151
R2005 B.n502 B.n501 10.6151
R2006 B.n503 B.n502 10.6151
R2007 B.n503 B.n150 10.6151
R2008 B.n513 B.n150 10.6151
R2009 B.n514 B.n513 10.6151
R2010 B.n515 B.n514 10.6151
R2011 B.n515 B.n142 10.6151
R2012 B.n525 B.n142 10.6151
R2013 B.n526 B.n525 10.6151
R2014 B.n527 B.n526 10.6151
R2015 B.n527 B.n135 10.6151
R2016 B.n538 B.n135 10.6151
R2017 B.n539 B.n538 10.6151
R2018 B.n541 B.n539 10.6151
R2019 B.n541 B.n540 10.6151
R2020 B.n540 B.n127 10.6151
R2021 B.n552 B.n127 10.6151
R2022 B.n553 B.n552 10.6151
R2023 B.n554 B.n553 10.6151
R2024 B.n555 B.n554 10.6151
R2025 B.n556 B.n555 10.6151
R2026 B.n559 B.n556 10.6151
R2027 B.n560 B.n559 10.6151
R2028 B.n561 B.n560 10.6151
R2029 B.n562 B.n561 10.6151
R2030 B.n564 B.n562 10.6151
R2031 B.n565 B.n564 10.6151
R2032 B.n566 B.n565 10.6151
R2033 B.n567 B.n566 10.6151
R2034 B.n569 B.n567 10.6151
R2035 B.n570 B.n569 10.6151
R2036 B.n571 B.n570 10.6151
R2037 B.n572 B.n571 10.6151
R2038 B.n574 B.n572 10.6151
R2039 B.n575 B.n574 10.6151
R2040 B.n576 B.n575 10.6151
R2041 B.n577 B.n576 10.6151
R2042 B.n579 B.n577 10.6151
R2043 B.n580 B.n579 10.6151
R2044 B.n581 B.n580 10.6151
R2045 B.n582 B.n581 10.6151
R2046 B.n584 B.n582 10.6151
R2047 B.n585 B.n584 10.6151
R2048 B.n586 B.n585 10.6151
R2049 B.n587 B.n586 10.6151
R2050 B.n589 B.n587 10.6151
R2051 B.n590 B.n589 10.6151
R2052 B.n591 B.n590 10.6151
R2053 B.n592 B.n591 10.6151
R2054 B.n594 B.n592 10.6151
R2055 B.n595 B.n594 10.6151
R2056 B.n596 B.n595 10.6151
R2057 B.n597 B.n596 10.6151
R2058 B.n599 B.n597 10.6151
R2059 B.n600 B.n599 10.6151
R2060 B.n601 B.n600 10.6151
R2061 B.n602 B.n601 10.6151
R2062 B.n604 B.n602 10.6151
R2063 B.n605 B.n604 10.6151
R2064 B.n606 B.n605 10.6151
R2065 B.n607 B.n606 10.6151
R2066 B.n859 B.n1 10.6151
R2067 B.n859 B.n858 10.6151
R2068 B.n858 B.n857 10.6151
R2069 B.n857 B.n10 10.6151
R2070 B.n851 B.n10 10.6151
R2071 B.n851 B.n850 10.6151
R2072 B.n850 B.n849 10.6151
R2073 B.n849 B.n17 10.6151
R2074 B.n843 B.n17 10.6151
R2075 B.n843 B.n842 10.6151
R2076 B.n842 B.n841 10.6151
R2077 B.n841 B.n25 10.6151
R2078 B.n835 B.n25 10.6151
R2079 B.n835 B.n834 10.6151
R2080 B.n834 B.n833 10.6151
R2081 B.n833 B.n32 10.6151
R2082 B.n827 B.n32 10.6151
R2083 B.n827 B.n826 10.6151
R2084 B.n826 B.n825 10.6151
R2085 B.n825 B.n38 10.6151
R2086 B.n819 B.n38 10.6151
R2087 B.n819 B.n818 10.6151
R2088 B.n818 B.n817 10.6151
R2089 B.n817 B.n46 10.6151
R2090 B.n811 B.n46 10.6151
R2091 B.n811 B.n810 10.6151
R2092 B.n810 B.n809 10.6151
R2093 B.n809 B.n53 10.6151
R2094 B.n803 B.n53 10.6151
R2095 B.n803 B.n802 10.6151
R2096 B.n802 B.n801 10.6151
R2097 B.n801 B.n60 10.6151
R2098 B.n795 B.n60 10.6151
R2099 B.n795 B.n794 10.6151
R2100 B.n794 B.n793 10.6151
R2101 B.n793 B.n67 10.6151
R2102 B.n787 B.n67 10.6151
R2103 B.n787 B.n786 10.6151
R2104 B.n786 B.n785 10.6151
R2105 B.n785 B.n74 10.6151
R2106 B.n779 B.n74 10.6151
R2107 B.n778 B.n777 10.6151
R2108 B.n777 B.n81 10.6151
R2109 B.n771 B.n81 10.6151
R2110 B.n771 B.n770 10.6151
R2111 B.n770 B.n769 10.6151
R2112 B.n769 B.n83 10.6151
R2113 B.n763 B.n83 10.6151
R2114 B.n763 B.n762 10.6151
R2115 B.n762 B.n761 10.6151
R2116 B.n761 B.n85 10.6151
R2117 B.n755 B.n85 10.6151
R2118 B.n755 B.n754 10.6151
R2119 B.n754 B.n753 10.6151
R2120 B.n753 B.n87 10.6151
R2121 B.n747 B.n87 10.6151
R2122 B.n747 B.n746 10.6151
R2123 B.n746 B.n745 10.6151
R2124 B.n745 B.n89 10.6151
R2125 B.n739 B.n89 10.6151
R2126 B.n739 B.n738 10.6151
R2127 B.n738 B.n737 10.6151
R2128 B.n737 B.n91 10.6151
R2129 B.n731 B.n91 10.6151
R2130 B.n731 B.n730 10.6151
R2131 B.n730 B.n729 10.6151
R2132 B.n729 B.n93 10.6151
R2133 B.n723 B.n93 10.6151
R2134 B.n723 B.n722 10.6151
R2135 B.n722 B.n721 10.6151
R2136 B.n721 B.n95 10.6151
R2137 B.n715 B.n95 10.6151
R2138 B.n715 B.n714 10.6151
R2139 B.n714 B.n713 10.6151
R2140 B.n713 B.n97 10.6151
R2141 B.n707 B.n97 10.6151
R2142 B.n707 B.n706 10.6151
R2143 B.n706 B.n705 10.6151
R2144 B.n701 B.n700 10.6151
R2145 B.n700 B.n103 10.6151
R2146 B.n695 B.n103 10.6151
R2147 B.n695 B.n694 10.6151
R2148 B.n694 B.n693 10.6151
R2149 B.n693 B.n105 10.6151
R2150 B.n687 B.n105 10.6151
R2151 B.n687 B.n686 10.6151
R2152 B.n684 B.n109 10.6151
R2153 B.n678 B.n109 10.6151
R2154 B.n678 B.n677 10.6151
R2155 B.n677 B.n676 10.6151
R2156 B.n676 B.n111 10.6151
R2157 B.n670 B.n111 10.6151
R2158 B.n670 B.n669 10.6151
R2159 B.n669 B.n668 10.6151
R2160 B.n668 B.n113 10.6151
R2161 B.n662 B.n113 10.6151
R2162 B.n662 B.n661 10.6151
R2163 B.n661 B.n660 10.6151
R2164 B.n660 B.n115 10.6151
R2165 B.n654 B.n115 10.6151
R2166 B.n654 B.n653 10.6151
R2167 B.n653 B.n652 10.6151
R2168 B.n652 B.n117 10.6151
R2169 B.n646 B.n117 10.6151
R2170 B.n646 B.n645 10.6151
R2171 B.n645 B.n644 10.6151
R2172 B.n644 B.n119 10.6151
R2173 B.n638 B.n119 10.6151
R2174 B.n638 B.n637 10.6151
R2175 B.n637 B.n636 10.6151
R2176 B.n636 B.n121 10.6151
R2177 B.n630 B.n121 10.6151
R2178 B.n630 B.n629 10.6151
R2179 B.n629 B.n628 10.6151
R2180 B.n628 B.n123 10.6151
R2181 B.n622 B.n123 10.6151
R2182 B.n622 B.n621 10.6151
R2183 B.n621 B.n620 10.6151
R2184 B.n620 B.n125 10.6151
R2185 B.n614 B.n125 10.6151
R2186 B.n614 B.n613 10.6151
R2187 B.n613 B.n612 10.6151
R2188 B.n612 B.n608 10.6151
R2189 B.n529 B.t1 8.31546
R2190 B.n19 B.t0 8.31546
R2191 B.n867 B.n0 8.11757
R2192 B.n867 B.n1 8.11757
R2193 B.n347 B.n231 6.5566
R2194 B.n331 B.n330 6.5566
R2195 B.n701 B.n101 6.5566
R2196 B.n686 B.n685 6.5566
R2197 B.n191 B.t5 4.15798
R2198 B.t12 B.n798 4.15798
R2199 B.n231 B.n227 4.05904
R2200 B.n330 B.n329 4.05904
R2201 B.n705 B.n101 4.05904
R2202 B.n685 B.n684 4.05904
R2203 VP.n19 VP.n18 161.3
R2204 VP.n17 VP.n1 161.3
R2205 VP.n16 VP.n15 161.3
R2206 VP.n14 VP.n2 161.3
R2207 VP.n13 VP.n12 161.3
R2208 VP.n11 VP.n3 161.3
R2209 VP.n10 VP.n9 161.3
R2210 VP.n8 VP.n4 161.3
R2211 VP.n5 VP.t2 106.547
R2212 VP.n5 VP.t0 105.311
R2213 VP.n7 VP.n6 80.6547
R2214 VP.n20 VP.n0 80.6547
R2215 VP.n6 VP.t1 71.7589
R2216 VP.n0 VP.t3 71.7589
R2217 VP.n12 VP.n2 56.5617
R2218 VP.n7 VP.n5 50.3945
R2219 VP.n10 VP.n4 24.5923
R2220 VP.n11 VP.n10 24.5923
R2221 VP.n12 VP.n11 24.5923
R2222 VP.n16 VP.n2 24.5923
R2223 VP.n17 VP.n16 24.5923
R2224 VP.n18 VP.n17 24.5923
R2225 VP.n6 VP.n4 9.59132
R2226 VP.n18 VP.n0 9.59132
R2227 VP.n8 VP.n7 0.354861
R2228 VP.n20 VP.n19 0.354861
R2229 VP VP.n20 0.267071
R2230 VP.n9 VP.n8 0.189894
R2231 VP.n9 VP.n3 0.189894
R2232 VP.n13 VP.n3 0.189894
R2233 VP.n14 VP.n13 0.189894
R2234 VP.n15 VP.n14 0.189894
R2235 VP.n15 VP.n1 0.189894
R2236 VP.n19 VP.n1 0.189894
R2237 VDD1 VDD1.n1 104.227
R2238 VDD1 VDD1.n0 60.8468
R2239 VDD1.n0 VDD1.t1 1.86842
R2240 VDD1.n0 VDD1.t3 1.86842
R2241 VDD1.n1 VDD1.t2 1.86842
R2242 VDD1.n1 VDD1.t0 1.86842
C0 VP VN 6.61882f
C1 VP VTAIL 4.57839f
C2 VP VDD1 4.74659f
C3 VP VDD2 0.455877f
C4 VN VTAIL 4.56429f
C5 VN VDD1 0.150352f
C6 VN VDD2 4.44204f
C7 VDD1 VTAIL 5.36383f
C8 VDD2 VTAIL 5.42447f
C9 VDD1 VDD2 1.25721f
C10 VDD2 B 4.208403f
C11 VDD1 B 8.57163f
C12 VTAIL B 9.754914f
C13 VN B 12.45034f
C14 VP B 10.88239f
C15 VDD1.t1 B 0.232252f
C16 VDD1.t3 B 0.232252f
C17 VDD1.n0 B 2.05191f
C18 VDD1.t2 B 0.232252f
C19 VDD1.t0 B 0.232252f
C20 VDD1.n1 B 2.78207f
C21 VP.t3 B 2.21835f
C22 VP.n0 B 0.867013f
C23 VP.n1 B 0.021658f
C24 VP.n2 B 0.031483f
C25 VP.n3 B 0.021658f
C26 VP.n4 B 0.028068f
C27 VP.t2 B 2.52957f
C28 VP.t0 B 2.51902f
C29 VP.n5 B 2.8403f
C30 VP.t1 B 2.21835f
C31 VP.n6 B 0.867013f
C32 VP.n7 B 1.25623f
C33 VP.n8 B 0.034949f
C34 VP.n9 B 0.021658f
C35 VP.n10 B 0.040162f
C36 VP.n11 B 0.040162f
C37 VP.n12 B 0.031483f
C38 VP.n13 B 0.021658f
C39 VP.n14 B 0.021658f
C40 VP.n15 B 0.021658f
C41 VP.n16 B 0.040162f
C42 VP.n17 B 0.040162f
C43 VP.n18 B 0.028068f
C44 VP.n19 B 0.034949f
C45 VP.n20 B 0.059071f
C46 VDD2.t0 B 0.227662f
C47 VDD2.t3 B 0.227662f
C48 VDD2.n0 B 2.69977f
C49 VDD2.t2 B 0.227662f
C50 VDD2.t1 B 0.227662f
C51 VDD2.n1 B 2.01084f
C52 VDD2.n2 B 3.87921f
C53 VTAIL.n0 B 0.022812f
C54 VTAIL.n1 B 0.017579f
C55 VTAIL.n2 B 0.009446f
C56 VTAIL.n3 B 0.022328f
C57 VTAIL.n4 B 0.010002f
C58 VTAIL.n5 B 0.017579f
C59 VTAIL.n6 B 0.009446f
C60 VTAIL.n7 B 0.022328f
C61 VTAIL.n8 B 0.010002f
C62 VTAIL.n9 B 0.017579f
C63 VTAIL.n10 B 0.009446f
C64 VTAIL.n11 B 0.022328f
C65 VTAIL.n12 B 0.010002f
C66 VTAIL.n13 B 0.017579f
C67 VTAIL.n14 B 0.009446f
C68 VTAIL.n15 B 0.022328f
C69 VTAIL.n16 B 0.010002f
C70 VTAIL.n17 B 0.117297f
C71 VTAIL.t3 B 0.037578f
C72 VTAIL.n18 B 0.016746f
C73 VTAIL.n19 B 0.015784f
C74 VTAIL.n20 B 0.009446f
C75 VTAIL.n21 B 0.777378f
C76 VTAIL.n22 B 0.017579f
C77 VTAIL.n23 B 0.009446f
C78 VTAIL.n24 B 0.010002f
C79 VTAIL.n25 B 0.022328f
C80 VTAIL.n26 B 0.022328f
C81 VTAIL.n27 B 0.010002f
C82 VTAIL.n28 B 0.009446f
C83 VTAIL.n29 B 0.017579f
C84 VTAIL.n30 B 0.017579f
C85 VTAIL.n31 B 0.009446f
C86 VTAIL.n32 B 0.010002f
C87 VTAIL.n33 B 0.022328f
C88 VTAIL.n34 B 0.022328f
C89 VTAIL.n35 B 0.022328f
C90 VTAIL.n36 B 0.010002f
C91 VTAIL.n37 B 0.009446f
C92 VTAIL.n38 B 0.017579f
C93 VTAIL.n39 B 0.017579f
C94 VTAIL.n40 B 0.009446f
C95 VTAIL.n41 B 0.009724f
C96 VTAIL.n42 B 0.009724f
C97 VTAIL.n43 B 0.022328f
C98 VTAIL.n44 B 0.022328f
C99 VTAIL.n45 B 0.010002f
C100 VTAIL.n46 B 0.009446f
C101 VTAIL.n47 B 0.017579f
C102 VTAIL.n48 B 0.017579f
C103 VTAIL.n49 B 0.009446f
C104 VTAIL.n50 B 0.010002f
C105 VTAIL.n51 B 0.022328f
C106 VTAIL.n52 B 0.04498f
C107 VTAIL.n53 B 0.010002f
C108 VTAIL.n54 B 0.009446f
C109 VTAIL.n55 B 0.038713f
C110 VTAIL.n56 B 0.024763f
C111 VTAIL.n57 B 0.138817f
C112 VTAIL.n58 B 0.022812f
C113 VTAIL.n59 B 0.017579f
C114 VTAIL.n60 B 0.009446f
C115 VTAIL.n61 B 0.022328f
C116 VTAIL.n62 B 0.010002f
C117 VTAIL.n63 B 0.017579f
C118 VTAIL.n64 B 0.009446f
C119 VTAIL.n65 B 0.022328f
C120 VTAIL.n66 B 0.010002f
C121 VTAIL.n67 B 0.017579f
C122 VTAIL.n68 B 0.009446f
C123 VTAIL.n69 B 0.022328f
C124 VTAIL.n70 B 0.010002f
C125 VTAIL.n71 B 0.017579f
C126 VTAIL.n72 B 0.009446f
C127 VTAIL.n73 B 0.022328f
C128 VTAIL.n74 B 0.010002f
C129 VTAIL.n75 B 0.117297f
C130 VTAIL.t5 B 0.037578f
C131 VTAIL.n76 B 0.016746f
C132 VTAIL.n77 B 0.015784f
C133 VTAIL.n78 B 0.009446f
C134 VTAIL.n79 B 0.777378f
C135 VTAIL.n80 B 0.017579f
C136 VTAIL.n81 B 0.009446f
C137 VTAIL.n82 B 0.010002f
C138 VTAIL.n83 B 0.022328f
C139 VTAIL.n84 B 0.022328f
C140 VTAIL.n85 B 0.010002f
C141 VTAIL.n86 B 0.009446f
C142 VTAIL.n87 B 0.017579f
C143 VTAIL.n88 B 0.017579f
C144 VTAIL.n89 B 0.009446f
C145 VTAIL.n90 B 0.010002f
C146 VTAIL.n91 B 0.022328f
C147 VTAIL.n92 B 0.022328f
C148 VTAIL.n93 B 0.022328f
C149 VTAIL.n94 B 0.010002f
C150 VTAIL.n95 B 0.009446f
C151 VTAIL.n96 B 0.017579f
C152 VTAIL.n97 B 0.017579f
C153 VTAIL.n98 B 0.009446f
C154 VTAIL.n99 B 0.009724f
C155 VTAIL.n100 B 0.009724f
C156 VTAIL.n101 B 0.022328f
C157 VTAIL.n102 B 0.022328f
C158 VTAIL.n103 B 0.010002f
C159 VTAIL.n104 B 0.009446f
C160 VTAIL.n105 B 0.017579f
C161 VTAIL.n106 B 0.017579f
C162 VTAIL.n107 B 0.009446f
C163 VTAIL.n108 B 0.010002f
C164 VTAIL.n109 B 0.022328f
C165 VTAIL.n110 B 0.04498f
C166 VTAIL.n111 B 0.010002f
C167 VTAIL.n112 B 0.009446f
C168 VTAIL.n113 B 0.038713f
C169 VTAIL.n114 B 0.024763f
C170 VTAIL.n115 B 0.230498f
C171 VTAIL.n116 B 0.022812f
C172 VTAIL.n117 B 0.017579f
C173 VTAIL.n118 B 0.009446f
C174 VTAIL.n119 B 0.022328f
C175 VTAIL.n120 B 0.010002f
C176 VTAIL.n121 B 0.017579f
C177 VTAIL.n122 B 0.009446f
C178 VTAIL.n123 B 0.022328f
C179 VTAIL.n124 B 0.010002f
C180 VTAIL.n125 B 0.017579f
C181 VTAIL.n126 B 0.009446f
C182 VTAIL.n127 B 0.022328f
C183 VTAIL.n128 B 0.010002f
C184 VTAIL.n129 B 0.017579f
C185 VTAIL.n130 B 0.009446f
C186 VTAIL.n131 B 0.022328f
C187 VTAIL.n132 B 0.010002f
C188 VTAIL.n133 B 0.117297f
C189 VTAIL.t6 B 0.037578f
C190 VTAIL.n134 B 0.016746f
C191 VTAIL.n135 B 0.015784f
C192 VTAIL.n136 B 0.009446f
C193 VTAIL.n137 B 0.777378f
C194 VTAIL.n138 B 0.017579f
C195 VTAIL.n139 B 0.009446f
C196 VTAIL.n140 B 0.010002f
C197 VTAIL.n141 B 0.022328f
C198 VTAIL.n142 B 0.022328f
C199 VTAIL.n143 B 0.010002f
C200 VTAIL.n144 B 0.009446f
C201 VTAIL.n145 B 0.017579f
C202 VTAIL.n146 B 0.017579f
C203 VTAIL.n147 B 0.009446f
C204 VTAIL.n148 B 0.010002f
C205 VTAIL.n149 B 0.022328f
C206 VTAIL.n150 B 0.022328f
C207 VTAIL.n151 B 0.022328f
C208 VTAIL.n152 B 0.010002f
C209 VTAIL.n153 B 0.009446f
C210 VTAIL.n154 B 0.017579f
C211 VTAIL.n155 B 0.017579f
C212 VTAIL.n156 B 0.009446f
C213 VTAIL.n157 B 0.009724f
C214 VTAIL.n158 B 0.009724f
C215 VTAIL.n159 B 0.022328f
C216 VTAIL.n160 B 0.022328f
C217 VTAIL.n161 B 0.010002f
C218 VTAIL.n162 B 0.009446f
C219 VTAIL.n163 B 0.017579f
C220 VTAIL.n164 B 0.017579f
C221 VTAIL.n165 B 0.009446f
C222 VTAIL.n166 B 0.010002f
C223 VTAIL.n167 B 0.022328f
C224 VTAIL.n168 B 0.04498f
C225 VTAIL.n169 B 0.010002f
C226 VTAIL.n170 B 0.009446f
C227 VTAIL.n171 B 0.038713f
C228 VTAIL.n172 B 0.024763f
C229 VTAIL.n173 B 1.15025f
C230 VTAIL.n174 B 0.022812f
C231 VTAIL.n175 B 0.017579f
C232 VTAIL.n176 B 0.009446f
C233 VTAIL.n177 B 0.022328f
C234 VTAIL.n178 B 0.010002f
C235 VTAIL.n179 B 0.017579f
C236 VTAIL.n180 B 0.009446f
C237 VTAIL.n181 B 0.022328f
C238 VTAIL.n182 B 0.010002f
C239 VTAIL.n183 B 0.017579f
C240 VTAIL.n184 B 0.009446f
C241 VTAIL.n185 B 0.022328f
C242 VTAIL.n186 B 0.022328f
C243 VTAIL.n187 B 0.010002f
C244 VTAIL.n188 B 0.017579f
C245 VTAIL.n189 B 0.009446f
C246 VTAIL.n190 B 0.022328f
C247 VTAIL.n191 B 0.010002f
C248 VTAIL.n192 B 0.117297f
C249 VTAIL.t2 B 0.037578f
C250 VTAIL.n193 B 0.016746f
C251 VTAIL.n194 B 0.015784f
C252 VTAIL.n195 B 0.009446f
C253 VTAIL.n196 B 0.777378f
C254 VTAIL.n197 B 0.017579f
C255 VTAIL.n198 B 0.009446f
C256 VTAIL.n199 B 0.010002f
C257 VTAIL.n200 B 0.022328f
C258 VTAIL.n201 B 0.022328f
C259 VTAIL.n202 B 0.010002f
C260 VTAIL.n203 B 0.009446f
C261 VTAIL.n204 B 0.017579f
C262 VTAIL.n205 B 0.017579f
C263 VTAIL.n206 B 0.009446f
C264 VTAIL.n207 B 0.010002f
C265 VTAIL.n208 B 0.022328f
C266 VTAIL.n209 B 0.022328f
C267 VTAIL.n210 B 0.010002f
C268 VTAIL.n211 B 0.009446f
C269 VTAIL.n212 B 0.017579f
C270 VTAIL.n213 B 0.017579f
C271 VTAIL.n214 B 0.009446f
C272 VTAIL.n215 B 0.009724f
C273 VTAIL.n216 B 0.009724f
C274 VTAIL.n217 B 0.022328f
C275 VTAIL.n218 B 0.022328f
C276 VTAIL.n219 B 0.010002f
C277 VTAIL.n220 B 0.009446f
C278 VTAIL.n221 B 0.017579f
C279 VTAIL.n222 B 0.017579f
C280 VTAIL.n223 B 0.009446f
C281 VTAIL.n224 B 0.010002f
C282 VTAIL.n225 B 0.022328f
C283 VTAIL.n226 B 0.04498f
C284 VTAIL.n227 B 0.010002f
C285 VTAIL.n228 B 0.009446f
C286 VTAIL.n229 B 0.038713f
C287 VTAIL.n230 B 0.024763f
C288 VTAIL.n231 B 1.15025f
C289 VTAIL.n232 B 0.022812f
C290 VTAIL.n233 B 0.017579f
C291 VTAIL.n234 B 0.009446f
C292 VTAIL.n235 B 0.022328f
C293 VTAIL.n236 B 0.010002f
C294 VTAIL.n237 B 0.017579f
C295 VTAIL.n238 B 0.009446f
C296 VTAIL.n239 B 0.022328f
C297 VTAIL.n240 B 0.010002f
C298 VTAIL.n241 B 0.017579f
C299 VTAIL.n242 B 0.009446f
C300 VTAIL.n243 B 0.022328f
C301 VTAIL.n244 B 0.022328f
C302 VTAIL.n245 B 0.010002f
C303 VTAIL.n246 B 0.017579f
C304 VTAIL.n247 B 0.009446f
C305 VTAIL.n248 B 0.022328f
C306 VTAIL.n249 B 0.010002f
C307 VTAIL.n250 B 0.117297f
C308 VTAIL.t0 B 0.037578f
C309 VTAIL.n251 B 0.016746f
C310 VTAIL.n252 B 0.015784f
C311 VTAIL.n253 B 0.009446f
C312 VTAIL.n254 B 0.777378f
C313 VTAIL.n255 B 0.017579f
C314 VTAIL.n256 B 0.009446f
C315 VTAIL.n257 B 0.010002f
C316 VTAIL.n258 B 0.022328f
C317 VTAIL.n259 B 0.022328f
C318 VTAIL.n260 B 0.010002f
C319 VTAIL.n261 B 0.009446f
C320 VTAIL.n262 B 0.017579f
C321 VTAIL.n263 B 0.017579f
C322 VTAIL.n264 B 0.009446f
C323 VTAIL.n265 B 0.010002f
C324 VTAIL.n266 B 0.022328f
C325 VTAIL.n267 B 0.022328f
C326 VTAIL.n268 B 0.010002f
C327 VTAIL.n269 B 0.009446f
C328 VTAIL.n270 B 0.017579f
C329 VTAIL.n271 B 0.017579f
C330 VTAIL.n272 B 0.009446f
C331 VTAIL.n273 B 0.009724f
C332 VTAIL.n274 B 0.009724f
C333 VTAIL.n275 B 0.022328f
C334 VTAIL.n276 B 0.022328f
C335 VTAIL.n277 B 0.010002f
C336 VTAIL.n278 B 0.009446f
C337 VTAIL.n279 B 0.017579f
C338 VTAIL.n280 B 0.017579f
C339 VTAIL.n281 B 0.009446f
C340 VTAIL.n282 B 0.010002f
C341 VTAIL.n283 B 0.022328f
C342 VTAIL.n284 B 0.04498f
C343 VTAIL.n285 B 0.010002f
C344 VTAIL.n286 B 0.009446f
C345 VTAIL.n287 B 0.038713f
C346 VTAIL.n288 B 0.024763f
C347 VTAIL.n289 B 0.230498f
C348 VTAIL.n290 B 0.022812f
C349 VTAIL.n291 B 0.017579f
C350 VTAIL.n292 B 0.009446f
C351 VTAIL.n293 B 0.022328f
C352 VTAIL.n294 B 0.010002f
C353 VTAIL.n295 B 0.017579f
C354 VTAIL.n296 B 0.009446f
C355 VTAIL.n297 B 0.022328f
C356 VTAIL.n298 B 0.010002f
C357 VTAIL.n299 B 0.017579f
C358 VTAIL.n300 B 0.009446f
C359 VTAIL.n301 B 0.022328f
C360 VTAIL.n302 B 0.022328f
C361 VTAIL.n303 B 0.010002f
C362 VTAIL.n304 B 0.017579f
C363 VTAIL.n305 B 0.009446f
C364 VTAIL.n306 B 0.022328f
C365 VTAIL.n307 B 0.010002f
C366 VTAIL.n308 B 0.117297f
C367 VTAIL.t4 B 0.037578f
C368 VTAIL.n309 B 0.016746f
C369 VTAIL.n310 B 0.015784f
C370 VTAIL.n311 B 0.009446f
C371 VTAIL.n312 B 0.777378f
C372 VTAIL.n313 B 0.017579f
C373 VTAIL.n314 B 0.009446f
C374 VTAIL.n315 B 0.010002f
C375 VTAIL.n316 B 0.022328f
C376 VTAIL.n317 B 0.022328f
C377 VTAIL.n318 B 0.010002f
C378 VTAIL.n319 B 0.009446f
C379 VTAIL.n320 B 0.017579f
C380 VTAIL.n321 B 0.017579f
C381 VTAIL.n322 B 0.009446f
C382 VTAIL.n323 B 0.010002f
C383 VTAIL.n324 B 0.022328f
C384 VTAIL.n325 B 0.022328f
C385 VTAIL.n326 B 0.010002f
C386 VTAIL.n327 B 0.009446f
C387 VTAIL.n328 B 0.017579f
C388 VTAIL.n329 B 0.017579f
C389 VTAIL.n330 B 0.009446f
C390 VTAIL.n331 B 0.009724f
C391 VTAIL.n332 B 0.009724f
C392 VTAIL.n333 B 0.022328f
C393 VTAIL.n334 B 0.022328f
C394 VTAIL.n335 B 0.010002f
C395 VTAIL.n336 B 0.009446f
C396 VTAIL.n337 B 0.017579f
C397 VTAIL.n338 B 0.017579f
C398 VTAIL.n339 B 0.009446f
C399 VTAIL.n340 B 0.010002f
C400 VTAIL.n341 B 0.022328f
C401 VTAIL.n342 B 0.04498f
C402 VTAIL.n343 B 0.010002f
C403 VTAIL.n344 B 0.009446f
C404 VTAIL.n345 B 0.038713f
C405 VTAIL.n346 B 0.024763f
C406 VTAIL.n347 B 0.230498f
C407 VTAIL.n348 B 0.022812f
C408 VTAIL.n349 B 0.017579f
C409 VTAIL.n350 B 0.009446f
C410 VTAIL.n351 B 0.022328f
C411 VTAIL.n352 B 0.010002f
C412 VTAIL.n353 B 0.017579f
C413 VTAIL.n354 B 0.009446f
C414 VTAIL.n355 B 0.022328f
C415 VTAIL.n356 B 0.010002f
C416 VTAIL.n357 B 0.017579f
C417 VTAIL.n358 B 0.009446f
C418 VTAIL.n359 B 0.022328f
C419 VTAIL.n360 B 0.022328f
C420 VTAIL.n361 B 0.010002f
C421 VTAIL.n362 B 0.017579f
C422 VTAIL.n363 B 0.009446f
C423 VTAIL.n364 B 0.022328f
C424 VTAIL.n365 B 0.010002f
C425 VTAIL.n366 B 0.117297f
C426 VTAIL.t7 B 0.037578f
C427 VTAIL.n367 B 0.016746f
C428 VTAIL.n368 B 0.015784f
C429 VTAIL.n369 B 0.009446f
C430 VTAIL.n370 B 0.777378f
C431 VTAIL.n371 B 0.017579f
C432 VTAIL.n372 B 0.009446f
C433 VTAIL.n373 B 0.010002f
C434 VTAIL.n374 B 0.022328f
C435 VTAIL.n375 B 0.022328f
C436 VTAIL.n376 B 0.010002f
C437 VTAIL.n377 B 0.009446f
C438 VTAIL.n378 B 0.017579f
C439 VTAIL.n379 B 0.017579f
C440 VTAIL.n380 B 0.009446f
C441 VTAIL.n381 B 0.010002f
C442 VTAIL.n382 B 0.022328f
C443 VTAIL.n383 B 0.022328f
C444 VTAIL.n384 B 0.010002f
C445 VTAIL.n385 B 0.009446f
C446 VTAIL.n386 B 0.017579f
C447 VTAIL.n387 B 0.017579f
C448 VTAIL.n388 B 0.009446f
C449 VTAIL.n389 B 0.009724f
C450 VTAIL.n390 B 0.009724f
C451 VTAIL.n391 B 0.022328f
C452 VTAIL.n392 B 0.022328f
C453 VTAIL.n393 B 0.010002f
C454 VTAIL.n394 B 0.009446f
C455 VTAIL.n395 B 0.017579f
C456 VTAIL.n396 B 0.017579f
C457 VTAIL.n397 B 0.009446f
C458 VTAIL.n398 B 0.010002f
C459 VTAIL.n399 B 0.022328f
C460 VTAIL.n400 B 0.04498f
C461 VTAIL.n401 B 0.010002f
C462 VTAIL.n402 B 0.009446f
C463 VTAIL.n403 B 0.038713f
C464 VTAIL.n404 B 0.024763f
C465 VTAIL.n405 B 1.15025f
C466 VTAIL.n406 B 0.022812f
C467 VTAIL.n407 B 0.017579f
C468 VTAIL.n408 B 0.009446f
C469 VTAIL.n409 B 0.022328f
C470 VTAIL.n410 B 0.010002f
C471 VTAIL.n411 B 0.017579f
C472 VTAIL.n412 B 0.009446f
C473 VTAIL.n413 B 0.022328f
C474 VTAIL.n414 B 0.010002f
C475 VTAIL.n415 B 0.017579f
C476 VTAIL.n416 B 0.009446f
C477 VTAIL.n417 B 0.022328f
C478 VTAIL.n418 B 0.010002f
C479 VTAIL.n419 B 0.017579f
C480 VTAIL.n420 B 0.009446f
C481 VTAIL.n421 B 0.022328f
C482 VTAIL.n422 B 0.010002f
C483 VTAIL.n423 B 0.117297f
C484 VTAIL.t1 B 0.037578f
C485 VTAIL.n424 B 0.016746f
C486 VTAIL.n425 B 0.015784f
C487 VTAIL.n426 B 0.009446f
C488 VTAIL.n427 B 0.777378f
C489 VTAIL.n428 B 0.017579f
C490 VTAIL.n429 B 0.009446f
C491 VTAIL.n430 B 0.010002f
C492 VTAIL.n431 B 0.022328f
C493 VTAIL.n432 B 0.022328f
C494 VTAIL.n433 B 0.010002f
C495 VTAIL.n434 B 0.009446f
C496 VTAIL.n435 B 0.017579f
C497 VTAIL.n436 B 0.017579f
C498 VTAIL.n437 B 0.009446f
C499 VTAIL.n438 B 0.010002f
C500 VTAIL.n439 B 0.022328f
C501 VTAIL.n440 B 0.022328f
C502 VTAIL.n441 B 0.022328f
C503 VTAIL.n442 B 0.010002f
C504 VTAIL.n443 B 0.009446f
C505 VTAIL.n444 B 0.017579f
C506 VTAIL.n445 B 0.017579f
C507 VTAIL.n446 B 0.009446f
C508 VTAIL.n447 B 0.009724f
C509 VTAIL.n448 B 0.009724f
C510 VTAIL.n449 B 0.022328f
C511 VTAIL.n450 B 0.022328f
C512 VTAIL.n451 B 0.010002f
C513 VTAIL.n452 B 0.009446f
C514 VTAIL.n453 B 0.017579f
C515 VTAIL.n454 B 0.017579f
C516 VTAIL.n455 B 0.009446f
C517 VTAIL.n456 B 0.010002f
C518 VTAIL.n457 B 0.022328f
C519 VTAIL.n458 B 0.04498f
C520 VTAIL.n459 B 0.010002f
C521 VTAIL.n460 B 0.009446f
C522 VTAIL.n461 B 0.038713f
C523 VTAIL.n462 B 0.024763f
C524 VTAIL.n463 B 1.05197f
C525 VN.t0 B 2.46677f
C526 VN.t3 B 2.4771f
C527 VN.n0 B 1.46644f
C528 VN.t2 B 2.4771f
C529 VN.t1 B 2.46677f
C530 VN.n1 B 2.78999f
.ends

