* NGSPICE file created from diff_pair_sample_0235.ext - technology: sky130A

.subckt diff_pair_sample_0235 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=2.9328 ps=15.82 w=7.52 l=2.45
X1 B.t11 B.t9 B.t10 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=0 ps=0 w=7.52 l=2.45
X2 VDD2.t1 VN.t0 VTAIL.t0 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=2.9328 ps=15.82 w=7.52 l=2.45
X3 B.t8 B.t6 B.t7 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=0 ps=0 w=7.52 l=2.45
X4 B.t5 B.t3 B.t4 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=0 ps=0 w=7.52 l=2.45
X5 B.t2 B.t0 B.t1 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=0 ps=0 w=7.52 l=2.45
X6 VDD1.t0 VP.t1 VTAIL.t3 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=2.9328 ps=15.82 w=7.52 l=2.45
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n2082_n2472# sky130_fd_pr__pfet_01v8 ad=2.9328 pd=15.82 as=2.9328 ps=15.82 w=7.52 l=2.45
R0 VP.n0 VP.t0 164.053
R1 VP.n0 VP.t1 123.188
R2 VP VP.n0 0.336784
R3 VTAIL.n1 VTAIL.t0 72.7354
R4 VTAIL.n3 VTAIL.t1 72.7352
R5 VTAIL.n0 VTAIL.t3 72.7352
R6 VTAIL.n2 VTAIL.t2 72.7352
R7 VTAIL.n1 VTAIL.n0 23.6427
R8 VTAIL.n3 VTAIL.n2 21.2462
R9 VTAIL.n2 VTAIL.n1 1.6686
R10 VTAIL VTAIL.n0 1.12766
R11 VTAIL VTAIL.n3 0.541448
R12 VDD1 VDD1.t0 125.474
R13 VDD1 VDD1.t1 90.0713
R14 B.n260 B.n259 585
R15 B.n258 B.n77 585
R16 B.n257 B.n256 585
R17 B.n255 B.n78 585
R18 B.n254 B.n253 585
R19 B.n252 B.n79 585
R20 B.n251 B.n250 585
R21 B.n249 B.n80 585
R22 B.n248 B.n247 585
R23 B.n246 B.n81 585
R24 B.n245 B.n244 585
R25 B.n243 B.n82 585
R26 B.n242 B.n241 585
R27 B.n240 B.n83 585
R28 B.n239 B.n238 585
R29 B.n237 B.n84 585
R30 B.n236 B.n235 585
R31 B.n234 B.n85 585
R32 B.n233 B.n232 585
R33 B.n231 B.n86 585
R34 B.n230 B.n229 585
R35 B.n228 B.n87 585
R36 B.n227 B.n226 585
R37 B.n225 B.n88 585
R38 B.n224 B.n223 585
R39 B.n222 B.n89 585
R40 B.n221 B.n220 585
R41 B.n219 B.n90 585
R42 B.n218 B.n217 585
R43 B.n213 B.n91 585
R44 B.n212 B.n211 585
R45 B.n210 B.n92 585
R46 B.n209 B.n208 585
R47 B.n207 B.n93 585
R48 B.n206 B.n205 585
R49 B.n204 B.n94 585
R50 B.n203 B.n202 585
R51 B.n201 B.n95 585
R52 B.n199 B.n198 585
R53 B.n197 B.n98 585
R54 B.n196 B.n195 585
R55 B.n194 B.n99 585
R56 B.n193 B.n192 585
R57 B.n191 B.n100 585
R58 B.n190 B.n189 585
R59 B.n188 B.n101 585
R60 B.n187 B.n186 585
R61 B.n185 B.n102 585
R62 B.n184 B.n183 585
R63 B.n182 B.n103 585
R64 B.n181 B.n180 585
R65 B.n179 B.n104 585
R66 B.n178 B.n177 585
R67 B.n176 B.n105 585
R68 B.n175 B.n174 585
R69 B.n173 B.n106 585
R70 B.n172 B.n171 585
R71 B.n170 B.n107 585
R72 B.n169 B.n168 585
R73 B.n167 B.n108 585
R74 B.n166 B.n165 585
R75 B.n164 B.n109 585
R76 B.n163 B.n162 585
R77 B.n161 B.n110 585
R78 B.n160 B.n159 585
R79 B.n158 B.n111 585
R80 B.n261 B.n76 585
R81 B.n263 B.n262 585
R82 B.n264 B.n75 585
R83 B.n266 B.n265 585
R84 B.n267 B.n74 585
R85 B.n269 B.n268 585
R86 B.n270 B.n73 585
R87 B.n272 B.n271 585
R88 B.n273 B.n72 585
R89 B.n275 B.n274 585
R90 B.n276 B.n71 585
R91 B.n278 B.n277 585
R92 B.n279 B.n70 585
R93 B.n281 B.n280 585
R94 B.n282 B.n69 585
R95 B.n284 B.n283 585
R96 B.n285 B.n68 585
R97 B.n287 B.n286 585
R98 B.n288 B.n67 585
R99 B.n290 B.n289 585
R100 B.n291 B.n66 585
R101 B.n293 B.n292 585
R102 B.n294 B.n65 585
R103 B.n296 B.n295 585
R104 B.n297 B.n64 585
R105 B.n299 B.n298 585
R106 B.n300 B.n63 585
R107 B.n302 B.n301 585
R108 B.n303 B.n62 585
R109 B.n305 B.n304 585
R110 B.n306 B.n61 585
R111 B.n308 B.n307 585
R112 B.n309 B.n60 585
R113 B.n311 B.n310 585
R114 B.n312 B.n59 585
R115 B.n314 B.n313 585
R116 B.n315 B.n58 585
R117 B.n317 B.n316 585
R118 B.n318 B.n57 585
R119 B.n320 B.n319 585
R120 B.n321 B.n56 585
R121 B.n323 B.n322 585
R122 B.n324 B.n55 585
R123 B.n326 B.n325 585
R124 B.n327 B.n54 585
R125 B.n329 B.n328 585
R126 B.n330 B.n53 585
R127 B.n332 B.n331 585
R128 B.n333 B.n52 585
R129 B.n335 B.n334 585
R130 B.n435 B.n14 585
R131 B.n434 B.n433 585
R132 B.n432 B.n15 585
R133 B.n431 B.n430 585
R134 B.n429 B.n16 585
R135 B.n428 B.n427 585
R136 B.n426 B.n17 585
R137 B.n425 B.n424 585
R138 B.n423 B.n18 585
R139 B.n422 B.n421 585
R140 B.n420 B.n19 585
R141 B.n419 B.n418 585
R142 B.n417 B.n20 585
R143 B.n416 B.n415 585
R144 B.n414 B.n21 585
R145 B.n413 B.n412 585
R146 B.n411 B.n22 585
R147 B.n410 B.n409 585
R148 B.n408 B.n23 585
R149 B.n407 B.n406 585
R150 B.n405 B.n24 585
R151 B.n404 B.n403 585
R152 B.n402 B.n25 585
R153 B.n401 B.n400 585
R154 B.n399 B.n26 585
R155 B.n398 B.n397 585
R156 B.n396 B.n27 585
R157 B.n395 B.n394 585
R158 B.n393 B.n392 585
R159 B.n391 B.n31 585
R160 B.n390 B.n389 585
R161 B.n388 B.n32 585
R162 B.n387 B.n386 585
R163 B.n385 B.n33 585
R164 B.n384 B.n383 585
R165 B.n382 B.n34 585
R166 B.n381 B.n380 585
R167 B.n379 B.n35 585
R168 B.n377 B.n376 585
R169 B.n375 B.n38 585
R170 B.n374 B.n373 585
R171 B.n372 B.n39 585
R172 B.n371 B.n370 585
R173 B.n369 B.n40 585
R174 B.n368 B.n367 585
R175 B.n366 B.n41 585
R176 B.n365 B.n364 585
R177 B.n363 B.n42 585
R178 B.n362 B.n361 585
R179 B.n360 B.n43 585
R180 B.n359 B.n358 585
R181 B.n357 B.n44 585
R182 B.n356 B.n355 585
R183 B.n354 B.n45 585
R184 B.n353 B.n352 585
R185 B.n351 B.n46 585
R186 B.n350 B.n349 585
R187 B.n348 B.n47 585
R188 B.n347 B.n346 585
R189 B.n345 B.n48 585
R190 B.n344 B.n343 585
R191 B.n342 B.n49 585
R192 B.n341 B.n340 585
R193 B.n339 B.n50 585
R194 B.n338 B.n337 585
R195 B.n336 B.n51 585
R196 B.n437 B.n436 585
R197 B.n438 B.n13 585
R198 B.n440 B.n439 585
R199 B.n441 B.n12 585
R200 B.n443 B.n442 585
R201 B.n444 B.n11 585
R202 B.n446 B.n445 585
R203 B.n447 B.n10 585
R204 B.n449 B.n448 585
R205 B.n450 B.n9 585
R206 B.n452 B.n451 585
R207 B.n453 B.n8 585
R208 B.n455 B.n454 585
R209 B.n456 B.n7 585
R210 B.n458 B.n457 585
R211 B.n459 B.n6 585
R212 B.n461 B.n460 585
R213 B.n462 B.n5 585
R214 B.n464 B.n463 585
R215 B.n465 B.n4 585
R216 B.n467 B.n466 585
R217 B.n468 B.n3 585
R218 B.n470 B.n469 585
R219 B.n471 B.n0 585
R220 B.n2 B.n1 585
R221 B.n124 B.n123 585
R222 B.n125 B.n122 585
R223 B.n127 B.n126 585
R224 B.n128 B.n121 585
R225 B.n130 B.n129 585
R226 B.n131 B.n120 585
R227 B.n133 B.n132 585
R228 B.n134 B.n119 585
R229 B.n136 B.n135 585
R230 B.n137 B.n118 585
R231 B.n139 B.n138 585
R232 B.n140 B.n117 585
R233 B.n142 B.n141 585
R234 B.n143 B.n116 585
R235 B.n145 B.n144 585
R236 B.n146 B.n115 585
R237 B.n148 B.n147 585
R238 B.n149 B.n114 585
R239 B.n151 B.n150 585
R240 B.n152 B.n113 585
R241 B.n154 B.n153 585
R242 B.n155 B.n112 585
R243 B.n157 B.n156 585
R244 B.n156 B.n111 530.939
R245 B.n261 B.n260 530.939
R246 B.n334 B.n51 530.939
R247 B.n436 B.n435 530.939
R248 B.n96 B.t9 281.781
R249 B.n214 B.t0 281.781
R250 B.n36 B.t3 281.781
R251 B.n28 B.t6 281.781
R252 B.n473 B.n472 256.663
R253 B.n472 B.n471 235.042
R254 B.n472 B.n2 235.042
R255 B.n214 B.t1 163.72
R256 B.n36 B.t5 163.72
R257 B.n96 B.t10 163.713
R258 B.n28 B.t8 163.713
R259 B.n160 B.n111 163.367
R260 B.n161 B.n160 163.367
R261 B.n162 B.n161 163.367
R262 B.n162 B.n109 163.367
R263 B.n166 B.n109 163.367
R264 B.n167 B.n166 163.367
R265 B.n168 B.n167 163.367
R266 B.n168 B.n107 163.367
R267 B.n172 B.n107 163.367
R268 B.n173 B.n172 163.367
R269 B.n174 B.n173 163.367
R270 B.n174 B.n105 163.367
R271 B.n178 B.n105 163.367
R272 B.n179 B.n178 163.367
R273 B.n180 B.n179 163.367
R274 B.n180 B.n103 163.367
R275 B.n184 B.n103 163.367
R276 B.n185 B.n184 163.367
R277 B.n186 B.n185 163.367
R278 B.n186 B.n101 163.367
R279 B.n190 B.n101 163.367
R280 B.n191 B.n190 163.367
R281 B.n192 B.n191 163.367
R282 B.n192 B.n99 163.367
R283 B.n196 B.n99 163.367
R284 B.n197 B.n196 163.367
R285 B.n198 B.n197 163.367
R286 B.n198 B.n95 163.367
R287 B.n203 B.n95 163.367
R288 B.n204 B.n203 163.367
R289 B.n205 B.n204 163.367
R290 B.n205 B.n93 163.367
R291 B.n209 B.n93 163.367
R292 B.n210 B.n209 163.367
R293 B.n211 B.n210 163.367
R294 B.n211 B.n91 163.367
R295 B.n218 B.n91 163.367
R296 B.n219 B.n218 163.367
R297 B.n220 B.n219 163.367
R298 B.n220 B.n89 163.367
R299 B.n224 B.n89 163.367
R300 B.n225 B.n224 163.367
R301 B.n226 B.n225 163.367
R302 B.n226 B.n87 163.367
R303 B.n230 B.n87 163.367
R304 B.n231 B.n230 163.367
R305 B.n232 B.n231 163.367
R306 B.n232 B.n85 163.367
R307 B.n236 B.n85 163.367
R308 B.n237 B.n236 163.367
R309 B.n238 B.n237 163.367
R310 B.n238 B.n83 163.367
R311 B.n242 B.n83 163.367
R312 B.n243 B.n242 163.367
R313 B.n244 B.n243 163.367
R314 B.n244 B.n81 163.367
R315 B.n248 B.n81 163.367
R316 B.n249 B.n248 163.367
R317 B.n250 B.n249 163.367
R318 B.n250 B.n79 163.367
R319 B.n254 B.n79 163.367
R320 B.n255 B.n254 163.367
R321 B.n256 B.n255 163.367
R322 B.n256 B.n77 163.367
R323 B.n260 B.n77 163.367
R324 B.n334 B.n333 163.367
R325 B.n333 B.n332 163.367
R326 B.n332 B.n53 163.367
R327 B.n328 B.n53 163.367
R328 B.n328 B.n327 163.367
R329 B.n327 B.n326 163.367
R330 B.n326 B.n55 163.367
R331 B.n322 B.n55 163.367
R332 B.n322 B.n321 163.367
R333 B.n321 B.n320 163.367
R334 B.n320 B.n57 163.367
R335 B.n316 B.n57 163.367
R336 B.n316 B.n315 163.367
R337 B.n315 B.n314 163.367
R338 B.n314 B.n59 163.367
R339 B.n310 B.n59 163.367
R340 B.n310 B.n309 163.367
R341 B.n309 B.n308 163.367
R342 B.n308 B.n61 163.367
R343 B.n304 B.n61 163.367
R344 B.n304 B.n303 163.367
R345 B.n303 B.n302 163.367
R346 B.n302 B.n63 163.367
R347 B.n298 B.n63 163.367
R348 B.n298 B.n297 163.367
R349 B.n297 B.n296 163.367
R350 B.n296 B.n65 163.367
R351 B.n292 B.n65 163.367
R352 B.n292 B.n291 163.367
R353 B.n291 B.n290 163.367
R354 B.n290 B.n67 163.367
R355 B.n286 B.n67 163.367
R356 B.n286 B.n285 163.367
R357 B.n285 B.n284 163.367
R358 B.n284 B.n69 163.367
R359 B.n280 B.n69 163.367
R360 B.n280 B.n279 163.367
R361 B.n279 B.n278 163.367
R362 B.n278 B.n71 163.367
R363 B.n274 B.n71 163.367
R364 B.n274 B.n273 163.367
R365 B.n273 B.n272 163.367
R366 B.n272 B.n73 163.367
R367 B.n268 B.n73 163.367
R368 B.n268 B.n267 163.367
R369 B.n267 B.n266 163.367
R370 B.n266 B.n75 163.367
R371 B.n262 B.n75 163.367
R372 B.n262 B.n261 163.367
R373 B.n435 B.n434 163.367
R374 B.n434 B.n15 163.367
R375 B.n430 B.n15 163.367
R376 B.n430 B.n429 163.367
R377 B.n429 B.n428 163.367
R378 B.n428 B.n17 163.367
R379 B.n424 B.n17 163.367
R380 B.n424 B.n423 163.367
R381 B.n423 B.n422 163.367
R382 B.n422 B.n19 163.367
R383 B.n418 B.n19 163.367
R384 B.n418 B.n417 163.367
R385 B.n417 B.n416 163.367
R386 B.n416 B.n21 163.367
R387 B.n412 B.n21 163.367
R388 B.n412 B.n411 163.367
R389 B.n411 B.n410 163.367
R390 B.n410 B.n23 163.367
R391 B.n406 B.n23 163.367
R392 B.n406 B.n405 163.367
R393 B.n405 B.n404 163.367
R394 B.n404 B.n25 163.367
R395 B.n400 B.n25 163.367
R396 B.n400 B.n399 163.367
R397 B.n399 B.n398 163.367
R398 B.n398 B.n27 163.367
R399 B.n394 B.n27 163.367
R400 B.n394 B.n393 163.367
R401 B.n393 B.n31 163.367
R402 B.n389 B.n31 163.367
R403 B.n389 B.n388 163.367
R404 B.n388 B.n387 163.367
R405 B.n387 B.n33 163.367
R406 B.n383 B.n33 163.367
R407 B.n383 B.n382 163.367
R408 B.n382 B.n381 163.367
R409 B.n381 B.n35 163.367
R410 B.n376 B.n35 163.367
R411 B.n376 B.n375 163.367
R412 B.n375 B.n374 163.367
R413 B.n374 B.n39 163.367
R414 B.n370 B.n39 163.367
R415 B.n370 B.n369 163.367
R416 B.n369 B.n368 163.367
R417 B.n368 B.n41 163.367
R418 B.n364 B.n41 163.367
R419 B.n364 B.n363 163.367
R420 B.n363 B.n362 163.367
R421 B.n362 B.n43 163.367
R422 B.n358 B.n43 163.367
R423 B.n358 B.n357 163.367
R424 B.n357 B.n356 163.367
R425 B.n356 B.n45 163.367
R426 B.n352 B.n45 163.367
R427 B.n352 B.n351 163.367
R428 B.n351 B.n350 163.367
R429 B.n350 B.n47 163.367
R430 B.n346 B.n47 163.367
R431 B.n346 B.n345 163.367
R432 B.n345 B.n344 163.367
R433 B.n344 B.n49 163.367
R434 B.n340 B.n49 163.367
R435 B.n340 B.n339 163.367
R436 B.n339 B.n338 163.367
R437 B.n338 B.n51 163.367
R438 B.n436 B.n13 163.367
R439 B.n440 B.n13 163.367
R440 B.n441 B.n440 163.367
R441 B.n442 B.n441 163.367
R442 B.n442 B.n11 163.367
R443 B.n446 B.n11 163.367
R444 B.n447 B.n446 163.367
R445 B.n448 B.n447 163.367
R446 B.n448 B.n9 163.367
R447 B.n452 B.n9 163.367
R448 B.n453 B.n452 163.367
R449 B.n454 B.n453 163.367
R450 B.n454 B.n7 163.367
R451 B.n458 B.n7 163.367
R452 B.n459 B.n458 163.367
R453 B.n460 B.n459 163.367
R454 B.n460 B.n5 163.367
R455 B.n464 B.n5 163.367
R456 B.n465 B.n464 163.367
R457 B.n466 B.n465 163.367
R458 B.n466 B.n3 163.367
R459 B.n470 B.n3 163.367
R460 B.n471 B.n470 163.367
R461 B.n124 B.n2 163.367
R462 B.n125 B.n124 163.367
R463 B.n126 B.n125 163.367
R464 B.n126 B.n121 163.367
R465 B.n130 B.n121 163.367
R466 B.n131 B.n130 163.367
R467 B.n132 B.n131 163.367
R468 B.n132 B.n119 163.367
R469 B.n136 B.n119 163.367
R470 B.n137 B.n136 163.367
R471 B.n138 B.n137 163.367
R472 B.n138 B.n117 163.367
R473 B.n142 B.n117 163.367
R474 B.n143 B.n142 163.367
R475 B.n144 B.n143 163.367
R476 B.n144 B.n115 163.367
R477 B.n148 B.n115 163.367
R478 B.n149 B.n148 163.367
R479 B.n150 B.n149 163.367
R480 B.n150 B.n113 163.367
R481 B.n154 B.n113 163.367
R482 B.n155 B.n154 163.367
R483 B.n156 B.n155 163.367
R484 B.n215 B.t2 109.805
R485 B.n37 B.t4 109.805
R486 B.n97 B.t11 109.797
R487 B.n29 B.t7 109.797
R488 B.n200 B.n97 59.5399
R489 B.n216 B.n215 59.5399
R490 B.n378 B.n37 59.5399
R491 B.n30 B.n29 59.5399
R492 B.n97 B.n96 53.9157
R493 B.n215 B.n214 53.9157
R494 B.n37 B.n36 53.9157
R495 B.n29 B.n28 53.9157
R496 B.n437 B.n14 34.4981
R497 B.n336 B.n335 34.4981
R498 B.n259 B.n76 34.4981
R499 B.n158 B.n157 34.4981
R500 B B.n473 18.0485
R501 B.n438 B.n437 10.6151
R502 B.n439 B.n438 10.6151
R503 B.n439 B.n12 10.6151
R504 B.n443 B.n12 10.6151
R505 B.n444 B.n443 10.6151
R506 B.n445 B.n444 10.6151
R507 B.n445 B.n10 10.6151
R508 B.n449 B.n10 10.6151
R509 B.n450 B.n449 10.6151
R510 B.n451 B.n450 10.6151
R511 B.n451 B.n8 10.6151
R512 B.n455 B.n8 10.6151
R513 B.n456 B.n455 10.6151
R514 B.n457 B.n456 10.6151
R515 B.n457 B.n6 10.6151
R516 B.n461 B.n6 10.6151
R517 B.n462 B.n461 10.6151
R518 B.n463 B.n462 10.6151
R519 B.n463 B.n4 10.6151
R520 B.n467 B.n4 10.6151
R521 B.n468 B.n467 10.6151
R522 B.n469 B.n468 10.6151
R523 B.n469 B.n0 10.6151
R524 B.n433 B.n14 10.6151
R525 B.n433 B.n432 10.6151
R526 B.n432 B.n431 10.6151
R527 B.n431 B.n16 10.6151
R528 B.n427 B.n16 10.6151
R529 B.n427 B.n426 10.6151
R530 B.n426 B.n425 10.6151
R531 B.n425 B.n18 10.6151
R532 B.n421 B.n18 10.6151
R533 B.n421 B.n420 10.6151
R534 B.n420 B.n419 10.6151
R535 B.n419 B.n20 10.6151
R536 B.n415 B.n20 10.6151
R537 B.n415 B.n414 10.6151
R538 B.n414 B.n413 10.6151
R539 B.n413 B.n22 10.6151
R540 B.n409 B.n22 10.6151
R541 B.n409 B.n408 10.6151
R542 B.n408 B.n407 10.6151
R543 B.n407 B.n24 10.6151
R544 B.n403 B.n24 10.6151
R545 B.n403 B.n402 10.6151
R546 B.n402 B.n401 10.6151
R547 B.n401 B.n26 10.6151
R548 B.n397 B.n26 10.6151
R549 B.n397 B.n396 10.6151
R550 B.n396 B.n395 10.6151
R551 B.n392 B.n391 10.6151
R552 B.n391 B.n390 10.6151
R553 B.n390 B.n32 10.6151
R554 B.n386 B.n32 10.6151
R555 B.n386 B.n385 10.6151
R556 B.n385 B.n384 10.6151
R557 B.n384 B.n34 10.6151
R558 B.n380 B.n34 10.6151
R559 B.n380 B.n379 10.6151
R560 B.n377 B.n38 10.6151
R561 B.n373 B.n38 10.6151
R562 B.n373 B.n372 10.6151
R563 B.n372 B.n371 10.6151
R564 B.n371 B.n40 10.6151
R565 B.n367 B.n40 10.6151
R566 B.n367 B.n366 10.6151
R567 B.n366 B.n365 10.6151
R568 B.n365 B.n42 10.6151
R569 B.n361 B.n42 10.6151
R570 B.n361 B.n360 10.6151
R571 B.n360 B.n359 10.6151
R572 B.n359 B.n44 10.6151
R573 B.n355 B.n44 10.6151
R574 B.n355 B.n354 10.6151
R575 B.n354 B.n353 10.6151
R576 B.n353 B.n46 10.6151
R577 B.n349 B.n46 10.6151
R578 B.n349 B.n348 10.6151
R579 B.n348 B.n347 10.6151
R580 B.n347 B.n48 10.6151
R581 B.n343 B.n48 10.6151
R582 B.n343 B.n342 10.6151
R583 B.n342 B.n341 10.6151
R584 B.n341 B.n50 10.6151
R585 B.n337 B.n50 10.6151
R586 B.n337 B.n336 10.6151
R587 B.n335 B.n52 10.6151
R588 B.n331 B.n52 10.6151
R589 B.n331 B.n330 10.6151
R590 B.n330 B.n329 10.6151
R591 B.n329 B.n54 10.6151
R592 B.n325 B.n54 10.6151
R593 B.n325 B.n324 10.6151
R594 B.n324 B.n323 10.6151
R595 B.n323 B.n56 10.6151
R596 B.n319 B.n56 10.6151
R597 B.n319 B.n318 10.6151
R598 B.n318 B.n317 10.6151
R599 B.n317 B.n58 10.6151
R600 B.n313 B.n58 10.6151
R601 B.n313 B.n312 10.6151
R602 B.n312 B.n311 10.6151
R603 B.n311 B.n60 10.6151
R604 B.n307 B.n60 10.6151
R605 B.n307 B.n306 10.6151
R606 B.n306 B.n305 10.6151
R607 B.n305 B.n62 10.6151
R608 B.n301 B.n62 10.6151
R609 B.n301 B.n300 10.6151
R610 B.n300 B.n299 10.6151
R611 B.n299 B.n64 10.6151
R612 B.n295 B.n64 10.6151
R613 B.n295 B.n294 10.6151
R614 B.n294 B.n293 10.6151
R615 B.n293 B.n66 10.6151
R616 B.n289 B.n66 10.6151
R617 B.n289 B.n288 10.6151
R618 B.n288 B.n287 10.6151
R619 B.n287 B.n68 10.6151
R620 B.n283 B.n68 10.6151
R621 B.n283 B.n282 10.6151
R622 B.n282 B.n281 10.6151
R623 B.n281 B.n70 10.6151
R624 B.n277 B.n70 10.6151
R625 B.n277 B.n276 10.6151
R626 B.n276 B.n275 10.6151
R627 B.n275 B.n72 10.6151
R628 B.n271 B.n72 10.6151
R629 B.n271 B.n270 10.6151
R630 B.n270 B.n269 10.6151
R631 B.n269 B.n74 10.6151
R632 B.n265 B.n74 10.6151
R633 B.n265 B.n264 10.6151
R634 B.n264 B.n263 10.6151
R635 B.n263 B.n76 10.6151
R636 B.n123 B.n1 10.6151
R637 B.n123 B.n122 10.6151
R638 B.n127 B.n122 10.6151
R639 B.n128 B.n127 10.6151
R640 B.n129 B.n128 10.6151
R641 B.n129 B.n120 10.6151
R642 B.n133 B.n120 10.6151
R643 B.n134 B.n133 10.6151
R644 B.n135 B.n134 10.6151
R645 B.n135 B.n118 10.6151
R646 B.n139 B.n118 10.6151
R647 B.n140 B.n139 10.6151
R648 B.n141 B.n140 10.6151
R649 B.n141 B.n116 10.6151
R650 B.n145 B.n116 10.6151
R651 B.n146 B.n145 10.6151
R652 B.n147 B.n146 10.6151
R653 B.n147 B.n114 10.6151
R654 B.n151 B.n114 10.6151
R655 B.n152 B.n151 10.6151
R656 B.n153 B.n152 10.6151
R657 B.n153 B.n112 10.6151
R658 B.n157 B.n112 10.6151
R659 B.n159 B.n158 10.6151
R660 B.n159 B.n110 10.6151
R661 B.n163 B.n110 10.6151
R662 B.n164 B.n163 10.6151
R663 B.n165 B.n164 10.6151
R664 B.n165 B.n108 10.6151
R665 B.n169 B.n108 10.6151
R666 B.n170 B.n169 10.6151
R667 B.n171 B.n170 10.6151
R668 B.n171 B.n106 10.6151
R669 B.n175 B.n106 10.6151
R670 B.n176 B.n175 10.6151
R671 B.n177 B.n176 10.6151
R672 B.n177 B.n104 10.6151
R673 B.n181 B.n104 10.6151
R674 B.n182 B.n181 10.6151
R675 B.n183 B.n182 10.6151
R676 B.n183 B.n102 10.6151
R677 B.n187 B.n102 10.6151
R678 B.n188 B.n187 10.6151
R679 B.n189 B.n188 10.6151
R680 B.n189 B.n100 10.6151
R681 B.n193 B.n100 10.6151
R682 B.n194 B.n193 10.6151
R683 B.n195 B.n194 10.6151
R684 B.n195 B.n98 10.6151
R685 B.n199 B.n98 10.6151
R686 B.n202 B.n201 10.6151
R687 B.n202 B.n94 10.6151
R688 B.n206 B.n94 10.6151
R689 B.n207 B.n206 10.6151
R690 B.n208 B.n207 10.6151
R691 B.n208 B.n92 10.6151
R692 B.n212 B.n92 10.6151
R693 B.n213 B.n212 10.6151
R694 B.n217 B.n213 10.6151
R695 B.n221 B.n90 10.6151
R696 B.n222 B.n221 10.6151
R697 B.n223 B.n222 10.6151
R698 B.n223 B.n88 10.6151
R699 B.n227 B.n88 10.6151
R700 B.n228 B.n227 10.6151
R701 B.n229 B.n228 10.6151
R702 B.n229 B.n86 10.6151
R703 B.n233 B.n86 10.6151
R704 B.n234 B.n233 10.6151
R705 B.n235 B.n234 10.6151
R706 B.n235 B.n84 10.6151
R707 B.n239 B.n84 10.6151
R708 B.n240 B.n239 10.6151
R709 B.n241 B.n240 10.6151
R710 B.n241 B.n82 10.6151
R711 B.n245 B.n82 10.6151
R712 B.n246 B.n245 10.6151
R713 B.n247 B.n246 10.6151
R714 B.n247 B.n80 10.6151
R715 B.n251 B.n80 10.6151
R716 B.n252 B.n251 10.6151
R717 B.n253 B.n252 10.6151
R718 B.n253 B.n78 10.6151
R719 B.n257 B.n78 10.6151
R720 B.n258 B.n257 10.6151
R721 B.n259 B.n258 10.6151
R722 B.n395 B.n30 9.36635
R723 B.n378 B.n377 9.36635
R724 B.n200 B.n199 9.36635
R725 B.n216 B.n90 9.36635
R726 B.n473 B.n0 8.11757
R727 B.n473 B.n1 8.11757
R728 B.n392 B.n30 1.24928
R729 B.n379 B.n378 1.24928
R730 B.n201 B.n200 1.24928
R731 B.n217 B.n216 1.24928
R732 VN VN.t0 164.149
R733 VN VN.t1 123.525
R734 VDD2.n0 VDD2.t0 124.35
R735 VDD2.n0 VDD2.t1 89.4139
R736 VDD2 VDD2.n0 0.657828
C0 VN VP 4.55161f
C1 VP VTAIL 1.68653f
C2 VP B 1.41052f
C3 w_n2082_n2472# VDD1 1.45225f
C4 VDD2 VP 0.326732f
C5 VN VDD1 0.148387f
C6 VDD1 VTAIL 3.85117f
C7 VDD1 B 1.33219f
C8 VDD2 VDD1 0.656092f
C9 w_n2082_n2472# VN 2.77708f
C10 w_n2082_n2472# VTAIL 2.12691f
C11 w_n2082_n2472# B 7.39135f
C12 VDD2 w_n2082_n2472# 1.47634f
C13 VN VTAIL 1.67231f
C14 VN B 0.975642f
C15 VDD2 VN 1.81794f
C16 VTAIL B 2.60344f
C17 VDD2 VTAIL 3.90172f
C18 VDD2 B 1.36094f
C19 VDD1 VP 1.9945f
C20 w_n2082_n2472# VP 3.04196f
C21 VDD2 VSUBS 0.698997f
C22 VDD1 VSUBS 2.91961f
C23 VTAIL VSUBS 0.784f
C24 VN VSUBS 5.4465f
C25 VP VSUBS 1.45367f
C26 B VSUBS 3.421083f
C27 w_n2082_n2472# VSUBS 63.9341f
C28 VDD2.t0 VSUBS 1.05846f
C29 VDD2.t1 VSUBS 0.791042f
C30 VDD2.n0 VSUBS 1.96574f
C31 VN.t1 VSUBS 1.84916f
C32 VN.t0 VSUBS 2.30379f
C33 B.n0 VSUBS 0.006402f
C34 B.n1 VSUBS 0.006402f
C35 B.n2 VSUBS 0.009468f
C36 B.n3 VSUBS 0.007255f
C37 B.n4 VSUBS 0.007255f
C38 B.n5 VSUBS 0.007255f
C39 B.n6 VSUBS 0.007255f
C40 B.n7 VSUBS 0.007255f
C41 B.n8 VSUBS 0.007255f
C42 B.n9 VSUBS 0.007255f
C43 B.n10 VSUBS 0.007255f
C44 B.n11 VSUBS 0.007255f
C45 B.n12 VSUBS 0.007255f
C46 B.n13 VSUBS 0.007255f
C47 B.n14 VSUBS 0.017813f
C48 B.n15 VSUBS 0.007255f
C49 B.n16 VSUBS 0.007255f
C50 B.n17 VSUBS 0.007255f
C51 B.n18 VSUBS 0.007255f
C52 B.n19 VSUBS 0.007255f
C53 B.n20 VSUBS 0.007255f
C54 B.n21 VSUBS 0.007255f
C55 B.n22 VSUBS 0.007255f
C56 B.n23 VSUBS 0.007255f
C57 B.n24 VSUBS 0.007255f
C58 B.n25 VSUBS 0.007255f
C59 B.n26 VSUBS 0.007255f
C60 B.n27 VSUBS 0.007255f
C61 B.t7 VSUBS 0.238007f
C62 B.t8 VSUBS 0.258709f
C63 B.t6 VSUBS 0.890241f
C64 B.n28 VSUBS 0.140377f
C65 B.n29 VSUBS 0.07321f
C66 B.n30 VSUBS 0.01681f
C67 B.n31 VSUBS 0.007255f
C68 B.n32 VSUBS 0.007255f
C69 B.n33 VSUBS 0.007255f
C70 B.n34 VSUBS 0.007255f
C71 B.n35 VSUBS 0.007255f
C72 B.t4 VSUBS 0.238005f
C73 B.t5 VSUBS 0.258707f
C74 B.t3 VSUBS 0.890241f
C75 B.n36 VSUBS 0.140379f
C76 B.n37 VSUBS 0.073212f
C77 B.n38 VSUBS 0.007255f
C78 B.n39 VSUBS 0.007255f
C79 B.n40 VSUBS 0.007255f
C80 B.n41 VSUBS 0.007255f
C81 B.n42 VSUBS 0.007255f
C82 B.n43 VSUBS 0.007255f
C83 B.n44 VSUBS 0.007255f
C84 B.n45 VSUBS 0.007255f
C85 B.n46 VSUBS 0.007255f
C86 B.n47 VSUBS 0.007255f
C87 B.n48 VSUBS 0.007255f
C88 B.n49 VSUBS 0.007255f
C89 B.n50 VSUBS 0.007255f
C90 B.n51 VSUBS 0.017813f
C91 B.n52 VSUBS 0.007255f
C92 B.n53 VSUBS 0.007255f
C93 B.n54 VSUBS 0.007255f
C94 B.n55 VSUBS 0.007255f
C95 B.n56 VSUBS 0.007255f
C96 B.n57 VSUBS 0.007255f
C97 B.n58 VSUBS 0.007255f
C98 B.n59 VSUBS 0.007255f
C99 B.n60 VSUBS 0.007255f
C100 B.n61 VSUBS 0.007255f
C101 B.n62 VSUBS 0.007255f
C102 B.n63 VSUBS 0.007255f
C103 B.n64 VSUBS 0.007255f
C104 B.n65 VSUBS 0.007255f
C105 B.n66 VSUBS 0.007255f
C106 B.n67 VSUBS 0.007255f
C107 B.n68 VSUBS 0.007255f
C108 B.n69 VSUBS 0.007255f
C109 B.n70 VSUBS 0.007255f
C110 B.n71 VSUBS 0.007255f
C111 B.n72 VSUBS 0.007255f
C112 B.n73 VSUBS 0.007255f
C113 B.n74 VSUBS 0.007255f
C114 B.n75 VSUBS 0.007255f
C115 B.n76 VSUBS 0.018209f
C116 B.n77 VSUBS 0.007255f
C117 B.n78 VSUBS 0.007255f
C118 B.n79 VSUBS 0.007255f
C119 B.n80 VSUBS 0.007255f
C120 B.n81 VSUBS 0.007255f
C121 B.n82 VSUBS 0.007255f
C122 B.n83 VSUBS 0.007255f
C123 B.n84 VSUBS 0.007255f
C124 B.n85 VSUBS 0.007255f
C125 B.n86 VSUBS 0.007255f
C126 B.n87 VSUBS 0.007255f
C127 B.n88 VSUBS 0.007255f
C128 B.n89 VSUBS 0.007255f
C129 B.n90 VSUBS 0.006829f
C130 B.n91 VSUBS 0.007255f
C131 B.n92 VSUBS 0.007255f
C132 B.n93 VSUBS 0.007255f
C133 B.n94 VSUBS 0.007255f
C134 B.n95 VSUBS 0.007255f
C135 B.t11 VSUBS 0.238007f
C136 B.t10 VSUBS 0.258709f
C137 B.t9 VSUBS 0.890241f
C138 B.n96 VSUBS 0.140377f
C139 B.n97 VSUBS 0.07321f
C140 B.n98 VSUBS 0.007255f
C141 B.n99 VSUBS 0.007255f
C142 B.n100 VSUBS 0.007255f
C143 B.n101 VSUBS 0.007255f
C144 B.n102 VSUBS 0.007255f
C145 B.n103 VSUBS 0.007255f
C146 B.n104 VSUBS 0.007255f
C147 B.n105 VSUBS 0.007255f
C148 B.n106 VSUBS 0.007255f
C149 B.n107 VSUBS 0.007255f
C150 B.n108 VSUBS 0.007255f
C151 B.n109 VSUBS 0.007255f
C152 B.n110 VSUBS 0.007255f
C153 B.n111 VSUBS 0.017813f
C154 B.n112 VSUBS 0.007255f
C155 B.n113 VSUBS 0.007255f
C156 B.n114 VSUBS 0.007255f
C157 B.n115 VSUBS 0.007255f
C158 B.n116 VSUBS 0.007255f
C159 B.n117 VSUBS 0.007255f
C160 B.n118 VSUBS 0.007255f
C161 B.n119 VSUBS 0.007255f
C162 B.n120 VSUBS 0.007255f
C163 B.n121 VSUBS 0.007255f
C164 B.n122 VSUBS 0.007255f
C165 B.n123 VSUBS 0.007255f
C166 B.n124 VSUBS 0.007255f
C167 B.n125 VSUBS 0.007255f
C168 B.n126 VSUBS 0.007255f
C169 B.n127 VSUBS 0.007255f
C170 B.n128 VSUBS 0.007255f
C171 B.n129 VSUBS 0.007255f
C172 B.n130 VSUBS 0.007255f
C173 B.n131 VSUBS 0.007255f
C174 B.n132 VSUBS 0.007255f
C175 B.n133 VSUBS 0.007255f
C176 B.n134 VSUBS 0.007255f
C177 B.n135 VSUBS 0.007255f
C178 B.n136 VSUBS 0.007255f
C179 B.n137 VSUBS 0.007255f
C180 B.n138 VSUBS 0.007255f
C181 B.n139 VSUBS 0.007255f
C182 B.n140 VSUBS 0.007255f
C183 B.n141 VSUBS 0.007255f
C184 B.n142 VSUBS 0.007255f
C185 B.n143 VSUBS 0.007255f
C186 B.n144 VSUBS 0.007255f
C187 B.n145 VSUBS 0.007255f
C188 B.n146 VSUBS 0.007255f
C189 B.n147 VSUBS 0.007255f
C190 B.n148 VSUBS 0.007255f
C191 B.n149 VSUBS 0.007255f
C192 B.n150 VSUBS 0.007255f
C193 B.n151 VSUBS 0.007255f
C194 B.n152 VSUBS 0.007255f
C195 B.n153 VSUBS 0.007255f
C196 B.n154 VSUBS 0.007255f
C197 B.n155 VSUBS 0.007255f
C198 B.n156 VSUBS 0.017397f
C199 B.n157 VSUBS 0.017397f
C200 B.n158 VSUBS 0.017813f
C201 B.n159 VSUBS 0.007255f
C202 B.n160 VSUBS 0.007255f
C203 B.n161 VSUBS 0.007255f
C204 B.n162 VSUBS 0.007255f
C205 B.n163 VSUBS 0.007255f
C206 B.n164 VSUBS 0.007255f
C207 B.n165 VSUBS 0.007255f
C208 B.n166 VSUBS 0.007255f
C209 B.n167 VSUBS 0.007255f
C210 B.n168 VSUBS 0.007255f
C211 B.n169 VSUBS 0.007255f
C212 B.n170 VSUBS 0.007255f
C213 B.n171 VSUBS 0.007255f
C214 B.n172 VSUBS 0.007255f
C215 B.n173 VSUBS 0.007255f
C216 B.n174 VSUBS 0.007255f
C217 B.n175 VSUBS 0.007255f
C218 B.n176 VSUBS 0.007255f
C219 B.n177 VSUBS 0.007255f
C220 B.n178 VSUBS 0.007255f
C221 B.n179 VSUBS 0.007255f
C222 B.n180 VSUBS 0.007255f
C223 B.n181 VSUBS 0.007255f
C224 B.n182 VSUBS 0.007255f
C225 B.n183 VSUBS 0.007255f
C226 B.n184 VSUBS 0.007255f
C227 B.n185 VSUBS 0.007255f
C228 B.n186 VSUBS 0.007255f
C229 B.n187 VSUBS 0.007255f
C230 B.n188 VSUBS 0.007255f
C231 B.n189 VSUBS 0.007255f
C232 B.n190 VSUBS 0.007255f
C233 B.n191 VSUBS 0.007255f
C234 B.n192 VSUBS 0.007255f
C235 B.n193 VSUBS 0.007255f
C236 B.n194 VSUBS 0.007255f
C237 B.n195 VSUBS 0.007255f
C238 B.n196 VSUBS 0.007255f
C239 B.n197 VSUBS 0.007255f
C240 B.n198 VSUBS 0.007255f
C241 B.n199 VSUBS 0.006829f
C242 B.n200 VSUBS 0.01681f
C243 B.n201 VSUBS 0.004054f
C244 B.n202 VSUBS 0.007255f
C245 B.n203 VSUBS 0.007255f
C246 B.n204 VSUBS 0.007255f
C247 B.n205 VSUBS 0.007255f
C248 B.n206 VSUBS 0.007255f
C249 B.n207 VSUBS 0.007255f
C250 B.n208 VSUBS 0.007255f
C251 B.n209 VSUBS 0.007255f
C252 B.n210 VSUBS 0.007255f
C253 B.n211 VSUBS 0.007255f
C254 B.n212 VSUBS 0.007255f
C255 B.n213 VSUBS 0.007255f
C256 B.t2 VSUBS 0.238005f
C257 B.t1 VSUBS 0.258707f
C258 B.t0 VSUBS 0.890241f
C259 B.n214 VSUBS 0.140379f
C260 B.n215 VSUBS 0.073212f
C261 B.n216 VSUBS 0.01681f
C262 B.n217 VSUBS 0.004054f
C263 B.n218 VSUBS 0.007255f
C264 B.n219 VSUBS 0.007255f
C265 B.n220 VSUBS 0.007255f
C266 B.n221 VSUBS 0.007255f
C267 B.n222 VSUBS 0.007255f
C268 B.n223 VSUBS 0.007255f
C269 B.n224 VSUBS 0.007255f
C270 B.n225 VSUBS 0.007255f
C271 B.n226 VSUBS 0.007255f
C272 B.n227 VSUBS 0.007255f
C273 B.n228 VSUBS 0.007255f
C274 B.n229 VSUBS 0.007255f
C275 B.n230 VSUBS 0.007255f
C276 B.n231 VSUBS 0.007255f
C277 B.n232 VSUBS 0.007255f
C278 B.n233 VSUBS 0.007255f
C279 B.n234 VSUBS 0.007255f
C280 B.n235 VSUBS 0.007255f
C281 B.n236 VSUBS 0.007255f
C282 B.n237 VSUBS 0.007255f
C283 B.n238 VSUBS 0.007255f
C284 B.n239 VSUBS 0.007255f
C285 B.n240 VSUBS 0.007255f
C286 B.n241 VSUBS 0.007255f
C287 B.n242 VSUBS 0.007255f
C288 B.n243 VSUBS 0.007255f
C289 B.n244 VSUBS 0.007255f
C290 B.n245 VSUBS 0.007255f
C291 B.n246 VSUBS 0.007255f
C292 B.n247 VSUBS 0.007255f
C293 B.n248 VSUBS 0.007255f
C294 B.n249 VSUBS 0.007255f
C295 B.n250 VSUBS 0.007255f
C296 B.n251 VSUBS 0.007255f
C297 B.n252 VSUBS 0.007255f
C298 B.n253 VSUBS 0.007255f
C299 B.n254 VSUBS 0.007255f
C300 B.n255 VSUBS 0.007255f
C301 B.n256 VSUBS 0.007255f
C302 B.n257 VSUBS 0.007255f
C303 B.n258 VSUBS 0.007255f
C304 B.n259 VSUBS 0.017001f
C305 B.n260 VSUBS 0.017813f
C306 B.n261 VSUBS 0.017397f
C307 B.n262 VSUBS 0.007255f
C308 B.n263 VSUBS 0.007255f
C309 B.n264 VSUBS 0.007255f
C310 B.n265 VSUBS 0.007255f
C311 B.n266 VSUBS 0.007255f
C312 B.n267 VSUBS 0.007255f
C313 B.n268 VSUBS 0.007255f
C314 B.n269 VSUBS 0.007255f
C315 B.n270 VSUBS 0.007255f
C316 B.n271 VSUBS 0.007255f
C317 B.n272 VSUBS 0.007255f
C318 B.n273 VSUBS 0.007255f
C319 B.n274 VSUBS 0.007255f
C320 B.n275 VSUBS 0.007255f
C321 B.n276 VSUBS 0.007255f
C322 B.n277 VSUBS 0.007255f
C323 B.n278 VSUBS 0.007255f
C324 B.n279 VSUBS 0.007255f
C325 B.n280 VSUBS 0.007255f
C326 B.n281 VSUBS 0.007255f
C327 B.n282 VSUBS 0.007255f
C328 B.n283 VSUBS 0.007255f
C329 B.n284 VSUBS 0.007255f
C330 B.n285 VSUBS 0.007255f
C331 B.n286 VSUBS 0.007255f
C332 B.n287 VSUBS 0.007255f
C333 B.n288 VSUBS 0.007255f
C334 B.n289 VSUBS 0.007255f
C335 B.n290 VSUBS 0.007255f
C336 B.n291 VSUBS 0.007255f
C337 B.n292 VSUBS 0.007255f
C338 B.n293 VSUBS 0.007255f
C339 B.n294 VSUBS 0.007255f
C340 B.n295 VSUBS 0.007255f
C341 B.n296 VSUBS 0.007255f
C342 B.n297 VSUBS 0.007255f
C343 B.n298 VSUBS 0.007255f
C344 B.n299 VSUBS 0.007255f
C345 B.n300 VSUBS 0.007255f
C346 B.n301 VSUBS 0.007255f
C347 B.n302 VSUBS 0.007255f
C348 B.n303 VSUBS 0.007255f
C349 B.n304 VSUBS 0.007255f
C350 B.n305 VSUBS 0.007255f
C351 B.n306 VSUBS 0.007255f
C352 B.n307 VSUBS 0.007255f
C353 B.n308 VSUBS 0.007255f
C354 B.n309 VSUBS 0.007255f
C355 B.n310 VSUBS 0.007255f
C356 B.n311 VSUBS 0.007255f
C357 B.n312 VSUBS 0.007255f
C358 B.n313 VSUBS 0.007255f
C359 B.n314 VSUBS 0.007255f
C360 B.n315 VSUBS 0.007255f
C361 B.n316 VSUBS 0.007255f
C362 B.n317 VSUBS 0.007255f
C363 B.n318 VSUBS 0.007255f
C364 B.n319 VSUBS 0.007255f
C365 B.n320 VSUBS 0.007255f
C366 B.n321 VSUBS 0.007255f
C367 B.n322 VSUBS 0.007255f
C368 B.n323 VSUBS 0.007255f
C369 B.n324 VSUBS 0.007255f
C370 B.n325 VSUBS 0.007255f
C371 B.n326 VSUBS 0.007255f
C372 B.n327 VSUBS 0.007255f
C373 B.n328 VSUBS 0.007255f
C374 B.n329 VSUBS 0.007255f
C375 B.n330 VSUBS 0.007255f
C376 B.n331 VSUBS 0.007255f
C377 B.n332 VSUBS 0.007255f
C378 B.n333 VSUBS 0.007255f
C379 B.n334 VSUBS 0.017397f
C380 B.n335 VSUBS 0.017397f
C381 B.n336 VSUBS 0.017813f
C382 B.n337 VSUBS 0.007255f
C383 B.n338 VSUBS 0.007255f
C384 B.n339 VSUBS 0.007255f
C385 B.n340 VSUBS 0.007255f
C386 B.n341 VSUBS 0.007255f
C387 B.n342 VSUBS 0.007255f
C388 B.n343 VSUBS 0.007255f
C389 B.n344 VSUBS 0.007255f
C390 B.n345 VSUBS 0.007255f
C391 B.n346 VSUBS 0.007255f
C392 B.n347 VSUBS 0.007255f
C393 B.n348 VSUBS 0.007255f
C394 B.n349 VSUBS 0.007255f
C395 B.n350 VSUBS 0.007255f
C396 B.n351 VSUBS 0.007255f
C397 B.n352 VSUBS 0.007255f
C398 B.n353 VSUBS 0.007255f
C399 B.n354 VSUBS 0.007255f
C400 B.n355 VSUBS 0.007255f
C401 B.n356 VSUBS 0.007255f
C402 B.n357 VSUBS 0.007255f
C403 B.n358 VSUBS 0.007255f
C404 B.n359 VSUBS 0.007255f
C405 B.n360 VSUBS 0.007255f
C406 B.n361 VSUBS 0.007255f
C407 B.n362 VSUBS 0.007255f
C408 B.n363 VSUBS 0.007255f
C409 B.n364 VSUBS 0.007255f
C410 B.n365 VSUBS 0.007255f
C411 B.n366 VSUBS 0.007255f
C412 B.n367 VSUBS 0.007255f
C413 B.n368 VSUBS 0.007255f
C414 B.n369 VSUBS 0.007255f
C415 B.n370 VSUBS 0.007255f
C416 B.n371 VSUBS 0.007255f
C417 B.n372 VSUBS 0.007255f
C418 B.n373 VSUBS 0.007255f
C419 B.n374 VSUBS 0.007255f
C420 B.n375 VSUBS 0.007255f
C421 B.n376 VSUBS 0.007255f
C422 B.n377 VSUBS 0.006829f
C423 B.n378 VSUBS 0.01681f
C424 B.n379 VSUBS 0.004054f
C425 B.n380 VSUBS 0.007255f
C426 B.n381 VSUBS 0.007255f
C427 B.n382 VSUBS 0.007255f
C428 B.n383 VSUBS 0.007255f
C429 B.n384 VSUBS 0.007255f
C430 B.n385 VSUBS 0.007255f
C431 B.n386 VSUBS 0.007255f
C432 B.n387 VSUBS 0.007255f
C433 B.n388 VSUBS 0.007255f
C434 B.n389 VSUBS 0.007255f
C435 B.n390 VSUBS 0.007255f
C436 B.n391 VSUBS 0.007255f
C437 B.n392 VSUBS 0.004054f
C438 B.n393 VSUBS 0.007255f
C439 B.n394 VSUBS 0.007255f
C440 B.n395 VSUBS 0.006829f
C441 B.n396 VSUBS 0.007255f
C442 B.n397 VSUBS 0.007255f
C443 B.n398 VSUBS 0.007255f
C444 B.n399 VSUBS 0.007255f
C445 B.n400 VSUBS 0.007255f
C446 B.n401 VSUBS 0.007255f
C447 B.n402 VSUBS 0.007255f
C448 B.n403 VSUBS 0.007255f
C449 B.n404 VSUBS 0.007255f
C450 B.n405 VSUBS 0.007255f
C451 B.n406 VSUBS 0.007255f
C452 B.n407 VSUBS 0.007255f
C453 B.n408 VSUBS 0.007255f
C454 B.n409 VSUBS 0.007255f
C455 B.n410 VSUBS 0.007255f
C456 B.n411 VSUBS 0.007255f
C457 B.n412 VSUBS 0.007255f
C458 B.n413 VSUBS 0.007255f
C459 B.n414 VSUBS 0.007255f
C460 B.n415 VSUBS 0.007255f
C461 B.n416 VSUBS 0.007255f
C462 B.n417 VSUBS 0.007255f
C463 B.n418 VSUBS 0.007255f
C464 B.n419 VSUBS 0.007255f
C465 B.n420 VSUBS 0.007255f
C466 B.n421 VSUBS 0.007255f
C467 B.n422 VSUBS 0.007255f
C468 B.n423 VSUBS 0.007255f
C469 B.n424 VSUBS 0.007255f
C470 B.n425 VSUBS 0.007255f
C471 B.n426 VSUBS 0.007255f
C472 B.n427 VSUBS 0.007255f
C473 B.n428 VSUBS 0.007255f
C474 B.n429 VSUBS 0.007255f
C475 B.n430 VSUBS 0.007255f
C476 B.n431 VSUBS 0.007255f
C477 B.n432 VSUBS 0.007255f
C478 B.n433 VSUBS 0.007255f
C479 B.n434 VSUBS 0.007255f
C480 B.n435 VSUBS 0.017813f
C481 B.n436 VSUBS 0.017397f
C482 B.n437 VSUBS 0.017397f
C483 B.n438 VSUBS 0.007255f
C484 B.n439 VSUBS 0.007255f
C485 B.n440 VSUBS 0.007255f
C486 B.n441 VSUBS 0.007255f
C487 B.n442 VSUBS 0.007255f
C488 B.n443 VSUBS 0.007255f
C489 B.n444 VSUBS 0.007255f
C490 B.n445 VSUBS 0.007255f
C491 B.n446 VSUBS 0.007255f
C492 B.n447 VSUBS 0.007255f
C493 B.n448 VSUBS 0.007255f
C494 B.n449 VSUBS 0.007255f
C495 B.n450 VSUBS 0.007255f
C496 B.n451 VSUBS 0.007255f
C497 B.n452 VSUBS 0.007255f
C498 B.n453 VSUBS 0.007255f
C499 B.n454 VSUBS 0.007255f
C500 B.n455 VSUBS 0.007255f
C501 B.n456 VSUBS 0.007255f
C502 B.n457 VSUBS 0.007255f
C503 B.n458 VSUBS 0.007255f
C504 B.n459 VSUBS 0.007255f
C505 B.n460 VSUBS 0.007255f
C506 B.n461 VSUBS 0.007255f
C507 B.n462 VSUBS 0.007255f
C508 B.n463 VSUBS 0.007255f
C509 B.n464 VSUBS 0.007255f
C510 B.n465 VSUBS 0.007255f
C511 B.n466 VSUBS 0.007255f
C512 B.n467 VSUBS 0.007255f
C513 B.n468 VSUBS 0.007255f
C514 B.n469 VSUBS 0.007255f
C515 B.n470 VSUBS 0.007255f
C516 B.n471 VSUBS 0.009468f
C517 B.n472 VSUBS 0.010086f
C518 B.n473 VSUBS 0.020056f
C519 VDD1.t1 VSUBS 0.782821f
C520 VDD1.t0 VSUBS 1.06342f
C521 VTAIL.t3 VSUBS 1.28853f
C522 VTAIL.n0 VSUBS 1.88927f
C523 VTAIL.t0 VSUBS 1.28853f
C524 VTAIL.n1 VSUBS 1.93271f
C525 VTAIL.t2 VSUBS 1.28853f
C526 VTAIL.n2 VSUBS 1.74022f
C527 VTAIL.t1 VSUBS 1.28853f
C528 VTAIL.n3 VSUBS 1.64969f
C529 VP.t0 VSUBS 2.37637f
C530 VP.t1 VSUBS 1.90882f
C531 VP.n0 VSUBS 3.24199f
.ends

