* NGSPICE file created from diff_pair_sample_0061.ext - technology: sky130A

.subckt diff_pair_sample_0061 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=0 ps=0 w=19.72 l=0.5
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=7.6908 ps=40.22 w=19.72 l=0.5
X2 B.t8 B.t6 B.t7 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=0 ps=0 w=19.72 l=0.5
X3 VDD1.t0 VP.t1 VTAIL.t3 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=7.6908 ps=40.22 w=19.72 l=0.5
X4 B.t5 B.t3 B.t4 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=0 ps=0 w=19.72 l=0.5
X5 VDD2.t1 VN.t0 VTAIL.t0 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=7.6908 ps=40.22 w=19.72 l=0.5
X6 B.t2 B.t0 B.t1 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=0 ps=0 w=19.72 l=0.5
X7 VDD2.t0 VN.t1 VTAIL.t1 w_n1302_n4916# sky130_fd_pr__pfet_01v8 ad=7.6908 pd=40.22 as=7.6908 ps=40.22 w=19.72 l=0.5
R0 B.n129 B.t6 1156.91
R1 B.n135 B.t0 1156.91
R2 B.n42 B.t9 1156.91
R3 B.n49 B.t3 1156.91
R4 B.n443 B.n82 585
R5 B.n445 B.n444 585
R6 B.n446 B.n81 585
R7 B.n448 B.n447 585
R8 B.n449 B.n80 585
R9 B.n451 B.n450 585
R10 B.n452 B.n79 585
R11 B.n454 B.n453 585
R12 B.n455 B.n78 585
R13 B.n457 B.n456 585
R14 B.n458 B.n77 585
R15 B.n460 B.n459 585
R16 B.n461 B.n76 585
R17 B.n463 B.n462 585
R18 B.n464 B.n75 585
R19 B.n466 B.n465 585
R20 B.n467 B.n74 585
R21 B.n469 B.n468 585
R22 B.n470 B.n73 585
R23 B.n472 B.n471 585
R24 B.n473 B.n72 585
R25 B.n475 B.n474 585
R26 B.n476 B.n71 585
R27 B.n478 B.n477 585
R28 B.n479 B.n70 585
R29 B.n481 B.n480 585
R30 B.n482 B.n69 585
R31 B.n484 B.n483 585
R32 B.n485 B.n68 585
R33 B.n487 B.n486 585
R34 B.n488 B.n67 585
R35 B.n490 B.n489 585
R36 B.n491 B.n66 585
R37 B.n493 B.n492 585
R38 B.n494 B.n65 585
R39 B.n496 B.n495 585
R40 B.n497 B.n64 585
R41 B.n499 B.n498 585
R42 B.n500 B.n63 585
R43 B.n502 B.n501 585
R44 B.n503 B.n62 585
R45 B.n505 B.n504 585
R46 B.n506 B.n61 585
R47 B.n508 B.n507 585
R48 B.n509 B.n60 585
R49 B.n511 B.n510 585
R50 B.n512 B.n59 585
R51 B.n514 B.n513 585
R52 B.n515 B.n58 585
R53 B.n517 B.n516 585
R54 B.n518 B.n57 585
R55 B.n520 B.n519 585
R56 B.n521 B.n56 585
R57 B.n523 B.n522 585
R58 B.n524 B.n55 585
R59 B.n526 B.n525 585
R60 B.n527 B.n54 585
R61 B.n529 B.n528 585
R62 B.n530 B.n53 585
R63 B.n532 B.n531 585
R64 B.n533 B.n52 585
R65 B.n535 B.n534 585
R66 B.n536 B.n51 585
R67 B.n538 B.n537 585
R68 B.n540 B.n48 585
R69 B.n542 B.n541 585
R70 B.n543 B.n47 585
R71 B.n545 B.n544 585
R72 B.n546 B.n46 585
R73 B.n548 B.n547 585
R74 B.n549 B.n45 585
R75 B.n551 B.n550 585
R76 B.n552 B.n41 585
R77 B.n554 B.n553 585
R78 B.n555 B.n40 585
R79 B.n557 B.n556 585
R80 B.n558 B.n39 585
R81 B.n560 B.n559 585
R82 B.n561 B.n38 585
R83 B.n563 B.n562 585
R84 B.n564 B.n37 585
R85 B.n566 B.n565 585
R86 B.n567 B.n36 585
R87 B.n569 B.n568 585
R88 B.n570 B.n35 585
R89 B.n572 B.n571 585
R90 B.n573 B.n34 585
R91 B.n575 B.n574 585
R92 B.n576 B.n33 585
R93 B.n578 B.n577 585
R94 B.n579 B.n32 585
R95 B.n581 B.n580 585
R96 B.n582 B.n31 585
R97 B.n584 B.n583 585
R98 B.n585 B.n30 585
R99 B.n587 B.n586 585
R100 B.n588 B.n29 585
R101 B.n590 B.n589 585
R102 B.n591 B.n28 585
R103 B.n593 B.n592 585
R104 B.n594 B.n27 585
R105 B.n596 B.n595 585
R106 B.n597 B.n26 585
R107 B.n599 B.n598 585
R108 B.n600 B.n25 585
R109 B.n602 B.n601 585
R110 B.n603 B.n24 585
R111 B.n605 B.n604 585
R112 B.n606 B.n23 585
R113 B.n608 B.n607 585
R114 B.n609 B.n22 585
R115 B.n611 B.n610 585
R116 B.n612 B.n21 585
R117 B.n614 B.n613 585
R118 B.n615 B.n20 585
R119 B.n617 B.n616 585
R120 B.n618 B.n19 585
R121 B.n620 B.n619 585
R122 B.n621 B.n18 585
R123 B.n623 B.n622 585
R124 B.n624 B.n17 585
R125 B.n626 B.n625 585
R126 B.n627 B.n16 585
R127 B.n629 B.n628 585
R128 B.n630 B.n15 585
R129 B.n632 B.n631 585
R130 B.n633 B.n14 585
R131 B.n635 B.n634 585
R132 B.n636 B.n13 585
R133 B.n638 B.n637 585
R134 B.n639 B.n12 585
R135 B.n641 B.n640 585
R136 B.n642 B.n11 585
R137 B.n644 B.n643 585
R138 B.n645 B.n10 585
R139 B.n647 B.n646 585
R140 B.n648 B.n9 585
R141 B.n650 B.n649 585
R142 B.n442 B.n441 585
R143 B.n440 B.n83 585
R144 B.n439 B.n438 585
R145 B.n437 B.n84 585
R146 B.n436 B.n435 585
R147 B.n434 B.n85 585
R148 B.n433 B.n432 585
R149 B.n431 B.n86 585
R150 B.n430 B.n429 585
R151 B.n428 B.n87 585
R152 B.n427 B.n426 585
R153 B.n425 B.n88 585
R154 B.n424 B.n423 585
R155 B.n422 B.n89 585
R156 B.n421 B.n420 585
R157 B.n419 B.n90 585
R158 B.n418 B.n417 585
R159 B.n416 B.n91 585
R160 B.n415 B.n414 585
R161 B.n413 B.n92 585
R162 B.n412 B.n411 585
R163 B.n410 B.n93 585
R164 B.n409 B.n408 585
R165 B.n407 B.n94 585
R166 B.n406 B.n405 585
R167 B.n404 B.n95 585
R168 B.n403 B.n402 585
R169 B.n194 B.n169 585
R170 B.n196 B.n195 585
R171 B.n197 B.n168 585
R172 B.n199 B.n198 585
R173 B.n200 B.n167 585
R174 B.n202 B.n201 585
R175 B.n203 B.n166 585
R176 B.n205 B.n204 585
R177 B.n206 B.n165 585
R178 B.n208 B.n207 585
R179 B.n209 B.n164 585
R180 B.n211 B.n210 585
R181 B.n212 B.n163 585
R182 B.n214 B.n213 585
R183 B.n215 B.n162 585
R184 B.n217 B.n216 585
R185 B.n218 B.n161 585
R186 B.n220 B.n219 585
R187 B.n221 B.n160 585
R188 B.n223 B.n222 585
R189 B.n224 B.n159 585
R190 B.n226 B.n225 585
R191 B.n227 B.n158 585
R192 B.n229 B.n228 585
R193 B.n230 B.n157 585
R194 B.n232 B.n231 585
R195 B.n233 B.n156 585
R196 B.n235 B.n234 585
R197 B.n236 B.n155 585
R198 B.n238 B.n237 585
R199 B.n239 B.n154 585
R200 B.n241 B.n240 585
R201 B.n242 B.n153 585
R202 B.n244 B.n243 585
R203 B.n245 B.n152 585
R204 B.n247 B.n246 585
R205 B.n248 B.n151 585
R206 B.n250 B.n249 585
R207 B.n251 B.n150 585
R208 B.n253 B.n252 585
R209 B.n254 B.n149 585
R210 B.n256 B.n255 585
R211 B.n257 B.n148 585
R212 B.n259 B.n258 585
R213 B.n260 B.n147 585
R214 B.n262 B.n261 585
R215 B.n263 B.n146 585
R216 B.n265 B.n264 585
R217 B.n266 B.n145 585
R218 B.n268 B.n267 585
R219 B.n269 B.n144 585
R220 B.n271 B.n270 585
R221 B.n272 B.n143 585
R222 B.n274 B.n273 585
R223 B.n275 B.n142 585
R224 B.n277 B.n276 585
R225 B.n278 B.n141 585
R226 B.n280 B.n279 585
R227 B.n281 B.n140 585
R228 B.n283 B.n282 585
R229 B.n284 B.n139 585
R230 B.n286 B.n285 585
R231 B.n287 B.n138 585
R232 B.n289 B.n288 585
R233 B.n291 B.n290 585
R234 B.n292 B.n134 585
R235 B.n294 B.n293 585
R236 B.n295 B.n133 585
R237 B.n297 B.n296 585
R238 B.n298 B.n132 585
R239 B.n300 B.n299 585
R240 B.n301 B.n131 585
R241 B.n303 B.n302 585
R242 B.n304 B.n128 585
R243 B.n307 B.n306 585
R244 B.n308 B.n127 585
R245 B.n310 B.n309 585
R246 B.n311 B.n126 585
R247 B.n313 B.n312 585
R248 B.n314 B.n125 585
R249 B.n316 B.n315 585
R250 B.n317 B.n124 585
R251 B.n319 B.n318 585
R252 B.n320 B.n123 585
R253 B.n322 B.n321 585
R254 B.n323 B.n122 585
R255 B.n325 B.n324 585
R256 B.n326 B.n121 585
R257 B.n328 B.n327 585
R258 B.n329 B.n120 585
R259 B.n331 B.n330 585
R260 B.n332 B.n119 585
R261 B.n334 B.n333 585
R262 B.n335 B.n118 585
R263 B.n337 B.n336 585
R264 B.n338 B.n117 585
R265 B.n340 B.n339 585
R266 B.n341 B.n116 585
R267 B.n343 B.n342 585
R268 B.n344 B.n115 585
R269 B.n346 B.n345 585
R270 B.n347 B.n114 585
R271 B.n349 B.n348 585
R272 B.n350 B.n113 585
R273 B.n352 B.n351 585
R274 B.n353 B.n112 585
R275 B.n355 B.n354 585
R276 B.n356 B.n111 585
R277 B.n358 B.n357 585
R278 B.n359 B.n110 585
R279 B.n361 B.n360 585
R280 B.n362 B.n109 585
R281 B.n364 B.n363 585
R282 B.n365 B.n108 585
R283 B.n367 B.n366 585
R284 B.n368 B.n107 585
R285 B.n370 B.n369 585
R286 B.n371 B.n106 585
R287 B.n373 B.n372 585
R288 B.n374 B.n105 585
R289 B.n376 B.n375 585
R290 B.n377 B.n104 585
R291 B.n379 B.n378 585
R292 B.n380 B.n103 585
R293 B.n382 B.n381 585
R294 B.n383 B.n102 585
R295 B.n385 B.n384 585
R296 B.n386 B.n101 585
R297 B.n388 B.n387 585
R298 B.n389 B.n100 585
R299 B.n391 B.n390 585
R300 B.n392 B.n99 585
R301 B.n394 B.n393 585
R302 B.n395 B.n98 585
R303 B.n397 B.n396 585
R304 B.n398 B.n97 585
R305 B.n400 B.n399 585
R306 B.n401 B.n96 585
R307 B.n193 B.n192 585
R308 B.n191 B.n170 585
R309 B.n190 B.n189 585
R310 B.n188 B.n171 585
R311 B.n187 B.n186 585
R312 B.n185 B.n172 585
R313 B.n184 B.n183 585
R314 B.n182 B.n173 585
R315 B.n181 B.n180 585
R316 B.n179 B.n174 585
R317 B.n178 B.n177 585
R318 B.n176 B.n175 585
R319 B.n2 B.n0 585
R320 B.n669 B.n1 585
R321 B.n668 B.n667 585
R322 B.n666 B.n3 585
R323 B.n665 B.n664 585
R324 B.n663 B.n4 585
R325 B.n662 B.n661 585
R326 B.n660 B.n5 585
R327 B.n659 B.n658 585
R328 B.n657 B.n6 585
R329 B.n656 B.n655 585
R330 B.n654 B.n7 585
R331 B.n653 B.n652 585
R332 B.n651 B.n8 585
R333 B.n671 B.n670 585
R334 B.n129 B.t8 531.01
R335 B.n49 B.t4 531.01
R336 B.n135 B.t2 531.01
R337 B.n42 B.t10 531.01
R338 B.n194 B.n193 526.135
R339 B.n651 B.n650 526.135
R340 B.n403 B.n96 526.135
R341 B.n441 B.n82 526.135
R342 B.n130 B.t7 514.913
R343 B.n50 B.t5 514.913
R344 B.n136 B.t1 514.913
R345 B.n43 B.t11 514.913
R346 B.n193 B.n170 163.367
R347 B.n189 B.n170 163.367
R348 B.n189 B.n188 163.367
R349 B.n188 B.n187 163.367
R350 B.n187 B.n172 163.367
R351 B.n183 B.n172 163.367
R352 B.n183 B.n182 163.367
R353 B.n182 B.n181 163.367
R354 B.n181 B.n174 163.367
R355 B.n177 B.n174 163.367
R356 B.n177 B.n176 163.367
R357 B.n176 B.n2 163.367
R358 B.n670 B.n2 163.367
R359 B.n670 B.n669 163.367
R360 B.n669 B.n668 163.367
R361 B.n668 B.n3 163.367
R362 B.n664 B.n3 163.367
R363 B.n664 B.n663 163.367
R364 B.n663 B.n662 163.367
R365 B.n662 B.n5 163.367
R366 B.n658 B.n5 163.367
R367 B.n658 B.n657 163.367
R368 B.n657 B.n656 163.367
R369 B.n656 B.n7 163.367
R370 B.n652 B.n7 163.367
R371 B.n652 B.n651 163.367
R372 B.n195 B.n194 163.367
R373 B.n195 B.n168 163.367
R374 B.n199 B.n168 163.367
R375 B.n200 B.n199 163.367
R376 B.n201 B.n200 163.367
R377 B.n201 B.n166 163.367
R378 B.n205 B.n166 163.367
R379 B.n206 B.n205 163.367
R380 B.n207 B.n206 163.367
R381 B.n207 B.n164 163.367
R382 B.n211 B.n164 163.367
R383 B.n212 B.n211 163.367
R384 B.n213 B.n212 163.367
R385 B.n213 B.n162 163.367
R386 B.n217 B.n162 163.367
R387 B.n218 B.n217 163.367
R388 B.n219 B.n218 163.367
R389 B.n219 B.n160 163.367
R390 B.n223 B.n160 163.367
R391 B.n224 B.n223 163.367
R392 B.n225 B.n224 163.367
R393 B.n225 B.n158 163.367
R394 B.n229 B.n158 163.367
R395 B.n230 B.n229 163.367
R396 B.n231 B.n230 163.367
R397 B.n231 B.n156 163.367
R398 B.n235 B.n156 163.367
R399 B.n236 B.n235 163.367
R400 B.n237 B.n236 163.367
R401 B.n237 B.n154 163.367
R402 B.n241 B.n154 163.367
R403 B.n242 B.n241 163.367
R404 B.n243 B.n242 163.367
R405 B.n243 B.n152 163.367
R406 B.n247 B.n152 163.367
R407 B.n248 B.n247 163.367
R408 B.n249 B.n248 163.367
R409 B.n249 B.n150 163.367
R410 B.n253 B.n150 163.367
R411 B.n254 B.n253 163.367
R412 B.n255 B.n254 163.367
R413 B.n255 B.n148 163.367
R414 B.n259 B.n148 163.367
R415 B.n260 B.n259 163.367
R416 B.n261 B.n260 163.367
R417 B.n261 B.n146 163.367
R418 B.n265 B.n146 163.367
R419 B.n266 B.n265 163.367
R420 B.n267 B.n266 163.367
R421 B.n267 B.n144 163.367
R422 B.n271 B.n144 163.367
R423 B.n272 B.n271 163.367
R424 B.n273 B.n272 163.367
R425 B.n273 B.n142 163.367
R426 B.n277 B.n142 163.367
R427 B.n278 B.n277 163.367
R428 B.n279 B.n278 163.367
R429 B.n279 B.n140 163.367
R430 B.n283 B.n140 163.367
R431 B.n284 B.n283 163.367
R432 B.n285 B.n284 163.367
R433 B.n285 B.n138 163.367
R434 B.n289 B.n138 163.367
R435 B.n290 B.n289 163.367
R436 B.n290 B.n134 163.367
R437 B.n294 B.n134 163.367
R438 B.n295 B.n294 163.367
R439 B.n296 B.n295 163.367
R440 B.n296 B.n132 163.367
R441 B.n300 B.n132 163.367
R442 B.n301 B.n300 163.367
R443 B.n302 B.n301 163.367
R444 B.n302 B.n128 163.367
R445 B.n307 B.n128 163.367
R446 B.n308 B.n307 163.367
R447 B.n309 B.n308 163.367
R448 B.n309 B.n126 163.367
R449 B.n313 B.n126 163.367
R450 B.n314 B.n313 163.367
R451 B.n315 B.n314 163.367
R452 B.n315 B.n124 163.367
R453 B.n319 B.n124 163.367
R454 B.n320 B.n319 163.367
R455 B.n321 B.n320 163.367
R456 B.n321 B.n122 163.367
R457 B.n325 B.n122 163.367
R458 B.n326 B.n325 163.367
R459 B.n327 B.n326 163.367
R460 B.n327 B.n120 163.367
R461 B.n331 B.n120 163.367
R462 B.n332 B.n331 163.367
R463 B.n333 B.n332 163.367
R464 B.n333 B.n118 163.367
R465 B.n337 B.n118 163.367
R466 B.n338 B.n337 163.367
R467 B.n339 B.n338 163.367
R468 B.n339 B.n116 163.367
R469 B.n343 B.n116 163.367
R470 B.n344 B.n343 163.367
R471 B.n345 B.n344 163.367
R472 B.n345 B.n114 163.367
R473 B.n349 B.n114 163.367
R474 B.n350 B.n349 163.367
R475 B.n351 B.n350 163.367
R476 B.n351 B.n112 163.367
R477 B.n355 B.n112 163.367
R478 B.n356 B.n355 163.367
R479 B.n357 B.n356 163.367
R480 B.n357 B.n110 163.367
R481 B.n361 B.n110 163.367
R482 B.n362 B.n361 163.367
R483 B.n363 B.n362 163.367
R484 B.n363 B.n108 163.367
R485 B.n367 B.n108 163.367
R486 B.n368 B.n367 163.367
R487 B.n369 B.n368 163.367
R488 B.n369 B.n106 163.367
R489 B.n373 B.n106 163.367
R490 B.n374 B.n373 163.367
R491 B.n375 B.n374 163.367
R492 B.n375 B.n104 163.367
R493 B.n379 B.n104 163.367
R494 B.n380 B.n379 163.367
R495 B.n381 B.n380 163.367
R496 B.n381 B.n102 163.367
R497 B.n385 B.n102 163.367
R498 B.n386 B.n385 163.367
R499 B.n387 B.n386 163.367
R500 B.n387 B.n100 163.367
R501 B.n391 B.n100 163.367
R502 B.n392 B.n391 163.367
R503 B.n393 B.n392 163.367
R504 B.n393 B.n98 163.367
R505 B.n397 B.n98 163.367
R506 B.n398 B.n397 163.367
R507 B.n399 B.n398 163.367
R508 B.n399 B.n96 163.367
R509 B.n404 B.n403 163.367
R510 B.n405 B.n404 163.367
R511 B.n405 B.n94 163.367
R512 B.n409 B.n94 163.367
R513 B.n410 B.n409 163.367
R514 B.n411 B.n410 163.367
R515 B.n411 B.n92 163.367
R516 B.n415 B.n92 163.367
R517 B.n416 B.n415 163.367
R518 B.n417 B.n416 163.367
R519 B.n417 B.n90 163.367
R520 B.n421 B.n90 163.367
R521 B.n422 B.n421 163.367
R522 B.n423 B.n422 163.367
R523 B.n423 B.n88 163.367
R524 B.n427 B.n88 163.367
R525 B.n428 B.n427 163.367
R526 B.n429 B.n428 163.367
R527 B.n429 B.n86 163.367
R528 B.n433 B.n86 163.367
R529 B.n434 B.n433 163.367
R530 B.n435 B.n434 163.367
R531 B.n435 B.n84 163.367
R532 B.n439 B.n84 163.367
R533 B.n440 B.n439 163.367
R534 B.n441 B.n440 163.367
R535 B.n650 B.n9 163.367
R536 B.n646 B.n9 163.367
R537 B.n646 B.n645 163.367
R538 B.n645 B.n644 163.367
R539 B.n644 B.n11 163.367
R540 B.n640 B.n11 163.367
R541 B.n640 B.n639 163.367
R542 B.n639 B.n638 163.367
R543 B.n638 B.n13 163.367
R544 B.n634 B.n13 163.367
R545 B.n634 B.n633 163.367
R546 B.n633 B.n632 163.367
R547 B.n632 B.n15 163.367
R548 B.n628 B.n15 163.367
R549 B.n628 B.n627 163.367
R550 B.n627 B.n626 163.367
R551 B.n626 B.n17 163.367
R552 B.n622 B.n17 163.367
R553 B.n622 B.n621 163.367
R554 B.n621 B.n620 163.367
R555 B.n620 B.n19 163.367
R556 B.n616 B.n19 163.367
R557 B.n616 B.n615 163.367
R558 B.n615 B.n614 163.367
R559 B.n614 B.n21 163.367
R560 B.n610 B.n21 163.367
R561 B.n610 B.n609 163.367
R562 B.n609 B.n608 163.367
R563 B.n608 B.n23 163.367
R564 B.n604 B.n23 163.367
R565 B.n604 B.n603 163.367
R566 B.n603 B.n602 163.367
R567 B.n602 B.n25 163.367
R568 B.n598 B.n25 163.367
R569 B.n598 B.n597 163.367
R570 B.n597 B.n596 163.367
R571 B.n596 B.n27 163.367
R572 B.n592 B.n27 163.367
R573 B.n592 B.n591 163.367
R574 B.n591 B.n590 163.367
R575 B.n590 B.n29 163.367
R576 B.n586 B.n29 163.367
R577 B.n586 B.n585 163.367
R578 B.n585 B.n584 163.367
R579 B.n584 B.n31 163.367
R580 B.n580 B.n31 163.367
R581 B.n580 B.n579 163.367
R582 B.n579 B.n578 163.367
R583 B.n578 B.n33 163.367
R584 B.n574 B.n33 163.367
R585 B.n574 B.n573 163.367
R586 B.n573 B.n572 163.367
R587 B.n572 B.n35 163.367
R588 B.n568 B.n35 163.367
R589 B.n568 B.n567 163.367
R590 B.n567 B.n566 163.367
R591 B.n566 B.n37 163.367
R592 B.n562 B.n37 163.367
R593 B.n562 B.n561 163.367
R594 B.n561 B.n560 163.367
R595 B.n560 B.n39 163.367
R596 B.n556 B.n39 163.367
R597 B.n556 B.n555 163.367
R598 B.n555 B.n554 163.367
R599 B.n554 B.n41 163.367
R600 B.n550 B.n41 163.367
R601 B.n550 B.n549 163.367
R602 B.n549 B.n548 163.367
R603 B.n548 B.n46 163.367
R604 B.n544 B.n46 163.367
R605 B.n544 B.n543 163.367
R606 B.n543 B.n542 163.367
R607 B.n542 B.n48 163.367
R608 B.n537 B.n48 163.367
R609 B.n537 B.n536 163.367
R610 B.n536 B.n535 163.367
R611 B.n535 B.n52 163.367
R612 B.n531 B.n52 163.367
R613 B.n531 B.n530 163.367
R614 B.n530 B.n529 163.367
R615 B.n529 B.n54 163.367
R616 B.n525 B.n54 163.367
R617 B.n525 B.n524 163.367
R618 B.n524 B.n523 163.367
R619 B.n523 B.n56 163.367
R620 B.n519 B.n56 163.367
R621 B.n519 B.n518 163.367
R622 B.n518 B.n517 163.367
R623 B.n517 B.n58 163.367
R624 B.n513 B.n58 163.367
R625 B.n513 B.n512 163.367
R626 B.n512 B.n511 163.367
R627 B.n511 B.n60 163.367
R628 B.n507 B.n60 163.367
R629 B.n507 B.n506 163.367
R630 B.n506 B.n505 163.367
R631 B.n505 B.n62 163.367
R632 B.n501 B.n62 163.367
R633 B.n501 B.n500 163.367
R634 B.n500 B.n499 163.367
R635 B.n499 B.n64 163.367
R636 B.n495 B.n64 163.367
R637 B.n495 B.n494 163.367
R638 B.n494 B.n493 163.367
R639 B.n493 B.n66 163.367
R640 B.n489 B.n66 163.367
R641 B.n489 B.n488 163.367
R642 B.n488 B.n487 163.367
R643 B.n487 B.n68 163.367
R644 B.n483 B.n68 163.367
R645 B.n483 B.n482 163.367
R646 B.n482 B.n481 163.367
R647 B.n481 B.n70 163.367
R648 B.n477 B.n70 163.367
R649 B.n477 B.n476 163.367
R650 B.n476 B.n475 163.367
R651 B.n475 B.n72 163.367
R652 B.n471 B.n72 163.367
R653 B.n471 B.n470 163.367
R654 B.n470 B.n469 163.367
R655 B.n469 B.n74 163.367
R656 B.n465 B.n74 163.367
R657 B.n465 B.n464 163.367
R658 B.n464 B.n463 163.367
R659 B.n463 B.n76 163.367
R660 B.n459 B.n76 163.367
R661 B.n459 B.n458 163.367
R662 B.n458 B.n457 163.367
R663 B.n457 B.n78 163.367
R664 B.n453 B.n78 163.367
R665 B.n453 B.n452 163.367
R666 B.n452 B.n451 163.367
R667 B.n451 B.n80 163.367
R668 B.n447 B.n80 163.367
R669 B.n447 B.n446 163.367
R670 B.n446 B.n445 163.367
R671 B.n445 B.n82 163.367
R672 B.n305 B.n130 59.5399
R673 B.n137 B.n136 59.5399
R674 B.n44 B.n43 59.5399
R675 B.n539 B.n50 59.5399
R676 B.n649 B.n8 34.1859
R677 B.n443 B.n442 34.1859
R678 B.n402 B.n401 34.1859
R679 B.n192 B.n169 34.1859
R680 B B.n671 18.0485
R681 B.n130 B.n129 16.0975
R682 B.n136 B.n135 16.0975
R683 B.n43 B.n42 16.0975
R684 B.n50 B.n49 16.0975
R685 B.n649 B.n648 10.6151
R686 B.n648 B.n647 10.6151
R687 B.n647 B.n10 10.6151
R688 B.n643 B.n10 10.6151
R689 B.n643 B.n642 10.6151
R690 B.n642 B.n641 10.6151
R691 B.n641 B.n12 10.6151
R692 B.n637 B.n12 10.6151
R693 B.n637 B.n636 10.6151
R694 B.n636 B.n635 10.6151
R695 B.n635 B.n14 10.6151
R696 B.n631 B.n14 10.6151
R697 B.n631 B.n630 10.6151
R698 B.n630 B.n629 10.6151
R699 B.n629 B.n16 10.6151
R700 B.n625 B.n16 10.6151
R701 B.n625 B.n624 10.6151
R702 B.n624 B.n623 10.6151
R703 B.n623 B.n18 10.6151
R704 B.n619 B.n18 10.6151
R705 B.n619 B.n618 10.6151
R706 B.n618 B.n617 10.6151
R707 B.n617 B.n20 10.6151
R708 B.n613 B.n20 10.6151
R709 B.n613 B.n612 10.6151
R710 B.n612 B.n611 10.6151
R711 B.n611 B.n22 10.6151
R712 B.n607 B.n22 10.6151
R713 B.n607 B.n606 10.6151
R714 B.n606 B.n605 10.6151
R715 B.n605 B.n24 10.6151
R716 B.n601 B.n24 10.6151
R717 B.n601 B.n600 10.6151
R718 B.n600 B.n599 10.6151
R719 B.n599 B.n26 10.6151
R720 B.n595 B.n26 10.6151
R721 B.n595 B.n594 10.6151
R722 B.n594 B.n593 10.6151
R723 B.n593 B.n28 10.6151
R724 B.n589 B.n28 10.6151
R725 B.n589 B.n588 10.6151
R726 B.n588 B.n587 10.6151
R727 B.n587 B.n30 10.6151
R728 B.n583 B.n30 10.6151
R729 B.n583 B.n582 10.6151
R730 B.n582 B.n581 10.6151
R731 B.n581 B.n32 10.6151
R732 B.n577 B.n32 10.6151
R733 B.n577 B.n576 10.6151
R734 B.n576 B.n575 10.6151
R735 B.n575 B.n34 10.6151
R736 B.n571 B.n34 10.6151
R737 B.n571 B.n570 10.6151
R738 B.n570 B.n569 10.6151
R739 B.n569 B.n36 10.6151
R740 B.n565 B.n36 10.6151
R741 B.n565 B.n564 10.6151
R742 B.n564 B.n563 10.6151
R743 B.n563 B.n38 10.6151
R744 B.n559 B.n38 10.6151
R745 B.n559 B.n558 10.6151
R746 B.n558 B.n557 10.6151
R747 B.n557 B.n40 10.6151
R748 B.n553 B.n552 10.6151
R749 B.n552 B.n551 10.6151
R750 B.n551 B.n45 10.6151
R751 B.n547 B.n45 10.6151
R752 B.n547 B.n546 10.6151
R753 B.n546 B.n545 10.6151
R754 B.n545 B.n47 10.6151
R755 B.n541 B.n47 10.6151
R756 B.n541 B.n540 10.6151
R757 B.n538 B.n51 10.6151
R758 B.n534 B.n51 10.6151
R759 B.n534 B.n533 10.6151
R760 B.n533 B.n532 10.6151
R761 B.n532 B.n53 10.6151
R762 B.n528 B.n53 10.6151
R763 B.n528 B.n527 10.6151
R764 B.n527 B.n526 10.6151
R765 B.n526 B.n55 10.6151
R766 B.n522 B.n55 10.6151
R767 B.n522 B.n521 10.6151
R768 B.n521 B.n520 10.6151
R769 B.n520 B.n57 10.6151
R770 B.n516 B.n57 10.6151
R771 B.n516 B.n515 10.6151
R772 B.n515 B.n514 10.6151
R773 B.n514 B.n59 10.6151
R774 B.n510 B.n59 10.6151
R775 B.n510 B.n509 10.6151
R776 B.n509 B.n508 10.6151
R777 B.n508 B.n61 10.6151
R778 B.n504 B.n61 10.6151
R779 B.n504 B.n503 10.6151
R780 B.n503 B.n502 10.6151
R781 B.n502 B.n63 10.6151
R782 B.n498 B.n63 10.6151
R783 B.n498 B.n497 10.6151
R784 B.n497 B.n496 10.6151
R785 B.n496 B.n65 10.6151
R786 B.n492 B.n65 10.6151
R787 B.n492 B.n491 10.6151
R788 B.n491 B.n490 10.6151
R789 B.n490 B.n67 10.6151
R790 B.n486 B.n67 10.6151
R791 B.n486 B.n485 10.6151
R792 B.n485 B.n484 10.6151
R793 B.n484 B.n69 10.6151
R794 B.n480 B.n69 10.6151
R795 B.n480 B.n479 10.6151
R796 B.n479 B.n478 10.6151
R797 B.n478 B.n71 10.6151
R798 B.n474 B.n71 10.6151
R799 B.n474 B.n473 10.6151
R800 B.n473 B.n472 10.6151
R801 B.n472 B.n73 10.6151
R802 B.n468 B.n73 10.6151
R803 B.n468 B.n467 10.6151
R804 B.n467 B.n466 10.6151
R805 B.n466 B.n75 10.6151
R806 B.n462 B.n75 10.6151
R807 B.n462 B.n461 10.6151
R808 B.n461 B.n460 10.6151
R809 B.n460 B.n77 10.6151
R810 B.n456 B.n77 10.6151
R811 B.n456 B.n455 10.6151
R812 B.n455 B.n454 10.6151
R813 B.n454 B.n79 10.6151
R814 B.n450 B.n79 10.6151
R815 B.n450 B.n449 10.6151
R816 B.n449 B.n448 10.6151
R817 B.n448 B.n81 10.6151
R818 B.n444 B.n81 10.6151
R819 B.n444 B.n443 10.6151
R820 B.n402 B.n95 10.6151
R821 B.n406 B.n95 10.6151
R822 B.n407 B.n406 10.6151
R823 B.n408 B.n407 10.6151
R824 B.n408 B.n93 10.6151
R825 B.n412 B.n93 10.6151
R826 B.n413 B.n412 10.6151
R827 B.n414 B.n413 10.6151
R828 B.n414 B.n91 10.6151
R829 B.n418 B.n91 10.6151
R830 B.n419 B.n418 10.6151
R831 B.n420 B.n419 10.6151
R832 B.n420 B.n89 10.6151
R833 B.n424 B.n89 10.6151
R834 B.n425 B.n424 10.6151
R835 B.n426 B.n425 10.6151
R836 B.n426 B.n87 10.6151
R837 B.n430 B.n87 10.6151
R838 B.n431 B.n430 10.6151
R839 B.n432 B.n431 10.6151
R840 B.n432 B.n85 10.6151
R841 B.n436 B.n85 10.6151
R842 B.n437 B.n436 10.6151
R843 B.n438 B.n437 10.6151
R844 B.n438 B.n83 10.6151
R845 B.n442 B.n83 10.6151
R846 B.n196 B.n169 10.6151
R847 B.n197 B.n196 10.6151
R848 B.n198 B.n197 10.6151
R849 B.n198 B.n167 10.6151
R850 B.n202 B.n167 10.6151
R851 B.n203 B.n202 10.6151
R852 B.n204 B.n203 10.6151
R853 B.n204 B.n165 10.6151
R854 B.n208 B.n165 10.6151
R855 B.n209 B.n208 10.6151
R856 B.n210 B.n209 10.6151
R857 B.n210 B.n163 10.6151
R858 B.n214 B.n163 10.6151
R859 B.n215 B.n214 10.6151
R860 B.n216 B.n215 10.6151
R861 B.n216 B.n161 10.6151
R862 B.n220 B.n161 10.6151
R863 B.n221 B.n220 10.6151
R864 B.n222 B.n221 10.6151
R865 B.n222 B.n159 10.6151
R866 B.n226 B.n159 10.6151
R867 B.n227 B.n226 10.6151
R868 B.n228 B.n227 10.6151
R869 B.n228 B.n157 10.6151
R870 B.n232 B.n157 10.6151
R871 B.n233 B.n232 10.6151
R872 B.n234 B.n233 10.6151
R873 B.n234 B.n155 10.6151
R874 B.n238 B.n155 10.6151
R875 B.n239 B.n238 10.6151
R876 B.n240 B.n239 10.6151
R877 B.n240 B.n153 10.6151
R878 B.n244 B.n153 10.6151
R879 B.n245 B.n244 10.6151
R880 B.n246 B.n245 10.6151
R881 B.n246 B.n151 10.6151
R882 B.n250 B.n151 10.6151
R883 B.n251 B.n250 10.6151
R884 B.n252 B.n251 10.6151
R885 B.n252 B.n149 10.6151
R886 B.n256 B.n149 10.6151
R887 B.n257 B.n256 10.6151
R888 B.n258 B.n257 10.6151
R889 B.n258 B.n147 10.6151
R890 B.n262 B.n147 10.6151
R891 B.n263 B.n262 10.6151
R892 B.n264 B.n263 10.6151
R893 B.n264 B.n145 10.6151
R894 B.n268 B.n145 10.6151
R895 B.n269 B.n268 10.6151
R896 B.n270 B.n269 10.6151
R897 B.n270 B.n143 10.6151
R898 B.n274 B.n143 10.6151
R899 B.n275 B.n274 10.6151
R900 B.n276 B.n275 10.6151
R901 B.n276 B.n141 10.6151
R902 B.n280 B.n141 10.6151
R903 B.n281 B.n280 10.6151
R904 B.n282 B.n281 10.6151
R905 B.n282 B.n139 10.6151
R906 B.n286 B.n139 10.6151
R907 B.n287 B.n286 10.6151
R908 B.n288 B.n287 10.6151
R909 B.n292 B.n291 10.6151
R910 B.n293 B.n292 10.6151
R911 B.n293 B.n133 10.6151
R912 B.n297 B.n133 10.6151
R913 B.n298 B.n297 10.6151
R914 B.n299 B.n298 10.6151
R915 B.n299 B.n131 10.6151
R916 B.n303 B.n131 10.6151
R917 B.n304 B.n303 10.6151
R918 B.n306 B.n127 10.6151
R919 B.n310 B.n127 10.6151
R920 B.n311 B.n310 10.6151
R921 B.n312 B.n311 10.6151
R922 B.n312 B.n125 10.6151
R923 B.n316 B.n125 10.6151
R924 B.n317 B.n316 10.6151
R925 B.n318 B.n317 10.6151
R926 B.n318 B.n123 10.6151
R927 B.n322 B.n123 10.6151
R928 B.n323 B.n322 10.6151
R929 B.n324 B.n323 10.6151
R930 B.n324 B.n121 10.6151
R931 B.n328 B.n121 10.6151
R932 B.n329 B.n328 10.6151
R933 B.n330 B.n329 10.6151
R934 B.n330 B.n119 10.6151
R935 B.n334 B.n119 10.6151
R936 B.n335 B.n334 10.6151
R937 B.n336 B.n335 10.6151
R938 B.n336 B.n117 10.6151
R939 B.n340 B.n117 10.6151
R940 B.n341 B.n340 10.6151
R941 B.n342 B.n341 10.6151
R942 B.n342 B.n115 10.6151
R943 B.n346 B.n115 10.6151
R944 B.n347 B.n346 10.6151
R945 B.n348 B.n347 10.6151
R946 B.n348 B.n113 10.6151
R947 B.n352 B.n113 10.6151
R948 B.n353 B.n352 10.6151
R949 B.n354 B.n353 10.6151
R950 B.n354 B.n111 10.6151
R951 B.n358 B.n111 10.6151
R952 B.n359 B.n358 10.6151
R953 B.n360 B.n359 10.6151
R954 B.n360 B.n109 10.6151
R955 B.n364 B.n109 10.6151
R956 B.n365 B.n364 10.6151
R957 B.n366 B.n365 10.6151
R958 B.n366 B.n107 10.6151
R959 B.n370 B.n107 10.6151
R960 B.n371 B.n370 10.6151
R961 B.n372 B.n371 10.6151
R962 B.n372 B.n105 10.6151
R963 B.n376 B.n105 10.6151
R964 B.n377 B.n376 10.6151
R965 B.n378 B.n377 10.6151
R966 B.n378 B.n103 10.6151
R967 B.n382 B.n103 10.6151
R968 B.n383 B.n382 10.6151
R969 B.n384 B.n383 10.6151
R970 B.n384 B.n101 10.6151
R971 B.n388 B.n101 10.6151
R972 B.n389 B.n388 10.6151
R973 B.n390 B.n389 10.6151
R974 B.n390 B.n99 10.6151
R975 B.n394 B.n99 10.6151
R976 B.n395 B.n394 10.6151
R977 B.n396 B.n395 10.6151
R978 B.n396 B.n97 10.6151
R979 B.n400 B.n97 10.6151
R980 B.n401 B.n400 10.6151
R981 B.n192 B.n191 10.6151
R982 B.n191 B.n190 10.6151
R983 B.n190 B.n171 10.6151
R984 B.n186 B.n171 10.6151
R985 B.n186 B.n185 10.6151
R986 B.n185 B.n184 10.6151
R987 B.n184 B.n173 10.6151
R988 B.n180 B.n173 10.6151
R989 B.n180 B.n179 10.6151
R990 B.n179 B.n178 10.6151
R991 B.n178 B.n175 10.6151
R992 B.n175 B.n0 10.6151
R993 B.n667 B.n1 10.6151
R994 B.n667 B.n666 10.6151
R995 B.n666 B.n665 10.6151
R996 B.n665 B.n4 10.6151
R997 B.n661 B.n4 10.6151
R998 B.n661 B.n660 10.6151
R999 B.n660 B.n659 10.6151
R1000 B.n659 B.n6 10.6151
R1001 B.n655 B.n6 10.6151
R1002 B.n655 B.n654 10.6151
R1003 B.n654 B.n653 10.6151
R1004 B.n653 B.n8 10.6151
R1005 B.n44 B.n40 8.74196
R1006 B.n539 B.n538 8.74196
R1007 B.n288 B.n137 8.74196
R1008 B.n306 B.n305 8.74196
R1009 B.n671 B.n0 2.81026
R1010 B.n671 B.n1 2.81026
R1011 B.n553 B.n44 1.87367
R1012 B.n540 B.n539 1.87367
R1013 B.n291 B.n137 1.87367
R1014 B.n305 B.n304 1.87367
R1015 VP.n0 VP.t0 1235.32
R1016 VP.n0 VP.t1 1190.37
R1017 VP VP.n0 0.0516364
R1018 VTAIL.n434 VTAIL.n330 756.745
R1019 VTAIL.n104 VTAIL.n0 756.745
R1020 VTAIL.n324 VTAIL.n220 756.745
R1021 VTAIL.n214 VTAIL.n110 756.745
R1022 VTAIL.n367 VTAIL.n366 585
R1023 VTAIL.n369 VTAIL.n368 585
R1024 VTAIL.n362 VTAIL.n361 585
R1025 VTAIL.n375 VTAIL.n374 585
R1026 VTAIL.n377 VTAIL.n376 585
R1027 VTAIL.n358 VTAIL.n357 585
R1028 VTAIL.n383 VTAIL.n382 585
R1029 VTAIL.n385 VTAIL.n384 585
R1030 VTAIL.n354 VTAIL.n353 585
R1031 VTAIL.n391 VTAIL.n390 585
R1032 VTAIL.n393 VTAIL.n392 585
R1033 VTAIL.n350 VTAIL.n349 585
R1034 VTAIL.n399 VTAIL.n398 585
R1035 VTAIL.n401 VTAIL.n400 585
R1036 VTAIL.n346 VTAIL.n345 585
R1037 VTAIL.n408 VTAIL.n407 585
R1038 VTAIL.n409 VTAIL.n344 585
R1039 VTAIL.n411 VTAIL.n410 585
R1040 VTAIL.n342 VTAIL.n341 585
R1041 VTAIL.n417 VTAIL.n416 585
R1042 VTAIL.n419 VTAIL.n418 585
R1043 VTAIL.n338 VTAIL.n337 585
R1044 VTAIL.n425 VTAIL.n424 585
R1045 VTAIL.n427 VTAIL.n426 585
R1046 VTAIL.n334 VTAIL.n333 585
R1047 VTAIL.n433 VTAIL.n432 585
R1048 VTAIL.n435 VTAIL.n434 585
R1049 VTAIL.n37 VTAIL.n36 585
R1050 VTAIL.n39 VTAIL.n38 585
R1051 VTAIL.n32 VTAIL.n31 585
R1052 VTAIL.n45 VTAIL.n44 585
R1053 VTAIL.n47 VTAIL.n46 585
R1054 VTAIL.n28 VTAIL.n27 585
R1055 VTAIL.n53 VTAIL.n52 585
R1056 VTAIL.n55 VTAIL.n54 585
R1057 VTAIL.n24 VTAIL.n23 585
R1058 VTAIL.n61 VTAIL.n60 585
R1059 VTAIL.n63 VTAIL.n62 585
R1060 VTAIL.n20 VTAIL.n19 585
R1061 VTAIL.n69 VTAIL.n68 585
R1062 VTAIL.n71 VTAIL.n70 585
R1063 VTAIL.n16 VTAIL.n15 585
R1064 VTAIL.n78 VTAIL.n77 585
R1065 VTAIL.n79 VTAIL.n14 585
R1066 VTAIL.n81 VTAIL.n80 585
R1067 VTAIL.n12 VTAIL.n11 585
R1068 VTAIL.n87 VTAIL.n86 585
R1069 VTAIL.n89 VTAIL.n88 585
R1070 VTAIL.n8 VTAIL.n7 585
R1071 VTAIL.n95 VTAIL.n94 585
R1072 VTAIL.n97 VTAIL.n96 585
R1073 VTAIL.n4 VTAIL.n3 585
R1074 VTAIL.n103 VTAIL.n102 585
R1075 VTAIL.n105 VTAIL.n104 585
R1076 VTAIL.n325 VTAIL.n324 585
R1077 VTAIL.n323 VTAIL.n322 585
R1078 VTAIL.n224 VTAIL.n223 585
R1079 VTAIL.n317 VTAIL.n316 585
R1080 VTAIL.n315 VTAIL.n314 585
R1081 VTAIL.n228 VTAIL.n227 585
R1082 VTAIL.n309 VTAIL.n308 585
R1083 VTAIL.n307 VTAIL.n306 585
R1084 VTAIL.n232 VTAIL.n231 585
R1085 VTAIL.n236 VTAIL.n234 585
R1086 VTAIL.n301 VTAIL.n300 585
R1087 VTAIL.n299 VTAIL.n298 585
R1088 VTAIL.n238 VTAIL.n237 585
R1089 VTAIL.n293 VTAIL.n292 585
R1090 VTAIL.n291 VTAIL.n290 585
R1091 VTAIL.n242 VTAIL.n241 585
R1092 VTAIL.n285 VTAIL.n284 585
R1093 VTAIL.n283 VTAIL.n282 585
R1094 VTAIL.n246 VTAIL.n245 585
R1095 VTAIL.n277 VTAIL.n276 585
R1096 VTAIL.n275 VTAIL.n274 585
R1097 VTAIL.n250 VTAIL.n249 585
R1098 VTAIL.n269 VTAIL.n268 585
R1099 VTAIL.n267 VTAIL.n266 585
R1100 VTAIL.n254 VTAIL.n253 585
R1101 VTAIL.n261 VTAIL.n260 585
R1102 VTAIL.n259 VTAIL.n258 585
R1103 VTAIL.n215 VTAIL.n214 585
R1104 VTAIL.n213 VTAIL.n212 585
R1105 VTAIL.n114 VTAIL.n113 585
R1106 VTAIL.n207 VTAIL.n206 585
R1107 VTAIL.n205 VTAIL.n204 585
R1108 VTAIL.n118 VTAIL.n117 585
R1109 VTAIL.n199 VTAIL.n198 585
R1110 VTAIL.n197 VTAIL.n196 585
R1111 VTAIL.n122 VTAIL.n121 585
R1112 VTAIL.n126 VTAIL.n124 585
R1113 VTAIL.n191 VTAIL.n190 585
R1114 VTAIL.n189 VTAIL.n188 585
R1115 VTAIL.n128 VTAIL.n127 585
R1116 VTAIL.n183 VTAIL.n182 585
R1117 VTAIL.n181 VTAIL.n180 585
R1118 VTAIL.n132 VTAIL.n131 585
R1119 VTAIL.n175 VTAIL.n174 585
R1120 VTAIL.n173 VTAIL.n172 585
R1121 VTAIL.n136 VTAIL.n135 585
R1122 VTAIL.n167 VTAIL.n166 585
R1123 VTAIL.n165 VTAIL.n164 585
R1124 VTAIL.n140 VTAIL.n139 585
R1125 VTAIL.n159 VTAIL.n158 585
R1126 VTAIL.n157 VTAIL.n156 585
R1127 VTAIL.n144 VTAIL.n143 585
R1128 VTAIL.n151 VTAIL.n150 585
R1129 VTAIL.n149 VTAIL.n148 585
R1130 VTAIL.n365 VTAIL.t1 327.466
R1131 VTAIL.n35 VTAIL.t3 327.466
R1132 VTAIL.n257 VTAIL.t2 327.466
R1133 VTAIL.n147 VTAIL.t0 327.466
R1134 VTAIL.n368 VTAIL.n367 171.744
R1135 VTAIL.n368 VTAIL.n361 171.744
R1136 VTAIL.n375 VTAIL.n361 171.744
R1137 VTAIL.n376 VTAIL.n375 171.744
R1138 VTAIL.n376 VTAIL.n357 171.744
R1139 VTAIL.n383 VTAIL.n357 171.744
R1140 VTAIL.n384 VTAIL.n383 171.744
R1141 VTAIL.n384 VTAIL.n353 171.744
R1142 VTAIL.n391 VTAIL.n353 171.744
R1143 VTAIL.n392 VTAIL.n391 171.744
R1144 VTAIL.n392 VTAIL.n349 171.744
R1145 VTAIL.n399 VTAIL.n349 171.744
R1146 VTAIL.n400 VTAIL.n399 171.744
R1147 VTAIL.n400 VTAIL.n345 171.744
R1148 VTAIL.n408 VTAIL.n345 171.744
R1149 VTAIL.n409 VTAIL.n408 171.744
R1150 VTAIL.n410 VTAIL.n409 171.744
R1151 VTAIL.n410 VTAIL.n341 171.744
R1152 VTAIL.n417 VTAIL.n341 171.744
R1153 VTAIL.n418 VTAIL.n417 171.744
R1154 VTAIL.n418 VTAIL.n337 171.744
R1155 VTAIL.n425 VTAIL.n337 171.744
R1156 VTAIL.n426 VTAIL.n425 171.744
R1157 VTAIL.n426 VTAIL.n333 171.744
R1158 VTAIL.n433 VTAIL.n333 171.744
R1159 VTAIL.n434 VTAIL.n433 171.744
R1160 VTAIL.n38 VTAIL.n37 171.744
R1161 VTAIL.n38 VTAIL.n31 171.744
R1162 VTAIL.n45 VTAIL.n31 171.744
R1163 VTAIL.n46 VTAIL.n45 171.744
R1164 VTAIL.n46 VTAIL.n27 171.744
R1165 VTAIL.n53 VTAIL.n27 171.744
R1166 VTAIL.n54 VTAIL.n53 171.744
R1167 VTAIL.n54 VTAIL.n23 171.744
R1168 VTAIL.n61 VTAIL.n23 171.744
R1169 VTAIL.n62 VTAIL.n61 171.744
R1170 VTAIL.n62 VTAIL.n19 171.744
R1171 VTAIL.n69 VTAIL.n19 171.744
R1172 VTAIL.n70 VTAIL.n69 171.744
R1173 VTAIL.n70 VTAIL.n15 171.744
R1174 VTAIL.n78 VTAIL.n15 171.744
R1175 VTAIL.n79 VTAIL.n78 171.744
R1176 VTAIL.n80 VTAIL.n79 171.744
R1177 VTAIL.n80 VTAIL.n11 171.744
R1178 VTAIL.n87 VTAIL.n11 171.744
R1179 VTAIL.n88 VTAIL.n87 171.744
R1180 VTAIL.n88 VTAIL.n7 171.744
R1181 VTAIL.n95 VTAIL.n7 171.744
R1182 VTAIL.n96 VTAIL.n95 171.744
R1183 VTAIL.n96 VTAIL.n3 171.744
R1184 VTAIL.n103 VTAIL.n3 171.744
R1185 VTAIL.n104 VTAIL.n103 171.744
R1186 VTAIL.n324 VTAIL.n323 171.744
R1187 VTAIL.n323 VTAIL.n223 171.744
R1188 VTAIL.n316 VTAIL.n223 171.744
R1189 VTAIL.n316 VTAIL.n315 171.744
R1190 VTAIL.n315 VTAIL.n227 171.744
R1191 VTAIL.n308 VTAIL.n227 171.744
R1192 VTAIL.n308 VTAIL.n307 171.744
R1193 VTAIL.n307 VTAIL.n231 171.744
R1194 VTAIL.n236 VTAIL.n231 171.744
R1195 VTAIL.n300 VTAIL.n236 171.744
R1196 VTAIL.n300 VTAIL.n299 171.744
R1197 VTAIL.n299 VTAIL.n237 171.744
R1198 VTAIL.n292 VTAIL.n237 171.744
R1199 VTAIL.n292 VTAIL.n291 171.744
R1200 VTAIL.n291 VTAIL.n241 171.744
R1201 VTAIL.n284 VTAIL.n241 171.744
R1202 VTAIL.n284 VTAIL.n283 171.744
R1203 VTAIL.n283 VTAIL.n245 171.744
R1204 VTAIL.n276 VTAIL.n245 171.744
R1205 VTAIL.n276 VTAIL.n275 171.744
R1206 VTAIL.n275 VTAIL.n249 171.744
R1207 VTAIL.n268 VTAIL.n249 171.744
R1208 VTAIL.n268 VTAIL.n267 171.744
R1209 VTAIL.n267 VTAIL.n253 171.744
R1210 VTAIL.n260 VTAIL.n253 171.744
R1211 VTAIL.n260 VTAIL.n259 171.744
R1212 VTAIL.n214 VTAIL.n213 171.744
R1213 VTAIL.n213 VTAIL.n113 171.744
R1214 VTAIL.n206 VTAIL.n113 171.744
R1215 VTAIL.n206 VTAIL.n205 171.744
R1216 VTAIL.n205 VTAIL.n117 171.744
R1217 VTAIL.n198 VTAIL.n117 171.744
R1218 VTAIL.n198 VTAIL.n197 171.744
R1219 VTAIL.n197 VTAIL.n121 171.744
R1220 VTAIL.n126 VTAIL.n121 171.744
R1221 VTAIL.n190 VTAIL.n126 171.744
R1222 VTAIL.n190 VTAIL.n189 171.744
R1223 VTAIL.n189 VTAIL.n127 171.744
R1224 VTAIL.n182 VTAIL.n127 171.744
R1225 VTAIL.n182 VTAIL.n181 171.744
R1226 VTAIL.n181 VTAIL.n131 171.744
R1227 VTAIL.n174 VTAIL.n131 171.744
R1228 VTAIL.n174 VTAIL.n173 171.744
R1229 VTAIL.n173 VTAIL.n135 171.744
R1230 VTAIL.n166 VTAIL.n135 171.744
R1231 VTAIL.n166 VTAIL.n165 171.744
R1232 VTAIL.n165 VTAIL.n139 171.744
R1233 VTAIL.n158 VTAIL.n139 171.744
R1234 VTAIL.n158 VTAIL.n157 171.744
R1235 VTAIL.n157 VTAIL.n143 171.744
R1236 VTAIL.n150 VTAIL.n143 171.744
R1237 VTAIL.n150 VTAIL.n149 171.744
R1238 VTAIL.n367 VTAIL.t1 85.8723
R1239 VTAIL.n37 VTAIL.t3 85.8723
R1240 VTAIL.n259 VTAIL.t2 85.8723
R1241 VTAIL.n149 VTAIL.t0 85.8723
R1242 VTAIL.n439 VTAIL.n438 32.9611
R1243 VTAIL.n109 VTAIL.n108 32.9611
R1244 VTAIL.n329 VTAIL.n328 32.9611
R1245 VTAIL.n219 VTAIL.n218 32.9611
R1246 VTAIL.n219 VTAIL.n109 30.8152
R1247 VTAIL.n439 VTAIL.n329 30.0996
R1248 VTAIL.n366 VTAIL.n365 16.3895
R1249 VTAIL.n36 VTAIL.n35 16.3895
R1250 VTAIL.n258 VTAIL.n257 16.3895
R1251 VTAIL.n148 VTAIL.n147 16.3895
R1252 VTAIL.n411 VTAIL.n342 13.1884
R1253 VTAIL.n81 VTAIL.n12 13.1884
R1254 VTAIL.n234 VTAIL.n232 13.1884
R1255 VTAIL.n124 VTAIL.n122 13.1884
R1256 VTAIL.n369 VTAIL.n364 12.8005
R1257 VTAIL.n412 VTAIL.n344 12.8005
R1258 VTAIL.n416 VTAIL.n415 12.8005
R1259 VTAIL.n39 VTAIL.n34 12.8005
R1260 VTAIL.n82 VTAIL.n14 12.8005
R1261 VTAIL.n86 VTAIL.n85 12.8005
R1262 VTAIL.n306 VTAIL.n305 12.8005
R1263 VTAIL.n302 VTAIL.n301 12.8005
R1264 VTAIL.n261 VTAIL.n256 12.8005
R1265 VTAIL.n196 VTAIL.n195 12.8005
R1266 VTAIL.n192 VTAIL.n191 12.8005
R1267 VTAIL.n151 VTAIL.n146 12.8005
R1268 VTAIL.n370 VTAIL.n362 12.0247
R1269 VTAIL.n407 VTAIL.n406 12.0247
R1270 VTAIL.n419 VTAIL.n340 12.0247
R1271 VTAIL.n40 VTAIL.n32 12.0247
R1272 VTAIL.n77 VTAIL.n76 12.0247
R1273 VTAIL.n89 VTAIL.n10 12.0247
R1274 VTAIL.n309 VTAIL.n230 12.0247
R1275 VTAIL.n298 VTAIL.n235 12.0247
R1276 VTAIL.n262 VTAIL.n254 12.0247
R1277 VTAIL.n199 VTAIL.n120 12.0247
R1278 VTAIL.n188 VTAIL.n125 12.0247
R1279 VTAIL.n152 VTAIL.n144 12.0247
R1280 VTAIL.n374 VTAIL.n373 11.249
R1281 VTAIL.n405 VTAIL.n346 11.249
R1282 VTAIL.n420 VTAIL.n338 11.249
R1283 VTAIL.n44 VTAIL.n43 11.249
R1284 VTAIL.n75 VTAIL.n16 11.249
R1285 VTAIL.n90 VTAIL.n8 11.249
R1286 VTAIL.n310 VTAIL.n228 11.249
R1287 VTAIL.n297 VTAIL.n238 11.249
R1288 VTAIL.n266 VTAIL.n265 11.249
R1289 VTAIL.n200 VTAIL.n118 11.249
R1290 VTAIL.n187 VTAIL.n128 11.249
R1291 VTAIL.n156 VTAIL.n155 11.249
R1292 VTAIL.n377 VTAIL.n360 10.4732
R1293 VTAIL.n402 VTAIL.n401 10.4732
R1294 VTAIL.n424 VTAIL.n423 10.4732
R1295 VTAIL.n47 VTAIL.n30 10.4732
R1296 VTAIL.n72 VTAIL.n71 10.4732
R1297 VTAIL.n94 VTAIL.n93 10.4732
R1298 VTAIL.n314 VTAIL.n313 10.4732
R1299 VTAIL.n294 VTAIL.n293 10.4732
R1300 VTAIL.n269 VTAIL.n252 10.4732
R1301 VTAIL.n204 VTAIL.n203 10.4732
R1302 VTAIL.n184 VTAIL.n183 10.4732
R1303 VTAIL.n159 VTAIL.n142 10.4732
R1304 VTAIL.n378 VTAIL.n358 9.69747
R1305 VTAIL.n398 VTAIL.n348 9.69747
R1306 VTAIL.n427 VTAIL.n336 9.69747
R1307 VTAIL.n48 VTAIL.n28 9.69747
R1308 VTAIL.n68 VTAIL.n18 9.69747
R1309 VTAIL.n97 VTAIL.n6 9.69747
R1310 VTAIL.n317 VTAIL.n226 9.69747
R1311 VTAIL.n290 VTAIL.n240 9.69747
R1312 VTAIL.n270 VTAIL.n250 9.69747
R1313 VTAIL.n207 VTAIL.n116 9.69747
R1314 VTAIL.n180 VTAIL.n130 9.69747
R1315 VTAIL.n160 VTAIL.n140 9.69747
R1316 VTAIL.n438 VTAIL.n437 9.45567
R1317 VTAIL.n108 VTAIL.n107 9.45567
R1318 VTAIL.n328 VTAIL.n327 9.45567
R1319 VTAIL.n218 VTAIL.n217 9.45567
R1320 VTAIL.n437 VTAIL.n436 9.3005
R1321 VTAIL.n431 VTAIL.n430 9.3005
R1322 VTAIL.n429 VTAIL.n428 9.3005
R1323 VTAIL.n336 VTAIL.n335 9.3005
R1324 VTAIL.n423 VTAIL.n422 9.3005
R1325 VTAIL.n421 VTAIL.n420 9.3005
R1326 VTAIL.n340 VTAIL.n339 9.3005
R1327 VTAIL.n415 VTAIL.n414 9.3005
R1328 VTAIL.n387 VTAIL.n386 9.3005
R1329 VTAIL.n356 VTAIL.n355 9.3005
R1330 VTAIL.n381 VTAIL.n380 9.3005
R1331 VTAIL.n379 VTAIL.n378 9.3005
R1332 VTAIL.n360 VTAIL.n359 9.3005
R1333 VTAIL.n373 VTAIL.n372 9.3005
R1334 VTAIL.n371 VTAIL.n370 9.3005
R1335 VTAIL.n364 VTAIL.n363 9.3005
R1336 VTAIL.n389 VTAIL.n388 9.3005
R1337 VTAIL.n352 VTAIL.n351 9.3005
R1338 VTAIL.n395 VTAIL.n394 9.3005
R1339 VTAIL.n397 VTAIL.n396 9.3005
R1340 VTAIL.n348 VTAIL.n347 9.3005
R1341 VTAIL.n403 VTAIL.n402 9.3005
R1342 VTAIL.n405 VTAIL.n404 9.3005
R1343 VTAIL.n406 VTAIL.n343 9.3005
R1344 VTAIL.n413 VTAIL.n412 9.3005
R1345 VTAIL.n332 VTAIL.n331 9.3005
R1346 VTAIL.n107 VTAIL.n106 9.3005
R1347 VTAIL.n101 VTAIL.n100 9.3005
R1348 VTAIL.n99 VTAIL.n98 9.3005
R1349 VTAIL.n6 VTAIL.n5 9.3005
R1350 VTAIL.n93 VTAIL.n92 9.3005
R1351 VTAIL.n91 VTAIL.n90 9.3005
R1352 VTAIL.n10 VTAIL.n9 9.3005
R1353 VTAIL.n85 VTAIL.n84 9.3005
R1354 VTAIL.n57 VTAIL.n56 9.3005
R1355 VTAIL.n26 VTAIL.n25 9.3005
R1356 VTAIL.n51 VTAIL.n50 9.3005
R1357 VTAIL.n49 VTAIL.n48 9.3005
R1358 VTAIL.n30 VTAIL.n29 9.3005
R1359 VTAIL.n43 VTAIL.n42 9.3005
R1360 VTAIL.n41 VTAIL.n40 9.3005
R1361 VTAIL.n34 VTAIL.n33 9.3005
R1362 VTAIL.n59 VTAIL.n58 9.3005
R1363 VTAIL.n22 VTAIL.n21 9.3005
R1364 VTAIL.n65 VTAIL.n64 9.3005
R1365 VTAIL.n67 VTAIL.n66 9.3005
R1366 VTAIL.n18 VTAIL.n17 9.3005
R1367 VTAIL.n73 VTAIL.n72 9.3005
R1368 VTAIL.n75 VTAIL.n74 9.3005
R1369 VTAIL.n76 VTAIL.n13 9.3005
R1370 VTAIL.n83 VTAIL.n82 9.3005
R1371 VTAIL.n2 VTAIL.n1 9.3005
R1372 VTAIL.n244 VTAIL.n243 9.3005
R1373 VTAIL.n287 VTAIL.n286 9.3005
R1374 VTAIL.n289 VTAIL.n288 9.3005
R1375 VTAIL.n240 VTAIL.n239 9.3005
R1376 VTAIL.n295 VTAIL.n294 9.3005
R1377 VTAIL.n297 VTAIL.n296 9.3005
R1378 VTAIL.n235 VTAIL.n233 9.3005
R1379 VTAIL.n303 VTAIL.n302 9.3005
R1380 VTAIL.n327 VTAIL.n326 9.3005
R1381 VTAIL.n222 VTAIL.n221 9.3005
R1382 VTAIL.n321 VTAIL.n320 9.3005
R1383 VTAIL.n319 VTAIL.n318 9.3005
R1384 VTAIL.n226 VTAIL.n225 9.3005
R1385 VTAIL.n313 VTAIL.n312 9.3005
R1386 VTAIL.n311 VTAIL.n310 9.3005
R1387 VTAIL.n230 VTAIL.n229 9.3005
R1388 VTAIL.n305 VTAIL.n304 9.3005
R1389 VTAIL.n281 VTAIL.n280 9.3005
R1390 VTAIL.n279 VTAIL.n278 9.3005
R1391 VTAIL.n248 VTAIL.n247 9.3005
R1392 VTAIL.n273 VTAIL.n272 9.3005
R1393 VTAIL.n271 VTAIL.n270 9.3005
R1394 VTAIL.n252 VTAIL.n251 9.3005
R1395 VTAIL.n265 VTAIL.n264 9.3005
R1396 VTAIL.n263 VTAIL.n262 9.3005
R1397 VTAIL.n256 VTAIL.n255 9.3005
R1398 VTAIL.n134 VTAIL.n133 9.3005
R1399 VTAIL.n177 VTAIL.n176 9.3005
R1400 VTAIL.n179 VTAIL.n178 9.3005
R1401 VTAIL.n130 VTAIL.n129 9.3005
R1402 VTAIL.n185 VTAIL.n184 9.3005
R1403 VTAIL.n187 VTAIL.n186 9.3005
R1404 VTAIL.n125 VTAIL.n123 9.3005
R1405 VTAIL.n193 VTAIL.n192 9.3005
R1406 VTAIL.n217 VTAIL.n216 9.3005
R1407 VTAIL.n112 VTAIL.n111 9.3005
R1408 VTAIL.n211 VTAIL.n210 9.3005
R1409 VTAIL.n209 VTAIL.n208 9.3005
R1410 VTAIL.n116 VTAIL.n115 9.3005
R1411 VTAIL.n203 VTAIL.n202 9.3005
R1412 VTAIL.n201 VTAIL.n200 9.3005
R1413 VTAIL.n120 VTAIL.n119 9.3005
R1414 VTAIL.n195 VTAIL.n194 9.3005
R1415 VTAIL.n171 VTAIL.n170 9.3005
R1416 VTAIL.n169 VTAIL.n168 9.3005
R1417 VTAIL.n138 VTAIL.n137 9.3005
R1418 VTAIL.n163 VTAIL.n162 9.3005
R1419 VTAIL.n161 VTAIL.n160 9.3005
R1420 VTAIL.n142 VTAIL.n141 9.3005
R1421 VTAIL.n155 VTAIL.n154 9.3005
R1422 VTAIL.n153 VTAIL.n152 9.3005
R1423 VTAIL.n146 VTAIL.n145 9.3005
R1424 VTAIL.n382 VTAIL.n381 8.92171
R1425 VTAIL.n397 VTAIL.n350 8.92171
R1426 VTAIL.n428 VTAIL.n334 8.92171
R1427 VTAIL.n52 VTAIL.n51 8.92171
R1428 VTAIL.n67 VTAIL.n20 8.92171
R1429 VTAIL.n98 VTAIL.n4 8.92171
R1430 VTAIL.n318 VTAIL.n224 8.92171
R1431 VTAIL.n289 VTAIL.n242 8.92171
R1432 VTAIL.n274 VTAIL.n273 8.92171
R1433 VTAIL.n208 VTAIL.n114 8.92171
R1434 VTAIL.n179 VTAIL.n132 8.92171
R1435 VTAIL.n164 VTAIL.n163 8.92171
R1436 VTAIL.n385 VTAIL.n356 8.14595
R1437 VTAIL.n394 VTAIL.n393 8.14595
R1438 VTAIL.n432 VTAIL.n431 8.14595
R1439 VTAIL.n55 VTAIL.n26 8.14595
R1440 VTAIL.n64 VTAIL.n63 8.14595
R1441 VTAIL.n102 VTAIL.n101 8.14595
R1442 VTAIL.n322 VTAIL.n321 8.14595
R1443 VTAIL.n286 VTAIL.n285 8.14595
R1444 VTAIL.n277 VTAIL.n248 8.14595
R1445 VTAIL.n212 VTAIL.n211 8.14595
R1446 VTAIL.n176 VTAIL.n175 8.14595
R1447 VTAIL.n167 VTAIL.n138 8.14595
R1448 VTAIL.n386 VTAIL.n354 7.3702
R1449 VTAIL.n390 VTAIL.n352 7.3702
R1450 VTAIL.n435 VTAIL.n332 7.3702
R1451 VTAIL.n438 VTAIL.n330 7.3702
R1452 VTAIL.n56 VTAIL.n24 7.3702
R1453 VTAIL.n60 VTAIL.n22 7.3702
R1454 VTAIL.n105 VTAIL.n2 7.3702
R1455 VTAIL.n108 VTAIL.n0 7.3702
R1456 VTAIL.n328 VTAIL.n220 7.3702
R1457 VTAIL.n325 VTAIL.n222 7.3702
R1458 VTAIL.n282 VTAIL.n244 7.3702
R1459 VTAIL.n278 VTAIL.n246 7.3702
R1460 VTAIL.n218 VTAIL.n110 7.3702
R1461 VTAIL.n215 VTAIL.n112 7.3702
R1462 VTAIL.n172 VTAIL.n134 7.3702
R1463 VTAIL.n168 VTAIL.n136 7.3702
R1464 VTAIL.n389 VTAIL.n354 6.59444
R1465 VTAIL.n390 VTAIL.n389 6.59444
R1466 VTAIL.n436 VTAIL.n435 6.59444
R1467 VTAIL.n436 VTAIL.n330 6.59444
R1468 VTAIL.n59 VTAIL.n24 6.59444
R1469 VTAIL.n60 VTAIL.n59 6.59444
R1470 VTAIL.n106 VTAIL.n105 6.59444
R1471 VTAIL.n106 VTAIL.n0 6.59444
R1472 VTAIL.n326 VTAIL.n220 6.59444
R1473 VTAIL.n326 VTAIL.n325 6.59444
R1474 VTAIL.n282 VTAIL.n281 6.59444
R1475 VTAIL.n281 VTAIL.n246 6.59444
R1476 VTAIL.n216 VTAIL.n110 6.59444
R1477 VTAIL.n216 VTAIL.n215 6.59444
R1478 VTAIL.n172 VTAIL.n171 6.59444
R1479 VTAIL.n171 VTAIL.n136 6.59444
R1480 VTAIL.n386 VTAIL.n385 5.81868
R1481 VTAIL.n393 VTAIL.n352 5.81868
R1482 VTAIL.n432 VTAIL.n332 5.81868
R1483 VTAIL.n56 VTAIL.n55 5.81868
R1484 VTAIL.n63 VTAIL.n22 5.81868
R1485 VTAIL.n102 VTAIL.n2 5.81868
R1486 VTAIL.n322 VTAIL.n222 5.81868
R1487 VTAIL.n285 VTAIL.n244 5.81868
R1488 VTAIL.n278 VTAIL.n277 5.81868
R1489 VTAIL.n212 VTAIL.n112 5.81868
R1490 VTAIL.n175 VTAIL.n134 5.81868
R1491 VTAIL.n168 VTAIL.n167 5.81868
R1492 VTAIL.n382 VTAIL.n356 5.04292
R1493 VTAIL.n394 VTAIL.n350 5.04292
R1494 VTAIL.n431 VTAIL.n334 5.04292
R1495 VTAIL.n52 VTAIL.n26 5.04292
R1496 VTAIL.n64 VTAIL.n20 5.04292
R1497 VTAIL.n101 VTAIL.n4 5.04292
R1498 VTAIL.n321 VTAIL.n224 5.04292
R1499 VTAIL.n286 VTAIL.n242 5.04292
R1500 VTAIL.n274 VTAIL.n248 5.04292
R1501 VTAIL.n211 VTAIL.n114 5.04292
R1502 VTAIL.n176 VTAIL.n132 5.04292
R1503 VTAIL.n164 VTAIL.n138 5.04292
R1504 VTAIL.n381 VTAIL.n358 4.26717
R1505 VTAIL.n398 VTAIL.n397 4.26717
R1506 VTAIL.n428 VTAIL.n427 4.26717
R1507 VTAIL.n51 VTAIL.n28 4.26717
R1508 VTAIL.n68 VTAIL.n67 4.26717
R1509 VTAIL.n98 VTAIL.n97 4.26717
R1510 VTAIL.n318 VTAIL.n317 4.26717
R1511 VTAIL.n290 VTAIL.n289 4.26717
R1512 VTAIL.n273 VTAIL.n250 4.26717
R1513 VTAIL.n208 VTAIL.n207 4.26717
R1514 VTAIL.n180 VTAIL.n179 4.26717
R1515 VTAIL.n163 VTAIL.n140 4.26717
R1516 VTAIL.n365 VTAIL.n363 3.70982
R1517 VTAIL.n35 VTAIL.n33 3.70982
R1518 VTAIL.n257 VTAIL.n255 3.70982
R1519 VTAIL.n147 VTAIL.n145 3.70982
R1520 VTAIL.n378 VTAIL.n377 3.49141
R1521 VTAIL.n401 VTAIL.n348 3.49141
R1522 VTAIL.n424 VTAIL.n336 3.49141
R1523 VTAIL.n48 VTAIL.n47 3.49141
R1524 VTAIL.n71 VTAIL.n18 3.49141
R1525 VTAIL.n94 VTAIL.n6 3.49141
R1526 VTAIL.n314 VTAIL.n226 3.49141
R1527 VTAIL.n293 VTAIL.n240 3.49141
R1528 VTAIL.n270 VTAIL.n269 3.49141
R1529 VTAIL.n204 VTAIL.n116 3.49141
R1530 VTAIL.n183 VTAIL.n130 3.49141
R1531 VTAIL.n160 VTAIL.n159 3.49141
R1532 VTAIL.n374 VTAIL.n360 2.71565
R1533 VTAIL.n402 VTAIL.n346 2.71565
R1534 VTAIL.n423 VTAIL.n338 2.71565
R1535 VTAIL.n44 VTAIL.n30 2.71565
R1536 VTAIL.n72 VTAIL.n16 2.71565
R1537 VTAIL.n93 VTAIL.n8 2.71565
R1538 VTAIL.n313 VTAIL.n228 2.71565
R1539 VTAIL.n294 VTAIL.n238 2.71565
R1540 VTAIL.n266 VTAIL.n252 2.71565
R1541 VTAIL.n203 VTAIL.n118 2.71565
R1542 VTAIL.n184 VTAIL.n128 2.71565
R1543 VTAIL.n156 VTAIL.n142 2.71565
R1544 VTAIL.n373 VTAIL.n362 1.93989
R1545 VTAIL.n407 VTAIL.n405 1.93989
R1546 VTAIL.n420 VTAIL.n419 1.93989
R1547 VTAIL.n43 VTAIL.n32 1.93989
R1548 VTAIL.n77 VTAIL.n75 1.93989
R1549 VTAIL.n90 VTAIL.n89 1.93989
R1550 VTAIL.n310 VTAIL.n309 1.93989
R1551 VTAIL.n298 VTAIL.n297 1.93989
R1552 VTAIL.n265 VTAIL.n254 1.93989
R1553 VTAIL.n200 VTAIL.n199 1.93989
R1554 VTAIL.n188 VTAIL.n187 1.93989
R1555 VTAIL.n155 VTAIL.n144 1.93989
R1556 VTAIL.n370 VTAIL.n369 1.16414
R1557 VTAIL.n406 VTAIL.n344 1.16414
R1558 VTAIL.n416 VTAIL.n340 1.16414
R1559 VTAIL.n40 VTAIL.n39 1.16414
R1560 VTAIL.n76 VTAIL.n14 1.16414
R1561 VTAIL.n86 VTAIL.n10 1.16414
R1562 VTAIL.n306 VTAIL.n230 1.16414
R1563 VTAIL.n301 VTAIL.n235 1.16414
R1564 VTAIL.n262 VTAIL.n261 1.16414
R1565 VTAIL.n196 VTAIL.n120 1.16414
R1566 VTAIL.n191 VTAIL.n125 1.16414
R1567 VTAIL.n152 VTAIL.n151 1.16414
R1568 VTAIL.n329 VTAIL.n219 0.828086
R1569 VTAIL VTAIL.n109 0.707397
R1570 VTAIL.n366 VTAIL.n364 0.388379
R1571 VTAIL.n412 VTAIL.n411 0.388379
R1572 VTAIL.n415 VTAIL.n342 0.388379
R1573 VTAIL.n36 VTAIL.n34 0.388379
R1574 VTAIL.n82 VTAIL.n81 0.388379
R1575 VTAIL.n85 VTAIL.n12 0.388379
R1576 VTAIL.n305 VTAIL.n232 0.388379
R1577 VTAIL.n302 VTAIL.n234 0.388379
R1578 VTAIL.n258 VTAIL.n256 0.388379
R1579 VTAIL.n195 VTAIL.n122 0.388379
R1580 VTAIL.n192 VTAIL.n124 0.388379
R1581 VTAIL.n148 VTAIL.n146 0.388379
R1582 VTAIL.n371 VTAIL.n363 0.155672
R1583 VTAIL.n372 VTAIL.n371 0.155672
R1584 VTAIL.n372 VTAIL.n359 0.155672
R1585 VTAIL.n379 VTAIL.n359 0.155672
R1586 VTAIL.n380 VTAIL.n379 0.155672
R1587 VTAIL.n380 VTAIL.n355 0.155672
R1588 VTAIL.n387 VTAIL.n355 0.155672
R1589 VTAIL.n388 VTAIL.n387 0.155672
R1590 VTAIL.n388 VTAIL.n351 0.155672
R1591 VTAIL.n395 VTAIL.n351 0.155672
R1592 VTAIL.n396 VTAIL.n395 0.155672
R1593 VTAIL.n396 VTAIL.n347 0.155672
R1594 VTAIL.n403 VTAIL.n347 0.155672
R1595 VTAIL.n404 VTAIL.n403 0.155672
R1596 VTAIL.n404 VTAIL.n343 0.155672
R1597 VTAIL.n413 VTAIL.n343 0.155672
R1598 VTAIL.n414 VTAIL.n413 0.155672
R1599 VTAIL.n414 VTAIL.n339 0.155672
R1600 VTAIL.n421 VTAIL.n339 0.155672
R1601 VTAIL.n422 VTAIL.n421 0.155672
R1602 VTAIL.n422 VTAIL.n335 0.155672
R1603 VTAIL.n429 VTAIL.n335 0.155672
R1604 VTAIL.n430 VTAIL.n429 0.155672
R1605 VTAIL.n430 VTAIL.n331 0.155672
R1606 VTAIL.n437 VTAIL.n331 0.155672
R1607 VTAIL.n41 VTAIL.n33 0.155672
R1608 VTAIL.n42 VTAIL.n41 0.155672
R1609 VTAIL.n42 VTAIL.n29 0.155672
R1610 VTAIL.n49 VTAIL.n29 0.155672
R1611 VTAIL.n50 VTAIL.n49 0.155672
R1612 VTAIL.n50 VTAIL.n25 0.155672
R1613 VTAIL.n57 VTAIL.n25 0.155672
R1614 VTAIL.n58 VTAIL.n57 0.155672
R1615 VTAIL.n58 VTAIL.n21 0.155672
R1616 VTAIL.n65 VTAIL.n21 0.155672
R1617 VTAIL.n66 VTAIL.n65 0.155672
R1618 VTAIL.n66 VTAIL.n17 0.155672
R1619 VTAIL.n73 VTAIL.n17 0.155672
R1620 VTAIL.n74 VTAIL.n73 0.155672
R1621 VTAIL.n74 VTAIL.n13 0.155672
R1622 VTAIL.n83 VTAIL.n13 0.155672
R1623 VTAIL.n84 VTAIL.n83 0.155672
R1624 VTAIL.n84 VTAIL.n9 0.155672
R1625 VTAIL.n91 VTAIL.n9 0.155672
R1626 VTAIL.n92 VTAIL.n91 0.155672
R1627 VTAIL.n92 VTAIL.n5 0.155672
R1628 VTAIL.n99 VTAIL.n5 0.155672
R1629 VTAIL.n100 VTAIL.n99 0.155672
R1630 VTAIL.n100 VTAIL.n1 0.155672
R1631 VTAIL.n107 VTAIL.n1 0.155672
R1632 VTAIL.n327 VTAIL.n221 0.155672
R1633 VTAIL.n320 VTAIL.n221 0.155672
R1634 VTAIL.n320 VTAIL.n319 0.155672
R1635 VTAIL.n319 VTAIL.n225 0.155672
R1636 VTAIL.n312 VTAIL.n225 0.155672
R1637 VTAIL.n312 VTAIL.n311 0.155672
R1638 VTAIL.n311 VTAIL.n229 0.155672
R1639 VTAIL.n304 VTAIL.n229 0.155672
R1640 VTAIL.n304 VTAIL.n303 0.155672
R1641 VTAIL.n303 VTAIL.n233 0.155672
R1642 VTAIL.n296 VTAIL.n233 0.155672
R1643 VTAIL.n296 VTAIL.n295 0.155672
R1644 VTAIL.n295 VTAIL.n239 0.155672
R1645 VTAIL.n288 VTAIL.n239 0.155672
R1646 VTAIL.n288 VTAIL.n287 0.155672
R1647 VTAIL.n287 VTAIL.n243 0.155672
R1648 VTAIL.n280 VTAIL.n243 0.155672
R1649 VTAIL.n280 VTAIL.n279 0.155672
R1650 VTAIL.n279 VTAIL.n247 0.155672
R1651 VTAIL.n272 VTAIL.n247 0.155672
R1652 VTAIL.n272 VTAIL.n271 0.155672
R1653 VTAIL.n271 VTAIL.n251 0.155672
R1654 VTAIL.n264 VTAIL.n251 0.155672
R1655 VTAIL.n264 VTAIL.n263 0.155672
R1656 VTAIL.n263 VTAIL.n255 0.155672
R1657 VTAIL.n217 VTAIL.n111 0.155672
R1658 VTAIL.n210 VTAIL.n111 0.155672
R1659 VTAIL.n210 VTAIL.n209 0.155672
R1660 VTAIL.n209 VTAIL.n115 0.155672
R1661 VTAIL.n202 VTAIL.n115 0.155672
R1662 VTAIL.n202 VTAIL.n201 0.155672
R1663 VTAIL.n201 VTAIL.n119 0.155672
R1664 VTAIL.n194 VTAIL.n119 0.155672
R1665 VTAIL.n194 VTAIL.n193 0.155672
R1666 VTAIL.n193 VTAIL.n123 0.155672
R1667 VTAIL.n186 VTAIL.n123 0.155672
R1668 VTAIL.n186 VTAIL.n185 0.155672
R1669 VTAIL.n185 VTAIL.n129 0.155672
R1670 VTAIL.n178 VTAIL.n129 0.155672
R1671 VTAIL.n178 VTAIL.n177 0.155672
R1672 VTAIL.n177 VTAIL.n133 0.155672
R1673 VTAIL.n170 VTAIL.n133 0.155672
R1674 VTAIL.n170 VTAIL.n169 0.155672
R1675 VTAIL.n169 VTAIL.n137 0.155672
R1676 VTAIL.n162 VTAIL.n137 0.155672
R1677 VTAIL.n162 VTAIL.n161 0.155672
R1678 VTAIL.n161 VTAIL.n141 0.155672
R1679 VTAIL.n154 VTAIL.n141 0.155672
R1680 VTAIL.n154 VTAIL.n153 0.155672
R1681 VTAIL.n153 VTAIL.n145 0.155672
R1682 VTAIL VTAIL.n439 0.12119
R1683 VDD1.n104 VDD1.n0 756.745
R1684 VDD1.n213 VDD1.n109 756.745
R1685 VDD1.n105 VDD1.n104 585
R1686 VDD1.n103 VDD1.n102 585
R1687 VDD1.n4 VDD1.n3 585
R1688 VDD1.n97 VDD1.n96 585
R1689 VDD1.n95 VDD1.n94 585
R1690 VDD1.n8 VDD1.n7 585
R1691 VDD1.n89 VDD1.n88 585
R1692 VDD1.n87 VDD1.n86 585
R1693 VDD1.n12 VDD1.n11 585
R1694 VDD1.n16 VDD1.n14 585
R1695 VDD1.n81 VDD1.n80 585
R1696 VDD1.n79 VDD1.n78 585
R1697 VDD1.n18 VDD1.n17 585
R1698 VDD1.n73 VDD1.n72 585
R1699 VDD1.n71 VDD1.n70 585
R1700 VDD1.n22 VDD1.n21 585
R1701 VDD1.n65 VDD1.n64 585
R1702 VDD1.n63 VDD1.n62 585
R1703 VDD1.n26 VDD1.n25 585
R1704 VDD1.n57 VDD1.n56 585
R1705 VDD1.n55 VDD1.n54 585
R1706 VDD1.n30 VDD1.n29 585
R1707 VDD1.n49 VDD1.n48 585
R1708 VDD1.n47 VDD1.n46 585
R1709 VDD1.n34 VDD1.n33 585
R1710 VDD1.n41 VDD1.n40 585
R1711 VDD1.n39 VDD1.n38 585
R1712 VDD1.n146 VDD1.n145 585
R1713 VDD1.n148 VDD1.n147 585
R1714 VDD1.n141 VDD1.n140 585
R1715 VDD1.n154 VDD1.n153 585
R1716 VDD1.n156 VDD1.n155 585
R1717 VDD1.n137 VDD1.n136 585
R1718 VDD1.n162 VDD1.n161 585
R1719 VDD1.n164 VDD1.n163 585
R1720 VDD1.n133 VDD1.n132 585
R1721 VDD1.n170 VDD1.n169 585
R1722 VDD1.n172 VDD1.n171 585
R1723 VDD1.n129 VDD1.n128 585
R1724 VDD1.n178 VDD1.n177 585
R1725 VDD1.n180 VDD1.n179 585
R1726 VDD1.n125 VDD1.n124 585
R1727 VDD1.n187 VDD1.n186 585
R1728 VDD1.n188 VDD1.n123 585
R1729 VDD1.n190 VDD1.n189 585
R1730 VDD1.n121 VDD1.n120 585
R1731 VDD1.n196 VDD1.n195 585
R1732 VDD1.n198 VDD1.n197 585
R1733 VDD1.n117 VDD1.n116 585
R1734 VDD1.n204 VDD1.n203 585
R1735 VDD1.n206 VDD1.n205 585
R1736 VDD1.n113 VDD1.n112 585
R1737 VDD1.n212 VDD1.n211 585
R1738 VDD1.n214 VDD1.n213 585
R1739 VDD1.n37 VDD1.t1 327.466
R1740 VDD1.n144 VDD1.t0 327.466
R1741 VDD1.n104 VDD1.n103 171.744
R1742 VDD1.n103 VDD1.n3 171.744
R1743 VDD1.n96 VDD1.n3 171.744
R1744 VDD1.n96 VDD1.n95 171.744
R1745 VDD1.n95 VDD1.n7 171.744
R1746 VDD1.n88 VDD1.n7 171.744
R1747 VDD1.n88 VDD1.n87 171.744
R1748 VDD1.n87 VDD1.n11 171.744
R1749 VDD1.n16 VDD1.n11 171.744
R1750 VDD1.n80 VDD1.n16 171.744
R1751 VDD1.n80 VDD1.n79 171.744
R1752 VDD1.n79 VDD1.n17 171.744
R1753 VDD1.n72 VDD1.n17 171.744
R1754 VDD1.n72 VDD1.n71 171.744
R1755 VDD1.n71 VDD1.n21 171.744
R1756 VDD1.n64 VDD1.n21 171.744
R1757 VDD1.n64 VDD1.n63 171.744
R1758 VDD1.n63 VDD1.n25 171.744
R1759 VDD1.n56 VDD1.n25 171.744
R1760 VDD1.n56 VDD1.n55 171.744
R1761 VDD1.n55 VDD1.n29 171.744
R1762 VDD1.n48 VDD1.n29 171.744
R1763 VDD1.n48 VDD1.n47 171.744
R1764 VDD1.n47 VDD1.n33 171.744
R1765 VDD1.n40 VDD1.n33 171.744
R1766 VDD1.n40 VDD1.n39 171.744
R1767 VDD1.n147 VDD1.n146 171.744
R1768 VDD1.n147 VDD1.n140 171.744
R1769 VDD1.n154 VDD1.n140 171.744
R1770 VDD1.n155 VDD1.n154 171.744
R1771 VDD1.n155 VDD1.n136 171.744
R1772 VDD1.n162 VDD1.n136 171.744
R1773 VDD1.n163 VDD1.n162 171.744
R1774 VDD1.n163 VDD1.n132 171.744
R1775 VDD1.n170 VDD1.n132 171.744
R1776 VDD1.n171 VDD1.n170 171.744
R1777 VDD1.n171 VDD1.n128 171.744
R1778 VDD1.n178 VDD1.n128 171.744
R1779 VDD1.n179 VDD1.n178 171.744
R1780 VDD1.n179 VDD1.n124 171.744
R1781 VDD1.n187 VDD1.n124 171.744
R1782 VDD1.n188 VDD1.n187 171.744
R1783 VDD1.n189 VDD1.n188 171.744
R1784 VDD1.n189 VDD1.n120 171.744
R1785 VDD1.n196 VDD1.n120 171.744
R1786 VDD1.n197 VDD1.n196 171.744
R1787 VDD1.n197 VDD1.n116 171.744
R1788 VDD1.n204 VDD1.n116 171.744
R1789 VDD1.n205 VDD1.n204 171.744
R1790 VDD1.n205 VDD1.n112 171.744
R1791 VDD1.n212 VDD1.n112 171.744
R1792 VDD1.n213 VDD1.n212 171.744
R1793 VDD1 VDD1.n217 92.4513
R1794 VDD1.n39 VDD1.t1 85.8723
R1795 VDD1.n146 VDD1.t0 85.8723
R1796 VDD1 VDD1.n108 49.877
R1797 VDD1.n38 VDD1.n37 16.3895
R1798 VDD1.n145 VDD1.n144 16.3895
R1799 VDD1.n14 VDD1.n12 13.1884
R1800 VDD1.n190 VDD1.n121 13.1884
R1801 VDD1.n86 VDD1.n85 12.8005
R1802 VDD1.n82 VDD1.n81 12.8005
R1803 VDD1.n41 VDD1.n36 12.8005
R1804 VDD1.n148 VDD1.n143 12.8005
R1805 VDD1.n191 VDD1.n123 12.8005
R1806 VDD1.n195 VDD1.n194 12.8005
R1807 VDD1.n89 VDD1.n10 12.0247
R1808 VDD1.n78 VDD1.n15 12.0247
R1809 VDD1.n42 VDD1.n34 12.0247
R1810 VDD1.n149 VDD1.n141 12.0247
R1811 VDD1.n186 VDD1.n185 12.0247
R1812 VDD1.n198 VDD1.n119 12.0247
R1813 VDD1.n90 VDD1.n8 11.249
R1814 VDD1.n77 VDD1.n18 11.249
R1815 VDD1.n46 VDD1.n45 11.249
R1816 VDD1.n153 VDD1.n152 11.249
R1817 VDD1.n184 VDD1.n125 11.249
R1818 VDD1.n199 VDD1.n117 11.249
R1819 VDD1.n94 VDD1.n93 10.4732
R1820 VDD1.n74 VDD1.n73 10.4732
R1821 VDD1.n49 VDD1.n32 10.4732
R1822 VDD1.n156 VDD1.n139 10.4732
R1823 VDD1.n181 VDD1.n180 10.4732
R1824 VDD1.n203 VDD1.n202 10.4732
R1825 VDD1.n97 VDD1.n6 9.69747
R1826 VDD1.n70 VDD1.n20 9.69747
R1827 VDD1.n50 VDD1.n30 9.69747
R1828 VDD1.n157 VDD1.n137 9.69747
R1829 VDD1.n177 VDD1.n127 9.69747
R1830 VDD1.n206 VDD1.n115 9.69747
R1831 VDD1.n108 VDD1.n107 9.45567
R1832 VDD1.n217 VDD1.n216 9.45567
R1833 VDD1.n24 VDD1.n23 9.3005
R1834 VDD1.n67 VDD1.n66 9.3005
R1835 VDD1.n69 VDD1.n68 9.3005
R1836 VDD1.n20 VDD1.n19 9.3005
R1837 VDD1.n75 VDD1.n74 9.3005
R1838 VDD1.n77 VDD1.n76 9.3005
R1839 VDD1.n15 VDD1.n13 9.3005
R1840 VDD1.n83 VDD1.n82 9.3005
R1841 VDD1.n107 VDD1.n106 9.3005
R1842 VDD1.n2 VDD1.n1 9.3005
R1843 VDD1.n101 VDD1.n100 9.3005
R1844 VDD1.n99 VDD1.n98 9.3005
R1845 VDD1.n6 VDD1.n5 9.3005
R1846 VDD1.n93 VDD1.n92 9.3005
R1847 VDD1.n91 VDD1.n90 9.3005
R1848 VDD1.n10 VDD1.n9 9.3005
R1849 VDD1.n85 VDD1.n84 9.3005
R1850 VDD1.n61 VDD1.n60 9.3005
R1851 VDD1.n59 VDD1.n58 9.3005
R1852 VDD1.n28 VDD1.n27 9.3005
R1853 VDD1.n53 VDD1.n52 9.3005
R1854 VDD1.n51 VDD1.n50 9.3005
R1855 VDD1.n32 VDD1.n31 9.3005
R1856 VDD1.n45 VDD1.n44 9.3005
R1857 VDD1.n43 VDD1.n42 9.3005
R1858 VDD1.n36 VDD1.n35 9.3005
R1859 VDD1.n216 VDD1.n215 9.3005
R1860 VDD1.n210 VDD1.n209 9.3005
R1861 VDD1.n208 VDD1.n207 9.3005
R1862 VDD1.n115 VDD1.n114 9.3005
R1863 VDD1.n202 VDD1.n201 9.3005
R1864 VDD1.n200 VDD1.n199 9.3005
R1865 VDD1.n119 VDD1.n118 9.3005
R1866 VDD1.n194 VDD1.n193 9.3005
R1867 VDD1.n166 VDD1.n165 9.3005
R1868 VDD1.n135 VDD1.n134 9.3005
R1869 VDD1.n160 VDD1.n159 9.3005
R1870 VDD1.n158 VDD1.n157 9.3005
R1871 VDD1.n139 VDD1.n138 9.3005
R1872 VDD1.n152 VDD1.n151 9.3005
R1873 VDD1.n150 VDD1.n149 9.3005
R1874 VDD1.n143 VDD1.n142 9.3005
R1875 VDD1.n168 VDD1.n167 9.3005
R1876 VDD1.n131 VDD1.n130 9.3005
R1877 VDD1.n174 VDD1.n173 9.3005
R1878 VDD1.n176 VDD1.n175 9.3005
R1879 VDD1.n127 VDD1.n126 9.3005
R1880 VDD1.n182 VDD1.n181 9.3005
R1881 VDD1.n184 VDD1.n183 9.3005
R1882 VDD1.n185 VDD1.n122 9.3005
R1883 VDD1.n192 VDD1.n191 9.3005
R1884 VDD1.n111 VDD1.n110 9.3005
R1885 VDD1.n98 VDD1.n4 8.92171
R1886 VDD1.n69 VDD1.n22 8.92171
R1887 VDD1.n54 VDD1.n53 8.92171
R1888 VDD1.n161 VDD1.n160 8.92171
R1889 VDD1.n176 VDD1.n129 8.92171
R1890 VDD1.n207 VDD1.n113 8.92171
R1891 VDD1.n102 VDD1.n101 8.14595
R1892 VDD1.n66 VDD1.n65 8.14595
R1893 VDD1.n57 VDD1.n28 8.14595
R1894 VDD1.n164 VDD1.n135 8.14595
R1895 VDD1.n173 VDD1.n172 8.14595
R1896 VDD1.n211 VDD1.n210 8.14595
R1897 VDD1.n108 VDD1.n0 7.3702
R1898 VDD1.n105 VDD1.n2 7.3702
R1899 VDD1.n62 VDD1.n24 7.3702
R1900 VDD1.n58 VDD1.n26 7.3702
R1901 VDD1.n165 VDD1.n133 7.3702
R1902 VDD1.n169 VDD1.n131 7.3702
R1903 VDD1.n214 VDD1.n111 7.3702
R1904 VDD1.n217 VDD1.n109 7.3702
R1905 VDD1.n106 VDD1.n0 6.59444
R1906 VDD1.n106 VDD1.n105 6.59444
R1907 VDD1.n62 VDD1.n61 6.59444
R1908 VDD1.n61 VDD1.n26 6.59444
R1909 VDD1.n168 VDD1.n133 6.59444
R1910 VDD1.n169 VDD1.n168 6.59444
R1911 VDD1.n215 VDD1.n214 6.59444
R1912 VDD1.n215 VDD1.n109 6.59444
R1913 VDD1.n102 VDD1.n2 5.81868
R1914 VDD1.n65 VDD1.n24 5.81868
R1915 VDD1.n58 VDD1.n57 5.81868
R1916 VDD1.n165 VDD1.n164 5.81868
R1917 VDD1.n172 VDD1.n131 5.81868
R1918 VDD1.n211 VDD1.n111 5.81868
R1919 VDD1.n101 VDD1.n4 5.04292
R1920 VDD1.n66 VDD1.n22 5.04292
R1921 VDD1.n54 VDD1.n28 5.04292
R1922 VDD1.n161 VDD1.n135 5.04292
R1923 VDD1.n173 VDD1.n129 5.04292
R1924 VDD1.n210 VDD1.n113 5.04292
R1925 VDD1.n98 VDD1.n97 4.26717
R1926 VDD1.n70 VDD1.n69 4.26717
R1927 VDD1.n53 VDD1.n30 4.26717
R1928 VDD1.n160 VDD1.n137 4.26717
R1929 VDD1.n177 VDD1.n176 4.26717
R1930 VDD1.n207 VDD1.n206 4.26717
R1931 VDD1.n37 VDD1.n35 3.70982
R1932 VDD1.n144 VDD1.n142 3.70982
R1933 VDD1.n94 VDD1.n6 3.49141
R1934 VDD1.n73 VDD1.n20 3.49141
R1935 VDD1.n50 VDD1.n49 3.49141
R1936 VDD1.n157 VDD1.n156 3.49141
R1937 VDD1.n180 VDD1.n127 3.49141
R1938 VDD1.n203 VDD1.n115 3.49141
R1939 VDD1.n93 VDD1.n8 2.71565
R1940 VDD1.n74 VDD1.n18 2.71565
R1941 VDD1.n46 VDD1.n32 2.71565
R1942 VDD1.n153 VDD1.n139 2.71565
R1943 VDD1.n181 VDD1.n125 2.71565
R1944 VDD1.n202 VDD1.n117 2.71565
R1945 VDD1.n90 VDD1.n89 1.93989
R1946 VDD1.n78 VDD1.n77 1.93989
R1947 VDD1.n45 VDD1.n34 1.93989
R1948 VDD1.n152 VDD1.n141 1.93989
R1949 VDD1.n186 VDD1.n184 1.93989
R1950 VDD1.n199 VDD1.n198 1.93989
R1951 VDD1.n86 VDD1.n10 1.16414
R1952 VDD1.n81 VDD1.n15 1.16414
R1953 VDD1.n42 VDD1.n41 1.16414
R1954 VDD1.n149 VDD1.n148 1.16414
R1955 VDD1.n185 VDD1.n123 1.16414
R1956 VDD1.n195 VDD1.n119 1.16414
R1957 VDD1.n85 VDD1.n12 0.388379
R1958 VDD1.n82 VDD1.n14 0.388379
R1959 VDD1.n38 VDD1.n36 0.388379
R1960 VDD1.n145 VDD1.n143 0.388379
R1961 VDD1.n191 VDD1.n190 0.388379
R1962 VDD1.n194 VDD1.n121 0.388379
R1963 VDD1.n107 VDD1.n1 0.155672
R1964 VDD1.n100 VDD1.n1 0.155672
R1965 VDD1.n100 VDD1.n99 0.155672
R1966 VDD1.n99 VDD1.n5 0.155672
R1967 VDD1.n92 VDD1.n5 0.155672
R1968 VDD1.n92 VDD1.n91 0.155672
R1969 VDD1.n91 VDD1.n9 0.155672
R1970 VDD1.n84 VDD1.n9 0.155672
R1971 VDD1.n84 VDD1.n83 0.155672
R1972 VDD1.n83 VDD1.n13 0.155672
R1973 VDD1.n76 VDD1.n13 0.155672
R1974 VDD1.n76 VDD1.n75 0.155672
R1975 VDD1.n75 VDD1.n19 0.155672
R1976 VDD1.n68 VDD1.n19 0.155672
R1977 VDD1.n68 VDD1.n67 0.155672
R1978 VDD1.n67 VDD1.n23 0.155672
R1979 VDD1.n60 VDD1.n23 0.155672
R1980 VDD1.n60 VDD1.n59 0.155672
R1981 VDD1.n59 VDD1.n27 0.155672
R1982 VDD1.n52 VDD1.n27 0.155672
R1983 VDD1.n52 VDD1.n51 0.155672
R1984 VDD1.n51 VDD1.n31 0.155672
R1985 VDD1.n44 VDD1.n31 0.155672
R1986 VDD1.n44 VDD1.n43 0.155672
R1987 VDD1.n43 VDD1.n35 0.155672
R1988 VDD1.n150 VDD1.n142 0.155672
R1989 VDD1.n151 VDD1.n150 0.155672
R1990 VDD1.n151 VDD1.n138 0.155672
R1991 VDD1.n158 VDD1.n138 0.155672
R1992 VDD1.n159 VDD1.n158 0.155672
R1993 VDD1.n159 VDD1.n134 0.155672
R1994 VDD1.n166 VDD1.n134 0.155672
R1995 VDD1.n167 VDD1.n166 0.155672
R1996 VDD1.n167 VDD1.n130 0.155672
R1997 VDD1.n174 VDD1.n130 0.155672
R1998 VDD1.n175 VDD1.n174 0.155672
R1999 VDD1.n175 VDD1.n126 0.155672
R2000 VDD1.n182 VDD1.n126 0.155672
R2001 VDD1.n183 VDD1.n182 0.155672
R2002 VDD1.n183 VDD1.n122 0.155672
R2003 VDD1.n192 VDD1.n122 0.155672
R2004 VDD1.n193 VDD1.n192 0.155672
R2005 VDD1.n193 VDD1.n118 0.155672
R2006 VDD1.n200 VDD1.n118 0.155672
R2007 VDD1.n201 VDD1.n200 0.155672
R2008 VDD1.n201 VDD1.n114 0.155672
R2009 VDD1.n208 VDD1.n114 0.155672
R2010 VDD1.n209 VDD1.n208 0.155672
R2011 VDD1.n209 VDD1.n110 0.155672
R2012 VDD1.n216 VDD1.n110 0.155672
R2013 VN VN.t0 1235.7
R2014 VN VN.t1 1190.42
R2015 VDD2.n213 VDD2.n109 756.745
R2016 VDD2.n104 VDD2.n0 756.745
R2017 VDD2.n214 VDD2.n213 585
R2018 VDD2.n212 VDD2.n211 585
R2019 VDD2.n113 VDD2.n112 585
R2020 VDD2.n206 VDD2.n205 585
R2021 VDD2.n204 VDD2.n203 585
R2022 VDD2.n117 VDD2.n116 585
R2023 VDD2.n198 VDD2.n197 585
R2024 VDD2.n196 VDD2.n195 585
R2025 VDD2.n121 VDD2.n120 585
R2026 VDD2.n125 VDD2.n123 585
R2027 VDD2.n190 VDD2.n189 585
R2028 VDD2.n188 VDD2.n187 585
R2029 VDD2.n127 VDD2.n126 585
R2030 VDD2.n182 VDD2.n181 585
R2031 VDD2.n180 VDD2.n179 585
R2032 VDD2.n131 VDD2.n130 585
R2033 VDD2.n174 VDD2.n173 585
R2034 VDD2.n172 VDD2.n171 585
R2035 VDD2.n135 VDD2.n134 585
R2036 VDD2.n166 VDD2.n165 585
R2037 VDD2.n164 VDD2.n163 585
R2038 VDD2.n139 VDD2.n138 585
R2039 VDD2.n158 VDD2.n157 585
R2040 VDD2.n156 VDD2.n155 585
R2041 VDD2.n143 VDD2.n142 585
R2042 VDD2.n150 VDD2.n149 585
R2043 VDD2.n148 VDD2.n147 585
R2044 VDD2.n37 VDD2.n36 585
R2045 VDD2.n39 VDD2.n38 585
R2046 VDD2.n32 VDD2.n31 585
R2047 VDD2.n45 VDD2.n44 585
R2048 VDD2.n47 VDD2.n46 585
R2049 VDD2.n28 VDD2.n27 585
R2050 VDD2.n53 VDD2.n52 585
R2051 VDD2.n55 VDD2.n54 585
R2052 VDD2.n24 VDD2.n23 585
R2053 VDD2.n61 VDD2.n60 585
R2054 VDD2.n63 VDD2.n62 585
R2055 VDD2.n20 VDD2.n19 585
R2056 VDD2.n69 VDD2.n68 585
R2057 VDD2.n71 VDD2.n70 585
R2058 VDD2.n16 VDD2.n15 585
R2059 VDD2.n78 VDD2.n77 585
R2060 VDD2.n79 VDD2.n14 585
R2061 VDD2.n81 VDD2.n80 585
R2062 VDD2.n12 VDD2.n11 585
R2063 VDD2.n87 VDD2.n86 585
R2064 VDD2.n89 VDD2.n88 585
R2065 VDD2.n8 VDD2.n7 585
R2066 VDD2.n95 VDD2.n94 585
R2067 VDD2.n97 VDD2.n96 585
R2068 VDD2.n4 VDD2.n3 585
R2069 VDD2.n103 VDD2.n102 585
R2070 VDD2.n105 VDD2.n104 585
R2071 VDD2.n146 VDD2.t1 327.466
R2072 VDD2.n35 VDD2.t0 327.466
R2073 VDD2.n213 VDD2.n212 171.744
R2074 VDD2.n212 VDD2.n112 171.744
R2075 VDD2.n205 VDD2.n112 171.744
R2076 VDD2.n205 VDD2.n204 171.744
R2077 VDD2.n204 VDD2.n116 171.744
R2078 VDD2.n197 VDD2.n116 171.744
R2079 VDD2.n197 VDD2.n196 171.744
R2080 VDD2.n196 VDD2.n120 171.744
R2081 VDD2.n125 VDD2.n120 171.744
R2082 VDD2.n189 VDD2.n125 171.744
R2083 VDD2.n189 VDD2.n188 171.744
R2084 VDD2.n188 VDD2.n126 171.744
R2085 VDD2.n181 VDD2.n126 171.744
R2086 VDD2.n181 VDD2.n180 171.744
R2087 VDD2.n180 VDD2.n130 171.744
R2088 VDD2.n173 VDD2.n130 171.744
R2089 VDD2.n173 VDD2.n172 171.744
R2090 VDD2.n172 VDD2.n134 171.744
R2091 VDD2.n165 VDD2.n134 171.744
R2092 VDD2.n165 VDD2.n164 171.744
R2093 VDD2.n164 VDD2.n138 171.744
R2094 VDD2.n157 VDD2.n138 171.744
R2095 VDD2.n157 VDD2.n156 171.744
R2096 VDD2.n156 VDD2.n142 171.744
R2097 VDD2.n149 VDD2.n142 171.744
R2098 VDD2.n149 VDD2.n148 171.744
R2099 VDD2.n38 VDD2.n37 171.744
R2100 VDD2.n38 VDD2.n31 171.744
R2101 VDD2.n45 VDD2.n31 171.744
R2102 VDD2.n46 VDD2.n45 171.744
R2103 VDD2.n46 VDD2.n27 171.744
R2104 VDD2.n53 VDD2.n27 171.744
R2105 VDD2.n54 VDD2.n53 171.744
R2106 VDD2.n54 VDD2.n23 171.744
R2107 VDD2.n61 VDD2.n23 171.744
R2108 VDD2.n62 VDD2.n61 171.744
R2109 VDD2.n62 VDD2.n19 171.744
R2110 VDD2.n69 VDD2.n19 171.744
R2111 VDD2.n70 VDD2.n69 171.744
R2112 VDD2.n70 VDD2.n15 171.744
R2113 VDD2.n78 VDD2.n15 171.744
R2114 VDD2.n79 VDD2.n78 171.744
R2115 VDD2.n80 VDD2.n79 171.744
R2116 VDD2.n80 VDD2.n11 171.744
R2117 VDD2.n87 VDD2.n11 171.744
R2118 VDD2.n88 VDD2.n87 171.744
R2119 VDD2.n88 VDD2.n7 171.744
R2120 VDD2.n95 VDD2.n7 171.744
R2121 VDD2.n96 VDD2.n95 171.744
R2122 VDD2.n96 VDD2.n3 171.744
R2123 VDD2.n103 VDD2.n3 171.744
R2124 VDD2.n104 VDD2.n103 171.744
R2125 VDD2.n218 VDD2.n108 91.7476
R2126 VDD2.n148 VDD2.t1 85.8723
R2127 VDD2.n37 VDD2.t0 85.8723
R2128 VDD2.n218 VDD2.n217 49.6399
R2129 VDD2.n147 VDD2.n146 16.3895
R2130 VDD2.n36 VDD2.n35 16.3895
R2131 VDD2.n123 VDD2.n121 13.1884
R2132 VDD2.n81 VDD2.n12 13.1884
R2133 VDD2.n195 VDD2.n194 12.8005
R2134 VDD2.n191 VDD2.n190 12.8005
R2135 VDD2.n150 VDD2.n145 12.8005
R2136 VDD2.n39 VDD2.n34 12.8005
R2137 VDD2.n82 VDD2.n14 12.8005
R2138 VDD2.n86 VDD2.n85 12.8005
R2139 VDD2.n198 VDD2.n119 12.0247
R2140 VDD2.n187 VDD2.n124 12.0247
R2141 VDD2.n151 VDD2.n143 12.0247
R2142 VDD2.n40 VDD2.n32 12.0247
R2143 VDD2.n77 VDD2.n76 12.0247
R2144 VDD2.n89 VDD2.n10 12.0247
R2145 VDD2.n199 VDD2.n117 11.249
R2146 VDD2.n186 VDD2.n127 11.249
R2147 VDD2.n155 VDD2.n154 11.249
R2148 VDD2.n44 VDD2.n43 11.249
R2149 VDD2.n75 VDD2.n16 11.249
R2150 VDD2.n90 VDD2.n8 11.249
R2151 VDD2.n203 VDD2.n202 10.4732
R2152 VDD2.n183 VDD2.n182 10.4732
R2153 VDD2.n158 VDD2.n141 10.4732
R2154 VDD2.n47 VDD2.n30 10.4732
R2155 VDD2.n72 VDD2.n71 10.4732
R2156 VDD2.n94 VDD2.n93 10.4732
R2157 VDD2.n206 VDD2.n115 9.69747
R2158 VDD2.n179 VDD2.n129 9.69747
R2159 VDD2.n159 VDD2.n139 9.69747
R2160 VDD2.n48 VDD2.n28 9.69747
R2161 VDD2.n68 VDD2.n18 9.69747
R2162 VDD2.n97 VDD2.n6 9.69747
R2163 VDD2.n217 VDD2.n216 9.45567
R2164 VDD2.n108 VDD2.n107 9.45567
R2165 VDD2.n133 VDD2.n132 9.3005
R2166 VDD2.n176 VDD2.n175 9.3005
R2167 VDD2.n178 VDD2.n177 9.3005
R2168 VDD2.n129 VDD2.n128 9.3005
R2169 VDD2.n184 VDD2.n183 9.3005
R2170 VDD2.n186 VDD2.n185 9.3005
R2171 VDD2.n124 VDD2.n122 9.3005
R2172 VDD2.n192 VDD2.n191 9.3005
R2173 VDD2.n216 VDD2.n215 9.3005
R2174 VDD2.n111 VDD2.n110 9.3005
R2175 VDD2.n210 VDD2.n209 9.3005
R2176 VDD2.n208 VDD2.n207 9.3005
R2177 VDD2.n115 VDD2.n114 9.3005
R2178 VDD2.n202 VDD2.n201 9.3005
R2179 VDD2.n200 VDD2.n199 9.3005
R2180 VDD2.n119 VDD2.n118 9.3005
R2181 VDD2.n194 VDD2.n193 9.3005
R2182 VDD2.n170 VDD2.n169 9.3005
R2183 VDD2.n168 VDD2.n167 9.3005
R2184 VDD2.n137 VDD2.n136 9.3005
R2185 VDD2.n162 VDD2.n161 9.3005
R2186 VDD2.n160 VDD2.n159 9.3005
R2187 VDD2.n141 VDD2.n140 9.3005
R2188 VDD2.n154 VDD2.n153 9.3005
R2189 VDD2.n152 VDD2.n151 9.3005
R2190 VDD2.n145 VDD2.n144 9.3005
R2191 VDD2.n107 VDD2.n106 9.3005
R2192 VDD2.n101 VDD2.n100 9.3005
R2193 VDD2.n99 VDD2.n98 9.3005
R2194 VDD2.n6 VDD2.n5 9.3005
R2195 VDD2.n93 VDD2.n92 9.3005
R2196 VDD2.n91 VDD2.n90 9.3005
R2197 VDD2.n10 VDD2.n9 9.3005
R2198 VDD2.n85 VDD2.n84 9.3005
R2199 VDD2.n57 VDD2.n56 9.3005
R2200 VDD2.n26 VDD2.n25 9.3005
R2201 VDD2.n51 VDD2.n50 9.3005
R2202 VDD2.n49 VDD2.n48 9.3005
R2203 VDD2.n30 VDD2.n29 9.3005
R2204 VDD2.n43 VDD2.n42 9.3005
R2205 VDD2.n41 VDD2.n40 9.3005
R2206 VDD2.n34 VDD2.n33 9.3005
R2207 VDD2.n59 VDD2.n58 9.3005
R2208 VDD2.n22 VDD2.n21 9.3005
R2209 VDD2.n65 VDD2.n64 9.3005
R2210 VDD2.n67 VDD2.n66 9.3005
R2211 VDD2.n18 VDD2.n17 9.3005
R2212 VDD2.n73 VDD2.n72 9.3005
R2213 VDD2.n75 VDD2.n74 9.3005
R2214 VDD2.n76 VDD2.n13 9.3005
R2215 VDD2.n83 VDD2.n82 9.3005
R2216 VDD2.n2 VDD2.n1 9.3005
R2217 VDD2.n207 VDD2.n113 8.92171
R2218 VDD2.n178 VDD2.n131 8.92171
R2219 VDD2.n163 VDD2.n162 8.92171
R2220 VDD2.n52 VDD2.n51 8.92171
R2221 VDD2.n67 VDD2.n20 8.92171
R2222 VDD2.n98 VDD2.n4 8.92171
R2223 VDD2.n211 VDD2.n210 8.14595
R2224 VDD2.n175 VDD2.n174 8.14595
R2225 VDD2.n166 VDD2.n137 8.14595
R2226 VDD2.n55 VDD2.n26 8.14595
R2227 VDD2.n64 VDD2.n63 8.14595
R2228 VDD2.n102 VDD2.n101 8.14595
R2229 VDD2.n217 VDD2.n109 7.3702
R2230 VDD2.n214 VDD2.n111 7.3702
R2231 VDD2.n171 VDD2.n133 7.3702
R2232 VDD2.n167 VDD2.n135 7.3702
R2233 VDD2.n56 VDD2.n24 7.3702
R2234 VDD2.n60 VDD2.n22 7.3702
R2235 VDD2.n105 VDD2.n2 7.3702
R2236 VDD2.n108 VDD2.n0 7.3702
R2237 VDD2.n215 VDD2.n109 6.59444
R2238 VDD2.n215 VDD2.n214 6.59444
R2239 VDD2.n171 VDD2.n170 6.59444
R2240 VDD2.n170 VDD2.n135 6.59444
R2241 VDD2.n59 VDD2.n24 6.59444
R2242 VDD2.n60 VDD2.n59 6.59444
R2243 VDD2.n106 VDD2.n105 6.59444
R2244 VDD2.n106 VDD2.n0 6.59444
R2245 VDD2.n211 VDD2.n111 5.81868
R2246 VDD2.n174 VDD2.n133 5.81868
R2247 VDD2.n167 VDD2.n166 5.81868
R2248 VDD2.n56 VDD2.n55 5.81868
R2249 VDD2.n63 VDD2.n22 5.81868
R2250 VDD2.n102 VDD2.n2 5.81868
R2251 VDD2.n210 VDD2.n113 5.04292
R2252 VDD2.n175 VDD2.n131 5.04292
R2253 VDD2.n163 VDD2.n137 5.04292
R2254 VDD2.n52 VDD2.n26 5.04292
R2255 VDD2.n64 VDD2.n20 5.04292
R2256 VDD2.n101 VDD2.n4 5.04292
R2257 VDD2.n207 VDD2.n206 4.26717
R2258 VDD2.n179 VDD2.n178 4.26717
R2259 VDD2.n162 VDD2.n139 4.26717
R2260 VDD2.n51 VDD2.n28 4.26717
R2261 VDD2.n68 VDD2.n67 4.26717
R2262 VDD2.n98 VDD2.n97 4.26717
R2263 VDD2.n146 VDD2.n144 3.70982
R2264 VDD2.n35 VDD2.n33 3.70982
R2265 VDD2.n203 VDD2.n115 3.49141
R2266 VDD2.n182 VDD2.n129 3.49141
R2267 VDD2.n159 VDD2.n158 3.49141
R2268 VDD2.n48 VDD2.n47 3.49141
R2269 VDD2.n71 VDD2.n18 3.49141
R2270 VDD2.n94 VDD2.n6 3.49141
R2271 VDD2.n202 VDD2.n117 2.71565
R2272 VDD2.n183 VDD2.n127 2.71565
R2273 VDD2.n155 VDD2.n141 2.71565
R2274 VDD2.n44 VDD2.n30 2.71565
R2275 VDD2.n72 VDD2.n16 2.71565
R2276 VDD2.n93 VDD2.n8 2.71565
R2277 VDD2.n199 VDD2.n198 1.93989
R2278 VDD2.n187 VDD2.n186 1.93989
R2279 VDD2.n154 VDD2.n143 1.93989
R2280 VDD2.n43 VDD2.n32 1.93989
R2281 VDD2.n77 VDD2.n75 1.93989
R2282 VDD2.n90 VDD2.n89 1.93989
R2283 VDD2.n195 VDD2.n119 1.16414
R2284 VDD2.n190 VDD2.n124 1.16414
R2285 VDD2.n151 VDD2.n150 1.16414
R2286 VDD2.n40 VDD2.n39 1.16414
R2287 VDD2.n76 VDD2.n14 1.16414
R2288 VDD2.n86 VDD2.n10 1.16414
R2289 VDD2.n194 VDD2.n121 0.388379
R2290 VDD2.n191 VDD2.n123 0.388379
R2291 VDD2.n147 VDD2.n145 0.388379
R2292 VDD2.n36 VDD2.n34 0.388379
R2293 VDD2.n82 VDD2.n81 0.388379
R2294 VDD2.n85 VDD2.n12 0.388379
R2295 VDD2 VDD2.n218 0.237569
R2296 VDD2.n216 VDD2.n110 0.155672
R2297 VDD2.n209 VDD2.n110 0.155672
R2298 VDD2.n209 VDD2.n208 0.155672
R2299 VDD2.n208 VDD2.n114 0.155672
R2300 VDD2.n201 VDD2.n114 0.155672
R2301 VDD2.n201 VDD2.n200 0.155672
R2302 VDD2.n200 VDD2.n118 0.155672
R2303 VDD2.n193 VDD2.n118 0.155672
R2304 VDD2.n193 VDD2.n192 0.155672
R2305 VDD2.n192 VDD2.n122 0.155672
R2306 VDD2.n185 VDD2.n122 0.155672
R2307 VDD2.n185 VDD2.n184 0.155672
R2308 VDD2.n184 VDD2.n128 0.155672
R2309 VDD2.n177 VDD2.n128 0.155672
R2310 VDD2.n177 VDD2.n176 0.155672
R2311 VDD2.n176 VDD2.n132 0.155672
R2312 VDD2.n169 VDD2.n132 0.155672
R2313 VDD2.n169 VDD2.n168 0.155672
R2314 VDD2.n168 VDD2.n136 0.155672
R2315 VDD2.n161 VDD2.n136 0.155672
R2316 VDD2.n161 VDD2.n160 0.155672
R2317 VDD2.n160 VDD2.n140 0.155672
R2318 VDD2.n153 VDD2.n140 0.155672
R2319 VDD2.n153 VDD2.n152 0.155672
R2320 VDD2.n152 VDD2.n144 0.155672
R2321 VDD2.n41 VDD2.n33 0.155672
R2322 VDD2.n42 VDD2.n41 0.155672
R2323 VDD2.n42 VDD2.n29 0.155672
R2324 VDD2.n49 VDD2.n29 0.155672
R2325 VDD2.n50 VDD2.n49 0.155672
R2326 VDD2.n50 VDD2.n25 0.155672
R2327 VDD2.n57 VDD2.n25 0.155672
R2328 VDD2.n58 VDD2.n57 0.155672
R2329 VDD2.n58 VDD2.n21 0.155672
R2330 VDD2.n65 VDD2.n21 0.155672
R2331 VDD2.n66 VDD2.n65 0.155672
R2332 VDD2.n66 VDD2.n17 0.155672
R2333 VDD2.n73 VDD2.n17 0.155672
R2334 VDD2.n74 VDD2.n73 0.155672
R2335 VDD2.n74 VDD2.n13 0.155672
R2336 VDD2.n83 VDD2.n13 0.155672
R2337 VDD2.n84 VDD2.n83 0.155672
R2338 VDD2.n84 VDD2.n9 0.155672
R2339 VDD2.n91 VDD2.n9 0.155672
R2340 VDD2.n92 VDD2.n91 0.155672
R2341 VDD2.n92 VDD2.n5 0.155672
R2342 VDD2.n99 VDD2.n5 0.155672
R2343 VDD2.n100 VDD2.n99 0.155672
R2344 VDD2.n100 VDD2.n1 0.155672
R2345 VDD2.n107 VDD2.n1 0.155672
C0 VN w_n1302_n4916# 1.7694f
C1 VDD2 VN 2.73241f
C2 VDD1 B 1.93083f
C3 B w_n1302_n4916# 8.707769f
C4 VDD1 VP 2.82428f
C5 VDD2 B 1.944f
C6 VP w_n1302_n4916# 1.93072f
C7 VDD2 VP 0.248312f
C8 VDD1 w_n1302_n4916# 2.12651f
C9 VN VTAIL 1.83521f
C10 VDD1 VDD2 0.4461f
C11 VDD2 w_n1302_n4916# 2.12915f
C12 VTAIL B 3.96618f
C13 VTAIL VP 1.85025f
C14 VN B 0.785398f
C15 VN VP 5.89891f
C16 VDD1 VTAIL 9.28388f
C17 VTAIL w_n1302_n4916# 4.28169f
C18 VDD2 VTAIL 9.31067f
C19 VDD1 VN 0.148831f
C20 B VP 1.04219f
C21 VDD2 VSUBS 1.006098f
C22 VDD1 VSUBS 4.70164f
C23 VTAIL VSUBS 0.258778f
C24 VN VSUBS 7.38771f
C25 VP VSUBS 1.340962f
C26 B VSUBS 3.003082f
C27 w_n1302_n4916# VSUBS 78.1669f
C28 VDD2.n0 VSUBS 0.029051f
C29 VDD2.n1 VSUBS 0.025362f
C30 VDD2.n2 VSUBS 0.013628f
C31 VDD2.n3 VSUBS 0.032212f
C32 VDD2.n4 VSUBS 0.01443f
C33 VDD2.n5 VSUBS 0.025362f
C34 VDD2.n6 VSUBS 0.013628f
C35 VDD2.n7 VSUBS 0.032212f
C36 VDD2.n8 VSUBS 0.01443f
C37 VDD2.n9 VSUBS 0.025362f
C38 VDD2.n10 VSUBS 0.013628f
C39 VDD2.n11 VSUBS 0.032212f
C40 VDD2.n12 VSUBS 0.014029f
C41 VDD2.n13 VSUBS 0.025362f
C42 VDD2.n14 VSUBS 0.01443f
C43 VDD2.n15 VSUBS 0.032212f
C44 VDD2.n16 VSUBS 0.01443f
C45 VDD2.n17 VSUBS 0.025362f
C46 VDD2.n18 VSUBS 0.013628f
C47 VDD2.n19 VSUBS 0.032212f
C48 VDD2.n20 VSUBS 0.01443f
C49 VDD2.n21 VSUBS 0.025362f
C50 VDD2.n22 VSUBS 0.013628f
C51 VDD2.n23 VSUBS 0.032212f
C52 VDD2.n24 VSUBS 0.01443f
C53 VDD2.n25 VSUBS 0.025362f
C54 VDD2.n26 VSUBS 0.013628f
C55 VDD2.n27 VSUBS 0.032212f
C56 VDD2.n28 VSUBS 0.01443f
C57 VDD2.n29 VSUBS 0.025362f
C58 VDD2.n30 VSUBS 0.013628f
C59 VDD2.n31 VSUBS 0.032212f
C60 VDD2.n32 VSUBS 0.01443f
C61 VDD2.n33 VSUBS 2.16284f
C62 VDD2.n34 VSUBS 0.013628f
C63 VDD2.t0 VSUBS 0.069258f
C64 VDD2.n35 VSUBS 0.214087f
C65 VDD2.n36 VSUBS 0.020492f
C66 VDD2.n37 VSUBS 0.024159f
C67 VDD2.n38 VSUBS 0.032212f
C68 VDD2.n39 VSUBS 0.01443f
C69 VDD2.n40 VSUBS 0.013628f
C70 VDD2.n41 VSUBS 0.025362f
C71 VDD2.n42 VSUBS 0.025362f
C72 VDD2.n43 VSUBS 0.013628f
C73 VDD2.n44 VSUBS 0.01443f
C74 VDD2.n45 VSUBS 0.032212f
C75 VDD2.n46 VSUBS 0.032212f
C76 VDD2.n47 VSUBS 0.01443f
C77 VDD2.n48 VSUBS 0.013628f
C78 VDD2.n49 VSUBS 0.025362f
C79 VDD2.n50 VSUBS 0.025362f
C80 VDD2.n51 VSUBS 0.013628f
C81 VDD2.n52 VSUBS 0.01443f
C82 VDD2.n53 VSUBS 0.032212f
C83 VDD2.n54 VSUBS 0.032212f
C84 VDD2.n55 VSUBS 0.01443f
C85 VDD2.n56 VSUBS 0.013628f
C86 VDD2.n57 VSUBS 0.025362f
C87 VDD2.n58 VSUBS 0.025362f
C88 VDD2.n59 VSUBS 0.013628f
C89 VDD2.n60 VSUBS 0.01443f
C90 VDD2.n61 VSUBS 0.032212f
C91 VDD2.n62 VSUBS 0.032212f
C92 VDD2.n63 VSUBS 0.01443f
C93 VDD2.n64 VSUBS 0.013628f
C94 VDD2.n65 VSUBS 0.025362f
C95 VDD2.n66 VSUBS 0.025362f
C96 VDD2.n67 VSUBS 0.013628f
C97 VDD2.n68 VSUBS 0.01443f
C98 VDD2.n69 VSUBS 0.032212f
C99 VDD2.n70 VSUBS 0.032212f
C100 VDD2.n71 VSUBS 0.01443f
C101 VDD2.n72 VSUBS 0.013628f
C102 VDD2.n73 VSUBS 0.025362f
C103 VDD2.n74 VSUBS 0.025362f
C104 VDD2.n75 VSUBS 0.013628f
C105 VDD2.n76 VSUBS 0.013628f
C106 VDD2.n77 VSUBS 0.01443f
C107 VDD2.n78 VSUBS 0.032212f
C108 VDD2.n79 VSUBS 0.032212f
C109 VDD2.n80 VSUBS 0.032212f
C110 VDD2.n81 VSUBS 0.014029f
C111 VDD2.n82 VSUBS 0.013628f
C112 VDD2.n83 VSUBS 0.025362f
C113 VDD2.n84 VSUBS 0.025362f
C114 VDD2.n85 VSUBS 0.013628f
C115 VDD2.n86 VSUBS 0.01443f
C116 VDD2.n87 VSUBS 0.032212f
C117 VDD2.n88 VSUBS 0.032212f
C118 VDD2.n89 VSUBS 0.01443f
C119 VDD2.n90 VSUBS 0.013628f
C120 VDD2.n91 VSUBS 0.025362f
C121 VDD2.n92 VSUBS 0.025362f
C122 VDD2.n93 VSUBS 0.013628f
C123 VDD2.n94 VSUBS 0.01443f
C124 VDD2.n95 VSUBS 0.032212f
C125 VDD2.n96 VSUBS 0.032212f
C126 VDD2.n97 VSUBS 0.01443f
C127 VDD2.n98 VSUBS 0.013628f
C128 VDD2.n99 VSUBS 0.025362f
C129 VDD2.n100 VSUBS 0.025362f
C130 VDD2.n101 VSUBS 0.013628f
C131 VDD2.n102 VSUBS 0.01443f
C132 VDD2.n103 VSUBS 0.032212f
C133 VDD2.n104 VSUBS 0.082016f
C134 VDD2.n105 VSUBS 0.01443f
C135 VDD2.n106 VSUBS 0.013628f
C136 VDD2.n107 VSUBS 0.060008f
C137 VDD2.n108 VSUBS 0.886719f
C138 VDD2.n109 VSUBS 0.029051f
C139 VDD2.n110 VSUBS 0.025362f
C140 VDD2.n111 VSUBS 0.013628f
C141 VDD2.n112 VSUBS 0.032212f
C142 VDD2.n113 VSUBS 0.01443f
C143 VDD2.n114 VSUBS 0.025362f
C144 VDD2.n115 VSUBS 0.013628f
C145 VDD2.n116 VSUBS 0.032212f
C146 VDD2.n117 VSUBS 0.01443f
C147 VDD2.n118 VSUBS 0.025362f
C148 VDD2.n119 VSUBS 0.013628f
C149 VDD2.n120 VSUBS 0.032212f
C150 VDD2.n121 VSUBS 0.014029f
C151 VDD2.n122 VSUBS 0.025362f
C152 VDD2.n123 VSUBS 0.014029f
C153 VDD2.n124 VSUBS 0.013628f
C154 VDD2.n125 VSUBS 0.032212f
C155 VDD2.n126 VSUBS 0.032212f
C156 VDD2.n127 VSUBS 0.01443f
C157 VDD2.n128 VSUBS 0.025362f
C158 VDD2.n129 VSUBS 0.013628f
C159 VDD2.n130 VSUBS 0.032212f
C160 VDD2.n131 VSUBS 0.01443f
C161 VDD2.n132 VSUBS 0.025362f
C162 VDD2.n133 VSUBS 0.013628f
C163 VDD2.n134 VSUBS 0.032212f
C164 VDD2.n135 VSUBS 0.01443f
C165 VDD2.n136 VSUBS 0.025362f
C166 VDD2.n137 VSUBS 0.013628f
C167 VDD2.n138 VSUBS 0.032212f
C168 VDD2.n139 VSUBS 0.01443f
C169 VDD2.n140 VSUBS 0.025362f
C170 VDD2.n141 VSUBS 0.013628f
C171 VDD2.n142 VSUBS 0.032212f
C172 VDD2.n143 VSUBS 0.01443f
C173 VDD2.n144 VSUBS 2.16284f
C174 VDD2.n145 VSUBS 0.013628f
C175 VDD2.t1 VSUBS 0.069258f
C176 VDD2.n146 VSUBS 0.214087f
C177 VDD2.n147 VSUBS 0.020492f
C178 VDD2.n148 VSUBS 0.024159f
C179 VDD2.n149 VSUBS 0.032212f
C180 VDD2.n150 VSUBS 0.01443f
C181 VDD2.n151 VSUBS 0.013628f
C182 VDD2.n152 VSUBS 0.025362f
C183 VDD2.n153 VSUBS 0.025362f
C184 VDD2.n154 VSUBS 0.013628f
C185 VDD2.n155 VSUBS 0.01443f
C186 VDD2.n156 VSUBS 0.032212f
C187 VDD2.n157 VSUBS 0.032212f
C188 VDD2.n158 VSUBS 0.01443f
C189 VDD2.n159 VSUBS 0.013628f
C190 VDD2.n160 VSUBS 0.025362f
C191 VDD2.n161 VSUBS 0.025362f
C192 VDD2.n162 VSUBS 0.013628f
C193 VDD2.n163 VSUBS 0.01443f
C194 VDD2.n164 VSUBS 0.032212f
C195 VDD2.n165 VSUBS 0.032212f
C196 VDD2.n166 VSUBS 0.01443f
C197 VDD2.n167 VSUBS 0.013628f
C198 VDD2.n168 VSUBS 0.025362f
C199 VDD2.n169 VSUBS 0.025362f
C200 VDD2.n170 VSUBS 0.013628f
C201 VDD2.n171 VSUBS 0.01443f
C202 VDD2.n172 VSUBS 0.032212f
C203 VDD2.n173 VSUBS 0.032212f
C204 VDD2.n174 VSUBS 0.01443f
C205 VDD2.n175 VSUBS 0.013628f
C206 VDD2.n176 VSUBS 0.025362f
C207 VDD2.n177 VSUBS 0.025362f
C208 VDD2.n178 VSUBS 0.013628f
C209 VDD2.n179 VSUBS 0.01443f
C210 VDD2.n180 VSUBS 0.032212f
C211 VDD2.n181 VSUBS 0.032212f
C212 VDD2.n182 VSUBS 0.01443f
C213 VDD2.n183 VSUBS 0.013628f
C214 VDD2.n184 VSUBS 0.025362f
C215 VDD2.n185 VSUBS 0.025362f
C216 VDD2.n186 VSUBS 0.013628f
C217 VDD2.n187 VSUBS 0.01443f
C218 VDD2.n188 VSUBS 0.032212f
C219 VDD2.n189 VSUBS 0.032212f
C220 VDD2.n190 VSUBS 0.01443f
C221 VDD2.n191 VSUBS 0.013628f
C222 VDD2.n192 VSUBS 0.025362f
C223 VDD2.n193 VSUBS 0.025362f
C224 VDD2.n194 VSUBS 0.013628f
C225 VDD2.n195 VSUBS 0.01443f
C226 VDD2.n196 VSUBS 0.032212f
C227 VDD2.n197 VSUBS 0.032212f
C228 VDD2.n198 VSUBS 0.01443f
C229 VDD2.n199 VSUBS 0.013628f
C230 VDD2.n200 VSUBS 0.025362f
C231 VDD2.n201 VSUBS 0.025362f
C232 VDD2.n202 VSUBS 0.013628f
C233 VDD2.n203 VSUBS 0.01443f
C234 VDD2.n204 VSUBS 0.032212f
C235 VDD2.n205 VSUBS 0.032212f
C236 VDD2.n206 VSUBS 0.01443f
C237 VDD2.n207 VSUBS 0.013628f
C238 VDD2.n208 VSUBS 0.025362f
C239 VDD2.n209 VSUBS 0.025362f
C240 VDD2.n210 VSUBS 0.013628f
C241 VDD2.n211 VSUBS 0.01443f
C242 VDD2.n212 VSUBS 0.032212f
C243 VDD2.n213 VSUBS 0.082016f
C244 VDD2.n214 VSUBS 0.01443f
C245 VDD2.n215 VSUBS 0.013628f
C246 VDD2.n216 VSUBS 0.060008f
C247 VDD2.n217 VSUBS 0.058967f
C248 VDD2.n218 VSUBS 3.49576f
C249 VN.t1 VSUBS 1.47574f
C250 VN.t0 VSUBS 1.57849f
C251 VDD1.n0 VSUBS 0.029064f
C252 VDD1.n1 VSUBS 0.025373f
C253 VDD1.n2 VSUBS 0.013634f
C254 VDD1.n3 VSUBS 0.032227f
C255 VDD1.n4 VSUBS 0.014436f
C256 VDD1.n5 VSUBS 0.025373f
C257 VDD1.n6 VSUBS 0.013634f
C258 VDD1.n7 VSUBS 0.032227f
C259 VDD1.n8 VSUBS 0.014436f
C260 VDD1.n9 VSUBS 0.025373f
C261 VDD1.n10 VSUBS 0.013634f
C262 VDD1.n11 VSUBS 0.032227f
C263 VDD1.n12 VSUBS 0.014035f
C264 VDD1.n13 VSUBS 0.025373f
C265 VDD1.n14 VSUBS 0.014035f
C266 VDD1.n15 VSUBS 0.013634f
C267 VDD1.n16 VSUBS 0.032227f
C268 VDD1.n17 VSUBS 0.032227f
C269 VDD1.n18 VSUBS 0.014436f
C270 VDD1.n19 VSUBS 0.025373f
C271 VDD1.n20 VSUBS 0.013634f
C272 VDD1.n21 VSUBS 0.032227f
C273 VDD1.n22 VSUBS 0.014436f
C274 VDD1.n23 VSUBS 0.025373f
C275 VDD1.n24 VSUBS 0.013634f
C276 VDD1.n25 VSUBS 0.032227f
C277 VDD1.n26 VSUBS 0.014436f
C278 VDD1.n27 VSUBS 0.025373f
C279 VDD1.n28 VSUBS 0.013634f
C280 VDD1.n29 VSUBS 0.032227f
C281 VDD1.n30 VSUBS 0.014436f
C282 VDD1.n31 VSUBS 0.025373f
C283 VDD1.n32 VSUBS 0.013634f
C284 VDD1.n33 VSUBS 0.032227f
C285 VDD1.n34 VSUBS 0.014436f
C286 VDD1.n35 VSUBS 2.1638f
C287 VDD1.n36 VSUBS 0.013634f
C288 VDD1.t1 VSUBS 0.069289f
C289 VDD1.n37 VSUBS 0.214183f
C290 VDD1.n38 VSUBS 0.020501f
C291 VDD1.n39 VSUBS 0.02417f
C292 VDD1.n40 VSUBS 0.032227f
C293 VDD1.n41 VSUBS 0.014436f
C294 VDD1.n42 VSUBS 0.013634f
C295 VDD1.n43 VSUBS 0.025373f
C296 VDD1.n44 VSUBS 0.025373f
C297 VDD1.n45 VSUBS 0.013634f
C298 VDD1.n46 VSUBS 0.014436f
C299 VDD1.n47 VSUBS 0.032227f
C300 VDD1.n48 VSUBS 0.032227f
C301 VDD1.n49 VSUBS 0.014436f
C302 VDD1.n50 VSUBS 0.013634f
C303 VDD1.n51 VSUBS 0.025373f
C304 VDD1.n52 VSUBS 0.025373f
C305 VDD1.n53 VSUBS 0.013634f
C306 VDD1.n54 VSUBS 0.014436f
C307 VDD1.n55 VSUBS 0.032227f
C308 VDD1.n56 VSUBS 0.032227f
C309 VDD1.n57 VSUBS 0.014436f
C310 VDD1.n58 VSUBS 0.013634f
C311 VDD1.n59 VSUBS 0.025373f
C312 VDD1.n60 VSUBS 0.025373f
C313 VDD1.n61 VSUBS 0.013634f
C314 VDD1.n62 VSUBS 0.014436f
C315 VDD1.n63 VSUBS 0.032227f
C316 VDD1.n64 VSUBS 0.032227f
C317 VDD1.n65 VSUBS 0.014436f
C318 VDD1.n66 VSUBS 0.013634f
C319 VDD1.n67 VSUBS 0.025373f
C320 VDD1.n68 VSUBS 0.025373f
C321 VDD1.n69 VSUBS 0.013634f
C322 VDD1.n70 VSUBS 0.014436f
C323 VDD1.n71 VSUBS 0.032227f
C324 VDD1.n72 VSUBS 0.032227f
C325 VDD1.n73 VSUBS 0.014436f
C326 VDD1.n74 VSUBS 0.013634f
C327 VDD1.n75 VSUBS 0.025373f
C328 VDD1.n76 VSUBS 0.025373f
C329 VDD1.n77 VSUBS 0.013634f
C330 VDD1.n78 VSUBS 0.014436f
C331 VDD1.n79 VSUBS 0.032227f
C332 VDD1.n80 VSUBS 0.032227f
C333 VDD1.n81 VSUBS 0.014436f
C334 VDD1.n82 VSUBS 0.013634f
C335 VDD1.n83 VSUBS 0.025373f
C336 VDD1.n84 VSUBS 0.025373f
C337 VDD1.n85 VSUBS 0.013634f
C338 VDD1.n86 VSUBS 0.014436f
C339 VDD1.n87 VSUBS 0.032227f
C340 VDD1.n88 VSUBS 0.032227f
C341 VDD1.n89 VSUBS 0.014436f
C342 VDD1.n90 VSUBS 0.013634f
C343 VDD1.n91 VSUBS 0.025373f
C344 VDD1.n92 VSUBS 0.025373f
C345 VDD1.n93 VSUBS 0.013634f
C346 VDD1.n94 VSUBS 0.014436f
C347 VDD1.n95 VSUBS 0.032227f
C348 VDD1.n96 VSUBS 0.032227f
C349 VDD1.n97 VSUBS 0.014436f
C350 VDD1.n98 VSUBS 0.013634f
C351 VDD1.n99 VSUBS 0.025373f
C352 VDD1.n100 VSUBS 0.025373f
C353 VDD1.n101 VSUBS 0.013634f
C354 VDD1.n102 VSUBS 0.014436f
C355 VDD1.n103 VSUBS 0.032227f
C356 VDD1.n104 VSUBS 0.082052f
C357 VDD1.n105 VSUBS 0.014436f
C358 VDD1.n106 VSUBS 0.013634f
C359 VDD1.n107 VSUBS 0.060035f
C360 VDD1.n108 VSUBS 0.059322f
C361 VDD1.n109 VSUBS 0.029064f
C362 VDD1.n110 VSUBS 0.025373f
C363 VDD1.n111 VSUBS 0.013634f
C364 VDD1.n112 VSUBS 0.032227f
C365 VDD1.n113 VSUBS 0.014436f
C366 VDD1.n114 VSUBS 0.025373f
C367 VDD1.n115 VSUBS 0.013634f
C368 VDD1.n116 VSUBS 0.032227f
C369 VDD1.n117 VSUBS 0.014436f
C370 VDD1.n118 VSUBS 0.025373f
C371 VDD1.n119 VSUBS 0.013634f
C372 VDD1.n120 VSUBS 0.032227f
C373 VDD1.n121 VSUBS 0.014035f
C374 VDD1.n122 VSUBS 0.025373f
C375 VDD1.n123 VSUBS 0.014436f
C376 VDD1.n124 VSUBS 0.032227f
C377 VDD1.n125 VSUBS 0.014436f
C378 VDD1.n126 VSUBS 0.025373f
C379 VDD1.n127 VSUBS 0.013634f
C380 VDD1.n128 VSUBS 0.032227f
C381 VDD1.n129 VSUBS 0.014436f
C382 VDD1.n130 VSUBS 0.025373f
C383 VDD1.n131 VSUBS 0.013634f
C384 VDD1.n132 VSUBS 0.032227f
C385 VDD1.n133 VSUBS 0.014436f
C386 VDD1.n134 VSUBS 0.025373f
C387 VDD1.n135 VSUBS 0.013634f
C388 VDD1.n136 VSUBS 0.032227f
C389 VDD1.n137 VSUBS 0.014436f
C390 VDD1.n138 VSUBS 0.025373f
C391 VDD1.n139 VSUBS 0.013634f
C392 VDD1.n140 VSUBS 0.032227f
C393 VDD1.n141 VSUBS 0.014436f
C394 VDD1.n142 VSUBS 2.1638f
C395 VDD1.n143 VSUBS 0.013634f
C396 VDD1.t0 VSUBS 0.069289f
C397 VDD1.n144 VSUBS 0.214183f
C398 VDD1.n145 VSUBS 0.020501f
C399 VDD1.n146 VSUBS 0.02417f
C400 VDD1.n147 VSUBS 0.032227f
C401 VDD1.n148 VSUBS 0.014436f
C402 VDD1.n149 VSUBS 0.013634f
C403 VDD1.n150 VSUBS 0.025373f
C404 VDD1.n151 VSUBS 0.025373f
C405 VDD1.n152 VSUBS 0.013634f
C406 VDD1.n153 VSUBS 0.014436f
C407 VDD1.n154 VSUBS 0.032227f
C408 VDD1.n155 VSUBS 0.032227f
C409 VDD1.n156 VSUBS 0.014436f
C410 VDD1.n157 VSUBS 0.013634f
C411 VDD1.n158 VSUBS 0.025373f
C412 VDD1.n159 VSUBS 0.025373f
C413 VDD1.n160 VSUBS 0.013634f
C414 VDD1.n161 VSUBS 0.014436f
C415 VDD1.n162 VSUBS 0.032227f
C416 VDD1.n163 VSUBS 0.032227f
C417 VDD1.n164 VSUBS 0.014436f
C418 VDD1.n165 VSUBS 0.013634f
C419 VDD1.n166 VSUBS 0.025373f
C420 VDD1.n167 VSUBS 0.025373f
C421 VDD1.n168 VSUBS 0.013634f
C422 VDD1.n169 VSUBS 0.014436f
C423 VDD1.n170 VSUBS 0.032227f
C424 VDD1.n171 VSUBS 0.032227f
C425 VDD1.n172 VSUBS 0.014436f
C426 VDD1.n173 VSUBS 0.013634f
C427 VDD1.n174 VSUBS 0.025373f
C428 VDD1.n175 VSUBS 0.025373f
C429 VDD1.n176 VSUBS 0.013634f
C430 VDD1.n177 VSUBS 0.014436f
C431 VDD1.n178 VSUBS 0.032227f
C432 VDD1.n179 VSUBS 0.032227f
C433 VDD1.n180 VSUBS 0.014436f
C434 VDD1.n181 VSUBS 0.013634f
C435 VDD1.n182 VSUBS 0.025373f
C436 VDD1.n183 VSUBS 0.025373f
C437 VDD1.n184 VSUBS 0.013634f
C438 VDD1.n185 VSUBS 0.013634f
C439 VDD1.n186 VSUBS 0.014436f
C440 VDD1.n187 VSUBS 0.032227f
C441 VDD1.n188 VSUBS 0.032227f
C442 VDD1.n189 VSUBS 0.032227f
C443 VDD1.n190 VSUBS 0.014035f
C444 VDD1.n191 VSUBS 0.013634f
C445 VDD1.n192 VSUBS 0.025373f
C446 VDD1.n193 VSUBS 0.025373f
C447 VDD1.n194 VSUBS 0.013634f
C448 VDD1.n195 VSUBS 0.014436f
C449 VDD1.n196 VSUBS 0.032227f
C450 VDD1.n197 VSUBS 0.032227f
C451 VDD1.n198 VSUBS 0.014436f
C452 VDD1.n199 VSUBS 0.013634f
C453 VDD1.n200 VSUBS 0.025373f
C454 VDD1.n201 VSUBS 0.025373f
C455 VDD1.n202 VSUBS 0.013634f
C456 VDD1.n203 VSUBS 0.014436f
C457 VDD1.n204 VSUBS 0.032227f
C458 VDD1.n205 VSUBS 0.032227f
C459 VDD1.n206 VSUBS 0.014436f
C460 VDD1.n207 VSUBS 0.013634f
C461 VDD1.n208 VSUBS 0.025373f
C462 VDD1.n209 VSUBS 0.025373f
C463 VDD1.n210 VSUBS 0.013634f
C464 VDD1.n211 VSUBS 0.014436f
C465 VDD1.n212 VSUBS 0.032227f
C466 VDD1.n213 VSUBS 0.082052f
C467 VDD1.n214 VSUBS 0.014436f
C468 VDD1.n215 VSUBS 0.013634f
C469 VDD1.n216 VSUBS 0.060035f
C470 VDD1.n217 VSUBS 0.9229f
C471 VTAIL.n0 VSUBS 0.028905f
C472 VTAIL.n1 VSUBS 0.025234f
C473 VTAIL.n2 VSUBS 0.01356f
C474 VTAIL.n3 VSUBS 0.03205f
C475 VTAIL.n4 VSUBS 0.014357f
C476 VTAIL.n5 VSUBS 0.025234f
C477 VTAIL.n6 VSUBS 0.01356f
C478 VTAIL.n7 VSUBS 0.03205f
C479 VTAIL.n8 VSUBS 0.014357f
C480 VTAIL.n9 VSUBS 0.025234f
C481 VTAIL.n10 VSUBS 0.01356f
C482 VTAIL.n11 VSUBS 0.03205f
C483 VTAIL.n12 VSUBS 0.013958f
C484 VTAIL.n13 VSUBS 0.025234f
C485 VTAIL.n14 VSUBS 0.014357f
C486 VTAIL.n15 VSUBS 0.03205f
C487 VTAIL.n16 VSUBS 0.014357f
C488 VTAIL.n17 VSUBS 0.025234f
C489 VTAIL.n18 VSUBS 0.01356f
C490 VTAIL.n19 VSUBS 0.03205f
C491 VTAIL.n20 VSUBS 0.014357f
C492 VTAIL.n21 VSUBS 0.025234f
C493 VTAIL.n22 VSUBS 0.01356f
C494 VTAIL.n23 VSUBS 0.03205f
C495 VTAIL.n24 VSUBS 0.014357f
C496 VTAIL.n25 VSUBS 0.025234f
C497 VTAIL.n26 VSUBS 0.01356f
C498 VTAIL.n27 VSUBS 0.03205f
C499 VTAIL.n28 VSUBS 0.014357f
C500 VTAIL.n29 VSUBS 0.025234f
C501 VTAIL.n30 VSUBS 0.01356f
C502 VTAIL.n31 VSUBS 0.03205f
C503 VTAIL.n32 VSUBS 0.014357f
C504 VTAIL.n33 VSUBS 2.15194f
C505 VTAIL.n34 VSUBS 0.01356f
C506 VTAIL.t3 VSUBS 0.068909f
C507 VTAIL.n35 VSUBS 0.213009f
C508 VTAIL.n36 VSUBS 0.020389f
C509 VTAIL.n37 VSUBS 0.024038f
C510 VTAIL.n38 VSUBS 0.03205f
C511 VTAIL.n39 VSUBS 0.014357f
C512 VTAIL.n40 VSUBS 0.01356f
C513 VTAIL.n41 VSUBS 0.025234f
C514 VTAIL.n42 VSUBS 0.025234f
C515 VTAIL.n43 VSUBS 0.01356f
C516 VTAIL.n44 VSUBS 0.014357f
C517 VTAIL.n45 VSUBS 0.03205f
C518 VTAIL.n46 VSUBS 0.03205f
C519 VTAIL.n47 VSUBS 0.014357f
C520 VTAIL.n48 VSUBS 0.01356f
C521 VTAIL.n49 VSUBS 0.025234f
C522 VTAIL.n50 VSUBS 0.025234f
C523 VTAIL.n51 VSUBS 0.01356f
C524 VTAIL.n52 VSUBS 0.014357f
C525 VTAIL.n53 VSUBS 0.03205f
C526 VTAIL.n54 VSUBS 0.03205f
C527 VTAIL.n55 VSUBS 0.014357f
C528 VTAIL.n56 VSUBS 0.01356f
C529 VTAIL.n57 VSUBS 0.025234f
C530 VTAIL.n58 VSUBS 0.025234f
C531 VTAIL.n59 VSUBS 0.01356f
C532 VTAIL.n60 VSUBS 0.014357f
C533 VTAIL.n61 VSUBS 0.03205f
C534 VTAIL.n62 VSUBS 0.03205f
C535 VTAIL.n63 VSUBS 0.014357f
C536 VTAIL.n64 VSUBS 0.01356f
C537 VTAIL.n65 VSUBS 0.025234f
C538 VTAIL.n66 VSUBS 0.025234f
C539 VTAIL.n67 VSUBS 0.01356f
C540 VTAIL.n68 VSUBS 0.014357f
C541 VTAIL.n69 VSUBS 0.03205f
C542 VTAIL.n70 VSUBS 0.03205f
C543 VTAIL.n71 VSUBS 0.014357f
C544 VTAIL.n72 VSUBS 0.01356f
C545 VTAIL.n73 VSUBS 0.025234f
C546 VTAIL.n74 VSUBS 0.025234f
C547 VTAIL.n75 VSUBS 0.01356f
C548 VTAIL.n76 VSUBS 0.01356f
C549 VTAIL.n77 VSUBS 0.014357f
C550 VTAIL.n78 VSUBS 0.03205f
C551 VTAIL.n79 VSUBS 0.03205f
C552 VTAIL.n80 VSUBS 0.03205f
C553 VTAIL.n81 VSUBS 0.013958f
C554 VTAIL.n82 VSUBS 0.01356f
C555 VTAIL.n83 VSUBS 0.025234f
C556 VTAIL.n84 VSUBS 0.025234f
C557 VTAIL.n85 VSUBS 0.01356f
C558 VTAIL.n86 VSUBS 0.014357f
C559 VTAIL.n87 VSUBS 0.03205f
C560 VTAIL.n88 VSUBS 0.03205f
C561 VTAIL.n89 VSUBS 0.014357f
C562 VTAIL.n90 VSUBS 0.01356f
C563 VTAIL.n91 VSUBS 0.025234f
C564 VTAIL.n92 VSUBS 0.025234f
C565 VTAIL.n93 VSUBS 0.01356f
C566 VTAIL.n94 VSUBS 0.014357f
C567 VTAIL.n95 VSUBS 0.03205f
C568 VTAIL.n96 VSUBS 0.03205f
C569 VTAIL.n97 VSUBS 0.014357f
C570 VTAIL.n98 VSUBS 0.01356f
C571 VTAIL.n99 VSUBS 0.025234f
C572 VTAIL.n100 VSUBS 0.025234f
C573 VTAIL.n101 VSUBS 0.01356f
C574 VTAIL.n102 VSUBS 0.014357f
C575 VTAIL.n103 VSUBS 0.03205f
C576 VTAIL.n104 VSUBS 0.081603f
C577 VTAIL.n105 VSUBS 0.014357f
C578 VTAIL.n106 VSUBS 0.01356f
C579 VTAIL.n107 VSUBS 0.059706f
C580 VTAIL.n108 VSUBS 0.041257f
C581 VTAIL.n109 VSUBS 1.9226f
C582 VTAIL.n110 VSUBS 0.028905f
C583 VTAIL.n111 VSUBS 0.025234f
C584 VTAIL.n112 VSUBS 0.01356f
C585 VTAIL.n113 VSUBS 0.03205f
C586 VTAIL.n114 VSUBS 0.014357f
C587 VTAIL.n115 VSUBS 0.025234f
C588 VTAIL.n116 VSUBS 0.01356f
C589 VTAIL.n117 VSUBS 0.03205f
C590 VTAIL.n118 VSUBS 0.014357f
C591 VTAIL.n119 VSUBS 0.025234f
C592 VTAIL.n120 VSUBS 0.01356f
C593 VTAIL.n121 VSUBS 0.03205f
C594 VTAIL.n122 VSUBS 0.013958f
C595 VTAIL.n123 VSUBS 0.025234f
C596 VTAIL.n124 VSUBS 0.013958f
C597 VTAIL.n125 VSUBS 0.01356f
C598 VTAIL.n126 VSUBS 0.03205f
C599 VTAIL.n127 VSUBS 0.03205f
C600 VTAIL.n128 VSUBS 0.014357f
C601 VTAIL.n129 VSUBS 0.025234f
C602 VTAIL.n130 VSUBS 0.01356f
C603 VTAIL.n131 VSUBS 0.03205f
C604 VTAIL.n132 VSUBS 0.014357f
C605 VTAIL.n133 VSUBS 0.025234f
C606 VTAIL.n134 VSUBS 0.01356f
C607 VTAIL.n135 VSUBS 0.03205f
C608 VTAIL.n136 VSUBS 0.014357f
C609 VTAIL.n137 VSUBS 0.025234f
C610 VTAIL.n138 VSUBS 0.01356f
C611 VTAIL.n139 VSUBS 0.03205f
C612 VTAIL.n140 VSUBS 0.014357f
C613 VTAIL.n141 VSUBS 0.025234f
C614 VTAIL.n142 VSUBS 0.01356f
C615 VTAIL.n143 VSUBS 0.03205f
C616 VTAIL.n144 VSUBS 0.014357f
C617 VTAIL.n145 VSUBS 2.15194f
C618 VTAIL.n146 VSUBS 0.01356f
C619 VTAIL.t0 VSUBS 0.068909f
C620 VTAIL.n147 VSUBS 0.213009f
C621 VTAIL.n148 VSUBS 0.020389f
C622 VTAIL.n149 VSUBS 0.024038f
C623 VTAIL.n150 VSUBS 0.03205f
C624 VTAIL.n151 VSUBS 0.014357f
C625 VTAIL.n152 VSUBS 0.01356f
C626 VTAIL.n153 VSUBS 0.025234f
C627 VTAIL.n154 VSUBS 0.025234f
C628 VTAIL.n155 VSUBS 0.01356f
C629 VTAIL.n156 VSUBS 0.014357f
C630 VTAIL.n157 VSUBS 0.03205f
C631 VTAIL.n158 VSUBS 0.03205f
C632 VTAIL.n159 VSUBS 0.014357f
C633 VTAIL.n160 VSUBS 0.01356f
C634 VTAIL.n161 VSUBS 0.025234f
C635 VTAIL.n162 VSUBS 0.025234f
C636 VTAIL.n163 VSUBS 0.01356f
C637 VTAIL.n164 VSUBS 0.014357f
C638 VTAIL.n165 VSUBS 0.03205f
C639 VTAIL.n166 VSUBS 0.03205f
C640 VTAIL.n167 VSUBS 0.014357f
C641 VTAIL.n168 VSUBS 0.01356f
C642 VTAIL.n169 VSUBS 0.025234f
C643 VTAIL.n170 VSUBS 0.025234f
C644 VTAIL.n171 VSUBS 0.01356f
C645 VTAIL.n172 VSUBS 0.014357f
C646 VTAIL.n173 VSUBS 0.03205f
C647 VTAIL.n174 VSUBS 0.03205f
C648 VTAIL.n175 VSUBS 0.014357f
C649 VTAIL.n176 VSUBS 0.01356f
C650 VTAIL.n177 VSUBS 0.025234f
C651 VTAIL.n178 VSUBS 0.025234f
C652 VTAIL.n179 VSUBS 0.01356f
C653 VTAIL.n180 VSUBS 0.014357f
C654 VTAIL.n181 VSUBS 0.03205f
C655 VTAIL.n182 VSUBS 0.03205f
C656 VTAIL.n183 VSUBS 0.014357f
C657 VTAIL.n184 VSUBS 0.01356f
C658 VTAIL.n185 VSUBS 0.025234f
C659 VTAIL.n186 VSUBS 0.025234f
C660 VTAIL.n187 VSUBS 0.01356f
C661 VTAIL.n188 VSUBS 0.014357f
C662 VTAIL.n189 VSUBS 0.03205f
C663 VTAIL.n190 VSUBS 0.03205f
C664 VTAIL.n191 VSUBS 0.014357f
C665 VTAIL.n192 VSUBS 0.01356f
C666 VTAIL.n193 VSUBS 0.025234f
C667 VTAIL.n194 VSUBS 0.025234f
C668 VTAIL.n195 VSUBS 0.01356f
C669 VTAIL.n196 VSUBS 0.014357f
C670 VTAIL.n197 VSUBS 0.03205f
C671 VTAIL.n198 VSUBS 0.03205f
C672 VTAIL.n199 VSUBS 0.014357f
C673 VTAIL.n200 VSUBS 0.01356f
C674 VTAIL.n201 VSUBS 0.025234f
C675 VTAIL.n202 VSUBS 0.025234f
C676 VTAIL.n203 VSUBS 0.01356f
C677 VTAIL.n204 VSUBS 0.014357f
C678 VTAIL.n205 VSUBS 0.03205f
C679 VTAIL.n206 VSUBS 0.03205f
C680 VTAIL.n207 VSUBS 0.014357f
C681 VTAIL.n208 VSUBS 0.01356f
C682 VTAIL.n209 VSUBS 0.025234f
C683 VTAIL.n210 VSUBS 0.025234f
C684 VTAIL.n211 VSUBS 0.01356f
C685 VTAIL.n212 VSUBS 0.014357f
C686 VTAIL.n213 VSUBS 0.03205f
C687 VTAIL.n214 VSUBS 0.081603f
C688 VTAIL.n215 VSUBS 0.014357f
C689 VTAIL.n216 VSUBS 0.01356f
C690 VTAIL.n217 VSUBS 0.059706f
C691 VTAIL.n218 VSUBS 0.041257f
C692 VTAIL.n219 VSUBS 1.93242f
C693 VTAIL.n220 VSUBS 0.028905f
C694 VTAIL.n221 VSUBS 0.025234f
C695 VTAIL.n222 VSUBS 0.01356f
C696 VTAIL.n223 VSUBS 0.03205f
C697 VTAIL.n224 VSUBS 0.014357f
C698 VTAIL.n225 VSUBS 0.025234f
C699 VTAIL.n226 VSUBS 0.01356f
C700 VTAIL.n227 VSUBS 0.03205f
C701 VTAIL.n228 VSUBS 0.014357f
C702 VTAIL.n229 VSUBS 0.025234f
C703 VTAIL.n230 VSUBS 0.01356f
C704 VTAIL.n231 VSUBS 0.03205f
C705 VTAIL.n232 VSUBS 0.013958f
C706 VTAIL.n233 VSUBS 0.025234f
C707 VTAIL.n234 VSUBS 0.013958f
C708 VTAIL.n235 VSUBS 0.01356f
C709 VTAIL.n236 VSUBS 0.03205f
C710 VTAIL.n237 VSUBS 0.03205f
C711 VTAIL.n238 VSUBS 0.014357f
C712 VTAIL.n239 VSUBS 0.025234f
C713 VTAIL.n240 VSUBS 0.01356f
C714 VTAIL.n241 VSUBS 0.03205f
C715 VTAIL.n242 VSUBS 0.014357f
C716 VTAIL.n243 VSUBS 0.025234f
C717 VTAIL.n244 VSUBS 0.01356f
C718 VTAIL.n245 VSUBS 0.03205f
C719 VTAIL.n246 VSUBS 0.014357f
C720 VTAIL.n247 VSUBS 0.025234f
C721 VTAIL.n248 VSUBS 0.01356f
C722 VTAIL.n249 VSUBS 0.03205f
C723 VTAIL.n250 VSUBS 0.014357f
C724 VTAIL.n251 VSUBS 0.025234f
C725 VTAIL.n252 VSUBS 0.01356f
C726 VTAIL.n253 VSUBS 0.03205f
C727 VTAIL.n254 VSUBS 0.014357f
C728 VTAIL.n255 VSUBS 2.15194f
C729 VTAIL.n256 VSUBS 0.01356f
C730 VTAIL.t2 VSUBS 0.068909f
C731 VTAIL.n257 VSUBS 0.213009f
C732 VTAIL.n258 VSUBS 0.020389f
C733 VTAIL.n259 VSUBS 0.024038f
C734 VTAIL.n260 VSUBS 0.03205f
C735 VTAIL.n261 VSUBS 0.014357f
C736 VTAIL.n262 VSUBS 0.01356f
C737 VTAIL.n263 VSUBS 0.025234f
C738 VTAIL.n264 VSUBS 0.025234f
C739 VTAIL.n265 VSUBS 0.01356f
C740 VTAIL.n266 VSUBS 0.014357f
C741 VTAIL.n267 VSUBS 0.03205f
C742 VTAIL.n268 VSUBS 0.03205f
C743 VTAIL.n269 VSUBS 0.014357f
C744 VTAIL.n270 VSUBS 0.01356f
C745 VTAIL.n271 VSUBS 0.025234f
C746 VTAIL.n272 VSUBS 0.025234f
C747 VTAIL.n273 VSUBS 0.01356f
C748 VTAIL.n274 VSUBS 0.014357f
C749 VTAIL.n275 VSUBS 0.03205f
C750 VTAIL.n276 VSUBS 0.03205f
C751 VTAIL.n277 VSUBS 0.014357f
C752 VTAIL.n278 VSUBS 0.01356f
C753 VTAIL.n279 VSUBS 0.025234f
C754 VTAIL.n280 VSUBS 0.025234f
C755 VTAIL.n281 VSUBS 0.01356f
C756 VTAIL.n282 VSUBS 0.014357f
C757 VTAIL.n283 VSUBS 0.03205f
C758 VTAIL.n284 VSUBS 0.03205f
C759 VTAIL.n285 VSUBS 0.014357f
C760 VTAIL.n286 VSUBS 0.01356f
C761 VTAIL.n287 VSUBS 0.025234f
C762 VTAIL.n288 VSUBS 0.025234f
C763 VTAIL.n289 VSUBS 0.01356f
C764 VTAIL.n290 VSUBS 0.014357f
C765 VTAIL.n291 VSUBS 0.03205f
C766 VTAIL.n292 VSUBS 0.03205f
C767 VTAIL.n293 VSUBS 0.014357f
C768 VTAIL.n294 VSUBS 0.01356f
C769 VTAIL.n295 VSUBS 0.025234f
C770 VTAIL.n296 VSUBS 0.025234f
C771 VTAIL.n297 VSUBS 0.01356f
C772 VTAIL.n298 VSUBS 0.014357f
C773 VTAIL.n299 VSUBS 0.03205f
C774 VTAIL.n300 VSUBS 0.03205f
C775 VTAIL.n301 VSUBS 0.014357f
C776 VTAIL.n302 VSUBS 0.01356f
C777 VTAIL.n303 VSUBS 0.025234f
C778 VTAIL.n304 VSUBS 0.025234f
C779 VTAIL.n305 VSUBS 0.01356f
C780 VTAIL.n306 VSUBS 0.014357f
C781 VTAIL.n307 VSUBS 0.03205f
C782 VTAIL.n308 VSUBS 0.03205f
C783 VTAIL.n309 VSUBS 0.014357f
C784 VTAIL.n310 VSUBS 0.01356f
C785 VTAIL.n311 VSUBS 0.025234f
C786 VTAIL.n312 VSUBS 0.025234f
C787 VTAIL.n313 VSUBS 0.01356f
C788 VTAIL.n314 VSUBS 0.014357f
C789 VTAIL.n315 VSUBS 0.03205f
C790 VTAIL.n316 VSUBS 0.03205f
C791 VTAIL.n317 VSUBS 0.014357f
C792 VTAIL.n318 VSUBS 0.01356f
C793 VTAIL.n319 VSUBS 0.025234f
C794 VTAIL.n320 VSUBS 0.025234f
C795 VTAIL.n321 VSUBS 0.01356f
C796 VTAIL.n322 VSUBS 0.014357f
C797 VTAIL.n323 VSUBS 0.03205f
C798 VTAIL.n324 VSUBS 0.081603f
C799 VTAIL.n325 VSUBS 0.014357f
C800 VTAIL.n326 VSUBS 0.01356f
C801 VTAIL.n327 VSUBS 0.059706f
C802 VTAIL.n328 VSUBS 0.041257f
C803 VTAIL.n329 VSUBS 1.87424f
C804 VTAIL.n330 VSUBS 0.028905f
C805 VTAIL.n331 VSUBS 0.025234f
C806 VTAIL.n332 VSUBS 0.01356f
C807 VTAIL.n333 VSUBS 0.03205f
C808 VTAIL.n334 VSUBS 0.014357f
C809 VTAIL.n335 VSUBS 0.025234f
C810 VTAIL.n336 VSUBS 0.01356f
C811 VTAIL.n337 VSUBS 0.03205f
C812 VTAIL.n338 VSUBS 0.014357f
C813 VTAIL.n339 VSUBS 0.025234f
C814 VTAIL.n340 VSUBS 0.01356f
C815 VTAIL.n341 VSUBS 0.03205f
C816 VTAIL.n342 VSUBS 0.013958f
C817 VTAIL.n343 VSUBS 0.025234f
C818 VTAIL.n344 VSUBS 0.014357f
C819 VTAIL.n345 VSUBS 0.03205f
C820 VTAIL.n346 VSUBS 0.014357f
C821 VTAIL.n347 VSUBS 0.025234f
C822 VTAIL.n348 VSUBS 0.01356f
C823 VTAIL.n349 VSUBS 0.03205f
C824 VTAIL.n350 VSUBS 0.014357f
C825 VTAIL.n351 VSUBS 0.025234f
C826 VTAIL.n352 VSUBS 0.01356f
C827 VTAIL.n353 VSUBS 0.03205f
C828 VTAIL.n354 VSUBS 0.014357f
C829 VTAIL.n355 VSUBS 0.025234f
C830 VTAIL.n356 VSUBS 0.01356f
C831 VTAIL.n357 VSUBS 0.03205f
C832 VTAIL.n358 VSUBS 0.014357f
C833 VTAIL.n359 VSUBS 0.025234f
C834 VTAIL.n360 VSUBS 0.01356f
C835 VTAIL.n361 VSUBS 0.03205f
C836 VTAIL.n362 VSUBS 0.014357f
C837 VTAIL.n363 VSUBS 2.15194f
C838 VTAIL.n364 VSUBS 0.01356f
C839 VTAIL.t1 VSUBS 0.068909f
C840 VTAIL.n365 VSUBS 0.213009f
C841 VTAIL.n366 VSUBS 0.020389f
C842 VTAIL.n367 VSUBS 0.024038f
C843 VTAIL.n368 VSUBS 0.03205f
C844 VTAIL.n369 VSUBS 0.014357f
C845 VTAIL.n370 VSUBS 0.01356f
C846 VTAIL.n371 VSUBS 0.025234f
C847 VTAIL.n372 VSUBS 0.025234f
C848 VTAIL.n373 VSUBS 0.01356f
C849 VTAIL.n374 VSUBS 0.014357f
C850 VTAIL.n375 VSUBS 0.03205f
C851 VTAIL.n376 VSUBS 0.03205f
C852 VTAIL.n377 VSUBS 0.014357f
C853 VTAIL.n378 VSUBS 0.01356f
C854 VTAIL.n379 VSUBS 0.025234f
C855 VTAIL.n380 VSUBS 0.025234f
C856 VTAIL.n381 VSUBS 0.01356f
C857 VTAIL.n382 VSUBS 0.014357f
C858 VTAIL.n383 VSUBS 0.03205f
C859 VTAIL.n384 VSUBS 0.03205f
C860 VTAIL.n385 VSUBS 0.014357f
C861 VTAIL.n386 VSUBS 0.01356f
C862 VTAIL.n387 VSUBS 0.025234f
C863 VTAIL.n388 VSUBS 0.025234f
C864 VTAIL.n389 VSUBS 0.01356f
C865 VTAIL.n390 VSUBS 0.014357f
C866 VTAIL.n391 VSUBS 0.03205f
C867 VTAIL.n392 VSUBS 0.03205f
C868 VTAIL.n393 VSUBS 0.014357f
C869 VTAIL.n394 VSUBS 0.01356f
C870 VTAIL.n395 VSUBS 0.025234f
C871 VTAIL.n396 VSUBS 0.025234f
C872 VTAIL.n397 VSUBS 0.01356f
C873 VTAIL.n398 VSUBS 0.014357f
C874 VTAIL.n399 VSUBS 0.03205f
C875 VTAIL.n400 VSUBS 0.03205f
C876 VTAIL.n401 VSUBS 0.014357f
C877 VTAIL.n402 VSUBS 0.01356f
C878 VTAIL.n403 VSUBS 0.025234f
C879 VTAIL.n404 VSUBS 0.025234f
C880 VTAIL.n405 VSUBS 0.01356f
C881 VTAIL.n406 VSUBS 0.01356f
C882 VTAIL.n407 VSUBS 0.014357f
C883 VTAIL.n408 VSUBS 0.03205f
C884 VTAIL.n409 VSUBS 0.03205f
C885 VTAIL.n410 VSUBS 0.03205f
C886 VTAIL.n411 VSUBS 0.013958f
C887 VTAIL.n412 VSUBS 0.01356f
C888 VTAIL.n413 VSUBS 0.025234f
C889 VTAIL.n414 VSUBS 0.025234f
C890 VTAIL.n415 VSUBS 0.01356f
C891 VTAIL.n416 VSUBS 0.014357f
C892 VTAIL.n417 VSUBS 0.03205f
C893 VTAIL.n418 VSUBS 0.03205f
C894 VTAIL.n419 VSUBS 0.014357f
C895 VTAIL.n420 VSUBS 0.01356f
C896 VTAIL.n421 VSUBS 0.025234f
C897 VTAIL.n422 VSUBS 0.025234f
C898 VTAIL.n423 VSUBS 0.01356f
C899 VTAIL.n424 VSUBS 0.014357f
C900 VTAIL.n425 VSUBS 0.03205f
C901 VTAIL.n426 VSUBS 0.03205f
C902 VTAIL.n427 VSUBS 0.014357f
C903 VTAIL.n428 VSUBS 0.01356f
C904 VTAIL.n429 VSUBS 0.025234f
C905 VTAIL.n430 VSUBS 0.025234f
C906 VTAIL.n431 VSUBS 0.01356f
C907 VTAIL.n432 VSUBS 0.014357f
C908 VTAIL.n433 VSUBS 0.03205f
C909 VTAIL.n434 VSUBS 0.081603f
C910 VTAIL.n435 VSUBS 0.014357f
C911 VTAIL.n436 VSUBS 0.01356f
C912 VTAIL.n437 VSUBS 0.059706f
C913 VTAIL.n438 VSUBS 0.041257f
C914 VTAIL.n439 VSUBS 1.81676f
C915 VP.t0 VSUBS 1.60802f
C916 VP.t1 VSUBS 1.50526f
C917 VP.n0 VSUBS 5.57517f
C918 B.n0 VSUBS 0.004427f
C919 B.n1 VSUBS 0.004427f
C920 B.n2 VSUBS 0.007001f
C921 B.n3 VSUBS 0.007001f
C922 B.n4 VSUBS 0.007001f
C923 B.n5 VSUBS 0.007001f
C924 B.n6 VSUBS 0.007001f
C925 B.n7 VSUBS 0.007001f
C926 B.n8 VSUBS 0.016625f
C927 B.n9 VSUBS 0.007001f
C928 B.n10 VSUBS 0.007001f
C929 B.n11 VSUBS 0.007001f
C930 B.n12 VSUBS 0.007001f
C931 B.n13 VSUBS 0.007001f
C932 B.n14 VSUBS 0.007001f
C933 B.n15 VSUBS 0.007001f
C934 B.n16 VSUBS 0.007001f
C935 B.n17 VSUBS 0.007001f
C936 B.n18 VSUBS 0.007001f
C937 B.n19 VSUBS 0.007001f
C938 B.n20 VSUBS 0.007001f
C939 B.n21 VSUBS 0.007001f
C940 B.n22 VSUBS 0.007001f
C941 B.n23 VSUBS 0.007001f
C942 B.n24 VSUBS 0.007001f
C943 B.n25 VSUBS 0.007001f
C944 B.n26 VSUBS 0.007001f
C945 B.n27 VSUBS 0.007001f
C946 B.n28 VSUBS 0.007001f
C947 B.n29 VSUBS 0.007001f
C948 B.n30 VSUBS 0.007001f
C949 B.n31 VSUBS 0.007001f
C950 B.n32 VSUBS 0.007001f
C951 B.n33 VSUBS 0.007001f
C952 B.n34 VSUBS 0.007001f
C953 B.n35 VSUBS 0.007001f
C954 B.n36 VSUBS 0.007001f
C955 B.n37 VSUBS 0.007001f
C956 B.n38 VSUBS 0.007001f
C957 B.n39 VSUBS 0.007001f
C958 B.n40 VSUBS 0.006384f
C959 B.n41 VSUBS 0.007001f
C960 B.t11 VSUBS 0.393292f
C961 B.t10 VSUBS 0.403299f
C962 B.t9 VSUBS 0.389021f
C963 B.n42 VSUBS 0.438662f
C964 B.n43 VSUBS 0.340118f
C965 B.n44 VSUBS 0.016221f
C966 B.n45 VSUBS 0.007001f
C967 B.n46 VSUBS 0.007001f
C968 B.n47 VSUBS 0.007001f
C969 B.n48 VSUBS 0.007001f
C970 B.t5 VSUBS 0.393295f
C971 B.t4 VSUBS 0.403303f
C972 B.t3 VSUBS 0.389021f
C973 B.n49 VSUBS 0.438658f
C974 B.n50 VSUBS 0.340115f
C975 B.n51 VSUBS 0.007001f
C976 B.n52 VSUBS 0.007001f
C977 B.n53 VSUBS 0.007001f
C978 B.n54 VSUBS 0.007001f
C979 B.n55 VSUBS 0.007001f
C980 B.n56 VSUBS 0.007001f
C981 B.n57 VSUBS 0.007001f
C982 B.n58 VSUBS 0.007001f
C983 B.n59 VSUBS 0.007001f
C984 B.n60 VSUBS 0.007001f
C985 B.n61 VSUBS 0.007001f
C986 B.n62 VSUBS 0.007001f
C987 B.n63 VSUBS 0.007001f
C988 B.n64 VSUBS 0.007001f
C989 B.n65 VSUBS 0.007001f
C990 B.n66 VSUBS 0.007001f
C991 B.n67 VSUBS 0.007001f
C992 B.n68 VSUBS 0.007001f
C993 B.n69 VSUBS 0.007001f
C994 B.n70 VSUBS 0.007001f
C995 B.n71 VSUBS 0.007001f
C996 B.n72 VSUBS 0.007001f
C997 B.n73 VSUBS 0.007001f
C998 B.n74 VSUBS 0.007001f
C999 B.n75 VSUBS 0.007001f
C1000 B.n76 VSUBS 0.007001f
C1001 B.n77 VSUBS 0.007001f
C1002 B.n78 VSUBS 0.007001f
C1003 B.n79 VSUBS 0.007001f
C1004 B.n80 VSUBS 0.007001f
C1005 B.n81 VSUBS 0.007001f
C1006 B.n82 VSUBS 0.017146f
C1007 B.n83 VSUBS 0.007001f
C1008 B.n84 VSUBS 0.007001f
C1009 B.n85 VSUBS 0.007001f
C1010 B.n86 VSUBS 0.007001f
C1011 B.n87 VSUBS 0.007001f
C1012 B.n88 VSUBS 0.007001f
C1013 B.n89 VSUBS 0.007001f
C1014 B.n90 VSUBS 0.007001f
C1015 B.n91 VSUBS 0.007001f
C1016 B.n92 VSUBS 0.007001f
C1017 B.n93 VSUBS 0.007001f
C1018 B.n94 VSUBS 0.007001f
C1019 B.n95 VSUBS 0.007001f
C1020 B.n96 VSUBS 0.017146f
C1021 B.n97 VSUBS 0.007001f
C1022 B.n98 VSUBS 0.007001f
C1023 B.n99 VSUBS 0.007001f
C1024 B.n100 VSUBS 0.007001f
C1025 B.n101 VSUBS 0.007001f
C1026 B.n102 VSUBS 0.007001f
C1027 B.n103 VSUBS 0.007001f
C1028 B.n104 VSUBS 0.007001f
C1029 B.n105 VSUBS 0.007001f
C1030 B.n106 VSUBS 0.007001f
C1031 B.n107 VSUBS 0.007001f
C1032 B.n108 VSUBS 0.007001f
C1033 B.n109 VSUBS 0.007001f
C1034 B.n110 VSUBS 0.007001f
C1035 B.n111 VSUBS 0.007001f
C1036 B.n112 VSUBS 0.007001f
C1037 B.n113 VSUBS 0.007001f
C1038 B.n114 VSUBS 0.007001f
C1039 B.n115 VSUBS 0.007001f
C1040 B.n116 VSUBS 0.007001f
C1041 B.n117 VSUBS 0.007001f
C1042 B.n118 VSUBS 0.007001f
C1043 B.n119 VSUBS 0.007001f
C1044 B.n120 VSUBS 0.007001f
C1045 B.n121 VSUBS 0.007001f
C1046 B.n122 VSUBS 0.007001f
C1047 B.n123 VSUBS 0.007001f
C1048 B.n124 VSUBS 0.007001f
C1049 B.n125 VSUBS 0.007001f
C1050 B.n126 VSUBS 0.007001f
C1051 B.n127 VSUBS 0.007001f
C1052 B.n128 VSUBS 0.007001f
C1053 B.t7 VSUBS 0.393295f
C1054 B.t8 VSUBS 0.403303f
C1055 B.t6 VSUBS 0.389021f
C1056 B.n129 VSUBS 0.438658f
C1057 B.n130 VSUBS 0.340115f
C1058 B.n131 VSUBS 0.007001f
C1059 B.n132 VSUBS 0.007001f
C1060 B.n133 VSUBS 0.007001f
C1061 B.n134 VSUBS 0.007001f
C1062 B.t1 VSUBS 0.393292f
C1063 B.t2 VSUBS 0.403299f
C1064 B.t0 VSUBS 0.389021f
C1065 B.n135 VSUBS 0.438662f
C1066 B.n136 VSUBS 0.340118f
C1067 B.n137 VSUBS 0.016221f
C1068 B.n138 VSUBS 0.007001f
C1069 B.n139 VSUBS 0.007001f
C1070 B.n140 VSUBS 0.007001f
C1071 B.n141 VSUBS 0.007001f
C1072 B.n142 VSUBS 0.007001f
C1073 B.n143 VSUBS 0.007001f
C1074 B.n144 VSUBS 0.007001f
C1075 B.n145 VSUBS 0.007001f
C1076 B.n146 VSUBS 0.007001f
C1077 B.n147 VSUBS 0.007001f
C1078 B.n148 VSUBS 0.007001f
C1079 B.n149 VSUBS 0.007001f
C1080 B.n150 VSUBS 0.007001f
C1081 B.n151 VSUBS 0.007001f
C1082 B.n152 VSUBS 0.007001f
C1083 B.n153 VSUBS 0.007001f
C1084 B.n154 VSUBS 0.007001f
C1085 B.n155 VSUBS 0.007001f
C1086 B.n156 VSUBS 0.007001f
C1087 B.n157 VSUBS 0.007001f
C1088 B.n158 VSUBS 0.007001f
C1089 B.n159 VSUBS 0.007001f
C1090 B.n160 VSUBS 0.007001f
C1091 B.n161 VSUBS 0.007001f
C1092 B.n162 VSUBS 0.007001f
C1093 B.n163 VSUBS 0.007001f
C1094 B.n164 VSUBS 0.007001f
C1095 B.n165 VSUBS 0.007001f
C1096 B.n166 VSUBS 0.007001f
C1097 B.n167 VSUBS 0.007001f
C1098 B.n168 VSUBS 0.007001f
C1099 B.n169 VSUBS 0.017146f
C1100 B.n170 VSUBS 0.007001f
C1101 B.n171 VSUBS 0.007001f
C1102 B.n172 VSUBS 0.007001f
C1103 B.n173 VSUBS 0.007001f
C1104 B.n174 VSUBS 0.007001f
C1105 B.n175 VSUBS 0.007001f
C1106 B.n176 VSUBS 0.007001f
C1107 B.n177 VSUBS 0.007001f
C1108 B.n178 VSUBS 0.007001f
C1109 B.n179 VSUBS 0.007001f
C1110 B.n180 VSUBS 0.007001f
C1111 B.n181 VSUBS 0.007001f
C1112 B.n182 VSUBS 0.007001f
C1113 B.n183 VSUBS 0.007001f
C1114 B.n184 VSUBS 0.007001f
C1115 B.n185 VSUBS 0.007001f
C1116 B.n186 VSUBS 0.007001f
C1117 B.n187 VSUBS 0.007001f
C1118 B.n188 VSUBS 0.007001f
C1119 B.n189 VSUBS 0.007001f
C1120 B.n190 VSUBS 0.007001f
C1121 B.n191 VSUBS 0.007001f
C1122 B.n192 VSUBS 0.016625f
C1123 B.n193 VSUBS 0.016625f
C1124 B.n194 VSUBS 0.017146f
C1125 B.n195 VSUBS 0.007001f
C1126 B.n196 VSUBS 0.007001f
C1127 B.n197 VSUBS 0.007001f
C1128 B.n198 VSUBS 0.007001f
C1129 B.n199 VSUBS 0.007001f
C1130 B.n200 VSUBS 0.007001f
C1131 B.n201 VSUBS 0.007001f
C1132 B.n202 VSUBS 0.007001f
C1133 B.n203 VSUBS 0.007001f
C1134 B.n204 VSUBS 0.007001f
C1135 B.n205 VSUBS 0.007001f
C1136 B.n206 VSUBS 0.007001f
C1137 B.n207 VSUBS 0.007001f
C1138 B.n208 VSUBS 0.007001f
C1139 B.n209 VSUBS 0.007001f
C1140 B.n210 VSUBS 0.007001f
C1141 B.n211 VSUBS 0.007001f
C1142 B.n212 VSUBS 0.007001f
C1143 B.n213 VSUBS 0.007001f
C1144 B.n214 VSUBS 0.007001f
C1145 B.n215 VSUBS 0.007001f
C1146 B.n216 VSUBS 0.007001f
C1147 B.n217 VSUBS 0.007001f
C1148 B.n218 VSUBS 0.007001f
C1149 B.n219 VSUBS 0.007001f
C1150 B.n220 VSUBS 0.007001f
C1151 B.n221 VSUBS 0.007001f
C1152 B.n222 VSUBS 0.007001f
C1153 B.n223 VSUBS 0.007001f
C1154 B.n224 VSUBS 0.007001f
C1155 B.n225 VSUBS 0.007001f
C1156 B.n226 VSUBS 0.007001f
C1157 B.n227 VSUBS 0.007001f
C1158 B.n228 VSUBS 0.007001f
C1159 B.n229 VSUBS 0.007001f
C1160 B.n230 VSUBS 0.007001f
C1161 B.n231 VSUBS 0.007001f
C1162 B.n232 VSUBS 0.007001f
C1163 B.n233 VSUBS 0.007001f
C1164 B.n234 VSUBS 0.007001f
C1165 B.n235 VSUBS 0.007001f
C1166 B.n236 VSUBS 0.007001f
C1167 B.n237 VSUBS 0.007001f
C1168 B.n238 VSUBS 0.007001f
C1169 B.n239 VSUBS 0.007001f
C1170 B.n240 VSUBS 0.007001f
C1171 B.n241 VSUBS 0.007001f
C1172 B.n242 VSUBS 0.007001f
C1173 B.n243 VSUBS 0.007001f
C1174 B.n244 VSUBS 0.007001f
C1175 B.n245 VSUBS 0.007001f
C1176 B.n246 VSUBS 0.007001f
C1177 B.n247 VSUBS 0.007001f
C1178 B.n248 VSUBS 0.007001f
C1179 B.n249 VSUBS 0.007001f
C1180 B.n250 VSUBS 0.007001f
C1181 B.n251 VSUBS 0.007001f
C1182 B.n252 VSUBS 0.007001f
C1183 B.n253 VSUBS 0.007001f
C1184 B.n254 VSUBS 0.007001f
C1185 B.n255 VSUBS 0.007001f
C1186 B.n256 VSUBS 0.007001f
C1187 B.n257 VSUBS 0.007001f
C1188 B.n258 VSUBS 0.007001f
C1189 B.n259 VSUBS 0.007001f
C1190 B.n260 VSUBS 0.007001f
C1191 B.n261 VSUBS 0.007001f
C1192 B.n262 VSUBS 0.007001f
C1193 B.n263 VSUBS 0.007001f
C1194 B.n264 VSUBS 0.007001f
C1195 B.n265 VSUBS 0.007001f
C1196 B.n266 VSUBS 0.007001f
C1197 B.n267 VSUBS 0.007001f
C1198 B.n268 VSUBS 0.007001f
C1199 B.n269 VSUBS 0.007001f
C1200 B.n270 VSUBS 0.007001f
C1201 B.n271 VSUBS 0.007001f
C1202 B.n272 VSUBS 0.007001f
C1203 B.n273 VSUBS 0.007001f
C1204 B.n274 VSUBS 0.007001f
C1205 B.n275 VSUBS 0.007001f
C1206 B.n276 VSUBS 0.007001f
C1207 B.n277 VSUBS 0.007001f
C1208 B.n278 VSUBS 0.007001f
C1209 B.n279 VSUBS 0.007001f
C1210 B.n280 VSUBS 0.007001f
C1211 B.n281 VSUBS 0.007001f
C1212 B.n282 VSUBS 0.007001f
C1213 B.n283 VSUBS 0.007001f
C1214 B.n284 VSUBS 0.007001f
C1215 B.n285 VSUBS 0.007001f
C1216 B.n286 VSUBS 0.007001f
C1217 B.n287 VSUBS 0.007001f
C1218 B.n288 VSUBS 0.006384f
C1219 B.n289 VSUBS 0.007001f
C1220 B.n290 VSUBS 0.007001f
C1221 B.n291 VSUBS 0.004118f
C1222 B.n292 VSUBS 0.007001f
C1223 B.n293 VSUBS 0.007001f
C1224 B.n294 VSUBS 0.007001f
C1225 B.n295 VSUBS 0.007001f
C1226 B.n296 VSUBS 0.007001f
C1227 B.n297 VSUBS 0.007001f
C1228 B.n298 VSUBS 0.007001f
C1229 B.n299 VSUBS 0.007001f
C1230 B.n300 VSUBS 0.007001f
C1231 B.n301 VSUBS 0.007001f
C1232 B.n302 VSUBS 0.007001f
C1233 B.n303 VSUBS 0.007001f
C1234 B.n304 VSUBS 0.004118f
C1235 B.n305 VSUBS 0.016221f
C1236 B.n306 VSUBS 0.006384f
C1237 B.n307 VSUBS 0.007001f
C1238 B.n308 VSUBS 0.007001f
C1239 B.n309 VSUBS 0.007001f
C1240 B.n310 VSUBS 0.007001f
C1241 B.n311 VSUBS 0.007001f
C1242 B.n312 VSUBS 0.007001f
C1243 B.n313 VSUBS 0.007001f
C1244 B.n314 VSUBS 0.007001f
C1245 B.n315 VSUBS 0.007001f
C1246 B.n316 VSUBS 0.007001f
C1247 B.n317 VSUBS 0.007001f
C1248 B.n318 VSUBS 0.007001f
C1249 B.n319 VSUBS 0.007001f
C1250 B.n320 VSUBS 0.007001f
C1251 B.n321 VSUBS 0.007001f
C1252 B.n322 VSUBS 0.007001f
C1253 B.n323 VSUBS 0.007001f
C1254 B.n324 VSUBS 0.007001f
C1255 B.n325 VSUBS 0.007001f
C1256 B.n326 VSUBS 0.007001f
C1257 B.n327 VSUBS 0.007001f
C1258 B.n328 VSUBS 0.007001f
C1259 B.n329 VSUBS 0.007001f
C1260 B.n330 VSUBS 0.007001f
C1261 B.n331 VSUBS 0.007001f
C1262 B.n332 VSUBS 0.007001f
C1263 B.n333 VSUBS 0.007001f
C1264 B.n334 VSUBS 0.007001f
C1265 B.n335 VSUBS 0.007001f
C1266 B.n336 VSUBS 0.007001f
C1267 B.n337 VSUBS 0.007001f
C1268 B.n338 VSUBS 0.007001f
C1269 B.n339 VSUBS 0.007001f
C1270 B.n340 VSUBS 0.007001f
C1271 B.n341 VSUBS 0.007001f
C1272 B.n342 VSUBS 0.007001f
C1273 B.n343 VSUBS 0.007001f
C1274 B.n344 VSUBS 0.007001f
C1275 B.n345 VSUBS 0.007001f
C1276 B.n346 VSUBS 0.007001f
C1277 B.n347 VSUBS 0.007001f
C1278 B.n348 VSUBS 0.007001f
C1279 B.n349 VSUBS 0.007001f
C1280 B.n350 VSUBS 0.007001f
C1281 B.n351 VSUBS 0.007001f
C1282 B.n352 VSUBS 0.007001f
C1283 B.n353 VSUBS 0.007001f
C1284 B.n354 VSUBS 0.007001f
C1285 B.n355 VSUBS 0.007001f
C1286 B.n356 VSUBS 0.007001f
C1287 B.n357 VSUBS 0.007001f
C1288 B.n358 VSUBS 0.007001f
C1289 B.n359 VSUBS 0.007001f
C1290 B.n360 VSUBS 0.007001f
C1291 B.n361 VSUBS 0.007001f
C1292 B.n362 VSUBS 0.007001f
C1293 B.n363 VSUBS 0.007001f
C1294 B.n364 VSUBS 0.007001f
C1295 B.n365 VSUBS 0.007001f
C1296 B.n366 VSUBS 0.007001f
C1297 B.n367 VSUBS 0.007001f
C1298 B.n368 VSUBS 0.007001f
C1299 B.n369 VSUBS 0.007001f
C1300 B.n370 VSUBS 0.007001f
C1301 B.n371 VSUBS 0.007001f
C1302 B.n372 VSUBS 0.007001f
C1303 B.n373 VSUBS 0.007001f
C1304 B.n374 VSUBS 0.007001f
C1305 B.n375 VSUBS 0.007001f
C1306 B.n376 VSUBS 0.007001f
C1307 B.n377 VSUBS 0.007001f
C1308 B.n378 VSUBS 0.007001f
C1309 B.n379 VSUBS 0.007001f
C1310 B.n380 VSUBS 0.007001f
C1311 B.n381 VSUBS 0.007001f
C1312 B.n382 VSUBS 0.007001f
C1313 B.n383 VSUBS 0.007001f
C1314 B.n384 VSUBS 0.007001f
C1315 B.n385 VSUBS 0.007001f
C1316 B.n386 VSUBS 0.007001f
C1317 B.n387 VSUBS 0.007001f
C1318 B.n388 VSUBS 0.007001f
C1319 B.n389 VSUBS 0.007001f
C1320 B.n390 VSUBS 0.007001f
C1321 B.n391 VSUBS 0.007001f
C1322 B.n392 VSUBS 0.007001f
C1323 B.n393 VSUBS 0.007001f
C1324 B.n394 VSUBS 0.007001f
C1325 B.n395 VSUBS 0.007001f
C1326 B.n396 VSUBS 0.007001f
C1327 B.n397 VSUBS 0.007001f
C1328 B.n398 VSUBS 0.007001f
C1329 B.n399 VSUBS 0.007001f
C1330 B.n400 VSUBS 0.007001f
C1331 B.n401 VSUBS 0.017146f
C1332 B.n402 VSUBS 0.016625f
C1333 B.n403 VSUBS 0.016625f
C1334 B.n404 VSUBS 0.007001f
C1335 B.n405 VSUBS 0.007001f
C1336 B.n406 VSUBS 0.007001f
C1337 B.n407 VSUBS 0.007001f
C1338 B.n408 VSUBS 0.007001f
C1339 B.n409 VSUBS 0.007001f
C1340 B.n410 VSUBS 0.007001f
C1341 B.n411 VSUBS 0.007001f
C1342 B.n412 VSUBS 0.007001f
C1343 B.n413 VSUBS 0.007001f
C1344 B.n414 VSUBS 0.007001f
C1345 B.n415 VSUBS 0.007001f
C1346 B.n416 VSUBS 0.007001f
C1347 B.n417 VSUBS 0.007001f
C1348 B.n418 VSUBS 0.007001f
C1349 B.n419 VSUBS 0.007001f
C1350 B.n420 VSUBS 0.007001f
C1351 B.n421 VSUBS 0.007001f
C1352 B.n422 VSUBS 0.007001f
C1353 B.n423 VSUBS 0.007001f
C1354 B.n424 VSUBS 0.007001f
C1355 B.n425 VSUBS 0.007001f
C1356 B.n426 VSUBS 0.007001f
C1357 B.n427 VSUBS 0.007001f
C1358 B.n428 VSUBS 0.007001f
C1359 B.n429 VSUBS 0.007001f
C1360 B.n430 VSUBS 0.007001f
C1361 B.n431 VSUBS 0.007001f
C1362 B.n432 VSUBS 0.007001f
C1363 B.n433 VSUBS 0.007001f
C1364 B.n434 VSUBS 0.007001f
C1365 B.n435 VSUBS 0.007001f
C1366 B.n436 VSUBS 0.007001f
C1367 B.n437 VSUBS 0.007001f
C1368 B.n438 VSUBS 0.007001f
C1369 B.n439 VSUBS 0.007001f
C1370 B.n440 VSUBS 0.007001f
C1371 B.n441 VSUBS 0.016625f
C1372 B.n442 VSUBS 0.017416f
C1373 B.n443 VSUBS 0.016355f
C1374 B.n444 VSUBS 0.007001f
C1375 B.n445 VSUBS 0.007001f
C1376 B.n446 VSUBS 0.007001f
C1377 B.n447 VSUBS 0.007001f
C1378 B.n448 VSUBS 0.007001f
C1379 B.n449 VSUBS 0.007001f
C1380 B.n450 VSUBS 0.007001f
C1381 B.n451 VSUBS 0.007001f
C1382 B.n452 VSUBS 0.007001f
C1383 B.n453 VSUBS 0.007001f
C1384 B.n454 VSUBS 0.007001f
C1385 B.n455 VSUBS 0.007001f
C1386 B.n456 VSUBS 0.007001f
C1387 B.n457 VSUBS 0.007001f
C1388 B.n458 VSUBS 0.007001f
C1389 B.n459 VSUBS 0.007001f
C1390 B.n460 VSUBS 0.007001f
C1391 B.n461 VSUBS 0.007001f
C1392 B.n462 VSUBS 0.007001f
C1393 B.n463 VSUBS 0.007001f
C1394 B.n464 VSUBS 0.007001f
C1395 B.n465 VSUBS 0.007001f
C1396 B.n466 VSUBS 0.007001f
C1397 B.n467 VSUBS 0.007001f
C1398 B.n468 VSUBS 0.007001f
C1399 B.n469 VSUBS 0.007001f
C1400 B.n470 VSUBS 0.007001f
C1401 B.n471 VSUBS 0.007001f
C1402 B.n472 VSUBS 0.007001f
C1403 B.n473 VSUBS 0.007001f
C1404 B.n474 VSUBS 0.007001f
C1405 B.n475 VSUBS 0.007001f
C1406 B.n476 VSUBS 0.007001f
C1407 B.n477 VSUBS 0.007001f
C1408 B.n478 VSUBS 0.007001f
C1409 B.n479 VSUBS 0.007001f
C1410 B.n480 VSUBS 0.007001f
C1411 B.n481 VSUBS 0.007001f
C1412 B.n482 VSUBS 0.007001f
C1413 B.n483 VSUBS 0.007001f
C1414 B.n484 VSUBS 0.007001f
C1415 B.n485 VSUBS 0.007001f
C1416 B.n486 VSUBS 0.007001f
C1417 B.n487 VSUBS 0.007001f
C1418 B.n488 VSUBS 0.007001f
C1419 B.n489 VSUBS 0.007001f
C1420 B.n490 VSUBS 0.007001f
C1421 B.n491 VSUBS 0.007001f
C1422 B.n492 VSUBS 0.007001f
C1423 B.n493 VSUBS 0.007001f
C1424 B.n494 VSUBS 0.007001f
C1425 B.n495 VSUBS 0.007001f
C1426 B.n496 VSUBS 0.007001f
C1427 B.n497 VSUBS 0.007001f
C1428 B.n498 VSUBS 0.007001f
C1429 B.n499 VSUBS 0.007001f
C1430 B.n500 VSUBS 0.007001f
C1431 B.n501 VSUBS 0.007001f
C1432 B.n502 VSUBS 0.007001f
C1433 B.n503 VSUBS 0.007001f
C1434 B.n504 VSUBS 0.007001f
C1435 B.n505 VSUBS 0.007001f
C1436 B.n506 VSUBS 0.007001f
C1437 B.n507 VSUBS 0.007001f
C1438 B.n508 VSUBS 0.007001f
C1439 B.n509 VSUBS 0.007001f
C1440 B.n510 VSUBS 0.007001f
C1441 B.n511 VSUBS 0.007001f
C1442 B.n512 VSUBS 0.007001f
C1443 B.n513 VSUBS 0.007001f
C1444 B.n514 VSUBS 0.007001f
C1445 B.n515 VSUBS 0.007001f
C1446 B.n516 VSUBS 0.007001f
C1447 B.n517 VSUBS 0.007001f
C1448 B.n518 VSUBS 0.007001f
C1449 B.n519 VSUBS 0.007001f
C1450 B.n520 VSUBS 0.007001f
C1451 B.n521 VSUBS 0.007001f
C1452 B.n522 VSUBS 0.007001f
C1453 B.n523 VSUBS 0.007001f
C1454 B.n524 VSUBS 0.007001f
C1455 B.n525 VSUBS 0.007001f
C1456 B.n526 VSUBS 0.007001f
C1457 B.n527 VSUBS 0.007001f
C1458 B.n528 VSUBS 0.007001f
C1459 B.n529 VSUBS 0.007001f
C1460 B.n530 VSUBS 0.007001f
C1461 B.n531 VSUBS 0.007001f
C1462 B.n532 VSUBS 0.007001f
C1463 B.n533 VSUBS 0.007001f
C1464 B.n534 VSUBS 0.007001f
C1465 B.n535 VSUBS 0.007001f
C1466 B.n536 VSUBS 0.007001f
C1467 B.n537 VSUBS 0.007001f
C1468 B.n538 VSUBS 0.006384f
C1469 B.n539 VSUBS 0.016221f
C1470 B.n540 VSUBS 0.004118f
C1471 B.n541 VSUBS 0.007001f
C1472 B.n542 VSUBS 0.007001f
C1473 B.n543 VSUBS 0.007001f
C1474 B.n544 VSUBS 0.007001f
C1475 B.n545 VSUBS 0.007001f
C1476 B.n546 VSUBS 0.007001f
C1477 B.n547 VSUBS 0.007001f
C1478 B.n548 VSUBS 0.007001f
C1479 B.n549 VSUBS 0.007001f
C1480 B.n550 VSUBS 0.007001f
C1481 B.n551 VSUBS 0.007001f
C1482 B.n552 VSUBS 0.007001f
C1483 B.n553 VSUBS 0.004118f
C1484 B.n554 VSUBS 0.007001f
C1485 B.n555 VSUBS 0.007001f
C1486 B.n556 VSUBS 0.007001f
C1487 B.n557 VSUBS 0.007001f
C1488 B.n558 VSUBS 0.007001f
C1489 B.n559 VSUBS 0.007001f
C1490 B.n560 VSUBS 0.007001f
C1491 B.n561 VSUBS 0.007001f
C1492 B.n562 VSUBS 0.007001f
C1493 B.n563 VSUBS 0.007001f
C1494 B.n564 VSUBS 0.007001f
C1495 B.n565 VSUBS 0.007001f
C1496 B.n566 VSUBS 0.007001f
C1497 B.n567 VSUBS 0.007001f
C1498 B.n568 VSUBS 0.007001f
C1499 B.n569 VSUBS 0.007001f
C1500 B.n570 VSUBS 0.007001f
C1501 B.n571 VSUBS 0.007001f
C1502 B.n572 VSUBS 0.007001f
C1503 B.n573 VSUBS 0.007001f
C1504 B.n574 VSUBS 0.007001f
C1505 B.n575 VSUBS 0.007001f
C1506 B.n576 VSUBS 0.007001f
C1507 B.n577 VSUBS 0.007001f
C1508 B.n578 VSUBS 0.007001f
C1509 B.n579 VSUBS 0.007001f
C1510 B.n580 VSUBS 0.007001f
C1511 B.n581 VSUBS 0.007001f
C1512 B.n582 VSUBS 0.007001f
C1513 B.n583 VSUBS 0.007001f
C1514 B.n584 VSUBS 0.007001f
C1515 B.n585 VSUBS 0.007001f
C1516 B.n586 VSUBS 0.007001f
C1517 B.n587 VSUBS 0.007001f
C1518 B.n588 VSUBS 0.007001f
C1519 B.n589 VSUBS 0.007001f
C1520 B.n590 VSUBS 0.007001f
C1521 B.n591 VSUBS 0.007001f
C1522 B.n592 VSUBS 0.007001f
C1523 B.n593 VSUBS 0.007001f
C1524 B.n594 VSUBS 0.007001f
C1525 B.n595 VSUBS 0.007001f
C1526 B.n596 VSUBS 0.007001f
C1527 B.n597 VSUBS 0.007001f
C1528 B.n598 VSUBS 0.007001f
C1529 B.n599 VSUBS 0.007001f
C1530 B.n600 VSUBS 0.007001f
C1531 B.n601 VSUBS 0.007001f
C1532 B.n602 VSUBS 0.007001f
C1533 B.n603 VSUBS 0.007001f
C1534 B.n604 VSUBS 0.007001f
C1535 B.n605 VSUBS 0.007001f
C1536 B.n606 VSUBS 0.007001f
C1537 B.n607 VSUBS 0.007001f
C1538 B.n608 VSUBS 0.007001f
C1539 B.n609 VSUBS 0.007001f
C1540 B.n610 VSUBS 0.007001f
C1541 B.n611 VSUBS 0.007001f
C1542 B.n612 VSUBS 0.007001f
C1543 B.n613 VSUBS 0.007001f
C1544 B.n614 VSUBS 0.007001f
C1545 B.n615 VSUBS 0.007001f
C1546 B.n616 VSUBS 0.007001f
C1547 B.n617 VSUBS 0.007001f
C1548 B.n618 VSUBS 0.007001f
C1549 B.n619 VSUBS 0.007001f
C1550 B.n620 VSUBS 0.007001f
C1551 B.n621 VSUBS 0.007001f
C1552 B.n622 VSUBS 0.007001f
C1553 B.n623 VSUBS 0.007001f
C1554 B.n624 VSUBS 0.007001f
C1555 B.n625 VSUBS 0.007001f
C1556 B.n626 VSUBS 0.007001f
C1557 B.n627 VSUBS 0.007001f
C1558 B.n628 VSUBS 0.007001f
C1559 B.n629 VSUBS 0.007001f
C1560 B.n630 VSUBS 0.007001f
C1561 B.n631 VSUBS 0.007001f
C1562 B.n632 VSUBS 0.007001f
C1563 B.n633 VSUBS 0.007001f
C1564 B.n634 VSUBS 0.007001f
C1565 B.n635 VSUBS 0.007001f
C1566 B.n636 VSUBS 0.007001f
C1567 B.n637 VSUBS 0.007001f
C1568 B.n638 VSUBS 0.007001f
C1569 B.n639 VSUBS 0.007001f
C1570 B.n640 VSUBS 0.007001f
C1571 B.n641 VSUBS 0.007001f
C1572 B.n642 VSUBS 0.007001f
C1573 B.n643 VSUBS 0.007001f
C1574 B.n644 VSUBS 0.007001f
C1575 B.n645 VSUBS 0.007001f
C1576 B.n646 VSUBS 0.007001f
C1577 B.n647 VSUBS 0.007001f
C1578 B.n648 VSUBS 0.007001f
C1579 B.n649 VSUBS 0.017146f
C1580 B.n650 VSUBS 0.017146f
C1581 B.n651 VSUBS 0.016625f
C1582 B.n652 VSUBS 0.007001f
C1583 B.n653 VSUBS 0.007001f
C1584 B.n654 VSUBS 0.007001f
C1585 B.n655 VSUBS 0.007001f
C1586 B.n656 VSUBS 0.007001f
C1587 B.n657 VSUBS 0.007001f
C1588 B.n658 VSUBS 0.007001f
C1589 B.n659 VSUBS 0.007001f
C1590 B.n660 VSUBS 0.007001f
C1591 B.n661 VSUBS 0.007001f
C1592 B.n662 VSUBS 0.007001f
C1593 B.n663 VSUBS 0.007001f
C1594 B.n664 VSUBS 0.007001f
C1595 B.n665 VSUBS 0.007001f
C1596 B.n666 VSUBS 0.007001f
C1597 B.n667 VSUBS 0.007001f
C1598 B.n668 VSUBS 0.007001f
C1599 B.n669 VSUBS 0.007001f
C1600 B.n670 VSUBS 0.007001f
C1601 B.n671 VSUBS 0.015853f
.ends

