* NGSPICE file created from diff_pair_sample_1000.ext - technology: sky130A

.subckt diff_pair_sample_1000 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t14 B.t5 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=4.3095 ps=22.88 w=11.05 l=2.53
X1 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=0 ps=0 w=11.05 l=2.53
X2 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=0 ps=0 w=11.05 l=2.53
X3 VTAIL.t1 VP.t0 VDD1.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=1.82325 ps=11.38 w=11.05 l=2.53
X4 VDD2.t6 VN.t1 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X5 VTAIL.t3 VP.t1 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=1.82325 ps=11.38 w=11.05 l=2.53
X6 VDD1.t5 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X7 VTAIL.t7 VP.t3 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X8 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=0 ps=0 w=11.05 l=2.53
X9 VDD1.t3 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=4.3095 ps=22.88 w=11.05 l=2.53
X10 VTAIL.t11 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=1.82325 ps=11.38 w=11.05 l=2.53
X11 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X12 VTAIL.t9 VN.t3 VDD2.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X13 VDD2.t3 VN.t4 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X14 VDD1.t1 VP.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X15 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=0 ps=0 w=11.05 l=2.53
X16 VDD2.t2 VN.t5 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=4.3095 ps=22.88 w=11.05 l=2.53
X17 VDD1.t0 VP.t7 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=4.3095 ps=22.88 w=11.05 l=2.53
X18 VTAIL.t15 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.82325 pd=11.38 as=1.82325 ps=11.38 w=11.05 l=2.53
X19 VTAIL.t13 VN.t7 VDD2.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=4.3095 pd=22.88 as=1.82325 ps=11.38 w=11.05 l=2.53
R0 VN.n51 VN.n27 161.3
R1 VN.n50 VN.n49 161.3
R2 VN.n48 VN.n28 161.3
R3 VN.n47 VN.n46 161.3
R4 VN.n45 VN.n29 161.3
R5 VN.n44 VN.n43 161.3
R6 VN.n42 VN.n41 161.3
R7 VN.n40 VN.n31 161.3
R8 VN.n39 VN.n38 161.3
R9 VN.n37 VN.n32 161.3
R10 VN.n36 VN.n35 161.3
R11 VN.n24 VN.n0 161.3
R12 VN.n23 VN.n22 161.3
R13 VN.n21 VN.n1 161.3
R14 VN.n20 VN.n19 161.3
R15 VN.n18 VN.n2 161.3
R16 VN.n17 VN.n16 161.3
R17 VN.n15 VN.n14 161.3
R18 VN.n13 VN.n4 161.3
R19 VN.n12 VN.n11 161.3
R20 VN.n10 VN.n5 161.3
R21 VN.n9 VN.n8 161.3
R22 VN.n6 VN.t7 140.048
R23 VN.n33 VN.t5 140.048
R24 VN.n7 VN.t4 105.26
R25 VN.n3 VN.t3 105.26
R26 VN.n25 VN.t0 105.26
R27 VN.n34 VN.t6 105.26
R28 VN.n30 VN.t1 105.26
R29 VN.n52 VN.t2 105.26
R30 VN.n26 VN.n25 96.5656
R31 VN.n53 VN.n52 96.5656
R32 VN.n19 VN.n1 54.0911
R33 VN.n46 VN.n28 54.0911
R34 VN.n7 VN.n6 51.6001
R35 VN.n34 VN.n33 51.6001
R36 VN VN.n53 50.1951
R37 VN.n12 VN.n5 40.4934
R38 VN.n13 VN.n12 40.4934
R39 VN.n39 VN.n32 40.4934
R40 VN.n40 VN.n39 40.4934
R41 VN.n23 VN.n1 26.8957
R42 VN.n50 VN.n28 26.8957
R43 VN.n8 VN.n5 24.4675
R44 VN.n14 VN.n13 24.4675
R45 VN.n18 VN.n17 24.4675
R46 VN.n19 VN.n18 24.4675
R47 VN.n24 VN.n23 24.4675
R48 VN.n35 VN.n32 24.4675
R49 VN.n46 VN.n45 24.4675
R50 VN.n45 VN.n44 24.4675
R51 VN.n41 VN.n40 24.4675
R52 VN.n51 VN.n50 24.4675
R53 VN.n8 VN.n7 21.0421
R54 VN.n14 VN.n3 21.0421
R55 VN.n35 VN.n34 21.0421
R56 VN.n41 VN.n30 21.0421
R57 VN.n25 VN.n24 14.1914
R58 VN.n52 VN.n51 14.1914
R59 VN.n36 VN.n33 6.57419
R60 VN.n9 VN.n6 6.57419
R61 VN.n17 VN.n3 3.42588
R62 VN.n44 VN.n30 3.42588
R63 VN.n53 VN.n27 0.278367
R64 VN.n26 VN.n0 0.278367
R65 VN.n49 VN.n27 0.189894
R66 VN.n49 VN.n48 0.189894
R67 VN.n48 VN.n47 0.189894
R68 VN.n47 VN.n29 0.189894
R69 VN.n43 VN.n29 0.189894
R70 VN.n43 VN.n42 0.189894
R71 VN.n42 VN.n31 0.189894
R72 VN.n38 VN.n31 0.189894
R73 VN.n38 VN.n37 0.189894
R74 VN.n37 VN.n36 0.189894
R75 VN.n10 VN.n9 0.189894
R76 VN.n11 VN.n10 0.189894
R77 VN.n11 VN.n4 0.189894
R78 VN.n15 VN.n4 0.189894
R79 VN.n16 VN.n15 0.189894
R80 VN.n16 VN.n2 0.189894
R81 VN.n20 VN.n2 0.189894
R82 VN.n21 VN.n20 0.189894
R83 VN.n22 VN.n21 0.189894
R84 VN.n22 VN.n0 0.189894
R85 VN VN.n26 0.153454
R86 VTAIL.n11 VTAIL.t1 47.5161
R87 VTAIL.n10 VTAIL.t10 47.5161
R88 VTAIL.n7 VTAIL.t11 47.5161
R89 VTAIL.n15 VTAIL.t14 47.516
R90 VTAIL.n2 VTAIL.t13 47.516
R91 VTAIL.n3 VTAIL.t4 47.516
R92 VTAIL.n6 VTAIL.t3 47.516
R93 VTAIL.n14 VTAIL.t5 47.516
R94 VTAIL.n13 VTAIL.n12 45.7243
R95 VTAIL.n9 VTAIL.n8 45.7243
R96 VTAIL.n1 VTAIL.n0 45.7241
R97 VTAIL.n5 VTAIL.n4 45.7241
R98 VTAIL.n15 VTAIL.n14 24.3583
R99 VTAIL.n7 VTAIL.n6 24.3583
R100 VTAIL.n9 VTAIL.n7 2.46602
R101 VTAIL.n10 VTAIL.n9 2.46602
R102 VTAIL.n13 VTAIL.n11 2.46602
R103 VTAIL.n14 VTAIL.n13 2.46602
R104 VTAIL.n6 VTAIL.n5 2.46602
R105 VTAIL.n5 VTAIL.n3 2.46602
R106 VTAIL.n2 VTAIL.n1 2.46602
R107 VTAIL VTAIL.n15 2.40783
R108 VTAIL.n0 VTAIL.t8 1.79236
R109 VTAIL.n0 VTAIL.t9 1.79236
R110 VTAIL.n4 VTAIL.t6 1.79236
R111 VTAIL.n4 VTAIL.t0 1.79236
R112 VTAIL.n12 VTAIL.t2 1.79236
R113 VTAIL.n12 VTAIL.t7 1.79236
R114 VTAIL.n8 VTAIL.t12 1.79236
R115 VTAIL.n8 VTAIL.t15 1.79236
R116 VTAIL.n11 VTAIL.n10 0.470328
R117 VTAIL.n3 VTAIL.n2 0.470328
R118 VTAIL VTAIL.n1 0.0586897
R119 VDD2.n2 VDD2.n1 63.5803
R120 VDD2.n2 VDD2.n0 63.5803
R121 VDD2 VDD2.n5 63.5775
R122 VDD2.n4 VDD2.n3 62.4031
R123 VDD2.n4 VDD2.n2 44.336
R124 VDD2.n5 VDD2.t1 1.79236
R125 VDD2.n5 VDD2.t2 1.79236
R126 VDD2.n3 VDD2.t5 1.79236
R127 VDD2.n3 VDD2.t6 1.79236
R128 VDD2.n1 VDD2.t4 1.79236
R129 VDD2.n1 VDD2.t7 1.79236
R130 VDD2.n0 VDD2.t0 1.79236
R131 VDD2.n0 VDD2.t3 1.79236
R132 VDD2 VDD2.n4 1.29145
R133 B.n676 B.n675 585
R134 B.n676 B.n92 585
R135 B.n679 B.n678 585
R136 B.n680 B.n140 585
R137 B.n682 B.n681 585
R138 B.n684 B.n139 585
R139 B.n687 B.n686 585
R140 B.n688 B.n138 585
R141 B.n690 B.n689 585
R142 B.n692 B.n137 585
R143 B.n695 B.n694 585
R144 B.n696 B.n136 585
R145 B.n698 B.n697 585
R146 B.n700 B.n135 585
R147 B.n703 B.n702 585
R148 B.n704 B.n134 585
R149 B.n706 B.n705 585
R150 B.n708 B.n133 585
R151 B.n711 B.n710 585
R152 B.n712 B.n132 585
R153 B.n714 B.n713 585
R154 B.n716 B.n131 585
R155 B.n719 B.n718 585
R156 B.n720 B.n130 585
R157 B.n722 B.n721 585
R158 B.n724 B.n129 585
R159 B.n727 B.n726 585
R160 B.n728 B.n128 585
R161 B.n730 B.n729 585
R162 B.n732 B.n127 585
R163 B.n735 B.n734 585
R164 B.n736 B.n126 585
R165 B.n738 B.n737 585
R166 B.n740 B.n125 585
R167 B.n743 B.n742 585
R168 B.n744 B.n124 585
R169 B.n746 B.n745 585
R170 B.n748 B.n123 585
R171 B.n751 B.n750 585
R172 B.n752 B.n120 585
R173 B.n755 B.n754 585
R174 B.n757 B.n119 585
R175 B.n760 B.n759 585
R176 B.n761 B.n118 585
R177 B.n763 B.n762 585
R178 B.n765 B.n117 585
R179 B.n768 B.n767 585
R180 B.n769 B.n113 585
R181 B.n771 B.n770 585
R182 B.n773 B.n112 585
R183 B.n776 B.n775 585
R184 B.n777 B.n111 585
R185 B.n779 B.n778 585
R186 B.n781 B.n110 585
R187 B.n784 B.n783 585
R188 B.n785 B.n109 585
R189 B.n787 B.n786 585
R190 B.n789 B.n108 585
R191 B.n792 B.n791 585
R192 B.n793 B.n107 585
R193 B.n795 B.n794 585
R194 B.n797 B.n106 585
R195 B.n800 B.n799 585
R196 B.n801 B.n105 585
R197 B.n803 B.n802 585
R198 B.n805 B.n104 585
R199 B.n808 B.n807 585
R200 B.n809 B.n103 585
R201 B.n811 B.n810 585
R202 B.n813 B.n102 585
R203 B.n816 B.n815 585
R204 B.n817 B.n101 585
R205 B.n819 B.n818 585
R206 B.n821 B.n100 585
R207 B.n824 B.n823 585
R208 B.n825 B.n99 585
R209 B.n827 B.n826 585
R210 B.n829 B.n98 585
R211 B.n832 B.n831 585
R212 B.n833 B.n97 585
R213 B.n835 B.n834 585
R214 B.n837 B.n96 585
R215 B.n840 B.n839 585
R216 B.n841 B.n95 585
R217 B.n843 B.n842 585
R218 B.n845 B.n94 585
R219 B.n848 B.n847 585
R220 B.n849 B.n93 585
R221 B.n674 B.n91 585
R222 B.n852 B.n91 585
R223 B.n673 B.n90 585
R224 B.n853 B.n90 585
R225 B.n672 B.n89 585
R226 B.n854 B.n89 585
R227 B.n671 B.n670 585
R228 B.n670 B.n85 585
R229 B.n669 B.n84 585
R230 B.n860 B.n84 585
R231 B.n668 B.n83 585
R232 B.n861 B.n83 585
R233 B.n667 B.n82 585
R234 B.n862 B.n82 585
R235 B.n666 B.n665 585
R236 B.n665 B.n81 585
R237 B.n664 B.n77 585
R238 B.n868 B.n77 585
R239 B.n663 B.n76 585
R240 B.n869 B.n76 585
R241 B.n662 B.n75 585
R242 B.n870 B.n75 585
R243 B.n661 B.n660 585
R244 B.n660 B.n71 585
R245 B.n659 B.n70 585
R246 B.n876 B.n70 585
R247 B.n658 B.n69 585
R248 B.n877 B.n69 585
R249 B.n657 B.n68 585
R250 B.n878 B.n68 585
R251 B.n656 B.n655 585
R252 B.n655 B.n64 585
R253 B.n654 B.n63 585
R254 B.n884 B.n63 585
R255 B.n653 B.n62 585
R256 B.n885 B.n62 585
R257 B.n652 B.n61 585
R258 B.n886 B.n61 585
R259 B.n651 B.n650 585
R260 B.n650 B.n57 585
R261 B.n649 B.n56 585
R262 B.n892 B.n56 585
R263 B.n648 B.n55 585
R264 B.n893 B.n55 585
R265 B.n647 B.n54 585
R266 B.n894 B.n54 585
R267 B.n646 B.n645 585
R268 B.n645 B.n50 585
R269 B.n644 B.n49 585
R270 B.n900 B.n49 585
R271 B.n643 B.n48 585
R272 B.n901 B.n48 585
R273 B.n642 B.n47 585
R274 B.n902 B.n47 585
R275 B.n641 B.n640 585
R276 B.n640 B.n46 585
R277 B.n639 B.n42 585
R278 B.n908 B.n42 585
R279 B.n638 B.n41 585
R280 B.n909 B.n41 585
R281 B.n637 B.n40 585
R282 B.n910 B.n40 585
R283 B.n636 B.n635 585
R284 B.n635 B.n36 585
R285 B.n634 B.n35 585
R286 B.n916 B.n35 585
R287 B.n633 B.n34 585
R288 B.n917 B.n34 585
R289 B.n632 B.n33 585
R290 B.n918 B.n33 585
R291 B.n631 B.n630 585
R292 B.n630 B.n32 585
R293 B.n629 B.n28 585
R294 B.n924 B.n28 585
R295 B.n628 B.n27 585
R296 B.n925 B.n27 585
R297 B.n627 B.n26 585
R298 B.n926 B.n26 585
R299 B.n626 B.n625 585
R300 B.n625 B.n22 585
R301 B.n624 B.n21 585
R302 B.n932 B.n21 585
R303 B.n623 B.n20 585
R304 B.n933 B.n20 585
R305 B.n622 B.n19 585
R306 B.n934 B.n19 585
R307 B.n621 B.n620 585
R308 B.n620 B.n15 585
R309 B.n619 B.n14 585
R310 B.n940 B.n14 585
R311 B.n618 B.n13 585
R312 B.n941 B.n13 585
R313 B.n617 B.n12 585
R314 B.n942 B.n12 585
R315 B.n616 B.n615 585
R316 B.n615 B.n8 585
R317 B.n614 B.n7 585
R318 B.n948 B.n7 585
R319 B.n613 B.n6 585
R320 B.n949 B.n6 585
R321 B.n612 B.n5 585
R322 B.n950 B.n5 585
R323 B.n611 B.n610 585
R324 B.n610 B.n4 585
R325 B.n609 B.n141 585
R326 B.n609 B.n608 585
R327 B.n599 B.n142 585
R328 B.n143 B.n142 585
R329 B.n601 B.n600 585
R330 B.n602 B.n601 585
R331 B.n598 B.n148 585
R332 B.n148 B.n147 585
R333 B.n597 B.n596 585
R334 B.n596 B.n595 585
R335 B.n150 B.n149 585
R336 B.n151 B.n150 585
R337 B.n588 B.n587 585
R338 B.n589 B.n588 585
R339 B.n586 B.n156 585
R340 B.n156 B.n155 585
R341 B.n585 B.n584 585
R342 B.n584 B.n583 585
R343 B.n158 B.n157 585
R344 B.n159 B.n158 585
R345 B.n576 B.n575 585
R346 B.n577 B.n576 585
R347 B.n574 B.n164 585
R348 B.n164 B.n163 585
R349 B.n573 B.n572 585
R350 B.n572 B.n571 585
R351 B.n166 B.n165 585
R352 B.n564 B.n166 585
R353 B.n563 B.n562 585
R354 B.n565 B.n563 585
R355 B.n561 B.n171 585
R356 B.n171 B.n170 585
R357 B.n560 B.n559 585
R358 B.n559 B.n558 585
R359 B.n173 B.n172 585
R360 B.n174 B.n173 585
R361 B.n551 B.n550 585
R362 B.n552 B.n551 585
R363 B.n549 B.n179 585
R364 B.n179 B.n178 585
R365 B.n548 B.n547 585
R366 B.n547 B.n546 585
R367 B.n181 B.n180 585
R368 B.n539 B.n181 585
R369 B.n538 B.n537 585
R370 B.n540 B.n538 585
R371 B.n536 B.n186 585
R372 B.n186 B.n185 585
R373 B.n535 B.n534 585
R374 B.n534 B.n533 585
R375 B.n188 B.n187 585
R376 B.n189 B.n188 585
R377 B.n526 B.n525 585
R378 B.n527 B.n526 585
R379 B.n524 B.n194 585
R380 B.n194 B.n193 585
R381 B.n523 B.n522 585
R382 B.n522 B.n521 585
R383 B.n196 B.n195 585
R384 B.n197 B.n196 585
R385 B.n514 B.n513 585
R386 B.n515 B.n514 585
R387 B.n512 B.n202 585
R388 B.n202 B.n201 585
R389 B.n511 B.n510 585
R390 B.n510 B.n509 585
R391 B.n204 B.n203 585
R392 B.n205 B.n204 585
R393 B.n502 B.n501 585
R394 B.n503 B.n502 585
R395 B.n500 B.n210 585
R396 B.n210 B.n209 585
R397 B.n499 B.n498 585
R398 B.n498 B.n497 585
R399 B.n212 B.n211 585
R400 B.n213 B.n212 585
R401 B.n490 B.n489 585
R402 B.n491 B.n490 585
R403 B.n488 B.n218 585
R404 B.n218 B.n217 585
R405 B.n487 B.n486 585
R406 B.n486 B.n485 585
R407 B.n220 B.n219 585
R408 B.n478 B.n220 585
R409 B.n477 B.n476 585
R410 B.n479 B.n477 585
R411 B.n475 B.n225 585
R412 B.n225 B.n224 585
R413 B.n474 B.n473 585
R414 B.n473 B.n472 585
R415 B.n227 B.n226 585
R416 B.n228 B.n227 585
R417 B.n465 B.n464 585
R418 B.n466 B.n465 585
R419 B.n463 B.n233 585
R420 B.n233 B.n232 585
R421 B.n462 B.n461 585
R422 B.n461 B.n460 585
R423 B.n457 B.n237 585
R424 B.n456 B.n455 585
R425 B.n453 B.n238 585
R426 B.n453 B.n236 585
R427 B.n452 B.n451 585
R428 B.n450 B.n449 585
R429 B.n448 B.n240 585
R430 B.n446 B.n445 585
R431 B.n444 B.n241 585
R432 B.n443 B.n442 585
R433 B.n440 B.n242 585
R434 B.n438 B.n437 585
R435 B.n436 B.n243 585
R436 B.n435 B.n434 585
R437 B.n432 B.n244 585
R438 B.n430 B.n429 585
R439 B.n428 B.n245 585
R440 B.n427 B.n426 585
R441 B.n424 B.n246 585
R442 B.n422 B.n421 585
R443 B.n420 B.n247 585
R444 B.n419 B.n418 585
R445 B.n416 B.n248 585
R446 B.n414 B.n413 585
R447 B.n412 B.n249 585
R448 B.n411 B.n410 585
R449 B.n408 B.n250 585
R450 B.n406 B.n405 585
R451 B.n404 B.n251 585
R452 B.n403 B.n402 585
R453 B.n400 B.n252 585
R454 B.n398 B.n397 585
R455 B.n396 B.n253 585
R456 B.n395 B.n394 585
R457 B.n392 B.n254 585
R458 B.n390 B.n389 585
R459 B.n388 B.n255 585
R460 B.n387 B.n386 585
R461 B.n384 B.n256 585
R462 B.n382 B.n381 585
R463 B.n379 B.n257 585
R464 B.n378 B.n377 585
R465 B.n375 B.n260 585
R466 B.n373 B.n372 585
R467 B.n371 B.n261 585
R468 B.n370 B.n369 585
R469 B.n367 B.n262 585
R470 B.n365 B.n364 585
R471 B.n363 B.n263 585
R472 B.n361 B.n360 585
R473 B.n358 B.n266 585
R474 B.n356 B.n355 585
R475 B.n354 B.n267 585
R476 B.n353 B.n352 585
R477 B.n350 B.n268 585
R478 B.n348 B.n347 585
R479 B.n346 B.n269 585
R480 B.n345 B.n344 585
R481 B.n342 B.n270 585
R482 B.n340 B.n339 585
R483 B.n338 B.n271 585
R484 B.n337 B.n336 585
R485 B.n334 B.n272 585
R486 B.n332 B.n331 585
R487 B.n330 B.n273 585
R488 B.n329 B.n328 585
R489 B.n326 B.n274 585
R490 B.n324 B.n323 585
R491 B.n322 B.n275 585
R492 B.n321 B.n320 585
R493 B.n318 B.n276 585
R494 B.n316 B.n315 585
R495 B.n314 B.n277 585
R496 B.n313 B.n312 585
R497 B.n310 B.n278 585
R498 B.n308 B.n307 585
R499 B.n306 B.n279 585
R500 B.n305 B.n304 585
R501 B.n302 B.n280 585
R502 B.n300 B.n299 585
R503 B.n298 B.n281 585
R504 B.n297 B.n296 585
R505 B.n294 B.n282 585
R506 B.n292 B.n291 585
R507 B.n290 B.n283 585
R508 B.n289 B.n288 585
R509 B.n286 B.n284 585
R510 B.n235 B.n234 585
R511 B.n459 B.n458 585
R512 B.n460 B.n459 585
R513 B.n231 B.n230 585
R514 B.n232 B.n231 585
R515 B.n468 B.n467 585
R516 B.n467 B.n466 585
R517 B.n469 B.n229 585
R518 B.n229 B.n228 585
R519 B.n471 B.n470 585
R520 B.n472 B.n471 585
R521 B.n223 B.n222 585
R522 B.n224 B.n223 585
R523 B.n481 B.n480 585
R524 B.n480 B.n479 585
R525 B.n482 B.n221 585
R526 B.n478 B.n221 585
R527 B.n484 B.n483 585
R528 B.n485 B.n484 585
R529 B.n216 B.n215 585
R530 B.n217 B.n216 585
R531 B.n493 B.n492 585
R532 B.n492 B.n491 585
R533 B.n494 B.n214 585
R534 B.n214 B.n213 585
R535 B.n496 B.n495 585
R536 B.n497 B.n496 585
R537 B.n208 B.n207 585
R538 B.n209 B.n208 585
R539 B.n505 B.n504 585
R540 B.n504 B.n503 585
R541 B.n506 B.n206 585
R542 B.n206 B.n205 585
R543 B.n508 B.n507 585
R544 B.n509 B.n508 585
R545 B.n200 B.n199 585
R546 B.n201 B.n200 585
R547 B.n517 B.n516 585
R548 B.n516 B.n515 585
R549 B.n518 B.n198 585
R550 B.n198 B.n197 585
R551 B.n520 B.n519 585
R552 B.n521 B.n520 585
R553 B.n192 B.n191 585
R554 B.n193 B.n192 585
R555 B.n529 B.n528 585
R556 B.n528 B.n527 585
R557 B.n530 B.n190 585
R558 B.n190 B.n189 585
R559 B.n532 B.n531 585
R560 B.n533 B.n532 585
R561 B.n184 B.n183 585
R562 B.n185 B.n184 585
R563 B.n542 B.n541 585
R564 B.n541 B.n540 585
R565 B.n543 B.n182 585
R566 B.n539 B.n182 585
R567 B.n545 B.n544 585
R568 B.n546 B.n545 585
R569 B.n177 B.n176 585
R570 B.n178 B.n177 585
R571 B.n554 B.n553 585
R572 B.n553 B.n552 585
R573 B.n555 B.n175 585
R574 B.n175 B.n174 585
R575 B.n557 B.n556 585
R576 B.n558 B.n557 585
R577 B.n169 B.n168 585
R578 B.n170 B.n169 585
R579 B.n567 B.n566 585
R580 B.n566 B.n565 585
R581 B.n568 B.n167 585
R582 B.n564 B.n167 585
R583 B.n570 B.n569 585
R584 B.n571 B.n570 585
R585 B.n162 B.n161 585
R586 B.n163 B.n162 585
R587 B.n579 B.n578 585
R588 B.n578 B.n577 585
R589 B.n580 B.n160 585
R590 B.n160 B.n159 585
R591 B.n582 B.n581 585
R592 B.n583 B.n582 585
R593 B.n154 B.n153 585
R594 B.n155 B.n154 585
R595 B.n591 B.n590 585
R596 B.n590 B.n589 585
R597 B.n592 B.n152 585
R598 B.n152 B.n151 585
R599 B.n594 B.n593 585
R600 B.n595 B.n594 585
R601 B.n146 B.n145 585
R602 B.n147 B.n146 585
R603 B.n604 B.n603 585
R604 B.n603 B.n602 585
R605 B.n605 B.n144 585
R606 B.n144 B.n143 585
R607 B.n607 B.n606 585
R608 B.n608 B.n607 585
R609 B.n2 B.n0 585
R610 B.n4 B.n2 585
R611 B.n3 B.n1 585
R612 B.n949 B.n3 585
R613 B.n947 B.n946 585
R614 B.n948 B.n947 585
R615 B.n945 B.n9 585
R616 B.n9 B.n8 585
R617 B.n944 B.n943 585
R618 B.n943 B.n942 585
R619 B.n11 B.n10 585
R620 B.n941 B.n11 585
R621 B.n939 B.n938 585
R622 B.n940 B.n939 585
R623 B.n937 B.n16 585
R624 B.n16 B.n15 585
R625 B.n936 B.n935 585
R626 B.n935 B.n934 585
R627 B.n18 B.n17 585
R628 B.n933 B.n18 585
R629 B.n931 B.n930 585
R630 B.n932 B.n931 585
R631 B.n929 B.n23 585
R632 B.n23 B.n22 585
R633 B.n928 B.n927 585
R634 B.n927 B.n926 585
R635 B.n25 B.n24 585
R636 B.n925 B.n25 585
R637 B.n923 B.n922 585
R638 B.n924 B.n923 585
R639 B.n921 B.n29 585
R640 B.n32 B.n29 585
R641 B.n920 B.n919 585
R642 B.n919 B.n918 585
R643 B.n31 B.n30 585
R644 B.n917 B.n31 585
R645 B.n915 B.n914 585
R646 B.n916 B.n915 585
R647 B.n913 B.n37 585
R648 B.n37 B.n36 585
R649 B.n912 B.n911 585
R650 B.n911 B.n910 585
R651 B.n39 B.n38 585
R652 B.n909 B.n39 585
R653 B.n907 B.n906 585
R654 B.n908 B.n907 585
R655 B.n905 B.n43 585
R656 B.n46 B.n43 585
R657 B.n904 B.n903 585
R658 B.n903 B.n902 585
R659 B.n45 B.n44 585
R660 B.n901 B.n45 585
R661 B.n899 B.n898 585
R662 B.n900 B.n899 585
R663 B.n897 B.n51 585
R664 B.n51 B.n50 585
R665 B.n896 B.n895 585
R666 B.n895 B.n894 585
R667 B.n53 B.n52 585
R668 B.n893 B.n53 585
R669 B.n891 B.n890 585
R670 B.n892 B.n891 585
R671 B.n889 B.n58 585
R672 B.n58 B.n57 585
R673 B.n888 B.n887 585
R674 B.n887 B.n886 585
R675 B.n60 B.n59 585
R676 B.n885 B.n60 585
R677 B.n883 B.n882 585
R678 B.n884 B.n883 585
R679 B.n881 B.n65 585
R680 B.n65 B.n64 585
R681 B.n880 B.n879 585
R682 B.n879 B.n878 585
R683 B.n67 B.n66 585
R684 B.n877 B.n67 585
R685 B.n875 B.n874 585
R686 B.n876 B.n875 585
R687 B.n873 B.n72 585
R688 B.n72 B.n71 585
R689 B.n872 B.n871 585
R690 B.n871 B.n870 585
R691 B.n74 B.n73 585
R692 B.n869 B.n74 585
R693 B.n867 B.n866 585
R694 B.n868 B.n867 585
R695 B.n865 B.n78 585
R696 B.n81 B.n78 585
R697 B.n864 B.n863 585
R698 B.n863 B.n862 585
R699 B.n80 B.n79 585
R700 B.n861 B.n80 585
R701 B.n859 B.n858 585
R702 B.n860 B.n859 585
R703 B.n857 B.n86 585
R704 B.n86 B.n85 585
R705 B.n856 B.n855 585
R706 B.n855 B.n854 585
R707 B.n88 B.n87 585
R708 B.n853 B.n88 585
R709 B.n851 B.n850 585
R710 B.n852 B.n851 585
R711 B.n952 B.n951 585
R712 B.n951 B.n950 585
R713 B.n459 B.n237 545.355
R714 B.n851 B.n93 545.355
R715 B.n461 B.n235 545.355
R716 B.n676 B.n91 545.355
R717 B.n264 B.t8 313.197
R718 B.n258 B.t19 313.197
R719 B.n114 B.t16 313.197
R720 B.n121 B.t12 313.197
R721 B.n677 B.n92 256.663
R722 B.n683 B.n92 256.663
R723 B.n685 B.n92 256.663
R724 B.n691 B.n92 256.663
R725 B.n693 B.n92 256.663
R726 B.n699 B.n92 256.663
R727 B.n701 B.n92 256.663
R728 B.n707 B.n92 256.663
R729 B.n709 B.n92 256.663
R730 B.n715 B.n92 256.663
R731 B.n717 B.n92 256.663
R732 B.n723 B.n92 256.663
R733 B.n725 B.n92 256.663
R734 B.n731 B.n92 256.663
R735 B.n733 B.n92 256.663
R736 B.n739 B.n92 256.663
R737 B.n741 B.n92 256.663
R738 B.n747 B.n92 256.663
R739 B.n749 B.n92 256.663
R740 B.n756 B.n92 256.663
R741 B.n758 B.n92 256.663
R742 B.n764 B.n92 256.663
R743 B.n766 B.n92 256.663
R744 B.n772 B.n92 256.663
R745 B.n774 B.n92 256.663
R746 B.n780 B.n92 256.663
R747 B.n782 B.n92 256.663
R748 B.n788 B.n92 256.663
R749 B.n790 B.n92 256.663
R750 B.n796 B.n92 256.663
R751 B.n798 B.n92 256.663
R752 B.n804 B.n92 256.663
R753 B.n806 B.n92 256.663
R754 B.n812 B.n92 256.663
R755 B.n814 B.n92 256.663
R756 B.n820 B.n92 256.663
R757 B.n822 B.n92 256.663
R758 B.n828 B.n92 256.663
R759 B.n830 B.n92 256.663
R760 B.n836 B.n92 256.663
R761 B.n838 B.n92 256.663
R762 B.n844 B.n92 256.663
R763 B.n846 B.n92 256.663
R764 B.n454 B.n236 256.663
R765 B.n239 B.n236 256.663
R766 B.n447 B.n236 256.663
R767 B.n441 B.n236 256.663
R768 B.n439 B.n236 256.663
R769 B.n433 B.n236 256.663
R770 B.n431 B.n236 256.663
R771 B.n425 B.n236 256.663
R772 B.n423 B.n236 256.663
R773 B.n417 B.n236 256.663
R774 B.n415 B.n236 256.663
R775 B.n409 B.n236 256.663
R776 B.n407 B.n236 256.663
R777 B.n401 B.n236 256.663
R778 B.n399 B.n236 256.663
R779 B.n393 B.n236 256.663
R780 B.n391 B.n236 256.663
R781 B.n385 B.n236 256.663
R782 B.n383 B.n236 256.663
R783 B.n376 B.n236 256.663
R784 B.n374 B.n236 256.663
R785 B.n368 B.n236 256.663
R786 B.n366 B.n236 256.663
R787 B.n359 B.n236 256.663
R788 B.n357 B.n236 256.663
R789 B.n351 B.n236 256.663
R790 B.n349 B.n236 256.663
R791 B.n343 B.n236 256.663
R792 B.n341 B.n236 256.663
R793 B.n335 B.n236 256.663
R794 B.n333 B.n236 256.663
R795 B.n327 B.n236 256.663
R796 B.n325 B.n236 256.663
R797 B.n319 B.n236 256.663
R798 B.n317 B.n236 256.663
R799 B.n311 B.n236 256.663
R800 B.n309 B.n236 256.663
R801 B.n303 B.n236 256.663
R802 B.n301 B.n236 256.663
R803 B.n295 B.n236 256.663
R804 B.n293 B.n236 256.663
R805 B.n287 B.n236 256.663
R806 B.n285 B.n236 256.663
R807 B.n459 B.n231 163.367
R808 B.n467 B.n231 163.367
R809 B.n467 B.n229 163.367
R810 B.n471 B.n229 163.367
R811 B.n471 B.n223 163.367
R812 B.n480 B.n223 163.367
R813 B.n480 B.n221 163.367
R814 B.n484 B.n221 163.367
R815 B.n484 B.n216 163.367
R816 B.n492 B.n216 163.367
R817 B.n492 B.n214 163.367
R818 B.n496 B.n214 163.367
R819 B.n496 B.n208 163.367
R820 B.n504 B.n208 163.367
R821 B.n504 B.n206 163.367
R822 B.n508 B.n206 163.367
R823 B.n508 B.n200 163.367
R824 B.n516 B.n200 163.367
R825 B.n516 B.n198 163.367
R826 B.n520 B.n198 163.367
R827 B.n520 B.n192 163.367
R828 B.n528 B.n192 163.367
R829 B.n528 B.n190 163.367
R830 B.n532 B.n190 163.367
R831 B.n532 B.n184 163.367
R832 B.n541 B.n184 163.367
R833 B.n541 B.n182 163.367
R834 B.n545 B.n182 163.367
R835 B.n545 B.n177 163.367
R836 B.n553 B.n177 163.367
R837 B.n553 B.n175 163.367
R838 B.n557 B.n175 163.367
R839 B.n557 B.n169 163.367
R840 B.n566 B.n169 163.367
R841 B.n566 B.n167 163.367
R842 B.n570 B.n167 163.367
R843 B.n570 B.n162 163.367
R844 B.n578 B.n162 163.367
R845 B.n578 B.n160 163.367
R846 B.n582 B.n160 163.367
R847 B.n582 B.n154 163.367
R848 B.n590 B.n154 163.367
R849 B.n590 B.n152 163.367
R850 B.n594 B.n152 163.367
R851 B.n594 B.n146 163.367
R852 B.n603 B.n146 163.367
R853 B.n603 B.n144 163.367
R854 B.n607 B.n144 163.367
R855 B.n607 B.n2 163.367
R856 B.n951 B.n2 163.367
R857 B.n951 B.n3 163.367
R858 B.n947 B.n3 163.367
R859 B.n947 B.n9 163.367
R860 B.n943 B.n9 163.367
R861 B.n943 B.n11 163.367
R862 B.n939 B.n11 163.367
R863 B.n939 B.n16 163.367
R864 B.n935 B.n16 163.367
R865 B.n935 B.n18 163.367
R866 B.n931 B.n18 163.367
R867 B.n931 B.n23 163.367
R868 B.n927 B.n23 163.367
R869 B.n927 B.n25 163.367
R870 B.n923 B.n25 163.367
R871 B.n923 B.n29 163.367
R872 B.n919 B.n29 163.367
R873 B.n919 B.n31 163.367
R874 B.n915 B.n31 163.367
R875 B.n915 B.n37 163.367
R876 B.n911 B.n37 163.367
R877 B.n911 B.n39 163.367
R878 B.n907 B.n39 163.367
R879 B.n907 B.n43 163.367
R880 B.n903 B.n43 163.367
R881 B.n903 B.n45 163.367
R882 B.n899 B.n45 163.367
R883 B.n899 B.n51 163.367
R884 B.n895 B.n51 163.367
R885 B.n895 B.n53 163.367
R886 B.n891 B.n53 163.367
R887 B.n891 B.n58 163.367
R888 B.n887 B.n58 163.367
R889 B.n887 B.n60 163.367
R890 B.n883 B.n60 163.367
R891 B.n883 B.n65 163.367
R892 B.n879 B.n65 163.367
R893 B.n879 B.n67 163.367
R894 B.n875 B.n67 163.367
R895 B.n875 B.n72 163.367
R896 B.n871 B.n72 163.367
R897 B.n871 B.n74 163.367
R898 B.n867 B.n74 163.367
R899 B.n867 B.n78 163.367
R900 B.n863 B.n78 163.367
R901 B.n863 B.n80 163.367
R902 B.n859 B.n80 163.367
R903 B.n859 B.n86 163.367
R904 B.n855 B.n86 163.367
R905 B.n855 B.n88 163.367
R906 B.n851 B.n88 163.367
R907 B.n455 B.n453 163.367
R908 B.n453 B.n452 163.367
R909 B.n449 B.n448 163.367
R910 B.n446 B.n241 163.367
R911 B.n442 B.n440 163.367
R912 B.n438 B.n243 163.367
R913 B.n434 B.n432 163.367
R914 B.n430 B.n245 163.367
R915 B.n426 B.n424 163.367
R916 B.n422 B.n247 163.367
R917 B.n418 B.n416 163.367
R918 B.n414 B.n249 163.367
R919 B.n410 B.n408 163.367
R920 B.n406 B.n251 163.367
R921 B.n402 B.n400 163.367
R922 B.n398 B.n253 163.367
R923 B.n394 B.n392 163.367
R924 B.n390 B.n255 163.367
R925 B.n386 B.n384 163.367
R926 B.n382 B.n257 163.367
R927 B.n377 B.n375 163.367
R928 B.n373 B.n261 163.367
R929 B.n369 B.n367 163.367
R930 B.n365 B.n263 163.367
R931 B.n360 B.n358 163.367
R932 B.n356 B.n267 163.367
R933 B.n352 B.n350 163.367
R934 B.n348 B.n269 163.367
R935 B.n344 B.n342 163.367
R936 B.n340 B.n271 163.367
R937 B.n336 B.n334 163.367
R938 B.n332 B.n273 163.367
R939 B.n328 B.n326 163.367
R940 B.n324 B.n275 163.367
R941 B.n320 B.n318 163.367
R942 B.n316 B.n277 163.367
R943 B.n312 B.n310 163.367
R944 B.n308 B.n279 163.367
R945 B.n304 B.n302 163.367
R946 B.n300 B.n281 163.367
R947 B.n296 B.n294 163.367
R948 B.n292 B.n283 163.367
R949 B.n288 B.n286 163.367
R950 B.n461 B.n233 163.367
R951 B.n465 B.n233 163.367
R952 B.n465 B.n227 163.367
R953 B.n473 B.n227 163.367
R954 B.n473 B.n225 163.367
R955 B.n477 B.n225 163.367
R956 B.n477 B.n220 163.367
R957 B.n486 B.n220 163.367
R958 B.n486 B.n218 163.367
R959 B.n490 B.n218 163.367
R960 B.n490 B.n212 163.367
R961 B.n498 B.n212 163.367
R962 B.n498 B.n210 163.367
R963 B.n502 B.n210 163.367
R964 B.n502 B.n204 163.367
R965 B.n510 B.n204 163.367
R966 B.n510 B.n202 163.367
R967 B.n514 B.n202 163.367
R968 B.n514 B.n196 163.367
R969 B.n522 B.n196 163.367
R970 B.n522 B.n194 163.367
R971 B.n526 B.n194 163.367
R972 B.n526 B.n188 163.367
R973 B.n534 B.n188 163.367
R974 B.n534 B.n186 163.367
R975 B.n538 B.n186 163.367
R976 B.n538 B.n181 163.367
R977 B.n547 B.n181 163.367
R978 B.n547 B.n179 163.367
R979 B.n551 B.n179 163.367
R980 B.n551 B.n173 163.367
R981 B.n559 B.n173 163.367
R982 B.n559 B.n171 163.367
R983 B.n563 B.n171 163.367
R984 B.n563 B.n166 163.367
R985 B.n572 B.n166 163.367
R986 B.n572 B.n164 163.367
R987 B.n576 B.n164 163.367
R988 B.n576 B.n158 163.367
R989 B.n584 B.n158 163.367
R990 B.n584 B.n156 163.367
R991 B.n588 B.n156 163.367
R992 B.n588 B.n150 163.367
R993 B.n596 B.n150 163.367
R994 B.n596 B.n148 163.367
R995 B.n601 B.n148 163.367
R996 B.n601 B.n142 163.367
R997 B.n609 B.n142 163.367
R998 B.n610 B.n609 163.367
R999 B.n610 B.n5 163.367
R1000 B.n6 B.n5 163.367
R1001 B.n7 B.n6 163.367
R1002 B.n615 B.n7 163.367
R1003 B.n615 B.n12 163.367
R1004 B.n13 B.n12 163.367
R1005 B.n14 B.n13 163.367
R1006 B.n620 B.n14 163.367
R1007 B.n620 B.n19 163.367
R1008 B.n20 B.n19 163.367
R1009 B.n21 B.n20 163.367
R1010 B.n625 B.n21 163.367
R1011 B.n625 B.n26 163.367
R1012 B.n27 B.n26 163.367
R1013 B.n28 B.n27 163.367
R1014 B.n630 B.n28 163.367
R1015 B.n630 B.n33 163.367
R1016 B.n34 B.n33 163.367
R1017 B.n35 B.n34 163.367
R1018 B.n635 B.n35 163.367
R1019 B.n635 B.n40 163.367
R1020 B.n41 B.n40 163.367
R1021 B.n42 B.n41 163.367
R1022 B.n640 B.n42 163.367
R1023 B.n640 B.n47 163.367
R1024 B.n48 B.n47 163.367
R1025 B.n49 B.n48 163.367
R1026 B.n645 B.n49 163.367
R1027 B.n645 B.n54 163.367
R1028 B.n55 B.n54 163.367
R1029 B.n56 B.n55 163.367
R1030 B.n650 B.n56 163.367
R1031 B.n650 B.n61 163.367
R1032 B.n62 B.n61 163.367
R1033 B.n63 B.n62 163.367
R1034 B.n655 B.n63 163.367
R1035 B.n655 B.n68 163.367
R1036 B.n69 B.n68 163.367
R1037 B.n70 B.n69 163.367
R1038 B.n660 B.n70 163.367
R1039 B.n660 B.n75 163.367
R1040 B.n76 B.n75 163.367
R1041 B.n77 B.n76 163.367
R1042 B.n665 B.n77 163.367
R1043 B.n665 B.n82 163.367
R1044 B.n83 B.n82 163.367
R1045 B.n84 B.n83 163.367
R1046 B.n670 B.n84 163.367
R1047 B.n670 B.n89 163.367
R1048 B.n90 B.n89 163.367
R1049 B.n91 B.n90 163.367
R1050 B.n847 B.n845 163.367
R1051 B.n843 B.n95 163.367
R1052 B.n839 B.n837 163.367
R1053 B.n835 B.n97 163.367
R1054 B.n831 B.n829 163.367
R1055 B.n827 B.n99 163.367
R1056 B.n823 B.n821 163.367
R1057 B.n819 B.n101 163.367
R1058 B.n815 B.n813 163.367
R1059 B.n811 B.n103 163.367
R1060 B.n807 B.n805 163.367
R1061 B.n803 B.n105 163.367
R1062 B.n799 B.n797 163.367
R1063 B.n795 B.n107 163.367
R1064 B.n791 B.n789 163.367
R1065 B.n787 B.n109 163.367
R1066 B.n783 B.n781 163.367
R1067 B.n779 B.n111 163.367
R1068 B.n775 B.n773 163.367
R1069 B.n771 B.n113 163.367
R1070 B.n767 B.n765 163.367
R1071 B.n763 B.n118 163.367
R1072 B.n759 B.n757 163.367
R1073 B.n755 B.n120 163.367
R1074 B.n750 B.n748 163.367
R1075 B.n746 B.n124 163.367
R1076 B.n742 B.n740 163.367
R1077 B.n738 B.n126 163.367
R1078 B.n734 B.n732 163.367
R1079 B.n730 B.n128 163.367
R1080 B.n726 B.n724 163.367
R1081 B.n722 B.n130 163.367
R1082 B.n718 B.n716 163.367
R1083 B.n714 B.n132 163.367
R1084 B.n710 B.n708 163.367
R1085 B.n706 B.n134 163.367
R1086 B.n702 B.n700 163.367
R1087 B.n698 B.n136 163.367
R1088 B.n694 B.n692 163.367
R1089 B.n690 B.n138 163.367
R1090 B.n686 B.n684 163.367
R1091 B.n682 B.n140 163.367
R1092 B.n678 B.n676 163.367
R1093 B.n264 B.t11 126.694
R1094 B.n121 B.t14 126.694
R1095 B.n258 B.t21 126.68
R1096 B.n114 B.t17 126.68
R1097 B.n460 B.n236 90.9653
R1098 B.n852 B.n92 90.9653
R1099 B.n454 B.n237 71.676
R1100 B.n452 B.n239 71.676
R1101 B.n448 B.n447 71.676
R1102 B.n441 B.n241 71.676
R1103 B.n440 B.n439 71.676
R1104 B.n433 B.n243 71.676
R1105 B.n432 B.n431 71.676
R1106 B.n425 B.n245 71.676
R1107 B.n424 B.n423 71.676
R1108 B.n417 B.n247 71.676
R1109 B.n416 B.n415 71.676
R1110 B.n409 B.n249 71.676
R1111 B.n408 B.n407 71.676
R1112 B.n401 B.n251 71.676
R1113 B.n400 B.n399 71.676
R1114 B.n393 B.n253 71.676
R1115 B.n392 B.n391 71.676
R1116 B.n385 B.n255 71.676
R1117 B.n384 B.n383 71.676
R1118 B.n376 B.n257 71.676
R1119 B.n375 B.n374 71.676
R1120 B.n368 B.n261 71.676
R1121 B.n367 B.n366 71.676
R1122 B.n359 B.n263 71.676
R1123 B.n358 B.n357 71.676
R1124 B.n351 B.n267 71.676
R1125 B.n350 B.n349 71.676
R1126 B.n343 B.n269 71.676
R1127 B.n342 B.n341 71.676
R1128 B.n335 B.n271 71.676
R1129 B.n334 B.n333 71.676
R1130 B.n327 B.n273 71.676
R1131 B.n326 B.n325 71.676
R1132 B.n319 B.n275 71.676
R1133 B.n318 B.n317 71.676
R1134 B.n311 B.n277 71.676
R1135 B.n310 B.n309 71.676
R1136 B.n303 B.n279 71.676
R1137 B.n302 B.n301 71.676
R1138 B.n295 B.n281 71.676
R1139 B.n294 B.n293 71.676
R1140 B.n287 B.n283 71.676
R1141 B.n286 B.n285 71.676
R1142 B.n846 B.n93 71.676
R1143 B.n845 B.n844 71.676
R1144 B.n838 B.n95 71.676
R1145 B.n837 B.n836 71.676
R1146 B.n830 B.n97 71.676
R1147 B.n829 B.n828 71.676
R1148 B.n822 B.n99 71.676
R1149 B.n821 B.n820 71.676
R1150 B.n814 B.n101 71.676
R1151 B.n813 B.n812 71.676
R1152 B.n806 B.n103 71.676
R1153 B.n805 B.n804 71.676
R1154 B.n798 B.n105 71.676
R1155 B.n797 B.n796 71.676
R1156 B.n790 B.n107 71.676
R1157 B.n789 B.n788 71.676
R1158 B.n782 B.n109 71.676
R1159 B.n781 B.n780 71.676
R1160 B.n774 B.n111 71.676
R1161 B.n773 B.n772 71.676
R1162 B.n766 B.n113 71.676
R1163 B.n765 B.n764 71.676
R1164 B.n758 B.n118 71.676
R1165 B.n757 B.n756 71.676
R1166 B.n749 B.n120 71.676
R1167 B.n748 B.n747 71.676
R1168 B.n741 B.n124 71.676
R1169 B.n740 B.n739 71.676
R1170 B.n733 B.n126 71.676
R1171 B.n732 B.n731 71.676
R1172 B.n725 B.n128 71.676
R1173 B.n724 B.n723 71.676
R1174 B.n717 B.n130 71.676
R1175 B.n716 B.n715 71.676
R1176 B.n709 B.n132 71.676
R1177 B.n708 B.n707 71.676
R1178 B.n701 B.n134 71.676
R1179 B.n700 B.n699 71.676
R1180 B.n693 B.n136 71.676
R1181 B.n692 B.n691 71.676
R1182 B.n685 B.n138 71.676
R1183 B.n684 B.n683 71.676
R1184 B.n677 B.n140 71.676
R1185 B.n678 B.n677 71.676
R1186 B.n683 B.n682 71.676
R1187 B.n686 B.n685 71.676
R1188 B.n691 B.n690 71.676
R1189 B.n694 B.n693 71.676
R1190 B.n699 B.n698 71.676
R1191 B.n702 B.n701 71.676
R1192 B.n707 B.n706 71.676
R1193 B.n710 B.n709 71.676
R1194 B.n715 B.n714 71.676
R1195 B.n718 B.n717 71.676
R1196 B.n723 B.n722 71.676
R1197 B.n726 B.n725 71.676
R1198 B.n731 B.n730 71.676
R1199 B.n734 B.n733 71.676
R1200 B.n739 B.n738 71.676
R1201 B.n742 B.n741 71.676
R1202 B.n747 B.n746 71.676
R1203 B.n750 B.n749 71.676
R1204 B.n756 B.n755 71.676
R1205 B.n759 B.n758 71.676
R1206 B.n764 B.n763 71.676
R1207 B.n767 B.n766 71.676
R1208 B.n772 B.n771 71.676
R1209 B.n775 B.n774 71.676
R1210 B.n780 B.n779 71.676
R1211 B.n783 B.n782 71.676
R1212 B.n788 B.n787 71.676
R1213 B.n791 B.n790 71.676
R1214 B.n796 B.n795 71.676
R1215 B.n799 B.n798 71.676
R1216 B.n804 B.n803 71.676
R1217 B.n807 B.n806 71.676
R1218 B.n812 B.n811 71.676
R1219 B.n815 B.n814 71.676
R1220 B.n820 B.n819 71.676
R1221 B.n823 B.n822 71.676
R1222 B.n828 B.n827 71.676
R1223 B.n831 B.n830 71.676
R1224 B.n836 B.n835 71.676
R1225 B.n839 B.n838 71.676
R1226 B.n844 B.n843 71.676
R1227 B.n847 B.n846 71.676
R1228 B.n455 B.n454 71.676
R1229 B.n449 B.n239 71.676
R1230 B.n447 B.n446 71.676
R1231 B.n442 B.n441 71.676
R1232 B.n439 B.n438 71.676
R1233 B.n434 B.n433 71.676
R1234 B.n431 B.n430 71.676
R1235 B.n426 B.n425 71.676
R1236 B.n423 B.n422 71.676
R1237 B.n418 B.n417 71.676
R1238 B.n415 B.n414 71.676
R1239 B.n410 B.n409 71.676
R1240 B.n407 B.n406 71.676
R1241 B.n402 B.n401 71.676
R1242 B.n399 B.n398 71.676
R1243 B.n394 B.n393 71.676
R1244 B.n391 B.n390 71.676
R1245 B.n386 B.n385 71.676
R1246 B.n383 B.n382 71.676
R1247 B.n377 B.n376 71.676
R1248 B.n374 B.n373 71.676
R1249 B.n369 B.n368 71.676
R1250 B.n366 B.n365 71.676
R1251 B.n360 B.n359 71.676
R1252 B.n357 B.n356 71.676
R1253 B.n352 B.n351 71.676
R1254 B.n349 B.n348 71.676
R1255 B.n344 B.n343 71.676
R1256 B.n341 B.n340 71.676
R1257 B.n336 B.n335 71.676
R1258 B.n333 B.n332 71.676
R1259 B.n328 B.n327 71.676
R1260 B.n325 B.n324 71.676
R1261 B.n320 B.n319 71.676
R1262 B.n317 B.n316 71.676
R1263 B.n312 B.n311 71.676
R1264 B.n309 B.n308 71.676
R1265 B.n304 B.n303 71.676
R1266 B.n301 B.n300 71.676
R1267 B.n296 B.n295 71.676
R1268 B.n293 B.n292 71.676
R1269 B.n288 B.n287 71.676
R1270 B.n285 B.n235 71.676
R1271 B.n265 B.t10 71.2272
R1272 B.n122 B.t15 71.2272
R1273 B.n259 B.t20 71.2135
R1274 B.n115 B.t18 71.2135
R1275 B.n362 B.n265 59.5399
R1276 B.n380 B.n259 59.5399
R1277 B.n116 B.n115 59.5399
R1278 B.n753 B.n122 59.5399
R1279 B.n265 B.n264 55.4672
R1280 B.n259 B.n258 55.4672
R1281 B.n115 B.n114 55.4672
R1282 B.n122 B.n121 55.4672
R1283 B.n460 B.n232 45.8198
R1284 B.n466 B.n232 45.8198
R1285 B.n466 B.n228 45.8198
R1286 B.n472 B.n228 45.8198
R1287 B.n472 B.n224 45.8198
R1288 B.n479 B.n224 45.8198
R1289 B.n479 B.n478 45.8198
R1290 B.n485 B.n217 45.8198
R1291 B.n491 B.n217 45.8198
R1292 B.n491 B.n213 45.8198
R1293 B.n497 B.n213 45.8198
R1294 B.n497 B.n209 45.8198
R1295 B.n503 B.n209 45.8198
R1296 B.n503 B.n205 45.8198
R1297 B.n509 B.n205 45.8198
R1298 B.n509 B.n201 45.8198
R1299 B.n515 B.n201 45.8198
R1300 B.n521 B.n197 45.8198
R1301 B.n521 B.n193 45.8198
R1302 B.n527 B.n193 45.8198
R1303 B.n527 B.n189 45.8198
R1304 B.n533 B.n189 45.8198
R1305 B.n533 B.n185 45.8198
R1306 B.n540 B.n185 45.8198
R1307 B.n540 B.n539 45.8198
R1308 B.n546 B.n178 45.8198
R1309 B.n552 B.n178 45.8198
R1310 B.n552 B.n174 45.8198
R1311 B.n558 B.n174 45.8198
R1312 B.n558 B.n170 45.8198
R1313 B.n565 B.n170 45.8198
R1314 B.n565 B.n564 45.8198
R1315 B.n571 B.n163 45.8198
R1316 B.n577 B.n163 45.8198
R1317 B.n577 B.n159 45.8198
R1318 B.n583 B.n159 45.8198
R1319 B.n583 B.n155 45.8198
R1320 B.n589 B.n155 45.8198
R1321 B.n589 B.n151 45.8198
R1322 B.n595 B.n151 45.8198
R1323 B.n602 B.n147 45.8198
R1324 B.n602 B.n143 45.8198
R1325 B.n608 B.n143 45.8198
R1326 B.n608 B.n4 45.8198
R1327 B.n950 B.n4 45.8198
R1328 B.n950 B.n949 45.8198
R1329 B.n949 B.n948 45.8198
R1330 B.n948 B.n8 45.8198
R1331 B.n942 B.n8 45.8198
R1332 B.n942 B.n941 45.8198
R1333 B.n940 B.n15 45.8198
R1334 B.n934 B.n15 45.8198
R1335 B.n934 B.n933 45.8198
R1336 B.n933 B.n932 45.8198
R1337 B.n932 B.n22 45.8198
R1338 B.n926 B.n22 45.8198
R1339 B.n926 B.n925 45.8198
R1340 B.n925 B.n924 45.8198
R1341 B.n918 B.n32 45.8198
R1342 B.n918 B.n917 45.8198
R1343 B.n917 B.n916 45.8198
R1344 B.n916 B.n36 45.8198
R1345 B.n910 B.n36 45.8198
R1346 B.n910 B.n909 45.8198
R1347 B.n909 B.n908 45.8198
R1348 B.n902 B.n46 45.8198
R1349 B.n902 B.n901 45.8198
R1350 B.n901 B.n900 45.8198
R1351 B.n900 B.n50 45.8198
R1352 B.n894 B.n50 45.8198
R1353 B.n894 B.n893 45.8198
R1354 B.n893 B.n892 45.8198
R1355 B.n892 B.n57 45.8198
R1356 B.n886 B.n885 45.8198
R1357 B.n885 B.n884 45.8198
R1358 B.n884 B.n64 45.8198
R1359 B.n878 B.n64 45.8198
R1360 B.n878 B.n877 45.8198
R1361 B.n877 B.n876 45.8198
R1362 B.n876 B.n71 45.8198
R1363 B.n870 B.n71 45.8198
R1364 B.n870 B.n869 45.8198
R1365 B.n869 B.n868 45.8198
R1366 B.n862 B.n81 45.8198
R1367 B.n862 B.n861 45.8198
R1368 B.n861 B.n860 45.8198
R1369 B.n860 B.n85 45.8198
R1370 B.n854 B.n85 45.8198
R1371 B.n854 B.n853 45.8198
R1372 B.n853 B.n852 45.8198
R1373 B.n515 B.t3 43.7984
R1374 B.n886 B.t5 43.7984
R1375 B.t4 B.n147 37.0602
R1376 B.n941 B.t1 37.0602
R1377 B.n564 B.t0 35.7126
R1378 B.n32 B.t2 35.7126
R1379 B.n675 B.n674 35.4346
R1380 B.n850 B.n849 35.4346
R1381 B.n462 B.n234 35.4346
R1382 B.n458 B.n457 35.4346
R1383 B.n485 B.t9 30.3221
R1384 B.n868 B.t13 30.3221
R1385 B.n546 B.t6 28.9745
R1386 B.n908 B.t7 28.9745
R1387 B B.n952 18.0485
R1388 B.n539 B.t6 16.8458
R1389 B.n46 B.t7 16.8458
R1390 B.n478 B.t9 15.4982
R1391 B.n81 B.t13 15.4982
R1392 B.n849 B.n848 10.6151
R1393 B.n848 B.n94 10.6151
R1394 B.n842 B.n94 10.6151
R1395 B.n842 B.n841 10.6151
R1396 B.n841 B.n840 10.6151
R1397 B.n840 B.n96 10.6151
R1398 B.n834 B.n96 10.6151
R1399 B.n834 B.n833 10.6151
R1400 B.n833 B.n832 10.6151
R1401 B.n832 B.n98 10.6151
R1402 B.n826 B.n98 10.6151
R1403 B.n826 B.n825 10.6151
R1404 B.n825 B.n824 10.6151
R1405 B.n824 B.n100 10.6151
R1406 B.n818 B.n100 10.6151
R1407 B.n818 B.n817 10.6151
R1408 B.n817 B.n816 10.6151
R1409 B.n816 B.n102 10.6151
R1410 B.n810 B.n102 10.6151
R1411 B.n810 B.n809 10.6151
R1412 B.n809 B.n808 10.6151
R1413 B.n808 B.n104 10.6151
R1414 B.n802 B.n104 10.6151
R1415 B.n802 B.n801 10.6151
R1416 B.n801 B.n800 10.6151
R1417 B.n800 B.n106 10.6151
R1418 B.n794 B.n106 10.6151
R1419 B.n794 B.n793 10.6151
R1420 B.n793 B.n792 10.6151
R1421 B.n792 B.n108 10.6151
R1422 B.n786 B.n108 10.6151
R1423 B.n786 B.n785 10.6151
R1424 B.n785 B.n784 10.6151
R1425 B.n784 B.n110 10.6151
R1426 B.n778 B.n110 10.6151
R1427 B.n778 B.n777 10.6151
R1428 B.n777 B.n776 10.6151
R1429 B.n776 B.n112 10.6151
R1430 B.n770 B.n769 10.6151
R1431 B.n769 B.n768 10.6151
R1432 B.n768 B.n117 10.6151
R1433 B.n762 B.n117 10.6151
R1434 B.n762 B.n761 10.6151
R1435 B.n761 B.n760 10.6151
R1436 B.n760 B.n119 10.6151
R1437 B.n754 B.n119 10.6151
R1438 B.n752 B.n751 10.6151
R1439 B.n751 B.n123 10.6151
R1440 B.n745 B.n123 10.6151
R1441 B.n745 B.n744 10.6151
R1442 B.n744 B.n743 10.6151
R1443 B.n743 B.n125 10.6151
R1444 B.n737 B.n125 10.6151
R1445 B.n737 B.n736 10.6151
R1446 B.n736 B.n735 10.6151
R1447 B.n735 B.n127 10.6151
R1448 B.n729 B.n127 10.6151
R1449 B.n729 B.n728 10.6151
R1450 B.n728 B.n727 10.6151
R1451 B.n727 B.n129 10.6151
R1452 B.n721 B.n129 10.6151
R1453 B.n721 B.n720 10.6151
R1454 B.n720 B.n719 10.6151
R1455 B.n719 B.n131 10.6151
R1456 B.n713 B.n131 10.6151
R1457 B.n713 B.n712 10.6151
R1458 B.n712 B.n711 10.6151
R1459 B.n711 B.n133 10.6151
R1460 B.n705 B.n133 10.6151
R1461 B.n705 B.n704 10.6151
R1462 B.n704 B.n703 10.6151
R1463 B.n703 B.n135 10.6151
R1464 B.n697 B.n135 10.6151
R1465 B.n697 B.n696 10.6151
R1466 B.n696 B.n695 10.6151
R1467 B.n695 B.n137 10.6151
R1468 B.n689 B.n137 10.6151
R1469 B.n689 B.n688 10.6151
R1470 B.n688 B.n687 10.6151
R1471 B.n687 B.n139 10.6151
R1472 B.n681 B.n139 10.6151
R1473 B.n681 B.n680 10.6151
R1474 B.n680 B.n679 10.6151
R1475 B.n679 B.n675 10.6151
R1476 B.n463 B.n462 10.6151
R1477 B.n464 B.n463 10.6151
R1478 B.n464 B.n226 10.6151
R1479 B.n474 B.n226 10.6151
R1480 B.n475 B.n474 10.6151
R1481 B.n476 B.n475 10.6151
R1482 B.n476 B.n219 10.6151
R1483 B.n487 B.n219 10.6151
R1484 B.n488 B.n487 10.6151
R1485 B.n489 B.n488 10.6151
R1486 B.n489 B.n211 10.6151
R1487 B.n499 B.n211 10.6151
R1488 B.n500 B.n499 10.6151
R1489 B.n501 B.n500 10.6151
R1490 B.n501 B.n203 10.6151
R1491 B.n511 B.n203 10.6151
R1492 B.n512 B.n511 10.6151
R1493 B.n513 B.n512 10.6151
R1494 B.n513 B.n195 10.6151
R1495 B.n523 B.n195 10.6151
R1496 B.n524 B.n523 10.6151
R1497 B.n525 B.n524 10.6151
R1498 B.n525 B.n187 10.6151
R1499 B.n535 B.n187 10.6151
R1500 B.n536 B.n535 10.6151
R1501 B.n537 B.n536 10.6151
R1502 B.n537 B.n180 10.6151
R1503 B.n548 B.n180 10.6151
R1504 B.n549 B.n548 10.6151
R1505 B.n550 B.n549 10.6151
R1506 B.n550 B.n172 10.6151
R1507 B.n560 B.n172 10.6151
R1508 B.n561 B.n560 10.6151
R1509 B.n562 B.n561 10.6151
R1510 B.n562 B.n165 10.6151
R1511 B.n573 B.n165 10.6151
R1512 B.n574 B.n573 10.6151
R1513 B.n575 B.n574 10.6151
R1514 B.n575 B.n157 10.6151
R1515 B.n585 B.n157 10.6151
R1516 B.n586 B.n585 10.6151
R1517 B.n587 B.n586 10.6151
R1518 B.n587 B.n149 10.6151
R1519 B.n597 B.n149 10.6151
R1520 B.n598 B.n597 10.6151
R1521 B.n600 B.n598 10.6151
R1522 B.n600 B.n599 10.6151
R1523 B.n599 B.n141 10.6151
R1524 B.n611 B.n141 10.6151
R1525 B.n612 B.n611 10.6151
R1526 B.n613 B.n612 10.6151
R1527 B.n614 B.n613 10.6151
R1528 B.n616 B.n614 10.6151
R1529 B.n617 B.n616 10.6151
R1530 B.n618 B.n617 10.6151
R1531 B.n619 B.n618 10.6151
R1532 B.n621 B.n619 10.6151
R1533 B.n622 B.n621 10.6151
R1534 B.n623 B.n622 10.6151
R1535 B.n624 B.n623 10.6151
R1536 B.n626 B.n624 10.6151
R1537 B.n627 B.n626 10.6151
R1538 B.n628 B.n627 10.6151
R1539 B.n629 B.n628 10.6151
R1540 B.n631 B.n629 10.6151
R1541 B.n632 B.n631 10.6151
R1542 B.n633 B.n632 10.6151
R1543 B.n634 B.n633 10.6151
R1544 B.n636 B.n634 10.6151
R1545 B.n637 B.n636 10.6151
R1546 B.n638 B.n637 10.6151
R1547 B.n639 B.n638 10.6151
R1548 B.n641 B.n639 10.6151
R1549 B.n642 B.n641 10.6151
R1550 B.n643 B.n642 10.6151
R1551 B.n644 B.n643 10.6151
R1552 B.n646 B.n644 10.6151
R1553 B.n647 B.n646 10.6151
R1554 B.n648 B.n647 10.6151
R1555 B.n649 B.n648 10.6151
R1556 B.n651 B.n649 10.6151
R1557 B.n652 B.n651 10.6151
R1558 B.n653 B.n652 10.6151
R1559 B.n654 B.n653 10.6151
R1560 B.n656 B.n654 10.6151
R1561 B.n657 B.n656 10.6151
R1562 B.n658 B.n657 10.6151
R1563 B.n659 B.n658 10.6151
R1564 B.n661 B.n659 10.6151
R1565 B.n662 B.n661 10.6151
R1566 B.n663 B.n662 10.6151
R1567 B.n664 B.n663 10.6151
R1568 B.n666 B.n664 10.6151
R1569 B.n667 B.n666 10.6151
R1570 B.n668 B.n667 10.6151
R1571 B.n669 B.n668 10.6151
R1572 B.n671 B.n669 10.6151
R1573 B.n672 B.n671 10.6151
R1574 B.n673 B.n672 10.6151
R1575 B.n674 B.n673 10.6151
R1576 B.n457 B.n456 10.6151
R1577 B.n456 B.n238 10.6151
R1578 B.n451 B.n238 10.6151
R1579 B.n451 B.n450 10.6151
R1580 B.n450 B.n240 10.6151
R1581 B.n445 B.n240 10.6151
R1582 B.n445 B.n444 10.6151
R1583 B.n444 B.n443 10.6151
R1584 B.n443 B.n242 10.6151
R1585 B.n437 B.n242 10.6151
R1586 B.n437 B.n436 10.6151
R1587 B.n436 B.n435 10.6151
R1588 B.n435 B.n244 10.6151
R1589 B.n429 B.n244 10.6151
R1590 B.n429 B.n428 10.6151
R1591 B.n428 B.n427 10.6151
R1592 B.n427 B.n246 10.6151
R1593 B.n421 B.n246 10.6151
R1594 B.n421 B.n420 10.6151
R1595 B.n420 B.n419 10.6151
R1596 B.n419 B.n248 10.6151
R1597 B.n413 B.n248 10.6151
R1598 B.n413 B.n412 10.6151
R1599 B.n412 B.n411 10.6151
R1600 B.n411 B.n250 10.6151
R1601 B.n405 B.n250 10.6151
R1602 B.n405 B.n404 10.6151
R1603 B.n404 B.n403 10.6151
R1604 B.n403 B.n252 10.6151
R1605 B.n397 B.n252 10.6151
R1606 B.n397 B.n396 10.6151
R1607 B.n396 B.n395 10.6151
R1608 B.n395 B.n254 10.6151
R1609 B.n389 B.n254 10.6151
R1610 B.n389 B.n388 10.6151
R1611 B.n388 B.n387 10.6151
R1612 B.n387 B.n256 10.6151
R1613 B.n381 B.n256 10.6151
R1614 B.n379 B.n378 10.6151
R1615 B.n378 B.n260 10.6151
R1616 B.n372 B.n260 10.6151
R1617 B.n372 B.n371 10.6151
R1618 B.n371 B.n370 10.6151
R1619 B.n370 B.n262 10.6151
R1620 B.n364 B.n262 10.6151
R1621 B.n364 B.n363 10.6151
R1622 B.n361 B.n266 10.6151
R1623 B.n355 B.n266 10.6151
R1624 B.n355 B.n354 10.6151
R1625 B.n354 B.n353 10.6151
R1626 B.n353 B.n268 10.6151
R1627 B.n347 B.n268 10.6151
R1628 B.n347 B.n346 10.6151
R1629 B.n346 B.n345 10.6151
R1630 B.n345 B.n270 10.6151
R1631 B.n339 B.n270 10.6151
R1632 B.n339 B.n338 10.6151
R1633 B.n338 B.n337 10.6151
R1634 B.n337 B.n272 10.6151
R1635 B.n331 B.n272 10.6151
R1636 B.n331 B.n330 10.6151
R1637 B.n330 B.n329 10.6151
R1638 B.n329 B.n274 10.6151
R1639 B.n323 B.n274 10.6151
R1640 B.n323 B.n322 10.6151
R1641 B.n322 B.n321 10.6151
R1642 B.n321 B.n276 10.6151
R1643 B.n315 B.n276 10.6151
R1644 B.n315 B.n314 10.6151
R1645 B.n314 B.n313 10.6151
R1646 B.n313 B.n278 10.6151
R1647 B.n307 B.n278 10.6151
R1648 B.n307 B.n306 10.6151
R1649 B.n306 B.n305 10.6151
R1650 B.n305 B.n280 10.6151
R1651 B.n299 B.n280 10.6151
R1652 B.n299 B.n298 10.6151
R1653 B.n298 B.n297 10.6151
R1654 B.n297 B.n282 10.6151
R1655 B.n291 B.n282 10.6151
R1656 B.n291 B.n290 10.6151
R1657 B.n290 B.n289 10.6151
R1658 B.n289 B.n284 10.6151
R1659 B.n284 B.n234 10.6151
R1660 B.n458 B.n230 10.6151
R1661 B.n468 B.n230 10.6151
R1662 B.n469 B.n468 10.6151
R1663 B.n470 B.n469 10.6151
R1664 B.n470 B.n222 10.6151
R1665 B.n481 B.n222 10.6151
R1666 B.n482 B.n481 10.6151
R1667 B.n483 B.n482 10.6151
R1668 B.n483 B.n215 10.6151
R1669 B.n493 B.n215 10.6151
R1670 B.n494 B.n493 10.6151
R1671 B.n495 B.n494 10.6151
R1672 B.n495 B.n207 10.6151
R1673 B.n505 B.n207 10.6151
R1674 B.n506 B.n505 10.6151
R1675 B.n507 B.n506 10.6151
R1676 B.n507 B.n199 10.6151
R1677 B.n517 B.n199 10.6151
R1678 B.n518 B.n517 10.6151
R1679 B.n519 B.n518 10.6151
R1680 B.n519 B.n191 10.6151
R1681 B.n529 B.n191 10.6151
R1682 B.n530 B.n529 10.6151
R1683 B.n531 B.n530 10.6151
R1684 B.n531 B.n183 10.6151
R1685 B.n542 B.n183 10.6151
R1686 B.n543 B.n542 10.6151
R1687 B.n544 B.n543 10.6151
R1688 B.n544 B.n176 10.6151
R1689 B.n554 B.n176 10.6151
R1690 B.n555 B.n554 10.6151
R1691 B.n556 B.n555 10.6151
R1692 B.n556 B.n168 10.6151
R1693 B.n567 B.n168 10.6151
R1694 B.n568 B.n567 10.6151
R1695 B.n569 B.n568 10.6151
R1696 B.n569 B.n161 10.6151
R1697 B.n579 B.n161 10.6151
R1698 B.n580 B.n579 10.6151
R1699 B.n581 B.n580 10.6151
R1700 B.n581 B.n153 10.6151
R1701 B.n591 B.n153 10.6151
R1702 B.n592 B.n591 10.6151
R1703 B.n593 B.n592 10.6151
R1704 B.n593 B.n145 10.6151
R1705 B.n604 B.n145 10.6151
R1706 B.n605 B.n604 10.6151
R1707 B.n606 B.n605 10.6151
R1708 B.n606 B.n0 10.6151
R1709 B.n946 B.n1 10.6151
R1710 B.n946 B.n945 10.6151
R1711 B.n945 B.n944 10.6151
R1712 B.n944 B.n10 10.6151
R1713 B.n938 B.n10 10.6151
R1714 B.n938 B.n937 10.6151
R1715 B.n937 B.n936 10.6151
R1716 B.n936 B.n17 10.6151
R1717 B.n930 B.n17 10.6151
R1718 B.n930 B.n929 10.6151
R1719 B.n929 B.n928 10.6151
R1720 B.n928 B.n24 10.6151
R1721 B.n922 B.n24 10.6151
R1722 B.n922 B.n921 10.6151
R1723 B.n921 B.n920 10.6151
R1724 B.n920 B.n30 10.6151
R1725 B.n914 B.n30 10.6151
R1726 B.n914 B.n913 10.6151
R1727 B.n913 B.n912 10.6151
R1728 B.n912 B.n38 10.6151
R1729 B.n906 B.n38 10.6151
R1730 B.n906 B.n905 10.6151
R1731 B.n905 B.n904 10.6151
R1732 B.n904 B.n44 10.6151
R1733 B.n898 B.n44 10.6151
R1734 B.n898 B.n897 10.6151
R1735 B.n897 B.n896 10.6151
R1736 B.n896 B.n52 10.6151
R1737 B.n890 B.n52 10.6151
R1738 B.n890 B.n889 10.6151
R1739 B.n889 B.n888 10.6151
R1740 B.n888 B.n59 10.6151
R1741 B.n882 B.n59 10.6151
R1742 B.n882 B.n881 10.6151
R1743 B.n881 B.n880 10.6151
R1744 B.n880 B.n66 10.6151
R1745 B.n874 B.n66 10.6151
R1746 B.n874 B.n873 10.6151
R1747 B.n873 B.n872 10.6151
R1748 B.n872 B.n73 10.6151
R1749 B.n866 B.n73 10.6151
R1750 B.n866 B.n865 10.6151
R1751 B.n865 B.n864 10.6151
R1752 B.n864 B.n79 10.6151
R1753 B.n858 B.n79 10.6151
R1754 B.n858 B.n857 10.6151
R1755 B.n857 B.n856 10.6151
R1756 B.n856 B.n87 10.6151
R1757 B.n850 B.n87 10.6151
R1758 B.n571 B.t0 10.1077
R1759 B.n924 B.t2 10.1077
R1760 B.n595 B.t4 8.76007
R1761 B.t1 B.n940 8.76007
R1762 B.n770 B.n116 6.5566
R1763 B.n754 B.n753 6.5566
R1764 B.n380 B.n379 6.5566
R1765 B.n363 B.n362 6.5566
R1766 B.n116 B.n112 4.05904
R1767 B.n753 B.n752 4.05904
R1768 B.n381 B.n380 4.05904
R1769 B.n362 B.n361 4.05904
R1770 B.n952 B.n0 2.81026
R1771 B.n952 B.n1 2.81026
R1772 B.t3 B.n197 2.02194
R1773 B.t5 B.n57 2.02194
R1774 VP.n19 VP.n18 161.3
R1775 VP.n20 VP.n15 161.3
R1776 VP.n22 VP.n21 161.3
R1777 VP.n23 VP.n14 161.3
R1778 VP.n25 VP.n24 161.3
R1779 VP.n27 VP.n26 161.3
R1780 VP.n28 VP.n12 161.3
R1781 VP.n30 VP.n29 161.3
R1782 VP.n31 VP.n11 161.3
R1783 VP.n33 VP.n32 161.3
R1784 VP.n34 VP.n10 161.3
R1785 VP.n64 VP.n0 161.3
R1786 VP.n63 VP.n62 161.3
R1787 VP.n61 VP.n1 161.3
R1788 VP.n60 VP.n59 161.3
R1789 VP.n58 VP.n2 161.3
R1790 VP.n57 VP.n56 161.3
R1791 VP.n55 VP.n54 161.3
R1792 VP.n53 VP.n4 161.3
R1793 VP.n52 VP.n51 161.3
R1794 VP.n50 VP.n5 161.3
R1795 VP.n49 VP.n48 161.3
R1796 VP.n46 VP.n6 161.3
R1797 VP.n45 VP.n44 161.3
R1798 VP.n43 VP.n7 161.3
R1799 VP.n42 VP.n41 161.3
R1800 VP.n40 VP.n8 161.3
R1801 VP.n39 VP.n38 161.3
R1802 VP.n16 VP.t0 140.048
R1803 VP.n9 VP.t1 105.26
R1804 VP.n47 VP.t6 105.26
R1805 VP.n3 VP.t5 105.26
R1806 VP.n65 VP.t7 105.26
R1807 VP.n35 VP.t4 105.26
R1808 VP.n13 VP.t3 105.26
R1809 VP.n17 VP.t2 105.26
R1810 VP.n37 VP.n9 96.5656
R1811 VP.n66 VP.n65 96.5656
R1812 VP.n36 VP.n35 96.5656
R1813 VP.n41 VP.n7 54.0911
R1814 VP.n59 VP.n1 54.0911
R1815 VP.n29 VP.n11 54.0911
R1816 VP.n17 VP.n16 51.6001
R1817 VP.n37 VP.n36 49.9163
R1818 VP.n52 VP.n5 40.4934
R1819 VP.n53 VP.n52 40.4934
R1820 VP.n23 VP.n22 40.4934
R1821 VP.n22 VP.n15 40.4934
R1822 VP.n41 VP.n40 26.8957
R1823 VP.n63 VP.n1 26.8957
R1824 VP.n33 VP.n11 26.8957
R1825 VP.n40 VP.n39 24.4675
R1826 VP.n45 VP.n7 24.4675
R1827 VP.n46 VP.n45 24.4675
R1828 VP.n48 VP.n5 24.4675
R1829 VP.n54 VP.n53 24.4675
R1830 VP.n58 VP.n57 24.4675
R1831 VP.n59 VP.n58 24.4675
R1832 VP.n64 VP.n63 24.4675
R1833 VP.n34 VP.n33 24.4675
R1834 VP.n24 VP.n23 24.4675
R1835 VP.n28 VP.n27 24.4675
R1836 VP.n29 VP.n28 24.4675
R1837 VP.n18 VP.n15 24.4675
R1838 VP.n48 VP.n47 21.0421
R1839 VP.n54 VP.n3 21.0421
R1840 VP.n24 VP.n13 21.0421
R1841 VP.n18 VP.n17 21.0421
R1842 VP.n39 VP.n9 14.1914
R1843 VP.n65 VP.n64 14.1914
R1844 VP.n35 VP.n34 14.1914
R1845 VP.n19 VP.n16 6.57419
R1846 VP.n47 VP.n46 3.42588
R1847 VP.n57 VP.n3 3.42588
R1848 VP.n27 VP.n13 3.42588
R1849 VP.n36 VP.n10 0.278367
R1850 VP.n38 VP.n37 0.278367
R1851 VP.n66 VP.n0 0.278367
R1852 VP.n20 VP.n19 0.189894
R1853 VP.n21 VP.n20 0.189894
R1854 VP.n21 VP.n14 0.189894
R1855 VP.n25 VP.n14 0.189894
R1856 VP.n26 VP.n25 0.189894
R1857 VP.n26 VP.n12 0.189894
R1858 VP.n30 VP.n12 0.189894
R1859 VP.n31 VP.n30 0.189894
R1860 VP.n32 VP.n31 0.189894
R1861 VP.n32 VP.n10 0.189894
R1862 VP.n38 VP.n8 0.189894
R1863 VP.n42 VP.n8 0.189894
R1864 VP.n43 VP.n42 0.189894
R1865 VP.n44 VP.n43 0.189894
R1866 VP.n44 VP.n6 0.189894
R1867 VP.n49 VP.n6 0.189894
R1868 VP.n50 VP.n49 0.189894
R1869 VP.n51 VP.n50 0.189894
R1870 VP.n51 VP.n4 0.189894
R1871 VP.n55 VP.n4 0.189894
R1872 VP.n56 VP.n55 0.189894
R1873 VP.n56 VP.n2 0.189894
R1874 VP.n60 VP.n2 0.189894
R1875 VP.n61 VP.n60 0.189894
R1876 VP.n62 VP.n61 0.189894
R1877 VP.n62 VP.n0 0.189894
R1878 VP VP.n66 0.153454
R1879 VDD1 VDD1.n0 63.694
R1880 VDD1.n3 VDD1.n2 63.5803
R1881 VDD1.n3 VDD1.n1 63.5803
R1882 VDD1.n5 VDD1.n4 62.4029
R1883 VDD1.n5 VDD1.n3 44.919
R1884 VDD1.n4 VDD1.t4 1.79236
R1885 VDD1.n4 VDD1.t3 1.79236
R1886 VDD1.n0 VDD1.t7 1.79236
R1887 VDD1.n0 VDD1.t5 1.79236
R1888 VDD1.n2 VDD1.t2 1.79236
R1889 VDD1.n2 VDD1.t0 1.79236
R1890 VDD1.n1 VDD1.t6 1.79236
R1891 VDD1.n1 VDD1.t1 1.79236
R1892 VDD1 VDD1.n5 1.17507
C0 VN VDD1 0.151599f
C1 VDD2 VTAIL 7.79626f
C2 VDD2 VP 0.512219f
C3 VDD2 VN 7.99455f
C4 VTAIL VP 8.42925f
C5 VDD2 VDD1 1.74091f
C6 VTAIL VN 8.415151f
C7 VN VP 7.39811f
C8 VTAIL VDD1 7.74232f
C9 VDD1 VP 8.35381f
C10 VDD2 B 5.205862f
C11 VDD1 B 5.635907f
C12 VTAIL B 9.864717f
C13 VN B 15.15201f
C14 VP B 13.745961f
C15 VDD1.t7 B 0.215143f
C16 VDD1.t5 B 0.215143f
C17 VDD1.n0 B 1.91765f
C18 VDD1.t6 B 0.215143f
C19 VDD1.t1 B 0.215143f
C20 VDD1.n1 B 1.91659f
C21 VDD1.t2 B 0.215143f
C22 VDD1.t0 B 0.215143f
C23 VDD1.n2 B 1.91659f
C24 VDD1.n3 B 3.18287f
C25 VDD1.t4 B 0.215143f
C26 VDD1.t3 B 0.215143f
C27 VDD1.n4 B 1.90729f
C28 VDD1.n5 B 2.84182f
C29 VP.n0 B 0.030561f
C30 VP.t7 B 1.76133f
C31 VP.n1 B 0.025316f
C32 VP.n2 B 0.02318f
C33 VP.t5 B 1.76133f
C34 VP.n3 B 0.626702f
C35 VP.n4 B 0.02318f
C36 VP.n5 B 0.046071f
C37 VP.n6 B 0.02318f
C38 VP.t6 B 1.76133f
C39 VP.n7 B 0.040631f
C40 VP.n8 B 0.02318f
C41 VP.t1 B 1.76133f
C42 VP.n9 B 0.707963f
C43 VP.n10 B 0.030561f
C44 VP.t4 B 1.76133f
C45 VP.n11 B 0.025316f
C46 VP.n12 B 0.02318f
C47 VP.t3 B 1.76133f
C48 VP.n13 B 0.626702f
C49 VP.n14 B 0.02318f
C50 VP.n15 B 0.046071f
C51 VP.t0 B 1.95278f
C52 VP.n16 B 0.669083f
C53 VP.t2 B 1.76133f
C54 VP.n17 B 0.701206f
C55 VP.n18 B 0.040216f
C56 VP.n19 B 0.222254f
C57 VP.n20 B 0.02318f
C58 VP.n21 B 0.02318f
C59 VP.n22 B 0.018739f
C60 VP.n23 B 0.046071f
C61 VP.n24 B 0.040216f
C62 VP.n25 B 0.02318f
C63 VP.n26 B 0.02318f
C64 VP.n27 B 0.024859f
C65 VP.n28 B 0.043202f
C66 VP.n29 B 0.040631f
C67 VP.n30 B 0.02318f
C68 VP.n31 B 0.02318f
C69 VP.n32 B 0.02318f
C70 VP.n33 B 0.044934f
C71 VP.n34 B 0.034244f
C72 VP.n35 B 0.707963f
C73 VP.n36 B 1.28398f
C74 VP.n37 B 1.30067f
C75 VP.n38 B 0.030561f
C76 VP.n39 B 0.034244f
C77 VP.n40 B 0.044934f
C78 VP.n41 B 0.025316f
C79 VP.n42 B 0.02318f
C80 VP.n43 B 0.02318f
C81 VP.n44 B 0.02318f
C82 VP.n45 B 0.043202f
C83 VP.n46 B 0.024859f
C84 VP.n47 B 0.626702f
C85 VP.n48 B 0.040216f
C86 VP.n49 B 0.02318f
C87 VP.n50 B 0.02318f
C88 VP.n51 B 0.02318f
C89 VP.n52 B 0.018739f
C90 VP.n53 B 0.046071f
C91 VP.n54 B 0.040216f
C92 VP.n55 B 0.02318f
C93 VP.n56 B 0.02318f
C94 VP.n57 B 0.024859f
C95 VP.n58 B 0.043202f
C96 VP.n59 B 0.040631f
C97 VP.n60 B 0.02318f
C98 VP.n61 B 0.02318f
C99 VP.n62 B 0.02318f
C100 VP.n63 B 0.044934f
C101 VP.n64 B 0.034244f
C102 VP.n65 B 0.707963f
C103 VP.n66 B 0.034531f
C104 VDD2.t0 B 0.212334f
C105 VDD2.t3 B 0.212334f
C106 VDD2.n0 B 1.89157f
C107 VDD2.t4 B 0.212334f
C108 VDD2.t7 B 0.212334f
C109 VDD2.n1 B 1.89157f
C110 VDD2.n2 B 3.0906f
C111 VDD2.t5 B 0.212334f
C112 VDD2.t6 B 0.212334f
C113 VDD2.n3 B 1.8824f
C114 VDD2.n4 B 2.77473f
C115 VDD2.t1 B 0.212334f
C116 VDD2.t2 B 0.212334f
C117 VDD2.n5 B 1.89153f
C118 VTAIL.t8 B 0.174782f
C119 VTAIL.t9 B 0.174782f
C120 VTAIL.n0 B 1.49086f
C121 VTAIL.n1 B 0.35871f
C122 VTAIL.t13 B 1.89993f
C123 VTAIL.n2 B 0.45287f
C124 VTAIL.t4 B 1.89993f
C125 VTAIL.n3 B 0.45287f
C126 VTAIL.t6 B 0.174782f
C127 VTAIL.t0 B 0.174782f
C128 VTAIL.n4 B 1.49086f
C129 VTAIL.n5 B 0.513975f
C130 VTAIL.t3 B 1.89993f
C131 VTAIL.n6 B 1.46787f
C132 VTAIL.t11 B 1.89994f
C133 VTAIL.n7 B 1.46785f
C134 VTAIL.t12 B 0.174782f
C135 VTAIL.t15 B 0.174782f
C136 VTAIL.n8 B 1.49087f
C137 VTAIL.n9 B 0.51397f
C138 VTAIL.t10 B 1.89994f
C139 VTAIL.n10 B 0.452858f
C140 VTAIL.t1 B 1.89994f
C141 VTAIL.n11 B 0.452858f
C142 VTAIL.t2 B 0.174782f
C143 VTAIL.t7 B 0.174782f
C144 VTAIL.n12 B 1.49087f
C145 VTAIL.n13 B 0.51397f
C146 VTAIL.t5 B 1.89993f
C147 VTAIL.n14 B 1.46787f
C148 VTAIL.t14 B 1.89993f
C149 VTAIL.n15 B 1.46411f
C150 VN.n0 B 0.030015f
C151 VN.t0 B 1.72989f
C152 VN.n1 B 0.024864f
C153 VN.n2 B 0.022767f
C154 VN.t3 B 1.72989f
C155 VN.n3 B 0.615515f
C156 VN.n4 B 0.022767f
C157 VN.n5 B 0.045248f
C158 VN.t7 B 1.91792f
C159 VN.n6 B 0.657139f
C160 VN.t4 B 1.72989f
C161 VN.n7 B 0.688689f
C162 VN.n8 B 0.039498f
C163 VN.n9 B 0.218287f
C164 VN.n10 B 0.022767f
C165 VN.n11 B 0.022767f
C166 VN.n12 B 0.018405f
C167 VN.n13 B 0.045248f
C168 VN.n14 B 0.039498f
C169 VN.n15 B 0.022767f
C170 VN.n16 B 0.022767f
C171 VN.n17 B 0.024416f
C172 VN.n18 B 0.042431f
C173 VN.n19 B 0.039905f
C174 VN.n20 B 0.022767f
C175 VN.n21 B 0.022767f
C176 VN.n22 B 0.022767f
C177 VN.n23 B 0.044132f
C178 VN.n24 B 0.033633f
C179 VN.n25 B 0.695325f
C180 VN.n26 B 0.033915f
C181 VN.n27 B 0.030015f
C182 VN.t2 B 1.72989f
C183 VN.n28 B 0.024864f
C184 VN.n29 B 0.022767f
C185 VN.t1 B 1.72989f
C186 VN.n30 B 0.615515f
C187 VN.n31 B 0.022767f
C188 VN.n32 B 0.045248f
C189 VN.t5 B 1.91792f
C190 VN.n33 B 0.657139f
C191 VN.t6 B 1.72989f
C192 VN.n34 B 0.688689f
C193 VN.n35 B 0.039498f
C194 VN.n36 B 0.218287f
C195 VN.n37 B 0.022767f
C196 VN.n38 B 0.022767f
C197 VN.n39 B 0.018405f
C198 VN.n40 B 0.045248f
C199 VN.n41 B 0.039498f
C200 VN.n42 B 0.022767f
C201 VN.n43 B 0.022767f
C202 VN.n44 B 0.024416f
C203 VN.n45 B 0.042431f
C204 VN.n46 B 0.039905f
C205 VN.n47 B 0.022767f
C206 VN.n48 B 0.022767f
C207 VN.n49 B 0.022767f
C208 VN.n50 B 0.044132f
C209 VN.n51 B 0.033633f
C210 VN.n52 B 0.695325f
C211 VN.n53 B 1.27329f
.ends

