* NGSPICE file created from diff_pair_sample_0483.ext - technology: sky130A

.subckt diff_pair_sample_0483 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t2 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X1 VDD2.t9 VN.t0 VTAIL.t18 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X2 VDD1.t4 VP.t1 VTAIL.t14 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X3 B.t11 B.t9 B.t10 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0 ps=0 w=2.62 l=3.65
X4 VTAIL.t2 VN.t1 VDD2.t8 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X5 VDD1.t0 VP.t2 VTAIL.t13 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=1.0218 ps=6.02 w=2.62 l=3.65
X6 VDD1.t7 VP.t3 VTAIL.t12 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=1.0218 ps=6.02 w=2.62 l=3.65
X7 VTAIL.t11 VP.t4 VDD1.t6 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X8 VTAIL.t4 VN.t2 VDD2.t7 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X9 VDD2.t6 VN.t3 VTAIL.t16 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X10 VDD2.t5 VN.t4 VTAIL.t5 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=1.0218 ps=6.02 w=2.62 l=3.65
X11 VDD1.t9 VP.t5 VTAIL.t10 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0.4323 ps=2.95 w=2.62 l=3.65
X12 B.t8 B.t6 B.t7 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0 ps=0 w=2.62 l=3.65
X13 VTAIL.t9 VP.t6 VDD1.t8 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X14 B.t5 B.t3 B.t4 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0 ps=0 w=2.62 l=3.65
X15 VTAIL.t8 VP.t7 VDD1.t3 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X16 VDD2.t4 VN.t5 VTAIL.t1 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0.4323 ps=2.95 w=2.62 l=3.65
X17 VDD2.t3 VN.t6 VTAIL.t19 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=1.0218 ps=6.02 w=2.62 l=3.65
X18 VTAIL.t0 VN.t7 VDD2.t2 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X19 VDD1.t5 VP.t8 VTAIL.t7 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0.4323 ps=2.95 w=2.62 l=3.65
X20 VDD2.t1 VN.t8 VTAIL.t3 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0.4323 ps=2.95 w=2.62 l=3.65
X21 B.t2 B.t0 B.t1 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=1.0218 pd=6.02 as=0 ps=0 w=2.62 l=3.65
X22 VDD1.t1 VP.t9 VTAIL.t6 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
X23 VTAIL.t17 VN.t9 VDD2.t0 w_n5746_n1492# sky130_fd_pr__pfet_01v8 ad=0.4323 pd=2.95 as=0.4323 ps=2.95 w=2.62 l=3.65
R0 VP.n32 VP.n29 161.3
R1 VP.n34 VP.n33 161.3
R2 VP.n35 VP.n28 161.3
R3 VP.n37 VP.n36 161.3
R4 VP.n38 VP.n27 161.3
R5 VP.n40 VP.n39 161.3
R6 VP.n41 VP.n26 161.3
R7 VP.n44 VP.n43 161.3
R8 VP.n45 VP.n25 161.3
R9 VP.n47 VP.n46 161.3
R10 VP.n48 VP.n24 161.3
R11 VP.n50 VP.n49 161.3
R12 VP.n51 VP.n23 161.3
R13 VP.n53 VP.n52 161.3
R14 VP.n54 VP.n22 161.3
R15 VP.n57 VP.n56 161.3
R16 VP.n58 VP.n21 161.3
R17 VP.n60 VP.n59 161.3
R18 VP.n61 VP.n20 161.3
R19 VP.n63 VP.n62 161.3
R20 VP.n64 VP.n19 161.3
R21 VP.n66 VP.n65 161.3
R22 VP.n67 VP.n18 161.3
R23 VP.n69 VP.n68 161.3
R24 VP.n123 VP.n122 161.3
R25 VP.n121 VP.n1 161.3
R26 VP.n120 VP.n119 161.3
R27 VP.n118 VP.n2 161.3
R28 VP.n117 VP.n116 161.3
R29 VP.n115 VP.n3 161.3
R30 VP.n114 VP.n113 161.3
R31 VP.n112 VP.n4 161.3
R32 VP.n111 VP.n110 161.3
R33 VP.n108 VP.n5 161.3
R34 VP.n107 VP.n106 161.3
R35 VP.n105 VP.n6 161.3
R36 VP.n104 VP.n103 161.3
R37 VP.n102 VP.n7 161.3
R38 VP.n101 VP.n100 161.3
R39 VP.n99 VP.n8 161.3
R40 VP.n98 VP.n97 161.3
R41 VP.n95 VP.n9 161.3
R42 VP.n94 VP.n93 161.3
R43 VP.n92 VP.n10 161.3
R44 VP.n91 VP.n90 161.3
R45 VP.n89 VP.n11 161.3
R46 VP.n88 VP.n87 161.3
R47 VP.n86 VP.n12 161.3
R48 VP.n85 VP.n84 161.3
R49 VP.n82 VP.n13 161.3
R50 VP.n81 VP.n80 161.3
R51 VP.n79 VP.n14 161.3
R52 VP.n78 VP.n77 161.3
R53 VP.n76 VP.n15 161.3
R54 VP.n75 VP.n74 161.3
R55 VP.n73 VP.n16 161.3
R56 VP.n72 VP.n71 79.917
R57 VP.n124 VP.n0 79.917
R58 VP.n70 VP.n17 79.917
R59 VP.n31 VP.n30 63.5339
R60 VP.n103 VP.n6 56.5617
R61 VP.n36 VP.n27 56.5617
R62 VP.n77 VP.n14 56.5617
R63 VP.n90 VP.n10 56.5617
R64 VP.n116 VP.n2 56.5617
R65 VP.n62 VP.n19 56.5617
R66 VP.n49 VP.n23 56.5617
R67 VP.n72 VP.n70 51.848
R68 VP.n31 VP.t5 50.8209
R69 VP.n75 VP.n16 24.5923
R70 VP.n76 VP.n75 24.5923
R71 VP.n77 VP.n76 24.5923
R72 VP.n81 VP.n14 24.5923
R73 VP.n82 VP.n81 24.5923
R74 VP.n84 VP.n82 24.5923
R75 VP.n88 VP.n12 24.5923
R76 VP.n89 VP.n88 24.5923
R77 VP.n90 VP.n89 24.5923
R78 VP.n94 VP.n10 24.5923
R79 VP.n95 VP.n94 24.5923
R80 VP.n97 VP.n95 24.5923
R81 VP.n101 VP.n8 24.5923
R82 VP.n102 VP.n101 24.5923
R83 VP.n103 VP.n102 24.5923
R84 VP.n107 VP.n6 24.5923
R85 VP.n108 VP.n107 24.5923
R86 VP.n110 VP.n108 24.5923
R87 VP.n114 VP.n4 24.5923
R88 VP.n115 VP.n114 24.5923
R89 VP.n116 VP.n115 24.5923
R90 VP.n120 VP.n2 24.5923
R91 VP.n121 VP.n120 24.5923
R92 VP.n122 VP.n121 24.5923
R93 VP.n66 VP.n19 24.5923
R94 VP.n67 VP.n66 24.5923
R95 VP.n68 VP.n67 24.5923
R96 VP.n53 VP.n23 24.5923
R97 VP.n54 VP.n53 24.5923
R98 VP.n56 VP.n54 24.5923
R99 VP.n60 VP.n21 24.5923
R100 VP.n61 VP.n60 24.5923
R101 VP.n62 VP.n61 24.5923
R102 VP.n40 VP.n27 24.5923
R103 VP.n41 VP.n40 24.5923
R104 VP.n43 VP.n41 24.5923
R105 VP.n47 VP.n25 24.5923
R106 VP.n48 VP.n47 24.5923
R107 VP.n49 VP.n48 24.5923
R108 VP.n34 VP.n29 24.5923
R109 VP.n35 VP.n34 24.5923
R110 VP.n36 VP.n35 24.5923
R111 VP.n71 VP.t8 17.2997
R112 VP.n83 VP.t6 17.2997
R113 VP.n96 VP.t1 17.2997
R114 VP.n109 VP.t0 17.2997
R115 VP.n0 VP.t2 17.2997
R116 VP.n17 VP.t3 17.2997
R117 VP.n55 VP.t7 17.2997
R118 VP.n42 VP.t9 17.2997
R119 VP.n30 VP.t4 17.2997
R120 VP.n84 VP.n83 13.2801
R121 VP.n109 VP.n4 13.2801
R122 VP.n55 VP.n21 13.2801
R123 VP.n97 VP.n96 12.2964
R124 VP.n96 VP.n8 12.2964
R125 VP.n43 VP.n42 12.2964
R126 VP.n42 VP.n25 12.2964
R127 VP.n83 VP.n12 11.3127
R128 VP.n110 VP.n109 11.3127
R129 VP.n56 VP.n55 11.3127
R130 VP.n30 VP.n29 11.3127
R131 VP.n71 VP.n16 10.3291
R132 VP.n122 VP.n0 10.3291
R133 VP.n68 VP.n17 10.3291
R134 VP.n32 VP.n31 3.13517
R135 VP.n70 VP.n69 0.354861
R136 VP.n73 VP.n72 0.354861
R137 VP.n124 VP.n123 0.354861
R138 VP VP.n124 0.267071
R139 VP.n33 VP.n32 0.189894
R140 VP.n33 VP.n28 0.189894
R141 VP.n37 VP.n28 0.189894
R142 VP.n38 VP.n37 0.189894
R143 VP.n39 VP.n38 0.189894
R144 VP.n39 VP.n26 0.189894
R145 VP.n44 VP.n26 0.189894
R146 VP.n45 VP.n44 0.189894
R147 VP.n46 VP.n45 0.189894
R148 VP.n46 VP.n24 0.189894
R149 VP.n50 VP.n24 0.189894
R150 VP.n51 VP.n50 0.189894
R151 VP.n52 VP.n51 0.189894
R152 VP.n52 VP.n22 0.189894
R153 VP.n57 VP.n22 0.189894
R154 VP.n58 VP.n57 0.189894
R155 VP.n59 VP.n58 0.189894
R156 VP.n59 VP.n20 0.189894
R157 VP.n63 VP.n20 0.189894
R158 VP.n64 VP.n63 0.189894
R159 VP.n65 VP.n64 0.189894
R160 VP.n65 VP.n18 0.189894
R161 VP.n69 VP.n18 0.189894
R162 VP.n74 VP.n73 0.189894
R163 VP.n74 VP.n15 0.189894
R164 VP.n78 VP.n15 0.189894
R165 VP.n79 VP.n78 0.189894
R166 VP.n80 VP.n79 0.189894
R167 VP.n80 VP.n13 0.189894
R168 VP.n85 VP.n13 0.189894
R169 VP.n86 VP.n85 0.189894
R170 VP.n87 VP.n86 0.189894
R171 VP.n87 VP.n11 0.189894
R172 VP.n91 VP.n11 0.189894
R173 VP.n92 VP.n91 0.189894
R174 VP.n93 VP.n92 0.189894
R175 VP.n93 VP.n9 0.189894
R176 VP.n98 VP.n9 0.189894
R177 VP.n99 VP.n98 0.189894
R178 VP.n100 VP.n99 0.189894
R179 VP.n100 VP.n7 0.189894
R180 VP.n104 VP.n7 0.189894
R181 VP.n105 VP.n104 0.189894
R182 VP.n106 VP.n105 0.189894
R183 VP.n106 VP.n5 0.189894
R184 VP.n111 VP.n5 0.189894
R185 VP.n112 VP.n111 0.189894
R186 VP.n113 VP.n112 0.189894
R187 VP.n113 VP.n3 0.189894
R188 VP.n117 VP.n3 0.189894
R189 VP.n118 VP.n117 0.189894
R190 VP.n119 VP.n118 0.189894
R191 VP.n119 VP.n1 0.189894
R192 VP.n123 VP.n1 0.189894
R193 VDD1.n6 VDD1.n0 756.745
R194 VDD1.n19 VDD1.n13 756.745
R195 VDD1.n7 VDD1.n6 585
R196 VDD1.n5 VDD1.n4 585
R197 VDD1.n18 VDD1.n17 585
R198 VDD1.n20 VDD1.n19 585
R199 VDD1.n3 VDD1.t9 355.474
R200 VDD1.n16 VDD1.t5 355.474
R201 VDD1.n6 VDD1.n5 171.744
R202 VDD1.n19 VDD1.n18 171.744
R203 VDD1.n27 VDD1.n26 158.505
R204 VDD1.n12 VDD1.n11 155.987
R205 VDD1.n29 VDD1.n28 155.987
R206 VDD1.n25 VDD1.n24 155.987
R207 VDD1.n5 VDD1.t9 85.8723
R208 VDD1.n18 VDD1.t5 85.8723
R209 VDD1.n12 VDD1.n10 56.5618
R210 VDD1.n25 VDD1.n23 56.5618
R211 VDD1.n29 VDD1.n27 44.5699
R212 VDD1.n4 VDD1.n3 15.8418
R213 VDD1.n17 VDD1.n16 15.8418
R214 VDD1.n7 VDD1.n2 12.8005
R215 VDD1.n20 VDD1.n15 12.8005
R216 VDD1.n28 VDD1.t3 12.407
R217 VDD1.n28 VDD1.t7 12.407
R218 VDD1.n11 VDD1.t6 12.407
R219 VDD1.n11 VDD1.t1 12.407
R220 VDD1.n26 VDD1.t2 12.407
R221 VDD1.n26 VDD1.t0 12.407
R222 VDD1.n24 VDD1.t8 12.407
R223 VDD1.n24 VDD1.t4 12.407
R224 VDD1.n8 VDD1.n0 12.0247
R225 VDD1.n21 VDD1.n13 12.0247
R226 VDD1.n10 VDD1.n9 9.45567
R227 VDD1.n23 VDD1.n22 9.45567
R228 VDD1.n9 VDD1.n8 9.3005
R229 VDD1.n2 VDD1.n1 9.3005
R230 VDD1.n22 VDD1.n21 9.3005
R231 VDD1.n15 VDD1.n14 9.3005
R232 VDD1.n3 VDD1.n1 4.29255
R233 VDD1.n16 VDD1.n14 4.29255
R234 VDD1 VDD1.n29 2.51559
R235 VDD1.n10 VDD1.n0 1.93989
R236 VDD1.n23 VDD1.n13 1.93989
R237 VDD1.n8 VDD1.n7 1.16414
R238 VDD1.n21 VDD1.n20 1.16414
R239 VDD1 VDD1.n12 0.916448
R240 VDD1.n27 VDD1.n25 0.802913
R241 VDD1.n4 VDD1.n2 0.388379
R242 VDD1.n17 VDD1.n15 0.388379
R243 VDD1.n9 VDD1.n1 0.155672
R244 VDD1.n22 VDD1.n14 0.155672
R245 VTAIL.n56 VTAIL.n50 756.745
R246 VTAIL.n8 VTAIL.n2 756.745
R247 VTAIL.n44 VTAIL.n38 756.745
R248 VTAIL.n28 VTAIL.n22 756.745
R249 VTAIL.n55 VTAIL.n54 585
R250 VTAIL.n57 VTAIL.n56 585
R251 VTAIL.n7 VTAIL.n6 585
R252 VTAIL.n9 VTAIL.n8 585
R253 VTAIL.n45 VTAIL.n44 585
R254 VTAIL.n43 VTAIL.n42 585
R255 VTAIL.n29 VTAIL.n28 585
R256 VTAIL.n27 VTAIL.n26 585
R257 VTAIL.n53 VTAIL.t19 355.474
R258 VTAIL.n5 VTAIL.t13 355.474
R259 VTAIL.n41 VTAIL.t12 355.474
R260 VTAIL.n25 VTAIL.t5 355.474
R261 VTAIL.n56 VTAIL.n55 171.744
R262 VTAIL.n8 VTAIL.n7 171.744
R263 VTAIL.n44 VTAIL.n43 171.744
R264 VTAIL.n28 VTAIL.n27 171.744
R265 VTAIL.n37 VTAIL.n36 139.309
R266 VTAIL.n35 VTAIL.n34 139.309
R267 VTAIL.n21 VTAIL.n20 139.309
R268 VTAIL.n19 VTAIL.n18 139.309
R269 VTAIL.n63 VTAIL.n62 139.309
R270 VTAIL.n1 VTAIL.n0 139.309
R271 VTAIL.n15 VTAIL.n14 139.309
R272 VTAIL.n17 VTAIL.n16 139.309
R273 VTAIL.n55 VTAIL.t19 85.8723
R274 VTAIL.n7 VTAIL.t13 85.8723
R275 VTAIL.n43 VTAIL.t12 85.8723
R276 VTAIL.n27 VTAIL.t5 85.8723
R277 VTAIL.n61 VTAIL.n60 36.452
R278 VTAIL.n13 VTAIL.n12 36.452
R279 VTAIL.n49 VTAIL.n48 36.452
R280 VTAIL.n33 VTAIL.n32 36.452
R281 VTAIL.n19 VTAIL.n17 21.4876
R282 VTAIL.n61 VTAIL.n49 18.0565
R283 VTAIL.n54 VTAIL.n53 15.8418
R284 VTAIL.n6 VTAIL.n5 15.8418
R285 VTAIL.n42 VTAIL.n41 15.8418
R286 VTAIL.n26 VTAIL.n25 15.8418
R287 VTAIL.n57 VTAIL.n52 12.8005
R288 VTAIL.n9 VTAIL.n4 12.8005
R289 VTAIL.n45 VTAIL.n40 12.8005
R290 VTAIL.n29 VTAIL.n24 12.8005
R291 VTAIL.n62 VTAIL.t18 12.407
R292 VTAIL.n62 VTAIL.t2 12.407
R293 VTAIL.n0 VTAIL.t3 12.407
R294 VTAIL.n0 VTAIL.t0 12.407
R295 VTAIL.n14 VTAIL.t14 12.407
R296 VTAIL.n14 VTAIL.t15 12.407
R297 VTAIL.n16 VTAIL.t7 12.407
R298 VTAIL.n16 VTAIL.t9 12.407
R299 VTAIL.n36 VTAIL.t6 12.407
R300 VTAIL.n36 VTAIL.t8 12.407
R301 VTAIL.n34 VTAIL.t10 12.407
R302 VTAIL.n34 VTAIL.t11 12.407
R303 VTAIL.n20 VTAIL.t16 12.407
R304 VTAIL.n20 VTAIL.t4 12.407
R305 VTAIL.n18 VTAIL.t1 12.407
R306 VTAIL.n18 VTAIL.t17 12.407
R307 VTAIL.n58 VTAIL.n50 12.0247
R308 VTAIL.n10 VTAIL.n2 12.0247
R309 VTAIL.n46 VTAIL.n38 12.0247
R310 VTAIL.n30 VTAIL.n22 12.0247
R311 VTAIL.n60 VTAIL.n59 9.45567
R312 VTAIL.n12 VTAIL.n11 9.45567
R313 VTAIL.n48 VTAIL.n47 9.45567
R314 VTAIL.n32 VTAIL.n31 9.45567
R315 VTAIL.n59 VTAIL.n58 9.3005
R316 VTAIL.n52 VTAIL.n51 9.3005
R317 VTAIL.n11 VTAIL.n10 9.3005
R318 VTAIL.n4 VTAIL.n3 9.3005
R319 VTAIL.n47 VTAIL.n46 9.3005
R320 VTAIL.n40 VTAIL.n39 9.3005
R321 VTAIL.n31 VTAIL.n30 9.3005
R322 VTAIL.n24 VTAIL.n23 9.3005
R323 VTAIL.n41 VTAIL.n39 4.29255
R324 VTAIL.n25 VTAIL.n23 4.29255
R325 VTAIL.n53 VTAIL.n51 4.29255
R326 VTAIL.n5 VTAIL.n3 4.29255
R327 VTAIL.n21 VTAIL.n19 3.43153
R328 VTAIL.n33 VTAIL.n21 3.43153
R329 VTAIL.n37 VTAIL.n35 3.43153
R330 VTAIL.n49 VTAIL.n37 3.43153
R331 VTAIL.n17 VTAIL.n15 3.43153
R332 VTAIL.n15 VTAIL.n13 3.43153
R333 VTAIL.n63 VTAIL.n61 3.43153
R334 VTAIL VTAIL.n1 2.63197
R335 VTAIL.n35 VTAIL.n33 2.18584
R336 VTAIL.n13 VTAIL.n1 2.18584
R337 VTAIL.n60 VTAIL.n50 1.93989
R338 VTAIL.n12 VTAIL.n2 1.93989
R339 VTAIL.n48 VTAIL.n38 1.93989
R340 VTAIL.n32 VTAIL.n22 1.93989
R341 VTAIL.n58 VTAIL.n57 1.16414
R342 VTAIL.n10 VTAIL.n9 1.16414
R343 VTAIL.n46 VTAIL.n45 1.16414
R344 VTAIL.n30 VTAIL.n29 1.16414
R345 VTAIL VTAIL.n63 0.800069
R346 VTAIL.n54 VTAIL.n52 0.388379
R347 VTAIL.n6 VTAIL.n4 0.388379
R348 VTAIL.n42 VTAIL.n40 0.388379
R349 VTAIL.n26 VTAIL.n24 0.388379
R350 VTAIL.n59 VTAIL.n51 0.155672
R351 VTAIL.n11 VTAIL.n3 0.155672
R352 VTAIL.n47 VTAIL.n39 0.155672
R353 VTAIL.n31 VTAIL.n23 0.155672
R354 VN.n106 VN.n105 161.3
R355 VN.n104 VN.n55 161.3
R356 VN.n103 VN.n102 161.3
R357 VN.n101 VN.n56 161.3
R358 VN.n100 VN.n99 161.3
R359 VN.n98 VN.n57 161.3
R360 VN.n97 VN.n96 161.3
R361 VN.n95 VN.n58 161.3
R362 VN.n94 VN.n93 161.3
R363 VN.n92 VN.n59 161.3
R364 VN.n91 VN.n90 161.3
R365 VN.n89 VN.n61 161.3
R366 VN.n88 VN.n87 161.3
R367 VN.n86 VN.n62 161.3
R368 VN.n85 VN.n84 161.3
R369 VN.n83 VN.n63 161.3
R370 VN.n82 VN.n81 161.3
R371 VN.n80 VN.n64 161.3
R372 VN.n79 VN.n78 161.3
R373 VN.n77 VN.n66 161.3
R374 VN.n76 VN.n75 161.3
R375 VN.n74 VN.n67 161.3
R376 VN.n73 VN.n72 161.3
R377 VN.n71 VN.n68 161.3
R378 VN.n52 VN.n51 161.3
R379 VN.n50 VN.n1 161.3
R380 VN.n49 VN.n48 161.3
R381 VN.n47 VN.n2 161.3
R382 VN.n46 VN.n45 161.3
R383 VN.n44 VN.n3 161.3
R384 VN.n43 VN.n42 161.3
R385 VN.n41 VN.n4 161.3
R386 VN.n40 VN.n39 161.3
R387 VN.n37 VN.n5 161.3
R388 VN.n36 VN.n35 161.3
R389 VN.n34 VN.n6 161.3
R390 VN.n33 VN.n32 161.3
R391 VN.n31 VN.n7 161.3
R392 VN.n30 VN.n29 161.3
R393 VN.n28 VN.n8 161.3
R394 VN.n27 VN.n26 161.3
R395 VN.n24 VN.n9 161.3
R396 VN.n23 VN.n22 161.3
R397 VN.n21 VN.n10 161.3
R398 VN.n20 VN.n19 161.3
R399 VN.n18 VN.n11 161.3
R400 VN.n17 VN.n16 161.3
R401 VN.n15 VN.n12 161.3
R402 VN.n53 VN.n0 79.917
R403 VN.n107 VN.n54 79.917
R404 VN.n14 VN.n13 63.5339
R405 VN.n70 VN.n69 63.5339
R406 VN.n32 VN.n6 56.5617
R407 VN.n87 VN.n61 56.5617
R408 VN.n19 VN.n10 56.5617
R409 VN.n45 VN.n2 56.5617
R410 VN.n75 VN.n66 56.5617
R411 VN.n99 VN.n56 56.5617
R412 VN VN.n107 52.0133
R413 VN.n70 VN.t4 50.8211
R414 VN.n14 VN.t8 50.8211
R415 VN.n17 VN.n12 24.5923
R416 VN.n18 VN.n17 24.5923
R417 VN.n19 VN.n18 24.5923
R418 VN.n23 VN.n10 24.5923
R419 VN.n24 VN.n23 24.5923
R420 VN.n26 VN.n24 24.5923
R421 VN.n30 VN.n8 24.5923
R422 VN.n31 VN.n30 24.5923
R423 VN.n32 VN.n31 24.5923
R424 VN.n36 VN.n6 24.5923
R425 VN.n37 VN.n36 24.5923
R426 VN.n39 VN.n37 24.5923
R427 VN.n43 VN.n4 24.5923
R428 VN.n44 VN.n43 24.5923
R429 VN.n45 VN.n44 24.5923
R430 VN.n49 VN.n2 24.5923
R431 VN.n50 VN.n49 24.5923
R432 VN.n51 VN.n50 24.5923
R433 VN.n75 VN.n74 24.5923
R434 VN.n74 VN.n73 24.5923
R435 VN.n73 VN.n68 24.5923
R436 VN.n87 VN.n86 24.5923
R437 VN.n86 VN.n85 24.5923
R438 VN.n85 VN.n63 24.5923
R439 VN.n81 VN.n80 24.5923
R440 VN.n80 VN.n79 24.5923
R441 VN.n79 VN.n66 24.5923
R442 VN.n99 VN.n98 24.5923
R443 VN.n98 VN.n97 24.5923
R444 VN.n97 VN.n58 24.5923
R445 VN.n93 VN.n92 24.5923
R446 VN.n92 VN.n91 24.5923
R447 VN.n91 VN.n61 24.5923
R448 VN.n105 VN.n104 24.5923
R449 VN.n104 VN.n103 24.5923
R450 VN.n103 VN.n56 24.5923
R451 VN.n13 VN.t7 17.2997
R452 VN.n25 VN.t0 17.2997
R453 VN.n38 VN.t1 17.2997
R454 VN.n0 VN.t6 17.2997
R455 VN.n69 VN.t2 17.2997
R456 VN.n65 VN.t3 17.2997
R457 VN.n60 VN.t9 17.2997
R458 VN.n54 VN.t5 17.2997
R459 VN.n38 VN.n4 13.2801
R460 VN.n60 VN.n58 13.2801
R461 VN.n26 VN.n25 12.2964
R462 VN.n25 VN.n8 12.2964
R463 VN.n65 VN.n63 12.2964
R464 VN.n81 VN.n65 12.2964
R465 VN.n13 VN.n12 11.3127
R466 VN.n39 VN.n38 11.3127
R467 VN.n69 VN.n68 11.3127
R468 VN.n93 VN.n60 11.3127
R469 VN.n51 VN.n0 10.3291
R470 VN.n105 VN.n54 10.3291
R471 VN.n71 VN.n70 3.13518
R472 VN.n15 VN.n14 3.13518
R473 VN.n107 VN.n106 0.354861
R474 VN.n53 VN.n52 0.354861
R475 VN VN.n53 0.267071
R476 VN.n106 VN.n55 0.189894
R477 VN.n102 VN.n55 0.189894
R478 VN.n102 VN.n101 0.189894
R479 VN.n101 VN.n100 0.189894
R480 VN.n100 VN.n57 0.189894
R481 VN.n96 VN.n57 0.189894
R482 VN.n96 VN.n95 0.189894
R483 VN.n95 VN.n94 0.189894
R484 VN.n94 VN.n59 0.189894
R485 VN.n90 VN.n59 0.189894
R486 VN.n90 VN.n89 0.189894
R487 VN.n89 VN.n88 0.189894
R488 VN.n88 VN.n62 0.189894
R489 VN.n84 VN.n62 0.189894
R490 VN.n84 VN.n83 0.189894
R491 VN.n83 VN.n82 0.189894
R492 VN.n82 VN.n64 0.189894
R493 VN.n78 VN.n64 0.189894
R494 VN.n78 VN.n77 0.189894
R495 VN.n77 VN.n76 0.189894
R496 VN.n76 VN.n67 0.189894
R497 VN.n72 VN.n67 0.189894
R498 VN.n72 VN.n71 0.189894
R499 VN.n16 VN.n15 0.189894
R500 VN.n16 VN.n11 0.189894
R501 VN.n20 VN.n11 0.189894
R502 VN.n21 VN.n20 0.189894
R503 VN.n22 VN.n21 0.189894
R504 VN.n22 VN.n9 0.189894
R505 VN.n27 VN.n9 0.189894
R506 VN.n28 VN.n27 0.189894
R507 VN.n29 VN.n28 0.189894
R508 VN.n29 VN.n7 0.189894
R509 VN.n33 VN.n7 0.189894
R510 VN.n34 VN.n33 0.189894
R511 VN.n35 VN.n34 0.189894
R512 VN.n35 VN.n5 0.189894
R513 VN.n40 VN.n5 0.189894
R514 VN.n41 VN.n40 0.189894
R515 VN.n42 VN.n41 0.189894
R516 VN.n42 VN.n3 0.189894
R517 VN.n46 VN.n3 0.189894
R518 VN.n47 VN.n46 0.189894
R519 VN.n48 VN.n47 0.189894
R520 VN.n48 VN.n1 0.189894
R521 VN.n52 VN.n1 0.189894
R522 VDD2.n21 VDD2.n15 756.745
R523 VDD2.n6 VDD2.n0 756.745
R524 VDD2.n22 VDD2.n21 585
R525 VDD2.n20 VDD2.n19 585
R526 VDD2.n5 VDD2.n4 585
R527 VDD2.n7 VDD2.n6 585
R528 VDD2.n18 VDD2.t4 355.474
R529 VDD2.n3 VDD2.t1 355.474
R530 VDD2.n21 VDD2.n20 171.744
R531 VDD2.n6 VDD2.n5 171.744
R532 VDD2.n14 VDD2.n13 158.505
R533 VDD2 VDD2.n29 158.501
R534 VDD2.n28 VDD2.n27 155.987
R535 VDD2.n12 VDD2.n11 155.987
R536 VDD2.n20 VDD2.t4 85.8723
R537 VDD2.n5 VDD2.t1 85.8723
R538 VDD2.n12 VDD2.n10 56.5618
R539 VDD2.n26 VDD2.n25 53.1308
R540 VDD2.n26 VDD2.n14 42.2713
R541 VDD2.n19 VDD2.n18 15.8418
R542 VDD2.n4 VDD2.n3 15.8418
R543 VDD2.n22 VDD2.n17 12.8005
R544 VDD2.n7 VDD2.n2 12.8005
R545 VDD2.n29 VDD2.t7 12.407
R546 VDD2.n29 VDD2.t5 12.407
R547 VDD2.n27 VDD2.t0 12.407
R548 VDD2.n27 VDD2.t6 12.407
R549 VDD2.n13 VDD2.t8 12.407
R550 VDD2.n13 VDD2.t3 12.407
R551 VDD2.n11 VDD2.t2 12.407
R552 VDD2.n11 VDD2.t9 12.407
R553 VDD2.n23 VDD2.n15 12.0247
R554 VDD2.n8 VDD2.n0 12.0247
R555 VDD2.n25 VDD2.n24 9.45567
R556 VDD2.n10 VDD2.n9 9.45567
R557 VDD2.n24 VDD2.n23 9.3005
R558 VDD2.n17 VDD2.n16 9.3005
R559 VDD2.n9 VDD2.n8 9.3005
R560 VDD2.n2 VDD2.n1 9.3005
R561 VDD2.n18 VDD2.n16 4.29255
R562 VDD2.n3 VDD2.n1 4.29255
R563 VDD2.n28 VDD2.n26 3.43153
R564 VDD2.n25 VDD2.n15 1.93989
R565 VDD2.n10 VDD2.n0 1.93989
R566 VDD2.n23 VDD2.n22 1.16414
R567 VDD2.n8 VDD2.n7 1.16414
R568 VDD2 VDD2.n28 0.916448
R569 VDD2.n14 VDD2.n12 0.802913
R570 VDD2.n19 VDD2.n17 0.388379
R571 VDD2.n4 VDD2.n2 0.388379
R572 VDD2.n24 VDD2.n16 0.155672
R573 VDD2.n9 VDD2.n1 0.155672
R574 B.n379 B.n378 585
R575 B.n377 B.n144 585
R576 B.n376 B.n375 585
R577 B.n374 B.n145 585
R578 B.n373 B.n372 585
R579 B.n371 B.n146 585
R580 B.n370 B.n369 585
R581 B.n368 B.n147 585
R582 B.n367 B.n366 585
R583 B.n365 B.n148 585
R584 B.n364 B.n363 585
R585 B.n362 B.n149 585
R586 B.n361 B.n360 585
R587 B.n359 B.n150 585
R588 B.n358 B.n357 585
R589 B.n353 B.n151 585
R590 B.n352 B.n351 585
R591 B.n350 B.n152 585
R592 B.n349 B.n348 585
R593 B.n347 B.n153 585
R594 B.n346 B.n345 585
R595 B.n344 B.n154 585
R596 B.n343 B.n342 585
R597 B.n341 B.n155 585
R598 B.n339 B.n338 585
R599 B.n337 B.n158 585
R600 B.n336 B.n335 585
R601 B.n334 B.n159 585
R602 B.n333 B.n332 585
R603 B.n331 B.n160 585
R604 B.n330 B.n329 585
R605 B.n328 B.n161 585
R606 B.n327 B.n326 585
R607 B.n325 B.n162 585
R608 B.n324 B.n323 585
R609 B.n322 B.n163 585
R610 B.n321 B.n320 585
R611 B.n319 B.n164 585
R612 B.n380 B.n143 585
R613 B.n382 B.n381 585
R614 B.n383 B.n142 585
R615 B.n385 B.n384 585
R616 B.n386 B.n141 585
R617 B.n388 B.n387 585
R618 B.n389 B.n140 585
R619 B.n391 B.n390 585
R620 B.n392 B.n139 585
R621 B.n394 B.n393 585
R622 B.n395 B.n138 585
R623 B.n397 B.n396 585
R624 B.n398 B.n137 585
R625 B.n400 B.n399 585
R626 B.n401 B.n136 585
R627 B.n403 B.n402 585
R628 B.n404 B.n135 585
R629 B.n406 B.n405 585
R630 B.n407 B.n134 585
R631 B.n409 B.n408 585
R632 B.n410 B.n133 585
R633 B.n412 B.n411 585
R634 B.n413 B.n132 585
R635 B.n415 B.n414 585
R636 B.n416 B.n131 585
R637 B.n418 B.n417 585
R638 B.n419 B.n130 585
R639 B.n421 B.n420 585
R640 B.n422 B.n129 585
R641 B.n424 B.n423 585
R642 B.n425 B.n128 585
R643 B.n427 B.n426 585
R644 B.n428 B.n127 585
R645 B.n430 B.n429 585
R646 B.n431 B.n126 585
R647 B.n433 B.n432 585
R648 B.n434 B.n125 585
R649 B.n436 B.n435 585
R650 B.n437 B.n124 585
R651 B.n439 B.n438 585
R652 B.n440 B.n123 585
R653 B.n442 B.n441 585
R654 B.n443 B.n122 585
R655 B.n445 B.n444 585
R656 B.n446 B.n121 585
R657 B.n448 B.n447 585
R658 B.n449 B.n120 585
R659 B.n451 B.n450 585
R660 B.n452 B.n119 585
R661 B.n454 B.n453 585
R662 B.n455 B.n118 585
R663 B.n457 B.n456 585
R664 B.n458 B.n117 585
R665 B.n460 B.n459 585
R666 B.n461 B.n116 585
R667 B.n463 B.n462 585
R668 B.n464 B.n115 585
R669 B.n466 B.n465 585
R670 B.n467 B.n114 585
R671 B.n469 B.n468 585
R672 B.n470 B.n113 585
R673 B.n472 B.n471 585
R674 B.n473 B.n112 585
R675 B.n475 B.n474 585
R676 B.n476 B.n111 585
R677 B.n478 B.n477 585
R678 B.n479 B.n110 585
R679 B.n481 B.n480 585
R680 B.n482 B.n109 585
R681 B.n484 B.n483 585
R682 B.n485 B.n108 585
R683 B.n487 B.n486 585
R684 B.n488 B.n107 585
R685 B.n490 B.n489 585
R686 B.n491 B.n106 585
R687 B.n493 B.n492 585
R688 B.n494 B.n105 585
R689 B.n496 B.n495 585
R690 B.n497 B.n104 585
R691 B.n499 B.n498 585
R692 B.n500 B.n103 585
R693 B.n502 B.n501 585
R694 B.n503 B.n102 585
R695 B.n505 B.n504 585
R696 B.n506 B.n101 585
R697 B.n508 B.n507 585
R698 B.n509 B.n100 585
R699 B.n511 B.n510 585
R700 B.n512 B.n99 585
R701 B.n514 B.n513 585
R702 B.n515 B.n98 585
R703 B.n517 B.n516 585
R704 B.n518 B.n97 585
R705 B.n520 B.n519 585
R706 B.n521 B.n96 585
R707 B.n523 B.n522 585
R708 B.n524 B.n95 585
R709 B.n526 B.n525 585
R710 B.n527 B.n94 585
R711 B.n529 B.n528 585
R712 B.n530 B.n93 585
R713 B.n532 B.n531 585
R714 B.n533 B.n92 585
R715 B.n535 B.n534 585
R716 B.n536 B.n91 585
R717 B.n538 B.n537 585
R718 B.n539 B.n90 585
R719 B.n541 B.n540 585
R720 B.n542 B.n89 585
R721 B.n544 B.n543 585
R722 B.n545 B.n88 585
R723 B.n547 B.n546 585
R724 B.n548 B.n87 585
R725 B.n550 B.n549 585
R726 B.n551 B.n86 585
R727 B.n553 B.n552 585
R728 B.n554 B.n85 585
R729 B.n556 B.n555 585
R730 B.n557 B.n84 585
R731 B.n559 B.n558 585
R732 B.n560 B.n83 585
R733 B.n562 B.n561 585
R734 B.n563 B.n82 585
R735 B.n565 B.n564 585
R736 B.n566 B.n81 585
R737 B.n568 B.n567 585
R738 B.n569 B.n80 585
R739 B.n571 B.n570 585
R740 B.n572 B.n79 585
R741 B.n574 B.n573 585
R742 B.n575 B.n78 585
R743 B.n577 B.n576 585
R744 B.n578 B.n77 585
R745 B.n580 B.n579 585
R746 B.n581 B.n76 585
R747 B.n583 B.n582 585
R748 B.n584 B.n75 585
R749 B.n586 B.n585 585
R750 B.n587 B.n74 585
R751 B.n589 B.n588 585
R752 B.n590 B.n73 585
R753 B.n592 B.n591 585
R754 B.n593 B.n72 585
R755 B.n595 B.n594 585
R756 B.n596 B.n71 585
R757 B.n598 B.n597 585
R758 B.n599 B.n70 585
R759 B.n601 B.n600 585
R760 B.n602 B.n69 585
R761 B.n604 B.n603 585
R762 B.n605 B.n68 585
R763 B.n607 B.n606 585
R764 B.n608 B.n67 585
R765 B.n610 B.n609 585
R766 B.n611 B.n66 585
R767 B.n613 B.n612 585
R768 B.n614 B.n65 585
R769 B.n616 B.n615 585
R770 B.n674 B.n41 585
R771 B.n673 B.n672 585
R772 B.n671 B.n42 585
R773 B.n670 B.n669 585
R774 B.n668 B.n43 585
R775 B.n667 B.n666 585
R776 B.n665 B.n44 585
R777 B.n664 B.n663 585
R778 B.n662 B.n45 585
R779 B.n661 B.n660 585
R780 B.n659 B.n46 585
R781 B.n658 B.n657 585
R782 B.n656 B.n47 585
R783 B.n655 B.n654 585
R784 B.n653 B.n652 585
R785 B.n651 B.n51 585
R786 B.n650 B.n649 585
R787 B.n648 B.n52 585
R788 B.n647 B.n646 585
R789 B.n645 B.n53 585
R790 B.n644 B.n643 585
R791 B.n642 B.n54 585
R792 B.n641 B.n640 585
R793 B.n639 B.n55 585
R794 B.n637 B.n636 585
R795 B.n635 B.n58 585
R796 B.n634 B.n633 585
R797 B.n632 B.n59 585
R798 B.n631 B.n630 585
R799 B.n629 B.n60 585
R800 B.n628 B.n627 585
R801 B.n626 B.n61 585
R802 B.n625 B.n624 585
R803 B.n623 B.n62 585
R804 B.n622 B.n621 585
R805 B.n620 B.n63 585
R806 B.n619 B.n618 585
R807 B.n617 B.n64 585
R808 B.n676 B.n675 585
R809 B.n677 B.n40 585
R810 B.n679 B.n678 585
R811 B.n680 B.n39 585
R812 B.n682 B.n681 585
R813 B.n683 B.n38 585
R814 B.n685 B.n684 585
R815 B.n686 B.n37 585
R816 B.n688 B.n687 585
R817 B.n689 B.n36 585
R818 B.n691 B.n690 585
R819 B.n692 B.n35 585
R820 B.n694 B.n693 585
R821 B.n695 B.n34 585
R822 B.n697 B.n696 585
R823 B.n698 B.n33 585
R824 B.n700 B.n699 585
R825 B.n701 B.n32 585
R826 B.n703 B.n702 585
R827 B.n704 B.n31 585
R828 B.n706 B.n705 585
R829 B.n707 B.n30 585
R830 B.n709 B.n708 585
R831 B.n710 B.n29 585
R832 B.n712 B.n711 585
R833 B.n713 B.n28 585
R834 B.n715 B.n714 585
R835 B.n716 B.n27 585
R836 B.n718 B.n717 585
R837 B.n719 B.n26 585
R838 B.n721 B.n720 585
R839 B.n722 B.n25 585
R840 B.n724 B.n723 585
R841 B.n725 B.n24 585
R842 B.n727 B.n726 585
R843 B.n728 B.n23 585
R844 B.n730 B.n729 585
R845 B.n731 B.n22 585
R846 B.n733 B.n732 585
R847 B.n734 B.n21 585
R848 B.n736 B.n735 585
R849 B.n737 B.n20 585
R850 B.n739 B.n738 585
R851 B.n740 B.n19 585
R852 B.n742 B.n741 585
R853 B.n743 B.n18 585
R854 B.n745 B.n744 585
R855 B.n746 B.n17 585
R856 B.n748 B.n747 585
R857 B.n749 B.n16 585
R858 B.n751 B.n750 585
R859 B.n752 B.n15 585
R860 B.n754 B.n753 585
R861 B.n755 B.n14 585
R862 B.n757 B.n756 585
R863 B.n758 B.n13 585
R864 B.n760 B.n759 585
R865 B.n761 B.n12 585
R866 B.n763 B.n762 585
R867 B.n764 B.n11 585
R868 B.n766 B.n765 585
R869 B.n767 B.n10 585
R870 B.n769 B.n768 585
R871 B.n770 B.n9 585
R872 B.n772 B.n771 585
R873 B.n773 B.n8 585
R874 B.n775 B.n774 585
R875 B.n776 B.n7 585
R876 B.n778 B.n777 585
R877 B.n779 B.n6 585
R878 B.n781 B.n780 585
R879 B.n782 B.n5 585
R880 B.n784 B.n783 585
R881 B.n785 B.n4 585
R882 B.n787 B.n786 585
R883 B.n788 B.n3 585
R884 B.n790 B.n789 585
R885 B.n791 B.n0 585
R886 B.n2 B.n1 585
R887 B.n204 B.n203 585
R888 B.n205 B.n202 585
R889 B.n207 B.n206 585
R890 B.n208 B.n201 585
R891 B.n210 B.n209 585
R892 B.n211 B.n200 585
R893 B.n213 B.n212 585
R894 B.n214 B.n199 585
R895 B.n216 B.n215 585
R896 B.n217 B.n198 585
R897 B.n219 B.n218 585
R898 B.n220 B.n197 585
R899 B.n222 B.n221 585
R900 B.n223 B.n196 585
R901 B.n225 B.n224 585
R902 B.n226 B.n195 585
R903 B.n228 B.n227 585
R904 B.n229 B.n194 585
R905 B.n231 B.n230 585
R906 B.n232 B.n193 585
R907 B.n234 B.n233 585
R908 B.n235 B.n192 585
R909 B.n237 B.n236 585
R910 B.n238 B.n191 585
R911 B.n240 B.n239 585
R912 B.n241 B.n190 585
R913 B.n243 B.n242 585
R914 B.n244 B.n189 585
R915 B.n246 B.n245 585
R916 B.n247 B.n188 585
R917 B.n249 B.n248 585
R918 B.n250 B.n187 585
R919 B.n252 B.n251 585
R920 B.n253 B.n186 585
R921 B.n255 B.n254 585
R922 B.n256 B.n185 585
R923 B.n258 B.n257 585
R924 B.n259 B.n184 585
R925 B.n261 B.n260 585
R926 B.n262 B.n183 585
R927 B.n264 B.n263 585
R928 B.n265 B.n182 585
R929 B.n267 B.n266 585
R930 B.n268 B.n181 585
R931 B.n270 B.n269 585
R932 B.n271 B.n180 585
R933 B.n273 B.n272 585
R934 B.n274 B.n179 585
R935 B.n276 B.n275 585
R936 B.n277 B.n178 585
R937 B.n279 B.n278 585
R938 B.n280 B.n177 585
R939 B.n282 B.n281 585
R940 B.n283 B.n176 585
R941 B.n285 B.n284 585
R942 B.n286 B.n175 585
R943 B.n288 B.n287 585
R944 B.n289 B.n174 585
R945 B.n291 B.n290 585
R946 B.n292 B.n173 585
R947 B.n294 B.n293 585
R948 B.n295 B.n172 585
R949 B.n297 B.n296 585
R950 B.n298 B.n171 585
R951 B.n300 B.n299 585
R952 B.n301 B.n170 585
R953 B.n303 B.n302 585
R954 B.n304 B.n169 585
R955 B.n306 B.n305 585
R956 B.n307 B.n168 585
R957 B.n309 B.n308 585
R958 B.n310 B.n167 585
R959 B.n312 B.n311 585
R960 B.n313 B.n166 585
R961 B.n315 B.n314 585
R962 B.n316 B.n165 585
R963 B.n318 B.n317 585
R964 B.n319 B.n318 444.452
R965 B.n378 B.n143 444.452
R966 B.n617 B.n616 444.452
R967 B.n676 B.n41 444.452
R968 B.n354 B.t10 303.767
R969 B.n56 B.t5 303.767
R970 B.n156 B.t7 303.767
R971 B.n48 B.t2 303.767
R972 B.n793 B.n792 256.663
R973 B.n792 B.n791 235.042
R974 B.n792 B.n2 235.042
R975 B.n355 B.t11 226.578
R976 B.n57 B.t4 226.578
R977 B.n157 B.t8 226.578
R978 B.n49 B.t1 226.578
R979 B.n156 B.t6 226.523
R980 B.n354 B.t9 226.523
R981 B.n56 B.t3 226.523
R982 B.n48 B.t0 226.523
R983 B.n320 B.n319 163.367
R984 B.n320 B.n163 163.367
R985 B.n324 B.n163 163.367
R986 B.n325 B.n324 163.367
R987 B.n326 B.n325 163.367
R988 B.n326 B.n161 163.367
R989 B.n330 B.n161 163.367
R990 B.n331 B.n330 163.367
R991 B.n332 B.n331 163.367
R992 B.n332 B.n159 163.367
R993 B.n336 B.n159 163.367
R994 B.n337 B.n336 163.367
R995 B.n338 B.n337 163.367
R996 B.n338 B.n155 163.367
R997 B.n343 B.n155 163.367
R998 B.n344 B.n343 163.367
R999 B.n345 B.n344 163.367
R1000 B.n345 B.n153 163.367
R1001 B.n349 B.n153 163.367
R1002 B.n350 B.n349 163.367
R1003 B.n351 B.n350 163.367
R1004 B.n351 B.n151 163.367
R1005 B.n358 B.n151 163.367
R1006 B.n359 B.n358 163.367
R1007 B.n360 B.n359 163.367
R1008 B.n360 B.n149 163.367
R1009 B.n364 B.n149 163.367
R1010 B.n365 B.n364 163.367
R1011 B.n366 B.n365 163.367
R1012 B.n366 B.n147 163.367
R1013 B.n370 B.n147 163.367
R1014 B.n371 B.n370 163.367
R1015 B.n372 B.n371 163.367
R1016 B.n372 B.n145 163.367
R1017 B.n376 B.n145 163.367
R1018 B.n377 B.n376 163.367
R1019 B.n378 B.n377 163.367
R1020 B.n616 B.n65 163.367
R1021 B.n612 B.n65 163.367
R1022 B.n612 B.n611 163.367
R1023 B.n611 B.n610 163.367
R1024 B.n610 B.n67 163.367
R1025 B.n606 B.n67 163.367
R1026 B.n606 B.n605 163.367
R1027 B.n605 B.n604 163.367
R1028 B.n604 B.n69 163.367
R1029 B.n600 B.n69 163.367
R1030 B.n600 B.n599 163.367
R1031 B.n599 B.n598 163.367
R1032 B.n598 B.n71 163.367
R1033 B.n594 B.n71 163.367
R1034 B.n594 B.n593 163.367
R1035 B.n593 B.n592 163.367
R1036 B.n592 B.n73 163.367
R1037 B.n588 B.n73 163.367
R1038 B.n588 B.n587 163.367
R1039 B.n587 B.n586 163.367
R1040 B.n586 B.n75 163.367
R1041 B.n582 B.n75 163.367
R1042 B.n582 B.n581 163.367
R1043 B.n581 B.n580 163.367
R1044 B.n580 B.n77 163.367
R1045 B.n576 B.n77 163.367
R1046 B.n576 B.n575 163.367
R1047 B.n575 B.n574 163.367
R1048 B.n574 B.n79 163.367
R1049 B.n570 B.n79 163.367
R1050 B.n570 B.n569 163.367
R1051 B.n569 B.n568 163.367
R1052 B.n568 B.n81 163.367
R1053 B.n564 B.n81 163.367
R1054 B.n564 B.n563 163.367
R1055 B.n563 B.n562 163.367
R1056 B.n562 B.n83 163.367
R1057 B.n558 B.n83 163.367
R1058 B.n558 B.n557 163.367
R1059 B.n557 B.n556 163.367
R1060 B.n556 B.n85 163.367
R1061 B.n552 B.n85 163.367
R1062 B.n552 B.n551 163.367
R1063 B.n551 B.n550 163.367
R1064 B.n550 B.n87 163.367
R1065 B.n546 B.n87 163.367
R1066 B.n546 B.n545 163.367
R1067 B.n545 B.n544 163.367
R1068 B.n544 B.n89 163.367
R1069 B.n540 B.n89 163.367
R1070 B.n540 B.n539 163.367
R1071 B.n539 B.n538 163.367
R1072 B.n538 B.n91 163.367
R1073 B.n534 B.n91 163.367
R1074 B.n534 B.n533 163.367
R1075 B.n533 B.n532 163.367
R1076 B.n532 B.n93 163.367
R1077 B.n528 B.n93 163.367
R1078 B.n528 B.n527 163.367
R1079 B.n527 B.n526 163.367
R1080 B.n526 B.n95 163.367
R1081 B.n522 B.n95 163.367
R1082 B.n522 B.n521 163.367
R1083 B.n521 B.n520 163.367
R1084 B.n520 B.n97 163.367
R1085 B.n516 B.n97 163.367
R1086 B.n516 B.n515 163.367
R1087 B.n515 B.n514 163.367
R1088 B.n514 B.n99 163.367
R1089 B.n510 B.n99 163.367
R1090 B.n510 B.n509 163.367
R1091 B.n509 B.n508 163.367
R1092 B.n508 B.n101 163.367
R1093 B.n504 B.n101 163.367
R1094 B.n504 B.n503 163.367
R1095 B.n503 B.n502 163.367
R1096 B.n502 B.n103 163.367
R1097 B.n498 B.n103 163.367
R1098 B.n498 B.n497 163.367
R1099 B.n497 B.n496 163.367
R1100 B.n496 B.n105 163.367
R1101 B.n492 B.n105 163.367
R1102 B.n492 B.n491 163.367
R1103 B.n491 B.n490 163.367
R1104 B.n490 B.n107 163.367
R1105 B.n486 B.n107 163.367
R1106 B.n486 B.n485 163.367
R1107 B.n485 B.n484 163.367
R1108 B.n484 B.n109 163.367
R1109 B.n480 B.n109 163.367
R1110 B.n480 B.n479 163.367
R1111 B.n479 B.n478 163.367
R1112 B.n478 B.n111 163.367
R1113 B.n474 B.n111 163.367
R1114 B.n474 B.n473 163.367
R1115 B.n473 B.n472 163.367
R1116 B.n472 B.n113 163.367
R1117 B.n468 B.n113 163.367
R1118 B.n468 B.n467 163.367
R1119 B.n467 B.n466 163.367
R1120 B.n466 B.n115 163.367
R1121 B.n462 B.n115 163.367
R1122 B.n462 B.n461 163.367
R1123 B.n461 B.n460 163.367
R1124 B.n460 B.n117 163.367
R1125 B.n456 B.n117 163.367
R1126 B.n456 B.n455 163.367
R1127 B.n455 B.n454 163.367
R1128 B.n454 B.n119 163.367
R1129 B.n450 B.n119 163.367
R1130 B.n450 B.n449 163.367
R1131 B.n449 B.n448 163.367
R1132 B.n448 B.n121 163.367
R1133 B.n444 B.n121 163.367
R1134 B.n444 B.n443 163.367
R1135 B.n443 B.n442 163.367
R1136 B.n442 B.n123 163.367
R1137 B.n438 B.n123 163.367
R1138 B.n438 B.n437 163.367
R1139 B.n437 B.n436 163.367
R1140 B.n436 B.n125 163.367
R1141 B.n432 B.n125 163.367
R1142 B.n432 B.n431 163.367
R1143 B.n431 B.n430 163.367
R1144 B.n430 B.n127 163.367
R1145 B.n426 B.n127 163.367
R1146 B.n426 B.n425 163.367
R1147 B.n425 B.n424 163.367
R1148 B.n424 B.n129 163.367
R1149 B.n420 B.n129 163.367
R1150 B.n420 B.n419 163.367
R1151 B.n419 B.n418 163.367
R1152 B.n418 B.n131 163.367
R1153 B.n414 B.n131 163.367
R1154 B.n414 B.n413 163.367
R1155 B.n413 B.n412 163.367
R1156 B.n412 B.n133 163.367
R1157 B.n408 B.n133 163.367
R1158 B.n408 B.n407 163.367
R1159 B.n407 B.n406 163.367
R1160 B.n406 B.n135 163.367
R1161 B.n402 B.n135 163.367
R1162 B.n402 B.n401 163.367
R1163 B.n401 B.n400 163.367
R1164 B.n400 B.n137 163.367
R1165 B.n396 B.n137 163.367
R1166 B.n396 B.n395 163.367
R1167 B.n395 B.n394 163.367
R1168 B.n394 B.n139 163.367
R1169 B.n390 B.n139 163.367
R1170 B.n390 B.n389 163.367
R1171 B.n389 B.n388 163.367
R1172 B.n388 B.n141 163.367
R1173 B.n384 B.n141 163.367
R1174 B.n384 B.n383 163.367
R1175 B.n383 B.n382 163.367
R1176 B.n382 B.n143 163.367
R1177 B.n672 B.n41 163.367
R1178 B.n672 B.n671 163.367
R1179 B.n671 B.n670 163.367
R1180 B.n670 B.n43 163.367
R1181 B.n666 B.n43 163.367
R1182 B.n666 B.n665 163.367
R1183 B.n665 B.n664 163.367
R1184 B.n664 B.n45 163.367
R1185 B.n660 B.n45 163.367
R1186 B.n660 B.n659 163.367
R1187 B.n659 B.n658 163.367
R1188 B.n658 B.n47 163.367
R1189 B.n654 B.n47 163.367
R1190 B.n654 B.n653 163.367
R1191 B.n653 B.n51 163.367
R1192 B.n649 B.n51 163.367
R1193 B.n649 B.n648 163.367
R1194 B.n648 B.n647 163.367
R1195 B.n647 B.n53 163.367
R1196 B.n643 B.n53 163.367
R1197 B.n643 B.n642 163.367
R1198 B.n642 B.n641 163.367
R1199 B.n641 B.n55 163.367
R1200 B.n636 B.n55 163.367
R1201 B.n636 B.n635 163.367
R1202 B.n635 B.n634 163.367
R1203 B.n634 B.n59 163.367
R1204 B.n630 B.n59 163.367
R1205 B.n630 B.n629 163.367
R1206 B.n629 B.n628 163.367
R1207 B.n628 B.n61 163.367
R1208 B.n624 B.n61 163.367
R1209 B.n624 B.n623 163.367
R1210 B.n623 B.n622 163.367
R1211 B.n622 B.n63 163.367
R1212 B.n618 B.n63 163.367
R1213 B.n618 B.n617 163.367
R1214 B.n677 B.n676 163.367
R1215 B.n678 B.n677 163.367
R1216 B.n678 B.n39 163.367
R1217 B.n682 B.n39 163.367
R1218 B.n683 B.n682 163.367
R1219 B.n684 B.n683 163.367
R1220 B.n684 B.n37 163.367
R1221 B.n688 B.n37 163.367
R1222 B.n689 B.n688 163.367
R1223 B.n690 B.n689 163.367
R1224 B.n690 B.n35 163.367
R1225 B.n694 B.n35 163.367
R1226 B.n695 B.n694 163.367
R1227 B.n696 B.n695 163.367
R1228 B.n696 B.n33 163.367
R1229 B.n700 B.n33 163.367
R1230 B.n701 B.n700 163.367
R1231 B.n702 B.n701 163.367
R1232 B.n702 B.n31 163.367
R1233 B.n706 B.n31 163.367
R1234 B.n707 B.n706 163.367
R1235 B.n708 B.n707 163.367
R1236 B.n708 B.n29 163.367
R1237 B.n712 B.n29 163.367
R1238 B.n713 B.n712 163.367
R1239 B.n714 B.n713 163.367
R1240 B.n714 B.n27 163.367
R1241 B.n718 B.n27 163.367
R1242 B.n719 B.n718 163.367
R1243 B.n720 B.n719 163.367
R1244 B.n720 B.n25 163.367
R1245 B.n724 B.n25 163.367
R1246 B.n725 B.n724 163.367
R1247 B.n726 B.n725 163.367
R1248 B.n726 B.n23 163.367
R1249 B.n730 B.n23 163.367
R1250 B.n731 B.n730 163.367
R1251 B.n732 B.n731 163.367
R1252 B.n732 B.n21 163.367
R1253 B.n736 B.n21 163.367
R1254 B.n737 B.n736 163.367
R1255 B.n738 B.n737 163.367
R1256 B.n738 B.n19 163.367
R1257 B.n742 B.n19 163.367
R1258 B.n743 B.n742 163.367
R1259 B.n744 B.n743 163.367
R1260 B.n744 B.n17 163.367
R1261 B.n748 B.n17 163.367
R1262 B.n749 B.n748 163.367
R1263 B.n750 B.n749 163.367
R1264 B.n750 B.n15 163.367
R1265 B.n754 B.n15 163.367
R1266 B.n755 B.n754 163.367
R1267 B.n756 B.n755 163.367
R1268 B.n756 B.n13 163.367
R1269 B.n760 B.n13 163.367
R1270 B.n761 B.n760 163.367
R1271 B.n762 B.n761 163.367
R1272 B.n762 B.n11 163.367
R1273 B.n766 B.n11 163.367
R1274 B.n767 B.n766 163.367
R1275 B.n768 B.n767 163.367
R1276 B.n768 B.n9 163.367
R1277 B.n772 B.n9 163.367
R1278 B.n773 B.n772 163.367
R1279 B.n774 B.n773 163.367
R1280 B.n774 B.n7 163.367
R1281 B.n778 B.n7 163.367
R1282 B.n779 B.n778 163.367
R1283 B.n780 B.n779 163.367
R1284 B.n780 B.n5 163.367
R1285 B.n784 B.n5 163.367
R1286 B.n785 B.n784 163.367
R1287 B.n786 B.n785 163.367
R1288 B.n786 B.n3 163.367
R1289 B.n790 B.n3 163.367
R1290 B.n791 B.n790 163.367
R1291 B.n204 B.n2 163.367
R1292 B.n205 B.n204 163.367
R1293 B.n206 B.n205 163.367
R1294 B.n206 B.n201 163.367
R1295 B.n210 B.n201 163.367
R1296 B.n211 B.n210 163.367
R1297 B.n212 B.n211 163.367
R1298 B.n212 B.n199 163.367
R1299 B.n216 B.n199 163.367
R1300 B.n217 B.n216 163.367
R1301 B.n218 B.n217 163.367
R1302 B.n218 B.n197 163.367
R1303 B.n222 B.n197 163.367
R1304 B.n223 B.n222 163.367
R1305 B.n224 B.n223 163.367
R1306 B.n224 B.n195 163.367
R1307 B.n228 B.n195 163.367
R1308 B.n229 B.n228 163.367
R1309 B.n230 B.n229 163.367
R1310 B.n230 B.n193 163.367
R1311 B.n234 B.n193 163.367
R1312 B.n235 B.n234 163.367
R1313 B.n236 B.n235 163.367
R1314 B.n236 B.n191 163.367
R1315 B.n240 B.n191 163.367
R1316 B.n241 B.n240 163.367
R1317 B.n242 B.n241 163.367
R1318 B.n242 B.n189 163.367
R1319 B.n246 B.n189 163.367
R1320 B.n247 B.n246 163.367
R1321 B.n248 B.n247 163.367
R1322 B.n248 B.n187 163.367
R1323 B.n252 B.n187 163.367
R1324 B.n253 B.n252 163.367
R1325 B.n254 B.n253 163.367
R1326 B.n254 B.n185 163.367
R1327 B.n258 B.n185 163.367
R1328 B.n259 B.n258 163.367
R1329 B.n260 B.n259 163.367
R1330 B.n260 B.n183 163.367
R1331 B.n264 B.n183 163.367
R1332 B.n265 B.n264 163.367
R1333 B.n266 B.n265 163.367
R1334 B.n266 B.n181 163.367
R1335 B.n270 B.n181 163.367
R1336 B.n271 B.n270 163.367
R1337 B.n272 B.n271 163.367
R1338 B.n272 B.n179 163.367
R1339 B.n276 B.n179 163.367
R1340 B.n277 B.n276 163.367
R1341 B.n278 B.n277 163.367
R1342 B.n278 B.n177 163.367
R1343 B.n282 B.n177 163.367
R1344 B.n283 B.n282 163.367
R1345 B.n284 B.n283 163.367
R1346 B.n284 B.n175 163.367
R1347 B.n288 B.n175 163.367
R1348 B.n289 B.n288 163.367
R1349 B.n290 B.n289 163.367
R1350 B.n290 B.n173 163.367
R1351 B.n294 B.n173 163.367
R1352 B.n295 B.n294 163.367
R1353 B.n296 B.n295 163.367
R1354 B.n296 B.n171 163.367
R1355 B.n300 B.n171 163.367
R1356 B.n301 B.n300 163.367
R1357 B.n302 B.n301 163.367
R1358 B.n302 B.n169 163.367
R1359 B.n306 B.n169 163.367
R1360 B.n307 B.n306 163.367
R1361 B.n308 B.n307 163.367
R1362 B.n308 B.n167 163.367
R1363 B.n312 B.n167 163.367
R1364 B.n313 B.n312 163.367
R1365 B.n314 B.n313 163.367
R1366 B.n314 B.n165 163.367
R1367 B.n318 B.n165 163.367
R1368 B.n157 B.n156 77.1884
R1369 B.n355 B.n354 77.1884
R1370 B.n57 B.n56 77.1884
R1371 B.n49 B.n48 77.1884
R1372 B.n340 B.n157 59.5399
R1373 B.n356 B.n355 59.5399
R1374 B.n638 B.n57 59.5399
R1375 B.n50 B.n49 59.5399
R1376 B.n675 B.n674 28.8785
R1377 B.n615 B.n64 28.8785
R1378 B.n380 B.n379 28.8785
R1379 B.n317 B.n164 28.8785
R1380 B B.n793 18.0485
R1381 B.n675 B.n40 10.6151
R1382 B.n679 B.n40 10.6151
R1383 B.n680 B.n679 10.6151
R1384 B.n681 B.n680 10.6151
R1385 B.n681 B.n38 10.6151
R1386 B.n685 B.n38 10.6151
R1387 B.n686 B.n685 10.6151
R1388 B.n687 B.n686 10.6151
R1389 B.n687 B.n36 10.6151
R1390 B.n691 B.n36 10.6151
R1391 B.n692 B.n691 10.6151
R1392 B.n693 B.n692 10.6151
R1393 B.n693 B.n34 10.6151
R1394 B.n697 B.n34 10.6151
R1395 B.n698 B.n697 10.6151
R1396 B.n699 B.n698 10.6151
R1397 B.n699 B.n32 10.6151
R1398 B.n703 B.n32 10.6151
R1399 B.n704 B.n703 10.6151
R1400 B.n705 B.n704 10.6151
R1401 B.n705 B.n30 10.6151
R1402 B.n709 B.n30 10.6151
R1403 B.n710 B.n709 10.6151
R1404 B.n711 B.n710 10.6151
R1405 B.n711 B.n28 10.6151
R1406 B.n715 B.n28 10.6151
R1407 B.n716 B.n715 10.6151
R1408 B.n717 B.n716 10.6151
R1409 B.n717 B.n26 10.6151
R1410 B.n721 B.n26 10.6151
R1411 B.n722 B.n721 10.6151
R1412 B.n723 B.n722 10.6151
R1413 B.n723 B.n24 10.6151
R1414 B.n727 B.n24 10.6151
R1415 B.n728 B.n727 10.6151
R1416 B.n729 B.n728 10.6151
R1417 B.n729 B.n22 10.6151
R1418 B.n733 B.n22 10.6151
R1419 B.n734 B.n733 10.6151
R1420 B.n735 B.n734 10.6151
R1421 B.n735 B.n20 10.6151
R1422 B.n739 B.n20 10.6151
R1423 B.n740 B.n739 10.6151
R1424 B.n741 B.n740 10.6151
R1425 B.n741 B.n18 10.6151
R1426 B.n745 B.n18 10.6151
R1427 B.n746 B.n745 10.6151
R1428 B.n747 B.n746 10.6151
R1429 B.n747 B.n16 10.6151
R1430 B.n751 B.n16 10.6151
R1431 B.n752 B.n751 10.6151
R1432 B.n753 B.n752 10.6151
R1433 B.n753 B.n14 10.6151
R1434 B.n757 B.n14 10.6151
R1435 B.n758 B.n757 10.6151
R1436 B.n759 B.n758 10.6151
R1437 B.n759 B.n12 10.6151
R1438 B.n763 B.n12 10.6151
R1439 B.n764 B.n763 10.6151
R1440 B.n765 B.n764 10.6151
R1441 B.n765 B.n10 10.6151
R1442 B.n769 B.n10 10.6151
R1443 B.n770 B.n769 10.6151
R1444 B.n771 B.n770 10.6151
R1445 B.n771 B.n8 10.6151
R1446 B.n775 B.n8 10.6151
R1447 B.n776 B.n775 10.6151
R1448 B.n777 B.n776 10.6151
R1449 B.n777 B.n6 10.6151
R1450 B.n781 B.n6 10.6151
R1451 B.n782 B.n781 10.6151
R1452 B.n783 B.n782 10.6151
R1453 B.n783 B.n4 10.6151
R1454 B.n787 B.n4 10.6151
R1455 B.n788 B.n787 10.6151
R1456 B.n789 B.n788 10.6151
R1457 B.n789 B.n0 10.6151
R1458 B.n674 B.n673 10.6151
R1459 B.n673 B.n42 10.6151
R1460 B.n669 B.n42 10.6151
R1461 B.n669 B.n668 10.6151
R1462 B.n668 B.n667 10.6151
R1463 B.n667 B.n44 10.6151
R1464 B.n663 B.n44 10.6151
R1465 B.n663 B.n662 10.6151
R1466 B.n662 B.n661 10.6151
R1467 B.n661 B.n46 10.6151
R1468 B.n657 B.n46 10.6151
R1469 B.n657 B.n656 10.6151
R1470 B.n656 B.n655 10.6151
R1471 B.n652 B.n651 10.6151
R1472 B.n651 B.n650 10.6151
R1473 B.n650 B.n52 10.6151
R1474 B.n646 B.n52 10.6151
R1475 B.n646 B.n645 10.6151
R1476 B.n645 B.n644 10.6151
R1477 B.n644 B.n54 10.6151
R1478 B.n640 B.n54 10.6151
R1479 B.n640 B.n639 10.6151
R1480 B.n637 B.n58 10.6151
R1481 B.n633 B.n58 10.6151
R1482 B.n633 B.n632 10.6151
R1483 B.n632 B.n631 10.6151
R1484 B.n631 B.n60 10.6151
R1485 B.n627 B.n60 10.6151
R1486 B.n627 B.n626 10.6151
R1487 B.n626 B.n625 10.6151
R1488 B.n625 B.n62 10.6151
R1489 B.n621 B.n62 10.6151
R1490 B.n621 B.n620 10.6151
R1491 B.n620 B.n619 10.6151
R1492 B.n619 B.n64 10.6151
R1493 B.n615 B.n614 10.6151
R1494 B.n614 B.n613 10.6151
R1495 B.n613 B.n66 10.6151
R1496 B.n609 B.n66 10.6151
R1497 B.n609 B.n608 10.6151
R1498 B.n608 B.n607 10.6151
R1499 B.n607 B.n68 10.6151
R1500 B.n603 B.n68 10.6151
R1501 B.n603 B.n602 10.6151
R1502 B.n602 B.n601 10.6151
R1503 B.n601 B.n70 10.6151
R1504 B.n597 B.n70 10.6151
R1505 B.n597 B.n596 10.6151
R1506 B.n596 B.n595 10.6151
R1507 B.n595 B.n72 10.6151
R1508 B.n591 B.n72 10.6151
R1509 B.n591 B.n590 10.6151
R1510 B.n590 B.n589 10.6151
R1511 B.n589 B.n74 10.6151
R1512 B.n585 B.n74 10.6151
R1513 B.n585 B.n584 10.6151
R1514 B.n584 B.n583 10.6151
R1515 B.n583 B.n76 10.6151
R1516 B.n579 B.n76 10.6151
R1517 B.n579 B.n578 10.6151
R1518 B.n578 B.n577 10.6151
R1519 B.n577 B.n78 10.6151
R1520 B.n573 B.n78 10.6151
R1521 B.n573 B.n572 10.6151
R1522 B.n572 B.n571 10.6151
R1523 B.n571 B.n80 10.6151
R1524 B.n567 B.n80 10.6151
R1525 B.n567 B.n566 10.6151
R1526 B.n566 B.n565 10.6151
R1527 B.n565 B.n82 10.6151
R1528 B.n561 B.n82 10.6151
R1529 B.n561 B.n560 10.6151
R1530 B.n560 B.n559 10.6151
R1531 B.n559 B.n84 10.6151
R1532 B.n555 B.n84 10.6151
R1533 B.n555 B.n554 10.6151
R1534 B.n554 B.n553 10.6151
R1535 B.n553 B.n86 10.6151
R1536 B.n549 B.n86 10.6151
R1537 B.n549 B.n548 10.6151
R1538 B.n548 B.n547 10.6151
R1539 B.n547 B.n88 10.6151
R1540 B.n543 B.n88 10.6151
R1541 B.n543 B.n542 10.6151
R1542 B.n542 B.n541 10.6151
R1543 B.n541 B.n90 10.6151
R1544 B.n537 B.n90 10.6151
R1545 B.n537 B.n536 10.6151
R1546 B.n536 B.n535 10.6151
R1547 B.n535 B.n92 10.6151
R1548 B.n531 B.n92 10.6151
R1549 B.n531 B.n530 10.6151
R1550 B.n530 B.n529 10.6151
R1551 B.n529 B.n94 10.6151
R1552 B.n525 B.n94 10.6151
R1553 B.n525 B.n524 10.6151
R1554 B.n524 B.n523 10.6151
R1555 B.n523 B.n96 10.6151
R1556 B.n519 B.n96 10.6151
R1557 B.n519 B.n518 10.6151
R1558 B.n518 B.n517 10.6151
R1559 B.n517 B.n98 10.6151
R1560 B.n513 B.n98 10.6151
R1561 B.n513 B.n512 10.6151
R1562 B.n512 B.n511 10.6151
R1563 B.n511 B.n100 10.6151
R1564 B.n507 B.n100 10.6151
R1565 B.n507 B.n506 10.6151
R1566 B.n506 B.n505 10.6151
R1567 B.n505 B.n102 10.6151
R1568 B.n501 B.n102 10.6151
R1569 B.n501 B.n500 10.6151
R1570 B.n500 B.n499 10.6151
R1571 B.n499 B.n104 10.6151
R1572 B.n495 B.n104 10.6151
R1573 B.n495 B.n494 10.6151
R1574 B.n494 B.n493 10.6151
R1575 B.n493 B.n106 10.6151
R1576 B.n489 B.n106 10.6151
R1577 B.n489 B.n488 10.6151
R1578 B.n488 B.n487 10.6151
R1579 B.n487 B.n108 10.6151
R1580 B.n483 B.n108 10.6151
R1581 B.n483 B.n482 10.6151
R1582 B.n482 B.n481 10.6151
R1583 B.n481 B.n110 10.6151
R1584 B.n477 B.n110 10.6151
R1585 B.n477 B.n476 10.6151
R1586 B.n476 B.n475 10.6151
R1587 B.n475 B.n112 10.6151
R1588 B.n471 B.n112 10.6151
R1589 B.n471 B.n470 10.6151
R1590 B.n470 B.n469 10.6151
R1591 B.n469 B.n114 10.6151
R1592 B.n465 B.n114 10.6151
R1593 B.n465 B.n464 10.6151
R1594 B.n464 B.n463 10.6151
R1595 B.n463 B.n116 10.6151
R1596 B.n459 B.n116 10.6151
R1597 B.n459 B.n458 10.6151
R1598 B.n458 B.n457 10.6151
R1599 B.n457 B.n118 10.6151
R1600 B.n453 B.n118 10.6151
R1601 B.n453 B.n452 10.6151
R1602 B.n452 B.n451 10.6151
R1603 B.n451 B.n120 10.6151
R1604 B.n447 B.n120 10.6151
R1605 B.n447 B.n446 10.6151
R1606 B.n446 B.n445 10.6151
R1607 B.n445 B.n122 10.6151
R1608 B.n441 B.n122 10.6151
R1609 B.n441 B.n440 10.6151
R1610 B.n440 B.n439 10.6151
R1611 B.n439 B.n124 10.6151
R1612 B.n435 B.n124 10.6151
R1613 B.n435 B.n434 10.6151
R1614 B.n434 B.n433 10.6151
R1615 B.n433 B.n126 10.6151
R1616 B.n429 B.n126 10.6151
R1617 B.n429 B.n428 10.6151
R1618 B.n428 B.n427 10.6151
R1619 B.n427 B.n128 10.6151
R1620 B.n423 B.n128 10.6151
R1621 B.n423 B.n422 10.6151
R1622 B.n422 B.n421 10.6151
R1623 B.n421 B.n130 10.6151
R1624 B.n417 B.n130 10.6151
R1625 B.n417 B.n416 10.6151
R1626 B.n416 B.n415 10.6151
R1627 B.n415 B.n132 10.6151
R1628 B.n411 B.n132 10.6151
R1629 B.n411 B.n410 10.6151
R1630 B.n410 B.n409 10.6151
R1631 B.n409 B.n134 10.6151
R1632 B.n405 B.n134 10.6151
R1633 B.n405 B.n404 10.6151
R1634 B.n404 B.n403 10.6151
R1635 B.n403 B.n136 10.6151
R1636 B.n399 B.n136 10.6151
R1637 B.n399 B.n398 10.6151
R1638 B.n398 B.n397 10.6151
R1639 B.n397 B.n138 10.6151
R1640 B.n393 B.n138 10.6151
R1641 B.n393 B.n392 10.6151
R1642 B.n392 B.n391 10.6151
R1643 B.n391 B.n140 10.6151
R1644 B.n387 B.n140 10.6151
R1645 B.n387 B.n386 10.6151
R1646 B.n386 B.n385 10.6151
R1647 B.n385 B.n142 10.6151
R1648 B.n381 B.n142 10.6151
R1649 B.n381 B.n380 10.6151
R1650 B.n203 B.n1 10.6151
R1651 B.n203 B.n202 10.6151
R1652 B.n207 B.n202 10.6151
R1653 B.n208 B.n207 10.6151
R1654 B.n209 B.n208 10.6151
R1655 B.n209 B.n200 10.6151
R1656 B.n213 B.n200 10.6151
R1657 B.n214 B.n213 10.6151
R1658 B.n215 B.n214 10.6151
R1659 B.n215 B.n198 10.6151
R1660 B.n219 B.n198 10.6151
R1661 B.n220 B.n219 10.6151
R1662 B.n221 B.n220 10.6151
R1663 B.n221 B.n196 10.6151
R1664 B.n225 B.n196 10.6151
R1665 B.n226 B.n225 10.6151
R1666 B.n227 B.n226 10.6151
R1667 B.n227 B.n194 10.6151
R1668 B.n231 B.n194 10.6151
R1669 B.n232 B.n231 10.6151
R1670 B.n233 B.n232 10.6151
R1671 B.n233 B.n192 10.6151
R1672 B.n237 B.n192 10.6151
R1673 B.n238 B.n237 10.6151
R1674 B.n239 B.n238 10.6151
R1675 B.n239 B.n190 10.6151
R1676 B.n243 B.n190 10.6151
R1677 B.n244 B.n243 10.6151
R1678 B.n245 B.n244 10.6151
R1679 B.n245 B.n188 10.6151
R1680 B.n249 B.n188 10.6151
R1681 B.n250 B.n249 10.6151
R1682 B.n251 B.n250 10.6151
R1683 B.n251 B.n186 10.6151
R1684 B.n255 B.n186 10.6151
R1685 B.n256 B.n255 10.6151
R1686 B.n257 B.n256 10.6151
R1687 B.n257 B.n184 10.6151
R1688 B.n261 B.n184 10.6151
R1689 B.n262 B.n261 10.6151
R1690 B.n263 B.n262 10.6151
R1691 B.n263 B.n182 10.6151
R1692 B.n267 B.n182 10.6151
R1693 B.n268 B.n267 10.6151
R1694 B.n269 B.n268 10.6151
R1695 B.n269 B.n180 10.6151
R1696 B.n273 B.n180 10.6151
R1697 B.n274 B.n273 10.6151
R1698 B.n275 B.n274 10.6151
R1699 B.n275 B.n178 10.6151
R1700 B.n279 B.n178 10.6151
R1701 B.n280 B.n279 10.6151
R1702 B.n281 B.n280 10.6151
R1703 B.n281 B.n176 10.6151
R1704 B.n285 B.n176 10.6151
R1705 B.n286 B.n285 10.6151
R1706 B.n287 B.n286 10.6151
R1707 B.n287 B.n174 10.6151
R1708 B.n291 B.n174 10.6151
R1709 B.n292 B.n291 10.6151
R1710 B.n293 B.n292 10.6151
R1711 B.n293 B.n172 10.6151
R1712 B.n297 B.n172 10.6151
R1713 B.n298 B.n297 10.6151
R1714 B.n299 B.n298 10.6151
R1715 B.n299 B.n170 10.6151
R1716 B.n303 B.n170 10.6151
R1717 B.n304 B.n303 10.6151
R1718 B.n305 B.n304 10.6151
R1719 B.n305 B.n168 10.6151
R1720 B.n309 B.n168 10.6151
R1721 B.n310 B.n309 10.6151
R1722 B.n311 B.n310 10.6151
R1723 B.n311 B.n166 10.6151
R1724 B.n315 B.n166 10.6151
R1725 B.n316 B.n315 10.6151
R1726 B.n317 B.n316 10.6151
R1727 B.n321 B.n164 10.6151
R1728 B.n322 B.n321 10.6151
R1729 B.n323 B.n322 10.6151
R1730 B.n323 B.n162 10.6151
R1731 B.n327 B.n162 10.6151
R1732 B.n328 B.n327 10.6151
R1733 B.n329 B.n328 10.6151
R1734 B.n329 B.n160 10.6151
R1735 B.n333 B.n160 10.6151
R1736 B.n334 B.n333 10.6151
R1737 B.n335 B.n334 10.6151
R1738 B.n335 B.n158 10.6151
R1739 B.n339 B.n158 10.6151
R1740 B.n342 B.n341 10.6151
R1741 B.n342 B.n154 10.6151
R1742 B.n346 B.n154 10.6151
R1743 B.n347 B.n346 10.6151
R1744 B.n348 B.n347 10.6151
R1745 B.n348 B.n152 10.6151
R1746 B.n352 B.n152 10.6151
R1747 B.n353 B.n352 10.6151
R1748 B.n357 B.n353 10.6151
R1749 B.n361 B.n150 10.6151
R1750 B.n362 B.n361 10.6151
R1751 B.n363 B.n362 10.6151
R1752 B.n363 B.n148 10.6151
R1753 B.n367 B.n148 10.6151
R1754 B.n368 B.n367 10.6151
R1755 B.n369 B.n368 10.6151
R1756 B.n369 B.n146 10.6151
R1757 B.n373 B.n146 10.6151
R1758 B.n374 B.n373 10.6151
R1759 B.n375 B.n374 10.6151
R1760 B.n375 B.n144 10.6151
R1761 B.n379 B.n144 10.6151
R1762 B.n655 B.n50 9.36635
R1763 B.n638 B.n637 9.36635
R1764 B.n340 B.n339 9.36635
R1765 B.n356 B.n150 9.36635
R1766 B.n793 B.n0 8.11757
R1767 B.n793 B.n1 8.11757
R1768 B.n652 B.n50 1.24928
R1769 B.n639 B.n638 1.24928
R1770 B.n341 B.n340 1.24928
R1771 B.n357 B.n356 1.24928
C0 VTAIL VN 4.82129f
C1 VN w_n5746_n1492# 12.448501f
C2 VDD2 VN 2.89727f
C3 VDD1 VTAIL 7.20644f
C4 VTAIL VP 4.83546f
C5 VDD1 w_n5746_n1492# 2.54427f
C6 w_n5746_n1492# VP 13.196799f
C7 VDD1 VDD2 2.85894f
C8 VDD2 VP 0.724373f
C9 VTAIL B 1.80668f
C10 VDD1 VN 0.161893f
C11 w_n5746_n1492# B 9.75085f
C12 VN VP 8.206019f
C13 VDD2 B 2.29051f
C14 VN B 1.47759f
C15 VDD1 VP 3.45533f
C16 VTAIL w_n5746_n1492# 2.066f
C17 VDD1 B 2.13137f
C18 B VP 2.74627f
C19 VDD2 VTAIL 7.26682f
C20 VDD2 w_n5746_n1492# 2.7418f
C21 VDD2 VSUBS 2.524359f
C22 VDD1 VSUBS 2.229961f
C23 VTAIL VSUBS 0.723386f
C24 VN VSUBS 9.587481f
C25 VP VSUBS 4.858373f
C26 B VSUBS 5.499282f
C27 w_n5746_n1492# VSUBS 0.108875p
C28 B.n0 VSUBS 0.011942f
C29 B.n1 VSUBS 0.011942f
C30 B.n2 VSUBS 0.017661f
C31 B.n3 VSUBS 0.013534f
C32 B.n4 VSUBS 0.013534f
C33 B.n5 VSUBS 0.013534f
C34 B.n6 VSUBS 0.013534f
C35 B.n7 VSUBS 0.013534f
C36 B.n8 VSUBS 0.013534f
C37 B.n9 VSUBS 0.013534f
C38 B.n10 VSUBS 0.013534f
C39 B.n11 VSUBS 0.013534f
C40 B.n12 VSUBS 0.013534f
C41 B.n13 VSUBS 0.013534f
C42 B.n14 VSUBS 0.013534f
C43 B.n15 VSUBS 0.013534f
C44 B.n16 VSUBS 0.013534f
C45 B.n17 VSUBS 0.013534f
C46 B.n18 VSUBS 0.013534f
C47 B.n19 VSUBS 0.013534f
C48 B.n20 VSUBS 0.013534f
C49 B.n21 VSUBS 0.013534f
C50 B.n22 VSUBS 0.013534f
C51 B.n23 VSUBS 0.013534f
C52 B.n24 VSUBS 0.013534f
C53 B.n25 VSUBS 0.013534f
C54 B.n26 VSUBS 0.013534f
C55 B.n27 VSUBS 0.013534f
C56 B.n28 VSUBS 0.013534f
C57 B.n29 VSUBS 0.013534f
C58 B.n30 VSUBS 0.013534f
C59 B.n31 VSUBS 0.013534f
C60 B.n32 VSUBS 0.013534f
C61 B.n33 VSUBS 0.013534f
C62 B.n34 VSUBS 0.013534f
C63 B.n35 VSUBS 0.013534f
C64 B.n36 VSUBS 0.013534f
C65 B.n37 VSUBS 0.013534f
C66 B.n38 VSUBS 0.013534f
C67 B.n39 VSUBS 0.013534f
C68 B.n40 VSUBS 0.013534f
C69 B.n41 VSUBS 0.030162f
C70 B.n42 VSUBS 0.013534f
C71 B.n43 VSUBS 0.013534f
C72 B.n44 VSUBS 0.013534f
C73 B.n45 VSUBS 0.013534f
C74 B.n46 VSUBS 0.013534f
C75 B.n47 VSUBS 0.013534f
C76 B.t1 VSUBS 0.078843f
C77 B.t2 VSUBS 0.116826f
C78 B.t0 VSUBS 0.909468f
C79 B.n48 VSUBS 0.204823f
C80 B.n49 VSUBS 0.168785f
C81 B.n50 VSUBS 0.031357f
C82 B.n51 VSUBS 0.013534f
C83 B.n52 VSUBS 0.013534f
C84 B.n53 VSUBS 0.013534f
C85 B.n54 VSUBS 0.013534f
C86 B.n55 VSUBS 0.013534f
C87 B.t4 VSUBS 0.078843f
C88 B.t5 VSUBS 0.116827f
C89 B.t3 VSUBS 0.909468f
C90 B.n56 VSUBS 0.204822f
C91 B.n57 VSUBS 0.168784f
C92 B.n58 VSUBS 0.013534f
C93 B.n59 VSUBS 0.013534f
C94 B.n60 VSUBS 0.013534f
C95 B.n61 VSUBS 0.013534f
C96 B.n62 VSUBS 0.013534f
C97 B.n63 VSUBS 0.013534f
C98 B.n64 VSUBS 0.030162f
C99 B.n65 VSUBS 0.013534f
C100 B.n66 VSUBS 0.013534f
C101 B.n67 VSUBS 0.013534f
C102 B.n68 VSUBS 0.013534f
C103 B.n69 VSUBS 0.013534f
C104 B.n70 VSUBS 0.013534f
C105 B.n71 VSUBS 0.013534f
C106 B.n72 VSUBS 0.013534f
C107 B.n73 VSUBS 0.013534f
C108 B.n74 VSUBS 0.013534f
C109 B.n75 VSUBS 0.013534f
C110 B.n76 VSUBS 0.013534f
C111 B.n77 VSUBS 0.013534f
C112 B.n78 VSUBS 0.013534f
C113 B.n79 VSUBS 0.013534f
C114 B.n80 VSUBS 0.013534f
C115 B.n81 VSUBS 0.013534f
C116 B.n82 VSUBS 0.013534f
C117 B.n83 VSUBS 0.013534f
C118 B.n84 VSUBS 0.013534f
C119 B.n85 VSUBS 0.013534f
C120 B.n86 VSUBS 0.013534f
C121 B.n87 VSUBS 0.013534f
C122 B.n88 VSUBS 0.013534f
C123 B.n89 VSUBS 0.013534f
C124 B.n90 VSUBS 0.013534f
C125 B.n91 VSUBS 0.013534f
C126 B.n92 VSUBS 0.013534f
C127 B.n93 VSUBS 0.013534f
C128 B.n94 VSUBS 0.013534f
C129 B.n95 VSUBS 0.013534f
C130 B.n96 VSUBS 0.013534f
C131 B.n97 VSUBS 0.013534f
C132 B.n98 VSUBS 0.013534f
C133 B.n99 VSUBS 0.013534f
C134 B.n100 VSUBS 0.013534f
C135 B.n101 VSUBS 0.013534f
C136 B.n102 VSUBS 0.013534f
C137 B.n103 VSUBS 0.013534f
C138 B.n104 VSUBS 0.013534f
C139 B.n105 VSUBS 0.013534f
C140 B.n106 VSUBS 0.013534f
C141 B.n107 VSUBS 0.013534f
C142 B.n108 VSUBS 0.013534f
C143 B.n109 VSUBS 0.013534f
C144 B.n110 VSUBS 0.013534f
C145 B.n111 VSUBS 0.013534f
C146 B.n112 VSUBS 0.013534f
C147 B.n113 VSUBS 0.013534f
C148 B.n114 VSUBS 0.013534f
C149 B.n115 VSUBS 0.013534f
C150 B.n116 VSUBS 0.013534f
C151 B.n117 VSUBS 0.013534f
C152 B.n118 VSUBS 0.013534f
C153 B.n119 VSUBS 0.013534f
C154 B.n120 VSUBS 0.013534f
C155 B.n121 VSUBS 0.013534f
C156 B.n122 VSUBS 0.013534f
C157 B.n123 VSUBS 0.013534f
C158 B.n124 VSUBS 0.013534f
C159 B.n125 VSUBS 0.013534f
C160 B.n126 VSUBS 0.013534f
C161 B.n127 VSUBS 0.013534f
C162 B.n128 VSUBS 0.013534f
C163 B.n129 VSUBS 0.013534f
C164 B.n130 VSUBS 0.013534f
C165 B.n131 VSUBS 0.013534f
C166 B.n132 VSUBS 0.013534f
C167 B.n133 VSUBS 0.013534f
C168 B.n134 VSUBS 0.013534f
C169 B.n135 VSUBS 0.013534f
C170 B.n136 VSUBS 0.013534f
C171 B.n137 VSUBS 0.013534f
C172 B.n138 VSUBS 0.013534f
C173 B.n139 VSUBS 0.013534f
C174 B.n140 VSUBS 0.013534f
C175 B.n141 VSUBS 0.013534f
C176 B.n142 VSUBS 0.013534f
C177 B.n143 VSUBS 0.028354f
C178 B.n144 VSUBS 0.013534f
C179 B.n145 VSUBS 0.013534f
C180 B.n146 VSUBS 0.013534f
C181 B.n147 VSUBS 0.013534f
C182 B.n148 VSUBS 0.013534f
C183 B.n149 VSUBS 0.013534f
C184 B.n150 VSUBS 0.012738f
C185 B.n151 VSUBS 0.013534f
C186 B.n152 VSUBS 0.013534f
C187 B.n153 VSUBS 0.013534f
C188 B.n154 VSUBS 0.013534f
C189 B.n155 VSUBS 0.013534f
C190 B.t8 VSUBS 0.078843f
C191 B.t7 VSUBS 0.116826f
C192 B.t6 VSUBS 0.909468f
C193 B.n156 VSUBS 0.204823f
C194 B.n157 VSUBS 0.168785f
C195 B.n158 VSUBS 0.013534f
C196 B.n159 VSUBS 0.013534f
C197 B.n160 VSUBS 0.013534f
C198 B.n161 VSUBS 0.013534f
C199 B.n162 VSUBS 0.013534f
C200 B.n163 VSUBS 0.013534f
C201 B.n164 VSUBS 0.030162f
C202 B.n165 VSUBS 0.013534f
C203 B.n166 VSUBS 0.013534f
C204 B.n167 VSUBS 0.013534f
C205 B.n168 VSUBS 0.013534f
C206 B.n169 VSUBS 0.013534f
C207 B.n170 VSUBS 0.013534f
C208 B.n171 VSUBS 0.013534f
C209 B.n172 VSUBS 0.013534f
C210 B.n173 VSUBS 0.013534f
C211 B.n174 VSUBS 0.013534f
C212 B.n175 VSUBS 0.013534f
C213 B.n176 VSUBS 0.013534f
C214 B.n177 VSUBS 0.013534f
C215 B.n178 VSUBS 0.013534f
C216 B.n179 VSUBS 0.013534f
C217 B.n180 VSUBS 0.013534f
C218 B.n181 VSUBS 0.013534f
C219 B.n182 VSUBS 0.013534f
C220 B.n183 VSUBS 0.013534f
C221 B.n184 VSUBS 0.013534f
C222 B.n185 VSUBS 0.013534f
C223 B.n186 VSUBS 0.013534f
C224 B.n187 VSUBS 0.013534f
C225 B.n188 VSUBS 0.013534f
C226 B.n189 VSUBS 0.013534f
C227 B.n190 VSUBS 0.013534f
C228 B.n191 VSUBS 0.013534f
C229 B.n192 VSUBS 0.013534f
C230 B.n193 VSUBS 0.013534f
C231 B.n194 VSUBS 0.013534f
C232 B.n195 VSUBS 0.013534f
C233 B.n196 VSUBS 0.013534f
C234 B.n197 VSUBS 0.013534f
C235 B.n198 VSUBS 0.013534f
C236 B.n199 VSUBS 0.013534f
C237 B.n200 VSUBS 0.013534f
C238 B.n201 VSUBS 0.013534f
C239 B.n202 VSUBS 0.013534f
C240 B.n203 VSUBS 0.013534f
C241 B.n204 VSUBS 0.013534f
C242 B.n205 VSUBS 0.013534f
C243 B.n206 VSUBS 0.013534f
C244 B.n207 VSUBS 0.013534f
C245 B.n208 VSUBS 0.013534f
C246 B.n209 VSUBS 0.013534f
C247 B.n210 VSUBS 0.013534f
C248 B.n211 VSUBS 0.013534f
C249 B.n212 VSUBS 0.013534f
C250 B.n213 VSUBS 0.013534f
C251 B.n214 VSUBS 0.013534f
C252 B.n215 VSUBS 0.013534f
C253 B.n216 VSUBS 0.013534f
C254 B.n217 VSUBS 0.013534f
C255 B.n218 VSUBS 0.013534f
C256 B.n219 VSUBS 0.013534f
C257 B.n220 VSUBS 0.013534f
C258 B.n221 VSUBS 0.013534f
C259 B.n222 VSUBS 0.013534f
C260 B.n223 VSUBS 0.013534f
C261 B.n224 VSUBS 0.013534f
C262 B.n225 VSUBS 0.013534f
C263 B.n226 VSUBS 0.013534f
C264 B.n227 VSUBS 0.013534f
C265 B.n228 VSUBS 0.013534f
C266 B.n229 VSUBS 0.013534f
C267 B.n230 VSUBS 0.013534f
C268 B.n231 VSUBS 0.013534f
C269 B.n232 VSUBS 0.013534f
C270 B.n233 VSUBS 0.013534f
C271 B.n234 VSUBS 0.013534f
C272 B.n235 VSUBS 0.013534f
C273 B.n236 VSUBS 0.013534f
C274 B.n237 VSUBS 0.013534f
C275 B.n238 VSUBS 0.013534f
C276 B.n239 VSUBS 0.013534f
C277 B.n240 VSUBS 0.013534f
C278 B.n241 VSUBS 0.013534f
C279 B.n242 VSUBS 0.013534f
C280 B.n243 VSUBS 0.013534f
C281 B.n244 VSUBS 0.013534f
C282 B.n245 VSUBS 0.013534f
C283 B.n246 VSUBS 0.013534f
C284 B.n247 VSUBS 0.013534f
C285 B.n248 VSUBS 0.013534f
C286 B.n249 VSUBS 0.013534f
C287 B.n250 VSUBS 0.013534f
C288 B.n251 VSUBS 0.013534f
C289 B.n252 VSUBS 0.013534f
C290 B.n253 VSUBS 0.013534f
C291 B.n254 VSUBS 0.013534f
C292 B.n255 VSUBS 0.013534f
C293 B.n256 VSUBS 0.013534f
C294 B.n257 VSUBS 0.013534f
C295 B.n258 VSUBS 0.013534f
C296 B.n259 VSUBS 0.013534f
C297 B.n260 VSUBS 0.013534f
C298 B.n261 VSUBS 0.013534f
C299 B.n262 VSUBS 0.013534f
C300 B.n263 VSUBS 0.013534f
C301 B.n264 VSUBS 0.013534f
C302 B.n265 VSUBS 0.013534f
C303 B.n266 VSUBS 0.013534f
C304 B.n267 VSUBS 0.013534f
C305 B.n268 VSUBS 0.013534f
C306 B.n269 VSUBS 0.013534f
C307 B.n270 VSUBS 0.013534f
C308 B.n271 VSUBS 0.013534f
C309 B.n272 VSUBS 0.013534f
C310 B.n273 VSUBS 0.013534f
C311 B.n274 VSUBS 0.013534f
C312 B.n275 VSUBS 0.013534f
C313 B.n276 VSUBS 0.013534f
C314 B.n277 VSUBS 0.013534f
C315 B.n278 VSUBS 0.013534f
C316 B.n279 VSUBS 0.013534f
C317 B.n280 VSUBS 0.013534f
C318 B.n281 VSUBS 0.013534f
C319 B.n282 VSUBS 0.013534f
C320 B.n283 VSUBS 0.013534f
C321 B.n284 VSUBS 0.013534f
C322 B.n285 VSUBS 0.013534f
C323 B.n286 VSUBS 0.013534f
C324 B.n287 VSUBS 0.013534f
C325 B.n288 VSUBS 0.013534f
C326 B.n289 VSUBS 0.013534f
C327 B.n290 VSUBS 0.013534f
C328 B.n291 VSUBS 0.013534f
C329 B.n292 VSUBS 0.013534f
C330 B.n293 VSUBS 0.013534f
C331 B.n294 VSUBS 0.013534f
C332 B.n295 VSUBS 0.013534f
C333 B.n296 VSUBS 0.013534f
C334 B.n297 VSUBS 0.013534f
C335 B.n298 VSUBS 0.013534f
C336 B.n299 VSUBS 0.013534f
C337 B.n300 VSUBS 0.013534f
C338 B.n301 VSUBS 0.013534f
C339 B.n302 VSUBS 0.013534f
C340 B.n303 VSUBS 0.013534f
C341 B.n304 VSUBS 0.013534f
C342 B.n305 VSUBS 0.013534f
C343 B.n306 VSUBS 0.013534f
C344 B.n307 VSUBS 0.013534f
C345 B.n308 VSUBS 0.013534f
C346 B.n309 VSUBS 0.013534f
C347 B.n310 VSUBS 0.013534f
C348 B.n311 VSUBS 0.013534f
C349 B.n312 VSUBS 0.013534f
C350 B.n313 VSUBS 0.013534f
C351 B.n314 VSUBS 0.013534f
C352 B.n315 VSUBS 0.013534f
C353 B.n316 VSUBS 0.013534f
C354 B.n317 VSUBS 0.028354f
C355 B.n318 VSUBS 0.028354f
C356 B.n319 VSUBS 0.030162f
C357 B.n320 VSUBS 0.013534f
C358 B.n321 VSUBS 0.013534f
C359 B.n322 VSUBS 0.013534f
C360 B.n323 VSUBS 0.013534f
C361 B.n324 VSUBS 0.013534f
C362 B.n325 VSUBS 0.013534f
C363 B.n326 VSUBS 0.013534f
C364 B.n327 VSUBS 0.013534f
C365 B.n328 VSUBS 0.013534f
C366 B.n329 VSUBS 0.013534f
C367 B.n330 VSUBS 0.013534f
C368 B.n331 VSUBS 0.013534f
C369 B.n332 VSUBS 0.013534f
C370 B.n333 VSUBS 0.013534f
C371 B.n334 VSUBS 0.013534f
C372 B.n335 VSUBS 0.013534f
C373 B.n336 VSUBS 0.013534f
C374 B.n337 VSUBS 0.013534f
C375 B.n338 VSUBS 0.013534f
C376 B.n339 VSUBS 0.012738f
C377 B.n340 VSUBS 0.031357f
C378 B.n341 VSUBS 0.007563f
C379 B.n342 VSUBS 0.013534f
C380 B.n343 VSUBS 0.013534f
C381 B.n344 VSUBS 0.013534f
C382 B.n345 VSUBS 0.013534f
C383 B.n346 VSUBS 0.013534f
C384 B.n347 VSUBS 0.013534f
C385 B.n348 VSUBS 0.013534f
C386 B.n349 VSUBS 0.013534f
C387 B.n350 VSUBS 0.013534f
C388 B.n351 VSUBS 0.013534f
C389 B.n352 VSUBS 0.013534f
C390 B.n353 VSUBS 0.013534f
C391 B.t11 VSUBS 0.078843f
C392 B.t10 VSUBS 0.116827f
C393 B.t9 VSUBS 0.909468f
C394 B.n354 VSUBS 0.204822f
C395 B.n355 VSUBS 0.168784f
C396 B.n356 VSUBS 0.031357f
C397 B.n357 VSUBS 0.007563f
C398 B.n358 VSUBS 0.013534f
C399 B.n359 VSUBS 0.013534f
C400 B.n360 VSUBS 0.013534f
C401 B.n361 VSUBS 0.013534f
C402 B.n362 VSUBS 0.013534f
C403 B.n363 VSUBS 0.013534f
C404 B.n364 VSUBS 0.013534f
C405 B.n365 VSUBS 0.013534f
C406 B.n366 VSUBS 0.013534f
C407 B.n367 VSUBS 0.013534f
C408 B.n368 VSUBS 0.013534f
C409 B.n369 VSUBS 0.013534f
C410 B.n370 VSUBS 0.013534f
C411 B.n371 VSUBS 0.013534f
C412 B.n372 VSUBS 0.013534f
C413 B.n373 VSUBS 0.013534f
C414 B.n374 VSUBS 0.013534f
C415 B.n375 VSUBS 0.013534f
C416 B.n376 VSUBS 0.013534f
C417 B.n377 VSUBS 0.013534f
C418 B.n378 VSUBS 0.030162f
C419 B.n379 VSUBS 0.028354f
C420 B.n380 VSUBS 0.030162f
C421 B.n381 VSUBS 0.013534f
C422 B.n382 VSUBS 0.013534f
C423 B.n383 VSUBS 0.013534f
C424 B.n384 VSUBS 0.013534f
C425 B.n385 VSUBS 0.013534f
C426 B.n386 VSUBS 0.013534f
C427 B.n387 VSUBS 0.013534f
C428 B.n388 VSUBS 0.013534f
C429 B.n389 VSUBS 0.013534f
C430 B.n390 VSUBS 0.013534f
C431 B.n391 VSUBS 0.013534f
C432 B.n392 VSUBS 0.013534f
C433 B.n393 VSUBS 0.013534f
C434 B.n394 VSUBS 0.013534f
C435 B.n395 VSUBS 0.013534f
C436 B.n396 VSUBS 0.013534f
C437 B.n397 VSUBS 0.013534f
C438 B.n398 VSUBS 0.013534f
C439 B.n399 VSUBS 0.013534f
C440 B.n400 VSUBS 0.013534f
C441 B.n401 VSUBS 0.013534f
C442 B.n402 VSUBS 0.013534f
C443 B.n403 VSUBS 0.013534f
C444 B.n404 VSUBS 0.013534f
C445 B.n405 VSUBS 0.013534f
C446 B.n406 VSUBS 0.013534f
C447 B.n407 VSUBS 0.013534f
C448 B.n408 VSUBS 0.013534f
C449 B.n409 VSUBS 0.013534f
C450 B.n410 VSUBS 0.013534f
C451 B.n411 VSUBS 0.013534f
C452 B.n412 VSUBS 0.013534f
C453 B.n413 VSUBS 0.013534f
C454 B.n414 VSUBS 0.013534f
C455 B.n415 VSUBS 0.013534f
C456 B.n416 VSUBS 0.013534f
C457 B.n417 VSUBS 0.013534f
C458 B.n418 VSUBS 0.013534f
C459 B.n419 VSUBS 0.013534f
C460 B.n420 VSUBS 0.013534f
C461 B.n421 VSUBS 0.013534f
C462 B.n422 VSUBS 0.013534f
C463 B.n423 VSUBS 0.013534f
C464 B.n424 VSUBS 0.013534f
C465 B.n425 VSUBS 0.013534f
C466 B.n426 VSUBS 0.013534f
C467 B.n427 VSUBS 0.013534f
C468 B.n428 VSUBS 0.013534f
C469 B.n429 VSUBS 0.013534f
C470 B.n430 VSUBS 0.013534f
C471 B.n431 VSUBS 0.013534f
C472 B.n432 VSUBS 0.013534f
C473 B.n433 VSUBS 0.013534f
C474 B.n434 VSUBS 0.013534f
C475 B.n435 VSUBS 0.013534f
C476 B.n436 VSUBS 0.013534f
C477 B.n437 VSUBS 0.013534f
C478 B.n438 VSUBS 0.013534f
C479 B.n439 VSUBS 0.013534f
C480 B.n440 VSUBS 0.013534f
C481 B.n441 VSUBS 0.013534f
C482 B.n442 VSUBS 0.013534f
C483 B.n443 VSUBS 0.013534f
C484 B.n444 VSUBS 0.013534f
C485 B.n445 VSUBS 0.013534f
C486 B.n446 VSUBS 0.013534f
C487 B.n447 VSUBS 0.013534f
C488 B.n448 VSUBS 0.013534f
C489 B.n449 VSUBS 0.013534f
C490 B.n450 VSUBS 0.013534f
C491 B.n451 VSUBS 0.013534f
C492 B.n452 VSUBS 0.013534f
C493 B.n453 VSUBS 0.013534f
C494 B.n454 VSUBS 0.013534f
C495 B.n455 VSUBS 0.013534f
C496 B.n456 VSUBS 0.013534f
C497 B.n457 VSUBS 0.013534f
C498 B.n458 VSUBS 0.013534f
C499 B.n459 VSUBS 0.013534f
C500 B.n460 VSUBS 0.013534f
C501 B.n461 VSUBS 0.013534f
C502 B.n462 VSUBS 0.013534f
C503 B.n463 VSUBS 0.013534f
C504 B.n464 VSUBS 0.013534f
C505 B.n465 VSUBS 0.013534f
C506 B.n466 VSUBS 0.013534f
C507 B.n467 VSUBS 0.013534f
C508 B.n468 VSUBS 0.013534f
C509 B.n469 VSUBS 0.013534f
C510 B.n470 VSUBS 0.013534f
C511 B.n471 VSUBS 0.013534f
C512 B.n472 VSUBS 0.013534f
C513 B.n473 VSUBS 0.013534f
C514 B.n474 VSUBS 0.013534f
C515 B.n475 VSUBS 0.013534f
C516 B.n476 VSUBS 0.013534f
C517 B.n477 VSUBS 0.013534f
C518 B.n478 VSUBS 0.013534f
C519 B.n479 VSUBS 0.013534f
C520 B.n480 VSUBS 0.013534f
C521 B.n481 VSUBS 0.013534f
C522 B.n482 VSUBS 0.013534f
C523 B.n483 VSUBS 0.013534f
C524 B.n484 VSUBS 0.013534f
C525 B.n485 VSUBS 0.013534f
C526 B.n486 VSUBS 0.013534f
C527 B.n487 VSUBS 0.013534f
C528 B.n488 VSUBS 0.013534f
C529 B.n489 VSUBS 0.013534f
C530 B.n490 VSUBS 0.013534f
C531 B.n491 VSUBS 0.013534f
C532 B.n492 VSUBS 0.013534f
C533 B.n493 VSUBS 0.013534f
C534 B.n494 VSUBS 0.013534f
C535 B.n495 VSUBS 0.013534f
C536 B.n496 VSUBS 0.013534f
C537 B.n497 VSUBS 0.013534f
C538 B.n498 VSUBS 0.013534f
C539 B.n499 VSUBS 0.013534f
C540 B.n500 VSUBS 0.013534f
C541 B.n501 VSUBS 0.013534f
C542 B.n502 VSUBS 0.013534f
C543 B.n503 VSUBS 0.013534f
C544 B.n504 VSUBS 0.013534f
C545 B.n505 VSUBS 0.013534f
C546 B.n506 VSUBS 0.013534f
C547 B.n507 VSUBS 0.013534f
C548 B.n508 VSUBS 0.013534f
C549 B.n509 VSUBS 0.013534f
C550 B.n510 VSUBS 0.013534f
C551 B.n511 VSUBS 0.013534f
C552 B.n512 VSUBS 0.013534f
C553 B.n513 VSUBS 0.013534f
C554 B.n514 VSUBS 0.013534f
C555 B.n515 VSUBS 0.013534f
C556 B.n516 VSUBS 0.013534f
C557 B.n517 VSUBS 0.013534f
C558 B.n518 VSUBS 0.013534f
C559 B.n519 VSUBS 0.013534f
C560 B.n520 VSUBS 0.013534f
C561 B.n521 VSUBS 0.013534f
C562 B.n522 VSUBS 0.013534f
C563 B.n523 VSUBS 0.013534f
C564 B.n524 VSUBS 0.013534f
C565 B.n525 VSUBS 0.013534f
C566 B.n526 VSUBS 0.013534f
C567 B.n527 VSUBS 0.013534f
C568 B.n528 VSUBS 0.013534f
C569 B.n529 VSUBS 0.013534f
C570 B.n530 VSUBS 0.013534f
C571 B.n531 VSUBS 0.013534f
C572 B.n532 VSUBS 0.013534f
C573 B.n533 VSUBS 0.013534f
C574 B.n534 VSUBS 0.013534f
C575 B.n535 VSUBS 0.013534f
C576 B.n536 VSUBS 0.013534f
C577 B.n537 VSUBS 0.013534f
C578 B.n538 VSUBS 0.013534f
C579 B.n539 VSUBS 0.013534f
C580 B.n540 VSUBS 0.013534f
C581 B.n541 VSUBS 0.013534f
C582 B.n542 VSUBS 0.013534f
C583 B.n543 VSUBS 0.013534f
C584 B.n544 VSUBS 0.013534f
C585 B.n545 VSUBS 0.013534f
C586 B.n546 VSUBS 0.013534f
C587 B.n547 VSUBS 0.013534f
C588 B.n548 VSUBS 0.013534f
C589 B.n549 VSUBS 0.013534f
C590 B.n550 VSUBS 0.013534f
C591 B.n551 VSUBS 0.013534f
C592 B.n552 VSUBS 0.013534f
C593 B.n553 VSUBS 0.013534f
C594 B.n554 VSUBS 0.013534f
C595 B.n555 VSUBS 0.013534f
C596 B.n556 VSUBS 0.013534f
C597 B.n557 VSUBS 0.013534f
C598 B.n558 VSUBS 0.013534f
C599 B.n559 VSUBS 0.013534f
C600 B.n560 VSUBS 0.013534f
C601 B.n561 VSUBS 0.013534f
C602 B.n562 VSUBS 0.013534f
C603 B.n563 VSUBS 0.013534f
C604 B.n564 VSUBS 0.013534f
C605 B.n565 VSUBS 0.013534f
C606 B.n566 VSUBS 0.013534f
C607 B.n567 VSUBS 0.013534f
C608 B.n568 VSUBS 0.013534f
C609 B.n569 VSUBS 0.013534f
C610 B.n570 VSUBS 0.013534f
C611 B.n571 VSUBS 0.013534f
C612 B.n572 VSUBS 0.013534f
C613 B.n573 VSUBS 0.013534f
C614 B.n574 VSUBS 0.013534f
C615 B.n575 VSUBS 0.013534f
C616 B.n576 VSUBS 0.013534f
C617 B.n577 VSUBS 0.013534f
C618 B.n578 VSUBS 0.013534f
C619 B.n579 VSUBS 0.013534f
C620 B.n580 VSUBS 0.013534f
C621 B.n581 VSUBS 0.013534f
C622 B.n582 VSUBS 0.013534f
C623 B.n583 VSUBS 0.013534f
C624 B.n584 VSUBS 0.013534f
C625 B.n585 VSUBS 0.013534f
C626 B.n586 VSUBS 0.013534f
C627 B.n587 VSUBS 0.013534f
C628 B.n588 VSUBS 0.013534f
C629 B.n589 VSUBS 0.013534f
C630 B.n590 VSUBS 0.013534f
C631 B.n591 VSUBS 0.013534f
C632 B.n592 VSUBS 0.013534f
C633 B.n593 VSUBS 0.013534f
C634 B.n594 VSUBS 0.013534f
C635 B.n595 VSUBS 0.013534f
C636 B.n596 VSUBS 0.013534f
C637 B.n597 VSUBS 0.013534f
C638 B.n598 VSUBS 0.013534f
C639 B.n599 VSUBS 0.013534f
C640 B.n600 VSUBS 0.013534f
C641 B.n601 VSUBS 0.013534f
C642 B.n602 VSUBS 0.013534f
C643 B.n603 VSUBS 0.013534f
C644 B.n604 VSUBS 0.013534f
C645 B.n605 VSUBS 0.013534f
C646 B.n606 VSUBS 0.013534f
C647 B.n607 VSUBS 0.013534f
C648 B.n608 VSUBS 0.013534f
C649 B.n609 VSUBS 0.013534f
C650 B.n610 VSUBS 0.013534f
C651 B.n611 VSUBS 0.013534f
C652 B.n612 VSUBS 0.013534f
C653 B.n613 VSUBS 0.013534f
C654 B.n614 VSUBS 0.013534f
C655 B.n615 VSUBS 0.028354f
C656 B.n616 VSUBS 0.028354f
C657 B.n617 VSUBS 0.030162f
C658 B.n618 VSUBS 0.013534f
C659 B.n619 VSUBS 0.013534f
C660 B.n620 VSUBS 0.013534f
C661 B.n621 VSUBS 0.013534f
C662 B.n622 VSUBS 0.013534f
C663 B.n623 VSUBS 0.013534f
C664 B.n624 VSUBS 0.013534f
C665 B.n625 VSUBS 0.013534f
C666 B.n626 VSUBS 0.013534f
C667 B.n627 VSUBS 0.013534f
C668 B.n628 VSUBS 0.013534f
C669 B.n629 VSUBS 0.013534f
C670 B.n630 VSUBS 0.013534f
C671 B.n631 VSUBS 0.013534f
C672 B.n632 VSUBS 0.013534f
C673 B.n633 VSUBS 0.013534f
C674 B.n634 VSUBS 0.013534f
C675 B.n635 VSUBS 0.013534f
C676 B.n636 VSUBS 0.013534f
C677 B.n637 VSUBS 0.012738f
C678 B.n638 VSUBS 0.031357f
C679 B.n639 VSUBS 0.007563f
C680 B.n640 VSUBS 0.013534f
C681 B.n641 VSUBS 0.013534f
C682 B.n642 VSUBS 0.013534f
C683 B.n643 VSUBS 0.013534f
C684 B.n644 VSUBS 0.013534f
C685 B.n645 VSUBS 0.013534f
C686 B.n646 VSUBS 0.013534f
C687 B.n647 VSUBS 0.013534f
C688 B.n648 VSUBS 0.013534f
C689 B.n649 VSUBS 0.013534f
C690 B.n650 VSUBS 0.013534f
C691 B.n651 VSUBS 0.013534f
C692 B.n652 VSUBS 0.007563f
C693 B.n653 VSUBS 0.013534f
C694 B.n654 VSUBS 0.013534f
C695 B.n655 VSUBS 0.012738f
C696 B.n656 VSUBS 0.013534f
C697 B.n657 VSUBS 0.013534f
C698 B.n658 VSUBS 0.013534f
C699 B.n659 VSUBS 0.013534f
C700 B.n660 VSUBS 0.013534f
C701 B.n661 VSUBS 0.013534f
C702 B.n662 VSUBS 0.013534f
C703 B.n663 VSUBS 0.013534f
C704 B.n664 VSUBS 0.013534f
C705 B.n665 VSUBS 0.013534f
C706 B.n666 VSUBS 0.013534f
C707 B.n667 VSUBS 0.013534f
C708 B.n668 VSUBS 0.013534f
C709 B.n669 VSUBS 0.013534f
C710 B.n670 VSUBS 0.013534f
C711 B.n671 VSUBS 0.013534f
C712 B.n672 VSUBS 0.013534f
C713 B.n673 VSUBS 0.013534f
C714 B.n674 VSUBS 0.030162f
C715 B.n675 VSUBS 0.028354f
C716 B.n676 VSUBS 0.028354f
C717 B.n677 VSUBS 0.013534f
C718 B.n678 VSUBS 0.013534f
C719 B.n679 VSUBS 0.013534f
C720 B.n680 VSUBS 0.013534f
C721 B.n681 VSUBS 0.013534f
C722 B.n682 VSUBS 0.013534f
C723 B.n683 VSUBS 0.013534f
C724 B.n684 VSUBS 0.013534f
C725 B.n685 VSUBS 0.013534f
C726 B.n686 VSUBS 0.013534f
C727 B.n687 VSUBS 0.013534f
C728 B.n688 VSUBS 0.013534f
C729 B.n689 VSUBS 0.013534f
C730 B.n690 VSUBS 0.013534f
C731 B.n691 VSUBS 0.013534f
C732 B.n692 VSUBS 0.013534f
C733 B.n693 VSUBS 0.013534f
C734 B.n694 VSUBS 0.013534f
C735 B.n695 VSUBS 0.013534f
C736 B.n696 VSUBS 0.013534f
C737 B.n697 VSUBS 0.013534f
C738 B.n698 VSUBS 0.013534f
C739 B.n699 VSUBS 0.013534f
C740 B.n700 VSUBS 0.013534f
C741 B.n701 VSUBS 0.013534f
C742 B.n702 VSUBS 0.013534f
C743 B.n703 VSUBS 0.013534f
C744 B.n704 VSUBS 0.013534f
C745 B.n705 VSUBS 0.013534f
C746 B.n706 VSUBS 0.013534f
C747 B.n707 VSUBS 0.013534f
C748 B.n708 VSUBS 0.013534f
C749 B.n709 VSUBS 0.013534f
C750 B.n710 VSUBS 0.013534f
C751 B.n711 VSUBS 0.013534f
C752 B.n712 VSUBS 0.013534f
C753 B.n713 VSUBS 0.013534f
C754 B.n714 VSUBS 0.013534f
C755 B.n715 VSUBS 0.013534f
C756 B.n716 VSUBS 0.013534f
C757 B.n717 VSUBS 0.013534f
C758 B.n718 VSUBS 0.013534f
C759 B.n719 VSUBS 0.013534f
C760 B.n720 VSUBS 0.013534f
C761 B.n721 VSUBS 0.013534f
C762 B.n722 VSUBS 0.013534f
C763 B.n723 VSUBS 0.013534f
C764 B.n724 VSUBS 0.013534f
C765 B.n725 VSUBS 0.013534f
C766 B.n726 VSUBS 0.013534f
C767 B.n727 VSUBS 0.013534f
C768 B.n728 VSUBS 0.013534f
C769 B.n729 VSUBS 0.013534f
C770 B.n730 VSUBS 0.013534f
C771 B.n731 VSUBS 0.013534f
C772 B.n732 VSUBS 0.013534f
C773 B.n733 VSUBS 0.013534f
C774 B.n734 VSUBS 0.013534f
C775 B.n735 VSUBS 0.013534f
C776 B.n736 VSUBS 0.013534f
C777 B.n737 VSUBS 0.013534f
C778 B.n738 VSUBS 0.013534f
C779 B.n739 VSUBS 0.013534f
C780 B.n740 VSUBS 0.013534f
C781 B.n741 VSUBS 0.013534f
C782 B.n742 VSUBS 0.013534f
C783 B.n743 VSUBS 0.013534f
C784 B.n744 VSUBS 0.013534f
C785 B.n745 VSUBS 0.013534f
C786 B.n746 VSUBS 0.013534f
C787 B.n747 VSUBS 0.013534f
C788 B.n748 VSUBS 0.013534f
C789 B.n749 VSUBS 0.013534f
C790 B.n750 VSUBS 0.013534f
C791 B.n751 VSUBS 0.013534f
C792 B.n752 VSUBS 0.013534f
C793 B.n753 VSUBS 0.013534f
C794 B.n754 VSUBS 0.013534f
C795 B.n755 VSUBS 0.013534f
C796 B.n756 VSUBS 0.013534f
C797 B.n757 VSUBS 0.013534f
C798 B.n758 VSUBS 0.013534f
C799 B.n759 VSUBS 0.013534f
C800 B.n760 VSUBS 0.013534f
C801 B.n761 VSUBS 0.013534f
C802 B.n762 VSUBS 0.013534f
C803 B.n763 VSUBS 0.013534f
C804 B.n764 VSUBS 0.013534f
C805 B.n765 VSUBS 0.013534f
C806 B.n766 VSUBS 0.013534f
C807 B.n767 VSUBS 0.013534f
C808 B.n768 VSUBS 0.013534f
C809 B.n769 VSUBS 0.013534f
C810 B.n770 VSUBS 0.013534f
C811 B.n771 VSUBS 0.013534f
C812 B.n772 VSUBS 0.013534f
C813 B.n773 VSUBS 0.013534f
C814 B.n774 VSUBS 0.013534f
C815 B.n775 VSUBS 0.013534f
C816 B.n776 VSUBS 0.013534f
C817 B.n777 VSUBS 0.013534f
C818 B.n778 VSUBS 0.013534f
C819 B.n779 VSUBS 0.013534f
C820 B.n780 VSUBS 0.013534f
C821 B.n781 VSUBS 0.013534f
C822 B.n782 VSUBS 0.013534f
C823 B.n783 VSUBS 0.013534f
C824 B.n784 VSUBS 0.013534f
C825 B.n785 VSUBS 0.013534f
C826 B.n786 VSUBS 0.013534f
C827 B.n787 VSUBS 0.013534f
C828 B.n788 VSUBS 0.013534f
C829 B.n789 VSUBS 0.013534f
C830 B.n790 VSUBS 0.013534f
C831 B.n791 VSUBS 0.017661f
C832 B.n792 VSUBS 0.018814f
C833 B.n793 VSUBS 0.037413f
C834 VDD2.n0 VSUBS 0.045341f
C835 VDD2.n1 VSUBS 0.305392f
C836 VDD2.n2 VSUBS 0.022088f
C837 VDD2.t1 VSUBS 0.119982f
C838 VDD2.n3 VSUBS 0.141667f
C839 VDD2.n4 VSUBS 0.030783f
C840 VDD2.n5 VSUBS 0.039155f
C841 VDD2.n6 VSUBS 0.12699f
C842 VDD2.n7 VSUBS 0.023387f
C843 VDD2.n8 VSUBS 0.022088f
C844 VDD2.n9 VSUBS 0.107364f
C845 VDD2.n10 VSUBS 0.125342f
C846 VDD2.t2 VSUBS 0.085102f
C847 VDD2.t9 VSUBS 0.085102f
C848 VDD2.n11 VSUBS 0.420119f
C849 VDD2.n12 VSUBS 1.56399f
C850 VDD2.t8 VSUBS 0.085102f
C851 VDD2.t3 VSUBS 0.085102f
C852 VDD2.n13 VSUBS 0.440756f
C853 VDD2.n14 VSUBS 4.91382f
C854 VDD2.n15 VSUBS 0.045341f
C855 VDD2.n16 VSUBS 0.305392f
C856 VDD2.n17 VSUBS 0.022088f
C857 VDD2.t4 VSUBS 0.119982f
C858 VDD2.n18 VSUBS 0.141667f
C859 VDD2.n19 VSUBS 0.030783f
C860 VDD2.n20 VSUBS 0.039155f
C861 VDD2.n21 VSUBS 0.12699f
C862 VDD2.n22 VSUBS 0.023387f
C863 VDD2.n23 VSUBS 0.022088f
C864 VDD2.n24 VSUBS 0.107364f
C865 VDD2.n25 VSUBS 0.092546f
C866 VDD2.n26 VSUBS 4.23114f
C867 VDD2.t0 VSUBS 0.085102f
C868 VDD2.t6 VSUBS 0.085102f
C869 VDD2.n27 VSUBS 0.420121f
C870 VDD2.n28 VSUBS 1.06998f
C871 VDD2.t7 VSUBS 0.085102f
C872 VDD2.t5 VSUBS 0.085102f
C873 VDD2.n29 VSUBS 0.440721f
C874 VN.t6 VSUBS 1.01509f
C875 VN.n0 VSUBS 0.60105f
C876 VN.n1 VSUBS 0.043398f
C877 VN.n2 VSUBS 0.066687f
C878 VN.n3 VSUBS 0.043398f
C879 VN.n4 VSUBS 0.062201f
C880 VN.n5 VSUBS 0.043398f
C881 VN.n6 VSUBS 0.064286f
C882 VN.n7 VSUBS 0.043398f
C883 VN.n8 VSUBS 0.060612f
C884 VN.n9 VSUBS 0.043398f
C885 VN.n10 VSUBS 0.061885f
C886 VN.n11 VSUBS 0.043398f
C887 VN.n12 VSUBS 0.059023f
C888 VN.t7 VSUBS 1.01509f
C889 VN.n13 VSUBS 0.576497f
C890 VN.t8 VSUBS 1.51583f
C891 VN.n14 VSUBS 0.607992f
C892 VN.n15 VSUBS 0.543376f
C893 VN.n16 VSUBS 0.043398f
C894 VN.n17 VSUBS 0.080477f
C895 VN.n18 VSUBS 0.080477f
C896 VN.n19 VSUBS 0.064286f
C897 VN.n20 VSUBS 0.043398f
C898 VN.n21 VSUBS 0.043398f
C899 VN.n22 VSUBS 0.043398f
C900 VN.n23 VSUBS 0.080477f
C901 VN.n24 VSUBS 0.080477f
C902 VN.t0 VSUBS 1.01509f
C903 VN.n25 VSUBS 0.427416f
C904 VN.n26 VSUBS 0.060612f
C905 VN.n27 VSUBS 0.043398f
C906 VN.n28 VSUBS 0.043398f
C907 VN.n29 VSUBS 0.043398f
C908 VN.n30 VSUBS 0.080477f
C909 VN.n31 VSUBS 0.080477f
C910 VN.n32 VSUBS 0.061885f
C911 VN.n33 VSUBS 0.043398f
C912 VN.n34 VSUBS 0.043398f
C913 VN.n35 VSUBS 0.043398f
C914 VN.n36 VSUBS 0.080477f
C915 VN.n37 VSUBS 0.080477f
C916 VN.t1 VSUBS 1.01509f
C917 VN.n38 VSUBS 0.427416f
C918 VN.n39 VSUBS 0.059023f
C919 VN.n40 VSUBS 0.043398f
C920 VN.n41 VSUBS 0.043398f
C921 VN.n42 VSUBS 0.043398f
C922 VN.n43 VSUBS 0.080477f
C923 VN.n44 VSUBS 0.080477f
C924 VN.n45 VSUBS 0.059483f
C925 VN.n46 VSUBS 0.043398f
C926 VN.n47 VSUBS 0.043398f
C927 VN.n48 VSUBS 0.043398f
C928 VN.n49 VSUBS 0.080477f
C929 VN.n50 VSUBS 0.080477f
C930 VN.n51 VSUBS 0.057434f
C931 VN.n52 VSUBS 0.070032f
C932 VN.n53 VSUBS 0.119049f
C933 VN.t5 VSUBS 1.01509f
C934 VN.n54 VSUBS 0.60105f
C935 VN.n55 VSUBS 0.043398f
C936 VN.n56 VSUBS 0.066687f
C937 VN.n57 VSUBS 0.043398f
C938 VN.n58 VSUBS 0.062201f
C939 VN.n59 VSUBS 0.043398f
C940 VN.t9 VSUBS 1.01509f
C941 VN.n60 VSUBS 0.427416f
C942 VN.n61 VSUBS 0.064286f
C943 VN.n62 VSUBS 0.043398f
C944 VN.n63 VSUBS 0.060612f
C945 VN.n64 VSUBS 0.043398f
C946 VN.t3 VSUBS 1.01509f
C947 VN.n65 VSUBS 0.427416f
C948 VN.n66 VSUBS 0.061885f
C949 VN.n67 VSUBS 0.043398f
C950 VN.n68 VSUBS 0.059023f
C951 VN.t4 VSUBS 1.51583f
C952 VN.t2 VSUBS 1.01509f
C953 VN.n69 VSUBS 0.576497f
C954 VN.n70 VSUBS 0.607992f
C955 VN.n71 VSUBS 0.543376f
C956 VN.n72 VSUBS 0.043398f
C957 VN.n73 VSUBS 0.080477f
C958 VN.n74 VSUBS 0.080477f
C959 VN.n75 VSUBS 0.064286f
C960 VN.n76 VSUBS 0.043398f
C961 VN.n77 VSUBS 0.043398f
C962 VN.n78 VSUBS 0.043398f
C963 VN.n79 VSUBS 0.080477f
C964 VN.n80 VSUBS 0.080477f
C965 VN.n81 VSUBS 0.060612f
C966 VN.n82 VSUBS 0.043398f
C967 VN.n83 VSUBS 0.043398f
C968 VN.n84 VSUBS 0.043398f
C969 VN.n85 VSUBS 0.080477f
C970 VN.n86 VSUBS 0.080477f
C971 VN.n87 VSUBS 0.061885f
C972 VN.n88 VSUBS 0.043398f
C973 VN.n89 VSUBS 0.043398f
C974 VN.n90 VSUBS 0.043398f
C975 VN.n91 VSUBS 0.080477f
C976 VN.n92 VSUBS 0.080477f
C977 VN.n93 VSUBS 0.059023f
C978 VN.n94 VSUBS 0.043398f
C979 VN.n95 VSUBS 0.043398f
C980 VN.n96 VSUBS 0.043398f
C981 VN.n97 VSUBS 0.080477f
C982 VN.n98 VSUBS 0.080477f
C983 VN.n99 VSUBS 0.059483f
C984 VN.n100 VSUBS 0.043398f
C985 VN.n101 VSUBS 0.043398f
C986 VN.n102 VSUBS 0.043398f
C987 VN.n103 VSUBS 0.080477f
C988 VN.n104 VSUBS 0.080477f
C989 VN.n105 VSUBS 0.057434f
C990 VN.n106 VSUBS 0.070032f
C991 VN.n107 VSUBS 2.63409f
C992 VTAIL.t3 VSUBS 0.082043f
C993 VTAIL.t0 VSUBS 0.082043f
C994 VTAIL.n0 VSUBS 0.348872f
C995 VTAIL.n1 VSUBS 1.09378f
C996 VTAIL.n2 VSUBS 0.043711f
C997 VTAIL.n3 VSUBS 0.294412f
C998 VTAIL.n4 VSUBS 0.021294f
C999 VTAIL.t13 VSUBS 0.115668f
C1000 VTAIL.n5 VSUBS 0.136574f
C1001 VTAIL.n6 VSUBS 0.029676f
C1002 VTAIL.n7 VSUBS 0.037748f
C1003 VTAIL.n8 VSUBS 0.122424f
C1004 VTAIL.n9 VSUBS 0.022546f
C1005 VTAIL.n10 VSUBS 0.021294f
C1006 VTAIL.n11 VSUBS 0.103504f
C1007 VTAIL.n12 VSUBS 0.061938f
C1008 VTAIL.n13 VSUBS 0.757714f
C1009 VTAIL.t14 VSUBS 0.082043f
C1010 VTAIL.t15 VSUBS 0.082043f
C1011 VTAIL.n14 VSUBS 0.348872f
C1012 VTAIL.n15 VSUBS 1.35493f
C1013 VTAIL.t7 VSUBS 0.082043f
C1014 VTAIL.t9 VSUBS 0.082043f
C1015 VTAIL.n16 VSUBS 0.348872f
C1016 VTAIL.n17 VSUBS 2.6197f
C1017 VTAIL.t1 VSUBS 0.082043f
C1018 VTAIL.t17 VSUBS 0.082043f
C1019 VTAIL.n18 VSUBS 0.348874f
C1020 VTAIL.n19 VSUBS 2.61969f
C1021 VTAIL.t16 VSUBS 0.082043f
C1022 VTAIL.t4 VSUBS 0.082043f
C1023 VTAIL.n20 VSUBS 0.348874f
C1024 VTAIL.n21 VSUBS 1.35493f
C1025 VTAIL.n22 VSUBS 0.043711f
C1026 VTAIL.n23 VSUBS 0.294412f
C1027 VTAIL.n24 VSUBS 0.021294f
C1028 VTAIL.t5 VSUBS 0.115668f
C1029 VTAIL.n25 VSUBS 0.136574f
C1030 VTAIL.n26 VSUBS 0.029676f
C1031 VTAIL.n27 VSUBS 0.037748f
C1032 VTAIL.n28 VSUBS 0.122424f
C1033 VTAIL.n29 VSUBS 0.022546f
C1034 VTAIL.n30 VSUBS 0.021294f
C1035 VTAIL.n31 VSUBS 0.103504f
C1036 VTAIL.n32 VSUBS 0.061938f
C1037 VTAIL.n33 VSUBS 0.757714f
C1038 VTAIL.t10 VSUBS 0.082043f
C1039 VTAIL.t11 VSUBS 0.082043f
C1040 VTAIL.n34 VSUBS 0.348874f
C1041 VTAIL.n35 VSUBS 1.19587f
C1042 VTAIL.t6 VSUBS 0.082043f
C1043 VTAIL.t8 VSUBS 0.082043f
C1044 VTAIL.n36 VSUBS 0.348874f
C1045 VTAIL.n37 VSUBS 1.35493f
C1046 VTAIL.n38 VSUBS 0.043711f
C1047 VTAIL.n39 VSUBS 0.294412f
C1048 VTAIL.n40 VSUBS 0.021294f
C1049 VTAIL.t12 VSUBS 0.115668f
C1050 VTAIL.n41 VSUBS 0.136574f
C1051 VTAIL.n42 VSUBS 0.029676f
C1052 VTAIL.n43 VSUBS 0.037748f
C1053 VTAIL.n44 VSUBS 0.122424f
C1054 VTAIL.n45 VSUBS 0.022546f
C1055 VTAIL.n46 VSUBS 0.021294f
C1056 VTAIL.n47 VSUBS 0.103504f
C1057 VTAIL.n48 VSUBS 0.061938f
C1058 VTAIL.n49 VSUBS 1.74344f
C1059 VTAIL.n50 VSUBS 0.043711f
C1060 VTAIL.n51 VSUBS 0.294412f
C1061 VTAIL.n52 VSUBS 0.021294f
C1062 VTAIL.t19 VSUBS 0.115668f
C1063 VTAIL.n53 VSUBS 0.136574f
C1064 VTAIL.n54 VSUBS 0.029676f
C1065 VTAIL.n55 VSUBS 0.037748f
C1066 VTAIL.n56 VSUBS 0.122424f
C1067 VTAIL.n57 VSUBS 0.022546f
C1068 VTAIL.n58 VSUBS 0.021294f
C1069 VTAIL.n59 VSUBS 0.103504f
C1070 VTAIL.n60 VSUBS 0.061938f
C1071 VTAIL.n61 VSUBS 1.74344f
C1072 VTAIL.t18 VSUBS 0.082043f
C1073 VTAIL.t2 VSUBS 0.082043f
C1074 VTAIL.n62 VSUBS 0.348872f
C1075 VTAIL.n63 VSUBS 1.01893f
C1076 VDD1.n0 VSUBS 0.045213f
C1077 VDD1.n1 VSUBS 0.304525f
C1078 VDD1.n2 VSUBS 0.022025f
C1079 VDD1.t9 VSUBS 0.119641f
C1080 VDD1.n3 VSUBS 0.141265f
C1081 VDD1.n4 VSUBS 0.030695f
C1082 VDD1.n5 VSUBS 0.039044f
C1083 VDD1.n6 VSUBS 0.126629f
C1084 VDD1.n7 VSUBS 0.023321f
C1085 VDD1.n8 VSUBS 0.022025f
C1086 VDD1.n9 VSUBS 0.107059f
C1087 VDD1.n10 VSUBS 0.124986f
C1088 VDD1.t6 VSUBS 0.084861f
C1089 VDD1.t1 VSUBS 0.084861f
C1090 VDD1.n11 VSUBS 0.418928f
C1091 VDD1.n12 VSUBS 1.57336f
C1092 VDD1.n13 VSUBS 0.045213f
C1093 VDD1.n14 VSUBS 0.304525f
C1094 VDD1.n15 VSUBS 0.022025f
C1095 VDD1.t5 VSUBS 0.119641f
C1096 VDD1.n16 VSUBS 0.141265f
C1097 VDD1.n17 VSUBS 0.030695f
C1098 VDD1.n18 VSUBS 0.039044f
C1099 VDD1.n19 VSUBS 0.126629f
C1100 VDD1.n20 VSUBS 0.023321f
C1101 VDD1.n21 VSUBS 0.022025f
C1102 VDD1.n22 VSUBS 0.107059f
C1103 VDD1.n23 VSUBS 0.124986f
C1104 VDD1.t8 VSUBS 0.084861f
C1105 VDD1.t4 VSUBS 0.084861f
C1106 VDD1.n24 VSUBS 0.418927f
C1107 VDD1.n25 VSUBS 1.55955f
C1108 VDD1.t2 VSUBS 0.084861f
C1109 VDD1.t0 VSUBS 0.084861f
C1110 VDD1.n26 VSUBS 0.439505f
C1111 VDD1.n27 VSUBS 5.1368f
C1112 VDD1.t3 VSUBS 0.084861f
C1113 VDD1.t7 VSUBS 0.084861f
C1114 VDD1.n28 VSUBS 0.418927f
C1115 VDD1.n29 VSUBS 4.88912f
C1116 VP.t2 VSUBS 1.16466f
C1117 VP.n0 VSUBS 0.689614f
C1118 VP.n1 VSUBS 0.049792f
C1119 VP.n2 VSUBS 0.076514f
C1120 VP.n3 VSUBS 0.049792f
C1121 VP.n4 VSUBS 0.071367f
C1122 VP.n5 VSUBS 0.049792f
C1123 VP.n6 VSUBS 0.073758f
C1124 VP.n7 VSUBS 0.049792f
C1125 VP.n8 VSUBS 0.069544f
C1126 VP.n9 VSUBS 0.049792f
C1127 VP.n10 VSUBS 0.071003f
C1128 VP.n11 VSUBS 0.049792f
C1129 VP.n12 VSUBS 0.06772f
C1130 VP.n13 VSUBS 0.049792f
C1131 VP.n14 VSUBS 0.068248f
C1132 VP.n15 VSUBS 0.049792f
C1133 VP.n16 VSUBS 0.065897f
C1134 VP.t3 VSUBS 1.16466f
C1135 VP.n17 VSUBS 0.689614f
C1136 VP.n18 VSUBS 0.049792f
C1137 VP.n19 VSUBS 0.076514f
C1138 VP.n20 VSUBS 0.049792f
C1139 VP.n21 VSUBS 0.071367f
C1140 VP.n22 VSUBS 0.049792f
C1141 VP.n23 VSUBS 0.073758f
C1142 VP.n24 VSUBS 0.049792f
C1143 VP.n25 VSUBS 0.069544f
C1144 VP.n26 VSUBS 0.049792f
C1145 VP.n27 VSUBS 0.071003f
C1146 VP.n28 VSUBS 0.049792f
C1147 VP.n29 VSUBS 0.06772f
C1148 VP.t5 VSUBS 1.73918f
C1149 VP.t4 VSUBS 1.16466f
C1150 VP.n30 VSUBS 0.661443f
C1151 VP.n31 VSUBS 0.69758f
C1152 VP.n32 VSUBS 0.623443f
C1153 VP.n33 VSUBS 0.049792f
C1154 VP.n34 VSUBS 0.092335f
C1155 VP.n35 VSUBS 0.092335f
C1156 VP.n36 VSUBS 0.073758f
C1157 VP.n37 VSUBS 0.049792f
C1158 VP.n38 VSUBS 0.049792f
C1159 VP.n39 VSUBS 0.049792f
C1160 VP.n40 VSUBS 0.092335f
C1161 VP.n41 VSUBS 0.092335f
C1162 VP.t9 VSUBS 1.16466f
C1163 VP.n42 VSUBS 0.490395f
C1164 VP.n43 VSUBS 0.069544f
C1165 VP.n44 VSUBS 0.049792f
C1166 VP.n45 VSUBS 0.049792f
C1167 VP.n46 VSUBS 0.049792f
C1168 VP.n47 VSUBS 0.092335f
C1169 VP.n48 VSUBS 0.092335f
C1170 VP.n49 VSUBS 0.071003f
C1171 VP.n50 VSUBS 0.049792f
C1172 VP.n51 VSUBS 0.049792f
C1173 VP.n52 VSUBS 0.049792f
C1174 VP.n53 VSUBS 0.092335f
C1175 VP.n54 VSUBS 0.092335f
C1176 VP.t7 VSUBS 1.16466f
C1177 VP.n55 VSUBS 0.490395f
C1178 VP.n56 VSUBS 0.06772f
C1179 VP.n57 VSUBS 0.049792f
C1180 VP.n58 VSUBS 0.049792f
C1181 VP.n59 VSUBS 0.049792f
C1182 VP.n60 VSUBS 0.092335f
C1183 VP.n61 VSUBS 0.092335f
C1184 VP.n62 VSUBS 0.068248f
C1185 VP.n63 VSUBS 0.049792f
C1186 VP.n64 VSUBS 0.049792f
C1187 VP.n65 VSUBS 0.049792f
C1188 VP.n66 VSUBS 0.092335f
C1189 VP.n67 VSUBS 0.092335f
C1190 VP.n68 VSUBS 0.065897f
C1191 VP.n69 VSUBS 0.080351f
C1192 VP.n70 VSUBS 3.00212f
C1193 VP.t8 VSUBS 1.16466f
C1194 VP.n71 VSUBS 0.689614f
C1195 VP.n72 VSUBS 3.03675f
C1196 VP.n73 VSUBS 0.080351f
C1197 VP.n74 VSUBS 0.049792f
C1198 VP.n75 VSUBS 0.092335f
C1199 VP.n76 VSUBS 0.092335f
C1200 VP.n77 VSUBS 0.076514f
C1201 VP.n78 VSUBS 0.049792f
C1202 VP.n79 VSUBS 0.049792f
C1203 VP.n80 VSUBS 0.049792f
C1204 VP.n81 VSUBS 0.092335f
C1205 VP.n82 VSUBS 0.092335f
C1206 VP.t6 VSUBS 1.16466f
C1207 VP.n83 VSUBS 0.490395f
C1208 VP.n84 VSUBS 0.071367f
C1209 VP.n85 VSUBS 0.049792f
C1210 VP.n86 VSUBS 0.049792f
C1211 VP.n87 VSUBS 0.049792f
C1212 VP.n88 VSUBS 0.092335f
C1213 VP.n89 VSUBS 0.092335f
C1214 VP.n90 VSUBS 0.073758f
C1215 VP.n91 VSUBS 0.049792f
C1216 VP.n92 VSUBS 0.049792f
C1217 VP.n93 VSUBS 0.049792f
C1218 VP.n94 VSUBS 0.092335f
C1219 VP.n95 VSUBS 0.092335f
C1220 VP.t1 VSUBS 1.16466f
C1221 VP.n96 VSUBS 0.490395f
C1222 VP.n97 VSUBS 0.069544f
C1223 VP.n98 VSUBS 0.049792f
C1224 VP.n99 VSUBS 0.049792f
C1225 VP.n100 VSUBS 0.049792f
C1226 VP.n101 VSUBS 0.092335f
C1227 VP.n102 VSUBS 0.092335f
C1228 VP.n103 VSUBS 0.071003f
C1229 VP.n104 VSUBS 0.049792f
C1230 VP.n105 VSUBS 0.049792f
C1231 VP.n106 VSUBS 0.049792f
C1232 VP.n107 VSUBS 0.092335f
C1233 VP.n108 VSUBS 0.092335f
C1234 VP.t0 VSUBS 1.16466f
C1235 VP.n109 VSUBS 0.490395f
C1236 VP.n110 VSUBS 0.06772f
C1237 VP.n111 VSUBS 0.049792f
C1238 VP.n112 VSUBS 0.049792f
C1239 VP.n113 VSUBS 0.049792f
C1240 VP.n114 VSUBS 0.092335f
C1241 VP.n115 VSUBS 0.092335f
C1242 VP.n116 VSUBS 0.068248f
C1243 VP.n117 VSUBS 0.049792f
C1244 VP.n118 VSUBS 0.049792f
C1245 VP.n119 VSUBS 0.049792f
C1246 VP.n120 VSUBS 0.092335f
C1247 VP.n121 VSUBS 0.092335f
C1248 VP.n122 VSUBS 0.065897f
C1249 VP.n123 VSUBS 0.080351f
C1250 VP.n124 VSUBS 0.136591f
.ends

