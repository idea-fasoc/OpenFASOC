* NGSPICE file created from diff_pair_sample_0644.ext - technology: sky130A

.subckt diff_pair_sample_0644 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=0 ps=0 w=14.83 l=0.57
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=2.44695 ps=15.16 w=14.83 l=0.57
X2 VDD2.t5 VN.t0 VTAIL.t11 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=2.44695 ps=15.16 w=14.83 l=0.57
X3 VDD2.t4 VN.t1 VTAIL.t0 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=2.44695 ps=15.16 w=14.83 l=0.57
X4 B.t8 B.t6 B.t7 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=0 ps=0 w=14.83 l=0.57
X5 VDD1.t4 VP.t1 VTAIL.t6 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=5.7837 ps=30.44 w=14.83 l=0.57
X6 VTAIL.t1 VN.t2 VDD2.t3 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=2.44695 ps=15.16 w=14.83 l=0.57
X7 VTAIL.t7 VP.t2 VDD1.t3 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=2.44695 ps=15.16 w=14.83 l=0.57
X8 VDD2.t2 VN.t3 VTAIL.t4 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=5.7837 ps=30.44 w=14.83 l=0.57
X9 VDD1.t2 VP.t3 VTAIL.t8 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=5.7837 ps=30.44 w=14.83 l=0.57
X10 VDD1.t1 VP.t4 VTAIL.t9 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=2.44695 ps=15.16 w=14.83 l=0.57
X11 VTAIL.t3 VN.t4 VDD2.t1 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=2.44695 ps=15.16 w=14.83 l=0.57
X12 B.t5 B.t3 B.t4 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=0 ps=0 w=14.83 l=0.57
X13 B.t2 B.t0 B.t1 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=5.7837 pd=30.44 as=0 ps=0 w=14.83 l=0.57
X14 VTAIL.t10 VP.t5 VDD1.t0 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=2.44695 ps=15.16 w=14.83 l=0.57
X15 VDD2.t0 VN.t5 VTAIL.t2 w_n1690_n3934# sky130_fd_pr__pfet_01v8 ad=2.44695 pd=15.16 as=5.7837 ps=30.44 w=14.83 l=0.57
R0 B.n122 B.t3 831.952
R1 B.n114 B.t9 831.952
R2 B.n44 B.t6 831.952
R3 B.n36 B.t0 831.952
R4 B.n346 B.n89 585
R5 B.n345 B.n344 585
R6 B.n343 B.n90 585
R7 B.n342 B.n341 585
R8 B.n340 B.n91 585
R9 B.n339 B.n338 585
R10 B.n337 B.n92 585
R11 B.n336 B.n335 585
R12 B.n334 B.n93 585
R13 B.n333 B.n332 585
R14 B.n331 B.n94 585
R15 B.n330 B.n329 585
R16 B.n328 B.n95 585
R17 B.n327 B.n326 585
R18 B.n325 B.n96 585
R19 B.n324 B.n323 585
R20 B.n322 B.n97 585
R21 B.n321 B.n320 585
R22 B.n319 B.n98 585
R23 B.n318 B.n317 585
R24 B.n316 B.n99 585
R25 B.n315 B.n314 585
R26 B.n313 B.n100 585
R27 B.n312 B.n311 585
R28 B.n310 B.n101 585
R29 B.n309 B.n308 585
R30 B.n307 B.n102 585
R31 B.n306 B.n305 585
R32 B.n304 B.n103 585
R33 B.n303 B.n302 585
R34 B.n301 B.n104 585
R35 B.n300 B.n299 585
R36 B.n298 B.n105 585
R37 B.n297 B.n296 585
R38 B.n295 B.n106 585
R39 B.n294 B.n293 585
R40 B.n292 B.n107 585
R41 B.n291 B.n290 585
R42 B.n289 B.n108 585
R43 B.n288 B.n287 585
R44 B.n286 B.n109 585
R45 B.n285 B.n284 585
R46 B.n283 B.n110 585
R47 B.n282 B.n281 585
R48 B.n280 B.n111 585
R49 B.n279 B.n278 585
R50 B.n277 B.n112 585
R51 B.n276 B.n275 585
R52 B.n274 B.n113 585
R53 B.n273 B.n272 585
R54 B.n271 B.n270 585
R55 B.n269 B.n117 585
R56 B.n268 B.n267 585
R57 B.n266 B.n118 585
R58 B.n265 B.n264 585
R59 B.n263 B.n119 585
R60 B.n262 B.n261 585
R61 B.n260 B.n120 585
R62 B.n259 B.n258 585
R63 B.n256 B.n121 585
R64 B.n255 B.n254 585
R65 B.n253 B.n124 585
R66 B.n252 B.n251 585
R67 B.n250 B.n125 585
R68 B.n249 B.n248 585
R69 B.n247 B.n126 585
R70 B.n246 B.n245 585
R71 B.n244 B.n127 585
R72 B.n243 B.n242 585
R73 B.n241 B.n128 585
R74 B.n240 B.n239 585
R75 B.n238 B.n129 585
R76 B.n237 B.n236 585
R77 B.n235 B.n130 585
R78 B.n234 B.n233 585
R79 B.n232 B.n131 585
R80 B.n231 B.n230 585
R81 B.n229 B.n132 585
R82 B.n228 B.n227 585
R83 B.n226 B.n133 585
R84 B.n225 B.n224 585
R85 B.n223 B.n134 585
R86 B.n222 B.n221 585
R87 B.n220 B.n135 585
R88 B.n219 B.n218 585
R89 B.n217 B.n136 585
R90 B.n216 B.n215 585
R91 B.n214 B.n137 585
R92 B.n213 B.n212 585
R93 B.n211 B.n138 585
R94 B.n210 B.n209 585
R95 B.n208 B.n139 585
R96 B.n207 B.n206 585
R97 B.n205 B.n140 585
R98 B.n204 B.n203 585
R99 B.n202 B.n141 585
R100 B.n201 B.n200 585
R101 B.n199 B.n142 585
R102 B.n198 B.n197 585
R103 B.n196 B.n143 585
R104 B.n195 B.n194 585
R105 B.n193 B.n144 585
R106 B.n192 B.n191 585
R107 B.n190 B.n145 585
R108 B.n189 B.n188 585
R109 B.n187 B.n146 585
R110 B.n186 B.n185 585
R111 B.n184 B.n147 585
R112 B.n183 B.n182 585
R113 B.n348 B.n347 585
R114 B.n349 B.n88 585
R115 B.n351 B.n350 585
R116 B.n352 B.n87 585
R117 B.n354 B.n353 585
R118 B.n355 B.n86 585
R119 B.n357 B.n356 585
R120 B.n358 B.n85 585
R121 B.n360 B.n359 585
R122 B.n361 B.n84 585
R123 B.n363 B.n362 585
R124 B.n364 B.n83 585
R125 B.n366 B.n365 585
R126 B.n367 B.n82 585
R127 B.n369 B.n368 585
R128 B.n370 B.n81 585
R129 B.n372 B.n371 585
R130 B.n373 B.n80 585
R131 B.n375 B.n374 585
R132 B.n376 B.n79 585
R133 B.n378 B.n377 585
R134 B.n379 B.n78 585
R135 B.n381 B.n380 585
R136 B.n382 B.n77 585
R137 B.n384 B.n383 585
R138 B.n385 B.n76 585
R139 B.n387 B.n386 585
R140 B.n388 B.n75 585
R141 B.n390 B.n389 585
R142 B.n391 B.n74 585
R143 B.n393 B.n392 585
R144 B.n394 B.n73 585
R145 B.n396 B.n395 585
R146 B.n397 B.n72 585
R147 B.n399 B.n398 585
R148 B.n400 B.n71 585
R149 B.n402 B.n401 585
R150 B.n403 B.n70 585
R151 B.n568 B.n11 585
R152 B.n567 B.n566 585
R153 B.n565 B.n12 585
R154 B.n564 B.n563 585
R155 B.n562 B.n13 585
R156 B.n561 B.n560 585
R157 B.n559 B.n14 585
R158 B.n558 B.n557 585
R159 B.n556 B.n15 585
R160 B.n555 B.n554 585
R161 B.n553 B.n16 585
R162 B.n552 B.n551 585
R163 B.n550 B.n17 585
R164 B.n549 B.n548 585
R165 B.n547 B.n18 585
R166 B.n546 B.n545 585
R167 B.n544 B.n19 585
R168 B.n543 B.n542 585
R169 B.n541 B.n20 585
R170 B.n540 B.n539 585
R171 B.n538 B.n21 585
R172 B.n537 B.n536 585
R173 B.n535 B.n22 585
R174 B.n534 B.n533 585
R175 B.n532 B.n23 585
R176 B.n531 B.n530 585
R177 B.n529 B.n24 585
R178 B.n528 B.n527 585
R179 B.n526 B.n25 585
R180 B.n525 B.n524 585
R181 B.n523 B.n26 585
R182 B.n522 B.n521 585
R183 B.n520 B.n27 585
R184 B.n519 B.n518 585
R185 B.n517 B.n28 585
R186 B.n516 B.n515 585
R187 B.n514 B.n29 585
R188 B.n513 B.n512 585
R189 B.n511 B.n30 585
R190 B.n510 B.n509 585
R191 B.n508 B.n31 585
R192 B.n507 B.n506 585
R193 B.n505 B.n32 585
R194 B.n504 B.n503 585
R195 B.n502 B.n33 585
R196 B.n501 B.n500 585
R197 B.n499 B.n34 585
R198 B.n498 B.n497 585
R199 B.n496 B.n35 585
R200 B.n495 B.n494 585
R201 B.n493 B.n492 585
R202 B.n491 B.n39 585
R203 B.n490 B.n489 585
R204 B.n488 B.n40 585
R205 B.n487 B.n486 585
R206 B.n485 B.n41 585
R207 B.n484 B.n483 585
R208 B.n482 B.n42 585
R209 B.n481 B.n480 585
R210 B.n478 B.n43 585
R211 B.n477 B.n476 585
R212 B.n475 B.n46 585
R213 B.n474 B.n473 585
R214 B.n472 B.n47 585
R215 B.n471 B.n470 585
R216 B.n469 B.n48 585
R217 B.n468 B.n467 585
R218 B.n466 B.n49 585
R219 B.n465 B.n464 585
R220 B.n463 B.n50 585
R221 B.n462 B.n461 585
R222 B.n460 B.n51 585
R223 B.n459 B.n458 585
R224 B.n457 B.n52 585
R225 B.n456 B.n455 585
R226 B.n454 B.n53 585
R227 B.n453 B.n452 585
R228 B.n451 B.n54 585
R229 B.n450 B.n449 585
R230 B.n448 B.n55 585
R231 B.n447 B.n446 585
R232 B.n445 B.n56 585
R233 B.n444 B.n443 585
R234 B.n442 B.n57 585
R235 B.n441 B.n440 585
R236 B.n439 B.n58 585
R237 B.n438 B.n437 585
R238 B.n436 B.n59 585
R239 B.n435 B.n434 585
R240 B.n433 B.n60 585
R241 B.n432 B.n431 585
R242 B.n430 B.n61 585
R243 B.n429 B.n428 585
R244 B.n427 B.n62 585
R245 B.n426 B.n425 585
R246 B.n424 B.n63 585
R247 B.n423 B.n422 585
R248 B.n421 B.n64 585
R249 B.n420 B.n419 585
R250 B.n418 B.n65 585
R251 B.n417 B.n416 585
R252 B.n415 B.n66 585
R253 B.n414 B.n413 585
R254 B.n412 B.n67 585
R255 B.n411 B.n410 585
R256 B.n409 B.n68 585
R257 B.n408 B.n407 585
R258 B.n406 B.n69 585
R259 B.n405 B.n404 585
R260 B.n570 B.n569 585
R261 B.n571 B.n10 585
R262 B.n573 B.n572 585
R263 B.n574 B.n9 585
R264 B.n576 B.n575 585
R265 B.n577 B.n8 585
R266 B.n579 B.n578 585
R267 B.n580 B.n7 585
R268 B.n582 B.n581 585
R269 B.n583 B.n6 585
R270 B.n585 B.n584 585
R271 B.n586 B.n5 585
R272 B.n588 B.n587 585
R273 B.n589 B.n4 585
R274 B.n591 B.n590 585
R275 B.n592 B.n3 585
R276 B.n594 B.n593 585
R277 B.n595 B.n0 585
R278 B.n2 B.n1 585
R279 B.n157 B.n156 585
R280 B.n159 B.n158 585
R281 B.n160 B.n155 585
R282 B.n162 B.n161 585
R283 B.n163 B.n154 585
R284 B.n165 B.n164 585
R285 B.n166 B.n153 585
R286 B.n168 B.n167 585
R287 B.n169 B.n152 585
R288 B.n171 B.n170 585
R289 B.n172 B.n151 585
R290 B.n174 B.n173 585
R291 B.n175 B.n150 585
R292 B.n177 B.n176 585
R293 B.n178 B.n149 585
R294 B.n180 B.n179 585
R295 B.n181 B.n148 585
R296 B.n182 B.n181 569.379
R297 B.n348 B.n89 569.379
R298 B.n404 B.n403 569.379
R299 B.n570 B.n11 569.379
R300 B.n114 B.t10 444.108
R301 B.n44 B.t8 444.108
R302 B.n122 B.t4 444.108
R303 B.n36 B.t2 444.108
R304 B.n115 B.t11 426.654
R305 B.n45 B.t7 426.654
R306 B.n123 B.t5 426.654
R307 B.n37 B.t1 426.654
R308 B.n597 B.n596 256.663
R309 B.n596 B.n595 235.042
R310 B.n596 B.n2 235.042
R311 B.n182 B.n147 163.367
R312 B.n186 B.n147 163.367
R313 B.n187 B.n186 163.367
R314 B.n188 B.n187 163.367
R315 B.n188 B.n145 163.367
R316 B.n192 B.n145 163.367
R317 B.n193 B.n192 163.367
R318 B.n194 B.n193 163.367
R319 B.n194 B.n143 163.367
R320 B.n198 B.n143 163.367
R321 B.n199 B.n198 163.367
R322 B.n200 B.n199 163.367
R323 B.n200 B.n141 163.367
R324 B.n204 B.n141 163.367
R325 B.n205 B.n204 163.367
R326 B.n206 B.n205 163.367
R327 B.n206 B.n139 163.367
R328 B.n210 B.n139 163.367
R329 B.n211 B.n210 163.367
R330 B.n212 B.n211 163.367
R331 B.n212 B.n137 163.367
R332 B.n216 B.n137 163.367
R333 B.n217 B.n216 163.367
R334 B.n218 B.n217 163.367
R335 B.n218 B.n135 163.367
R336 B.n222 B.n135 163.367
R337 B.n223 B.n222 163.367
R338 B.n224 B.n223 163.367
R339 B.n224 B.n133 163.367
R340 B.n228 B.n133 163.367
R341 B.n229 B.n228 163.367
R342 B.n230 B.n229 163.367
R343 B.n230 B.n131 163.367
R344 B.n234 B.n131 163.367
R345 B.n235 B.n234 163.367
R346 B.n236 B.n235 163.367
R347 B.n236 B.n129 163.367
R348 B.n240 B.n129 163.367
R349 B.n241 B.n240 163.367
R350 B.n242 B.n241 163.367
R351 B.n242 B.n127 163.367
R352 B.n246 B.n127 163.367
R353 B.n247 B.n246 163.367
R354 B.n248 B.n247 163.367
R355 B.n248 B.n125 163.367
R356 B.n252 B.n125 163.367
R357 B.n253 B.n252 163.367
R358 B.n254 B.n253 163.367
R359 B.n254 B.n121 163.367
R360 B.n259 B.n121 163.367
R361 B.n260 B.n259 163.367
R362 B.n261 B.n260 163.367
R363 B.n261 B.n119 163.367
R364 B.n265 B.n119 163.367
R365 B.n266 B.n265 163.367
R366 B.n267 B.n266 163.367
R367 B.n267 B.n117 163.367
R368 B.n271 B.n117 163.367
R369 B.n272 B.n271 163.367
R370 B.n272 B.n113 163.367
R371 B.n276 B.n113 163.367
R372 B.n277 B.n276 163.367
R373 B.n278 B.n277 163.367
R374 B.n278 B.n111 163.367
R375 B.n282 B.n111 163.367
R376 B.n283 B.n282 163.367
R377 B.n284 B.n283 163.367
R378 B.n284 B.n109 163.367
R379 B.n288 B.n109 163.367
R380 B.n289 B.n288 163.367
R381 B.n290 B.n289 163.367
R382 B.n290 B.n107 163.367
R383 B.n294 B.n107 163.367
R384 B.n295 B.n294 163.367
R385 B.n296 B.n295 163.367
R386 B.n296 B.n105 163.367
R387 B.n300 B.n105 163.367
R388 B.n301 B.n300 163.367
R389 B.n302 B.n301 163.367
R390 B.n302 B.n103 163.367
R391 B.n306 B.n103 163.367
R392 B.n307 B.n306 163.367
R393 B.n308 B.n307 163.367
R394 B.n308 B.n101 163.367
R395 B.n312 B.n101 163.367
R396 B.n313 B.n312 163.367
R397 B.n314 B.n313 163.367
R398 B.n314 B.n99 163.367
R399 B.n318 B.n99 163.367
R400 B.n319 B.n318 163.367
R401 B.n320 B.n319 163.367
R402 B.n320 B.n97 163.367
R403 B.n324 B.n97 163.367
R404 B.n325 B.n324 163.367
R405 B.n326 B.n325 163.367
R406 B.n326 B.n95 163.367
R407 B.n330 B.n95 163.367
R408 B.n331 B.n330 163.367
R409 B.n332 B.n331 163.367
R410 B.n332 B.n93 163.367
R411 B.n336 B.n93 163.367
R412 B.n337 B.n336 163.367
R413 B.n338 B.n337 163.367
R414 B.n338 B.n91 163.367
R415 B.n342 B.n91 163.367
R416 B.n343 B.n342 163.367
R417 B.n344 B.n343 163.367
R418 B.n344 B.n89 163.367
R419 B.n403 B.n402 163.367
R420 B.n402 B.n71 163.367
R421 B.n398 B.n71 163.367
R422 B.n398 B.n397 163.367
R423 B.n397 B.n396 163.367
R424 B.n396 B.n73 163.367
R425 B.n392 B.n73 163.367
R426 B.n392 B.n391 163.367
R427 B.n391 B.n390 163.367
R428 B.n390 B.n75 163.367
R429 B.n386 B.n75 163.367
R430 B.n386 B.n385 163.367
R431 B.n385 B.n384 163.367
R432 B.n384 B.n77 163.367
R433 B.n380 B.n77 163.367
R434 B.n380 B.n379 163.367
R435 B.n379 B.n378 163.367
R436 B.n378 B.n79 163.367
R437 B.n374 B.n79 163.367
R438 B.n374 B.n373 163.367
R439 B.n373 B.n372 163.367
R440 B.n372 B.n81 163.367
R441 B.n368 B.n81 163.367
R442 B.n368 B.n367 163.367
R443 B.n367 B.n366 163.367
R444 B.n366 B.n83 163.367
R445 B.n362 B.n83 163.367
R446 B.n362 B.n361 163.367
R447 B.n361 B.n360 163.367
R448 B.n360 B.n85 163.367
R449 B.n356 B.n85 163.367
R450 B.n356 B.n355 163.367
R451 B.n355 B.n354 163.367
R452 B.n354 B.n87 163.367
R453 B.n350 B.n87 163.367
R454 B.n350 B.n349 163.367
R455 B.n349 B.n348 163.367
R456 B.n566 B.n11 163.367
R457 B.n566 B.n565 163.367
R458 B.n565 B.n564 163.367
R459 B.n564 B.n13 163.367
R460 B.n560 B.n13 163.367
R461 B.n560 B.n559 163.367
R462 B.n559 B.n558 163.367
R463 B.n558 B.n15 163.367
R464 B.n554 B.n15 163.367
R465 B.n554 B.n553 163.367
R466 B.n553 B.n552 163.367
R467 B.n552 B.n17 163.367
R468 B.n548 B.n17 163.367
R469 B.n548 B.n547 163.367
R470 B.n547 B.n546 163.367
R471 B.n546 B.n19 163.367
R472 B.n542 B.n19 163.367
R473 B.n542 B.n541 163.367
R474 B.n541 B.n540 163.367
R475 B.n540 B.n21 163.367
R476 B.n536 B.n21 163.367
R477 B.n536 B.n535 163.367
R478 B.n535 B.n534 163.367
R479 B.n534 B.n23 163.367
R480 B.n530 B.n23 163.367
R481 B.n530 B.n529 163.367
R482 B.n529 B.n528 163.367
R483 B.n528 B.n25 163.367
R484 B.n524 B.n25 163.367
R485 B.n524 B.n523 163.367
R486 B.n523 B.n522 163.367
R487 B.n522 B.n27 163.367
R488 B.n518 B.n27 163.367
R489 B.n518 B.n517 163.367
R490 B.n517 B.n516 163.367
R491 B.n516 B.n29 163.367
R492 B.n512 B.n29 163.367
R493 B.n512 B.n511 163.367
R494 B.n511 B.n510 163.367
R495 B.n510 B.n31 163.367
R496 B.n506 B.n31 163.367
R497 B.n506 B.n505 163.367
R498 B.n505 B.n504 163.367
R499 B.n504 B.n33 163.367
R500 B.n500 B.n33 163.367
R501 B.n500 B.n499 163.367
R502 B.n499 B.n498 163.367
R503 B.n498 B.n35 163.367
R504 B.n494 B.n35 163.367
R505 B.n494 B.n493 163.367
R506 B.n493 B.n39 163.367
R507 B.n489 B.n39 163.367
R508 B.n489 B.n488 163.367
R509 B.n488 B.n487 163.367
R510 B.n487 B.n41 163.367
R511 B.n483 B.n41 163.367
R512 B.n483 B.n482 163.367
R513 B.n482 B.n481 163.367
R514 B.n481 B.n43 163.367
R515 B.n476 B.n43 163.367
R516 B.n476 B.n475 163.367
R517 B.n475 B.n474 163.367
R518 B.n474 B.n47 163.367
R519 B.n470 B.n47 163.367
R520 B.n470 B.n469 163.367
R521 B.n469 B.n468 163.367
R522 B.n468 B.n49 163.367
R523 B.n464 B.n49 163.367
R524 B.n464 B.n463 163.367
R525 B.n463 B.n462 163.367
R526 B.n462 B.n51 163.367
R527 B.n458 B.n51 163.367
R528 B.n458 B.n457 163.367
R529 B.n457 B.n456 163.367
R530 B.n456 B.n53 163.367
R531 B.n452 B.n53 163.367
R532 B.n452 B.n451 163.367
R533 B.n451 B.n450 163.367
R534 B.n450 B.n55 163.367
R535 B.n446 B.n55 163.367
R536 B.n446 B.n445 163.367
R537 B.n445 B.n444 163.367
R538 B.n444 B.n57 163.367
R539 B.n440 B.n57 163.367
R540 B.n440 B.n439 163.367
R541 B.n439 B.n438 163.367
R542 B.n438 B.n59 163.367
R543 B.n434 B.n59 163.367
R544 B.n434 B.n433 163.367
R545 B.n433 B.n432 163.367
R546 B.n432 B.n61 163.367
R547 B.n428 B.n61 163.367
R548 B.n428 B.n427 163.367
R549 B.n427 B.n426 163.367
R550 B.n426 B.n63 163.367
R551 B.n422 B.n63 163.367
R552 B.n422 B.n421 163.367
R553 B.n421 B.n420 163.367
R554 B.n420 B.n65 163.367
R555 B.n416 B.n65 163.367
R556 B.n416 B.n415 163.367
R557 B.n415 B.n414 163.367
R558 B.n414 B.n67 163.367
R559 B.n410 B.n67 163.367
R560 B.n410 B.n409 163.367
R561 B.n409 B.n408 163.367
R562 B.n408 B.n69 163.367
R563 B.n404 B.n69 163.367
R564 B.n571 B.n570 163.367
R565 B.n572 B.n571 163.367
R566 B.n572 B.n9 163.367
R567 B.n576 B.n9 163.367
R568 B.n577 B.n576 163.367
R569 B.n578 B.n577 163.367
R570 B.n578 B.n7 163.367
R571 B.n582 B.n7 163.367
R572 B.n583 B.n582 163.367
R573 B.n584 B.n583 163.367
R574 B.n584 B.n5 163.367
R575 B.n588 B.n5 163.367
R576 B.n589 B.n588 163.367
R577 B.n590 B.n589 163.367
R578 B.n590 B.n3 163.367
R579 B.n594 B.n3 163.367
R580 B.n595 B.n594 163.367
R581 B.n157 B.n2 163.367
R582 B.n158 B.n157 163.367
R583 B.n158 B.n155 163.367
R584 B.n162 B.n155 163.367
R585 B.n163 B.n162 163.367
R586 B.n164 B.n163 163.367
R587 B.n164 B.n153 163.367
R588 B.n168 B.n153 163.367
R589 B.n169 B.n168 163.367
R590 B.n170 B.n169 163.367
R591 B.n170 B.n151 163.367
R592 B.n174 B.n151 163.367
R593 B.n175 B.n174 163.367
R594 B.n176 B.n175 163.367
R595 B.n176 B.n149 163.367
R596 B.n180 B.n149 163.367
R597 B.n181 B.n180 163.367
R598 B.n257 B.n123 59.5399
R599 B.n116 B.n115 59.5399
R600 B.n479 B.n45 59.5399
R601 B.n38 B.n37 59.5399
R602 B.n569 B.n568 36.9956
R603 B.n405 B.n70 36.9956
R604 B.n347 B.n346 36.9956
R605 B.n183 B.n148 36.9956
R606 B B.n597 18.0485
R607 B.n123 B.n122 17.455
R608 B.n115 B.n114 17.455
R609 B.n45 B.n44 17.455
R610 B.n37 B.n36 17.455
R611 B.n569 B.n10 10.6151
R612 B.n573 B.n10 10.6151
R613 B.n574 B.n573 10.6151
R614 B.n575 B.n574 10.6151
R615 B.n575 B.n8 10.6151
R616 B.n579 B.n8 10.6151
R617 B.n580 B.n579 10.6151
R618 B.n581 B.n580 10.6151
R619 B.n581 B.n6 10.6151
R620 B.n585 B.n6 10.6151
R621 B.n586 B.n585 10.6151
R622 B.n587 B.n586 10.6151
R623 B.n587 B.n4 10.6151
R624 B.n591 B.n4 10.6151
R625 B.n592 B.n591 10.6151
R626 B.n593 B.n592 10.6151
R627 B.n593 B.n0 10.6151
R628 B.n568 B.n567 10.6151
R629 B.n567 B.n12 10.6151
R630 B.n563 B.n12 10.6151
R631 B.n563 B.n562 10.6151
R632 B.n562 B.n561 10.6151
R633 B.n561 B.n14 10.6151
R634 B.n557 B.n14 10.6151
R635 B.n557 B.n556 10.6151
R636 B.n556 B.n555 10.6151
R637 B.n555 B.n16 10.6151
R638 B.n551 B.n16 10.6151
R639 B.n551 B.n550 10.6151
R640 B.n550 B.n549 10.6151
R641 B.n549 B.n18 10.6151
R642 B.n545 B.n18 10.6151
R643 B.n545 B.n544 10.6151
R644 B.n544 B.n543 10.6151
R645 B.n543 B.n20 10.6151
R646 B.n539 B.n20 10.6151
R647 B.n539 B.n538 10.6151
R648 B.n538 B.n537 10.6151
R649 B.n537 B.n22 10.6151
R650 B.n533 B.n22 10.6151
R651 B.n533 B.n532 10.6151
R652 B.n532 B.n531 10.6151
R653 B.n531 B.n24 10.6151
R654 B.n527 B.n24 10.6151
R655 B.n527 B.n526 10.6151
R656 B.n526 B.n525 10.6151
R657 B.n525 B.n26 10.6151
R658 B.n521 B.n26 10.6151
R659 B.n521 B.n520 10.6151
R660 B.n520 B.n519 10.6151
R661 B.n519 B.n28 10.6151
R662 B.n515 B.n28 10.6151
R663 B.n515 B.n514 10.6151
R664 B.n514 B.n513 10.6151
R665 B.n513 B.n30 10.6151
R666 B.n509 B.n30 10.6151
R667 B.n509 B.n508 10.6151
R668 B.n508 B.n507 10.6151
R669 B.n507 B.n32 10.6151
R670 B.n503 B.n32 10.6151
R671 B.n503 B.n502 10.6151
R672 B.n502 B.n501 10.6151
R673 B.n501 B.n34 10.6151
R674 B.n497 B.n34 10.6151
R675 B.n497 B.n496 10.6151
R676 B.n496 B.n495 10.6151
R677 B.n492 B.n491 10.6151
R678 B.n491 B.n490 10.6151
R679 B.n490 B.n40 10.6151
R680 B.n486 B.n40 10.6151
R681 B.n486 B.n485 10.6151
R682 B.n485 B.n484 10.6151
R683 B.n484 B.n42 10.6151
R684 B.n480 B.n42 10.6151
R685 B.n478 B.n477 10.6151
R686 B.n477 B.n46 10.6151
R687 B.n473 B.n46 10.6151
R688 B.n473 B.n472 10.6151
R689 B.n472 B.n471 10.6151
R690 B.n471 B.n48 10.6151
R691 B.n467 B.n48 10.6151
R692 B.n467 B.n466 10.6151
R693 B.n466 B.n465 10.6151
R694 B.n465 B.n50 10.6151
R695 B.n461 B.n50 10.6151
R696 B.n461 B.n460 10.6151
R697 B.n460 B.n459 10.6151
R698 B.n459 B.n52 10.6151
R699 B.n455 B.n52 10.6151
R700 B.n455 B.n454 10.6151
R701 B.n454 B.n453 10.6151
R702 B.n453 B.n54 10.6151
R703 B.n449 B.n54 10.6151
R704 B.n449 B.n448 10.6151
R705 B.n448 B.n447 10.6151
R706 B.n447 B.n56 10.6151
R707 B.n443 B.n56 10.6151
R708 B.n443 B.n442 10.6151
R709 B.n442 B.n441 10.6151
R710 B.n441 B.n58 10.6151
R711 B.n437 B.n58 10.6151
R712 B.n437 B.n436 10.6151
R713 B.n436 B.n435 10.6151
R714 B.n435 B.n60 10.6151
R715 B.n431 B.n60 10.6151
R716 B.n431 B.n430 10.6151
R717 B.n430 B.n429 10.6151
R718 B.n429 B.n62 10.6151
R719 B.n425 B.n62 10.6151
R720 B.n425 B.n424 10.6151
R721 B.n424 B.n423 10.6151
R722 B.n423 B.n64 10.6151
R723 B.n419 B.n64 10.6151
R724 B.n419 B.n418 10.6151
R725 B.n418 B.n417 10.6151
R726 B.n417 B.n66 10.6151
R727 B.n413 B.n66 10.6151
R728 B.n413 B.n412 10.6151
R729 B.n412 B.n411 10.6151
R730 B.n411 B.n68 10.6151
R731 B.n407 B.n68 10.6151
R732 B.n407 B.n406 10.6151
R733 B.n406 B.n405 10.6151
R734 B.n401 B.n70 10.6151
R735 B.n401 B.n400 10.6151
R736 B.n400 B.n399 10.6151
R737 B.n399 B.n72 10.6151
R738 B.n395 B.n72 10.6151
R739 B.n395 B.n394 10.6151
R740 B.n394 B.n393 10.6151
R741 B.n393 B.n74 10.6151
R742 B.n389 B.n74 10.6151
R743 B.n389 B.n388 10.6151
R744 B.n388 B.n387 10.6151
R745 B.n387 B.n76 10.6151
R746 B.n383 B.n76 10.6151
R747 B.n383 B.n382 10.6151
R748 B.n382 B.n381 10.6151
R749 B.n381 B.n78 10.6151
R750 B.n377 B.n78 10.6151
R751 B.n377 B.n376 10.6151
R752 B.n376 B.n375 10.6151
R753 B.n375 B.n80 10.6151
R754 B.n371 B.n80 10.6151
R755 B.n371 B.n370 10.6151
R756 B.n370 B.n369 10.6151
R757 B.n369 B.n82 10.6151
R758 B.n365 B.n82 10.6151
R759 B.n365 B.n364 10.6151
R760 B.n364 B.n363 10.6151
R761 B.n363 B.n84 10.6151
R762 B.n359 B.n84 10.6151
R763 B.n359 B.n358 10.6151
R764 B.n358 B.n357 10.6151
R765 B.n357 B.n86 10.6151
R766 B.n353 B.n86 10.6151
R767 B.n353 B.n352 10.6151
R768 B.n352 B.n351 10.6151
R769 B.n351 B.n88 10.6151
R770 B.n347 B.n88 10.6151
R771 B.n156 B.n1 10.6151
R772 B.n159 B.n156 10.6151
R773 B.n160 B.n159 10.6151
R774 B.n161 B.n160 10.6151
R775 B.n161 B.n154 10.6151
R776 B.n165 B.n154 10.6151
R777 B.n166 B.n165 10.6151
R778 B.n167 B.n166 10.6151
R779 B.n167 B.n152 10.6151
R780 B.n171 B.n152 10.6151
R781 B.n172 B.n171 10.6151
R782 B.n173 B.n172 10.6151
R783 B.n173 B.n150 10.6151
R784 B.n177 B.n150 10.6151
R785 B.n178 B.n177 10.6151
R786 B.n179 B.n178 10.6151
R787 B.n179 B.n148 10.6151
R788 B.n184 B.n183 10.6151
R789 B.n185 B.n184 10.6151
R790 B.n185 B.n146 10.6151
R791 B.n189 B.n146 10.6151
R792 B.n190 B.n189 10.6151
R793 B.n191 B.n190 10.6151
R794 B.n191 B.n144 10.6151
R795 B.n195 B.n144 10.6151
R796 B.n196 B.n195 10.6151
R797 B.n197 B.n196 10.6151
R798 B.n197 B.n142 10.6151
R799 B.n201 B.n142 10.6151
R800 B.n202 B.n201 10.6151
R801 B.n203 B.n202 10.6151
R802 B.n203 B.n140 10.6151
R803 B.n207 B.n140 10.6151
R804 B.n208 B.n207 10.6151
R805 B.n209 B.n208 10.6151
R806 B.n209 B.n138 10.6151
R807 B.n213 B.n138 10.6151
R808 B.n214 B.n213 10.6151
R809 B.n215 B.n214 10.6151
R810 B.n215 B.n136 10.6151
R811 B.n219 B.n136 10.6151
R812 B.n220 B.n219 10.6151
R813 B.n221 B.n220 10.6151
R814 B.n221 B.n134 10.6151
R815 B.n225 B.n134 10.6151
R816 B.n226 B.n225 10.6151
R817 B.n227 B.n226 10.6151
R818 B.n227 B.n132 10.6151
R819 B.n231 B.n132 10.6151
R820 B.n232 B.n231 10.6151
R821 B.n233 B.n232 10.6151
R822 B.n233 B.n130 10.6151
R823 B.n237 B.n130 10.6151
R824 B.n238 B.n237 10.6151
R825 B.n239 B.n238 10.6151
R826 B.n239 B.n128 10.6151
R827 B.n243 B.n128 10.6151
R828 B.n244 B.n243 10.6151
R829 B.n245 B.n244 10.6151
R830 B.n245 B.n126 10.6151
R831 B.n249 B.n126 10.6151
R832 B.n250 B.n249 10.6151
R833 B.n251 B.n250 10.6151
R834 B.n251 B.n124 10.6151
R835 B.n255 B.n124 10.6151
R836 B.n256 B.n255 10.6151
R837 B.n258 B.n120 10.6151
R838 B.n262 B.n120 10.6151
R839 B.n263 B.n262 10.6151
R840 B.n264 B.n263 10.6151
R841 B.n264 B.n118 10.6151
R842 B.n268 B.n118 10.6151
R843 B.n269 B.n268 10.6151
R844 B.n270 B.n269 10.6151
R845 B.n274 B.n273 10.6151
R846 B.n275 B.n274 10.6151
R847 B.n275 B.n112 10.6151
R848 B.n279 B.n112 10.6151
R849 B.n280 B.n279 10.6151
R850 B.n281 B.n280 10.6151
R851 B.n281 B.n110 10.6151
R852 B.n285 B.n110 10.6151
R853 B.n286 B.n285 10.6151
R854 B.n287 B.n286 10.6151
R855 B.n287 B.n108 10.6151
R856 B.n291 B.n108 10.6151
R857 B.n292 B.n291 10.6151
R858 B.n293 B.n292 10.6151
R859 B.n293 B.n106 10.6151
R860 B.n297 B.n106 10.6151
R861 B.n298 B.n297 10.6151
R862 B.n299 B.n298 10.6151
R863 B.n299 B.n104 10.6151
R864 B.n303 B.n104 10.6151
R865 B.n304 B.n303 10.6151
R866 B.n305 B.n304 10.6151
R867 B.n305 B.n102 10.6151
R868 B.n309 B.n102 10.6151
R869 B.n310 B.n309 10.6151
R870 B.n311 B.n310 10.6151
R871 B.n311 B.n100 10.6151
R872 B.n315 B.n100 10.6151
R873 B.n316 B.n315 10.6151
R874 B.n317 B.n316 10.6151
R875 B.n317 B.n98 10.6151
R876 B.n321 B.n98 10.6151
R877 B.n322 B.n321 10.6151
R878 B.n323 B.n322 10.6151
R879 B.n323 B.n96 10.6151
R880 B.n327 B.n96 10.6151
R881 B.n328 B.n327 10.6151
R882 B.n329 B.n328 10.6151
R883 B.n329 B.n94 10.6151
R884 B.n333 B.n94 10.6151
R885 B.n334 B.n333 10.6151
R886 B.n335 B.n334 10.6151
R887 B.n335 B.n92 10.6151
R888 B.n339 B.n92 10.6151
R889 B.n340 B.n339 10.6151
R890 B.n341 B.n340 10.6151
R891 B.n341 B.n90 10.6151
R892 B.n345 B.n90 10.6151
R893 B.n346 B.n345 10.6151
R894 B.n597 B.n0 8.11757
R895 B.n597 B.n1 8.11757
R896 B.n492 B.n38 6.5566
R897 B.n480 B.n479 6.5566
R898 B.n258 B.n257 6.5566
R899 B.n270 B.n116 6.5566
R900 B.n495 B.n38 4.05904
R901 B.n479 B.n478 4.05904
R902 B.n257 B.n256 4.05904
R903 B.n273 B.n116 4.05904
R904 VP.n1 VP.t4 723.184
R905 VP.n6 VP.t0 696.364
R906 VP.n7 VP.t5 696.364
R907 VP.n8 VP.t3 696.364
R908 VP.n3 VP.t1 696.364
R909 VP.n2 VP.t2 696.364
R910 VP.n9 VP.n8 161.3
R911 VP.n4 VP.n3 161.3
R912 VP.n6 VP.n5 161.3
R913 VP.n7 VP.n0 80.6037
R914 VP.n7 VP.n6 48.2005
R915 VP.n8 VP.n7 48.2005
R916 VP.n3 VP.n2 48.2005
R917 VP.n4 VP.n1 45.1367
R918 VP.n5 VP.n4 42.8944
R919 VP.n2 VP.n1 13.3799
R920 VP.n5 VP.n0 0.285035
R921 VP.n9 VP.n0 0.285035
R922 VP VP.n9 0.0516364
R923 VTAIL.n330 VTAIL.n254 756.745
R924 VTAIL.n78 VTAIL.n2 756.745
R925 VTAIL.n248 VTAIL.n172 756.745
R926 VTAIL.n164 VTAIL.n88 756.745
R927 VTAIL.n281 VTAIL.n280 585
R928 VTAIL.n278 VTAIL.n277 585
R929 VTAIL.n287 VTAIL.n286 585
R930 VTAIL.n289 VTAIL.n288 585
R931 VTAIL.n274 VTAIL.n273 585
R932 VTAIL.n295 VTAIL.n294 585
R933 VTAIL.n297 VTAIL.n296 585
R934 VTAIL.n270 VTAIL.n269 585
R935 VTAIL.n303 VTAIL.n302 585
R936 VTAIL.n305 VTAIL.n304 585
R937 VTAIL.n266 VTAIL.n265 585
R938 VTAIL.n311 VTAIL.n310 585
R939 VTAIL.n313 VTAIL.n312 585
R940 VTAIL.n262 VTAIL.n261 585
R941 VTAIL.n319 VTAIL.n318 585
R942 VTAIL.n322 VTAIL.n321 585
R943 VTAIL.n320 VTAIL.n258 585
R944 VTAIL.n327 VTAIL.n257 585
R945 VTAIL.n329 VTAIL.n328 585
R946 VTAIL.n331 VTAIL.n330 585
R947 VTAIL.n29 VTAIL.n28 585
R948 VTAIL.n26 VTAIL.n25 585
R949 VTAIL.n35 VTAIL.n34 585
R950 VTAIL.n37 VTAIL.n36 585
R951 VTAIL.n22 VTAIL.n21 585
R952 VTAIL.n43 VTAIL.n42 585
R953 VTAIL.n45 VTAIL.n44 585
R954 VTAIL.n18 VTAIL.n17 585
R955 VTAIL.n51 VTAIL.n50 585
R956 VTAIL.n53 VTAIL.n52 585
R957 VTAIL.n14 VTAIL.n13 585
R958 VTAIL.n59 VTAIL.n58 585
R959 VTAIL.n61 VTAIL.n60 585
R960 VTAIL.n10 VTAIL.n9 585
R961 VTAIL.n67 VTAIL.n66 585
R962 VTAIL.n70 VTAIL.n69 585
R963 VTAIL.n68 VTAIL.n6 585
R964 VTAIL.n75 VTAIL.n5 585
R965 VTAIL.n77 VTAIL.n76 585
R966 VTAIL.n79 VTAIL.n78 585
R967 VTAIL.n249 VTAIL.n248 585
R968 VTAIL.n247 VTAIL.n246 585
R969 VTAIL.n245 VTAIL.n175 585
R970 VTAIL.n179 VTAIL.n176 585
R971 VTAIL.n240 VTAIL.n239 585
R972 VTAIL.n238 VTAIL.n237 585
R973 VTAIL.n181 VTAIL.n180 585
R974 VTAIL.n232 VTAIL.n231 585
R975 VTAIL.n230 VTAIL.n229 585
R976 VTAIL.n185 VTAIL.n184 585
R977 VTAIL.n224 VTAIL.n223 585
R978 VTAIL.n222 VTAIL.n221 585
R979 VTAIL.n189 VTAIL.n188 585
R980 VTAIL.n216 VTAIL.n215 585
R981 VTAIL.n214 VTAIL.n213 585
R982 VTAIL.n193 VTAIL.n192 585
R983 VTAIL.n208 VTAIL.n207 585
R984 VTAIL.n206 VTAIL.n205 585
R985 VTAIL.n197 VTAIL.n196 585
R986 VTAIL.n200 VTAIL.n199 585
R987 VTAIL.n165 VTAIL.n164 585
R988 VTAIL.n163 VTAIL.n162 585
R989 VTAIL.n161 VTAIL.n91 585
R990 VTAIL.n95 VTAIL.n92 585
R991 VTAIL.n156 VTAIL.n155 585
R992 VTAIL.n154 VTAIL.n153 585
R993 VTAIL.n97 VTAIL.n96 585
R994 VTAIL.n148 VTAIL.n147 585
R995 VTAIL.n146 VTAIL.n145 585
R996 VTAIL.n101 VTAIL.n100 585
R997 VTAIL.n140 VTAIL.n139 585
R998 VTAIL.n138 VTAIL.n137 585
R999 VTAIL.n105 VTAIL.n104 585
R1000 VTAIL.n132 VTAIL.n131 585
R1001 VTAIL.n130 VTAIL.n129 585
R1002 VTAIL.n109 VTAIL.n108 585
R1003 VTAIL.n124 VTAIL.n123 585
R1004 VTAIL.n122 VTAIL.n121 585
R1005 VTAIL.n113 VTAIL.n112 585
R1006 VTAIL.n116 VTAIL.n115 585
R1007 VTAIL.t6 VTAIL.n198 327.466
R1008 VTAIL.t4 VTAIL.n114 327.466
R1009 VTAIL.t2 VTAIL.n279 327.466
R1010 VTAIL.t8 VTAIL.n27 327.466
R1011 VTAIL.n280 VTAIL.n277 171.744
R1012 VTAIL.n287 VTAIL.n277 171.744
R1013 VTAIL.n288 VTAIL.n287 171.744
R1014 VTAIL.n288 VTAIL.n273 171.744
R1015 VTAIL.n295 VTAIL.n273 171.744
R1016 VTAIL.n296 VTAIL.n295 171.744
R1017 VTAIL.n296 VTAIL.n269 171.744
R1018 VTAIL.n303 VTAIL.n269 171.744
R1019 VTAIL.n304 VTAIL.n303 171.744
R1020 VTAIL.n304 VTAIL.n265 171.744
R1021 VTAIL.n311 VTAIL.n265 171.744
R1022 VTAIL.n312 VTAIL.n311 171.744
R1023 VTAIL.n312 VTAIL.n261 171.744
R1024 VTAIL.n319 VTAIL.n261 171.744
R1025 VTAIL.n321 VTAIL.n319 171.744
R1026 VTAIL.n321 VTAIL.n320 171.744
R1027 VTAIL.n320 VTAIL.n257 171.744
R1028 VTAIL.n329 VTAIL.n257 171.744
R1029 VTAIL.n330 VTAIL.n329 171.744
R1030 VTAIL.n28 VTAIL.n25 171.744
R1031 VTAIL.n35 VTAIL.n25 171.744
R1032 VTAIL.n36 VTAIL.n35 171.744
R1033 VTAIL.n36 VTAIL.n21 171.744
R1034 VTAIL.n43 VTAIL.n21 171.744
R1035 VTAIL.n44 VTAIL.n43 171.744
R1036 VTAIL.n44 VTAIL.n17 171.744
R1037 VTAIL.n51 VTAIL.n17 171.744
R1038 VTAIL.n52 VTAIL.n51 171.744
R1039 VTAIL.n52 VTAIL.n13 171.744
R1040 VTAIL.n59 VTAIL.n13 171.744
R1041 VTAIL.n60 VTAIL.n59 171.744
R1042 VTAIL.n60 VTAIL.n9 171.744
R1043 VTAIL.n67 VTAIL.n9 171.744
R1044 VTAIL.n69 VTAIL.n67 171.744
R1045 VTAIL.n69 VTAIL.n68 171.744
R1046 VTAIL.n68 VTAIL.n5 171.744
R1047 VTAIL.n77 VTAIL.n5 171.744
R1048 VTAIL.n78 VTAIL.n77 171.744
R1049 VTAIL.n248 VTAIL.n247 171.744
R1050 VTAIL.n247 VTAIL.n175 171.744
R1051 VTAIL.n179 VTAIL.n175 171.744
R1052 VTAIL.n239 VTAIL.n179 171.744
R1053 VTAIL.n239 VTAIL.n238 171.744
R1054 VTAIL.n238 VTAIL.n180 171.744
R1055 VTAIL.n231 VTAIL.n180 171.744
R1056 VTAIL.n231 VTAIL.n230 171.744
R1057 VTAIL.n230 VTAIL.n184 171.744
R1058 VTAIL.n223 VTAIL.n184 171.744
R1059 VTAIL.n223 VTAIL.n222 171.744
R1060 VTAIL.n222 VTAIL.n188 171.744
R1061 VTAIL.n215 VTAIL.n188 171.744
R1062 VTAIL.n215 VTAIL.n214 171.744
R1063 VTAIL.n214 VTAIL.n192 171.744
R1064 VTAIL.n207 VTAIL.n192 171.744
R1065 VTAIL.n207 VTAIL.n206 171.744
R1066 VTAIL.n206 VTAIL.n196 171.744
R1067 VTAIL.n199 VTAIL.n196 171.744
R1068 VTAIL.n164 VTAIL.n163 171.744
R1069 VTAIL.n163 VTAIL.n91 171.744
R1070 VTAIL.n95 VTAIL.n91 171.744
R1071 VTAIL.n155 VTAIL.n95 171.744
R1072 VTAIL.n155 VTAIL.n154 171.744
R1073 VTAIL.n154 VTAIL.n96 171.744
R1074 VTAIL.n147 VTAIL.n96 171.744
R1075 VTAIL.n147 VTAIL.n146 171.744
R1076 VTAIL.n146 VTAIL.n100 171.744
R1077 VTAIL.n139 VTAIL.n100 171.744
R1078 VTAIL.n139 VTAIL.n138 171.744
R1079 VTAIL.n138 VTAIL.n104 171.744
R1080 VTAIL.n131 VTAIL.n104 171.744
R1081 VTAIL.n131 VTAIL.n130 171.744
R1082 VTAIL.n130 VTAIL.n108 171.744
R1083 VTAIL.n123 VTAIL.n108 171.744
R1084 VTAIL.n123 VTAIL.n122 171.744
R1085 VTAIL.n122 VTAIL.n112 171.744
R1086 VTAIL.n115 VTAIL.n112 171.744
R1087 VTAIL.n280 VTAIL.t2 85.8723
R1088 VTAIL.n28 VTAIL.t8 85.8723
R1089 VTAIL.n199 VTAIL.t6 85.8723
R1090 VTAIL.n115 VTAIL.t4 85.8723
R1091 VTAIL.n171 VTAIL.n170 57.7726
R1092 VTAIL.n87 VTAIL.n86 57.7726
R1093 VTAIL.n1 VTAIL.n0 57.7724
R1094 VTAIL.n85 VTAIL.n84 57.7724
R1095 VTAIL.n335 VTAIL.n334 35.8702
R1096 VTAIL.n83 VTAIL.n82 35.8702
R1097 VTAIL.n253 VTAIL.n252 35.8702
R1098 VTAIL.n169 VTAIL.n168 35.8702
R1099 VTAIL.n87 VTAIL.n85 26.7031
R1100 VTAIL.n335 VTAIL.n253 25.9272
R1101 VTAIL.n281 VTAIL.n279 16.3895
R1102 VTAIL.n29 VTAIL.n27 16.3895
R1103 VTAIL.n200 VTAIL.n198 16.3895
R1104 VTAIL.n116 VTAIL.n114 16.3895
R1105 VTAIL.n328 VTAIL.n327 13.1884
R1106 VTAIL.n76 VTAIL.n75 13.1884
R1107 VTAIL.n246 VTAIL.n245 13.1884
R1108 VTAIL.n162 VTAIL.n161 13.1884
R1109 VTAIL.n282 VTAIL.n278 12.8005
R1110 VTAIL.n326 VTAIL.n258 12.8005
R1111 VTAIL.n331 VTAIL.n256 12.8005
R1112 VTAIL.n30 VTAIL.n26 12.8005
R1113 VTAIL.n74 VTAIL.n6 12.8005
R1114 VTAIL.n79 VTAIL.n4 12.8005
R1115 VTAIL.n249 VTAIL.n174 12.8005
R1116 VTAIL.n244 VTAIL.n176 12.8005
R1117 VTAIL.n201 VTAIL.n197 12.8005
R1118 VTAIL.n165 VTAIL.n90 12.8005
R1119 VTAIL.n160 VTAIL.n92 12.8005
R1120 VTAIL.n117 VTAIL.n113 12.8005
R1121 VTAIL.n286 VTAIL.n285 12.0247
R1122 VTAIL.n323 VTAIL.n322 12.0247
R1123 VTAIL.n332 VTAIL.n254 12.0247
R1124 VTAIL.n34 VTAIL.n33 12.0247
R1125 VTAIL.n71 VTAIL.n70 12.0247
R1126 VTAIL.n80 VTAIL.n2 12.0247
R1127 VTAIL.n250 VTAIL.n172 12.0247
R1128 VTAIL.n241 VTAIL.n240 12.0247
R1129 VTAIL.n205 VTAIL.n204 12.0247
R1130 VTAIL.n166 VTAIL.n88 12.0247
R1131 VTAIL.n157 VTAIL.n156 12.0247
R1132 VTAIL.n121 VTAIL.n120 12.0247
R1133 VTAIL.n289 VTAIL.n276 11.249
R1134 VTAIL.n318 VTAIL.n260 11.249
R1135 VTAIL.n37 VTAIL.n24 11.249
R1136 VTAIL.n66 VTAIL.n8 11.249
R1137 VTAIL.n237 VTAIL.n178 11.249
R1138 VTAIL.n208 VTAIL.n195 11.249
R1139 VTAIL.n153 VTAIL.n94 11.249
R1140 VTAIL.n124 VTAIL.n111 11.249
R1141 VTAIL.n290 VTAIL.n274 10.4732
R1142 VTAIL.n317 VTAIL.n262 10.4732
R1143 VTAIL.n38 VTAIL.n22 10.4732
R1144 VTAIL.n65 VTAIL.n10 10.4732
R1145 VTAIL.n236 VTAIL.n181 10.4732
R1146 VTAIL.n209 VTAIL.n193 10.4732
R1147 VTAIL.n152 VTAIL.n97 10.4732
R1148 VTAIL.n125 VTAIL.n109 10.4732
R1149 VTAIL.n294 VTAIL.n293 9.69747
R1150 VTAIL.n314 VTAIL.n313 9.69747
R1151 VTAIL.n42 VTAIL.n41 9.69747
R1152 VTAIL.n62 VTAIL.n61 9.69747
R1153 VTAIL.n233 VTAIL.n232 9.69747
R1154 VTAIL.n213 VTAIL.n212 9.69747
R1155 VTAIL.n149 VTAIL.n148 9.69747
R1156 VTAIL.n129 VTAIL.n128 9.69747
R1157 VTAIL.n334 VTAIL.n333 9.45567
R1158 VTAIL.n82 VTAIL.n81 9.45567
R1159 VTAIL.n252 VTAIL.n251 9.45567
R1160 VTAIL.n168 VTAIL.n167 9.45567
R1161 VTAIL.n333 VTAIL.n332 9.3005
R1162 VTAIL.n256 VTAIL.n255 9.3005
R1163 VTAIL.n301 VTAIL.n300 9.3005
R1164 VTAIL.n299 VTAIL.n298 9.3005
R1165 VTAIL.n272 VTAIL.n271 9.3005
R1166 VTAIL.n293 VTAIL.n292 9.3005
R1167 VTAIL.n291 VTAIL.n290 9.3005
R1168 VTAIL.n276 VTAIL.n275 9.3005
R1169 VTAIL.n285 VTAIL.n284 9.3005
R1170 VTAIL.n283 VTAIL.n282 9.3005
R1171 VTAIL.n268 VTAIL.n267 9.3005
R1172 VTAIL.n307 VTAIL.n306 9.3005
R1173 VTAIL.n309 VTAIL.n308 9.3005
R1174 VTAIL.n264 VTAIL.n263 9.3005
R1175 VTAIL.n315 VTAIL.n314 9.3005
R1176 VTAIL.n317 VTAIL.n316 9.3005
R1177 VTAIL.n260 VTAIL.n259 9.3005
R1178 VTAIL.n324 VTAIL.n323 9.3005
R1179 VTAIL.n326 VTAIL.n325 9.3005
R1180 VTAIL.n81 VTAIL.n80 9.3005
R1181 VTAIL.n4 VTAIL.n3 9.3005
R1182 VTAIL.n49 VTAIL.n48 9.3005
R1183 VTAIL.n47 VTAIL.n46 9.3005
R1184 VTAIL.n20 VTAIL.n19 9.3005
R1185 VTAIL.n41 VTAIL.n40 9.3005
R1186 VTAIL.n39 VTAIL.n38 9.3005
R1187 VTAIL.n24 VTAIL.n23 9.3005
R1188 VTAIL.n33 VTAIL.n32 9.3005
R1189 VTAIL.n31 VTAIL.n30 9.3005
R1190 VTAIL.n16 VTAIL.n15 9.3005
R1191 VTAIL.n55 VTAIL.n54 9.3005
R1192 VTAIL.n57 VTAIL.n56 9.3005
R1193 VTAIL.n12 VTAIL.n11 9.3005
R1194 VTAIL.n63 VTAIL.n62 9.3005
R1195 VTAIL.n65 VTAIL.n64 9.3005
R1196 VTAIL.n8 VTAIL.n7 9.3005
R1197 VTAIL.n72 VTAIL.n71 9.3005
R1198 VTAIL.n74 VTAIL.n73 9.3005
R1199 VTAIL.n226 VTAIL.n225 9.3005
R1200 VTAIL.n228 VTAIL.n227 9.3005
R1201 VTAIL.n183 VTAIL.n182 9.3005
R1202 VTAIL.n234 VTAIL.n233 9.3005
R1203 VTAIL.n236 VTAIL.n235 9.3005
R1204 VTAIL.n178 VTAIL.n177 9.3005
R1205 VTAIL.n242 VTAIL.n241 9.3005
R1206 VTAIL.n244 VTAIL.n243 9.3005
R1207 VTAIL.n251 VTAIL.n250 9.3005
R1208 VTAIL.n174 VTAIL.n173 9.3005
R1209 VTAIL.n187 VTAIL.n186 9.3005
R1210 VTAIL.n220 VTAIL.n219 9.3005
R1211 VTAIL.n218 VTAIL.n217 9.3005
R1212 VTAIL.n191 VTAIL.n190 9.3005
R1213 VTAIL.n212 VTAIL.n211 9.3005
R1214 VTAIL.n210 VTAIL.n209 9.3005
R1215 VTAIL.n195 VTAIL.n194 9.3005
R1216 VTAIL.n204 VTAIL.n203 9.3005
R1217 VTAIL.n202 VTAIL.n201 9.3005
R1218 VTAIL.n142 VTAIL.n141 9.3005
R1219 VTAIL.n144 VTAIL.n143 9.3005
R1220 VTAIL.n99 VTAIL.n98 9.3005
R1221 VTAIL.n150 VTAIL.n149 9.3005
R1222 VTAIL.n152 VTAIL.n151 9.3005
R1223 VTAIL.n94 VTAIL.n93 9.3005
R1224 VTAIL.n158 VTAIL.n157 9.3005
R1225 VTAIL.n160 VTAIL.n159 9.3005
R1226 VTAIL.n167 VTAIL.n166 9.3005
R1227 VTAIL.n90 VTAIL.n89 9.3005
R1228 VTAIL.n103 VTAIL.n102 9.3005
R1229 VTAIL.n136 VTAIL.n135 9.3005
R1230 VTAIL.n134 VTAIL.n133 9.3005
R1231 VTAIL.n107 VTAIL.n106 9.3005
R1232 VTAIL.n128 VTAIL.n127 9.3005
R1233 VTAIL.n126 VTAIL.n125 9.3005
R1234 VTAIL.n111 VTAIL.n110 9.3005
R1235 VTAIL.n120 VTAIL.n119 9.3005
R1236 VTAIL.n118 VTAIL.n117 9.3005
R1237 VTAIL.n297 VTAIL.n272 8.92171
R1238 VTAIL.n310 VTAIL.n264 8.92171
R1239 VTAIL.n45 VTAIL.n20 8.92171
R1240 VTAIL.n58 VTAIL.n12 8.92171
R1241 VTAIL.n229 VTAIL.n183 8.92171
R1242 VTAIL.n216 VTAIL.n191 8.92171
R1243 VTAIL.n145 VTAIL.n99 8.92171
R1244 VTAIL.n132 VTAIL.n107 8.92171
R1245 VTAIL.n298 VTAIL.n270 8.14595
R1246 VTAIL.n309 VTAIL.n266 8.14595
R1247 VTAIL.n46 VTAIL.n18 8.14595
R1248 VTAIL.n57 VTAIL.n14 8.14595
R1249 VTAIL.n228 VTAIL.n185 8.14595
R1250 VTAIL.n217 VTAIL.n189 8.14595
R1251 VTAIL.n144 VTAIL.n101 8.14595
R1252 VTAIL.n133 VTAIL.n105 8.14595
R1253 VTAIL.n302 VTAIL.n301 7.3702
R1254 VTAIL.n306 VTAIL.n305 7.3702
R1255 VTAIL.n50 VTAIL.n49 7.3702
R1256 VTAIL.n54 VTAIL.n53 7.3702
R1257 VTAIL.n225 VTAIL.n224 7.3702
R1258 VTAIL.n221 VTAIL.n220 7.3702
R1259 VTAIL.n141 VTAIL.n140 7.3702
R1260 VTAIL.n137 VTAIL.n136 7.3702
R1261 VTAIL.n302 VTAIL.n268 6.59444
R1262 VTAIL.n305 VTAIL.n268 6.59444
R1263 VTAIL.n50 VTAIL.n16 6.59444
R1264 VTAIL.n53 VTAIL.n16 6.59444
R1265 VTAIL.n224 VTAIL.n187 6.59444
R1266 VTAIL.n221 VTAIL.n187 6.59444
R1267 VTAIL.n140 VTAIL.n103 6.59444
R1268 VTAIL.n137 VTAIL.n103 6.59444
R1269 VTAIL.n301 VTAIL.n270 5.81868
R1270 VTAIL.n306 VTAIL.n266 5.81868
R1271 VTAIL.n49 VTAIL.n18 5.81868
R1272 VTAIL.n54 VTAIL.n14 5.81868
R1273 VTAIL.n225 VTAIL.n185 5.81868
R1274 VTAIL.n220 VTAIL.n189 5.81868
R1275 VTAIL.n141 VTAIL.n101 5.81868
R1276 VTAIL.n136 VTAIL.n105 5.81868
R1277 VTAIL.n298 VTAIL.n297 5.04292
R1278 VTAIL.n310 VTAIL.n309 5.04292
R1279 VTAIL.n46 VTAIL.n45 5.04292
R1280 VTAIL.n58 VTAIL.n57 5.04292
R1281 VTAIL.n229 VTAIL.n228 5.04292
R1282 VTAIL.n217 VTAIL.n216 5.04292
R1283 VTAIL.n145 VTAIL.n144 5.04292
R1284 VTAIL.n133 VTAIL.n132 5.04292
R1285 VTAIL.n294 VTAIL.n272 4.26717
R1286 VTAIL.n313 VTAIL.n264 4.26717
R1287 VTAIL.n42 VTAIL.n20 4.26717
R1288 VTAIL.n61 VTAIL.n12 4.26717
R1289 VTAIL.n232 VTAIL.n183 4.26717
R1290 VTAIL.n213 VTAIL.n191 4.26717
R1291 VTAIL.n148 VTAIL.n99 4.26717
R1292 VTAIL.n129 VTAIL.n107 4.26717
R1293 VTAIL.n283 VTAIL.n279 3.70982
R1294 VTAIL.n31 VTAIL.n27 3.70982
R1295 VTAIL.n202 VTAIL.n198 3.70982
R1296 VTAIL.n118 VTAIL.n114 3.70982
R1297 VTAIL.n293 VTAIL.n274 3.49141
R1298 VTAIL.n314 VTAIL.n262 3.49141
R1299 VTAIL.n41 VTAIL.n22 3.49141
R1300 VTAIL.n62 VTAIL.n10 3.49141
R1301 VTAIL.n233 VTAIL.n181 3.49141
R1302 VTAIL.n212 VTAIL.n193 3.49141
R1303 VTAIL.n149 VTAIL.n97 3.49141
R1304 VTAIL.n128 VTAIL.n109 3.49141
R1305 VTAIL.n290 VTAIL.n289 2.71565
R1306 VTAIL.n318 VTAIL.n317 2.71565
R1307 VTAIL.n38 VTAIL.n37 2.71565
R1308 VTAIL.n66 VTAIL.n65 2.71565
R1309 VTAIL.n237 VTAIL.n236 2.71565
R1310 VTAIL.n209 VTAIL.n208 2.71565
R1311 VTAIL.n153 VTAIL.n152 2.71565
R1312 VTAIL.n125 VTAIL.n124 2.71565
R1313 VTAIL.n0 VTAIL.t11 2.19234
R1314 VTAIL.n0 VTAIL.t3 2.19234
R1315 VTAIL.n84 VTAIL.t5 2.19234
R1316 VTAIL.n84 VTAIL.t10 2.19234
R1317 VTAIL.n170 VTAIL.t9 2.19234
R1318 VTAIL.n170 VTAIL.t7 2.19234
R1319 VTAIL.n86 VTAIL.t0 2.19234
R1320 VTAIL.n86 VTAIL.t1 2.19234
R1321 VTAIL.n286 VTAIL.n276 1.93989
R1322 VTAIL.n322 VTAIL.n260 1.93989
R1323 VTAIL.n334 VTAIL.n254 1.93989
R1324 VTAIL.n34 VTAIL.n24 1.93989
R1325 VTAIL.n70 VTAIL.n8 1.93989
R1326 VTAIL.n82 VTAIL.n2 1.93989
R1327 VTAIL.n252 VTAIL.n172 1.93989
R1328 VTAIL.n240 VTAIL.n178 1.93989
R1329 VTAIL.n205 VTAIL.n195 1.93989
R1330 VTAIL.n168 VTAIL.n88 1.93989
R1331 VTAIL.n156 VTAIL.n94 1.93989
R1332 VTAIL.n121 VTAIL.n111 1.93989
R1333 VTAIL.n285 VTAIL.n278 1.16414
R1334 VTAIL.n323 VTAIL.n258 1.16414
R1335 VTAIL.n332 VTAIL.n331 1.16414
R1336 VTAIL.n33 VTAIL.n26 1.16414
R1337 VTAIL.n71 VTAIL.n6 1.16414
R1338 VTAIL.n80 VTAIL.n79 1.16414
R1339 VTAIL.n250 VTAIL.n249 1.16414
R1340 VTAIL.n241 VTAIL.n176 1.16414
R1341 VTAIL.n204 VTAIL.n197 1.16414
R1342 VTAIL.n166 VTAIL.n165 1.16414
R1343 VTAIL.n157 VTAIL.n92 1.16414
R1344 VTAIL.n120 VTAIL.n113 1.16414
R1345 VTAIL.n171 VTAIL.n169 0.858259
R1346 VTAIL.n83 VTAIL.n1 0.858259
R1347 VTAIL.n169 VTAIL.n87 0.776362
R1348 VTAIL.n253 VTAIL.n171 0.776362
R1349 VTAIL.n85 VTAIL.n83 0.776362
R1350 VTAIL VTAIL.n335 0.524207
R1351 VTAIL.n282 VTAIL.n281 0.388379
R1352 VTAIL.n327 VTAIL.n326 0.388379
R1353 VTAIL.n328 VTAIL.n256 0.388379
R1354 VTAIL.n30 VTAIL.n29 0.388379
R1355 VTAIL.n75 VTAIL.n74 0.388379
R1356 VTAIL.n76 VTAIL.n4 0.388379
R1357 VTAIL.n246 VTAIL.n174 0.388379
R1358 VTAIL.n245 VTAIL.n244 0.388379
R1359 VTAIL.n201 VTAIL.n200 0.388379
R1360 VTAIL.n162 VTAIL.n90 0.388379
R1361 VTAIL.n161 VTAIL.n160 0.388379
R1362 VTAIL.n117 VTAIL.n116 0.388379
R1363 VTAIL VTAIL.n1 0.252655
R1364 VTAIL.n284 VTAIL.n283 0.155672
R1365 VTAIL.n284 VTAIL.n275 0.155672
R1366 VTAIL.n291 VTAIL.n275 0.155672
R1367 VTAIL.n292 VTAIL.n291 0.155672
R1368 VTAIL.n292 VTAIL.n271 0.155672
R1369 VTAIL.n299 VTAIL.n271 0.155672
R1370 VTAIL.n300 VTAIL.n299 0.155672
R1371 VTAIL.n300 VTAIL.n267 0.155672
R1372 VTAIL.n307 VTAIL.n267 0.155672
R1373 VTAIL.n308 VTAIL.n307 0.155672
R1374 VTAIL.n308 VTAIL.n263 0.155672
R1375 VTAIL.n315 VTAIL.n263 0.155672
R1376 VTAIL.n316 VTAIL.n315 0.155672
R1377 VTAIL.n316 VTAIL.n259 0.155672
R1378 VTAIL.n324 VTAIL.n259 0.155672
R1379 VTAIL.n325 VTAIL.n324 0.155672
R1380 VTAIL.n325 VTAIL.n255 0.155672
R1381 VTAIL.n333 VTAIL.n255 0.155672
R1382 VTAIL.n32 VTAIL.n31 0.155672
R1383 VTAIL.n32 VTAIL.n23 0.155672
R1384 VTAIL.n39 VTAIL.n23 0.155672
R1385 VTAIL.n40 VTAIL.n39 0.155672
R1386 VTAIL.n40 VTAIL.n19 0.155672
R1387 VTAIL.n47 VTAIL.n19 0.155672
R1388 VTAIL.n48 VTAIL.n47 0.155672
R1389 VTAIL.n48 VTAIL.n15 0.155672
R1390 VTAIL.n55 VTAIL.n15 0.155672
R1391 VTAIL.n56 VTAIL.n55 0.155672
R1392 VTAIL.n56 VTAIL.n11 0.155672
R1393 VTAIL.n63 VTAIL.n11 0.155672
R1394 VTAIL.n64 VTAIL.n63 0.155672
R1395 VTAIL.n64 VTAIL.n7 0.155672
R1396 VTAIL.n72 VTAIL.n7 0.155672
R1397 VTAIL.n73 VTAIL.n72 0.155672
R1398 VTAIL.n73 VTAIL.n3 0.155672
R1399 VTAIL.n81 VTAIL.n3 0.155672
R1400 VTAIL.n251 VTAIL.n173 0.155672
R1401 VTAIL.n243 VTAIL.n173 0.155672
R1402 VTAIL.n243 VTAIL.n242 0.155672
R1403 VTAIL.n242 VTAIL.n177 0.155672
R1404 VTAIL.n235 VTAIL.n177 0.155672
R1405 VTAIL.n235 VTAIL.n234 0.155672
R1406 VTAIL.n234 VTAIL.n182 0.155672
R1407 VTAIL.n227 VTAIL.n182 0.155672
R1408 VTAIL.n227 VTAIL.n226 0.155672
R1409 VTAIL.n226 VTAIL.n186 0.155672
R1410 VTAIL.n219 VTAIL.n186 0.155672
R1411 VTAIL.n219 VTAIL.n218 0.155672
R1412 VTAIL.n218 VTAIL.n190 0.155672
R1413 VTAIL.n211 VTAIL.n190 0.155672
R1414 VTAIL.n211 VTAIL.n210 0.155672
R1415 VTAIL.n210 VTAIL.n194 0.155672
R1416 VTAIL.n203 VTAIL.n194 0.155672
R1417 VTAIL.n203 VTAIL.n202 0.155672
R1418 VTAIL.n167 VTAIL.n89 0.155672
R1419 VTAIL.n159 VTAIL.n89 0.155672
R1420 VTAIL.n159 VTAIL.n158 0.155672
R1421 VTAIL.n158 VTAIL.n93 0.155672
R1422 VTAIL.n151 VTAIL.n93 0.155672
R1423 VTAIL.n151 VTAIL.n150 0.155672
R1424 VTAIL.n150 VTAIL.n98 0.155672
R1425 VTAIL.n143 VTAIL.n98 0.155672
R1426 VTAIL.n143 VTAIL.n142 0.155672
R1427 VTAIL.n142 VTAIL.n102 0.155672
R1428 VTAIL.n135 VTAIL.n102 0.155672
R1429 VTAIL.n135 VTAIL.n134 0.155672
R1430 VTAIL.n134 VTAIL.n106 0.155672
R1431 VTAIL.n127 VTAIL.n106 0.155672
R1432 VTAIL.n127 VTAIL.n126 0.155672
R1433 VTAIL.n126 VTAIL.n110 0.155672
R1434 VTAIL.n119 VTAIL.n110 0.155672
R1435 VTAIL.n119 VTAIL.n118 0.155672
R1436 VDD1.n76 VDD1.n0 756.745
R1437 VDD1.n157 VDD1.n81 756.745
R1438 VDD1.n77 VDD1.n76 585
R1439 VDD1.n75 VDD1.n74 585
R1440 VDD1.n73 VDD1.n3 585
R1441 VDD1.n7 VDD1.n4 585
R1442 VDD1.n68 VDD1.n67 585
R1443 VDD1.n66 VDD1.n65 585
R1444 VDD1.n9 VDD1.n8 585
R1445 VDD1.n60 VDD1.n59 585
R1446 VDD1.n58 VDD1.n57 585
R1447 VDD1.n13 VDD1.n12 585
R1448 VDD1.n52 VDD1.n51 585
R1449 VDD1.n50 VDD1.n49 585
R1450 VDD1.n17 VDD1.n16 585
R1451 VDD1.n44 VDD1.n43 585
R1452 VDD1.n42 VDD1.n41 585
R1453 VDD1.n21 VDD1.n20 585
R1454 VDD1.n36 VDD1.n35 585
R1455 VDD1.n34 VDD1.n33 585
R1456 VDD1.n25 VDD1.n24 585
R1457 VDD1.n28 VDD1.n27 585
R1458 VDD1.n108 VDD1.n107 585
R1459 VDD1.n105 VDD1.n104 585
R1460 VDD1.n114 VDD1.n113 585
R1461 VDD1.n116 VDD1.n115 585
R1462 VDD1.n101 VDD1.n100 585
R1463 VDD1.n122 VDD1.n121 585
R1464 VDD1.n124 VDD1.n123 585
R1465 VDD1.n97 VDD1.n96 585
R1466 VDD1.n130 VDD1.n129 585
R1467 VDD1.n132 VDD1.n131 585
R1468 VDD1.n93 VDD1.n92 585
R1469 VDD1.n138 VDD1.n137 585
R1470 VDD1.n140 VDD1.n139 585
R1471 VDD1.n89 VDD1.n88 585
R1472 VDD1.n146 VDD1.n145 585
R1473 VDD1.n149 VDD1.n148 585
R1474 VDD1.n147 VDD1.n85 585
R1475 VDD1.n154 VDD1.n84 585
R1476 VDD1.n156 VDD1.n155 585
R1477 VDD1.n158 VDD1.n157 585
R1478 VDD1.t1 VDD1.n26 327.466
R1479 VDD1.t5 VDD1.n106 327.466
R1480 VDD1.n76 VDD1.n75 171.744
R1481 VDD1.n75 VDD1.n3 171.744
R1482 VDD1.n7 VDD1.n3 171.744
R1483 VDD1.n67 VDD1.n7 171.744
R1484 VDD1.n67 VDD1.n66 171.744
R1485 VDD1.n66 VDD1.n8 171.744
R1486 VDD1.n59 VDD1.n8 171.744
R1487 VDD1.n59 VDD1.n58 171.744
R1488 VDD1.n58 VDD1.n12 171.744
R1489 VDD1.n51 VDD1.n12 171.744
R1490 VDD1.n51 VDD1.n50 171.744
R1491 VDD1.n50 VDD1.n16 171.744
R1492 VDD1.n43 VDD1.n16 171.744
R1493 VDD1.n43 VDD1.n42 171.744
R1494 VDD1.n42 VDD1.n20 171.744
R1495 VDD1.n35 VDD1.n20 171.744
R1496 VDD1.n35 VDD1.n34 171.744
R1497 VDD1.n34 VDD1.n24 171.744
R1498 VDD1.n27 VDD1.n24 171.744
R1499 VDD1.n107 VDD1.n104 171.744
R1500 VDD1.n114 VDD1.n104 171.744
R1501 VDD1.n115 VDD1.n114 171.744
R1502 VDD1.n115 VDD1.n100 171.744
R1503 VDD1.n122 VDD1.n100 171.744
R1504 VDD1.n123 VDD1.n122 171.744
R1505 VDD1.n123 VDD1.n96 171.744
R1506 VDD1.n130 VDD1.n96 171.744
R1507 VDD1.n131 VDD1.n130 171.744
R1508 VDD1.n131 VDD1.n92 171.744
R1509 VDD1.n138 VDD1.n92 171.744
R1510 VDD1.n139 VDD1.n138 171.744
R1511 VDD1.n139 VDD1.n88 171.744
R1512 VDD1.n146 VDD1.n88 171.744
R1513 VDD1.n148 VDD1.n146 171.744
R1514 VDD1.n148 VDD1.n147 171.744
R1515 VDD1.n147 VDD1.n84 171.744
R1516 VDD1.n156 VDD1.n84 171.744
R1517 VDD1.n157 VDD1.n156 171.744
R1518 VDD1.n27 VDD1.t1 85.8723
R1519 VDD1.n107 VDD1.t5 85.8723
R1520 VDD1.n163 VDD1.n162 74.5898
R1521 VDD1.n165 VDD1.n164 74.4512
R1522 VDD1 VDD1.n80 53.1891
R1523 VDD1.n163 VDD1.n161 53.0755
R1524 VDD1.n165 VDD1.n163 39.9923
R1525 VDD1.n28 VDD1.n26 16.3895
R1526 VDD1.n108 VDD1.n106 16.3895
R1527 VDD1.n74 VDD1.n73 13.1884
R1528 VDD1.n155 VDD1.n154 13.1884
R1529 VDD1.n77 VDD1.n2 12.8005
R1530 VDD1.n72 VDD1.n4 12.8005
R1531 VDD1.n29 VDD1.n25 12.8005
R1532 VDD1.n109 VDD1.n105 12.8005
R1533 VDD1.n153 VDD1.n85 12.8005
R1534 VDD1.n158 VDD1.n83 12.8005
R1535 VDD1.n78 VDD1.n0 12.0247
R1536 VDD1.n69 VDD1.n68 12.0247
R1537 VDD1.n33 VDD1.n32 12.0247
R1538 VDD1.n113 VDD1.n112 12.0247
R1539 VDD1.n150 VDD1.n149 12.0247
R1540 VDD1.n159 VDD1.n81 12.0247
R1541 VDD1.n65 VDD1.n6 11.249
R1542 VDD1.n36 VDD1.n23 11.249
R1543 VDD1.n116 VDD1.n103 11.249
R1544 VDD1.n145 VDD1.n87 11.249
R1545 VDD1.n64 VDD1.n9 10.4732
R1546 VDD1.n37 VDD1.n21 10.4732
R1547 VDD1.n117 VDD1.n101 10.4732
R1548 VDD1.n144 VDD1.n89 10.4732
R1549 VDD1.n61 VDD1.n60 9.69747
R1550 VDD1.n41 VDD1.n40 9.69747
R1551 VDD1.n121 VDD1.n120 9.69747
R1552 VDD1.n141 VDD1.n140 9.69747
R1553 VDD1.n80 VDD1.n79 9.45567
R1554 VDD1.n161 VDD1.n160 9.45567
R1555 VDD1.n54 VDD1.n53 9.3005
R1556 VDD1.n56 VDD1.n55 9.3005
R1557 VDD1.n11 VDD1.n10 9.3005
R1558 VDD1.n62 VDD1.n61 9.3005
R1559 VDD1.n64 VDD1.n63 9.3005
R1560 VDD1.n6 VDD1.n5 9.3005
R1561 VDD1.n70 VDD1.n69 9.3005
R1562 VDD1.n72 VDD1.n71 9.3005
R1563 VDD1.n79 VDD1.n78 9.3005
R1564 VDD1.n2 VDD1.n1 9.3005
R1565 VDD1.n15 VDD1.n14 9.3005
R1566 VDD1.n48 VDD1.n47 9.3005
R1567 VDD1.n46 VDD1.n45 9.3005
R1568 VDD1.n19 VDD1.n18 9.3005
R1569 VDD1.n40 VDD1.n39 9.3005
R1570 VDD1.n38 VDD1.n37 9.3005
R1571 VDD1.n23 VDD1.n22 9.3005
R1572 VDD1.n32 VDD1.n31 9.3005
R1573 VDD1.n30 VDD1.n29 9.3005
R1574 VDD1.n160 VDD1.n159 9.3005
R1575 VDD1.n83 VDD1.n82 9.3005
R1576 VDD1.n128 VDD1.n127 9.3005
R1577 VDD1.n126 VDD1.n125 9.3005
R1578 VDD1.n99 VDD1.n98 9.3005
R1579 VDD1.n120 VDD1.n119 9.3005
R1580 VDD1.n118 VDD1.n117 9.3005
R1581 VDD1.n103 VDD1.n102 9.3005
R1582 VDD1.n112 VDD1.n111 9.3005
R1583 VDD1.n110 VDD1.n109 9.3005
R1584 VDD1.n95 VDD1.n94 9.3005
R1585 VDD1.n134 VDD1.n133 9.3005
R1586 VDD1.n136 VDD1.n135 9.3005
R1587 VDD1.n91 VDD1.n90 9.3005
R1588 VDD1.n142 VDD1.n141 9.3005
R1589 VDD1.n144 VDD1.n143 9.3005
R1590 VDD1.n87 VDD1.n86 9.3005
R1591 VDD1.n151 VDD1.n150 9.3005
R1592 VDD1.n153 VDD1.n152 9.3005
R1593 VDD1.n57 VDD1.n11 8.92171
R1594 VDD1.n44 VDD1.n19 8.92171
R1595 VDD1.n124 VDD1.n99 8.92171
R1596 VDD1.n137 VDD1.n91 8.92171
R1597 VDD1.n56 VDD1.n13 8.14595
R1598 VDD1.n45 VDD1.n17 8.14595
R1599 VDD1.n125 VDD1.n97 8.14595
R1600 VDD1.n136 VDD1.n93 8.14595
R1601 VDD1.n53 VDD1.n52 7.3702
R1602 VDD1.n49 VDD1.n48 7.3702
R1603 VDD1.n129 VDD1.n128 7.3702
R1604 VDD1.n133 VDD1.n132 7.3702
R1605 VDD1.n52 VDD1.n15 6.59444
R1606 VDD1.n49 VDD1.n15 6.59444
R1607 VDD1.n129 VDD1.n95 6.59444
R1608 VDD1.n132 VDD1.n95 6.59444
R1609 VDD1.n53 VDD1.n13 5.81868
R1610 VDD1.n48 VDD1.n17 5.81868
R1611 VDD1.n128 VDD1.n97 5.81868
R1612 VDD1.n133 VDD1.n93 5.81868
R1613 VDD1.n57 VDD1.n56 5.04292
R1614 VDD1.n45 VDD1.n44 5.04292
R1615 VDD1.n125 VDD1.n124 5.04292
R1616 VDD1.n137 VDD1.n136 5.04292
R1617 VDD1.n60 VDD1.n11 4.26717
R1618 VDD1.n41 VDD1.n19 4.26717
R1619 VDD1.n121 VDD1.n99 4.26717
R1620 VDD1.n140 VDD1.n91 4.26717
R1621 VDD1.n30 VDD1.n26 3.70982
R1622 VDD1.n110 VDD1.n106 3.70982
R1623 VDD1.n61 VDD1.n9 3.49141
R1624 VDD1.n40 VDD1.n21 3.49141
R1625 VDD1.n120 VDD1.n101 3.49141
R1626 VDD1.n141 VDD1.n89 3.49141
R1627 VDD1.n65 VDD1.n64 2.71565
R1628 VDD1.n37 VDD1.n36 2.71565
R1629 VDD1.n117 VDD1.n116 2.71565
R1630 VDD1.n145 VDD1.n144 2.71565
R1631 VDD1.n164 VDD1.t3 2.19234
R1632 VDD1.n164 VDD1.t4 2.19234
R1633 VDD1.n162 VDD1.t0 2.19234
R1634 VDD1.n162 VDD1.t2 2.19234
R1635 VDD1.n80 VDD1.n0 1.93989
R1636 VDD1.n68 VDD1.n6 1.93989
R1637 VDD1.n33 VDD1.n23 1.93989
R1638 VDD1.n113 VDD1.n103 1.93989
R1639 VDD1.n149 VDD1.n87 1.93989
R1640 VDD1.n161 VDD1.n81 1.93989
R1641 VDD1.n78 VDD1.n77 1.16414
R1642 VDD1.n69 VDD1.n4 1.16414
R1643 VDD1.n32 VDD1.n25 1.16414
R1644 VDD1.n112 VDD1.n105 1.16414
R1645 VDD1.n150 VDD1.n85 1.16414
R1646 VDD1.n159 VDD1.n158 1.16414
R1647 VDD1.n74 VDD1.n2 0.388379
R1648 VDD1.n73 VDD1.n72 0.388379
R1649 VDD1.n29 VDD1.n28 0.388379
R1650 VDD1.n109 VDD1.n108 0.388379
R1651 VDD1.n154 VDD1.n153 0.388379
R1652 VDD1.n155 VDD1.n83 0.388379
R1653 VDD1.n79 VDD1.n1 0.155672
R1654 VDD1.n71 VDD1.n1 0.155672
R1655 VDD1.n71 VDD1.n70 0.155672
R1656 VDD1.n70 VDD1.n5 0.155672
R1657 VDD1.n63 VDD1.n5 0.155672
R1658 VDD1.n63 VDD1.n62 0.155672
R1659 VDD1.n62 VDD1.n10 0.155672
R1660 VDD1.n55 VDD1.n10 0.155672
R1661 VDD1.n55 VDD1.n54 0.155672
R1662 VDD1.n54 VDD1.n14 0.155672
R1663 VDD1.n47 VDD1.n14 0.155672
R1664 VDD1.n47 VDD1.n46 0.155672
R1665 VDD1.n46 VDD1.n18 0.155672
R1666 VDD1.n39 VDD1.n18 0.155672
R1667 VDD1.n39 VDD1.n38 0.155672
R1668 VDD1.n38 VDD1.n22 0.155672
R1669 VDD1.n31 VDD1.n22 0.155672
R1670 VDD1.n31 VDD1.n30 0.155672
R1671 VDD1.n111 VDD1.n110 0.155672
R1672 VDD1.n111 VDD1.n102 0.155672
R1673 VDD1.n118 VDD1.n102 0.155672
R1674 VDD1.n119 VDD1.n118 0.155672
R1675 VDD1.n119 VDD1.n98 0.155672
R1676 VDD1.n126 VDD1.n98 0.155672
R1677 VDD1.n127 VDD1.n126 0.155672
R1678 VDD1.n127 VDD1.n94 0.155672
R1679 VDD1.n134 VDD1.n94 0.155672
R1680 VDD1.n135 VDD1.n134 0.155672
R1681 VDD1.n135 VDD1.n90 0.155672
R1682 VDD1.n142 VDD1.n90 0.155672
R1683 VDD1.n143 VDD1.n142 0.155672
R1684 VDD1.n143 VDD1.n86 0.155672
R1685 VDD1.n151 VDD1.n86 0.155672
R1686 VDD1.n152 VDD1.n151 0.155672
R1687 VDD1.n152 VDD1.n82 0.155672
R1688 VDD1.n160 VDD1.n82 0.155672
R1689 VDD1 VDD1.n165 0.136276
R1690 VN.n0 VN.t0 723.184
R1691 VN.n4 VN.t3 723.184
R1692 VN.n1 VN.t4 696.364
R1693 VN.n2 VN.t5 696.364
R1694 VN.n5 VN.t2 696.364
R1695 VN.n6 VN.t1 696.364
R1696 VN.n3 VN.n2 161.3
R1697 VN.n7 VN.n6 161.3
R1698 VN.n2 VN.n1 48.2005
R1699 VN.n6 VN.n5 48.2005
R1700 VN.n7 VN.n4 45.1367
R1701 VN.n3 VN.n0 45.1367
R1702 VN VN.n7 43.2751
R1703 VN.n5 VN.n4 13.3799
R1704 VN.n1 VN.n0 13.3799
R1705 VN VN.n3 0.0516364
R1706 VDD2.n159 VDD2.n83 756.745
R1707 VDD2.n76 VDD2.n0 756.745
R1708 VDD2.n160 VDD2.n159 585
R1709 VDD2.n158 VDD2.n157 585
R1710 VDD2.n156 VDD2.n86 585
R1711 VDD2.n90 VDD2.n87 585
R1712 VDD2.n151 VDD2.n150 585
R1713 VDD2.n149 VDD2.n148 585
R1714 VDD2.n92 VDD2.n91 585
R1715 VDD2.n143 VDD2.n142 585
R1716 VDD2.n141 VDD2.n140 585
R1717 VDD2.n96 VDD2.n95 585
R1718 VDD2.n135 VDD2.n134 585
R1719 VDD2.n133 VDD2.n132 585
R1720 VDD2.n100 VDD2.n99 585
R1721 VDD2.n127 VDD2.n126 585
R1722 VDD2.n125 VDD2.n124 585
R1723 VDD2.n104 VDD2.n103 585
R1724 VDD2.n119 VDD2.n118 585
R1725 VDD2.n117 VDD2.n116 585
R1726 VDD2.n108 VDD2.n107 585
R1727 VDD2.n111 VDD2.n110 585
R1728 VDD2.n27 VDD2.n26 585
R1729 VDD2.n24 VDD2.n23 585
R1730 VDD2.n33 VDD2.n32 585
R1731 VDD2.n35 VDD2.n34 585
R1732 VDD2.n20 VDD2.n19 585
R1733 VDD2.n41 VDD2.n40 585
R1734 VDD2.n43 VDD2.n42 585
R1735 VDD2.n16 VDD2.n15 585
R1736 VDD2.n49 VDD2.n48 585
R1737 VDD2.n51 VDD2.n50 585
R1738 VDD2.n12 VDD2.n11 585
R1739 VDD2.n57 VDD2.n56 585
R1740 VDD2.n59 VDD2.n58 585
R1741 VDD2.n8 VDD2.n7 585
R1742 VDD2.n65 VDD2.n64 585
R1743 VDD2.n68 VDD2.n67 585
R1744 VDD2.n66 VDD2.n4 585
R1745 VDD2.n73 VDD2.n3 585
R1746 VDD2.n75 VDD2.n74 585
R1747 VDD2.n77 VDD2.n76 585
R1748 VDD2.t4 VDD2.n109 327.466
R1749 VDD2.t5 VDD2.n25 327.466
R1750 VDD2.n159 VDD2.n158 171.744
R1751 VDD2.n158 VDD2.n86 171.744
R1752 VDD2.n90 VDD2.n86 171.744
R1753 VDD2.n150 VDD2.n90 171.744
R1754 VDD2.n150 VDD2.n149 171.744
R1755 VDD2.n149 VDD2.n91 171.744
R1756 VDD2.n142 VDD2.n91 171.744
R1757 VDD2.n142 VDD2.n141 171.744
R1758 VDD2.n141 VDD2.n95 171.744
R1759 VDD2.n134 VDD2.n95 171.744
R1760 VDD2.n134 VDD2.n133 171.744
R1761 VDD2.n133 VDD2.n99 171.744
R1762 VDD2.n126 VDD2.n99 171.744
R1763 VDD2.n126 VDD2.n125 171.744
R1764 VDD2.n125 VDD2.n103 171.744
R1765 VDD2.n118 VDD2.n103 171.744
R1766 VDD2.n118 VDD2.n117 171.744
R1767 VDD2.n117 VDD2.n107 171.744
R1768 VDD2.n110 VDD2.n107 171.744
R1769 VDD2.n26 VDD2.n23 171.744
R1770 VDD2.n33 VDD2.n23 171.744
R1771 VDD2.n34 VDD2.n33 171.744
R1772 VDD2.n34 VDD2.n19 171.744
R1773 VDD2.n41 VDD2.n19 171.744
R1774 VDD2.n42 VDD2.n41 171.744
R1775 VDD2.n42 VDD2.n15 171.744
R1776 VDD2.n49 VDD2.n15 171.744
R1777 VDD2.n50 VDD2.n49 171.744
R1778 VDD2.n50 VDD2.n11 171.744
R1779 VDD2.n57 VDD2.n11 171.744
R1780 VDD2.n58 VDD2.n57 171.744
R1781 VDD2.n58 VDD2.n7 171.744
R1782 VDD2.n65 VDD2.n7 171.744
R1783 VDD2.n67 VDD2.n65 171.744
R1784 VDD2.n67 VDD2.n66 171.744
R1785 VDD2.n66 VDD2.n3 171.744
R1786 VDD2.n75 VDD2.n3 171.744
R1787 VDD2.n76 VDD2.n75 171.744
R1788 VDD2.n110 VDD2.t4 85.8723
R1789 VDD2.n26 VDD2.t5 85.8723
R1790 VDD2.n82 VDD2.n81 74.5898
R1791 VDD2 VDD2.n165 74.587
R1792 VDD2.n82 VDD2.n80 53.0755
R1793 VDD2.n164 VDD2.n163 52.549
R1794 VDD2.n164 VDD2.n82 39.0213
R1795 VDD2.n111 VDD2.n109 16.3895
R1796 VDD2.n27 VDD2.n25 16.3895
R1797 VDD2.n157 VDD2.n156 13.1884
R1798 VDD2.n74 VDD2.n73 13.1884
R1799 VDD2.n160 VDD2.n85 12.8005
R1800 VDD2.n155 VDD2.n87 12.8005
R1801 VDD2.n112 VDD2.n108 12.8005
R1802 VDD2.n28 VDD2.n24 12.8005
R1803 VDD2.n72 VDD2.n4 12.8005
R1804 VDD2.n77 VDD2.n2 12.8005
R1805 VDD2.n161 VDD2.n83 12.0247
R1806 VDD2.n152 VDD2.n151 12.0247
R1807 VDD2.n116 VDD2.n115 12.0247
R1808 VDD2.n32 VDD2.n31 12.0247
R1809 VDD2.n69 VDD2.n68 12.0247
R1810 VDD2.n78 VDD2.n0 12.0247
R1811 VDD2.n148 VDD2.n89 11.249
R1812 VDD2.n119 VDD2.n106 11.249
R1813 VDD2.n35 VDD2.n22 11.249
R1814 VDD2.n64 VDD2.n6 11.249
R1815 VDD2.n147 VDD2.n92 10.4732
R1816 VDD2.n120 VDD2.n104 10.4732
R1817 VDD2.n36 VDD2.n20 10.4732
R1818 VDD2.n63 VDD2.n8 10.4732
R1819 VDD2.n144 VDD2.n143 9.69747
R1820 VDD2.n124 VDD2.n123 9.69747
R1821 VDD2.n40 VDD2.n39 9.69747
R1822 VDD2.n60 VDD2.n59 9.69747
R1823 VDD2.n163 VDD2.n162 9.45567
R1824 VDD2.n80 VDD2.n79 9.45567
R1825 VDD2.n137 VDD2.n136 9.3005
R1826 VDD2.n139 VDD2.n138 9.3005
R1827 VDD2.n94 VDD2.n93 9.3005
R1828 VDD2.n145 VDD2.n144 9.3005
R1829 VDD2.n147 VDD2.n146 9.3005
R1830 VDD2.n89 VDD2.n88 9.3005
R1831 VDD2.n153 VDD2.n152 9.3005
R1832 VDD2.n155 VDD2.n154 9.3005
R1833 VDD2.n162 VDD2.n161 9.3005
R1834 VDD2.n85 VDD2.n84 9.3005
R1835 VDD2.n98 VDD2.n97 9.3005
R1836 VDD2.n131 VDD2.n130 9.3005
R1837 VDD2.n129 VDD2.n128 9.3005
R1838 VDD2.n102 VDD2.n101 9.3005
R1839 VDD2.n123 VDD2.n122 9.3005
R1840 VDD2.n121 VDD2.n120 9.3005
R1841 VDD2.n106 VDD2.n105 9.3005
R1842 VDD2.n115 VDD2.n114 9.3005
R1843 VDD2.n113 VDD2.n112 9.3005
R1844 VDD2.n79 VDD2.n78 9.3005
R1845 VDD2.n2 VDD2.n1 9.3005
R1846 VDD2.n47 VDD2.n46 9.3005
R1847 VDD2.n45 VDD2.n44 9.3005
R1848 VDD2.n18 VDD2.n17 9.3005
R1849 VDD2.n39 VDD2.n38 9.3005
R1850 VDD2.n37 VDD2.n36 9.3005
R1851 VDD2.n22 VDD2.n21 9.3005
R1852 VDD2.n31 VDD2.n30 9.3005
R1853 VDD2.n29 VDD2.n28 9.3005
R1854 VDD2.n14 VDD2.n13 9.3005
R1855 VDD2.n53 VDD2.n52 9.3005
R1856 VDD2.n55 VDD2.n54 9.3005
R1857 VDD2.n10 VDD2.n9 9.3005
R1858 VDD2.n61 VDD2.n60 9.3005
R1859 VDD2.n63 VDD2.n62 9.3005
R1860 VDD2.n6 VDD2.n5 9.3005
R1861 VDD2.n70 VDD2.n69 9.3005
R1862 VDD2.n72 VDD2.n71 9.3005
R1863 VDD2.n140 VDD2.n94 8.92171
R1864 VDD2.n127 VDD2.n102 8.92171
R1865 VDD2.n43 VDD2.n18 8.92171
R1866 VDD2.n56 VDD2.n10 8.92171
R1867 VDD2.n139 VDD2.n96 8.14595
R1868 VDD2.n128 VDD2.n100 8.14595
R1869 VDD2.n44 VDD2.n16 8.14595
R1870 VDD2.n55 VDD2.n12 8.14595
R1871 VDD2.n136 VDD2.n135 7.3702
R1872 VDD2.n132 VDD2.n131 7.3702
R1873 VDD2.n48 VDD2.n47 7.3702
R1874 VDD2.n52 VDD2.n51 7.3702
R1875 VDD2.n135 VDD2.n98 6.59444
R1876 VDD2.n132 VDD2.n98 6.59444
R1877 VDD2.n48 VDD2.n14 6.59444
R1878 VDD2.n51 VDD2.n14 6.59444
R1879 VDD2.n136 VDD2.n96 5.81868
R1880 VDD2.n131 VDD2.n100 5.81868
R1881 VDD2.n47 VDD2.n16 5.81868
R1882 VDD2.n52 VDD2.n12 5.81868
R1883 VDD2.n140 VDD2.n139 5.04292
R1884 VDD2.n128 VDD2.n127 5.04292
R1885 VDD2.n44 VDD2.n43 5.04292
R1886 VDD2.n56 VDD2.n55 5.04292
R1887 VDD2.n143 VDD2.n94 4.26717
R1888 VDD2.n124 VDD2.n102 4.26717
R1889 VDD2.n40 VDD2.n18 4.26717
R1890 VDD2.n59 VDD2.n10 4.26717
R1891 VDD2.n113 VDD2.n109 3.70982
R1892 VDD2.n29 VDD2.n25 3.70982
R1893 VDD2.n144 VDD2.n92 3.49141
R1894 VDD2.n123 VDD2.n104 3.49141
R1895 VDD2.n39 VDD2.n20 3.49141
R1896 VDD2.n60 VDD2.n8 3.49141
R1897 VDD2.n148 VDD2.n147 2.71565
R1898 VDD2.n120 VDD2.n119 2.71565
R1899 VDD2.n36 VDD2.n35 2.71565
R1900 VDD2.n64 VDD2.n63 2.71565
R1901 VDD2.n165 VDD2.t3 2.19234
R1902 VDD2.n165 VDD2.t2 2.19234
R1903 VDD2.n81 VDD2.t1 2.19234
R1904 VDD2.n81 VDD2.t0 2.19234
R1905 VDD2.n163 VDD2.n83 1.93989
R1906 VDD2.n151 VDD2.n89 1.93989
R1907 VDD2.n116 VDD2.n106 1.93989
R1908 VDD2.n32 VDD2.n22 1.93989
R1909 VDD2.n68 VDD2.n6 1.93989
R1910 VDD2.n80 VDD2.n0 1.93989
R1911 VDD2.n161 VDD2.n160 1.16414
R1912 VDD2.n152 VDD2.n87 1.16414
R1913 VDD2.n115 VDD2.n108 1.16414
R1914 VDD2.n31 VDD2.n24 1.16414
R1915 VDD2.n69 VDD2.n4 1.16414
R1916 VDD2.n78 VDD2.n77 1.16414
R1917 VDD2 VDD2.n164 0.640586
R1918 VDD2.n157 VDD2.n85 0.388379
R1919 VDD2.n156 VDD2.n155 0.388379
R1920 VDD2.n112 VDD2.n111 0.388379
R1921 VDD2.n28 VDD2.n27 0.388379
R1922 VDD2.n73 VDD2.n72 0.388379
R1923 VDD2.n74 VDD2.n2 0.388379
R1924 VDD2.n162 VDD2.n84 0.155672
R1925 VDD2.n154 VDD2.n84 0.155672
R1926 VDD2.n154 VDD2.n153 0.155672
R1927 VDD2.n153 VDD2.n88 0.155672
R1928 VDD2.n146 VDD2.n88 0.155672
R1929 VDD2.n146 VDD2.n145 0.155672
R1930 VDD2.n145 VDD2.n93 0.155672
R1931 VDD2.n138 VDD2.n93 0.155672
R1932 VDD2.n138 VDD2.n137 0.155672
R1933 VDD2.n137 VDD2.n97 0.155672
R1934 VDD2.n130 VDD2.n97 0.155672
R1935 VDD2.n130 VDD2.n129 0.155672
R1936 VDD2.n129 VDD2.n101 0.155672
R1937 VDD2.n122 VDD2.n101 0.155672
R1938 VDD2.n122 VDD2.n121 0.155672
R1939 VDD2.n121 VDD2.n105 0.155672
R1940 VDD2.n114 VDD2.n105 0.155672
R1941 VDD2.n114 VDD2.n113 0.155672
R1942 VDD2.n30 VDD2.n29 0.155672
R1943 VDD2.n30 VDD2.n21 0.155672
R1944 VDD2.n37 VDD2.n21 0.155672
R1945 VDD2.n38 VDD2.n37 0.155672
R1946 VDD2.n38 VDD2.n17 0.155672
R1947 VDD2.n45 VDD2.n17 0.155672
R1948 VDD2.n46 VDD2.n45 0.155672
R1949 VDD2.n46 VDD2.n13 0.155672
R1950 VDD2.n53 VDD2.n13 0.155672
R1951 VDD2.n54 VDD2.n53 0.155672
R1952 VDD2.n54 VDD2.n9 0.155672
R1953 VDD2.n61 VDD2.n9 0.155672
R1954 VDD2.n62 VDD2.n61 0.155672
R1955 VDD2.n62 VDD2.n5 0.155672
R1956 VDD2.n70 VDD2.n5 0.155672
R1957 VDD2.n71 VDD2.n70 0.155672
R1958 VDD2.n71 VDD2.n1 0.155672
R1959 VDD2.n79 VDD2.n1 0.155672
C0 B VP 1.11448f
C1 B VTAIL 3.11021f
C2 VDD2 VN 4.74636f
C3 VDD1 VP 4.87977f
C4 VDD1 VTAIL 12.862599f
C5 VDD1 B 1.7229f
C6 VN w_n1690_n3934# 2.75949f
C7 VDD2 VP 0.287181f
C8 VDD2 VTAIL 12.8935f
C9 VDD2 B 1.74882f
C10 VP w_n1690_n3934# 2.97233f
C11 VTAIL w_n1690_n3934# 3.40529f
C12 VDD2 VDD1 0.665581f
C13 VP VN 5.47787f
C14 VN VTAIL 4.28f
C15 B w_n1690_n3934# 7.66813f
C16 VDD1 w_n1690_n3934# 1.98615f
C17 B VN 0.769349f
C18 VDD1 VN 0.14802f
C19 VP VTAIL 4.29478f
C20 VDD2 w_n1690_n3934# 2.00618f
C21 VDD2 VSUBS 1.463378f
C22 VDD1 VSUBS 1.203877f
C23 VTAIL VSUBS 0.794408f
C24 VN VSUBS 4.671071f
C25 VP VSUBS 1.478588f
C26 B VSUBS 2.864439f
C27 w_n1690_n3934# VSUBS 81.5459f
C28 VDD2.n0 VSUBS 0.029294f
C29 VDD2.n1 VSUBS 0.026867f
C30 VDD2.n2 VSUBS 0.014437f
C31 VDD2.n3 VSUBS 0.034124f
C32 VDD2.n4 VSUBS 0.015286f
C33 VDD2.n5 VSUBS 0.026867f
C34 VDD2.n6 VSUBS 0.014437f
C35 VDD2.n7 VSUBS 0.034124f
C36 VDD2.n8 VSUBS 0.015286f
C37 VDD2.n9 VSUBS 0.026867f
C38 VDD2.n10 VSUBS 0.014437f
C39 VDD2.n11 VSUBS 0.034124f
C40 VDD2.n12 VSUBS 0.015286f
C41 VDD2.n13 VSUBS 0.026867f
C42 VDD2.n14 VSUBS 0.014437f
C43 VDD2.n15 VSUBS 0.034124f
C44 VDD2.n16 VSUBS 0.015286f
C45 VDD2.n17 VSUBS 0.026867f
C46 VDD2.n18 VSUBS 0.014437f
C47 VDD2.n19 VSUBS 0.034124f
C48 VDD2.n20 VSUBS 0.015286f
C49 VDD2.n21 VSUBS 0.026867f
C50 VDD2.n22 VSUBS 0.014437f
C51 VDD2.n23 VSUBS 0.034124f
C52 VDD2.n24 VSUBS 0.015286f
C53 VDD2.n25 VSUBS 0.188039f
C54 VDD2.t5 VSUBS 0.073041f
C55 VDD2.n26 VSUBS 0.025593f
C56 VDD2.n27 VSUBS 0.021708f
C57 VDD2.n28 VSUBS 0.014437f
C58 VDD2.n29 VSUBS 1.69475f
C59 VDD2.n30 VSUBS 0.026867f
C60 VDD2.n31 VSUBS 0.014437f
C61 VDD2.n32 VSUBS 0.015286f
C62 VDD2.n33 VSUBS 0.034124f
C63 VDD2.n34 VSUBS 0.034124f
C64 VDD2.n35 VSUBS 0.015286f
C65 VDD2.n36 VSUBS 0.014437f
C66 VDD2.n37 VSUBS 0.026867f
C67 VDD2.n38 VSUBS 0.026867f
C68 VDD2.n39 VSUBS 0.014437f
C69 VDD2.n40 VSUBS 0.015286f
C70 VDD2.n41 VSUBS 0.034124f
C71 VDD2.n42 VSUBS 0.034124f
C72 VDD2.n43 VSUBS 0.015286f
C73 VDD2.n44 VSUBS 0.014437f
C74 VDD2.n45 VSUBS 0.026867f
C75 VDD2.n46 VSUBS 0.026867f
C76 VDD2.n47 VSUBS 0.014437f
C77 VDD2.n48 VSUBS 0.015286f
C78 VDD2.n49 VSUBS 0.034124f
C79 VDD2.n50 VSUBS 0.034124f
C80 VDD2.n51 VSUBS 0.015286f
C81 VDD2.n52 VSUBS 0.014437f
C82 VDD2.n53 VSUBS 0.026867f
C83 VDD2.n54 VSUBS 0.026867f
C84 VDD2.n55 VSUBS 0.014437f
C85 VDD2.n56 VSUBS 0.015286f
C86 VDD2.n57 VSUBS 0.034124f
C87 VDD2.n58 VSUBS 0.034124f
C88 VDD2.n59 VSUBS 0.015286f
C89 VDD2.n60 VSUBS 0.014437f
C90 VDD2.n61 VSUBS 0.026867f
C91 VDD2.n62 VSUBS 0.026867f
C92 VDD2.n63 VSUBS 0.014437f
C93 VDD2.n64 VSUBS 0.015286f
C94 VDD2.n65 VSUBS 0.034124f
C95 VDD2.n66 VSUBS 0.034124f
C96 VDD2.n67 VSUBS 0.034124f
C97 VDD2.n68 VSUBS 0.015286f
C98 VDD2.n69 VSUBS 0.014437f
C99 VDD2.n70 VSUBS 0.026867f
C100 VDD2.n71 VSUBS 0.026867f
C101 VDD2.n72 VSUBS 0.014437f
C102 VDD2.n73 VSUBS 0.014861f
C103 VDD2.n74 VSUBS 0.014861f
C104 VDD2.n75 VSUBS 0.034124f
C105 VDD2.n76 VSUBS 0.081839f
C106 VDD2.n77 VSUBS 0.015286f
C107 VDD2.n78 VSUBS 0.014437f
C108 VDD2.n79 VSUBS 0.069074f
C109 VDD2.n80 VSUBS 0.060845f
C110 VDD2.t1 VSUBS 0.314852f
C111 VDD2.t0 VSUBS 0.314852f
C112 VDD2.n81 VSUBS 2.56624f
C113 VDD2.n82 VSUBS 2.39734f
C114 VDD2.n83 VSUBS 0.029294f
C115 VDD2.n84 VSUBS 0.026867f
C116 VDD2.n85 VSUBS 0.014437f
C117 VDD2.n86 VSUBS 0.034124f
C118 VDD2.n87 VSUBS 0.015286f
C119 VDD2.n88 VSUBS 0.026867f
C120 VDD2.n89 VSUBS 0.014437f
C121 VDD2.n90 VSUBS 0.034124f
C122 VDD2.n91 VSUBS 0.034124f
C123 VDD2.n92 VSUBS 0.015286f
C124 VDD2.n93 VSUBS 0.026867f
C125 VDD2.n94 VSUBS 0.014437f
C126 VDD2.n95 VSUBS 0.034124f
C127 VDD2.n96 VSUBS 0.015286f
C128 VDD2.n97 VSUBS 0.026867f
C129 VDD2.n98 VSUBS 0.014437f
C130 VDD2.n99 VSUBS 0.034124f
C131 VDD2.n100 VSUBS 0.015286f
C132 VDD2.n101 VSUBS 0.026867f
C133 VDD2.n102 VSUBS 0.014437f
C134 VDD2.n103 VSUBS 0.034124f
C135 VDD2.n104 VSUBS 0.015286f
C136 VDD2.n105 VSUBS 0.026867f
C137 VDD2.n106 VSUBS 0.014437f
C138 VDD2.n107 VSUBS 0.034124f
C139 VDD2.n108 VSUBS 0.015286f
C140 VDD2.n109 VSUBS 0.188039f
C141 VDD2.t4 VSUBS 0.073041f
C142 VDD2.n110 VSUBS 0.025593f
C143 VDD2.n111 VSUBS 0.021708f
C144 VDD2.n112 VSUBS 0.014437f
C145 VDD2.n113 VSUBS 1.69475f
C146 VDD2.n114 VSUBS 0.026867f
C147 VDD2.n115 VSUBS 0.014437f
C148 VDD2.n116 VSUBS 0.015286f
C149 VDD2.n117 VSUBS 0.034124f
C150 VDD2.n118 VSUBS 0.034124f
C151 VDD2.n119 VSUBS 0.015286f
C152 VDD2.n120 VSUBS 0.014437f
C153 VDD2.n121 VSUBS 0.026867f
C154 VDD2.n122 VSUBS 0.026867f
C155 VDD2.n123 VSUBS 0.014437f
C156 VDD2.n124 VSUBS 0.015286f
C157 VDD2.n125 VSUBS 0.034124f
C158 VDD2.n126 VSUBS 0.034124f
C159 VDD2.n127 VSUBS 0.015286f
C160 VDD2.n128 VSUBS 0.014437f
C161 VDD2.n129 VSUBS 0.026867f
C162 VDD2.n130 VSUBS 0.026867f
C163 VDD2.n131 VSUBS 0.014437f
C164 VDD2.n132 VSUBS 0.015286f
C165 VDD2.n133 VSUBS 0.034124f
C166 VDD2.n134 VSUBS 0.034124f
C167 VDD2.n135 VSUBS 0.015286f
C168 VDD2.n136 VSUBS 0.014437f
C169 VDD2.n137 VSUBS 0.026867f
C170 VDD2.n138 VSUBS 0.026867f
C171 VDD2.n139 VSUBS 0.014437f
C172 VDD2.n140 VSUBS 0.015286f
C173 VDD2.n141 VSUBS 0.034124f
C174 VDD2.n142 VSUBS 0.034124f
C175 VDD2.n143 VSUBS 0.015286f
C176 VDD2.n144 VSUBS 0.014437f
C177 VDD2.n145 VSUBS 0.026867f
C178 VDD2.n146 VSUBS 0.026867f
C179 VDD2.n147 VSUBS 0.014437f
C180 VDD2.n148 VSUBS 0.015286f
C181 VDD2.n149 VSUBS 0.034124f
C182 VDD2.n150 VSUBS 0.034124f
C183 VDD2.n151 VSUBS 0.015286f
C184 VDD2.n152 VSUBS 0.014437f
C185 VDD2.n153 VSUBS 0.026867f
C186 VDD2.n154 VSUBS 0.026867f
C187 VDD2.n155 VSUBS 0.014437f
C188 VDD2.n156 VSUBS 0.014861f
C189 VDD2.n157 VSUBS 0.014861f
C190 VDD2.n158 VSUBS 0.034124f
C191 VDD2.n159 VSUBS 0.081839f
C192 VDD2.n160 VSUBS 0.015286f
C193 VDD2.n161 VSUBS 0.014437f
C194 VDD2.n162 VSUBS 0.069074f
C195 VDD2.n163 VSUBS 0.059828f
C196 VDD2.n164 VSUBS 2.39884f
C197 VDD2.t3 VSUBS 0.314852f
C198 VDD2.t2 VSUBS 0.314852f
C199 VDD2.n165 VSUBS 2.5662f
C200 VN.t0 VSUBS 1.43002f
C201 VN.n0 VSUBS 0.529269f
C202 VN.t4 VSUBS 1.40968f
C203 VN.n1 VSUBS 0.561694f
C204 VN.t5 VSUBS 1.40968f
C205 VN.n2 VSUBS 0.548383f
C206 VN.n3 VSUBS 0.2336f
C207 VN.t3 VSUBS 1.43002f
C208 VN.n4 VSUBS 0.529269f
C209 VN.t2 VSUBS 1.40968f
C210 VN.n5 VSUBS 0.561694f
C211 VN.t1 VSUBS 1.40968f
C212 VN.n6 VSUBS 0.548383f
C213 VN.n7 VSUBS 2.73393f
C214 VDD1.n0 VSUBS 0.02647f
C215 VDD1.n1 VSUBS 0.024276f
C216 VDD1.n2 VSUBS 0.013045f
C217 VDD1.n3 VSUBS 0.030834f
C218 VDD1.n4 VSUBS 0.013812f
C219 VDD1.n5 VSUBS 0.024276f
C220 VDD1.n6 VSUBS 0.013045f
C221 VDD1.n7 VSUBS 0.030834f
C222 VDD1.n8 VSUBS 0.030834f
C223 VDD1.n9 VSUBS 0.013812f
C224 VDD1.n10 VSUBS 0.024276f
C225 VDD1.n11 VSUBS 0.013045f
C226 VDD1.n12 VSUBS 0.030834f
C227 VDD1.n13 VSUBS 0.013812f
C228 VDD1.n14 VSUBS 0.024276f
C229 VDD1.n15 VSUBS 0.013045f
C230 VDD1.n16 VSUBS 0.030834f
C231 VDD1.n17 VSUBS 0.013812f
C232 VDD1.n18 VSUBS 0.024276f
C233 VDD1.n19 VSUBS 0.013045f
C234 VDD1.n20 VSUBS 0.030834f
C235 VDD1.n21 VSUBS 0.013812f
C236 VDD1.n22 VSUBS 0.024276f
C237 VDD1.n23 VSUBS 0.013045f
C238 VDD1.n24 VSUBS 0.030834f
C239 VDD1.n25 VSUBS 0.013812f
C240 VDD1.n26 VSUBS 0.16991f
C241 VDD1.t1 VSUBS 0.065999f
C242 VDD1.n27 VSUBS 0.023125f
C243 VDD1.n28 VSUBS 0.019615f
C244 VDD1.n29 VSUBS 0.013045f
C245 VDD1.n30 VSUBS 1.53135f
C246 VDD1.n31 VSUBS 0.024276f
C247 VDD1.n32 VSUBS 0.013045f
C248 VDD1.n33 VSUBS 0.013812f
C249 VDD1.n34 VSUBS 0.030834f
C250 VDD1.n35 VSUBS 0.030834f
C251 VDD1.n36 VSUBS 0.013812f
C252 VDD1.n37 VSUBS 0.013045f
C253 VDD1.n38 VSUBS 0.024276f
C254 VDD1.n39 VSUBS 0.024276f
C255 VDD1.n40 VSUBS 0.013045f
C256 VDD1.n41 VSUBS 0.013812f
C257 VDD1.n42 VSUBS 0.030834f
C258 VDD1.n43 VSUBS 0.030834f
C259 VDD1.n44 VSUBS 0.013812f
C260 VDD1.n45 VSUBS 0.013045f
C261 VDD1.n46 VSUBS 0.024276f
C262 VDD1.n47 VSUBS 0.024276f
C263 VDD1.n48 VSUBS 0.013045f
C264 VDD1.n49 VSUBS 0.013812f
C265 VDD1.n50 VSUBS 0.030834f
C266 VDD1.n51 VSUBS 0.030834f
C267 VDD1.n52 VSUBS 0.013812f
C268 VDD1.n53 VSUBS 0.013045f
C269 VDD1.n54 VSUBS 0.024276f
C270 VDD1.n55 VSUBS 0.024276f
C271 VDD1.n56 VSUBS 0.013045f
C272 VDD1.n57 VSUBS 0.013812f
C273 VDD1.n58 VSUBS 0.030834f
C274 VDD1.n59 VSUBS 0.030834f
C275 VDD1.n60 VSUBS 0.013812f
C276 VDD1.n61 VSUBS 0.013045f
C277 VDD1.n62 VSUBS 0.024276f
C278 VDD1.n63 VSUBS 0.024276f
C279 VDD1.n64 VSUBS 0.013045f
C280 VDD1.n65 VSUBS 0.013812f
C281 VDD1.n66 VSUBS 0.030834f
C282 VDD1.n67 VSUBS 0.030834f
C283 VDD1.n68 VSUBS 0.013812f
C284 VDD1.n69 VSUBS 0.013045f
C285 VDD1.n70 VSUBS 0.024276f
C286 VDD1.n71 VSUBS 0.024276f
C287 VDD1.n72 VSUBS 0.013045f
C288 VDD1.n73 VSUBS 0.013429f
C289 VDD1.n74 VSUBS 0.013429f
C290 VDD1.n75 VSUBS 0.030834f
C291 VDD1.n76 VSUBS 0.073949f
C292 VDD1.n77 VSUBS 0.013812f
C293 VDD1.n78 VSUBS 0.013045f
C294 VDD1.n79 VSUBS 0.062415f
C295 VDD1.n80 VSUBS 0.055269f
C296 VDD1.n81 VSUBS 0.02647f
C297 VDD1.n82 VSUBS 0.024276f
C298 VDD1.n83 VSUBS 0.013045f
C299 VDD1.n84 VSUBS 0.030834f
C300 VDD1.n85 VSUBS 0.013812f
C301 VDD1.n86 VSUBS 0.024276f
C302 VDD1.n87 VSUBS 0.013045f
C303 VDD1.n88 VSUBS 0.030834f
C304 VDD1.n89 VSUBS 0.013812f
C305 VDD1.n90 VSUBS 0.024276f
C306 VDD1.n91 VSUBS 0.013045f
C307 VDD1.n92 VSUBS 0.030834f
C308 VDD1.n93 VSUBS 0.013812f
C309 VDD1.n94 VSUBS 0.024276f
C310 VDD1.n95 VSUBS 0.013045f
C311 VDD1.n96 VSUBS 0.030834f
C312 VDD1.n97 VSUBS 0.013812f
C313 VDD1.n98 VSUBS 0.024276f
C314 VDD1.n99 VSUBS 0.013045f
C315 VDD1.n100 VSUBS 0.030834f
C316 VDD1.n101 VSUBS 0.013812f
C317 VDD1.n102 VSUBS 0.024276f
C318 VDD1.n103 VSUBS 0.013045f
C319 VDD1.n104 VSUBS 0.030834f
C320 VDD1.n105 VSUBS 0.013812f
C321 VDD1.n106 VSUBS 0.16991f
C322 VDD1.t5 VSUBS 0.065999f
C323 VDD1.n107 VSUBS 0.023125f
C324 VDD1.n108 VSUBS 0.019615f
C325 VDD1.n109 VSUBS 0.013045f
C326 VDD1.n110 VSUBS 1.53135f
C327 VDD1.n111 VSUBS 0.024276f
C328 VDD1.n112 VSUBS 0.013045f
C329 VDD1.n113 VSUBS 0.013812f
C330 VDD1.n114 VSUBS 0.030834f
C331 VDD1.n115 VSUBS 0.030834f
C332 VDD1.n116 VSUBS 0.013812f
C333 VDD1.n117 VSUBS 0.013045f
C334 VDD1.n118 VSUBS 0.024276f
C335 VDD1.n119 VSUBS 0.024276f
C336 VDD1.n120 VSUBS 0.013045f
C337 VDD1.n121 VSUBS 0.013812f
C338 VDD1.n122 VSUBS 0.030834f
C339 VDD1.n123 VSUBS 0.030834f
C340 VDD1.n124 VSUBS 0.013812f
C341 VDD1.n125 VSUBS 0.013045f
C342 VDD1.n126 VSUBS 0.024276f
C343 VDD1.n127 VSUBS 0.024276f
C344 VDD1.n128 VSUBS 0.013045f
C345 VDD1.n129 VSUBS 0.013812f
C346 VDD1.n130 VSUBS 0.030834f
C347 VDD1.n131 VSUBS 0.030834f
C348 VDD1.n132 VSUBS 0.013812f
C349 VDD1.n133 VSUBS 0.013045f
C350 VDD1.n134 VSUBS 0.024276f
C351 VDD1.n135 VSUBS 0.024276f
C352 VDD1.n136 VSUBS 0.013045f
C353 VDD1.n137 VSUBS 0.013812f
C354 VDD1.n138 VSUBS 0.030834f
C355 VDD1.n139 VSUBS 0.030834f
C356 VDD1.n140 VSUBS 0.013812f
C357 VDD1.n141 VSUBS 0.013045f
C358 VDD1.n142 VSUBS 0.024276f
C359 VDD1.n143 VSUBS 0.024276f
C360 VDD1.n144 VSUBS 0.013045f
C361 VDD1.n145 VSUBS 0.013812f
C362 VDD1.n146 VSUBS 0.030834f
C363 VDD1.n147 VSUBS 0.030834f
C364 VDD1.n148 VSUBS 0.030834f
C365 VDD1.n149 VSUBS 0.013812f
C366 VDD1.n150 VSUBS 0.013045f
C367 VDD1.n151 VSUBS 0.024276f
C368 VDD1.n152 VSUBS 0.024276f
C369 VDD1.n153 VSUBS 0.013045f
C370 VDD1.n154 VSUBS 0.013429f
C371 VDD1.n155 VSUBS 0.013429f
C372 VDD1.n156 VSUBS 0.030834f
C373 VDD1.n157 VSUBS 0.073949f
C374 VDD1.n158 VSUBS 0.013812f
C375 VDD1.n159 VSUBS 0.013045f
C376 VDD1.n160 VSUBS 0.062415f
C377 VDD1.n161 VSUBS 0.054979f
C378 VDD1.t0 VSUBS 0.284497f
C379 VDD1.t2 VSUBS 0.284497f
C380 VDD1.n162 VSUBS 2.31882f
C381 VDD1.n163 VSUBS 2.23888f
C382 VDD1.t3 VSUBS 0.284497f
C383 VDD1.t4 VSUBS 0.284497f
C384 VDD1.n164 VSUBS 2.31782f
C385 VDD1.n165 VSUBS 2.6162f
C386 VTAIL.t11 VSUBS 0.345245f
C387 VTAIL.t3 VSUBS 0.345245f
C388 VTAIL.n0 VSUBS 2.65637f
C389 VTAIL.n1 VSUBS 0.76897f
C390 VTAIL.n2 VSUBS 0.032122f
C391 VTAIL.n3 VSUBS 0.02946f
C392 VTAIL.n4 VSUBS 0.015831f
C393 VTAIL.n5 VSUBS 0.037418f
C394 VTAIL.n6 VSUBS 0.016762f
C395 VTAIL.n7 VSUBS 0.02946f
C396 VTAIL.n8 VSUBS 0.015831f
C397 VTAIL.n9 VSUBS 0.037418f
C398 VTAIL.n10 VSUBS 0.016762f
C399 VTAIL.n11 VSUBS 0.02946f
C400 VTAIL.n12 VSUBS 0.015831f
C401 VTAIL.n13 VSUBS 0.037418f
C402 VTAIL.n14 VSUBS 0.016762f
C403 VTAIL.n15 VSUBS 0.02946f
C404 VTAIL.n16 VSUBS 0.015831f
C405 VTAIL.n17 VSUBS 0.037418f
C406 VTAIL.n18 VSUBS 0.016762f
C407 VTAIL.n19 VSUBS 0.02946f
C408 VTAIL.n20 VSUBS 0.015831f
C409 VTAIL.n21 VSUBS 0.037418f
C410 VTAIL.n22 VSUBS 0.016762f
C411 VTAIL.n23 VSUBS 0.02946f
C412 VTAIL.n24 VSUBS 0.015831f
C413 VTAIL.n25 VSUBS 0.037418f
C414 VTAIL.n26 VSUBS 0.016762f
C415 VTAIL.n27 VSUBS 0.206191f
C416 VTAIL.t8 VSUBS 0.080092f
C417 VTAIL.n28 VSUBS 0.028063f
C418 VTAIL.n29 VSUBS 0.023803f
C419 VTAIL.n30 VSUBS 0.015831f
C420 VTAIL.n31 VSUBS 1.85834f
C421 VTAIL.n32 VSUBS 0.02946f
C422 VTAIL.n33 VSUBS 0.015831f
C423 VTAIL.n34 VSUBS 0.016762f
C424 VTAIL.n35 VSUBS 0.037418f
C425 VTAIL.n36 VSUBS 0.037418f
C426 VTAIL.n37 VSUBS 0.016762f
C427 VTAIL.n38 VSUBS 0.015831f
C428 VTAIL.n39 VSUBS 0.02946f
C429 VTAIL.n40 VSUBS 0.02946f
C430 VTAIL.n41 VSUBS 0.015831f
C431 VTAIL.n42 VSUBS 0.016762f
C432 VTAIL.n43 VSUBS 0.037418f
C433 VTAIL.n44 VSUBS 0.037418f
C434 VTAIL.n45 VSUBS 0.016762f
C435 VTAIL.n46 VSUBS 0.015831f
C436 VTAIL.n47 VSUBS 0.02946f
C437 VTAIL.n48 VSUBS 0.02946f
C438 VTAIL.n49 VSUBS 0.015831f
C439 VTAIL.n50 VSUBS 0.016762f
C440 VTAIL.n51 VSUBS 0.037418f
C441 VTAIL.n52 VSUBS 0.037418f
C442 VTAIL.n53 VSUBS 0.016762f
C443 VTAIL.n54 VSUBS 0.015831f
C444 VTAIL.n55 VSUBS 0.02946f
C445 VTAIL.n56 VSUBS 0.02946f
C446 VTAIL.n57 VSUBS 0.015831f
C447 VTAIL.n58 VSUBS 0.016762f
C448 VTAIL.n59 VSUBS 0.037418f
C449 VTAIL.n60 VSUBS 0.037418f
C450 VTAIL.n61 VSUBS 0.016762f
C451 VTAIL.n62 VSUBS 0.015831f
C452 VTAIL.n63 VSUBS 0.02946f
C453 VTAIL.n64 VSUBS 0.02946f
C454 VTAIL.n65 VSUBS 0.015831f
C455 VTAIL.n66 VSUBS 0.016762f
C456 VTAIL.n67 VSUBS 0.037418f
C457 VTAIL.n68 VSUBS 0.037418f
C458 VTAIL.n69 VSUBS 0.037418f
C459 VTAIL.n70 VSUBS 0.016762f
C460 VTAIL.n71 VSUBS 0.015831f
C461 VTAIL.n72 VSUBS 0.02946f
C462 VTAIL.n73 VSUBS 0.02946f
C463 VTAIL.n74 VSUBS 0.015831f
C464 VTAIL.n75 VSUBS 0.016296f
C465 VTAIL.n76 VSUBS 0.016296f
C466 VTAIL.n77 VSUBS 0.037418f
C467 VTAIL.n78 VSUBS 0.089739f
C468 VTAIL.n79 VSUBS 0.016762f
C469 VTAIL.n80 VSUBS 0.015831f
C470 VTAIL.n81 VSUBS 0.075742f
C471 VTAIL.n82 VSUBS 0.045315f
C472 VTAIL.n83 VSUBS 0.184562f
C473 VTAIL.t5 VSUBS 0.345245f
C474 VTAIL.t10 VSUBS 0.345245f
C475 VTAIL.n84 VSUBS 2.65637f
C476 VTAIL.n85 VSUBS 2.49833f
C477 VTAIL.t0 VSUBS 0.345245f
C478 VTAIL.t1 VSUBS 0.345245f
C479 VTAIL.n86 VSUBS 2.65639f
C480 VTAIL.n87 VSUBS 2.49831f
C481 VTAIL.n88 VSUBS 0.032122f
C482 VTAIL.n89 VSUBS 0.02946f
C483 VTAIL.n90 VSUBS 0.015831f
C484 VTAIL.n91 VSUBS 0.037418f
C485 VTAIL.n92 VSUBS 0.016762f
C486 VTAIL.n93 VSUBS 0.02946f
C487 VTAIL.n94 VSUBS 0.015831f
C488 VTAIL.n95 VSUBS 0.037418f
C489 VTAIL.n96 VSUBS 0.037418f
C490 VTAIL.n97 VSUBS 0.016762f
C491 VTAIL.n98 VSUBS 0.02946f
C492 VTAIL.n99 VSUBS 0.015831f
C493 VTAIL.n100 VSUBS 0.037418f
C494 VTAIL.n101 VSUBS 0.016762f
C495 VTAIL.n102 VSUBS 0.02946f
C496 VTAIL.n103 VSUBS 0.015831f
C497 VTAIL.n104 VSUBS 0.037418f
C498 VTAIL.n105 VSUBS 0.016762f
C499 VTAIL.n106 VSUBS 0.02946f
C500 VTAIL.n107 VSUBS 0.015831f
C501 VTAIL.n108 VSUBS 0.037418f
C502 VTAIL.n109 VSUBS 0.016762f
C503 VTAIL.n110 VSUBS 0.02946f
C504 VTAIL.n111 VSUBS 0.015831f
C505 VTAIL.n112 VSUBS 0.037418f
C506 VTAIL.n113 VSUBS 0.016762f
C507 VTAIL.n114 VSUBS 0.206191f
C508 VTAIL.t4 VSUBS 0.080092f
C509 VTAIL.n115 VSUBS 0.028063f
C510 VTAIL.n116 VSUBS 0.023803f
C511 VTAIL.n117 VSUBS 0.015831f
C512 VTAIL.n118 VSUBS 1.85834f
C513 VTAIL.n119 VSUBS 0.02946f
C514 VTAIL.n120 VSUBS 0.015831f
C515 VTAIL.n121 VSUBS 0.016762f
C516 VTAIL.n122 VSUBS 0.037418f
C517 VTAIL.n123 VSUBS 0.037418f
C518 VTAIL.n124 VSUBS 0.016762f
C519 VTAIL.n125 VSUBS 0.015831f
C520 VTAIL.n126 VSUBS 0.02946f
C521 VTAIL.n127 VSUBS 0.02946f
C522 VTAIL.n128 VSUBS 0.015831f
C523 VTAIL.n129 VSUBS 0.016762f
C524 VTAIL.n130 VSUBS 0.037418f
C525 VTAIL.n131 VSUBS 0.037418f
C526 VTAIL.n132 VSUBS 0.016762f
C527 VTAIL.n133 VSUBS 0.015831f
C528 VTAIL.n134 VSUBS 0.02946f
C529 VTAIL.n135 VSUBS 0.02946f
C530 VTAIL.n136 VSUBS 0.015831f
C531 VTAIL.n137 VSUBS 0.016762f
C532 VTAIL.n138 VSUBS 0.037418f
C533 VTAIL.n139 VSUBS 0.037418f
C534 VTAIL.n140 VSUBS 0.016762f
C535 VTAIL.n141 VSUBS 0.015831f
C536 VTAIL.n142 VSUBS 0.02946f
C537 VTAIL.n143 VSUBS 0.02946f
C538 VTAIL.n144 VSUBS 0.015831f
C539 VTAIL.n145 VSUBS 0.016762f
C540 VTAIL.n146 VSUBS 0.037418f
C541 VTAIL.n147 VSUBS 0.037418f
C542 VTAIL.n148 VSUBS 0.016762f
C543 VTAIL.n149 VSUBS 0.015831f
C544 VTAIL.n150 VSUBS 0.02946f
C545 VTAIL.n151 VSUBS 0.02946f
C546 VTAIL.n152 VSUBS 0.015831f
C547 VTAIL.n153 VSUBS 0.016762f
C548 VTAIL.n154 VSUBS 0.037418f
C549 VTAIL.n155 VSUBS 0.037418f
C550 VTAIL.n156 VSUBS 0.016762f
C551 VTAIL.n157 VSUBS 0.015831f
C552 VTAIL.n158 VSUBS 0.02946f
C553 VTAIL.n159 VSUBS 0.02946f
C554 VTAIL.n160 VSUBS 0.015831f
C555 VTAIL.n161 VSUBS 0.016296f
C556 VTAIL.n162 VSUBS 0.016296f
C557 VTAIL.n163 VSUBS 0.037418f
C558 VTAIL.n164 VSUBS 0.089739f
C559 VTAIL.n165 VSUBS 0.016762f
C560 VTAIL.n166 VSUBS 0.015831f
C561 VTAIL.n167 VSUBS 0.075742f
C562 VTAIL.n168 VSUBS 0.045315f
C563 VTAIL.n169 VSUBS 0.184562f
C564 VTAIL.t9 VSUBS 0.345245f
C565 VTAIL.t7 VSUBS 0.345245f
C566 VTAIL.n170 VSUBS 2.65639f
C567 VTAIL.n171 VSUBS 0.818668f
C568 VTAIL.n172 VSUBS 0.032122f
C569 VTAIL.n173 VSUBS 0.02946f
C570 VTAIL.n174 VSUBS 0.015831f
C571 VTAIL.n175 VSUBS 0.037418f
C572 VTAIL.n176 VSUBS 0.016762f
C573 VTAIL.n177 VSUBS 0.02946f
C574 VTAIL.n178 VSUBS 0.015831f
C575 VTAIL.n179 VSUBS 0.037418f
C576 VTAIL.n180 VSUBS 0.037418f
C577 VTAIL.n181 VSUBS 0.016762f
C578 VTAIL.n182 VSUBS 0.02946f
C579 VTAIL.n183 VSUBS 0.015831f
C580 VTAIL.n184 VSUBS 0.037418f
C581 VTAIL.n185 VSUBS 0.016762f
C582 VTAIL.n186 VSUBS 0.02946f
C583 VTAIL.n187 VSUBS 0.015831f
C584 VTAIL.n188 VSUBS 0.037418f
C585 VTAIL.n189 VSUBS 0.016762f
C586 VTAIL.n190 VSUBS 0.02946f
C587 VTAIL.n191 VSUBS 0.015831f
C588 VTAIL.n192 VSUBS 0.037418f
C589 VTAIL.n193 VSUBS 0.016762f
C590 VTAIL.n194 VSUBS 0.02946f
C591 VTAIL.n195 VSUBS 0.015831f
C592 VTAIL.n196 VSUBS 0.037418f
C593 VTAIL.n197 VSUBS 0.016762f
C594 VTAIL.n198 VSUBS 0.206191f
C595 VTAIL.t6 VSUBS 0.080092f
C596 VTAIL.n199 VSUBS 0.028063f
C597 VTAIL.n200 VSUBS 0.023803f
C598 VTAIL.n201 VSUBS 0.015831f
C599 VTAIL.n202 VSUBS 1.85834f
C600 VTAIL.n203 VSUBS 0.02946f
C601 VTAIL.n204 VSUBS 0.015831f
C602 VTAIL.n205 VSUBS 0.016762f
C603 VTAIL.n206 VSUBS 0.037418f
C604 VTAIL.n207 VSUBS 0.037418f
C605 VTAIL.n208 VSUBS 0.016762f
C606 VTAIL.n209 VSUBS 0.015831f
C607 VTAIL.n210 VSUBS 0.02946f
C608 VTAIL.n211 VSUBS 0.02946f
C609 VTAIL.n212 VSUBS 0.015831f
C610 VTAIL.n213 VSUBS 0.016762f
C611 VTAIL.n214 VSUBS 0.037418f
C612 VTAIL.n215 VSUBS 0.037418f
C613 VTAIL.n216 VSUBS 0.016762f
C614 VTAIL.n217 VSUBS 0.015831f
C615 VTAIL.n218 VSUBS 0.02946f
C616 VTAIL.n219 VSUBS 0.02946f
C617 VTAIL.n220 VSUBS 0.015831f
C618 VTAIL.n221 VSUBS 0.016762f
C619 VTAIL.n222 VSUBS 0.037418f
C620 VTAIL.n223 VSUBS 0.037418f
C621 VTAIL.n224 VSUBS 0.016762f
C622 VTAIL.n225 VSUBS 0.015831f
C623 VTAIL.n226 VSUBS 0.02946f
C624 VTAIL.n227 VSUBS 0.02946f
C625 VTAIL.n228 VSUBS 0.015831f
C626 VTAIL.n229 VSUBS 0.016762f
C627 VTAIL.n230 VSUBS 0.037418f
C628 VTAIL.n231 VSUBS 0.037418f
C629 VTAIL.n232 VSUBS 0.016762f
C630 VTAIL.n233 VSUBS 0.015831f
C631 VTAIL.n234 VSUBS 0.02946f
C632 VTAIL.n235 VSUBS 0.02946f
C633 VTAIL.n236 VSUBS 0.015831f
C634 VTAIL.n237 VSUBS 0.016762f
C635 VTAIL.n238 VSUBS 0.037418f
C636 VTAIL.n239 VSUBS 0.037418f
C637 VTAIL.n240 VSUBS 0.016762f
C638 VTAIL.n241 VSUBS 0.015831f
C639 VTAIL.n242 VSUBS 0.02946f
C640 VTAIL.n243 VSUBS 0.02946f
C641 VTAIL.n244 VSUBS 0.015831f
C642 VTAIL.n245 VSUBS 0.016296f
C643 VTAIL.n246 VSUBS 0.016296f
C644 VTAIL.n247 VSUBS 0.037418f
C645 VTAIL.n248 VSUBS 0.089739f
C646 VTAIL.n249 VSUBS 0.016762f
C647 VTAIL.n250 VSUBS 0.015831f
C648 VTAIL.n251 VSUBS 0.075742f
C649 VTAIL.n252 VSUBS 0.045315f
C650 VTAIL.n253 VSUBS 1.79056f
C651 VTAIL.n254 VSUBS 0.032122f
C652 VTAIL.n255 VSUBS 0.02946f
C653 VTAIL.n256 VSUBS 0.015831f
C654 VTAIL.n257 VSUBS 0.037418f
C655 VTAIL.n258 VSUBS 0.016762f
C656 VTAIL.n259 VSUBS 0.02946f
C657 VTAIL.n260 VSUBS 0.015831f
C658 VTAIL.n261 VSUBS 0.037418f
C659 VTAIL.n262 VSUBS 0.016762f
C660 VTAIL.n263 VSUBS 0.02946f
C661 VTAIL.n264 VSUBS 0.015831f
C662 VTAIL.n265 VSUBS 0.037418f
C663 VTAIL.n266 VSUBS 0.016762f
C664 VTAIL.n267 VSUBS 0.02946f
C665 VTAIL.n268 VSUBS 0.015831f
C666 VTAIL.n269 VSUBS 0.037418f
C667 VTAIL.n270 VSUBS 0.016762f
C668 VTAIL.n271 VSUBS 0.02946f
C669 VTAIL.n272 VSUBS 0.015831f
C670 VTAIL.n273 VSUBS 0.037418f
C671 VTAIL.n274 VSUBS 0.016762f
C672 VTAIL.n275 VSUBS 0.02946f
C673 VTAIL.n276 VSUBS 0.015831f
C674 VTAIL.n277 VSUBS 0.037418f
C675 VTAIL.n278 VSUBS 0.016762f
C676 VTAIL.n279 VSUBS 0.206191f
C677 VTAIL.t2 VSUBS 0.080092f
C678 VTAIL.n280 VSUBS 0.028063f
C679 VTAIL.n281 VSUBS 0.023803f
C680 VTAIL.n282 VSUBS 0.015831f
C681 VTAIL.n283 VSUBS 1.85834f
C682 VTAIL.n284 VSUBS 0.02946f
C683 VTAIL.n285 VSUBS 0.015831f
C684 VTAIL.n286 VSUBS 0.016762f
C685 VTAIL.n287 VSUBS 0.037418f
C686 VTAIL.n288 VSUBS 0.037418f
C687 VTAIL.n289 VSUBS 0.016762f
C688 VTAIL.n290 VSUBS 0.015831f
C689 VTAIL.n291 VSUBS 0.02946f
C690 VTAIL.n292 VSUBS 0.02946f
C691 VTAIL.n293 VSUBS 0.015831f
C692 VTAIL.n294 VSUBS 0.016762f
C693 VTAIL.n295 VSUBS 0.037418f
C694 VTAIL.n296 VSUBS 0.037418f
C695 VTAIL.n297 VSUBS 0.016762f
C696 VTAIL.n298 VSUBS 0.015831f
C697 VTAIL.n299 VSUBS 0.02946f
C698 VTAIL.n300 VSUBS 0.02946f
C699 VTAIL.n301 VSUBS 0.015831f
C700 VTAIL.n302 VSUBS 0.016762f
C701 VTAIL.n303 VSUBS 0.037418f
C702 VTAIL.n304 VSUBS 0.037418f
C703 VTAIL.n305 VSUBS 0.016762f
C704 VTAIL.n306 VSUBS 0.015831f
C705 VTAIL.n307 VSUBS 0.02946f
C706 VTAIL.n308 VSUBS 0.02946f
C707 VTAIL.n309 VSUBS 0.015831f
C708 VTAIL.n310 VSUBS 0.016762f
C709 VTAIL.n311 VSUBS 0.037418f
C710 VTAIL.n312 VSUBS 0.037418f
C711 VTAIL.n313 VSUBS 0.016762f
C712 VTAIL.n314 VSUBS 0.015831f
C713 VTAIL.n315 VSUBS 0.02946f
C714 VTAIL.n316 VSUBS 0.02946f
C715 VTAIL.n317 VSUBS 0.015831f
C716 VTAIL.n318 VSUBS 0.016762f
C717 VTAIL.n319 VSUBS 0.037418f
C718 VTAIL.n320 VSUBS 0.037418f
C719 VTAIL.n321 VSUBS 0.037418f
C720 VTAIL.n322 VSUBS 0.016762f
C721 VTAIL.n323 VSUBS 0.015831f
C722 VTAIL.n324 VSUBS 0.02946f
C723 VTAIL.n325 VSUBS 0.02946f
C724 VTAIL.n326 VSUBS 0.015831f
C725 VTAIL.n327 VSUBS 0.016296f
C726 VTAIL.n328 VSUBS 0.016296f
C727 VTAIL.n329 VSUBS 0.037418f
C728 VTAIL.n330 VSUBS 0.089739f
C729 VTAIL.n331 VSUBS 0.016762f
C730 VTAIL.n332 VSUBS 0.015831f
C731 VTAIL.n333 VSUBS 0.075742f
C732 VTAIL.n334 VSUBS 0.045315f
C733 VTAIL.n335 VSUBS 1.76662f
C734 VP.n0 VSUBS 0.080283f
C735 VP.t4 VSUBS 1.47009f
C736 VP.n1 VSUBS 0.5441f
C737 VP.t1 VSUBS 1.44918f
C738 VP.t2 VSUBS 1.44918f
C739 VP.n2 VSUBS 0.577434f
C740 VP.n3 VSUBS 0.563749f
C741 VP.n4 VSUBS 2.771f
C742 VP.n5 VSUBS 2.64829f
C743 VP.t0 VSUBS 1.44918f
C744 VP.n6 VSUBS 0.563749f
C745 VP.t5 VSUBS 1.44918f
C746 VP.n7 VSUBS 0.577434f
C747 VP.t3 VSUBS 1.44918f
C748 VP.n8 VSUBS 0.563749f
C749 VP.n9 VSUBS 0.0669f
C750 B.n0 VSUBS 0.006343f
C751 B.n1 VSUBS 0.006343f
C752 B.n2 VSUBS 0.009381f
C753 B.n3 VSUBS 0.007189f
C754 B.n4 VSUBS 0.007189f
C755 B.n5 VSUBS 0.007189f
C756 B.n6 VSUBS 0.007189f
C757 B.n7 VSUBS 0.007189f
C758 B.n8 VSUBS 0.007189f
C759 B.n9 VSUBS 0.007189f
C760 B.n10 VSUBS 0.007189f
C761 B.n11 VSUBS 0.018628f
C762 B.n12 VSUBS 0.007189f
C763 B.n13 VSUBS 0.007189f
C764 B.n14 VSUBS 0.007189f
C765 B.n15 VSUBS 0.007189f
C766 B.n16 VSUBS 0.007189f
C767 B.n17 VSUBS 0.007189f
C768 B.n18 VSUBS 0.007189f
C769 B.n19 VSUBS 0.007189f
C770 B.n20 VSUBS 0.007189f
C771 B.n21 VSUBS 0.007189f
C772 B.n22 VSUBS 0.007189f
C773 B.n23 VSUBS 0.007189f
C774 B.n24 VSUBS 0.007189f
C775 B.n25 VSUBS 0.007189f
C776 B.n26 VSUBS 0.007189f
C777 B.n27 VSUBS 0.007189f
C778 B.n28 VSUBS 0.007189f
C779 B.n29 VSUBS 0.007189f
C780 B.n30 VSUBS 0.007189f
C781 B.n31 VSUBS 0.007189f
C782 B.n32 VSUBS 0.007189f
C783 B.n33 VSUBS 0.007189f
C784 B.n34 VSUBS 0.007189f
C785 B.n35 VSUBS 0.007189f
C786 B.t1 VSUBS 0.283147f
C787 B.t2 VSUBS 0.294089f
C788 B.t0 VSUBS 0.349228f
C789 B.n36 VSUBS 0.367429f
C790 B.n37 VSUBS 0.288647f
C791 B.n38 VSUBS 0.016656f
C792 B.n39 VSUBS 0.007189f
C793 B.n40 VSUBS 0.007189f
C794 B.n41 VSUBS 0.007189f
C795 B.n42 VSUBS 0.007189f
C796 B.n43 VSUBS 0.007189f
C797 B.t7 VSUBS 0.283151f
C798 B.t8 VSUBS 0.294092f
C799 B.t6 VSUBS 0.349228f
C800 B.n44 VSUBS 0.367426f
C801 B.n45 VSUBS 0.288644f
C802 B.n46 VSUBS 0.007189f
C803 B.n47 VSUBS 0.007189f
C804 B.n48 VSUBS 0.007189f
C805 B.n49 VSUBS 0.007189f
C806 B.n50 VSUBS 0.007189f
C807 B.n51 VSUBS 0.007189f
C808 B.n52 VSUBS 0.007189f
C809 B.n53 VSUBS 0.007189f
C810 B.n54 VSUBS 0.007189f
C811 B.n55 VSUBS 0.007189f
C812 B.n56 VSUBS 0.007189f
C813 B.n57 VSUBS 0.007189f
C814 B.n58 VSUBS 0.007189f
C815 B.n59 VSUBS 0.007189f
C816 B.n60 VSUBS 0.007189f
C817 B.n61 VSUBS 0.007189f
C818 B.n62 VSUBS 0.007189f
C819 B.n63 VSUBS 0.007189f
C820 B.n64 VSUBS 0.007189f
C821 B.n65 VSUBS 0.007189f
C822 B.n66 VSUBS 0.007189f
C823 B.n67 VSUBS 0.007189f
C824 B.n68 VSUBS 0.007189f
C825 B.n69 VSUBS 0.007189f
C826 B.n70 VSUBS 0.017951f
C827 B.n71 VSUBS 0.007189f
C828 B.n72 VSUBS 0.007189f
C829 B.n73 VSUBS 0.007189f
C830 B.n74 VSUBS 0.007189f
C831 B.n75 VSUBS 0.007189f
C832 B.n76 VSUBS 0.007189f
C833 B.n77 VSUBS 0.007189f
C834 B.n78 VSUBS 0.007189f
C835 B.n79 VSUBS 0.007189f
C836 B.n80 VSUBS 0.007189f
C837 B.n81 VSUBS 0.007189f
C838 B.n82 VSUBS 0.007189f
C839 B.n83 VSUBS 0.007189f
C840 B.n84 VSUBS 0.007189f
C841 B.n85 VSUBS 0.007189f
C842 B.n86 VSUBS 0.007189f
C843 B.n87 VSUBS 0.007189f
C844 B.n88 VSUBS 0.007189f
C845 B.n89 VSUBS 0.018628f
C846 B.n90 VSUBS 0.007189f
C847 B.n91 VSUBS 0.007189f
C848 B.n92 VSUBS 0.007189f
C849 B.n93 VSUBS 0.007189f
C850 B.n94 VSUBS 0.007189f
C851 B.n95 VSUBS 0.007189f
C852 B.n96 VSUBS 0.007189f
C853 B.n97 VSUBS 0.007189f
C854 B.n98 VSUBS 0.007189f
C855 B.n99 VSUBS 0.007189f
C856 B.n100 VSUBS 0.007189f
C857 B.n101 VSUBS 0.007189f
C858 B.n102 VSUBS 0.007189f
C859 B.n103 VSUBS 0.007189f
C860 B.n104 VSUBS 0.007189f
C861 B.n105 VSUBS 0.007189f
C862 B.n106 VSUBS 0.007189f
C863 B.n107 VSUBS 0.007189f
C864 B.n108 VSUBS 0.007189f
C865 B.n109 VSUBS 0.007189f
C866 B.n110 VSUBS 0.007189f
C867 B.n111 VSUBS 0.007189f
C868 B.n112 VSUBS 0.007189f
C869 B.n113 VSUBS 0.007189f
C870 B.t11 VSUBS 0.283151f
C871 B.t10 VSUBS 0.294092f
C872 B.t9 VSUBS 0.349228f
C873 B.n114 VSUBS 0.367426f
C874 B.n115 VSUBS 0.288644f
C875 B.n116 VSUBS 0.016656f
C876 B.n117 VSUBS 0.007189f
C877 B.n118 VSUBS 0.007189f
C878 B.n119 VSUBS 0.007189f
C879 B.n120 VSUBS 0.007189f
C880 B.n121 VSUBS 0.007189f
C881 B.t5 VSUBS 0.283147f
C882 B.t4 VSUBS 0.294089f
C883 B.t3 VSUBS 0.349228f
C884 B.n122 VSUBS 0.367429f
C885 B.n123 VSUBS 0.288647f
C886 B.n124 VSUBS 0.007189f
C887 B.n125 VSUBS 0.007189f
C888 B.n126 VSUBS 0.007189f
C889 B.n127 VSUBS 0.007189f
C890 B.n128 VSUBS 0.007189f
C891 B.n129 VSUBS 0.007189f
C892 B.n130 VSUBS 0.007189f
C893 B.n131 VSUBS 0.007189f
C894 B.n132 VSUBS 0.007189f
C895 B.n133 VSUBS 0.007189f
C896 B.n134 VSUBS 0.007189f
C897 B.n135 VSUBS 0.007189f
C898 B.n136 VSUBS 0.007189f
C899 B.n137 VSUBS 0.007189f
C900 B.n138 VSUBS 0.007189f
C901 B.n139 VSUBS 0.007189f
C902 B.n140 VSUBS 0.007189f
C903 B.n141 VSUBS 0.007189f
C904 B.n142 VSUBS 0.007189f
C905 B.n143 VSUBS 0.007189f
C906 B.n144 VSUBS 0.007189f
C907 B.n145 VSUBS 0.007189f
C908 B.n146 VSUBS 0.007189f
C909 B.n147 VSUBS 0.007189f
C910 B.n148 VSUBS 0.017951f
C911 B.n149 VSUBS 0.007189f
C912 B.n150 VSUBS 0.007189f
C913 B.n151 VSUBS 0.007189f
C914 B.n152 VSUBS 0.007189f
C915 B.n153 VSUBS 0.007189f
C916 B.n154 VSUBS 0.007189f
C917 B.n155 VSUBS 0.007189f
C918 B.n156 VSUBS 0.007189f
C919 B.n157 VSUBS 0.007189f
C920 B.n158 VSUBS 0.007189f
C921 B.n159 VSUBS 0.007189f
C922 B.n160 VSUBS 0.007189f
C923 B.n161 VSUBS 0.007189f
C924 B.n162 VSUBS 0.007189f
C925 B.n163 VSUBS 0.007189f
C926 B.n164 VSUBS 0.007189f
C927 B.n165 VSUBS 0.007189f
C928 B.n166 VSUBS 0.007189f
C929 B.n167 VSUBS 0.007189f
C930 B.n168 VSUBS 0.007189f
C931 B.n169 VSUBS 0.007189f
C932 B.n170 VSUBS 0.007189f
C933 B.n171 VSUBS 0.007189f
C934 B.n172 VSUBS 0.007189f
C935 B.n173 VSUBS 0.007189f
C936 B.n174 VSUBS 0.007189f
C937 B.n175 VSUBS 0.007189f
C938 B.n176 VSUBS 0.007189f
C939 B.n177 VSUBS 0.007189f
C940 B.n178 VSUBS 0.007189f
C941 B.n179 VSUBS 0.007189f
C942 B.n180 VSUBS 0.007189f
C943 B.n181 VSUBS 0.017951f
C944 B.n182 VSUBS 0.018628f
C945 B.n183 VSUBS 0.018628f
C946 B.n184 VSUBS 0.007189f
C947 B.n185 VSUBS 0.007189f
C948 B.n186 VSUBS 0.007189f
C949 B.n187 VSUBS 0.007189f
C950 B.n188 VSUBS 0.007189f
C951 B.n189 VSUBS 0.007189f
C952 B.n190 VSUBS 0.007189f
C953 B.n191 VSUBS 0.007189f
C954 B.n192 VSUBS 0.007189f
C955 B.n193 VSUBS 0.007189f
C956 B.n194 VSUBS 0.007189f
C957 B.n195 VSUBS 0.007189f
C958 B.n196 VSUBS 0.007189f
C959 B.n197 VSUBS 0.007189f
C960 B.n198 VSUBS 0.007189f
C961 B.n199 VSUBS 0.007189f
C962 B.n200 VSUBS 0.007189f
C963 B.n201 VSUBS 0.007189f
C964 B.n202 VSUBS 0.007189f
C965 B.n203 VSUBS 0.007189f
C966 B.n204 VSUBS 0.007189f
C967 B.n205 VSUBS 0.007189f
C968 B.n206 VSUBS 0.007189f
C969 B.n207 VSUBS 0.007189f
C970 B.n208 VSUBS 0.007189f
C971 B.n209 VSUBS 0.007189f
C972 B.n210 VSUBS 0.007189f
C973 B.n211 VSUBS 0.007189f
C974 B.n212 VSUBS 0.007189f
C975 B.n213 VSUBS 0.007189f
C976 B.n214 VSUBS 0.007189f
C977 B.n215 VSUBS 0.007189f
C978 B.n216 VSUBS 0.007189f
C979 B.n217 VSUBS 0.007189f
C980 B.n218 VSUBS 0.007189f
C981 B.n219 VSUBS 0.007189f
C982 B.n220 VSUBS 0.007189f
C983 B.n221 VSUBS 0.007189f
C984 B.n222 VSUBS 0.007189f
C985 B.n223 VSUBS 0.007189f
C986 B.n224 VSUBS 0.007189f
C987 B.n225 VSUBS 0.007189f
C988 B.n226 VSUBS 0.007189f
C989 B.n227 VSUBS 0.007189f
C990 B.n228 VSUBS 0.007189f
C991 B.n229 VSUBS 0.007189f
C992 B.n230 VSUBS 0.007189f
C993 B.n231 VSUBS 0.007189f
C994 B.n232 VSUBS 0.007189f
C995 B.n233 VSUBS 0.007189f
C996 B.n234 VSUBS 0.007189f
C997 B.n235 VSUBS 0.007189f
C998 B.n236 VSUBS 0.007189f
C999 B.n237 VSUBS 0.007189f
C1000 B.n238 VSUBS 0.007189f
C1001 B.n239 VSUBS 0.007189f
C1002 B.n240 VSUBS 0.007189f
C1003 B.n241 VSUBS 0.007189f
C1004 B.n242 VSUBS 0.007189f
C1005 B.n243 VSUBS 0.007189f
C1006 B.n244 VSUBS 0.007189f
C1007 B.n245 VSUBS 0.007189f
C1008 B.n246 VSUBS 0.007189f
C1009 B.n247 VSUBS 0.007189f
C1010 B.n248 VSUBS 0.007189f
C1011 B.n249 VSUBS 0.007189f
C1012 B.n250 VSUBS 0.007189f
C1013 B.n251 VSUBS 0.007189f
C1014 B.n252 VSUBS 0.007189f
C1015 B.n253 VSUBS 0.007189f
C1016 B.n254 VSUBS 0.007189f
C1017 B.n255 VSUBS 0.007189f
C1018 B.n256 VSUBS 0.004969f
C1019 B.n257 VSUBS 0.016656f
C1020 B.n258 VSUBS 0.005815f
C1021 B.n259 VSUBS 0.007189f
C1022 B.n260 VSUBS 0.007189f
C1023 B.n261 VSUBS 0.007189f
C1024 B.n262 VSUBS 0.007189f
C1025 B.n263 VSUBS 0.007189f
C1026 B.n264 VSUBS 0.007189f
C1027 B.n265 VSUBS 0.007189f
C1028 B.n266 VSUBS 0.007189f
C1029 B.n267 VSUBS 0.007189f
C1030 B.n268 VSUBS 0.007189f
C1031 B.n269 VSUBS 0.007189f
C1032 B.n270 VSUBS 0.005815f
C1033 B.n271 VSUBS 0.007189f
C1034 B.n272 VSUBS 0.007189f
C1035 B.n273 VSUBS 0.004969f
C1036 B.n274 VSUBS 0.007189f
C1037 B.n275 VSUBS 0.007189f
C1038 B.n276 VSUBS 0.007189f
C1039 B.n277 VSUBS 0.007189f
C1040 B.n278 VSUBS 0.007189f
C1041 B.n279 VSUBS 0.007189f
C1042 B.n280 VSUBS 0.007189f
C1043 B.n281 VSUBS 0.007189f
C1044 B.n282 VSUBS 0.007189f
C1045 B.n283 VSUBS 0.007189f
C1046 B.n284 VSUBS 0.007189f
C1047 B.n285 VSUBS 0.007189f
C1048 B.n286 VSUBS 0.007189f
C1049 B.n287 VSUBS 0.007189f
C1050 B.n288 VSUBS 0.007189f
C1051 B.n289 VSUBS 0.007189f
C1052 B.n290 VSUBS 0.007189f
C1053 B.n291 VSUBS 0.007189f
C1054 B.n292 VSUBS 0.007189f
C1055 B.n293 VSUBS 0.007189f
C1056 B.n294 VSUBS 0.007189f
C1057 B.n295 VSUBS 0.007189f
C1058 B.n296 VSUBS 0.007189f
C1059 B.n297 VSUBS 0.007189f
C1060 B.n298 VSUBS 0.007189f
C1061 B.n299 VSUBS 0.007189f
C1062 B.n300 VSUBS 0.007189f
C1063 B.n301 VSUBS 0.007189f
C1064 B.n302 VSUBS 0.007189f
C1065 B.n303 VSUBS 0.007189f
C1066 B.n304 VSUBS 0.007189f
C1067 B.n305 VSUBS 0.007189f
C1068 B.n306 VSUBS 0.007189f
C1069 B.n307 VSUBS 0.007189f
C1070 B.n308 VSUBS 0.007189f
C1071 B.n309 VSUBS 0.007189f
C1072 B.n310 VSUBS 0.007189f
C1073 B.n311 VSUBS 0.007189f
C1074 B.n312 VSUBS 0.007189f
C1075 B.n313 VSUBS 0.007189f
C1076 B.n314 VSUBS 0.007189f
C1077 B.n315 VSUBS 0.007189f
C1078 B.n316 VSUBS 0.007189f
C1079 B.n317 VSUBS 0.007189f
C1080 B.n318 VSUBS 0.007189f
C1081 B.n319 VSUBS 0.007189f
C1082 B.n320 VSUBS 0.007189f
C1083 B.n321 VSUBS 0.007189f
C1084 B.n322 VSUBS 0.007189f
C1085 B.n323 VSUBS 0.007189f
C1086 B.n324 VSUBS 0.007189f
C1087 B.n325 VSUBS 0.007189f
C1088 B.n326 VSUBS 0.007189f
C1089 B.n327 VSUBS 0.007189f
C1090 B.n328 VSUBS 0.007189f
C1091 B.n329 VSUBS 0.007189f
C1092 B.n330 VSUBS 0.007189f
C1093 B.n331 VSUBS 0.007189f
C1094 B.n332 VSUBS 0.007189f
C1095 B.n333 VSUBS 0.007189f
C1096 B.n334 VSUBS 0.007189f
C1097 B.n335 VSUBS 0.007189f
C1098 B.n336 VSUBS 0.007189f
C1099 B.n337 VSUBS 0.007189f
C1100 B.n338 VSUBS 0.007189f
C1101 B.n339 VSUBS 0.007189f
C1102 B.n340 VSUBS 0.007189f
C1103 B.n341 VSUBS 0.007189f
C1104 B.n342 VSUBS 0.007189f
C1105 B.n343 VSUBS 0.007189f
C1106 B.n344 VSUBS 0.007189f
C1107 B.n345 VSUBS 0.007189f
C1108 B.n346 VSUBS 0.017878f
C1109 B.n347 VSUBS 0.018701f
C1110 B.n348 VSUBS 0.017951f
C1111 B.n349 VSUBS 0.007189f
C1112 B.n350 VSUBS 0.007189f
C1113 B.n351 VSUBS 0.007189f
C1114 B.n352 VSUBS 0.007189f
C1115 B.n353 VSUBS 0.007189f
C1116 B.n354 VSUBS 0.007189f
C1117 B.n355 VSUBS 0.007189f
C1118 B.n356 VSUBS 0.007189f
C1119 B.n357 VSUBS 0.007189f
C1120 B.n358 VSUBS 0.007189f
C1121 B.n359 VSUBS 0.007189f
C1122 B.n360 VSUBS 0.007189f
C1123 B.n361 VSUBS 0.007189f
C1124 B.n362 VSUBS 0.007189f
C1125 B.n363 VSUBS 0.007189f
C1126 B.n364 VSUBS 0.007189f
C1127 B.n365 VSUBS 0.007189f
C1128 B.n366 VSUBS 0.007189f
C1129 B.n367 VSUBS 0.007189f
C1130 B.n368 VSUBS 0.007189f
C1131 B.n369 VSUBS 0.007189f
C1132 B.n370 VSUBS 0.007189f
C1133 B.n371 VSUBS 0.007189f
C1134 B.n372 VSUBS 0.007189f
C1135 B.n373 VSUBS 0.007189f
C1136 B.n374 VSUBS 0.007189f
C1137 B.n375 VSUBS 0.007189f
C1138 B.n376 VSUBS 0.007189f
C1139 B.n377 VSUBS 0.007189f
C1140 B.n378 VSUBS 0.007189f
C1141 B.n379 VSUBS 0.007189f
C1142 B.n380 VSUBS 0.007189f
C1143 B.n381 VSUBS 0.007189f
C1144 B.n382 VSUBS 0.007189f
C1145 B.n383 VSUBS 0.007189f
C1146 B.n384 VSUBS 0.007189f
C1147 B.n385 VSUBS 0.007189f
C1148 B.n386 VSUBS 0.007189f
C1149 B.n387 VSUBS 0.007189f
C1150 B.n388 VSUBS 0.007189f
C1151 B.n389 VSUBS 0.007189f
C1152 B.n390 VSUBS 0.007189f
C1153 B.n391 VSUBS 0.007189f
C1154 B.n392 VSUBS 0.007189f
C1155 B.n393 VSUBS 0.007189f
C1156 B.n394 VSUBS 0.007189f
C1157 B.n395 VSUBS 0.007189f
C1158 B.n396 VSUBS 0.007189f
C1159 B.n397 VSUBS 0.007189f
C1160 B.n398 VSUBS 0.007189f
C1161 B.n399 VSUBS 0.007189f
C1162 B.n400 VSUBS 0.007189f
C1163 B.n401 VSUBS 0.007189f
C1164 B.n402 VSUBS 0.007189f
C1165 B.n403 VSUBS 0.017951f
C1166 B.n404 VSUBS 0.018628f
C1167 B.n405 VSUBS 0.018628f
C1168 B.n406 VSUBS 0.007189f
C1169 B.n407 VSUBS 0.007189f
C1170 B.n408 VSUBS 0.007189f
C1171 B.n409 VSUBS 0.007189f
C1172 B.n410 VSUBS 0.007189f
C1173 B.n411 VSUBS 0.007189f
C1174 B.n412 VSUBS 0.007189f
C1175 B.n413 VSUBS 0.007189f
C1176 B.n414 VSUBS 0.007189f
C1177 B.n415 VSUBS 0.007189f
C1178 B.n416 VSUBS 0.007189f
C1179 B.n417 VSUBS 0.007189f
C1180 B.n418 VSUBS 0.007189f
C1181 B.n419 VSUBS 0.007189f
C1182 B.n420 VSUBS 0.007189f
C1183 B.n421 VSUBS 0.007189f
C1184 B.n422 VSUBS 0.007189f
C1185 B.n423 VSUBS 0.007189f
C1186 B.n424 VSUBS 0.007189f
C1187 B.n425 VSUBS 0.007189f
C1188 B.n426 VSUBS 0.007189f
C1189 B.n427 VSUBS 0.007189f
C1190 B.n428 VSUBS 0.007189f
C1191 B.n429 VSUBS 0.007189f
C1192 B.n430 VSUBS 0.007189f
C1193 B.n431 VSUBS 0.007189f
C1194 B.n432 VSUBS 0.007189f
C1195 B.n433 VSUBS 0.007189f
C1196 B.n434 VSUBS 0.007189f
C1197 B.n435 VSUBS 0.007189f
C1198 B.n436 VSUBS 0.007189f
C1199 B.n437 VSUBS 0.007189f
C1200 B.n438 VSUBS 0.007189f
C1201 B.n439 VSUBS 0.007189f
C1202 B.n440 VSUBS 0.007189f
C1203 B.n441 VSUBS 0.007189f
C1204 B.n442 VSUBS 0.007189f
C1205 B.n443 VSUBS 0.007189f
C1206 B.n444 VSUBS 0.007189f
C1207 B.n445 VSUBS 0.007189f
C1208 B.n446 VSUBS 0.007189f
C1209 B.n447 VSUBS 0.007189f
C1210 B.n448 VSUBS 0.007189f
C1211 B.n449 VSUBS 0.007189f
C1212 B.n450 VSUBS 0.007189f
C1213 B.n451 VSUBS 0.007189f
C1214 B.n452 VSUBS 0.007189f
C1215 B.n453 VSUBS 0.007189f
C1216 B.n454 VSUBS 0.007189f
C1217 B.n455 VSUBS 0.007189f
C1218 B.n456 VSUBS 0.007189f
C1219 B.n457 VSUBS 0.007189f
C1220 B.n458 VSUBS 0.007189f
C1221 B.n459 VSUBS 0.007189f
C1222 B.n460 VSUBS 0.007189f
C1223 B.n461 VSUBS 0.007189f
C1224 B.n462 VSUBS 0.007189f
C1225 B.n463 VSUBS 0.007189f
C1226 B.n464 VSUBS 0.007189f
C1227 B.n465 VSUBS 0.007189f
C1228 B.n466 VSUBS 0.007189f
C1229 B.n467 VSUBS 0.007189f
C1230 B.n468 VSUBS 0.007189f
C1231 B.n469 VSUBS 0.007189f
C1232 B.n470 VSUBS 0.007189f
C1233 B.n471 VSUBS 0.007189f
C1234 B.n472 VSUBS 0.007189f
C1235 B.n473 VSUBS 0.007189f
C1236 B.n474 VSUBS 0.007189f
C1237 B.n475 VSUBS 0.007189f
C1238 B.n476 VSUBS 0.007189f
C1239 B.n477 VSUBS 0.007189f
C1240 B.n478 VSUBS 0.004969f
C1241 B.n479 VSUBS 0.016656f
C1242 B.n480 VSUBS 0.005815f
C1243 B.n481 VSUBS 0.007189f
C1244 B.n482 VSUBS 0.007189f
C1245 B.n483 VSUBS 0.007189f
C1246 B.n484 VSUBS 0.007189f
C1247 B.n485 VSUBS 0.007189f
C1248 B.n486 VSUBS 0.007189f
C1249 B.n487 VSUBS 0.007189f
C1250 B.n488 VSUBS 0.007189f
C1251 B.n489 VSUBS 0.007189f
C1252 B.n490 VSUBS 0.007189f
C1253 B.n491 VSUBS 0.007189f
C1254 B.n492 VSUBS 0.005815f
C1255 B.n493 VSUBS 0.007189f
C1256 B.n494 VSUBS 0.007189f
C1257 B.n495 VSUBS 0.004969f
C1258 B.n496 VSUBS 0.007189f
C1259 B.n497 VSUBS 0.007189f
C1260 B.n498 VSUBS 0.007189f
C1261 B.n499 VSUBS 0.007189f
C1262 B.n500 VSUBS 0.007189f
C1263 B.n501 VSUBS 0.007189f
C1264 B.n502 VSUBS 0.007189f
C1265 B.n503 VSUBS 0.007189f
C1266 B.n504 VSUBS 0.007189f
C1267 B.n505 VSUBS 0.007189f
C1268 B.n506 VSUBS 0.007189f
C1269 B.n507 VSUBS 0.007189f
C1270 B.n508 VSUBS 0.007189f
C1271 B.n509 VSUBS 0.007189f
C1272 B.n510 VSUBS 0.007189f
C1273 B.n511 VSUBS 0.007189f
C1274 B.n512 VSUBS 0.007189f
C1275 B.n513 VSUBS 0.007189f
C1276 B.n514 VSUBS 0.007189f
C1277 B.n515 VSUBS 0.007189f
C1278 B.n516 VSUBS 0.007189f
C1279 B.n517 VSUBS 0.007189f
C1280 B.n518 VSUBS 0.007189f
C1281 B.n519 VSUBS 0.007189f
C1282 B.n520 VSUBS 0.007189f
C1283 B.n521 VSUBS 0.007189f
C1284 B.n522 VSUBS 0.007189f
C1285 B.n523 VSUBS 0.007189f
C1286 B.n524 VSUBS 0.007189f
C1287 B.n525 VSUBS 0.007189f
C1288 B.n526 VSUBS 0.007189f
C1289 B.n527 VSUBS 0.007189f
C1290 B.n528 VSUBS 0.007189f
C1291 B.n529 VSUBS 0.007189f
C1292 B.n530 VSUBS 0.007189f
C1293 B.n531 VSUBS 0.007189f
C1294 B.n532 VSUBS 0.007189f
C1295 B.n533 VSUBS 0.007189f
C1296 B.n534 VSUBS 0.007189f
C1297 B.n535 VSUBS 0.007189f
C1298 B.n536 VSUBS 0.007189f
C1299 B.n537 VSUBS 0.007189f
C1300 B.n538 VSUBS 0.007189f
C1301 B.n539 VSUBS 0.007189f
C1302 B.n540 VSUBS 0.007189f
C1303 B.n541 VSUBS 0.007189f
C1304 B.n542 VSUBS 0.007189f
C1305 B.n543 VSUBS 0.007189f
C1306 B.n544 VSUBS 0.007189f
C1307 B.n545 VSUBS 0.007189f
C1308 B.n546 VSUBS 0.007189f
C1309 B.n547 VSUBS 0.007189f
C1310 B.n548 VSUBS 0.007189f
C1311 B.n549 VSUBS 0.007189f
C1312 B.n550 VSUBS 0.007189f
C1313 B.n551 VSUBS 0.007189f
C1314 B.n552 VSUBS 0.007189f
C1315 B.n553 VSUBS 0.007189f
C1316 B.n554 VSUBS 0.007189f
C1317 B.n555 VSUBS 0.007189f
C1318 B.n556 VSUBS 0.007189f
C1319 B.n557 VSUBS 0.007189f
C1320 B.n558 VSUBS 0.007189f
C1321 B.n559 VSUBS 0.007189f
C1322 B.n560 VSUBS 0.007189f
C1323 B.n561 VSUBS 0.007189f
C1324 B.n562 VSUBS 0.007189f
C1325 B.n563 VSUBS 0.007189f
C1326 B.n564 VSUBS 0.007189f
C1327 B.n565 VSUBS 0.007189f
C1328 B.n566 VSUBS 0.007189f
C1329 B.n567 VSUBS 0.007189f
C1330 B.n568 VSUBS 0.018628f
C1331 B.n569 VSUBS 0.017951f
C1332 B.n570 VSUBS 0.017951f
C1333 B.n571 VSUBS 0.007189f
C1334 B.n572 VSUBS 0.007189f
C1335 B.n573 VSUBS 0.007189f
C1336 B.n574 VSUBS 0.007189f
C1337 B.n575 VSUBS 0.007189f
C1338 B.n576 VSUBS 0.007189f
C1339 B.n577 VSUBS 0.007189f
C1340 B.n578 VSUBS 0.007189f
C1341 B.n579 VSUBS 0.007189f
C1342 B.n580 VSUBS 0.007189f
C1343 B.n581 VSUBS 0.007189f
C1344 B.n582 VSUBS 0.007189f
C1345 B.n583 VSUBS 0.007189f
C1346 B.n584 VSUBS 0.007189f
C1347 B.n585 VSUBS 0.007189f
C1348 B.n586 VSUBS 0.007189f
C1349 B.n587 VSUBS 0.007189f
C1350 B.n588 VSUBS 0.007189f
C1351 B.n589 VSUBS 0.007189f
C1352 B.n590 VSUBS 0.007189f
C1353 B.n591 VSUBS 0.007189f
C1354 B.n592 VSUBS 0.007189f
C1355 B.n593 VSUBS 0.007189f
C1356 B.n594 VSUBS 0.007189f
C1357 B.n595 VSUBS 0.009381f
C1358 B.n596 VSUBS 0.009993f
C1359 B.n597 VSUBS 0.019873f
.ends

