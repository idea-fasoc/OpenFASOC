* NGSPICE file created from tg_sample_0005.ext - technology: sky130A

.subckt tg_sample_0005 VIN VGN VGP VSS VCC VOUT
X0 VSS.t17 VSS.t15 VSS.t16 VSS.t9 sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.28
X1 VCC.t17 VCC.t15 VCC.t16 VCC.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.28
X2 VOUT.t35 VOUT.t34 VOUT.t35 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=0 ps=0 w=8 l=0.28
X3 VOUT.t33 VOUT.t32 VOUT.t33 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=0 ps=0 w=8 l=0.28
X4 VOUT.t31 VOUT.t29 VOUT.t30 VCC.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.28
X5 VOUT.t28 VOUT.t27 VOUT.t28 VCC.t3 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=0 ps=0 w=8 l=0.28
X6 VOUT.t26 VOUT.t24 VOUT.t25 VSS.t1 sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.28
X7 VOUT.t23 VOUT.t22 VOUT.t23 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=0 ps=0 w=8 l=0.28
X8 VOUT.t21 VOUT.t20 VOUT.t21 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=0 ps=0 w=8 l=0.28
X9 VOUT.t19 VOUT.t17 VOUT.t18 VSS.t1 sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.28
X10 VOUT.t16 VOUT.t15 VOUT.t16 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0 ps=0 w=4 l=0.28
X11 VOUT.t14 VOUT.t13 VOUT.t14 VCC.t3 sky130_fd_pr__pfet_01v8 ad=1.32 pd=8.33 as=0 ps=0 w=8 l=0.28
X12 VSS.t14 VSS.t12 VSS.t13 VSS.t5 sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.28
X13 VSS.t11 VSS.t8 VSS.t10 VSS.t9 sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.28
X14 VOUT.t12 VOUT.t11 VOUT.t12 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0 ps=0 w=4 l=0.28
X15 VOUT.t10 VOUT.t9 VOUT.t10 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0 ps=0 w=4 l=0.28
X16 VSS.t7 VSS.t4 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=1.56 pd=8.78 as=0 ps=0 w=4 l=0.28
X17 VOUT.t8 VOUT.t7 VOUT.t8 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0 ps=0 w=4 l=0.28
X18 VOUT.t6 VOUT.t5 VOUT.t6 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0 ps=0 w=4 l=0.28
X19 VCC.t14 VCC.t12 VCC.t13 VCC.t5 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.28
X20 VCC.t11 VCC.t8 VCC.t10 VCC.t9 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.28
X21 VOUT.t4 VOUT.t3 VOUT.t4 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.66 pd=4.33 as=0 ps=0 w=4 l=0.28
X22 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.28
X23 VOUT.t2 VOUT.t0 VOUT.t1 VCC.t2 sky130_fd_pr__pfet_01v8 ad=3.12 pd=16.78 as=0 ps=0 w=8 l=0.28
R0 VSS.n764 VSS.n150 4974.43
R1 VSS.n812 VSS.n811 4974.43
R2 VSS.n771 VSS.n150 2972.97
R3 VSS.n772 VSS.n771 2972.97
R4 VSS.n773 VSS.n772 2972.97
R5 VSS.n773 VSS.n144 2972.97
R6 VSS.n781 VSS.n144 2972.97
R7 VSS.n782 VSS.n781 2972.97
R8 VSS.n783 VSS.n782 2972.97
R9 VSS.n783 VSS.n138 2972.97
R10 VSS.n791 VSS.n138 2972.97
R11 VSS.n792 VSS.n791 2972.97
R12 VSS.n793 VSS.n792 2972.97
R13 VSS.n793 VSS.n132 2972.97
R14 VSS.n801 VSS.n132 2972.97
R15 VSS.n802 VSS.n801 2972.97
R16 VSS.n803 VSS.n802 2972.97
R17 VSS.n803 VSS.n126 2972.97
R18 VSS.n811 VSS.n126 2972.97
R19 VSS.n764 VSS.n763 1719.54
R20 VSS.n763 VSS.n762 1719.54
R21 VSS.n762 VSS.n155 1719.54
R22 VSS.n756 VSS.n155 1719.54
R23 VSS.n756 VSS.n755 1719.54
R24 VSS.n755 VSS.n754 1719.54
R25 VSS.n754 VSS.n159 1719.54
R26 VSS.n748 VSS.n159 1719.54
R27 VSS.n748 VSS.n747 1719.54
R28 VSS.n747 VSS.n746 1719.54
R29 VSS.n746 VSS.n163 1719.54
R30 VSS.n740 VSS.n163 1719.54
R31 VSS.n740 VSS.n739 1719.54
R32 VSS.n739 VSS.n738 1719.54
R33 VSS.n738 VSS.n167 1719.54
R34 VSS.n732 VSS.n167 1719.54
R35 VSS.n732 VSS.n731 1719.54
R36 VSS.n731 VSS.n730 1719.54
R37 VSS.n730 VSS.n171 1719.54
R38 VSS.n724 VSS.n171 1719.54
R39 VSS.n724 VSS.n723 1719.54
R40 VSS.n723 VSS.n722 1719.54
R41 VSS.n722 VSS.n175 1719.54
R42 VSS.n716 VSS.n175 1719.54
R43 VSS.n716 VSS.n715 1719.54
R44 VSS.n715 VSS.n714 1719.54
R45 VSS.n714 VSS.n179 1719.54
R46 VSS.n708 VSS.n179 1719.54
R47 VSS.n708 VSS.n707 1719.54
R48 VSS.n707 VSS.n706 1719.54
R49 VSS.n706 VSS.n183 1719.54
R50 VSS.n700 VSS.n183 1719.54
R51 VSS.n700 VSS.n699 1719.54
R52 VSS.n699 VSS.n698 1719.54
R53 VSS.n698 VSS.n187 1719.54
R54 VSS.n692 VSS.n187 1719.54
R55 VSS.n692 VSS.n691 1719.54
R56 VSS.n691 VSS.n690 1719.54
R57 VSS.n690 VSS.n191 1719.54
R58 VSS.n684 VSS.n191 1719.54
R59 VSS.n684 VSS.n683 1719.54
R60 VSS.n683 VSS.n682 1719.54
R61 VSS.n682 VSS.n195 1719.54
R62 VSS.n676 VSS.n195 1719.54
R63 VSS.n676 VSS.n675 1719.54
R64 VSS.n675 VSS.n674 1719.54
R65 VSS.n674 VSS.n199 1719.54
R66 VSS.n668 VSS.n199 1719.54
R67 VSS.n668 VSS.n667 1719.54
R68 VSS.n667 VSS.n666 1719.54
R69 VSS.n666 VSS.n203 1719.54
R70 VSS.n660 VSS.n203 1719.54
R71 VSS.n660 VSS.n659 1719.54
R72 VSS.n659 VSS.n658 1719.54
R73 VSS.n658 VSS.n207 1719.54
R74 VSS.n652 VSS.n207 1719.54
R75 VSS.n652 VSS.n651 1719.54
R76 VSS.n651 VSS.n650 1719.54
R77 VSS.n650 VSS.n211 1719.54
R78 VSS.n644 VSS.n211 1719.54
R79 VSS.n644 VSS.n643 1719.54
R80 VSS.n643 VSS.n642 1719.54
R81 VSS.n642 VSS.n215 1719.54
R82 VSS.n636 VSS.n215 1719.54
R83 VSS.n636 VSS.n635 1719.54
R84 VSS.n813 VSS.n812 1719.54
R85 VSS.n813 VSS.n122 1719.54
R86 VSS.n819 VSS.n122 1719.54
R87 VSS.n820 VSS.n819 1719.54
R88 VSS.n821 VSS.n820 1719.54
R89 VSS.n821 VSS.n118 1719.54
R90 VSS.n827 VSS.n118 1719.54
R91 VSS.n828 VSS.n827 1719.54
R92 VSS.n829 VSS.n828 1719.54
R93 VSS.n829 VSS.n114 1719.54
R94 VSS.n835 VSS.n114 1719.54
R95 VSS.n836 VSS.n835 1719.54
R96 VSS.n837 VSS.n836 1719.54
R97 VSS.n837 VSS.n110 1719.54
R98 VSS.n843 VSS.n110 1719.54
R99 VSS.n844 VSS.n843 1719.54
R100 VSS.n845 VSS.n844 1719.54
R101 VSS.n845 VSS.n106 1719.54
R102 VSS.n851 VSS.n106 1719.54
R103 VSS.n852 VSS.n851 1719.54
R104 VSS.n853 VSS.n852 1719.54
R105 VSS.n853 VSS.n102 1719.54
R106 VSS.n859 VSS.n102 1719.54
R107 VSS.n860 VSS.n859 1719.54
R108 VSS.n861 VSS.n860 1719.54
R109 VSS.n861 VSS.n98 1719.54
R110 VSS.n867 VSS.n98 1719.54
R111 VSS.n868 VSS.n867 1719.54
R112 VSS.n869 VSS.n868 1719.54
R113 VSS.n869 VSS.n94 1719.54
R114 VSS.n875 VSS.n94 1719.54
R115 VSS.n876 VSS.n875 1719.54
R116 VSS.n877 VSS.n876 1719.54
R117 VSS.n877 VSS.n90 1719.54
R118 VSS.n883 VSS.n90 1719.54
R119 VSS.n884 VSS.n883 1719.54
R120 VSS.n885 VSS.n884 1719.54
R121 VSS.n885 VSS.n86 1719.54
R122 VSS.n891 VSS.n86 1719.54
R123 VSS.n892 VSS.n891 1719.54
R124 VSS.n893 VSS.n892 1719.54
R125 VSS.n893 VSS.n82 1719.54
R126 VSS.n899 VSS.n82 1719.54
R127 VSS.n900 VSS.n899 1719.54
R128 VSS.n901 VSS.n900 1719.54
R129 VSS.n901 VSS.n78 1719.54
R130 VSS.n907 VSS.n78 1719.54
R131 VSS.n908 VSS.n907 1719.54
R132 VSS.n909 VSS.n908 1719.54
R133 VSS.n909 VSS.n74 1719.54
R134 VSS.n915 VSS.n74 1719.54
R135 VSS.n916 VSS.n915 1719.54
R136 VSS.n917 VSS.n916 1719.54
R137 VSS.n917 VSS.n70 1719.54
R138 VSS.n923 VSS.n70 1719.54
R139 VSS.n924 VSS.n923 1719.54
R140 VSS.n925 VSS.n924 1719.54
R141 VSS.n925 VSS.n66 1719.54
R142 VSS.n931 VSS.n66 1719.54
R143 VSS.n932 VSS.n931 1719.54
R144 VSS.n933 VSS.n932 1719.54
R145 VSS.n933 VSS.n62 1719.54
R146 VSS.n940 VSS.n62 1719.54
R147 VSS.n941 VSS.n940 1719.54
R148 VSS.n942 VSS.n941 1719.54
R149 VSS.n765 VSS.n151 622.232
R150 VSS.n810 VSS.n125 622.232
R151 VSS.n1033 VSS.n34 622.232
R152 VSS.n632 VSS.n221 622.232
R153 VSS.n480 VSS.n339 610.22
R154 VSS.n557 VSS.n554 610.22
R155 VSS.n603 VSS.n435 610.22
R156 VSS.n1037 VSS.n10 610.22
R157 VSS.n766 VSS.n765 585
R158 VSS.n765 VSS.n764 585
R159 VSS.n154 VSS.n153 585
R160 VSS.n763 VSS.n154 585
R161 VSS.n761 VSS.n760 585
R162 VSS.n762 VSS.n761 585
R163 VSS.n759 VSS.n156 585
R164 VSS.n156 VSS.n155 585
R165 VSS.n758 VSS.n757 585
R166 VSS.n757 VSS.n756 585
R167 VSS.n158 VSS.n157 585
R168 VSS.n755 VSS.n158 585
R169 VSS.n753 VSS.n752 585
R170 VSS.n754 VSS.n753 585
R171 VSS.n751 VSS.n160 585
R172 VSS.n160 VSS.n159 585
R173 VSS.n750 VSS.n749 585
R174 VSS.n749 VSS.n748 585
R175 VSS.n162 VSS.n161 585
R176 VSS.n747 VSS.n162 585
R177 VSS.n745 VSS.n744 585
R178 VSS.n746 VSS.n745 585
R179 VSS.n743 VSS.n164 585
R180 VSS.n164 VSS.n163 585
R181 VSS.n742 VSS.n741 585
R182 VSS.n741 VSS.n740 585
R183 VSS.n166 VSS.n165 585
R184 VSS.n739 VSS.n166 585
R185 VSS.n737 VSS.n736 585
R186 VSS.n738 VSS.n737 585
R187 VSS.n735 VSS.n168 585
R188 VSS.n168 VSS.n167 585
R189 VSS.n734 VSS.n733 585
R190 VSS.n733 VSS.n732 585
R191 VSS.n170 VSS.n169 585
R192 VSS.n731 VSS.n170 585
R193 VSS.n729 VSS.n728 585
R194 VSS.n730 VSS.n729 585
R195 VSS.n727 VSS.n172 585
R196 VSS.n172 VSS.n171 585
R197 VSS.n726 VSS.n725 585
R198 VSS.n725 VSS.n724 585
R199 VSS.n174 VSS.n173 585
R200 VSS.n723 VSS.n174 585
R201 VSS.n721 VSS.n720 585
R202 VSS.n722 VSS.n721 585
R203 VSS.n719 VSS.n176 585
R204 VSS.n176 VSS.n175 585
R205 VSS.n718 VSS.n717 585
R206 VSS.n717 VSS.n716 585
R207 VSS.n178 VSS.n177 585
R208 VSS.n715 VSS.n178 585
R209 VSS.n713 VSS.n712 585
R210 VSS.n714 VSS.n713 585
R211 VSS.n711 VSS.n180 585
R212 VSS.n180 VSS.n179 585
R213 VSS.n710 VSS.n709 585
R214 VSS.n709 VSS.n708 585
R215 VSS.n182 VSS.n181 585
R216 VSS.n707 VSS.n182 585
R217 VSS.n705 VSS.n704 585
R218 VSS.n706 VSS.n705 585
R219 VSS.n703 VSS.n184 585
R220 VSS.n184 VSS.n183 585
R221 VSS.n702 VSS.n701 585
R222 VSS.n701 VSS.n700 585
R223 VSS.n186 VSS.n185 585
R224 VSS.n699 VSS.n186 585
R225 VSS.n697 VSS.n696 585
R226 VSS.n698 VSS.n697 585
R227 VSS.n695 VSS.n188 585
R228 VSS.n188 VSS.n187 585
R229 VSS.n694 VSS.n693 585
R230 VSS.n693 VSS.n692 585
R231 VSS.n190 VSS.n189 585
R232 VSS.n691 VSS.n190 585
R233 VSS.n689 VSS.n688 585
R234 VSS.n690 VSS.n689 585
R235 VSS.n687 VSS.n192 585
R236 VSS.n192 VSS.n191 585
R237 VSS.n686 VSS.n685 585
R238 VSS.n685 VSS.n684 585
R239 VSS.n194 VSS.n193 585
R240 VSS.n683 VSS.n194 585
R241 VSS.n681 VSS.n680 585
R242 VSS.n682 VSS.n681 585
R243 VSS.n679 VSS.n196 585
R244 VSS.n196 VSS.n195 585
R245 VSS.n678 VSS.n677 585
R246 VSS.n677 VSS.n676 585
R247 VSS.n198 VSS.n197 585
R248 VSS.n675 VSS.n198 585
R249 VSS.n673 VSS.n672 585
R250 VSS.n674 VSS.n673 585
R251 VSS.n671 VSS.n200 585
R252 VSS.n200 VSS.n199 585
R253 VSS.n670 VSS.n669 585
R254 VSS.n669 VSS.n668 585
R255 VSS.n202 VSS.n201 585
R256 VSS.n667 VSS.n202 585
R257 VSS.n665 VSS.n664 585
R258 VSS.n666 VSS.n665 585
R259 VSS.n663 VSS.n204 585
R260 VSS.n204 VSS.n203 585
R261 VSS.n662 VSS.n661 585
R262 VSS.n661 VSS.n660 585
R263 VSS.n206 VSS.n205 585
R264 VSS.n659 VSS.n206 585
R265 VSS.n657 VSS.n656 585
R266 VSS.n658 VSS.n657 585
R267 VSS.n655 VSS.n208 585
R268 VSS.n208 VSS.n207 585
R269 VSS.n654 VSS.n653 585
R270 VSS.n653 VSS.n652 585
R271 VSS.n210 VSS.n209 585
R272 VSS.n651 VSS.n210 585
R273 VSS.n649 VSS.n648 585
R274 VSS.n650 VSS.n649 585
R275 VSS.n647 VSS.n212 585
R276 VSS.n212 VSS.n211 585
R277 VSS.n646 VSS.n645 585
R278 VSS.n645 VSS.n644 585
R279 VSS.n214 VSS.n213 585
R280 VSS.n643 VSS.n214 585
R281 VSS.n641 VSS.n640 585
R282 VSS.n642 VSS.n641 585
R283 VSS.n639 VSS.n216 585
R284 VSS.n216 VSS.n215 585
R285 VSS.n638 VSS.n637 585
R286 VSS.n637 VSS.n636 585
R287 VSS.n218 VSS.n217 585
R288 VSS.n635 VSS.n218 585
R289 VSS.n152 VSS.n151 585
R290 VSS.n151 VSS.n150 585
R291 VSS.n770 VSS.n769 585
R292 VSS.n771 VSS.n770 585
R293 VSS.n149 VSS.n148 585
R294 VSS.n772 VSS.n149 585
R295 VSS.n775 VSS.n774 585
R296 VSS.n774 VSS.n773 585
R297 VSS.n146 VSS.n145 585
R298 VSS.n145 VSS.n144 585
R299 VSS.n780 VSS.n779 585
R300 VSS.n781 VSS.n780 585
R301 VSS.n143 VSS.n142 585
R302 VSS.n782 VSS.n143 585
R303 VSS.n785 VSS.n784 585
R304 VSS.n784 VSS.n783 585
R305 VSS.n140 VSS.n139 585
R306 VSS.n139 VSS.n138 585
R307 VSS.n790 VSS.n789 585
R308 VSS.n791 VSS.n790 585
R309 VSS.n137 VSS.n136 585
R310 VSS.n792 VSS.n137 585
R311 VSS.n795 VSS.n794 585
R312 VSS.n794 VSS.n793 585
R313 VSS.n134 VSS.n133 585
R314 VSS.n133 VSS.n132 585
R315 VSS.n800 VSS.n799 585
R316 VSS.n801 VSS.n800 585
R317 VSS.n131 VSS.n130 585
R318 VSS.n802 VSS.n131 585
R319 VSS.n805 VSS.n804 585
R320 VSS.n804 VSS.n803 585
R321 VSS.n128 VSS.n127 585
R322 VSS.n127 VSS.n126 585
R323 VSS.n810 VSS.n809 585
R324 VSS.n811 VSS.n810 585
R325 VSS.n943 VSS.n60 585
R326 VSS.n943 VSS.n942 585
R327 VSS.n937 VSS.n61 585
R328 VSS.n941 VSS.n61 585
R329 VSS.n939 VSS.n938 585
R330 VSS.n940 VSS.n939 585
R331 VSS.n936 VSS.n63 585
R332 VSS.n63 VSS.n62 585
R333 VSS.n935 VSS.n934 585
R334 VSS.n934 VSS.n933 585
R335 VSS.n65 VSS.n64 585
R336 VSS.n932 VSS.n65 585
R337 VSS.n930 VSS.n929 585
R338 VSS.n931 VSS.n930 585
R339 VSS.n928 VSS.n67 585
R340 VSS.n67 VSS.n66 585
R341 VSS.n927 VSS.n926 585
R342 VSS.n926 VSS.n925 585
R343 VSS.n69 VSS.n68 585
R344 VSS.n924 VSS.n69 585
R345 VSS.n922 VSS.n921 585
R346 VSS.n923 VSS.n922 585
R347 VSS.n920 VSS.n71 585
R348 VSS.n71 VSS.n70 585
R349 VSS.n919 VSS.n918 585
R350 VSS.n918 VSS.n917 585
R351 VSS.n73 VSS.n72 585
R352 VSS.n916 VSS.n73 585
R353 VSS.n914 VSS.n913 585
R354 VSS.n915 VSS.n914 585
R355 VSS.n912 VSS.n75 585
R356 VSS.n75 VSS.n74 585
R357 VSS.n911 VSS.n910 585
R358 VSS.n910 VSS.n909 585
R359 VSS.n77 VSS.n76 585
R360 VSS.n908 VSS.n77 585
R361 VSS.n906 VSS.n905 585
R362 VSS.n907 VSS.n906 585
R363 VSS.n904 VSS.n79 585
R364 VSS.n79 VSS.n78 585
R365 VSS.n903 VSS.n902 585
R366 VSS.n902 VSS.n901 585
R367 VSS.n81 VSS.n80 585
R368 VSS.n900 VSS.n81 585
R369 VSS.n898 VSS.n897 585
R370 VSS.n899 VSS.n898 585
R371 VSS.n896 VSS.n83 585
R372 VSS.n83 VSS.n82 585
R373 VSS.n895 VSS.n894 585
R374 VSS.n894 VSS.n893 585
R375 VSS.n85 VSS.n84 585
R376 VSS.n892 VSS.n85 585
R377 VSS.n890 VSS.n889 585
R378 VSS.n891 VSS.n890 585
R379 VSS.n888 VSS.n87 585
R380 VSS.n87 VSS.n86 585
R381 VSS.n887 VSS.n886 585
R382 VSS.n886 VSS.n885 585
R383 VSS.n89 VSS.n88 585
R384 VSS.n884 VSS.n89 585
R385 VSS.n882 VSS.n881 585
R386 VSS.n883 VSS.n882 585
R387 VSS.n880 VSS.n91 585
R388 VSS.n91 VSS.n90 585
R389 VSS.n879 VSS.n878 585
R390 VSS.n878 VSS.n877 585
R391 VSS.n93 VSS.n92 585
R392 VSS.n876 VSS.n93 585
R393 VSS.n874 VSS.n873 585
R394 VSS.n875 VSS.n874 585
R395 VSS.n872 VSS.n95 585
R396 VSS.n95 VSS.n94 585
R397 VSS.n871 VSS.n870 585
R398 VSS.n870 VSS.n869 585
R399 VSS.n97 VSS.n96 585
R400 VSS.n868 VSS.n97 585
R401 VSS.n866 VSS.n865 585
R402 VSS.n867 VSS.n866 585
R403 VSS.n864 VSS.n99 585
R404 VSS.n99 VSS.n98 585
R405 VSS.n863 VSS.n862 585
R406 VSS.n862 VSS.n861 585
R407 VSS.n101 VSS.n100 585
R408 VSS.n860 VSS.n101 585
R409 VSS.n858 VSS.n857 585
R410 VSS.n859 VSS.n858 585
R411 VSS.n856 VSS.n103 585
R412 VSS.n103 VSS.n102 585
R413 VSS.n855 VSS.n854 585
R414 VSS.n854 VSS.n853 585
R415 VSS.n105 VSS.n104 585
R416 VSS.n852 VSS.n105 585
R417 VSS.n850 VSS.n849 585
R418 VSS.n851 VSS.n850 585
R419 VSS.n848 VSS.n107 585
R420 VSS.n107 VSS.n106 585
R421 VSS.n847 VSS.n846 585
R422 VSS.n846 VSS.n845 585
R423 VSS.n109 VSS.n108 585
R424 VSS.n844 VSS.n109 585
R425 VSS.n842 VSS.n841 585
R426 VSS.n843 VSS.n842 585
R427 VSS.n840 VSS.n111 585
R428 VSS.n111 VSS.n110 585
R429 VSS.n839 VSS.n838 585
R430 VSS.n838 VSS.n837 585
R431 VSS.n113 VSS.n112 585
R432 VSS.n836 VSS.n113 585
R433 VSS.n834 VSS.n833 585
R434 VSS.n835 VSS.n834 585
R435 VSS.n832 VSS.n115 585
R436 VSS.n115 VSS.n114 585
R437 VSS.n831 VSS.n830 585
R438 VSS.n830 VSS.n829 585
R439 VSS.n117 VSS.n116 585
R440 VSS.n828 VSS.n117 585
R441 VSS.n826 VSS.n825 585
R442 VSS.n827 VSS.n826 585
R443 VSS.n824 VSS.n119 585
R444 VSS.n119 VSS.n118 585
R445 VSS.n823 VSS.n822 585
R446 VSS.n822 VSS.n821 585
R447 VSS.n121 VSS.n120 585
R448 VSS.n820 VSS.n121 585
R449 VSS.n818 VSS.n817 585
R450 VSS.n819 VSS.n818 585
R451 VSS.n816 VSS.n123 585
R452 VSS.n123 VSS.n122 585
R453 VSS.n815 VSS.n814 585
R454 VSS.n814 VSS.n813 585
R455 VSS.n125 VSS.n124 585
R456 VSS.n812 VSS.n125 585
R457 VSS.n245 VSS.n244 585
R458 VSS.n248 VSS.n247 585
R459 VSS.n249 VSS.n243 585
R460 VSS.n243 VSS.n219 585
R461 VSS.n251 VSS.n250 585
R462 VSS.n253 VSS.n242 585
R463 VSS.n256 VSS.n255 585
R464 VSS.n257 VSS.n241 585
R465 VSS.n259 VSS.n258 585
R466 VSS.n261 VSS.n240 585
R467 VSS.n264 VSS.n263 585
R468 VSS.n265 VSS.n239 585
R469 VSS.n267 VSS.n266 585
R470 VSS.n269 VSS.n238 585
R471 VSS.n272 VSS.n271 585
R472 VSS.n273 VSS.n237 585
R473 VSS.n275 VSS.n274 585
R474 VSS.n277 VSS.n236 585
R475 VSS.n280 VSS.n279 585
R476 VSS.n281 VSS.n235 585
R477 VSS.n283 VSS.n282 585
R478 VSS.n285 VSS.n234 585
R479 VSS.n288 VSS.n287 585
R480 VSS.n289 VSS.n233 585
R481 VSS.n291 VSS.n290 585
R482 VSS.n293 VSS.n232 585
R483 VSS.n296 VSS.n295 585
R484 VSS.n297 VSS.n231 585
R485 VSS.n299 VSS.n298 585
R486 VSS.n301 VSS.n230 585
R487 VSS.n304 VSS.n303 585
R488 VSS.n305 VSS.n229 585
R489 VSS.n307 VSS.n306 585
R490 VSS.n309 VSS.n228 585
R491 VSS.n312 VSS.n311 585
R492 VSS.n313 VSS.n227 585
R493 VSS.n315 VSS.n314 585
R494 VSS.n317 VSS.n226 585
R495 VSS.n320 VSS.n319 585
R496 VSS.n321 VSS.n225 585
R497 VSS.n323 VSS.n322 585
R498 VSS.n325 VSS.n224 585
R499 VSS.n326 VSS.n223 585
R500 VSS.n329 VSS.n328 585
R501 VSS.n330 VSS.n221 585
R502 VSS.n221 VSS.n219 585
R503 VSS.n1030 VSS.n34 585
R504 VSS.n1029 VSS.n1028 585
R505 VSS.n38 VSS.n37 585
R506 VSS.n1024 VSS.n1023 585
R507 VSS.n1022 VSS.n59 585
R508 VSS.n1021 VSS.n1020 585
R509 VSS.n1019 VSS.n1018 585
R510 VSS.n1017 VSS.n1016 585
R511 VSS.n1015 VSS.n1014 585
R512 VSS.n1013 VSS.n1012 585
R513 VSS.n1011 VSS.n1010 585
R514 VSS.n1009 VSS.n1008 585
R515 VSS.n1007 VSS.n1006 585
R516 VSS.n1005 VSS.n1004 585
R517 VSS.n1003 VSS.n1002 585
R518 VSS.n1001 VSS.n1000 585
R519 VSS.n999 VSS.n998 585
R520 VSS.n997 VSS.n996 585
R521 VSS.n995 VSS.n994 585
R522 VSS.n993 VSS.n992 585
R523 VSS.n991 VSS.n990 585
R524 VSS.n989 VSS.n988 585
R525 VSS.n987 VSS.n986 585
R526 VSS.n985 VSS.n984 585
R527 VSS.n983 VSS.n982 585
R528 VSS.n981 VSS.n980 585
R529 VSS.n979 VSS.n978 585
R530 VSS.n977 VSS.n976 585
R531 VSS.n975 VSS.n974 585
R532 VSS.n973 VSS.n972 585
R533 VSS.n971 VSS.n970 585
R534 VSS.n969 VSS.n968 585
R535 VSS.n967 VSS.n966 585
R536 VSS.n965 VSS.n964 585
R537 VSS.n963 VSS.n962 585
R538 VSS.n961 VSS.n960 585
R539 VSS.n959 VSS.n958 585
R540 VSS.n957 VSS.n956 585
R541 VSS.n955 VSS.n954 585
R542 VSS.n953 VSS.n952 585
R543 VSS.n951 VSS.n950 585
R544 VSS.n949 VSS.n948 585
R545 VSS.n947 VSS.n946 585
R546 VSS.n945 VSS.n944 585
R547 VSS.n1033 VSS.n1032 585
R548 VSS.n1034 VSS.n1033 585
R549 VSS.n35 VSS.n33 585
R550 VSS.n33 VSS.n13 585
R551 VSS.n601 VSS.n600 585
R552 VSS.n602 VSS.n601 585
R553 VSS.n438 VSS.n437 585
R554 VSS.n437 VSS.n436 585
R555 VSS.n596 VSS.n595 585
R556 VSS.n595 VSS.n594 585
R557 VSS.n441 VSS.n440 585
R558 VSS.n593 VSS.n441 585
R559 VSS.n589 VSS.n588 585
R560 VSS.n590 VSS.n589 585
R561 VSS.n443 VSS.n442 585
R562 VSS.n581 VSS.n442 585
R563 VSS.n584 VSS.n583 585
R564 VSS.n583 VSS.n582 585
R565 VSS.n446 VSS.n445 585
R566 VSS.n580 VSS.n446 585
R567 VSS.n575 VSS.n574 585
R568 VSS.n576 VSS.n575 585
R569 VSS.n450 VSS.n449 585
R570 VSS.n567 VSS.n449 585
R571 VSS.n570 VSS.n569 585
R572 VSS.n569 VSS.n568 585
R573 VSS.n336 VSS.n334 585
R574 VSS.n338 VSS.n336 585
R575 VSS.n626 VSS.n625 585
R576 VSS.n625 VSS.n624 585
R577 VSS.n335 VSS.n332 585
R578 VSS.n556 VSS.n335 585
R579 VSS.n630 VSS.n222 585
R580 VSS.n555 VSS.n222 585
R581 VSS.n632 VSS.n631 585
R582 VSS.n633 VSS.n632 585
R583 VSS.n604 VSS.n603 585
R584 VSS.n603 VSS.n602 585
R585 VSS.n605 VSS.n356 585
R586 VSS.n436 VSS.n356 585
R587 VSS.n606 VSS.n355 585
R588 VSS.n594 VSS.n355 585
R589 VSS.n592 VSS.n353 585
R590 VSS.n593 VSS.n592 585
R591 VSS.n610 VSS.n352 585
R592 VSS.n590 VSS.n352 585
R593 VSS.n611 VSS.n351 585
R594 VSS.n581 VSS.n351 585
R595 VSS.n612 VSS.n350 585
R596 VSS.n582 VSS.n350 585
R597 VSS.n579 VSS.n348 585
R598 VSS.n580 VSS.n579 585
R599 VSS.n616 VSS.n347 585
R600 VSS.n576 VSS.n347 585
R601 VSS.n617 VSS.n346 585
R602 VSS.n567 VSS.n346 585
R603 VSS.n618 VSS.n345 585
R604 VSS.n568 VSS.n345 585
R605 VSS.n342 VSS.n340 585
R606 VSS.n340 VSS.n338 585
R607 VSS.n623 VSS.n622 585
R608 VSS.n624 VSS.n623 585
R609 VSS.n341 VSS.n339 585
R610 VSS.n556 VSS.n339 585
R611 VSS.n1040 VSS.n10 585
R612 VSS.n602 VSS.n10 585
R613 VSS.n1041 VSS.n9 585
R614 VSS.n436 VSS.n9 585
R615 VSS.n1042 VSS.n8 585
R616 VSS.n594 VSS.n8 585
R617 VSS.n591 VSS.n6 585
R618 VSS.n593 VSS.n591 585
R619 VSS.n1046 VSS.n5 585
R620 VSS.n590 VSS.n5 585
R621 VSS.n1047 VSS.n4 585
R622 VSS.n581 VSS.n4 585
R623 VSS.n1048 VSS.n3 585
R624 VSS.n582 VSS.n3 585
R625 VSS.n578 VSS.n2 585
R626 VSS.n580 VSS.n578 585
R627 VSS.n577 VSS.n448 585
R628 VSS.n577 VSS.n576 585
R629 VSS.n453 VSS.n447 585
R630 VSS.n567 VSS.n447 585
R631 VSS.n566 VSS.n565 585
R632 VSS.n568 VSS.n566 585
R633 VSS.n452 VSS.n451 585
R634 VSS.n451 VSS.n338 585
R635 VSS.n559 VSS.n337 585
R636 VSS.n624 VSS.n337 585
R637 VSS.n558 VSS.n557 585
R638 VSS.n557 VSS.n556 585
R639 VSS.n1038 VSS.n1037 585
R640 VSS.n12 VSS.n11 585
R641 VSS.n363 VSS.n362 585
R642 VSS.n366 VSS.n365 585
R643 VSS.n368 VSS.n367 585
R644 VSS.n370 VSS.n369 585
R645 VSS.n372 VSS.n371 585
R646 VSS.n374 VSS.n373 585
R647 VSS.n376 VSS.n375 585
R648 VSS.n378 VSS.n377 585
R649 VSS.n380 VSS.n379 585
R650 VSS.n382 VSS.n381 585
R651 VSS.n384 VSS.n383 585
R652 VSS.n386 VSS.n385 585
R653 VSS.n388 VSS.n387 585
R654 VSS.n390 VSS.n389 585
R655 VSS.n392 VSS.n391 585
R656 VSS.n394 VSS.n393 585
R657 VSS.n396 VSS.n395 585
R658 VSS.n398 VSS.n397 585
R659 VSS.n400 VSS.n399 585
R660 VSS.n403 VSS.n402 585
R661 VSS.n405 VSS.n404 585
R662 VSS.n407 VSS.n406 585
R663 VSS.n409 VSS.n408 585
R664 VSS.n411 VSS.n410 585
R665 VSS.n413 VSS.n412 585
R666 VSS.n415 VSS.n414 585
R667 VSS.n417 VSS.n416 585
R668 VSS.n419 VSS.n418 585
R669 VSS.n421 VSS.n420 585
R670 VSS.n423 VSS.n422 585
R671 VSS.n425 VSS.n424 585
R672 VSS.n427 VSS.n426 585
R673 VSS.n429 VSS.n428 585
R674 VSS.n431 VSS.n430 585
R675 VSS.n433 VSS.n432 585
R676 VSS.n435 VSS.n434 585
R677 VSS.n480 VSS.n479 585
R678 VSS.n482 VSS.n478 585
R679 VSS.n483 VSS.n477 585
R680 VSS.n483 VSS.n220 585
R681 VSS.n486 VSS.n485 585
R682 VSS.n487 VSS.n476 585
R683 VSS.n489 VSS.n488 585
R684 VSS.n491 VSS.n475 585
R685 VSS.n494 VSS.n493 585
R686 VSS.n495 VSS.n474 585
R687 VSS.n497 VSS.n496 585
R688 VSS.n499 VSS.n473 585
R689 VSS.n502 VSS.n501 585
R690 VSS.n503 VSS.n472 585
R691 VSS.n505 VSS.n504 585
R692 VSS.n507 VSS.n471 585
R693 VSS.n510 VSS.n509 585
R694 VSS.n511 VSS.n468 585
R695 VSS.n514 VSS.n513 585
R696 VSS.n516 VSS.n467 585
R697 VSS.n519 VSS.n518 585
R698 VSS.n520 VSS.n466 585
R699 VSS.n522 VSS.n521 585
R700 VSS.n524 VSS.n465 585
R701 VSS.n527 VSS.n526 585
R702 VSS.n528 VSS.n464 585
R703 VSS.n530 VSS.n529 585
R704 VSS.n532 VSS.n463 585
R705 VSS.n535 VSS.n534 585
R706 VSS.n536 VSS.n462 585
R707 VSS.n538 VSS.n537 585
R708 VSS.n540 VSS.n461 585
R709 VSS.n543 VSS.n542 585
R710 VSS.n544 VSS.n460 585
R711 VSS.n546 VSS.n545 585
R712 VSS.n548 VSS.n459 585
R713 VSS.n551 VSS.n550 585
R714 VSS.n552 VSS.n455 585
R715 VSS.n554 VSS.n553 585
R716 VSS.n554 VSS.n220 585
R717 VSS.n358 VSS.t4 563.422
R718 VSS.n360 VSS.t12 563.422
R719 VSS.n456 VSS.t8 563.422
R720 VSS.n469 VSS.t15 563.422
R721 VSS.n635 VSS.n634 480.461
R722 VSS.n942 VSS.n32 480.461
R723 VSS.n246 VSS.n219 256.663
R724 VSS.n252 VSS.n219 256.663
R725 VSS.n254 VSS.n219 256.663
R726 VSS.n260 VSS.n219 256.663
R727 VSS.n262 VSS.n219 256.663
R728 VSS.n268 VSS.n219 256.663
R729 VSS.n270 VSS.n219 256.663
R730 VSS.n276 VSS.n219 256.663
R731 VSS.n278 VSS.n219 256.663
R732 VSS.n284 VSS.n219 256.663
R733 VSS.n286 VSS.n219 256.663
R734 VSS.n292 VSS.n219 256.663
R735 VSS.n294 VSS.n219 256.663
R736 VSS.n300 VSS.n219 256.663
R737 VSS.n302 VSS.n219 256.663
R738 VSS.n308 VSS.n219 256.663
R739 VSS.n310 VSS.n219 256.663
R740 VSS.n316 VSS.n219 256.663
R741 VSS.n318 VSS.n219 256.663
R742 VSS.n324 VSS.n219 256.663
R743 VSS.n327 VSS.n219 256.663
R744 VSS.n1027 VSS.n1026 256.663
R745 VSS.n1026 VSS.n1025 256.663
R746 VSS.n1026 VSS.n58 256.663
R747 VSS.n1026 VSS.n57 256.663
R748 VSS.n1026 VSS.n56 256.663
R749 VSS.n1026 VSS.n55 256.663
R750 VSS.n1026 VSS.n54 256.663
R751 VSS.n1026 VSS.n53 256.663
R752 VSS.n1026 VSS.n52 256.663
R753 VSS.n1026 VSS.n51 256.663
R754 VSS.n1026 VSS.n50 256.663
R755 VSS.n1026 VSS.n49 256.663
R756 VSS.n1026 VSS.n48 256.663
R757 VSS.n1026 VSS.n47 256.663
R758 VSS.n1026 VSS.n46 256.663
R759 VSS.n1026 VSS.n45 256.663
R760 VSS.n1026 VSS.n44 256.663
R761 VSS.n1026 VSS.n43 256.663
R762 VSS.n1026 VSS.n42 256.663
R763 VSS.n1026 VSS.n41 256.663
R764 VSS.n1026 VSS.n40 256.663
R765 VSS.n1026 VSS.n39 256.663
R766 VSS.n1036 VSS.n1035 256.663
R767 VSS.n1035 VSS.n31 256.663
R768 VSS.n1035 VSS.n30 256.663
R769 VSS.n1035 VSS.n29 256.663
R770 VSS.n1035 VSS.n28 256.663
R771 VSS.n1035 VSS.n27 256.663
R772 VSS.n1035 VSS.n26 256.663
R773 VSS.n1035 VSS.n25 256.663
R774 VSS.n1035 VSS.n24 256.663
R775 VSS.n1035 VSS.n23 256.663
R776 VSS.n1035 VSS.n22 256.663
R777 VSS.n1035 VSS.n21 256.663
R778 VSS.n1035 VSS.n20 256.663
R779 VSS.n1035 VSS.n19 256.663
R780 VSS.n1035 VSS.n18 256.663
R781 VSS.n1035 VSS.n17 256.663
R782 VSS.n1035 VSS.n16 256.663
R783 VSS.n1035 VSS.n15 256.663
R784 VSS.n1035 VSS.n14 256.663
R785 VSS.n481 VSS.n220 256.663
R786 VSS.n484 VSS.n220 256.663
R787 VSS.n490 VSS.n220 256.663
R788 VSS.n492 VSS.n220 256.663
R789 VSS.n498 VSS.n220 256.663
R790 VSS.n500 VSS.n220 256.663
R791 VSS.n506 VSS.n220 256.663
R792 VSS.n508 VSS.n220 256.663
R793 VSS.n515 VSS.n220 256.663
R794 VSS.n517 VSS.n220 256.663
R795 VSS.n523 VSS.n220 256.663
R796 VSS.n525 VSS.n220 256.663
R797 VSS.n531 VSS.n220 256.663
R798 VSS.n533 VSS.n220 256.663
R799 VSS.n539 VSS.n220 256.663
R800 VSS.n541 VSS.n220 256.663
R801 VSS.n547 VSS.n220 256.663
R802 VSS.n549 VSS.n220 256.663
R803 VSS.n770 VSS.n151 240.244
R804 VSS.n770 VSS.n149 240.244
R805 VSS.n774 VSS.n149 240.244
R806 VSS.n774 VSS.n145 240.244
R807 VSS.n780 VSS.n145 240.244
R808 VSS.n780 VSS.n143 240.244
R809 VSS.n784 VSS.n143 240.244
R810 VSS.n784 VSS.n139 240.244
R811 VSS.n790 VSS.n139 240.244
R812 VSS.n790 VSS.n137 240.244
R813 VSS.n794 VSS.n137 240.244
R814 VSS.n794 VSS.n133 240.244
R815 VSS.n800 VSS.n133 240.244
R816 VSS.n800 VSS.n131 240.244
R817 VSS.n804 VSS.n131 240.244
R818 VSS.n804 VSS.n127 240.244
R819 VSS.n810 VSS.n127 240.244
R820 VSS.n632 VSS.n222 240.244
R821 VSS.n335 VSS.n222 240.244
R822 VSS.n625 VSS.n335 240.244
R823 VSS.n625 VSS.n336 240.244
R824 VSS.n569 VSS.n336 240.244
R825 VSS.n569 VSS.n449 240.244
R826 VSS.n575 VSS.n449 240.244
R827 VSS.n575 VSS.n446 240.244
R828 VSS.n583 VSS.n446 240.244
R829 VSS.n583 VSS.n442 240.244
R830 VSS.n589 VSS.n442 240.244
R831 VSS.n589 VSS.n441 240.244
R832 VSS.n595 VSS.n441 240.244
R833 VSS.n595 VSS.n437 240.244
R834 VSS.n601 VSS.n437 240.244
R835 VSS.n601 VSS.n33 240.244
R836 VSS.n1033 VSS.n33 240.244
R837 VSS.n623 VSS.n339 240.244
R838 VSS.n623 VSS.n340 240.244
R839 VSS.n345 VSS.n340 240.244
R840 VSS.n346 VSS.n345 240.244
R841 VSS.n347 VSS.n346 240.244
R842 VSS.n579 VSS.n347 240.244
R843 VSS.n579 VSS.n350 240.244
R844 VSS.n351 VSS.n350 240.244
R845 VSS.n352 VSS.n351 240.244
R846 VSS.n592 VSS.n352 240.244
R847 VSS.n592 VSS.n355 240.244
R848 VSS.n356 VSS.n355 240.244
R849 VSS.n603 VSS.n356 240.244
R850 VSS.n557 VSS.n337 240.244
R851 VSS.n451 VSS.n337 240.244
R852 VSS.n566 VSS.n451 240.244
R853 VSS.n566 VSS.n447 240.244
R854 VSS.n577 VSS.n447 240.244
R855 VSS.n578 VSS.n577 240.244
R856 VSS.n578 VSS.n3 240.244
R857 VSS.n4 VSS.n3 240.244
R858 VSS.n5 VSS.n4 240.244
R859 VSS.n591 VSS.n5 240.244
R860 VSS.n591 VSS.n8 240.244
R861 VSS.n9 VSS.n8 240.244
R862 VSS.n10 VSS.n9 240.244
R863 VSS.n634 VSS.n633 205.297
R864 VSS.n1034 VSS.n32 205.297
R865 VSS.n814 VSS.n125 163.367
R866 VSS.n814 VSS.n123 163.367
R867 VSS.n818 VSS.n123 163.367
R868 VSS.n818 VSS.n121 163.367
R869 VSS.n822 VSS.n121 163.367
R870 VSS.n822 VSS.n119 163.367
R871 VSS.n826 VSS.n119 163.367
R872 VSS.n826 VSS.n117 163.367
R873 VSS.n830 VSS.n117 163.367
R874 VSS.n830 VSS.n115 163.367
R875 VSS.n834 VSS.n115 163.367
R876 VSS.n834 VSS.n113 163.367
R877 VSS.n838 VSS.n113 163.367
R878 VSS.n838 VSS.n111 163.367
R879 VSS.n842 VSS.n111 163.367
R880 VSS.n842 VSS.n109 163.367
R881 VSS.n846 VSS.n109 163.367
R882 VSS.n846 VSS.n107 163.367
R883 VSS.n850 VSS.n107 163.367
R884 VSS.n850 VSS.n105 163.367
R885 VSS.n854 VSS.n105 163.367
R886 VSS.n854 VSS.n103 163.367
R887 VSS.n858 VSS.n103 163.367
R888 VSS.n858 VSS.n101 163.367
R889 VSS.n862 VSS.n101 163.367
R890 VSS.n862 VSS.n99 163.367
R891 VSS.n866 VSS.n99 163.367
R892 VSS.n866 VSS.n97 163.367
R893 VSS.n870 VSS.n97 163.367
R894 VSS.n870 VSS.n95 163.367
R895 VSS.n874 VSS.n95 163.367
R896 VSS.n874 VSS.n93 163.367
R897 VSS.n878 VSS.n93 163.367
R898 VSS.n878 VSS.n91 163.367
R899 VSS.n882 VSS.n91 163.367
R900 VSS.n882 VSS.n89 163.367
R901 VSS.n886 VSS.n89 163.367
R902 VSS.n886 VSS.n87 163.367
R903 VSS.n890 VSS.n87 163.367
R904 VSS.n890 VSS.n85 163.367
R905 VSS.n894 VSS.n85 163.367
R906 VSS.n894 VSS.n83 163.367
R907 VSS.n898 VSS.n83 163.367
R908 VSS.n898 VSS.n81 163.367
R909 VSS.n902 VSS.n81 163.367
R910 VSS.n902 VSS.n79 163.367
R911 VSS.n906 VSS.n79 163.367
R912 VSS.n906 VSS.n77 163.367
R913 VSS.n910 VSS.n77 163.367
R914 VSS.n910 VSS.n75 163.367
R915 VSS.n914 VSS.n75 163.367
R916 VSS.n914 VSS.n73 163.367
R917 VSS.n918 VSS.n73 163.367
R918 VSS.n918 VSS.n71 163.367
R919 VSS.n922 VSS.n71 163.367
R920 VSS.n922 VSS.n69 163.367
R921 VSS.n926 VSS.n69 163.367
R922 VSS.n926 VSS.n67 163.367
R923 VSS.n930 VSS.n67 163.367
R924 VSS.n930 VSS.n65 163.367
R925 VSS.n934 VSS.n65 163.367
R926 VSS.n934 VSS.n63 163.367
R927 VSS.n939 VSS.n63 163.367
R928 VSS.n939 VSS.n61 163.367
R929 VSS.n943 VSS.n61 163.367
R930 VSS.n944 VSS.n943 163.367
R931 VSS.n948 VSS.n947 163.367
R932 VSS.n952 VSS.n951 163.367
R933 VSS.n956 VSS.n955 163.367
R934 VSS.n960 VSS.n959 163.367
R935 VSS.n964 VSS.n963 163.367
R936 VSS.n968 VSS.n967 163.367
R937 VSS.n972 VSS.n971 163.367
R938 VSS.n976 VSS.n975 163.367
R939 VSS.n980 VSS.n979 163.367
R940 VSS.n984 VSS.n983 163.367
R941 VSS.n988 VSS.n987 163.367
R942 VSS.n992 VSS.n991 163.367
R943 VSS.n996 VSS.n995 163.367
R944 VSS.n1000 VSS.n999 163.367
R945 VSS.n1004 VSS.n1003 163.367
R946 VSS.n1008 VSS.n1007 163.367
R947 VSS.n1012 VSS.n1011 163.367
R948 VSS.n1016 VSS.n1015 163.367
R949 VSS.n1020 VSS.n1019 163.367
R950 VSS.n1024 VSS.n59 163.367
R951 VSS.n1028 VSS.n38 163.367
R952 VSS.n765 VSS.n154 163.367
R953 VSS.n761 VSS.n154 163.367
R954 VSS.n761 VSS.n156 163.367
R955 VSS.n757 VSS.n156 163.367
R956 VSS.n757 VSS.n158 163.367
R957 VSS.n753 VSS.n158 163.367
R958 VSS.n753 VSS.n160 163.367
R959 VSS.n749 VSS.n160 163.367
R960 VSS.n749 VSS.n162 163.367
R961 VSS.n745 VSS.n162 163.367
R962 VSS.n745 VSS.n164 163.367
R963 VSS.n741 VSS.n164 163.367
R964 VSS.n741 VSS.n166 163.367
R965 VSS.n737 VSS.n166 163.367
R966 VSS.n737 VSS.n168 163.367
R967 VSS.n733 VSS.n168 163.367
R968 VSS.n733 VSS.n170 163.367
R969 VSS.n729 VSS.n170 163.367
R970 VSS.n729 VSS.n172 163.367
R971 VSS.n725 VSS.n172 163.367
R972 VSS.n725 VSS.n174 163.367
R973 VSS.n721 VSS.n174 163.367
R974 VSS.n721 VSS.n176 163.367
R975 VSS.n717 VSS.n176 163.367
R976 VSS.n717 VSS.n178 163.367
R977 VSS.n713 VSS.n178 163.367
R978 VSS.n713 VSS.n180 163.367
R979 VSS.n709 VSS.n180 163.367
R980 VSS.n709 VSS.n182 163.367
R981 VSS.n705 VSS.n182 163.367
R982 VSS.n705 VSS.n184 163.367
R983 VSS.n701 VSS.n184 163.367
R984 VSS.n701 VSS.n186 163.367
R985 VSS.n697 VSS.n186 163.367
R986 VSS.n697 VSS.n188 163.367
R987 VSS.n693 VSS.n188 163.367
R988 VSS.n693 VSS.n190 163.367
R989 VSS.n689 VSS.n190 163.367
R990 VSS.n689 VSS.n192 163.367
R991 VSS.n685 VSS.n192 163.367
R992 VSS.n685 VSS.n194 163.367
R993 VSS.n681 VSS.n194 163.367
R994 VSS.n681 VSS.n196 163.367
R995 VSS.n677 VSS.n196 163.367
R996 VSS.n677 VSS.n198 163.367
R997 VSS.n673 VSS.n198 163.367
R998 VSS.n673 VSS.n200 163.367
R999 VSS.n669 VSS.n200 163.367
R1000 VSS.n669 VSS.n202 163.367
R1001 VSS.n665 VSS.n202 163.367
R1002 VSS.n665 VSS.n204 163.367
R1003 VSS.n661 VSS.n204 163.367
R1004 VSS.n661 VSS.n206 163.367
R1005 VSS.n657 VSS.n206 163.367
R1006 VSS.n657 VSS.n208 163.367
R1007 VSS.n653 VSS.n208 163.367
R1008 VSS.n653 VSS.n210 163.367
R1009 VSS.n649 VSS.n210 163.367
R1010 VSS.n649 VSS.n212 163.367
R1011 VSS.n645 VSS.n212 163.367
R1012 VSS.n645 VSS.n214 163.367
R1013 VSS.n641 VSS.n214 163.367
R1014 VSS.n641 VSS.n216 163.367
R1015 VSS.n637 VSS.n216 163.367
R1016 VSS.n637 VSS.n218 163.367
R1017 VSS.n245 VSS.n218 163.367
R1018 VSS.n247 VSS.n243 163.367
R1019 VSS.n251 VSS.n243 163.367
R1020 VSS.n255 VSS.n253 163.367
R1021 VSS.n259 VSS.n241 163.367
R1022 VSS.n263 VSS.n261 163.367
R1023 VSS.n267 VSS.n239 163.367
R1024 VSS.n271 VSS.n269 163.367
R1025 VSS.n275 VSS.n237 163.367
R1026 VSS.n279 VSS.n277 163.367
R1027 VSS.n283 VSS.n235 163.367
R1028 VSS.n287 VSS.n285 163.367
R1029 VSS.n291 VSS.n233 163.367
R1030 VSS.n295 VSS.n293 163.367
R1031 VSS.n299 VSS.n231 163.367
R1032 VSS.n303 VSS.n301 163.367
R1033 VSS.n307 VSS.n229 163.367
R1034 VSS.n311 VSS.n309 163.367
R1035 VSS.n315 VSS.n227 163.367
R1036 VSS.n319 VSS.n317 163.367
R1037 VSS.n323 VSS.n225 163.367
R1038 VSS.n326 VSS.n325 163.367
R1039 VSS.n328 VSS.n221 163.367
R1040 VSS.n483 VSS.n482 163.367
R1041 VSS.n485 VSS.n483 163.367
R1042 VSS.n489 VSS.n476 163.367
R1043 VSS.n493 VSS.n491 163.367
R1044 VSS.n497 VSS.n474 163.367
R1045 VSS.n501 VSS.n499 163.367
R1046 VSS.n505 VSS.n472 163.367
R1047 VSS.n509 VSS.n507 163.367
R1048 VSS.n514 VSS.n468 163.367
R1049 VSS.n518 VSS.n516 163.367
R1050 VSS.n522 VSS.n466 163.367
R1051 VSS.n526 VSS.n524 163.367
R1052 VSS.n530 VSS.n464 163.367
R1053 VSS.n534 VSS.n532 163.367
R1054 VSS.n538 VSS.n462 163.367
R1055 VSS.n542 VSS.n540 163.367
R1056 VSS.n546 VSS.n460 163.367
R1057 VSS.n550 VSS.n548 163.367
R1058 VSS.n554 VSS.n455 163.367
R1059 VSS.n432 VSS.n431 163.367
R1060 VSS.n428 VSS.n427 163.367
R1061 VSS.n424 VSS.n423 163.367
R1062 VSS.n420 VSS.n419 163.367
R1063 VSS.n416 VSS.n415 163.367
R1064 VSS.n412 VSS.n411 163.367
R1065 VSS.n408 VSS.n407 163.367
R1066 VSS.n404 VSS.n403 163.367
R1067 VSS.n399 VSS.n398 163.367
R1068 VSS.n395 VSS.n394 163.367
R1069 VSS.n391 VSS.n390 163.367
R1070 VSS.n387 VSS.n386 163.367
R1071 VSS.n383 VSS.n382 163.367
R1072 VSS.n379 VSS.n378 163.367
R1073 VSS.n375 VSS.n374 163.367
R1074 VSS.n371 VSS.n370 163.367
R1075 VSS.n367 VSS.n366 163.367
R1076 VSS.n362 VSS.n12 163.367
R1077 VSS.n358 VSS.t6 157.09
R1078 VSS.n360 VSS.t13 157.09
R1079 VSS.n456 VSS.t11 157.09
R1080 VSS.n469 VSS.t17 157.09
R1081 VSS.n359 VSS.t7 145.261
R1082 VSS.n361 VSS.t14 145.261
R1083 VSS.n457 VSS.t10 145.261
R1084 VSS.n470 VSS.t16 145.261
R1085 VSS.n556 VSS.n555 138.714
R1086 VSS.n624 VSS.n338 138.714
R1087 VSS.n568 VSS.n338 138.714
R1088 VSS.n568 VSS.n567 138.714
R1089 VSS.n582 VSS.n581 138.714
R1090 VSS.n593 VSS.n590 138.714
R1091 VSS.n594 VSS.n593 138.714
R1092 VSS.n602 VSS.n436 138.714
R1093 VSS.n602 VSS.n13 138.714
R1094 VSS.n590 VSS.t1 137.327
R1095 VSS.n556 VSS.t9 131.779
R1096 VSS.n555 VSS.n220 116.52
R1097 VSS.n1035 VSS.n13 116.52
R1098 VSS.t2 VSS.n580 109.585
R1099 VSS.n576 VSS.t0 90.1644
R1100 VSS.t5 VSS.n436 81.8416
R1101 VSS.n576 VSS.t3 79.0673
R1102 VSS.n947 VSS.n39 71.676
R1103 VSS.n951 VSS.n40 71.676
R1104 VSS.n955 VSS.n41 71.676
R1105 VSS.n959 VSS.n42 71.676
R1106 VSS.n963 VSS.n43 71.676
R1107 VSS.n967 VSS.n44 71.676
R1108 VSS.n971 VSS.n45 71.676
R1109 VSS.n975 VSS.n46 71.676
R1110 VSS.n979 VSS.n47 71.676
R1111 VSS.n983 VSS.n48 71.676
R1112 VSS.n987 VSS.n49 71.676
R1113 VSS.n991 VSS.n50 71.676
R1114 VSS.n995 VSS.n51 71.676
R1115 VSS.n999 VSS.n52 71.676
R1116 VSS.n1003 VSS.n53 71.676
R1117 VSS.n1007 VSS.n54 71.676
R1118 VSS.n1011 VSS.n55 71.676
R1119 VSS.n1015 VSS.n56 71.676
R1120 VSS.n1019 VSS.n57 71.676
R1121 VSS.n59 VSS.n58 71.676
R1122 VSS.n1025 VSS.n38 71.676
R1123 VSS.n1027 VSS.n34 71.676
R1124 VSS.n246 VSS.n245 71.676
R1125 VSS.n252 VSS.n251 71.676
R1126 VSS.n255 VSS.n254 71.676
R1127 VSS.n260 VSS.n259 71.676
R1128 VSS.n263 VSS.n262 71.676
R1129 VSS.n268 VSS.n267 71.676
R1130 VSS.n271 VSS.n270 71.676
R1131 VSS.n276 VSS.n275 71.676
R1132 VSS.n279 VSS.n278 71.676
R1133 VSS.n284 VSS.n283 71.676
R1134 VSS.n287 VSS.n286 71.676
R1135 VSS.n292 VSS.n291 71.676
R1136 VSS.n295 VSS.n294 71.676
R1137 VSS.n300 VSS.n299 71.676
R1138 VSS.n303 VSS.n302 71.676
R1139 VSS.n308 VSS.n307 71.676
R1140 VSS.n311 VSS.n310 71.676
R1141 VSS.n316 VSS.n315 71.676
R1142 VSS.n319 VSS.n318 71.676
R1143 VSS.n324 VSS.n323 71.676
R1144 VSS.n327 VSS.n326 71.676
R1145 VSS.n247 VSS.n246 71.676
R1146 VSS.n253 VSS.n252 71.676
R1147 VSS.n254 VSS.n241 71.676
R1148 VSS.n261 VSS.n260 71.676
R1149 VSS.n262 VSS.n239 71.676
R1150 VSS.n269 VSS.n268 71.676
R1151 VSS.n270 VSS.n237 71.676
R1152 VSS.n277 VSS.n276 71.676
R1153 VSS.n278 VSS.n235 71.676
R1154 VSS.n285 VSS.n284 71.676
R1155 VSS.n286 VSS.n233 71.676
R1156 VSS.n293 VSS.n292 71.676
R1157 VSS.n294 VSS.n231 71.676
R1158 VSS.n301 VSS.n300 71.676
R1159 VSS.n302 VSS.n229 71.676
R1160 VSS.n309 VSS.n308 71.676
R1161 VSS.n310 VSS.n227 71.676
R1162 VSS.n317 VSS.n316 71.676
R1163 VSS.n318 VSS.n225 71.676
R1164 VSS.n325 VSS.n324 71.676
R1165 VSS.n328 VSS.n327 71.676
R1166 VSS.n1028 VSS.n1027 71.676
R1167 VSS.n1025 VSS.n1024 71.676
R1168 VSS.n1020 VSS.n58 71.676
R1169 VSS.n1016 VSS.n57 71.676
R1170 VSS.n1012 VSS.n56 71.676
R1171 VSS.n1008 VSS.n55 71.676
R1172 VSS.n1004 VSS.n54 71.676
R1173 VSS.n1000 VSS.n53 71.676
R1174 VSS.n996 VSS.n52 71.676
R1175 VSS.n992 VSS.n51 71.676
R1176 VSS.n988 VSS.n50 71.676
R1177 VSS.n984 VSS.n49 71.676
R1178 VSS.n980 VSS.n48 71.676
R1179 VSS.n976 VSS.n47 71.676
R1180 VSS.n972 VSS.n46 71.676
R1181 VSS.n968 VSS.n45 71.676
R1182 VSS.n964 VSS.n44 71.676
R1183 VSS.n960 VSS.n43 71.676
R1184 VSS.n956 VSS.n42 71.676
R1185 VSS.n952 VSS.n41 71.676
R1186 VSS.n948 VSS.n40 71.676
R1187 VSS.n944 VSS.n39 71.676
R1188 VSS.n481 VSS.n480 71.676
R1189 VSS.n485 VSS.n484 71.676
R1190 VSS.n490 VSS.n489 71.676
R1191 VSS.n493 VSS.n492 71.676
R1192 VSS.n498 VSS.n497 71.676
R1193 VSS.n501 VSS.n500 71.676
R1194 VSS.n506 VSS.n505 71.676
R1195 VSS.n509 VSS.n508 71.676
R1196 VSS.n515 VSS.n514 71.676
R1197 VSS.n518 VSS.n517 71.676
R1198 VSS.n523 VSS.n522 71.676
R1199 VSS.n526 VSS.n525 71.676
R1200 VSS.n531 VSS.n530 71.676
R1201 VSS.n534 VSS.n533 71.676
R1202 VSS.n539 VSS.n538 71.676
R1203 VSS.n542 VSS.n541 71.676
R1204 VSS.n547 VSS.n546 71.676
R1205 VSS.n550 VSS.n549 71.676
R1206 VSS.n432 VSS.n14 71.676
R1207 VSS.n428 VSS.n15 71.676
R1208 VSS.n424 VSS.n16 71.676
R1209 VSS.n420 VSS.n17 71.676
R1210 VSS.n416 VSS.n18 71.676
R1211 VSS.n412 VSS.n19 71.676
R1212 VSS.n408 VSS.n20 71.676
R1213 VSS.n404 VSS.n21 71.676
R1214 VSS.n399 VSS.n22 71.676
R1215 VSS.n395 VSS.n23 71.676
R1216 VSS.n391 VSS.n24 71.676
R1217 VSS.n387 VSS.n25 71.676
R1218 VSS.n383 VSS.n26 71.676
R1219 VSS.n379 VSS.n27 71.676
R1220 VSS.n375 VSS.n28 71.676
R1221 VSS.n371 VSS.n29 71.676
R1222 VSS.n367 VSS.n30 71.676
R1223 VSS.n362 VSS.n31 71.676
R1224 VSS.n1037 VSS.n1036 71.676
R1225 VSS.n1036 VSS.n12 71.676
R1226 VSS.n366 VSS.n31 71.676
R1227 VSS.n370 VSS.n30 71.676
R1228 VSS.n374 VSS.n29 71.676
R1229 VSS.n378 VSS.n28 71.676
R1230 VSS.n382 VSS.n27 71.676
R1231 VSS.n386 VSS.n26 71.676
R1232 VSS.n390 VSS.n25 71.676
R1233 VSS.n394 VSS.n24 71.676
R1234 VSS.n398 VSS.n23 71.676
R1235 VSS.n403 VSS.n22 71.676
R1236 VSS.n407 VSS.n21 71.676
R1237 VSS.n411 VSS.n20 71.676
R1238 VSS.n415 VSS.n19 71.676
R1239 VSS.n419 VSS.n18 71.676
R1240 VSS.n423 VSS.n17 71.676
R1241 VSS.n427 VSS.n16 71.676
R1242 VSS.n431 VSS.n15 71.676
R1243 VSS.n435 VSS.n14 71.676
R1244 VSS.n482 VSS.n481 71.676
R1245 VSS.n484 VSS.n476 71.676
R1246 VSS.n491 VSS.n490 71.676
R1247 VSS.n492 VSS.n474 71.676
R1248 VSS.n499 VSS.n498 71.676
R1249 VSS.n500 VSS.n472 71.676
R1250 VSS.n507 VSS.n506 71.676
R1251 VSS.n508 VSS.n468 71.676
R1252 VSS.n516 VSS.n515 71.676
R1253 VSS.n517 VSS.n466 71.676
R1254 VSS.n524 VSS.n523 71.676
R1255 VSS.n525 VSS.n464 71.676
R1256 VSS.n532 VSS.n531 71.676
R1257 VSS.n533 VSS.n462 71.676
R1258 VSS.n540 VSS.n539 71.676
R1259 VSS.n541 VSS.n460 71.676
R1260 VSS.n548 VSS.n547 71.676
R1261 VSS.n549 VSS.n455 71.676
R1262 VSS.n580 VSS.t3 59.6474
R1263 VSS.n594 VSS.t5 56.8731
R1264 VSS.n567 VSS.t0 48.5503
R1265 VSS.n401 VSS.n359 46.7399
R1266 VSS.n364 VSS.n361 46.7399
R1267 VSS.n458 VSS.n457 34.3278
R1268 VSS.n512 VSS.n470 34.3278
R1269 VSS.n808 VSS.n124 30.1615
R1270 VSS.n1031 VSS.n1030 30.1615
R1271 VSS.n767 VSS.n766 30.1615
R1272 VSS.n331 VSS.n330 30.1615
R1273 VSS.n582 VSS.t2 29.1304
R1274 VSS.n634 VSS.n219 27.7433
R1275 VSS.n1026 VSS.n32 27.7433
R1276 VSS.n434 VSS.n357 26.9078
R1277 VSS.n1039 VSS.n1038 26.9078
R1278 VSS.n479 VSS.n343 26.9078
R1279 VSS.n553 VSS.n454 26.9078
R1280 VSS.n633 VSS.n220 22.1947
R1281 VSS.n1035 VSS.n1034 22.1947
R1282 VSS.n769 VSS.n152 19.3944
R1283 VSS.n769 VSS.n148 19.3944
R1284 VSS.n775 VSS.n148 19.3944
R1285 VSS.n775 VSS.n146 19.3944
R1286 VSS.n779 VSS.n146 19.3944
R1287 VSS.n779 VSS.n142 19.3944
R1288 VSS.n785 VSS.n142 19.3944
R1289 VSS.n785 VSS.n140 19.3944
R1290 VSS.n789 VSS.n140 19.3944
R1291 VSS.n789 VSS.n136 19.3944
R1292 VSS.n795 VSS.n136 19.3944
R1293 VSS.n795 VSS.n134 19.3944
R1294 VSS.n799 VSS.n134 19.3944
R1295 VSS.n799 VSS.n130 19.3944
R1296 VSS.n805 VSS.n130 19.3944
R1297 VSS.n805 VSS.n128 19.3944
R1298 VSS.n809 VSS.n128 19.3944
R1299 VSS.n631 VSS.n630 19.3944
R1300 VSS.n630 VSS.n332 19.3944
R1301 VSS.n626 VSS.n332 19.3944
R1302 VSS.n626 VSS.n334 19.3944
R1303 VSS.n570 VSS.n334 19.3944
R1304 VSS.n570 VSS.n450 19.3944
R1305 VSS.n574 VSS.n450 19.3944
R1306 VSS.n574 VSS.n445 19.3944
R1307 VSS.n584 VSS.n445 19.3944
R1308 VSS.n584 VSS.n443 19.3944
R1309 VSS.n588 VSS.n443 19.3944
R1310 VSS.n588 VSS.n440 19.3944
R1311 VSS.n596 VSS.n440 19.3944
R1312 VSS.n596 VSS.n438 19.3944
R1313 VSS.n600 VSS.n438 19.3944
R1314 VSS.n600 VSS.n35 19.3944
R1315 VSS.n1032 VSS.n35 19.3944
R1316 VSS.n622 VSS.n341 19.3944
R1317 VSS.n622 VSS.n342 19.3944
R1318 VSS.n618 VSS.n342 19.3944
R1319 VSS.n618 VSS.n617 19.3944
R1320 VSS.n617 VSS.n616 19.3944
R1321 VSS.n616 VSS.n348 19.3944
R1322 VSS.n612 VSS.n348 19.3944
R1323 VSS.n612 VSS.n611 19.3944
R1324 VSS.n611 VSS.n610 19.3944
R1325 VSS.n610 VSS.n353 19.3944
R1326 VSS.n606 VSS.n353 19.3944
R1327 VSS.n606 VSS.n605 19.3944
R1328 VSS.n605 VSS.n604 19.3944
R1329 VSS.n559 VSS.n558 19.3944
R1330 VSS.n559 VSS.n452 19.3944
R1331 VSS.n565 VSS.n452 19.3944
R1332 VSS.n565 VSS.n453 19.3944
R1333 VSS.n453 VSS.n448 19.3944
R1334 VSS.n448 VSS.n2 19.3944
R1335 VSS.n1048 VSS.n2 19.3944
R1336 VSS.n1048 VSS.n1047 19.3944
R1337 VSS.n1047 VSS.n1046 19.3944
R1338 VSS.n1046 VSS.n6 19.3944
R1339 VSS.n1042 VSS.n6 19.3944
R1340 VSS.n1042 VSS.n1041 19.3944
R1341 VSS.n1041 VSS.n1040 19.3944
R1342 VSS.n359 VSS.n358 11.8308
R1343 VSS.n361 VSS.n360 11.8308
R1344 VSS.n457 VSS.n456 11.8308
R1345 VSS.n470 VSS.n469 11.8308
R1346 VSS.n815 VSS.n124 10.6151
R1347 VSS.n816 VSS.n815 10.6151
R1348 VSS.n817 VSS.n816 10.6151
R1349 VSS.n817 VSS.n120 10.6151
R1350 VSS.n823 VSS.n120 10.6151
R1351 VSS.n824 VSS.n823 10.6151
R1352 VSS.n825 VSS.n824 10.6151
R1353 VSS.n825 VSS.n116 10.6151
R1354 VSS.n831 VSS.n116 10.6151
R1355 VSS.n832 VSS.n831 10.6151
R1356 VSS.n833 VSS.n832 10.6151
R1357 VSS.n833 VSS.n112 10.6151
R1358 VSS.n839 VSS.n112 10.6151
R1359 VSS.n840 VSS.n839 10.6151
R1360 VSS.n841 VSS.n840 10.6151
R1361 VSS.n841 VSS.n108 10.6151
R1362 VSS.n847 VSS.n108 10.6151
R1363 VSS.n848 VSS.n847 10.6151
R1364 VSS.n849 VSS.n848 10.6151
R1365 VSS.n849 VSS.n104 10.6151
R1366 VSS.n855 VSS.n104 10.6151
R1367 VSS.n856 VSS.n855 10.6151
R1368 VSS.n857 VSS.n856 10.6151
R1369 VSS.n857 VSS.n100 10.6151
R1370 VSS.n863 VSS.n100 10.6151
R1371 VSS.n864 VSS.n863 10.6151
R1372 VSS.n865 VSS.n864 10.6151
R1373 VSS.n865 VSS.n96 10.6151
R1374 VSS.n871 VSS.n96 10.6151
R1375 VSS.n872 VSS.n871 10.6151
R1376 VSS.n873 VSS.n872 10.6151
R1377 VSS.n873 VSS.n92 10.6151
R1378 VSS.n879 VSS.n92 10.6151
R1379 VSS.n880 VSS.n879 10.6151
R1380 VSS.n881 VSS.n880 10.6151
R1381 VSS.n881 VSS.n88 10.6151
R1382 VSS.n887 VSS.n88 10.6151
R1383 VSS.n888 VSS.n887 10.6151
R1384 VSS.n889 VSS.n888 10.6151
R1385 VSS.n889 VSS.n84 10.6151
R1386 VSS.n895 VSS.n84 10.6151
R1387 VSS.n896 VSS.n895 10.6151
R1388 VSS.n897 VSS.n896 10.6151
R1389 VSS.n897 VSS.n80 10.6151
R1390 VSS.n903 VSS.n80 10.6151
R1391 VSS.n904 VSS.n903 10.6151
R1392 VSS.n905 VSS.n904 10.6151
R1393 VSS.n905 VSS.n76 10.6151
R1394 VSS.n911 VSS.n76 10.6151
R1395 VSS.n912 VSS.n911 10.6151
R1396 VSS.n913 VSS.n912 10.6151
R1397 VSS.n913 VSS.n72 10.6151
R1398 VSS.n919 VSS.n72 10.6151
R1399 VSS.n920 VSS.n919 10.6151
R1400 VSS.n921 VSS.n920 10.6151
R1401 VSS.n921 VSS.n68 10.6151
R1402 VSS.n927 VSS.n68 10.6151
R1403 VSS.n928 VSS.n927 10.6151
R1404 VSS.n929 VSS.n928 10.6151
R1405 VSS.n929 VSS.n64 10.6151
R1406 VSS.n935 VSS.n64 10.6151
R1407 VSS.n936 VSS.n935 10.6151
R1408 VSS.n938 VSS.n936 10.6151
R1409 VSS.n938 VSS.n937 10.6151
R1410 VSS.n937 VSS.n60 10.6151
R1411 VSS.n945 VSS.n60 10.6151
R1412 VSS.n946 VSS.n945 10.6151
R1413 VSS.n949 VSS.n946 10.6151
R1414 VSS.n950 VSS.n949 10.6151
R1415 VSS.n953 VSS.n950 10.6151
R1416 VSS.n954 VSS.n953 10.6151
R1417 VSS.n957 VSS.n954 10.6151
R1418 VSS.n958 VSS.n957 10.6151
R1419 VSS.n961 VSS.n958 10.6151
R1420 VSS.n962 VSS.n961 10.6151
R1421 VSS.n965 VSS.n962 10.6151
R1422 VSS.n966 VSS.n965 10.6151
R1423 VSS.n969 VSS.n966 10.6151
R1424 VSS.n970 VSS.n969 10.6151
R1425 VSS.n973 VSS.n970 10.6151
R1426 VSS.n974 VSS.n973 10.6151
R1427 VSS.n977 VSS.n974 10.6151
R1428 VSS.n978 VSS.n977 10.6151
R1429 VSS.n981 VSS.n978 10.6151
R1430 VSS.n982 VSS.n981 10.6151
R1431 VSS.n985 VSS.n982 10.6151
R1432 VSS.n986 VSS.n985 10.6151
R1433 VSS.n989 VSS.n986 10.6151
R1434 VSS.n990 VSS.n989 10.6151
R1435 VSS.n993 VSS.n990 10.6151
R1436 VSS.n994 VSS.n993 10.6151
R1437 VSS.n997 VSS.n994 10.6151
R1438 VSS.n998 VSS.n997 10.6151
R1439 VSS.n1001 VSS.n998 10.6151
R1440 VSS.n1002 VSS.n1001 10.6151
R1441 VSS.n1005 VSS.n1002 10.6151
R1442 VSS.n1006 VSS.n1005 10.6151
R1443 VSS.n1009 VSS.n1006 10.6151
R1444 VSS.n1010 VSS.n1009 10.6151
R1445 VSS.n1013 VSS.n1010 10.6151
R1446 VSS.n1014 VSS.n1013 10.6151
R1447 VSS.n1017 VSS.n1014 10.6151
R1448 VSS.n1018 VSS.n1017 10.6151
R1449 VSS.n1021 VSS.n1018 10.6151
R1450 VSS.n1022 VSS.n1021 10.6151
R1451 VSS.n1023 VSS.n1022 10.6151
R1452 VSS.n1023 VSS.n37 10.6151
R1453 VSS.n1029 VSS.n37 10.6151
R1454 VSS.n1030 VSS.n1029 10.6151
R1455 VSS.n766 VSS.n153 10.6151
R1456 VSS.n760 VSS.n153 10.6151
R1457 VSS.n760 VSS.n759 10.6151
R1458 VSS.n759 VSS.n758 10.6151
R1459 VSS.n758 VSS.n157 10.6151
R1460 VSS.n752 VSS.n157 10.6151
R1461 VSS.n752 VSS.n751 10.6151
R1462 VSS.n751 VSS.n750 10.6151
R1463 VSS.n750 VSS.n161 10.6151
R1464 VSS.n744 VSS.n161 10.6151
R1465 VSS.n744 VSS.n743 10.6151
R1466 VSS.n743 VSS.n742 10.6151
R1467 VSS.n742 VSS.n165 10.6151
R1468 VSS.n736 VSS.n165 10.6151
R1469 VSS.n736 VSS.n735 10.6151
R1470 VSS.n735 VSS.n734 10.6151
R1471 VSS.n734 VSS.n169 10.6151
R1472 VSS.n728 VSS.n169 10.6151
R1473 VSS.n728 VSS.n727 10.6151
R1474 VSS.n727 VSS.n726 10.6151
R1475 VSS.n726 VSS.n173 10.6151
R1476 VSS.n720 VSS.n173 10.6151
R1477 VSS.n720 VSS.n719 10.6151
R1478 VSS.n719 VSS.n718 10.6151
R1479 VSS.n718 VSS.n177 10.6151
R1480 VSS.n712 VSS.n177 10.6151
R1481 VSS.n712 VSS.n711 10.6151
R1482 VSS.n711 VSS.n710 10.6151
R1483 VSS.n710 VSS.n181 10.6151
R1484 VSS.n704 VSS.n181 10.6151
R1485 VSS.n704 VSS.n703 10.6151
R1486 VSS.n703 VSS.n702 10.6151
R1487 VSS.n702 VSS.n185 10.6151
R1488 VSS.n696 VSS.n185 10.6151
R1489 VSS.n696 VSS.n695 10.6151
R1490 VSS.n695 VSS.n694 10.6151
R1491 VSS.n694 VSS.n189 10.6151
R1492 VSS.n688 VSS.n189 10.6151
R1493 VSS.n688 VSS.n687 10.6151
R1494 VSS.n687 VSS.n686 10.6151
R1495 VSS.n686 VSS.n193 10.6151
R1496 VSS.n680 VSS.n193 10.6151
R1497 VSS.n680 VSS.n679 10.6151
R1498 VSS.n679 VSS.n678 10.6151
R1499 VSS.n678 VSS.n197 10.6151
R1500 VSS.n672 VSS.n197 10.6151
R1501 VSS.n672 VSS.n671 10.6151
R1502 VSS.n671 VSS.n670 10.6151
R1503 VSS.n670 VSS.n201 10.6151
R1504 VSS.n664 VSS.n201 10.6151
R1505 VSS.n664 VSS.n663 10.6151
R1506 VSS.n663 VSS.n662 10.6151
R1507 VSS.n662 VSS.n205 10.6151
R1508 VSS.n656 VSS.n205 10.6151
R1509 VSS.n656 VSS.n655 10.6151
R1510 VSS.n655 VSS.n654 10.6151
R1511 VSS.n654 VSS.n209 10.6151
R1512 VSS.n648 VSS.n209 10.6151
R1513 VSS.n648 VSS.n647 10.6151
R1514 VSS.n647 VSS.n646 10.6151
R1515 VSS.n646 VSS.n213 10.6151
R1516 VSS.n640 VSS.n213 10.6151
R1517 VSS.n640 VSS.n639 10.6151
R1518 VSS.n639 VSS.n638 10.6151
R1519 VSS.n638 VSS.n217 10.6151
R1520 VSS.n244 VSS.n217 10.6151
R1521 VSS.n248 VSS.n244 10.6151
R1522 VSS.n249 VSS.n248 10.6151
R1523 VSS.n250 VSS.n249 10.6151
R1524 VSS.n250 VSS.n242 10.6151
R1525 VSS.n256 VSS.n242 10.6151
R1526 VSS.n257 VSS.n256 10.6151
R1527 VSS.n258 VSS.n257 10.6151
R1528 VSS.n258 VSS.n240 10.6151
R1529 VSS.n264 VSS.n240 10.6151
R1530 VSS.n265 VSS.n264 10.6151
R1531 VSS.n266 VSS.n265 10.6151
R1532 VSS.n266 VSS.n238 10.6151
R1533 VSS.n272 VSS.n238 10.6151
R1534 VSS.n273 VSS.n272 10.6151
R1535 VSS.n274 VSS.n273 10.6151
R1536 VSS.n274 VSS.n236 10.6151
R1537 VSS.n280 VSS.n236 10.6151
R1538 VSS.n281 VSS.n280 10.6151
R1539 VSS.n282 VSS.n281 10.6151
R1540 VSS.n282 VSS.n234 10.6151
R1541 VSS.n288 VSS.n234 10.6151
R1542 VSS.n289 VSS.n288 10.6151
R1543 VSS.n290 VSS.n289 10.6151
R1544 VSS.n290 VSS.n232 10.6151
R1545 VSS.n296 VSS.n232 10.6151
R1546 VSS.n297 VSS.n296 10.6151
R1547 VSS.n298 VSS.n297 10.6151
R1548 VSS.n298 VSS.n230 10.6151
R1549 VSS.n304 VSS.n230 10.6151
R1550 VSS.n305 VSS.n304 10.6151
R1551 VSS.n306 VSS.n305 10.6151
R1552 VSS.n306 VSS.n228 10.6151
R1553 VSS.n312 VSS.n228 10.6151
R1554 VSS.n313 VSS.n312 10.6151
R1555 VSS.n314 VSS.n313 10.6151
R1556 VSS.n314 VSS.n226 10.6151
R1557 VSS.n320 VSS.n226 10.6151
R1558 VSS.n321 VSS.n320 10.6151
R1559 VSS.n322 VSS.n321 10.6151
R1560 VSS.n322 VSS.n224 10.6151
R1561 VSS.n224 VSS.n223 10.6151
R1562 VSS.n329 VSS.n223 10.6151
R1563 VSS.n330 VSS.n329 10.6151
R1564 VSS.n434 VSS.n433 10.6151
R1565 VSS.n433 VSS.n430 10.6151
R1566 VSS.n430 VSS.n429 10.6151
R1567 VSS.n429 VSS.n426 10.6151
R1568 VSS.n426 VSS.n425 10.6151
R1569 VSS.n425 VSS.n422 10.6151
R1570 VSS.n422 VSS.n421 10.6151
R1571 VSS.n421 VSS.n418 10.6151
R1572 VSS.n418 VSS.n417 10.6151
R1573 VSS.n417 VSS.n414 10.6151
R1574 VSS.n414 VSS.n413 10.6151
R1575 VSS.n413 VSS.n410 10.6151
R1576 VSS.n410 VSS.n409 10.6151
R1577 VSS.n409 VSS.n406 10.6151
R1578 VSS.n406 VSS.n405 10.6151
R1579 VSS.n405 VSS.n402 10.6151
R1580 VSS.n400 VSS.n397 10.6151
R1581 VSS.n397 VSS.n396 10.6151
R1582 VSS.n396 VSS.n393 10.6151
R1583 VSS.n393 VSS.n392 10.6151
R1584 VSS.n392 VSS.n389 10.6151
R1585 VSS.n389 VSS.n388 10.6151
R1586 VSS.n388 VSS.n385 10.6151
R1587 VSS.n385 VSS.n384 10.6151
R1588 VSS.n384 VSS.n381 10.6151
R1589 VSS.n381 VSS.n380 10.6151
R1590 VSS.n380 VSS.n377 10.6151
R1591 VSS.n377 VSS.n376 10.6151
R1592 VSS.n376 VSS.n373 10.6151
R1593 VSS.n373 VSS.n372 10.6151
R1594 VSS.n372 VSS.n369 10.6151
R1595 VSS.n369 VSS.n368 10.6151
R1596 VSS.n368 VSS.n365 10.6151
R1597 VSS.n363 VSS.n11 10.6151
R1598 VSS.n1038 VSS.n11 10.6151
R1599 VSS.n479 VSS.n478 10.6151
R1600 VSS.n478 VSS.n477 10.6151
R1601 VSS.n486 VSS.n477 10.6151
R1602 VSS.n487 VSS.n486 10.6151
R1603 VSS.n488 VSS.n487 10.6151
R1604 VSS.n488 VSS.n475 10.6151
R1605 VSS.n494 VSS.n475 10.6151
R1606 VSS.n495 VSS.n494 10.6151
R1607 VSS.n496 VSS.n495 10.6151
R1608 VSS.n496 VSS.n473 10.6151
R1609 VSS.n502 VSS.n473 10.6151
R1610 VSS.n503 VSS.n502 10.6151
R1611 VSS.n504 VSS.n503 10.6151
R1612 VSS.n504 VSS.n471 10.6151
R1613 VSS.n510 VSS.n471 10.6151
R1614 VSS.n511 VSS.n510 10.6151
R1615 VSS.n513 VSS.n467 10.6151
R1616 VSS.n519 VSS.n467 10.6151
R1617 VSS.n520 VSS.n519 10.6151
R1618 VSS.n521 VSS.n520 10.6151
R1619 VSS.n521 VSS.n465 10.6151
R1620 VSS.n527 VSS.n465 10.6151
R1621 VSS.n528 VSS.n527 10.6151
R1622 VSS.n529 VSS.n528 10.6151
R1623 VSS.n529 VSS.n463 10.6151
R1624 VSS.n535 VSS.n463 10.6151
R1625 VSS.n536 VSS.n535 10.6151
R1626 VSS.n537 VSS.n536 10.6151
R1627 VSS.n537 VSS.n461 10.6151
R1628 VSS.n543 VSS.n461 10.6151
R1629 VSS.n544 VSS.n543 10.6151
R1630 VSS.n545 VSS.n544 10.6151
R1631 VSS.n545 VSS.n459 10.6151
R1632 VSS.n552 VSS.n551 10.6151
R1633 VSS.n553 VSS.n552 10.6151
R1634 VSS.n401 VSS.n400 9.83465
R1635 VSS.n513 VSS.n512 9.83465
R1636 VSS.n630 VSS.n629 9.3005
R1637 VSS.n628 VSS.n332 9.3005
R1638 VSS.n627 VSS.n626 9.3005
R1639 VSS.n334 VSS.n333 9.3005
R1640 VSS.n571 VSS.n570 9.3005
R1641 VSS.n572 VSS.n450 9.3005
R1642 VSS.n574 VSS.n573 9.3005
R1643 VSS.n445 VSS.n444 9.3005
R1644 VSS.n585 VSS.n584 9.3005
R1645 VSS.n586 VSS.n443 9.3005
R1646 VSS.n588 VSS.n587 9.3005
R1647 VSS.n440 VSS.n439 9.3005
R1648 VSS.n597 VSS.n596 9.3005
R1649 VSS.n598 VSS.n438 9.3005
R1650 VSS.n600 VSS.n599 9.3005
R1651 VSS.n36 VSS.n35 9.3005
R1652 VSS.n1032 VSS.n1031 9.3005
R1653 VSS.n631 VSS.n331 9.3005
R1654 VSS.n767 VSS.n152 9.3005
R1655 VSS.n769 VSS.n768 9.3005
R1656 VSS.n148 VSS.n147 9.3005
R1657 VSS.n776 VSS.n775 9.3005
R1658 VSS.n777 VSS.n146 9.3005
R1659 VSS.n779 VSS.n778 9.3005
R1660 VSS.n142 VSS.n141 9.3005
R1661 VSS.n786 VSS.n785 9.3005
R1662 VSS.n787 VSS.n140 9.3005
R1663 VSS.n789 VSS.n788 9.3005
R1664 VSS.n136 VSS.n135 9.3005
R1665 VSS.n796 VSS.n795 9.3005
R1666 VSS.n797 VSS.n134 9.3005
R1667 VSS.n799 VSS.n798 9.3005
R1668 VSS.n130 VSS.n129 9.3005
R1669 VSS.n806 VSS.n805 9.3005
R1670 VSS.n807 VSS.n128 9.3005
R1671 VSS.n809 VSS.n808 9.3005
R1672 VSS.n1047 VSS.n0 9.3005
R1673 VSS.n1046 VSS.n1045 9.3005
R1674 VSS.n1044 VSS.n6 9.3005
R1675 VSS.n1043 VSS.n1042 9.3005
R1676 VSS.n1041 VSS.n7 9.3005
R1677 VSS.n1040 VSS.n1039 9.3005
R1678 VSS.n622 VSS.n621 9.3005
R1679 VSS.n620 VSS.n342 9.3005
R1680 VSS.n619 VSS.n618 9.3005
R1681 VSS.n617 VSS.n344 9.3005
R1682 VSS.n616 VSS.n615 9.3005
R1683 VSS.n614 VSS.n348 9.3005
R1684 VSS.n613 VSS.n612 9.3005
R1685 VSS.n611 VSS.n349 9.3005
R1686 VSS.n610 VSS.n609 9.3005
R1687 VSS.n608 VSS.n353 9.3005
R1688 VSS.n607 VSS.n606 9.3005
R1689 VSS.n605 VSS.n354 9.3005
R1690 VSS.n604 VSS.n357 9.3005
R1691 VSS.n343 VSS.n341 9.3005
R1692 VSS.n560 VSS.n559 9.3005
R1693 VSS.n561 VSS.n452 9.3005
R1694 VSS.n565 VSS.n564 9.3005
R1695 VSS.n563 VSS.n453 9.3005
R1696 VSS.n562 VSS.n448 9.3005
R1697 VSS.n2 VSS.n1 9.3005
R1698 VSS.n558 VSS.n454 9.3005
R1699 VSS VSS.n1048 9.3005
R1700 VSS.n624 VSS.t9 6.93619
R1701 VSS.n364 VSS.n363 5.46391
R1702 VSS.n551 VSS.n458 5.46391
R1703 VSS.n365 VSS.n364 5.15172
R1704 VSS.n459 VSS.n458 5.15172
R1705 VSS.n581 VSS.t1 1.38764
R1706 VSS.n402 VSS.n401 0.780988
R1707 VSS.n512 VSS.n511 0.780988
R1708 VSS.n629 VSS.n331 0.152939
R1709 VSS.n629 VSS.n628 0.152939
R1710 VSS.n628 VSS.n627 0.152939
R1711 VSS.n627 VSS.n333 0.152939
R1712 VSS.n571 VSS.n333 0.152939
R1713 VSS.n572 VSS.n571 0.152939
R1714 VSS.n573 VSS.n572 0.152939
R1715 VSS.n573 VSS.n444 0.152939
R1716 VSS.n585 VSS.n444 0.152939
R1717 VSS.n586 VSS.n585 0.152939
R1718 VSS.n587 VSS.n586 0.152939
R1719 VSS.n587 VSS.n439 0.152939
R1720 VSS.n597 VSS.n439 0.152939
R1721 VSS.n598 VSS.n597 0.152939
R1722 VSS.n599 VSS.n598 0.152939
R1723 VSS.n599 VSS.n36 0.152939
R1724 VSS.n1031 VSS.n36 0.152939
R1725 VSS.n768 VSS.n767 0.152939
R1726 VSS.n768 VSS.n147 0.152939
R1727 VSS.n776 VSS.n147 0.152939
R1728 VSS.n777 VSS.n776 0.152939
R1729 VSS.n778 VSS.n777 0.152939
R1730 VSS.n778 VSS.n141 0.152939
R1731 VSS.n786 VSS.n141 0.152939
R1732 VSS.n787 VSS.n786 0.152939
R1733 VSS.n788 VSS.n787 0.152939
R1734 VSS.n788 VSS.n135 0.152939
R1735 VSS.n796 VSS.n135 0.152939
R1736 VSS.n797 VSS.n796 0.152939
R1737 VSS.n798 VSS.n797 0.152939
R1738 VSS.n798 VSS.n129 0.152939
R1739 VSS.n806 VSS.n129 0.152939
R1740 VSS.n807 VSS.n806 0.152939
R1741 VSS.n808 VSS.n807 0.152939
R1742 VSS VSS.n0 0.152939
R1743 VSS.n1045 VSS.n0 0.152939
R1744 VSS.n1045 VSS.n1044 0.152939
R1745 VSS.n1044 VSS.n1043 0.152939
R1746 VSS.n1043 VSS.n7 0.152939
R1747 VSS.n1039 VSS.n7 0.152939
R1748 VSS.n621 VSS.n343 0.152939
R1749 VSS.n621 VSS.n620 0.152939
R1750 VSS.n620 VSS.n619 0.152939
R1751 VSS.n619 VSS.n344 0.152939
R1752 VSS.n615 VSS.n344 0.152939
R1753 VSS.n615 VSS.n614 0.152939
R1754 VSS.n614 VSS.n613 0.152939
R1755 VSS.n613 VSS.n349 0.152939
R1756 VSS.n609 VSS.n349 0.152939
R1757 VSS.n609 VSS.n608 0.152939
R1758 VSS.n608 VSS.n607 0.152939
R1759 VSS.n607 VSS.n354 0.152939
R1760 VSS.n357 VSS.n354 0.152939
R1761 VSS.n560 VSS.n454 0.152939
R1762 VSS.n561 VSS.n560 0.152939
R1763 VSS.n564 VSS.n561 0.152939
R1764 VSS.n564 VSS.n563 0.152939
R1765 VSS.n563 VSS.n562 0.152939
R1766 VSS.n562 VSS.n1 0.152939
R1767 VSS VSS.n1 0.1255
R1768 VCC.n13 VCC.t4 907.707
R1769 VCC.n39 VCC.t12 907.707
R1770 VCC.n125 VCC.t8 907.707
R1771 VCC.n123 VCC.t15 907.707
R1772 VCC.n398 VCC.n10 370.245
R1773 VCC.n294 VCC.n61 370.245
R1774 VCC.n245 VCC.n88 370.245
R1775 VCC.n242 VCC.n87 370.245
R1776 VCC.n13 VCC.t6 315.521
R1777 VCC.n39 VCC.t13 315.521
R1778 VCC.n125 VCC.t11 315.521
R1779 VCC.n123 VCC.t17 315.521
R1780 VCC.n14 VCC.t7 303.69
R1781 VCC.n40 VCC.t14 303.69
R1782 VCC.n126 VCC.t10 303.69
R1783 VCC.n124 VCC.t16 303.69
R1784 VCC.n291 VCC.n61 185
R1785 VCC.n287 VCC.n61 185
R1786 VCC.n290 VCC.n289 185
R1787 VCC.n289 VCC.n288 185
R1788 VCC.n64 VCC.n63 185
R1789 VCC.n286 VCC.n64 185
R1790 VCC.n283 VCC.n282 185
R1791 VCC.n285 VCC.n283 185
R1792 VCC.n67 VCC.n66 185
R1793 VCC.n66 VCC.n65 185
R1794 VCC.n277 VCC.n276 185
R1795 VCC.n276 VCC.n275 185
R1796 VCC.n70 VCC.n69 185
R1797 VCC.n274 VCC.n70 185
R1798 VCC.n76 VCC.n71 185
R1799 VCC.n273 VCC.n71 185
R1800 VCC.n269 VCC.n268 185
R1801 VCC.n270 VCC.n269 185
R1802 VCC.n75 VCC.n74 185
R1803 VCC.n81 VCC.n74 185
R1804 VCC.n263 VCC.n262 185
R1805 VCC.n262 VCC.n261 185
R1806 VCC.n79 VCC.n78 185
R1807 VCC.n80 VCC.n79 185
R1808 VCC.n250 VCC.n249 185
R1809 VCC.n251 VCC.n250 185
R1810 VCC.n89 VCC.n88 185
R1811 VCC.n120 VCC.n88 185
R1812 VCC.n87 VCC.n86 185
R1813 VCC.n120 VCC.n87 185
R1814 VCC.n253 VCC.n252 185
R1815 VCC.n252 VCC.n251 185
R1816 VCC.n83 VCC.n82 185
R1817 VCC.n82 VCC.n80 185
R1818 VCC.n260 VCC.n259 185
R1819 VCC.n261 VCC.n260 185
R1820 VCC.n84 VCC.n72 185
R1821 VCC.n81 VCC.n72 185
R1822 VCC.n271 VCC.n73 185
R1823 VCC.n271 VCC.n270 185
R1824 VCC.n272 VCC.n2 185
R1825 VCC.n273 VCC.n272 185
R1826 VCC.n409 VCC.n3 185
R1827 VCC.n274 VCC.n3 185
R1828 VCC.n408 VCC.n4 185
R1829 VCC.n275 VCC.n4 185
R1830 VCC.n407 VCC.n5 185
R1831 VCC.n65 VCC.n5 185
R1832 VCC.n284 VCC.n6 185
R1833 VCC.n285 VCC.n284 185
R1834 VCC.n403 VCC.n8 185
R1835 VCC.n286 VCC.n8 185
R1836 VCC.n402 VCC.n9 185
R1837 VCC.n288 VCC.n9 185
R1838 VCC.n401 VCC.n10 185
R1839 VCC.n287 VCC.n10 185
R1840 VCC.n294 VCC.n293 185
R1841 VCC.n296 VCC.n59 185
R1842 VCC.n298 VCC.n297 185
R1843 VCC.n299 VCC.n58 185
R1844 VCC.n301 VCC.n300 185
R1845 VCC.n303 VCC.n56 185
R1846 VCC.n305 VCC.n304 185
R1847 VCC.n306 VCC.n55 185
R1848 VCC.n308 VCC.n307 185
R1849 VCC.n310 VCC.n53 185
R1850 VCC.n312 VCC.n311 185
R1851 VCC.n313 VCC.n52 185
R1852 VCC.n315 VCC.n314 185
R1853 VCC.n317 VCC.n50 185
R1854 VCC.n319 VCC.n318 185
R1855 VCC.n320 VCC.n49 185
R1856 VCC.n322 VCC.n321 185
R1857 VCC.n324 VCC.n47 185
R1858 VCC.n326 VCC.n325 185
R1859 VCC.n327 VCC.n46 185
R1860 VCC.n329 VCC.n328 185
R1861 VCC.n331 VCC.n44 185
R1862 VCC.n333 VCC.n332 185
R1863 VCC.n334 VCC.n43 185
R1864 VCC.n336 VCC.n335 185
R1865 VCC.n338 VCC.n41 185
R1866 VCC.n340 VCC.n339 185
R1867 VCC.n341 VCC.n38 185
R1868 VCC.n344 VCC.n343 185
R1869 VCC.n346 VCC.n36 185
R1870 VCC.n348 VCC.n347 185
R1871 VCC.n349 VCC.n35 185
R1872 VCC.n351 VCC.n350 185
R1873 VCC.n353 VCC.n33 185
R1874 VCC.n355 VCC.n354 185
R1875 VCC.n356 VCC.n32 185
R1876 VCC.n358 VCC.n357 185
R1877 VCC.n360 VCC.n30 185
R1878 VCC.n362 VCC.n361 185
R1879 VCC.n363 VCC.n29 185
R1880 VCC.n365 VCC.n364 185
R1881 VCC.n367 VCC.n27 185
R1882 VCC.n369 VCC.n368 185
R1883 VCC.n370 VCC.n26 185
R1884 VCC.n372 VCC.n371 185
R1885 VCC.n374 VCC.n24 185
R1886 VCC.n376 VCC.n375 185
R1887 VCC.n377 VCC.n23 185
R1888 VCC.n379 VCC.n378 185
R1889 VCC.n381 VCC.n21 185
R1890 VCC.n383 VCC.n382 185
R1891 VCC.n384 VCC.n20 185
R1892 VCC.n386 VCC.n385 185
R1893 VCC.n388 VCC.n18 185
R1894 VCC.n390 VCC.n389 185
R1895 VCC.n391 VCC.n17 185
R1896 VCC.n393 VCC.n392 185
R1897 VCC.n395 VCC.n16 185
R1898 VCC.n396 VCC.n11 185
R1899 VCC.n399 VCC.n398 185
R1900 VCC.n242 VCC.n241 185
R1901 VCC.n240 VCC.n122 185
R1902 VCC.n238 VCC.n121 185
R1903 VCC.n244 VCC.n121 185
R1904 VCC.n237 VCC.n236 185
R1905 VCC.n235 VCC.n234 185
R1906 VCC.n233 VCC.n232 185
R1907 VCC.n231 VCC.n230 185
R1908 VCC.n229 VCC.n228 185
R1909 VCC.n227 VCC.n226 185
R1910 VCC.n225 VCC.n224 185
R1911 VCC.n223 VCC.n222 185
R1912 VCC.n221 VCC.n220 185
R1913 VCC.n219 VCC.n218 185
R1914 VCC.n217 VCC.n216 185
R1915 VCC.n215 VCC.n214 185
R1916 VCC.n213 VCC.n212 185
R1917 VCC.n211 VCC.n210 185
R1918 VCC.n209 VCC.n208 185
R1919 VCC.n207 VCC.n206 185
R1920 VCC.n205 VCC.n204 185
R1921 VCC.n203 VCC.n202 185
R1922 VCC.n201 VCC.n200 185
R1923 VCC.n199 VCC.n198 185
R1924 VCC.n197 VCC.n196 185
R1925 VCC.n195 VCC.n194 185
R1926 VCC.n193 VCC.n192 185
R1927 VCC.n191 VCC.n190 185
R1928 VCC.n189 VCC.n188 185
R1929 VCC.n187 VCC.n186 185
R1930 VCC.n185 VCC.n184 185
R1931 VCC.n183 VCC.n182 185
R1932 VCC.n181 VCC.n180 185
R1933 VCC.n178 VCC.n177 185
R1934 VCC.n176 VCC.n175 185
R1935 VCC.n174 VCC.n173 185
R1936 VCC.n172 VCC.n171 185
R1937 VCC.n170 VCC.n169 185
R1938 VCC.n168 VCC.n167 185
R1939 VCC.n166 VCC.n165 185
R1940 VCC.n164 VCC.n163 185
R1941 VCC.n162 VCC.n161 185
R1942 VCC.n160 VCC.n159 185
R1943 VCC.n158 VCC.n157 185
R1944 VCC.n156 VCC.n155 185
R1945 VCC.n154 VCC.n153 185
R1946 VCC.n152 VCC.n151 185
R1947 VCC.n150 VCC.n149 185
R1948 VCC.n148 VCC.n147 185
R1949 VCC.n146 VCC.n145 185
R1950 VCC.n144 VCC.n143 185
R1951 VCC.n142 VCC.n141 185
R1952 VCC.n140 VCC.n139 185
R1953 VCC.n138 VCC.n137 185
R1954 VCC.n136 VCC.n135 185
R1955 VCC.n134 VCC.n133 185
R1956 VCC.n132 VCC.n131 185
R1957 VCC.n130 VCC.n129 185
R1958 VCC.n128 VCC.n127 185
R1959 VCC.n91 VCC.n90 185
R1960 VCC.n246 VCC.n245 185
R1961 VCC.n245 VCC.n244 185
R1962 VCC.n250 VCC.n88 146.341
R1963 VCC.n250 VCC.n79 146.341
R1964 VCC.n262 VCC.n79 146.341
R1965 VCC.n262 VCC.n74 146.341
R1966 VCC.n269 VCC.n74 146.341
R1967 VCC.n269 VCC.n71 146.341
R1968 VCC.n71 VCC.n70 146.341
R1969 VCC.n276 VCC.n70 146.341
R1970 VCC.n276 VCC.n66 146.341
R1971 VCC.n283 VCC.n66 146.341
R1972 VCC.n283 VCC.n64 146.341
R1973 VCC.n289 VCC.n64 146.341
R1974 VCC.n289 VCC.n61 146.341
R1975 VCC.n252 VCC.n87 146.341
R1976 VCC.n252 VCC.n82 146.341
R1977 VCC.n260 VCC.n82 146.341
R1978 VCC.n260 VCC.n72 146.341
R1979 VCC.n271 VCC.n72 146.341
R1980 VCC.n272 VCC.n271 146.341
R1981 VCC.n272 VCC.n3 146.341
R1982 VCC.n4 VCC.n3 146.341
R1983 VCC.n5 VCC.n4 146.341
R1984 VCC.n284 VCC.n5 146.341
R1985 VCC.n284 VCC.n8 146.341
R1986 VCC.n9 VCC.n8 146.341
R1987 VCC.n10 VCC.n9 146.341
R1988 VCC.n396 VCC.n395 99.5127
R1989 VCC.n393 VCC.n17 99.5127
R1990 VCC.n389 VCC.n388 99.5127
R1991 VCC.n386 VCC.n20 99.5127
R1992 VCC.n382 VCC.n381 99.5127
R1993 VCC.n379 VCC.n23 99.5127
R1994 VCC.n375 VCC.n374 99.5127
R1995 VCC.n372 VCC.n26 99.5127
R1996 VCC.n368 VCC.n367 99.5127
R1997 VCC.n365 VCC.n29 99.5127
R1998 VCC.n361 VCC.n360 99.5127
R1999 VCC.n358 VCC.n32 99.5127
R2000 VCC.n354 VCC.n353 99.5127
R2001 VCC.n351 VCC.n35 99.5127
R2002 VCC.n347 VCC.n346 99.5127
R2003 VCC.n344 VCC.n38 99.5127
R2004 VCC.n339 VCC.n338 99.5127
R2005 VCC.n336 VCC.n43 99.5127
R2006 VCC.n332 VCC.n331 99.5127
R2007 VCC.n329 VCC.n46 99.5127
R2008 VCC.n325 VCC.n324 99.5127
R2009 VCC.n322 VCC.n49 99.5127
R2010 VCC.n318 VCC.n317 99.5127
R2011 VCC.n315 VCC.n52 99.5127
R2012 VCC.n311 VCC.n310 99.5127
R2013 VCC.n308 VCC.n55 99.5127
R2014 VCC.n304 VCC.n303 99.5127
R2015 VCC.n301 VCC.n58 99.5127
R2016 VCC.n297 VCC.n296 99.5127
R2017 VCC.n122 VCC.n121 99.5127
R2018 VCC.n236 VCC.n121 99.5127
R2019 VCC.n234 VCC.n233 99.5127
R2020 VCC.n230 VCC.n229 99.5127
R2021 VCC.n226 VCC.n225 99.5127
R2022 VCC.n222 VCC.n221 99.5127
R2023 VCC.n218 VCC.n217 99.5127
R2024 VCC.n214 VCC.n213 99.5127
R2025 VCC.n210 VCC.n209 99.5127
R2026 VCC.n206 VCC.n205 99.5127
R2027 VCC.n202 VCC.n201 99.5127
R2028 VCC.n198 VCC.n197 99.5127
R2029 VCC.n194 VCC.n193 99.5127
R2030 VCC.n190 VCC.n189 99.5127
R2031 VCC.n186 VCC.n185 99.5127
R2032 VCC.n182 VCC.n181 99.5127
R2033 VCC.n177 VCC.n176 99.5127
R2034 VCC.n173 VCC.n172 99.5127
R2035 VCC.n169 VCC.n168 99.5127
R2036 VCC.n165 VCC.n164 99.5127
R2037 VCC.n161 VCC.n160 99.5127
R2038 VCC.n157 VCC.n156 99.5127
R2039 VCC.n153 VCC.n152 99.5127
R2040 VCC.n149 VCC.n148 99.5127
R2041 VCC.n145 VCC.n144 99.5127
R2042 VCC.n141 VCC.n140 99.5127
R2043 VCC.n137 VCC.n136 99.5127
R2044 VCC.n133 VCC.n132 99.5127
R2045 VCC.n129 VCC.n128 99.5127
R2046 VCC.n245 VCC.n91 99.5127
R2047 VCC.n295 VCC.n12 72.8958
R2048 VCC.n60 VCC.n12 72.8958
R2049 VCC.n302 VCC.n12 72.8958
R2050 VCC.n57 VCC.n12 72.8958
R2051 VCC.n309 VCC.n12 72.8958
R2052 VCC.n54 VCC.n12 72.8958
R2053 VCC.n316 VCC.n12 72.8958
R2054 VCC.n51 VCC.n12 72.8958
R2055 VCC.n323 VCC.n12 72.8958
R2056 VCC.n48 VCC.n12 72.8958
R2057 VCC.n330 VCC.n12 72.8958
R2058 VCC.n45 VCC.n12 72.8958
R2059 VCC.n337 VCC.n12 72.8958
R2060 VCC.n42 VCC.n12 72.8958
R2061 VCC.n345 VCC.n12 72.8958
R2062 VCC.n37 VCC.n12 72.8958
R2063 VCC.n352 VCC.n12 72.8958
R2064 VCC.n34 VCC.n12 72.8958
R2065 VCC.n359 VCC.n12 72.8958
R2066 VCC.n31 VCC.n12 72.8958
R2067 VCC.n366 VCC.n12 72.8958
R2068 VCC.n28 VCC.n12 72.8958
R2069 VCC.n373 VCC.n12 72.8958
R2070 VCC.n25 VCC.n12 72.8958
R2071 VCC.n380 VCC.n12 72.8958
R2072 VCC.n22 VCC.n12 72.8958
R2073 VCC.n387 VCC.n12 72.8958
R2074 VCC.n19 VCC.n12 72.8958
R2075 VCC.n394 VCC.n12 72.8958
R2076 VCC.n397 VCC.n12 72.8958
R2077 VCC.n244 VCC.n243 72.8958
R2078 VCC.n244 VCC.n92 72.8958
R2079 VCC.n244 VCC.n93 72.8958
R2080 VCC.n244 VCC.n94 72.8958
R2081 VCC.n244 VCC.n95 72.8958
R2082 VCC.n244 VCC.n96 72.8958
R2083 VCC.n244 VCC.n97 72.8958
R2084 VCC.n244 VCC.n98 72.8958
R2085 VCC.n244 VCC.n99 72.8958
R2086 VCC.n244 VCC.n100 72.8958
R2087 VCC.n244 VCC.n101 72.8958
R2088 VCC.n244 VCC.n102 72.8958
R2089 VCC.n244 VCC.n103 72.8958
R2090 VCC.n244 VCC.n104 72.8958
R2091 VCC.n244 VCC.n105 72.8958
R2092 VCC.n244 VCC.n106 72.8958
R2093 VCC.n244 VCC.n107 72.8958
R2094 VCC.n244 VCC.n108 72.8958
R2095 VCC.n244 VCC.n109 72.8958
R2096 VCC.n244 VCC.n110 72.8958
R2097 VCC.n244 VCC.n111 72.8958
R2098 VCC.n244 VCC.n112 72.8958
R2099 VCC.n244 VCC.n113 72.8958
R2100 VCC.n244 VCC.n114 72.8958
R2101 VCC.n244 VCC.n115 72.8958
R2102 VCC.n244 VCC.n116 72.8958
R2103 VCC.n244 VCC.n117 72.8958
R2104 VCC.n244 VCC.n118 72.8958
R2105 VCC.n244 VCC.n119 72.8958
R2106 VCC.n15 VCC.n14 41.6975
R2107 VCC.n342 VCC.n40 41.6975
R2108 VCC.n397 VCC.n396 39.2114
R2109 VCC.n394 VCC.n393 39.2114
R2110 VCC.n389 VCC.n19 39.2114
R2111 VCC.n387 VCC.n386 39.2114
R2112 VCC.n382 VCC.n22 39.2114
R2113 VCC.n380 VCC.n379 39.2114
R2114 VCC.n375 VCC.n25 39.2114
R2115 VCC.n373 VCC.n372 39.2114
R2116 VCC.n368 VCC.n28 39.2114
R2117 VCC.n366 VCC.n365 39.2114
R2118 VCC.n361 VCC.n31 39.2114
R2119 VCC.n359 VCC.n358 39.2114
R2120 VCC.n354 VCC.n34 39.2114
R2121 VCC.n352 VCC.n351 39.2114
R2122 VCC.n347 VCC.n37 39.2114
R2123 VCC.n345 VCC.n344 39.2114
R2124 VCC.n339 VCC.n42 39.2114
R2125 VCC.n337 VCC.n336 39.2114
R2126 VCC.n332 VCC.n45 39.2114
R2127 VCC.n330 VCC.n329 39.2114
R2128 VCC.n325 VCC.n48 39.2114
R2129 VCC.n323 VCC.n322 39.2114
R2130 VCC.n318 VCC.n51 39.2114
R2131 VCC.n316 VCC.n315 39.2114
R2132 VCC.n311 VCC.n54 39.2114
R2133 VCC.n309 VCC.n308 39.2114
R2134 VCC.n304 VCC.n57 39.2114
R2135 VCC.n302 VCC.n301 39.2114
R2136 VCC.n297 VCC.n60 39.2114
R2137 VCC.n295 VCC.n294 39.2114
R2138 VCC.n243 VCC.n242 39.2114
R2139 VCC.n236 VCC.n92 39.2114
R2140 VCC.n233 VCC.n93 39.2114
R2141 VCC.n229 VCC.n94 39.2114
R2142 VCC.n225 VCC.n95 39.2114
R2143 VCC.n221 VCC.n96 39.2114
R2144 VCC.n217 VCC.n97 39.2114
R2145 VCC.n213 VCC.n98 39.2114
R2146 VCC.n209 VCC.n99 39.2114
R2147 VCC.n205 VCC.n100 39.2114
R2148 VCC.n201 VCC.n101 39.2114
R2149 VCC.n197 VCC.n102 39.2114
R2150 VCC.n193 VCC.n103 39.2114
R2151 VCC.n189 VCC.n104 39.2114
R2152 VCC.n185 VCC.n105 39.2114
R2153 VCC.n181 VCC.n106 39.2114
R2154 VCC.n176 VCC.n107 39.2114
R2155 VCC.n172 VCC.n108 39.2114
R2156 VCC.n168 VCC.n109 39.2114
R2157 VCC.n164 VCC.n110 39.2114
R2158 VCC.n160 VCC.n111 39.2114
R2159 VCC.n156 VCC.n112 39.2114
R2160 VCC.n152 VCC.n113 39.2114
R2161 VCC.n148 VCC.n114 39.2114
R2162 VCC.n144 VCC.n115 39.2114
R2163 VCC.n140 VCC.n116 39.2114
R2164 VCC.n136 VCC.n117 39.2114
R2165 VCC.n132 VCC.n118 39.2114
R2166 VCC.n128 VCC.n119 39.2114
R2167 VCC.n296 VCC.n295 39.2114
R2168 VCC.n60 VCC.n58 39.2114
R2169 VCC.n303 VCC.n302 39.2114
R2170 VCC.n57 VCC.n55 39.2114
R2171 VCC.n310 VCC.n309 39.2114
R2172 VCC.n54 VCC.n52 39.2114
R2173 VCC.n317 VCC.n316 39.2114
R2174 VCC.n51 VCC.n49 39.2114
R2175 VCC.n324 VCC.n323 39.2114
R2176 VCC.n48 VCC.n46 39.2114
R2177 VCC.n331 VCC.n330 39.2114
R2178 VCC.n45 VCC.n43 39.2114
R2179 VCC.n338 VCC.n337 39.2114
R2180 VCC.n42 VCC.n38 39.2114
R2181 VCC.n346 VCC.n345 39.2114
R2182 VCC.n37 VCC.n35 39.2114
R2183 VCC.n353 VCC.n352 39.2114
R2184 VCC.n34 VCC.n32 39.2114
R2185 VCC.n360 VCC.n359 39.2114
R2186 VCC.n31 VCC.n29 39.2114
R2187 VCC.n367 VCC.n366 39.2114
R2188 VCC.n28 VCC.n26 39.2114
R2189 VCC.n374 VCC.n373 39.2114
R2190 VCC.n25 VCC.n23 39.2114
R2191 VCC.n381 VCC.n380 39.2114
R2192 VCC.n22 VCC.n20 39.2114
R2193 VCC.n388 VCC.n387 39.2114
R2194 VCC.n19 VCC.n17 39.2114
R2195 VCC.n395 VCC.n394 39.2114
R2196 VCC.n398 VCC.n397 39.2114
R2197 VCC.n243 VCC.n122 39.2114
R2198 VCC.n234 VCC.n92 39.2114
R2199 VCC.n230 VCC.n93 39.2114
R2200 VCC.n226 VCC.n94 39.2114
R2201 VCC.n222 VCC.n95 39.2114
R2202 VCC.n218 VCC.n96 39.2114
R2203 VCC.n214 VCC.n97 39.2114
R2204 VCC.n210 VCC.n98 39.2114
R2205 VCC.n206 VCC.n99 39.2114
R2206 VCC.n202 VCC.n100 39.2114
R2207 VCC.n198 VCC.n101 39.2114
R2208 VCC.n194 VCC.n102 39.2114
R2209 VCC.n190 VCC.n103 39.2114
R2210 VCC.n186 VCC.n104 39.2114
R2211 VCC.n182 VCC.n105 39.2114
R2212 VCC.n177 VCC.n106 39.2114
R2213 VCC.n173 VCC.n107 39.2114
R2214 VCC.n169 VCC.n108 39.2114
R2215 VCC.n165 VCC.n109 39.2114
R2216 VCC.n161 VCC.n110 39.2114
R2217 VCC.n157 VCC.n111 39.2114
R2218 VCC.n153 VCC.n112 39.2114
R2219 VCC.n149 VCC.n113 39.2114
R2220 VCC.n145 VCC.n114 39.2114
R2221 VCC.n141 VCC.n115 39.2114
R2222 VCC.n137 VCC.n116 39.2114
R2223 VCC.n133 VCC.n117 39.2114
R2224 VCC.n129 VCC.n118 39.2114
R2225 VCC.n119 VCC.n91 39.2114
R2226 VCC.n244 VCC.n120 33.4303
R2227 VCC.n287 VCC.n12 33.4303
R2228 VCC.n400 VCC.n399 30.7706
R2229 VCC.n293 VCC.n292 30.7706
R2230 VCC.n241 VCC.n85 30.7706
R2231 VCC.n247 VCC.n246 30.7706
R2232 VCC.n179 VCC.n126 29.2853
R2233 VCC.n239 VCC.n124 29.2853
R2234 VCC.n251 VCC.n80 21.1586
R2235 VCC.n261 VCC.n80 21.1586
R2236 VCC.n261 VCC.n81 21.1586
R2237 VCC.n275 VCC.n274 21.1586
R2238 VCC.n285 VCC.n65 21.1586
R2239 VCC.n286 VCC.n285 21.1586
R2240 VCC.n288 VCC.n287 21.1586
R2241 VCC.t2 VCC.n65 20.947
R2242 VCC.n120 VCC.t9 20.1007
R2243 VCC.n249 VCC.n89 19.3944
R2244 VCC.n249 VCC.n78 19.3944
R2245 VCC.n263 VCC.n78 19.3944
R2246 VCC.n263 VCC.n75 19.3944
R2247 VCC.n268 VCC.n75 19.3944
R2248 VCC.n268 VCC.n76 19.3944
R2249 VCC.n76 VCC.n69 19.3944
R2250 VCC.n277 VCC.n69 19.3944
R2251 VCC.n277 VCC.n67 19.3944
R2252 VCC.n282 VCC.n67 19.3944
R2253 VCC.n282 VCC.n63 19.3944
R2254 VCC.n290 VCC.n63 19.3944
R2255 VCC.n291 VCC.n290 19.3944
R2256 VCC.n253 VCC.n86 19.3944
R2257 VCC.n253 VCC.n83 19.3944
R2258 VCC.n259 VCC.n83 19.3944
R2259 VCC.n259 VCC.n84 19.3944
R2260 VCC.n84 VCC.n73 19.3944
R2261 VCC.n73 VCC.n2 19.3944
R2262 VCC.n409 VCC.n2 19.3944
R2263 VCC.n409 VCC.n408 19.3944
R2264 VCC.n408 VCC.n407 19.3944
R2265 VCC.n407 VCC.n6 19.3944
R2266 VCC.n403 VCC.n6 19.3944
R2267 VCC.n403 VCC.n402 19.3944
R2268 VCC.n402 VCC.n401 19.3944
R2269 VCC.t3 VCC.n273 16.7154
R2270 VCC.n270 VCC.t0 13.7533
R2271 VCC.n288 VCC.t5 12.4838
R2272 VCC.n270 VCC.t1 12.0606
R2273 VCC.n14 VCC.n13 11.8308
R2274 VCC.n40 VCC.n39 11.8308
R2275 VCC.n126 VCC.n125 11.8308
R2276 VCC.n124 VCC.n123 11.8308
R2277 VCC.n399 VCC.n11 10.6151
R2278 VCC.n392 VCC.n16 10.6151
R2279 VCC.n392 VCC.n391 10.6151
R2280 VCC.n391 VCC.n390 10.6151
R2281 VCC.n390 VCC.n18 10.6151
R2282 VCC.n385 VCC.n18 10.6151
R2283 VCC.n385 VCC.n384 10.6151
R2284 VCC.n384 VCC.n383 10.6151
R2285 VCC.n383 VCC.n21 10.6151
R2286 VCC.n378 VCC.n21 10.6151
R2287 VCC.n378 VCC.n377 10.6151
R2288 VCC.n377 VCC.n376 10.6151
R2289 VCC.n376 VCC.n24 10.6151
R2290 VCC.n371 VCC.n24 10.6151
R2291 VCC.n371 VCC.n370 10.6151
R2292 VCC.n370 VCC.n369 10.6151
R2293 VCC.n369 VCC.n27 10.6151
R2294 VCC.n364 VCC.n27 10.6151
R2295 VCC.n364 VCC.n363 10.6151
R2296 VCC.n363 VCC.n362 10.6151
R2297 VCC.n362 VCC.n30 10.6151
R2298 VCC.n357 VCC.n30 10.6151
R2299 VCC.n357 VCC.n356 10.6151
R2300 VCC.n356 VCC.n355 10.6151
R2301 VCC.n355 VCC.n33 10.6151
R2302 VCC.n350 VCC.n33 10.6151
R2303 VCC.n350 VCC.n349 10.6151
R2304 VCC.n349 VCC.n348 10.6151
R2305 VCC.n348 VCC.n36 10.6151
R2306 VCC.n343 VCC.n36 10.6151
R2307 VCC.n341 VCC.n340 10.6151
R2308 VCC.n340 VCC.n41 10.6151
R2309 VCC.n335 VCC.n41 10.6151
R2310 VCC.n335 VCC.n334 10.6151
R2311 VCC.n334 VCC.n333 10.6151
R2312 VCC.n333 VCC.n44 10.6151
R2313 VCC.n328 VCC.n44 10.6151
R2314 VCC.n328 VCC.n327 10.6151
R2315 VCC.n327 VCC.n326 10.6151
R2316 VCC.n326 VCC.n47 10.6151
R2317 VCC.n321 VCC.n47 10.6151
R2318 VCC.n321 VCC.n320 10.6151
R2319 VCC.n320 VCC.n319 10.6151
R2320 VCC.n319 VCC.n50 10.6151
R2321 VCC.n314 VCC.n50 10.6151
R2322 VCC.n314 VCC.n313 10.6151
R2323 VCC.n313 VCC.n312 10.6151
R2324 VCC.n312 VCC.n53 10.6151
R2325 VCC.n307 VCC.n53 10.6151
R2326 VCC.n307 VCC.n306 10.6151
R2327 VCC.n306 VCC.n305 10.6151
R2328 VCC.n305 VCC.n56 10.6151
R2329 VCC.n300 VCC.n56 10.6151
R2330 VCC.n300 VCC.n299 10.6151
R2331 VCC.n299 VCC.n298 10.6151
R2332 VCC.n298 VCC.n59 10.6151
R2333 VCC.n293 VCC.n59 10.6151
R2334 VCC.n241 VCC.n240 10.6151
R2335 VCC.n238 VCC.n237 10.6151
R2336 VCC.n237 VCC.n235 10.6151
R2337 VCC.n235 VCC.n232 10.6151
R2338 VCC.n232 VCC.n231 10.6151
R2339 VCC.n231 VCC.n228 10.6151
R2340 VCC.n228 VCC.n227 10.6151
R2341 VCC.n227 VCC.n224 10.6151
R2342 VCC.n224 VCC.n223 10.6151
R2343 VCC.n223 VCC.n220 10.6151
R2344 VCC.n220 VCC.n219 10.6151
R2345 VCC.n219 VCC.n216 10.6151
R2346 VCC.n216 VCC.n215 10.6151
R2347 VCC.n215 VCC.n212 10.6151
R2348 VCC.n212 VCC.n211 10.6151
R2349 VCC.n211 VCC.n208 10.6151
R2350 VCC.n208 VCC.n207 10.6151
R2351 VCC.n207 VCC.n204 10.6151
R2352 VCC.n204 VCC.n203 10.6151
R2353 VCC.n203 VCC.n200 10.6151
R2354 VCC.n200 VCC.n199 10.6151
R2355 VCC.n199 VCC.n196 10.6151
R2356 VCC.n196 VCC.n195 10.6151
R2357 VCC.n195 VCC.n192 10.6151
R2358 VCC.n192 VCC.n191 10.6151
R2359 VCC.n191 VCC.n188 10.6151
R2360 VCC.n188 VCC.n187 10.6151
R2361 VCC.n187 VCC.n184 10.6151
R2362 VCC.n184 VCC.n183 10.6151
R2363 VCC.n183 VCC.n180 10.6151
R2364 VCC.n178 VCC.n175 10.6151
R2365 VCC.n175 VCC.n174 10.6151
R2366 VCC.n174 VCC.n171 10.6151
R2367 VCC.n171 VCC.n170 10.6151
R2368 VCC.n170 VCC.n167 10.6151
R2369 VCC.n167 VCC.n166 10.6151
R2370 VCC.n166 VCC.n163 10.6151
R2371 VCC.n163 VCC.n162 10.6151
R2372 VCC.n162 VCC.n159 10.6151
R2373 VCC.n159 VCC.n158 10.6151
R2374 VCC.n158 VCC.n155 10.6151
R2375 VCC.n155 VCC.n154 10.6151
R2376 VCC.n154 VCC.n151 10.6151
R2377 VCC.n151 VCC.n150 10.6151
R2378 VCC.n150 VCC.n147 10.6151
R2379 VCC.n147 VCC.n146 10.6151
R2380 VCC.n146 VCC.n143 10.6151
R2381 VCC.n143 VCC.n142 10.6151
R2382 VCC.n142 VCC.n139 10.6151
R2383 VCC.n139 VCC.n138 10.6151
R2384 VCC.n138 VCC.n135 10.6151
R2385 VCC.n135 VCC.n134 10.6151
R2386 VCC.n134 VCC.n131 10.6151
R2387 VCC.n131 VCC.n130 10.6151
R2388 VCC.n130 VCC.n127 10.6151
R2389 VCC.n127 VCC.n90 10.6151
R2390 VCC.n246 VCC.n90 10.6151
R2391 VCC.n343 VCC.n342 9.83465
R2392 VCC.n180 VCC.n179 9.83465
R2393 VCC.n408 VCC.n0 9.3005
R2394 VCC.n407 VCC.n406 9.3005
R2395 VCC.n405 VCC.n6 9.3005
R2396 VCC.n404 VCC.n403 9.3005
R2397 VCC.n402 VCC.n7 9.3005
R2398 VCC.n401 VCC.n400 9.3005
R2399 VCC.n249 VCC.n248 9.3005
R2400 VCC.n78 VCC.n77 9.3005
R2401 VCC.n264 VCC.n263 9.3005
R2402 VCC.n265 VCC.n75 9.3005
R2403 VCC.n268 VCC.n267 9.3005
R2404 VCC.n266 VCC.n76 9.3005
R2405 VCC.n69 VCC.n68 9.3005
R2406 VCC.n278 VCC.n277 9.3005
R2407 VCC.n279 VCC.n67 9.3005
R2408 VCC.n282 VCC.n281 9.3005
R2409 VCC.n280 VCC.n63 9.3005
R2410 VCC.n290 VCC.n62 9.3005
R2411 VCC.n292 VCC.n291 9.3005
R2412 VCC.n247 VCC.n89 9.3005
R2413 VCC.n86 VCC.n85 9.3005
R2414 VCC.n254 VCC.n253 9.3005
R2415 VCC.n255 VCC.n83 9.3005
R2416 VCC.n259 VCC.n258 9.3005
R2417 VCC.n257 VCC.n84 9.3005
R2418 VCC.n256 VCC.n73 9.3005
R2419 VCC.n2 VCC.n1 9.3005
R2420 VCC VCC.n409 9.3005
R2421 VCC.n273 VCC.t1 9.09849
R2422 VCC.t5 VCC.n286 8.67533
R2423 VCC.n15 VCC.n11 7.96148
R2424 VCC.n240 VCC.n239 7.96148
R2425 VCC.n81 VCC.t0 7.40585
R2426 VCC.n274 VCC.t3 4.44371
R2427 VCC.n16 VCC.n15 2.65416
R2428 VCC.n239 VCC.n238 2.65416
R2429 VCC.n251 VCC.t9 1.05841
R2430 VCC.n342 VCC.n341 0.780988
R2431 VCC.n179 VCC.n178 0.780988
R2432 VCC.n275 VCC.t2 0.212081
R2433 VCC VCC.n0 0.152939
R2434 VCC.n406 VCC.n0 0.152939
R2435 VCC.n406 VCC.n405 0.152939
R2436 VCC.n405 VCC.n404 0.152939
R2437 VCC.n404 VCC.n7 0.152939
R2438 VCC.n400 VCC.n7 0.152939
R2439 VCC.n248 VCC.n247 0.152939
R2440 VCC.n248 VCC.n77 0.152939
R2441 VCC.n264 VCC.n77 0.152939
R2442 VCC.n265 VCC.n264 0.152939
R2443 VCC.n267 VCC.n265 0.152939
R2444 VCC.n267 VCC.n266 0.152939
R2445 VCC.n266 VCC.n68 0.152939
R2446 VCC.n278 VCC.n68 0.152939
R2447 VCC.n279 VCC.n278 0.152939
R2448 VCC.n281 VCC.n279 0.152939
R2449 VCC.n281 VCC.n280 0.152939
R2450 VCC.n280 VCC.n62 0.152939
R2451 VCC.n292 VCC.n62 0.152939
R2452 VCC.n254 VCC.n85 0.152939
R2453 VCC.n255 VCC.n254 0.152939
R2454 VCC.n258 VCC.n255 0.152939
R2455 VCC.n258 VCC.n257 0.152939
R2456 VCC.n257 VCC.n256 0.152939
R2457 VCC.n256 VCC.n1 0.152939
R2458 VCC VCC.n1 0.1255
R2459 VOUT.n83 VOUT.t0 824.564
R2460 VOUT.n88 VOUT.t32 824.564
R2461 VOUT.n64 VOUT.t29 824.564
R2462 VOUT.n69 VOUT.t20 824.564
R2463 VOUT.n82 VOUT.t27 800.465
R2464 VOUT.n87 VOUT.t34 800.465
R2465 VOUT.n63 VOUT.t13 800.465
R2466 VOUT.n68 VOUT.t22 800.465
R2467 VOUT.n221 VOUT.n185 756.745
R2468 VOUT.n35 VOUT.n34 756.745
R2469 VOUT.n170 VOUT.n134 756.745
R2470 VOUT.n128 VOUT.n92 756.745
R2471 VOUT.n197 VOUT.n196 585
R2472 VOUT.n202 VOUT.n201 585
R2473 VOUT.n204 VOUT.n203 585
R2474 VOUT.n193 VOUT.n192 585
R2475 VOUT.n210 VOUT.n209 585
R2476 VOUT.n212 VOUT.n211 585
R2477 VOUT.n189 VOUT.n188 585
R2478 VOUT.n219 VOUT.n218 585
R2479 VOUT.n220 VOUT.n187 585
R2480 VOUT.n222 VOUT.n221 585
R2481 VOUT.n59 VOUT.n58 585
R2482 VOUT.n22 VOUT.n21 585
R2483 VOUT.n53 VOUT.n52 585
R2484 VOUT.n51 VOUT.n50 585
R2485 VOUT.n26 VOUT.n25 585
R2486 VOUT.n45 VOUT.n44 585
R2487 VOUT.n43 VOUT.n42 585
R2488 VOUT.n30 VOUT.n29 585
R2489 VOUT.n37 VOUT.n36 585
R2490 VOUT.n35 VOUT.n32 585
R2491 VOUT.n146 VOUT.n145 585
R2492 VOUT.n151 VOUT.n150 585
R2493 VOUT.n153 VOUT.n152 585
R2494 VOUT.n142 VOUT.n141 585
R2495 VOUT.n159 VOUT.n158 585
R2496 VOUT.n161 VOUT.n160 585
R2497 VOUT.n138 VOUT.n137 585
R2498 VOUT.n168 VOUT.n167 585
R2499 VOUT.n169 VOUT.n136 585
R2500 VOUT.n171 VOUT.n170 585
R2501 VOUT.n104 VOUT.n103 585
R2502 VOUT.n109 VOUT.n108 585
R2503 VOUT.n111 VOUT.n110 585
R2504 VOUT.n100 VOUT.n99 585
R2505 VOUT.n117 VOUT.n116 585
R2506 VOUT.n119 VOUT.n118 585
R2507 VOUT.n96 VOUT.n95 585
R2508 VOUT.n126 VOUT.n125 585
R2509 VOUT.n127 VOUT.n94 585
R2510 VOUT.n129 VOUT.n128 585
R2511 VOUT.n78 VOUT.t7 480.279
R2512 VOUT.n73 VOUT.t24 480.279
R2513 VOUT.n7 VOUT.t15 480.279
R2514 VOUT.n2 VOUT.t17 480.279
R2515 VOUT.n77 VOUT.t9 456.18
R2516 VOUT.n72 VOUT.t11 456.18
R2517 VOUT.n6 VOUT.t3 456.18
R2518 VOUT.n1 VOUT.t5 456.18
R2519 VOUT.n198 VOUT.t2 329.043
R2520 VOUT.t33 VOUT.n20 329.043
R2521 VOUT.n147 VOUT.t31 329.043
R2522 VOUT.n105 VOUT.t21 329.043
R2523 VOUT.n265 VOUT.n251 289.615
R2524 VOUT.n234 VOUT.n232 289.615
R2525 VOUT.n286 VOUT.n272 289.615
R2526 VOUT.n306 VOUT.n11 289.615
R2527 VOUT.n266 VOUT.n265 185
R2528 VOUT.n264 VOUT.n263 185
R2529 VOUT.n255 VOUT.n254 185
R2530 VOUT.n258 VOUT.n257 185
R2531 VOUT.n233 VOUT.n232 185
R2532 VOUT.n241 VOUT.n240 185
R2533 VOUT.n243 VOUT.n242 185
R2534 VOUT.n245 VOUT.n229 185
R2535 VOUT.n287 VOUT.n286 185
R2536 VOUT.n285 VOUT.n284 185
R2537 VOUT.n276 VOUT.n275 185
R2538 VOUT.n279 VOUT.n278 185
R2539 VOUT.n307 VOUT.n306 185
R2540 VOUT.n305 VOUT.n304 185
R2541 VOUT.n15 VOUT.n14 185
R2542 VOUT.n299 VOUT.n298 185
R2543 VOUT.n202 VOUT.n196 171.744
R2544 VOUT.n203 VOUT.n202 171.744
R2545 VOUT.n203 VOUT.n192 171.744
R2546 VOUT.n210 VOUT.n192 171.744
R2547 VOUT.n211 VOUT.n210 171.744
R2548 VOUT.n211 VOUT.n188 171.744
R2549 VOUT.n219 VOUT.n188 171.744
R2550 VOUT.n220 VOUT.n219 171.744
R2551 VOUT.n221 VOUT.n220 171.744
R2552 VOUT.n59 VOUT.n21 171.744
R2553 VOUT.n52 VOUT.n21 171.744
R2554 VOUT.n52 VOUT.n51 171.744
R2555 VOUT.n51 VOUT.n25 171.744
R2556 VOUT.n44 VOUT.n25 171.744
R2557 VOUT.n44 VOUT.n43 171.744
R2558 VOUT.n43 VOUT.n29 171.744
R2559 VOUT.n36 VOUT.n29 171.744
R2560 VOUT.n36 VOUT.n35 171.744
R2561 VOUT.n151 VOUT.n145 171.744
R2562 VOUT.n152 VOUT.n151 171.744
R2563 VOUT.n152 VOUT.n141 171.744
R2564 VOUT.n159 VOUT.n141 171.744
R2565 VOUT.n160 VOUT.n159 171.744
R2566 VOUT.n160 VOUT.n137 171.744
R2567 VOUT.n168 VOUT.n137 171.744
R2568 VOUT.n169 VOUT.n168 171.744
R2569 VOUT.n170 VOUT.n169 171.744
R2570 VOUT.n109 VOUT.n103 171.744
R2571 VOUT.n110 VOUT.n109 171.744
R2572 VOUT.n110 VOUT.n99 171.744
R2573 VOUT.n117 VOUT.n99 171.744
R2574 VOUT.n118 VOUT.n117 171.744
R2575 VOUT.n118 VOUT.n95 171.744
R2576 VOUT.n126 VOUT.n95 171.744
R2577 VOUT.n127 VOUT.n126 171.744
R2578 VOUT.n128 VOUT.n127 171.744
R2579 VOUT.n74 VOUT.n73 161.489
R2580 VOUT.n84 VOUT.n83 161.489
R2581 VOUT.n65 VOUT.n64 161.489
R2582 VOUT.n3 VOUT.n2 161.489
R2583 VOUT.n75 VOUT.n74 161.3
R2584 VOUT.n76 VOUT.n71 161.3
R2585 VOUT.n79 VOUT.n78 161.3
R2586 VOUT.n85 VOUT.n84 161.3
R2587 VOUT.n86 VOUT.n81 161.3
R2588 VOUT.n89 VOUT.n88 161.3
R2589 VOUT.n70 VOUT.n69 161.3
R2590 VOUT.n67 VOUT.n62 161.3
R2591 VOUT.n66 VOUT.n65 161.3
R2592 VOUT.n4 VOUT.n3 161.3
R2593 VOUT.n5 VOUT.n0 161.3
R2594 VOUT.n8 VOUT.n7 161.3
R2595 VOUT.t26 VOUT.n256 147.888
R2596 VOUT.t8 VOUT.n246 147.888
R2597 VOUT.t19 VOUT.n277 147.888
R2598 VOUT.t16 VOUT.n16 147.888
R2599 VOUT.n265 VOUT.n264 104.615
R2600 VOUT.n264 VOUT.n254 104.615
R2601 VOUT.n257 VOUT.n254 104.615
R2602 VOUT.n241 VOUT.n232 104.615
R2603 VOUT.n242 VOUT.n241 104.615
R2604 VOUT.n242 VOUT.n229 104.615
R2605 VOUT.n286 VOUT.n285 104.615
R2606 VOUT.n285 VOUT.n275 104.615
R2607 VOUT.n278 VOUT.n275 104.615
R2608 VOUT.n306 VOUT.n305 104.615
R2609 VOUT.n305 VOUT.n14 104.615
R2610 VOUT.n298 VOUT.n14 104.615
R2611 VOUT.n179 VOUT.n61 86.7637
R2612 VOUT.n181 VOUT.n60 86.7637
R2613 VOUT.n179 VOUT.n178 86.2379
R2614 VOUT.n182 VOUT.n181 86.2379
R2615 VOUT.t2 VOUT.n196 85.8723
R2616 VOUT.t33 VOUT.n59 85.8723
R2617 VOUT.t31 VOUT.n145 85.8723
R2618 VOUT.t21 VOUT.n103 85.8723
R2619 VOUT.n247 VOUT.n17 77.093
R2620 VOUT.n297 VOUT.n296 77.093
R2621 VOUT.n248 VOUT.n17 76.5671
R2622 VOUT.n296 VOUT.n295 76.5671
R2623 VOUT.n76 VOUT.n75 73.0308
R2624 VOUT.n86 VOUT.n85 73.0308
R2625 VOUT.n67 VOUT.n66 73.0308
R2626 VOUT.n5 VOUT.n4 73.0308
R2627 VOUT.n184 VOUT.n183 69.5591
R2628 VOUT.n177 VOUT.n176 69.5591
R2629 VOUT.n78 VOUT.n77 64.9975
R2630 VOUT.n73 VOUT.n72 64.9975
R2631 VOUT.n88 VOUT.n87 64.9975
R2632 VOUT.n83 VOUT.n82 64.9975
R2633 VOUT.n69 VOUT.n68 64.9975
R2634 VOUT.n64 VOUT.n63 64.9975
R2635 VOUT.n7 VOUT.n6 64.9975
R2636 VOUT.n2 VOUT.n1 64.9975
R2637 VOUT.n250 VOUT.n249 59.8883
R2638 VOUT.n294 VOUT.n10 59.8883
R2639 VOUT.n257 VOUT.t26 52.3082
R2640 VOUT.t8 VOUT.n229 52.3082
R2641 VOUT.n278 VOUT.t19 52.3082
R2642 VOUT.n298 VOUT.t16 52.3082
R2643 VOUT.n184 VOUT.n19 36.59
R2644 VOUT.n226 VOUT.n225 36.0641
R2645 VOUT.n175 VOUT.n174 36.0641
R2646 VOUT.n133 VOUT.n132 36.0641
R2647 VOUT.n250 VOUT.n228 35.8142
R2648 VOUT.n270 VOUT.n269 35.2884
R2649 VOUT.n291 VOUT.n290 35.2884
R2650 VOUT.n311 VOUT.n310 35.2884
R2651 VOUT.n258 VOUT.n256 15.6496
R2652 VOUT.n246 VOUT.n245 15.6496
R2653 VOUT.n279 VOUT.n277 15.6496
R2654 VOUT.n299 VOUT.n16 15.6496
R2655 VOUT.n181 VOUT.n180 15.0264
R2656 VOUT.n293 VOUT.n17 13.3022
R2657 VOUT.n222 VOUT.n187 13.1884
R2658 VOUT.n37 VOUT.n32 13.1884
R2659 VOUT.n171 VOUT.n136 13.1884
R2660 VOUT.n129 VOUT.n94 13.1884
R2661 VOUT.n218 VOUT.n217 12.8005
R2662 VOUT.n223 VOUT.n185 12.8005
R2663 VOUT.n38 VOUT.n30 12.8005
R2664 VOUT.n34 VOUT.n33 12.8005
R2665 VOUT.n259 VOUT.n255 12.8005
R2666 VOUT.n244 VOUT.n243 12.8005
R2667 VOUT.n280 VOUT.n276 12.8005
R2668 VOUT.n300 VOUT.n15 12.8005
R2669 VOUT.n167 VOUT.n166 12.8005
R2670 VOUT.n172 VOUT.n134 12.8005
R2671 VOUT.n125 VOUT.n124 12.8005
R2672 VOUT.n130 VOUT.n92 12.8005
R2673 VOUT.n216 VOUT.n189 12.0247
R2674 VOUT.n42 VOUT.n41 12.0247
R2675 VOUT.n263 VOUT.n262 12.0247
R2676 VOUT.n240 VOUT.n231 12.0247
R2677 VOUT.n284 VOUT.n283 12.0247
R2678 VOUT.n304 VOUT.n303 12.0247
R2679 VOUT.n165 VOUT.n138 12.0247
R2680 VOUT.n123 VOUT.n96 12.0247
R2681 VOUT.n213 VOUT.n212 11.249
R2682 VOUT.n45 VOUT.n28 11.249
R2683 VOUT.n266 VOUT.n253 11.249
R2684 VOUT.n239 VOUT.n233 11.249
R2685 VOUT.n287 VOUT.n274 11.249
R2686 VOUT.n307 VOUT.n13 11.249
R2687 VOUT.n162 VOUT.n161 11.249
R2688 VOUT.n120 VOUT.n119 11.249
R2689 VOUT.n198 VOUT.n197 10.7238
R2690 VOUT.n58 VOUT.n20 10.7238
R2691 VOUT.n147 VOUT.n146 10.7238
R2692 VOUT.n105 VOUT.n104 10.7238
R2693 VOUT.n209 VOUT.n191 10.4732
R2694 VOUT.n46 VOUT.n26 10.4732
R2695 VOUT.n267 VOUT.n251 10.4732
R2696 VOUT.n235 VOUT.n234 10.4732
R2697 VOUT.n288 VOUT.n272 10.4732
R2698 VOUT.n308 VOUT.n11 10.4732
R2699 VOUT.n158 VOUT.n140 10.4732
R2700 VOUT.n116 VOUT.n98 10.4732
R2701 VOUT.n208 VOUT.n193 9.69747
R2702 VOUT.n50 VOUT.n49 9.69747
R2703 VOUT.n157 VOUT.n142 9.69747
R2704 VOUT.n115 VOUT.n100 9.69747
R2705 VOUT.n225 VOUT.n224 9.45567
R2706 VOUT.n31 VOUT.n19 9.45567
R2707 VOUT.n269 VOUT.n268 9.45567
R2708 VOUT.n236 VOUT.n228 9.45567
R2709 VOUT.n290 VOUT.n289 9.45567
R2710 VOUT.n310 VOUT.n309 9.45567
R2711 VOUT.n174 VOUT.n173 9.45567
R2712 VOUT.n132 VOUT.n131 9.45567
R2713 VOUT.n224 VOUT.n223 9.3005
R2714 VOUT.n200 VOUT.n199 9.3005
R2715 VOUT.n195 VOUT.n194 9.3005
R2716 VOUT.n206 VOUT.n205 9.3005
R2717 VOUT.n208 VOUT.n207 9.3005
R2718 VOUT.n191 VOUT.n190 9.3005
R2719 VOUT.n214 VOUT.n213 9.3005
R2720 VOUT.n216 VOUT.n215 9.3005
R2721 VOUT.n217 VOUT.n186 9.3005
R2722 VOUT.n33 VOUT.n31 9.3005
R2723 VOUT.n57 VOUT.n56 9.3005
R2724 VOUT.n55 VOUT.n54 9.3005
R2725 VOUT.n24 VOUT.n23 9.3005
R2726 VOUT.n49 VOUT.n48 9.3005
R2727 VOUT.n47 VOUT.n46 9.3005
R2728 VOUT.n28 VOUT.n27 9.3005
R2729 VOUT.n41 VOUT.n40 9.3005
R2730 VOUT.n39 VOUT.n38 9.3005
R2731 VOUT.n268 VOUT.n267 9.3005
R2732 VOUT.n253 VOUT.n252 9.3005
R2733 VOUT.n262 VOUT.n261 9.3005
R2734 VOUT.n260 VOUT.n259 9.3005
R2735 VOUT.n236 VOUT.n235 9.3005
R2736 VOUT.n239 VOUT.n238 9.3005
R2737 VOUT.n237 VOUT.n231 9.3005
R2738 VOUT.n244 VOUT.n230 9.3005
R2739 VOUT.n289 VOUT.n288 9.3005
R2740 VOUT.n274 VOUT.n273 9.3005
R2741 VOUT.n283 VOUT.n282 9.3005
R2742 VOUT.n281 VOUT.n280 9.3005
R2743 VOUT.n309 VOUT.n308 9.3005
R2744 VOUT.n13 VOUT.n12 9.3005
R2745 VOUT.n303 VOUT.n302 9.3005
R2746 VOUT.n301 VOUT.n300 9.3005
R2747 VOUT.n173 VOUT.n172 9.3005
R2748 VOUT.n149 VOUT.n148 9.3005
R2749 VOUT.n144 VOUT.n143 9.3005
R2750 VOUT.n155 VOUT.n154 9.3005
R2751 VOUT.n157 VOUT.n156 9.3005
R2752 VOUT.n140 VOUT.n139 9.3005
R2753 VOUT.n163 VOUT.n162 9.3005
R2754 VOUT.n165 VOUT.n164 9.3005
R2755 VOUT.n166 VOUT.n135 9.3005
R2756 VOUT.n131 VOUT.n130 9.3005
R2757 VOUT.n107 VOUT.n106 9.3005
R2758 VOUT.n102 VOUT.n101 9.3005
R2759 VOUT.n113 VOUT.n112 9.3005
R2760 VOUT.n115 VOUT.n114 9.3005
R2761 VOUT.n98 VOUT.n97 9.3005
R2762 VOUT.n121 VOUT.n120 9.3005
R2763 VOUT.n123 VOUT.n122 9.3005
R2764 VOUT.n124 VOUT.n93 9.3005
R2765 VOUT.n205 VOUT.n204 8.92171
R2766 VOUT.n53 VOUT.n24 8.92171
R2767 VOUT.n154 VOUT.n153 8.92171
R2768 VOUT.n112 VOUT.n111 8.92171
R2769 VOUT.n91 VGP 8.234
R2770 VOUT.n201 VOUT.n195 8.14595
R2771 VOUT.n54 VOUT.n22 8.14595
R2772 VOUT.n150 VOUT.n144 8.14595
R2773 VOUT.n108 VOUT.n102 8.14595
R2774 VOUT.n77 VOUT.n76 8.03383
R2775 VOUT.n75 VOUT.n72 8.03383
R2776 VOUT.n87 VOUT.n86 8.03383
R2777 VOUT.n85 VOUT.n82 8.03383
R2778 VOUT.n68 VOUT.n67 8.03383
R2779 VOUT.n66 VOUT.n63 8.03383
R2780 VOUT.n6 VOUT.n5 8.03383
R2781 VOUT.n4 VOUT.n1 8.03383
R2782 VOUT.n90 VOUT.n80 7.77843
R2783 VOUT.n200 VOUT.n197 7.3702
R2784 VOUT.n58 VOUT.n57 7.3702
R2785 VOUT.n149 VOUT.n146 7.3702
R2786 VOUT.n107 VOUT.n104 7.3702
R2787 VOUT.n9 VGN 6.71885
R2788 VOUT.n201 VOUT.n200 5.81868
R2789 VOUT.n57 VOUT.n22 5.81868
R2790 VOUT.n150 VOUT.n149 5.81868
R2791 VOUT.n108 VOUT.n107 5.81868
R2792 VOUT.n175 VOUT.n18 5.06539
R2793 VOUT.n292 VOUT.n291 5.06539
R2794 VOUT.n204 VOUT.n195 5.04292
R2795 VOUT.n54 VOUT.n53 5.04292
R2796 VOUT.n153 VOUT.n144 5.04292
R2797 VOUT.n111 VOUT.n102 5.04292
R2798 VOUT.n249 VOUT.t10 4.9505
R2799 VOUT.n249 VOUT.t12 4.9505
R2800 VOUT.t12 VOUT.n248 4.9505
R2801 VOUT.n248 VOUT.t25 4.9505
R2802 VOUT.n247 VOUT.t8 4.9505
R2803 VOUT.t10 VOUT.n247 4.9505
R2804 VOUT.n295 VOUT.t6 4.9505
R2805 VOUT.n295 VOUT.t18 4.9505
R2806 VOUT.t16 VOUT.n297 4.9505
R2807 VOUT.n297 VOUT.t4 4.9505
R2808 VOUT.n294 VOUT.t4 4.9505
R2809 VOUT.t6 VOUT.n294 4.9505
R2810 VOUT.n80 VOUT.n79 4.9058
R2811 VOUT.n90 VOUT.n89 4.9058
R2812 VOUT.n227 VOUT.n226 4.88412
R2813 VOUT.n271 VOUT.n270 4.88412
R2814 VOUT.n133 VOUT.n91 4.84102
R2815 VIN VOUT.n9 4.83671
R2816 VOUT.n293 VOUT.n292 4.5005
R2817 VOUT.n180 VOUT.n18 4.5005
R2818 VOUT.n260 VOUT.n256 4.40546
R2819 VOUT.n246 VOUT.n230 4.40546
R2820 VOUT.n281 VOUT.n277 4.40546
R2821 VOUT.n301 VOUT.n16 4.40546
R2822 VOUT.n205 VOUT.n193 4.26717
R2823 VOUT.n50 VOUT.n24 4.26717
R2824 VOUT.n154 VOUT.n142 4.26717
R2825 VOUT.n112 VOUT.n100 4.26717
R2826 VOUT.n178 VOUT.t14 4.06363
R2827 VOUT.n178 VOUT.t30 4.06363
R2828 VOUT.t21 VOUT.n61 4.06363
R2829 VOUT.t23 VOUT.n61 4.06363
R2830 VOUT.n183 VOUT.t35 4.06363
R2831 VOUT.n183 VOUT.t28 4.06363
R2832 VOUT.n177 VOUT.t23 4.06363
R2833 VOUT.t14 VOUT.n177 4.06363
R2834 VOUT.t28 VOUT.n182 4.06363
R2835 VOUT.n182 VOUT.t1 4.06363
R2836 VOUT.n60 VOUT.t33 4.06363
R2837 VOUT.n60 VOUT.t35 4.06363
R2838 VOUT.n209 VOUT.n208 3.49141
R2839 VOUT.n49 VOUT.n26 3.49141
R2840 VOUT.n269 VOUT.n251 3.49141
R2841 VOUT.n234 VOUT.n228 3.49141
R2842 VOUT.n290 VOUT.n272 3.49141
R2843 VOUT.n310 VOUT.n11 3.49141
R2844 VOUT.n158 VOUT.n157 3.49141
R2845 VOUT.n116 VOUT.n115 3.49141
R2846 VOUT.n227 VOUT.n18 3.0853
R2847 VOUT.n212 VOUT.n191 2.71565
R2848 VOUT.n46 VOUT.n45 2.71565
R2849 VOUT.n267 VOUT.n266 2.71565
R2850 VOUT.n235 VOUT.n233 2.71565
R2851 VOUT.n288 VOUT.n287 2.71565
R2852 VOUT.n308 VOUT.n307 2.71565
R2853 VOUT.n161 VOUT.n140 2.71565
R2854 VOUT.n119 VOUT.n98 2.71565
R2855 VOUT.n199 VOUT.n198 2.4129
R2856 VOUT.n56 VOUT.n20 2.4129
R2857 VOUT.n148 VOUT.n147 2.4129
R2858 VOUT.n106 VOUT.n105 2.4129
R2859 VOUT.n213 VOUT.n189 1.93989
R2860 VOUT.n42 VOUT.n28 1.93989
R2861 VOUT.n263 VOUT.n253 1.93989
R2862 VOUT.n240 VOUT.n239 1.93989
R2863 VOUT.n284 VOUT.n274 1.93989
R2864 VOUT.n304 VOUT.n13 1.93989
R2865 VOUT.n162 VOUT.n138 1.93989
R2866 VOUT.n120 VOUT.n96 1.93989
R2867 VOUT.n292 VOUT.n271 1.80325
R2868 VOUT.n271 VOUT.n227 1.68416
R2869 VOUT.n218 VOUT.n216 1.16414
R2870 VOUT.n225 VOUT.n185 1.16414
R2871 VOUT.n41 VOUT.n30 1.16414
R2872 VOUT.n34 VOUT.n19 1.16414
R2873 VOUT.n262 VOUT.n255 1.16414
R2874 VOUT.n243 VOUT.n231 1.16414
R2875 VOUT.n283 VOUT.n276 1.16414
R2876 VOUT.n303 VOUT.n15 1.16414
R2877 VOUT.n167 VOUT.n165 1.16414
R2878 VOUT.n174 VOUT.n134 1.16414
R2879 VOUT.n125 VOUT.n123 1.16414
R2880 VOUT.n132 VOUT.n92 1.16414
R2881 VOUT.n296 VOUT.n293 0.603948
R2882 VOUT.n226 VOUT.n184 0.526362
R2883 VOUT.n270 VOUT.n250 0.526362
R2884 VOUT.n176 VOUT.n133 0.526362
R2885 VOUT.n176 VOUT.n175 0.526362
R2886 VOUT.n311 VOUT.n10 0.526362
R2887 VOUT.n291 VOUT.n10 0.526362
R2888 VOUT.n217 VOUT.n187 0.388379
R2889 VOUT.n223 VOUT.n222 0.388379
R2890 VOUT.n38 VOUT.n37 0.388379
R2891 VOUT.n33 VOUT.n32 0.388379
R2892 VOUT.n259 VOUT.n258 0.388379
R2893 VOUT.n245 VOUT.n244 0.388379
R2894 VOUT.n280 VOUT.n279 0.388379
R2895 VOUT.n300 VOUT.n299 0.388379
R2896 VOUT.n166 VOUT.n136 0.388379
R2897 VOUT.n172 VOUT.n171 0.388379
R2898 VOUT.n124 VOUT.n94 0.388379
R2899 VOUT.n130 VOUT.n129 0.388379
R2900 VOUT VOUT.n179 0.384121
R2901 VOUT.n91 VOUT.n90 0.282952
R2902 VOUT.n80 VOUT.n9 0.282952
R2903 VOUT.n180 VOUT 0.220328
R2904 VOUT.n79 VOUT.n71 0.189894
R2905 VOUT.n74 VOUT.n71 0.189894
R2906 VOUT.n89 VOUT.n81 0.189894
R2907 VOUT.n84 VOUT.n81 0.189894
R2908 VOUT.n70 VOUT.n62 0.189894
R2909 VOUT.n65 VOUT.n62 0.189894
R2910 VOUT.n8 VOUT.n0 0.189894
R2911 VOUT.n3 VOUT.n0 0.189894
R2912 VOUT.n199 VOUT.n194 0.155672
R2913 VOUT.n206 VOUT.n194 0.155672
R2914 VOUT.n207 VOUT.n206 0.155672
R2915 VOUT.n207 VOUT.n190 0.155672
R2916 VOUT.n214 VOUT.n190 0.155672
R2917 VOUT.n215 VOUT.n214 0.155672
R2918 VOUT.n215 VOUT.n186 0.155672
R2919 VOUT.n224 VOUT.n186 0.155672
R2920 VOUT.n56 VOUT.n55 0.155672
R2921 VOUT.n55 VOUT.n23 0.155672
R2922 VOUT.n48 VOUT.n23 0.155672
R2923 VOUT.n48 VOUT.n47 0.155672
R2924 VOUT.n47 VOUT.n27 0.155672
R2925 VOUT.n40 VOUT.n27 0.155672
R2926 VOUT.n40 VOUT.n39 0.155672
R2927 VOUT.n39 VOUT.n31 0.155672
R2928 VOUT.n268 VOUT.n252 0.155672
R2929 VOUT.n261 VOUT.n252 0.155672
R2930 VOUT.n261 VOUT.n260 0.155672
R2931 VOUT.n238 VOUT.n236 0.155672
R2932 VOUT.n238 VOUT.n237 0.155672
R2933 VOUT.n237 VOUT.n230 0.155672
R2934 VOUT.n289 VOUT.n273 0.155672
R2935 VOUT.n282 VOUT.n273 0.155672
R2936 VOUT.n282 VOUT.n281 0.155672
R2937 VOUT.n309 VOUT.n12 0.155672
R2938 VOUT.n302 VOUT.n12 0.155672
R2939 VOUT.n302 VOUT.n301 0.155672
R2940 VOUT.n148 VOUT.n143 0.155672
R2941 VOUT.n155 VOUT.n143 0.155672
R2942 VOUT.n156 VOUT.n155 0.155672
R2943 VOUT.n156 VOUT.n139 0.155672
R2944 VOUT.n163 VOUT.n139 0.155672
R2945 VOUT.n164 VOUT.n163 0.155672
R2946 VOUT.n164 VOUT.n135 0.155672
R2947 VOUT.n173 VOUT.n135 0.155672
R2948 VOUT.n106 VOUT.n101 0.155672
R2949 VOUT.n113 VOUT.n101 0.155672
R2950 VOUT.n114 VOUT.n113 0.155672
R2951 VOUT.n114 VOUT.n97 0.155672
R2952 VOUT.n121 VOUT.n97 0.155672
R2953 VOUT.n122 VOUT.n121 0.155672
R2954 VOUT.n122 VOUT.n93 0.155672
R2955 VOUT.n131 VOUT.n93 0.155672
R2956 VGP VOUT.n70 0.0648939
R2957 VGN VOUT.n8 0.0648939
R2958 VIN VOUT.n311 0.00481034
C0 VCC VOUT 7.274621f
C1 VOUT VSS 7.721633f
C2 VGP VSS 0.041624f
C3 VGN VSS 0.026573f
C4 VIN VSS 0.013276f
C5 VCC VSS 27.592247f
C6 VOUT.n0 VSS 0.010064f
C7 VOUT.t15 VSS 0.033218f
C8 VOUT.t3 VSS 0.032379f
C9 VOUT.t5 VSS 0.032379f
C10 VOUT.n1 VSS 0.017055f
C11 VOUT.t17 VSS 0.033218f
C12 VOUT.n2 VSS 0.019908f
C13 VOUT.n3 VSS 0.020799f
C14 VOUT.n4 VSS 0.00368f
C15 VOUT.n5 VSS 0.00368f
C16 VOUT.n6 VSS 0.017055f
C17 VOUT.n7 VSS 0.019896f
C18 VOUT.n8 VSS 0.008017f
C19 VOUT.n9 VSS 0.070498f
C20 VOUT.n10 VSS 0.04693f
C21 VOUT.n11 VSS 0.005624f
C22 VOUT.n12 VSS 0.003926f
C23 VOUT.n13 VSS 0.00211f
C24 VOUT.n14 VSS 0.004987f
C25 VOUT.n15 VSS 0.002234f
C26 VOUT.n16 VSS 0.015191f
C27 VOUT.t4 VSS 0.02482f
C28 VOUT.n17 VSS 0.152818f
C29 VOUT.n18 VSS 0.084312f
C30 VOUT.n19 VSS 0.006123f
C31 VOUT.t35 VSS 0.049641f
C32 VOUT.n20 VSS 0.023837f
C33 VOUT.n21 VSS 0.004987f
C34 VOUT.n22 VSS 0.002234f
C35 VOUT.n23 VSS 0.003926f
C36 VOUT.n24 VSS 0.00211f
C37 VOUT.n25 VSS 0.004987f
C38 VOUT.n26 VSS 0.002234f
C39 VOUT.n27 VSS 0.003926f
C40 VOUT.n28 VSS 0.00211f
C41 VOUT.n29 VSS 0.004987f
C42 VOUT.n30 VSS 0.002234f
C43 VOUT.n31 VSS 0.010148f
C44 VOUT.n32 VSS 0.002172f
C45 VOUT.n33 VSS 0.00211f
C46 VOUT.n34 VSS 0.004231f
C47 VOUT.n35 VSS 0.011789f
C48 VOUT.n36 VSS 0.004987f
C49 VOUT.n37 VSS 0.002172f
C50 VOUT.n38 VSS 0.00211f
C51 VOUT.n39 VSS 0.003926f
C52 VOUT.n40 VSS 0.003926f
C53 VOUT.n41 VSS 0.00211f
C54 VOUT.n42 VSS 0.002234f
C55 VOUT.n43 VSS 0.004987f
C56 VOUT.n44 VSS 0.004987f
C57 VOUT.n45 VSS 0.002234f
C58 VOUT.n46 VSS 0.00211f
C59 VOUT.n47 VSS 0.003926f
C60 VOUT.n48 VSS 0.003926f
C61 VOUT.n49 VSS 0.00211f
C62 VOUT.n50 VSS 0.002234f
C63 VOUT.n51 VSS 0.004987f
C64 VOUT.n52 VSS 0.004987f
C65 VOUT.n53 VSS 0.002234f
C66 VOUT.n54 VSS 0.00211f
C67 VOUT.n55 VSS 0.003926f
C68 VOUT.n56 VSS 0.124053f
C69 VOUT.n57 VSS 0.00211f
C70 VOUT.n58 VSS 0.003751f
C71 VOUT.n59 VSS 0.00374f
C72 VOUT.t33 VSS 0.035534f
C73 VOUT.n60 VSS 0.180778f
C74 VOUT.n61 VSS 0.180778f
C75 VOUT.t23 VSS 0.049641f
C76 VOUT.n62 VSS 0.010064f
C77 VOUT.t20 VSS 0.064765f
C78 VOUT.t22 VSS 0.063969f
C79 VOUT.t13 VSS 0.063969f
C80 VOUT.n63 VSS 0.027584f
C81 VOUT.t29 VSS 0.064765f
C82 VOUT.n64 VSS 0.030481f
C83 VOUT.n65 VSS 0.020799f
C84 VOUT.n66 VSS 0.00368f
C85 VOUT.n67 VSS 0.00368f
C86 VOUT.n68 VSS 0.027584f
C87 VOUT.n69 VSS 0.030468f
C88 VOUT.n70 VSS 0.008017f
C89 VOUT.n71 VSS 0.010064f
C90 VOUT.t7 VSS 0.033218f
C91 VOUT.t9 VSS 0.032379f
C92 VOUT.t11 VSS 0.032379f
C93 VOUT.n72 VSS 0.017055f
C94 VOUT.t24 VSS 0.033218f
C95 VOUT.n73 VSS 0.019908f
C96 VOUT.n74 VSS 0.020799f
C97 VOUT.n75 VSS 0.00368f
C98 VOUT.n76 VSS 0.00368f
C99 VOUT.n77 VSS 0.017055f
C100 VOUT.n78 VSS 0.019896f
C101 VOUT.n79 VSS 0.024202f
C102 VOUT.n80 VSS 0.112919f
C103 VOUT.n81 VSS 0.010064f
C104 VOUT.t32 VSS 0.064765f
C105 VOUT.t34 VSS 0.063969f
C106 VOUT.t27 VSS 0.063969f
C107 VOUT.n82 VSS 0.027584f
C108 VOUT.t0 VSS 0.064765f
C109 VOUT.n83 VSS 0.030481f
C110 VOUT.n84 VSS 0.020799f
C111 VOUT.n85 VSS 0.00368f
C112 VOUT.n86 VSS 0.00368f
C113 VOUT.n87 VSS 0.027584f
C114 VOUT.n88 VSS 0.030468f
C115 VOUT.n89 VSS 0.024202f
C116 VOUT.n90 VSS 0.112919f
C117 VOUT.n91 VSS 0.105099f
C118 VOUT.n92 VSS 0.004231f
C119 VOUT.n93 VSS 0.003926f
C120 VOUT.n94 VSS 0.002172f
C121 VOUT.n95 VSS 0.004987f
C122 VOUT.n96 VSS 0.002234f
C123 VOUT.n97 VSS 0.003926f
C124 VOUT.n98 VSS 0.00211f
C125 VOUT.n99 VSS 0.004987f
C126 VOUT.n100 VSS 0.002234f
C127 VOUT.n101 VSS 0.003926f
C128 VOUT.n102 VSS 0.00211f
C129 VOUT.n103 VSS 0.00374f
C130 VOUT.n104 VSS 0.003751f
C131 VOUT.t21 VSS 0.035534f
C132 VOUT.n105 VSS 0.023837f
C133 VOUT.n106 VSS 0.124053f
C134 VOUT.n107 VSS 0.00211f
C135 VOUT.n108 VSS 0.002234f
C136 VOUT.n109 VSS 0.004987f
C137 VOUT.n110 VSS 0.004987f
C138 VOUT.n111 VSS 0.002234f
C139 VOUT.n112 VSS 0.00211f
C140 VOUT.n113 VSS 0.003926f
C141 VOUT.n114 VSS 0.003926f
C142 VOUT.n115 VSS 0.00211f
C143 VOUT.n116 VSS 0.002234f
C144 VOUT.n117 VSS 0.004987f
C145 VOUT.n118 VSS 0.004987f
C146 VOUT.n119 VSS 0.002234f
C147 VOUT.n120 VSS 0.00211f
C148 VOUT.n121 VSS 0.003926f
C149 VOUT.n122 VSS 0.003926f
C150 VOUT.n123 VSS 0.00211f
C151 VOUT.n124 VSS 0.00211f
C152 VOUT.n125 VSS 0.002234f
C153 VOUT.n126 VSS 0.004987f
C154 VOUT.n127 VSS 0.004987f
C155 VOUT.n128 VSS 0.011789f
C156 VOUT.n129 VSS 0.002172f
C157 VOUT.n130 VSS 0.00211f
C158 VOUT.n131 VSS 0.010148f
C159 VOUT.n132 VSS 0.005948f
C160 VOUT.n133 VSS 0.023932f
C161 VOUT.n134 VSS 0.004231f
C162 VOUT.n135 VSS 0.003926f
C163 VOUT.n136 VSS 0.002172f
C164 VOUT.n137 VSS 0.004987f
C165 VOUT.n138 VSS 0.002234f
C166 VOUT.n139 VSS 0.003926f
C167 VOUT.n140 VSS 0.00211f
C168 VOUT.n141 VSS 0.004987f
C169 VOUT.n142 VSS 0.002234f
C170 VOUT.n143 VSS 0.003926f
C171 VOUT.n144 VSS 0.00211f
C172 VOUT.n145 VSS 0.00374f
C173 VOUT.n146 VSS 0.003751f
C174 VOUT.t31 VSS 0.010713f
C175 VOUT.n147 VSS 0.023837f
C176 VOUT.n148 VSS 0.124053f
C177 VOUT.n149 VSS 0.00211f
C178 VOUT.n150 VSS 0.002234f
C179 VOUT.n151 VSS 0.004987f
C180 VOUT.n152 VSS 0.004987f
C181 VOUT.n153 VSS 0.002234f
C182 VOUT.n154 VSS 0.00211f
C183 VOUT.n155 VSS 0.003926f
C184 VOUT.n156 VSS 0.003926f
C185 VOUT.n157 VSS 0.00211f
C186 VOUT.n158 VSS 0.002234f
C187 VOUT.n159 VSS 0.004987f
C188 VOUT.n160 VSS 0.004987f
C189 VOUT.n161 VSS 0.002234f
C190 VOUT.n162 VSS 0.00211f
C191 VOUT.n163 VSS 0.003926f
C192 VOUT.n164 VSS 0.003926f
C193 VOUT.n165 VSS 0.00211f
C194 VOUT.n166 VSS 0.00211f
C195 VOUT.n167 VSS 0.002234f
C196 VOUT.n168 VSS 0.004987f
C197 VOUT.n169 VSS 0.004987f
C198 VOUT.n170 VSS 0.011789f
C199 VOUT.n171 VSS 0.002172f
C200 VOUT.n172 VSS 0.00211f
C201 VOUT.n173 VSS 0.010148f
C202 VOUT.n174 VSS 0.005948f
C203 VOUT.n175 VSS 0.025204f
C204 VOUT.n176 VSS 0.089454f
C205 VOUT.n177 VSS 0.164674f
C206 VOUT.t14 VSS 0.049641f
C207 VOUT.t30 VSS 0.02482f
C208 VOUT.n178 VSS 0.180289f
C209 VOUT.n179 VSS 0.157643f
C210 VOUT.n180 VSS 0.088719f
C211 VOUT.n181 VSS 0.244326f
C212 VOUT.t1 VSS 0.02482f
C213 VOUT.n182 VSS 0.180289f
C214 VOUT.t28 VSS 0.049641f
C215 VOUT.n183 VSS 0.164674f
C216 VOUT.n184 VSS 0.101473f
C217 VOUT.n185 VSS 0.004231f
C218 VOUT.n186 VSS 0.003926f
C219 VOUT.n187 VSS 0.002172f
C220 VOUT.n188 VSS 0.004987f
C221 VOUT.n189 VSS 0.002234f
C222 VOUT.n190 VSS 0.003926f
C223 VOUT.n191 VSS 0.00211f
C224 VOUT.n192 VSS 0.004987f
C225 VOUT.n193 VSS 0.002234f
C226 VOUT.n194 VSS 0.003926f
C227 VOUT.n195 VSS 0.00211f
C228 VOUT.n196 VSS 0.00374f
C229 VOUT.n197 VSS 0.003751f
C230 VOUT.t2 VSS 0.010713f
C231 VOUT.n198 VSS 0.023837f
C232 VOUT.n199 VSS 0.124053f
C233 VOUT.n200 VSS 0.00211f
C234 VOUT.n201 VSS 0.002234f
C235 VOUT.n202 VSS 0.004987f
C236 VOUT.n203 VSS 0.004987f
C237 VOUT.n204 VSS 0.002234f
C238 VOUT.n205 VSS 0.00211f
C239 VOUT.n206 VSS 0.003926f
C240 VOUT.n207 VSS 0.003926f
C241 VOUT.n208 VSS 0.00211f
C242 VOUT.n209 VSS 0.002234f
C243 VOUT.n210 VSS 0.004987f
C244 VOUT.n211 VSS 0.004987f
C245 VOUT.n212 VSS 0.002234f
C246 VOUT.n213 VSS 0.00211f
C247 VOUT.n214 VSS 0.003926f
C248 VOUT.n215 VSS 0.003926f
C249 VOUT.n216 VSS 0.00211f
C250 VOUT.n217 VSS 0.00211f
C251 VOUT.n218 VSS 0.002234f
C252 VOUT.n219 VSS 0.004987f
C253 VOUT.n220 VSS 0.004987f
C254 VOUT.n221 VSS 0.011789f
C255 VOUT.n222 VSS 0.002172f
C256 VOUT.n223 VSS 0.00211f
C257 VOUT.n224 VSS 0.010148f
C258 VOUT.n225 VSS 0.005948f
C259 VOUT.n226 VSS 0.0249f
C260 VOUT.n227 VSS 0.095957f
C261 VOUT.n228 VSS 0.006367f
C262 VOUT.n229 VSS 0.00374f
C263 VOUT.n230 VSS 0.056882f
C264 VOUT.n231 VSS 0.00211f
C265 VOUT.n232 VSS 0.010983f
C266 VOUT.n233 VSS 0.002234f
C267 VOUT.n234 VSS 0.005624f
C268 VOUT.n235 VSS 0.00211f
C269 VOUT.n236 VSS 0.009933f
C270 VOUT.n237 VSS 0.003926f
C271 VOUT.n238 VSS 0.003926f
C272 VOUT.n239 VSS 0.00211f
C273 VOUT.n240 VSS 0.002234f
C274 VOUT.n241 VSS 0.004987f
C275 VOUT.n242 VSS 0.004987f
C276 VOUT.n243 VSS 0.002234f
C277 VOUT.n244 VSS 0.00211f
C278 VOUT.n245 VSS 0.002935f
C279 VOUT.n246 VSS 0.015191f
C280 VOUT.t8 VSS 0.020712f
C281 VOUT.n247 VSS 0.097748f
C282 VOUT.t10 VSS 0.02482f
C283 VOUT.t25 VSS 0.01241f
C284 VOUT.n248 VSS 0.097438f
C285 VOUT.t12 VSS 0.02482f
C286 VOUT.n249 VSS 0.089113f
C287 VOUT.n250 VSS 0.058826f
C288 VOUT.n251 VSS 0.005624f
C289 VOUT.n252 VSS 0.003926f
C290 VOUT.n253 VSS 0.00211f
C291 VOUT.n254 VSS 0.004987f
C292 VOUT.n255 VSS 0.002234f
C293 VOUT.n256 VSS 0.015191f
C294 VOUT.t26 VSS 0.008302f
C295 VOUT.n257 VSS 0.00374f
C296 VOUT.n258 VSS 0.002935f
C297 VOUT.n259 VSS 0.00211f
C298 VOUT.n260 VSS 0.056882f
C299 VOUT.n261 VSS 0.003926f
C300 VOUT.n262 VSS 0.00211f
C301 VOUT.n263 VSS 0.002234f
C302 VOUT.n264 VSS 0.004987f
C303 VOUT.n265 VSS 0.010983f
C304 VOUT.n266 VSS 0.002234f
C305 VOUT.n267 VSS 0.00211f
C306 VOUT.n268 VSS 0.009933f
C307 VOUT.n269 VSS 0.00619f
C308 VOUT.n270 VSS 0.024778f
C309 VOUT.n271 VSS 0.066624f
C310 VOUT.n272 VSS 0.005624f
C311 VOUT.n273 VSS 0.003926f
C312 VOUT.n274 VSS 0.00211f
C313 VOUT.n275 VSS 0.004987f
C314 VOUT.n276 VSS 0.002234f
C315 VOUT.n277 VSS 0.015191f
C316 VOUT.t19 VSS 0.008302f
C317 VOUT.n278 VSS 0.00374f
C318 VOUT.n279 VSS 0.002935f
C319 VOUT.n280 VSS 0.00211f
C320 VOUT.n281 VSS 0.056882f
C321 VOUT.n282 VSS 0.003926f
C322 VOUT.n283 VSS 0.00211f
C323 VOUT.n284 VSS 0.002234f
C324 VOUT.n285 VSS 0.004987f
C325 VOUT.n286 VSS 0.010983f
C326 VOUT.n287 VSS 0.002234f
C327 VOUT.n288 VSS 0.00211f
C328 VOUT.n289 VSS 0.009933f
C329 VOUT.n290 VSS 0.00619f
C330 VOUT.n291 VSS 0.025082f
C331 VOUT.n292 VSS 0.054979f
C332 VOUT.n293 VSS 0.071341f
C333 VOUT.n294 VSS 0.089113f
C334 VOUT.t6 VSS 0.02482f
C335 VOUT.t18 VSS 0.01241f
C336 VOUT.n295 VSS 0.097438f
C337 VOUT.n296 VSS 0.090235f
C338 VOUT.n297 VSS 0.097748f
C339 VOUT.t16 VSS 0.020712f
C340 VOUT.n298 VSS 0.00374f
C341 VOUT.n299 VSS 0.002935f
C342 VOUT.n300 VSS 0.00211f
C343 VOUT.n301 VSS 0.056882f
C344 VOUT.n302 VSS 0.003926f
C345 VOUT.n303 VSS 0.00211f
C346 VOUT.n304 VSS 0.002234f
C347 VOUT.n305 VSS 0.004987f
C348 VOUT.n306 VSS 0.010983f
C349 VOUT.n307 VSS 0.002234f
C350 VOUT.n308 VSS 0.00211f
C351 VOUT.n309 VSS 0.009933f
C352 VOUT.n310 VSS 0.00619f
C353 VOUT.n311 VSS 0.010546f
C354 VCC.n0 VSS 0.004728f
C355 VCC.n1 VSS 0.005247f
C356 VCC.n2 VSS 0.003806f
C357 VCC.n3 VSS 0.004728f
C358 VCC.n4 VSS 0.004728f
C359 VCC.n5 VSS 0.004728f
C360 VCC.n6 VSS 0.003806f
C361 VCC.n7 VSS 0.004728f
C362 VCC.n8 VSS 0.004728f
C363 VCC.n9 VSS 0.004728f
C364 VCC.n10 VSS 0.009074f
C365 VCC.n11 VSS 0.002813f
C366 VCC.n12 VSS 0.471215f
C367 VCC.t7 VSS 0.058173f
C368 VCC.t6 VSS 0.061135f
C369 VCC.t4 VSS 0.041042f
C370 VCC.n13 VSS 0.091499f
C371 VCC.n14 VSS 0.081839f
C372 VCC.n15 VSS 0.005699f
C373 VCC.n16 VSS 0.00201f
C374 VCC.n17 VSS 0.003215f
C375 VCC.n18 VSS 0.003215f
C376 VCC.n20 VSS 0.003215f
C377 VCC.n21 VSS 0.003215f
C378 VCC.n23 VSS 0.003215f
C379 VCC.n24 VSS 0.003215f
C380 VCC.n26 VSS 0.003215f
C381 VCC.n27 VSS 0.003215f
C382 VCC.n29 VSS 0.003215f
C383 VCC.n30 VSS 0.003215f
C384 VCC.n32 VSS 0.003215f
C385 VCC.n33 VSS 0.003215f
C386 VCC.n35 VSS 0.003215f
C387 VCC.n36 VSS 0.003215f
C388 VCC.n38 VSS 0.003215f
C389 VCC.t14 VSS 0.058173f
C390 VCC.t13 VSS 0.061135f
C391 VCC.t12 VSS 0.041042f
C392 VCC.n39 VSS 0.091499f
C393 VCC.n40 VSS 0.081839f
C394 VCC.n41 VSS 0.003215f
C395 VCC.n43 VSS 0.003215f
C396 VCC.n44 VSS 0.003215f
C397 VCC.n46 VSS 0.003215f
C398 VCC.n47 VSS 0.003215f
C399 VCC.n49 VSS 0.003215f
C400 VCC.n50 VSS 0.003215f
C401 VCC.n52 VSS 0.003215f
C402 VCC.n53 VSS 0.003215f
C403 VCC.n55 VSS 0.003215f
C404 VCC.n56 VSS 0.003215f
C405 VCC.n58 VSS 0.003215f
C406 VCC.n59 VSS 0.003215f
C407 VCC.n61 VSS 0.009074f
C408 VCC.n62 VSS 0.004728f
C409 VCC.n63 VSS 0.003806f
C410 VCC.n64 VSS 0.004728f
C411 VCC.n65 VSS 0.257615f
C412 VCC.n66 VSS 0.004728f
C413 VCC.n67 VSS 0.003806f
C414 VCC.n68 VSS 0.004728f
C415 VCC.n69 VSS 0.003806f
C416 VCC.n70 VSS 0.004728f
C417 VCC.t1 VSS 0.129455f
C418 VCC.n71 VSS 0.004728f
C419 VCC.n72 VSS 0.004728f
C420 VCC.n73 VSS 0.003806f
C421 VCC.t0 VSS 0.129455f
C422 VCC.n74 VSS 0.004728f
C423 VCC.n75 VSS 0.003806f
C424 VCC.n76 VSS 0.003806f
C425 VCC.n77 VSS 0.004728f
C426 VCC.n78 VSS 0.003806f
C427 VCC.n79 VSS 0.004728f
C428 VCC.n80 VSS 0.258909f
C429 VCC.n81 VSS 0.174764f
C430 VCC.n82 VSS 0.004728f
C431 VCC.n83 VSS 0.003806f
C432 VCC.n84 VSS 0.003806f
C433 VCC.n85 VSS 0.015285f
C434 VCC.n86 VSS 0.003159f
C435 VCC.n87 VSS 0.009074f
C436 VCC.t9 VSS 0.129455f
C437 VCC.n88 VSS 0.009074f
C438 VCC.n89 VSS 0.003159f
C439 VCC.n90 VSS 0.003215f
C440 VCC.n91 VSS 0.003215f
C441 VCC.n120 VSS 0.32752f
C442 VCC.n121 VSS 0.003215f
C443 VCC.n122 VSS 0.003215f
C444 VCC.t16 VSS 0.058173f
C445 VCC.t17 VSS 0.061135f
C446 VCC.t15 VSS 0.041042f
C447 VCC.n123 VSS 0.091499f
C448 VCC.n124 VSS 0.080621f
C449 VCC.t10 VSS 0.058173f
C450 VCC.t11 VSS 0.061135f
C451 VCC.t8 VSS 0.041042f
C452 VCC.n125 VSS 0.091499f
C453 VCC.n126 VSS 0.080621f
C454 VCC.n127 VSS 0.003215f
C455 VCC.n128 VSS 0.003215f
C456 VCC.n129 VSS 0.003215f
C457 VCC.n130 VSS 0.003215f
C458 VCC.n131 VSS 0.003215f
C459 VCC.n132 VSS 0.003215f
C460 VCC.n133 VSS 0.003215f
C461 VCC.n134 VSS 0.003215f
C462 VCC.n135 VSS 0.003215f
C463 VCC.n136 VSS 0.003215f
C464 VCC.n137 VSS 0.003215f
C465 VCC.n138 VSS 0.003215f
C466 VCC.n139 VSS 0.003215f
C467 VCC.n140 VSS 0.003215f
C468 VCC.n141 VSS 0.003215f
C469 VCC.n142 VSS 0.003215f
C470 VCC.n143 VSS 0.003215f
C471 VCC.n144 VSS 0.003215f
C472 VCC.n145 VSS 0.003215f
C473 VCC.n146 VSS 0.003215f
C474 VCC.n147 VSS 0.003215f
C475 VCC.n148 VSS 0.003215f
C476 VCC.n149 VSS 0.003215f
C477 VCC.n150 VSS 0.003215f
C478 VCC.n151 VSS 0.003215f
C479 VCC.n152 VSS 0.003215f
C480 VCC.n153 VSS 0.003215f
C481 VCC.n154 VSS 0.003215f
C482 VCC.n155 VSS 0.003215f
C483 VCC.n156 VSS 0.003215f
C484 VCC.n157 VSS 0.003215f
C485 VCC.n158 VSS 0.003215f
C486 VCC.n159 VSS 0.003215f
C487 VCC.n160 VSS 0.003215f
C488 VCC.n161 VSS 0.003215f
C489 VCC.n162 VSS 0.003215f
C490 VCC.n163 VSS 0.003215f
C491 VCC.n164 VSS 0.003215f
C492 VCC.n165 VSS 0.003215f
C493 VCC.n166 VSS 0.003215f
C494 VCC.n167 VSS 0.003215f
C495 VCC.n168 VSS 0.003215f
C496 VCC.n169 VSS 0.003215f
C497 VCC.n170 VSS 0.003215f
C498 VCC.n171 VSS 0.003215f
C499 VCC.n172 VSS 0.003215f
C500 VCC.n173 VSS 0.003215f
C501 VCC.n174 VSS 0.003215f
C502 VCC.n175 VSS 0.003215f
C503 VCC.n176 VSS 0.003215f
C504 VCC.n177 VSS 0.003215f
C505 VCC.n178 VSS 0.001726f
C506 VCC.n179 VSS 0.004481f
C507 VCC.n180 VSS 0.003097f
C508 VCC.n181 VSS 0.003215f
C509 VCC.n182 VSS 0.003215f
C510 VCC.n183 VSS 0.003215f
C511 VCC.n184 VSS 0.003215f
C512 VCC.n185 VSS 0.003215f
C513 VCC.n186 VSS 0.003215f
C514 VCC.n187 VSS 0.003215f
C515 VCC.n188 VSS 0.003215f
C516 VCC.n189 VSS 0.003215f
C517 VCC.n190 VSS 0.003215f
C518 VCC.n191 VSS 0.003215f
C519 VCC.n192 VSS 0.003215f
C520 VCC.n193 VSS 0.003215f
C521 VCC.n194 VSS 0.003215f
C522 VCC.n195 VSS 0.003215f
C523 VCC.n196 VSS 0.003215f
C524 VCC.n197 VSS 0.003215f
C525 VCC.n198 VSS 0.003215f
C526 VCC.n199 VSS 0.003215f
C527 VCC.n200 VSS 0.003215f
C528 VCC.n201 VSS 0.003215f
C529 VCC.n202 VSS 0.003215f
C530 VCC.n203 VSS 0.003215f
C531 VCC.n204 VSS 0.003215f
C532 VCC.n205 VSS 0.003215f
C533 VCC.n206 VSS 0.003215f
C534 VCC.n207 VSS 0.003215f
C535 VCC.n208 VSS 0.003215f
C536 VCC.n209 VSS 0.003215f
C537 VCC.n210 VSS 0.003215f
C538 VCC.n211 VSS 0.003215f
C539 VCC.n212 VSS 0.003215f
C540 VCC.n213 VSS 0.003215f
C541 VCC.n214 VSS 0.003215f
C542 VCC.n215 VSS 0.003215f
C543 VCC.n216 VSS 0.003215f
C544 VCC.n217 VSS 0.003215f
C545 VCC.n218 VSS 0.003215f
C546 VCC.n219 VSS 0.003215f
C547 VCC.n220 VSS 0.003215f
C548 VCC.n221 VSS 0.003215f
C549 VCC.n222 VSS 0.003215f
C550 VCC.n223 VSS 0.003215f
C551 VCC.n224 VSS 0.003215f
C552 VCC.n225 VSS 0.003215f
C553 VCC.n226 VSS 0.003215f
C554 VCC.n227 VSS 0.003215f
C555 VCC.n228 VSS 0.003215f
C556 VCC.n229 VSS 0.003215f
C557 VCC.n230 VSS 0.003215f
C558 VCC.n231 VSS 0.003215f
C559 VCC.n232 VSS 0.003215f
C560 VCC.n233 VSS 0.003215f
C561 VCC.n234 VSS 0.003215f
C562 VCC.n235 VSS 0.003215f
C563 VCC.n236 VSS 0.003215f
C564 VCC.n237 VSS 0.003215f
C565 VCC.n238 VSS 0.00201f
C566 VCC.n239 VSS 0.004481f
C567 VCC.n240 VSS 0.002813f
C568 VCC.n241 VSS 0.006465f
C569 VCC.n242 VSS 0.0088f
C570 VCC.n244 VSS 0.471215f
C571 VCC.n245 VSS 0.0088f
C572 VCC.n246 VSS 0.006465f
C573 VCC.n247 VSS 0.015285f
C574 VCC.n248 VSS 0.004728f
C575 VCC.n249 VSS 0.003806f
C576 VCC.n250 VSS 0.004728f
C577 VCC.n251 VSS 0.135927f
C578 VCC.n252 VSS 0.004728f
C579 VCC.n253 VSS 0.003806f
C580 VCC.n254 VSS 0.004728f
C581 VCC.n255 VSS 0.004728f
C582 VCC.n256 VSS 0.004728f
C583 VCC.n257 VSS 0.004728f
C584 VCC.n258 VSS 0.004728f
C585 VCC.n259 VSS 0.003806f
C586 VCC.n260 VSS 0.004728f
C587 VCC.n261 VSS 0.258909f
C588 VCC.n262 VSS 0.004728f
C589 VCC.n263 VSS 0.003806f
C590 VCC.n264 VSS 0.004728f
C591 VCC.n265 VSS 0.004728f
C592 VCC.n266 VSS 0.004728f
C593 VCC.n267 VSS 0.004728f
C594 VCC.n268 VSS 0.003806f
C595 VCC.n269 VSS 0.004728f
C596 VCC.n270 VSS 0.157935f
C597 VCC.n271 VSS 0.004728f
C598 VCC.n272 VSS 0.004728f
C599 VCC.n273 VSS 0.157935f
C600 VCC.t3 VSS 0.129455f
C601 VCC.n274 VSS 0.15664f
C602 VCC.t2 VSS 0.129455f
C603 VCC.n275 VSS 0.130749f
C604 VCC.n276 VSS 0.004728f
C605 VCC.n277 VSS 0.003806f
C606 VCC.n278 VSS 0.004728f
C607 VCC.n279 VSS 0.004728f
C608 VCC.n280 VSS 0.004728f
C609 VCC.n281 VSS 0.004728f
C610 VCC.n282 VSS 0.003806f
C611 VCC.n283 VSS 0.004728f
C612 VCC.n284 VSS 0.004728f
C613 VCC.n285 VSS 0.258909f
C614 VCC.n286 VSS 0.182531f
C615 VCC.t5 VSS 0.129455f
C616 VCC.n287 VSS 0.333993f
C617 VCC.n288 VSS 0.205833f
C618 VCC.n289 VSS 0.004728f
C619 VCC.n290 VSS 0.003806f
C620 VCC.n291 VSS 0.003159f
C621 VCC.n292 VSS 0.015285f
C622 VCC.n293 VSS 0.006465f
C623 VCC.n294 VSS 0.0088f
C624 VCC.n296 VSS 0.003215f
C625 VCC.n297 VSS 0.003215f
C626 VCC.n298 VSS 0.003215f
C627 VCC.n299 VSS 0.003215f
C628 VCC.n300 VSS 0.003215f
C629 VCC.n301 VSS 0.003215f
C630 VCC.n303 VSS 0.003215f
C631 VCC.n304 VSS 0.003215f
C632 VCC.n305 VSS 0.003215f
C633 VCC.n306 VSS 0.003215f
C634 VCC.n307 VSS 0.003215f
C635 VCC.n308 VSS 0.003215f
C636 VCC.n310 VSS 0.003215f
C637 VCC.n311 VSS 0.003215f
C638 VCC.n312 VSS 0.003215f
C639 VCC.n313 VSS 0.003215f
C640 VCC.n314 VSS 0.003215f
C641 VCC.n315 VSS 0.003215f
C642 VCC.n317 VSS 0.003215f
C643 VCC.n318 VSS 0.003215f
C644 VCC.n319 VSS 0.003215f
C645 VCC.n320 VSS 0.003215f
C646 VCC.n321 VSS 0.003215f
C647 VCC.n322 VSS 0.003215f
C648 VCC.n324 VSS 0.003215f
C649 VCC.n325 VSS 0.003215f
C650 VCC.n326 VSS 0.003215f
C651 VCC.n327 VSS 0.003215f
C652 VCC.n328 VSS 0.003215f
C653 VCC.n329 VSS 0.003215f
C654 VCC.n331 VSS 0.003215f
C655 VCC.n332 VSS 0.003215f
C656 VCC.n333 VSS 0.003215f
C657 VCC.n334 VSS 0.003215f
C658 VCC.n335 VSS 0.003215f
C659 VCC.n336 VSS 0.003215f
C660 VCC.n338 VSS 0.003215f
C661 VCC.n339 VSS 0.003215f
C662 VCC.n340 VSS 0.003215f
C663 VCC.n341 VSS 0.001726f
C664 VCC.n342 VSS 0.005699f
C665 VCC.n343 VSS 0.003097f
C666 VCC.n344 VSS 0.003215f
C667 VCC.n346 VSS 0.003215f
C668 VCC.n347 VSS 0.003215f
C669 VCC.n348 VSS 0.003215f
C670 VCC.n349 VSS 0.003215f
C671 VCC.n350 VSS 0.003215f
C672 VCC.n351 VSS 0.003215f
C673 VCC.n353 VSS 0.003215f
C674 VCC.n354 VSS 0.003215f
C675 VCC.n355 VSS 0.003215f
C676 VCC.n356 VSS 0.003215f
C677 VCC.n357 VSS 0.003215f
C678 VCC.n358 VSS 0.003215f
C679 VCC.n360 VSS 0.003215f
C680 VCC.n361 VSS 0.003215f
C681 VCC.n362 VSS 0.003215f
C682 VCC.n363 VSS 0.003215f
C683 VCC.n364 VSS 0.003215f
C684 VCC.n365 VSS 0.003215f
C685 VCC.n367 VSS 0.003215f
C686 VCC.n368 VSS 0.003215f
C687 VCC.n369 VSS 0.003215f
C688 VCC.n370 VSS 0.003215f
C689 VCC.n371 VSS 0.003215f
C690 VCC.n372 VSS 0.003215f
C691 VCC.n374 VSS 0.003215f
C692 VCC.n375 VSS 0.003215f
C693 VCC.n376 VSS 0.003215f
C694 VCC.n377 VSS 0.003215f
C695 VCC.n378 VSS 0.003215f
C696 VCC.n379 VSS 0.003215f
C697 VCC.n381 VSS 0.003215f
C698 VCC.n382 VSS 0.003215f
C699 VCC.n383 VSS 0.003215f
C700 VCC.n384 VSS 0.003215f
C701 VCC.n385 VSS 0.003215f
C702 VCC.n386 VSS 0.003215f
C703 VCC.n388 VSS 0.003215f
C704 VCC.n389 VSS 0.003215f
C705 VCC.n390 VSS 0.003215f
C706 VCC.n391 VSS 0.003215f
C707 VCC.n392 VSS 0.003215f
C708 VCC.n393 VSS 0.003215f
C709 VCC.n395 VSS 0.003215f
C710 VCC.n396 VSS 0.003215f
C711 VCC.n398 VSS 0.0088f
C712 VCC.n399 VSS 0.006465f
C713 VCC.n400 VSS 0.015285f
C714 VCC.n401 VSS 0.003159f
C715 VCC.n402 VSS 0.003806f
C716 VCC.n403 VSS 0.003806f
C717 VCC.n404 VSS 0.004728f
C718 VCC.n405 VSS 0.004728f
C719 VCC.n406 VSS 0.004728f
C720 VCC.n407 VSS 0.003806f
C721 VCC.n408 VSS 0.003806f
C722 VCC.n409 VSS 0.003806f
.ends

