* NGSPICE file created from diff_pair_sample_0352.ext - technology: sky130A

.subckt diff_pair_sample_0352 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t17 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=2.55255 ps=15.8 w=15.47 l=1.93
X1 B.t11 B.t9 B.t10 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=0 ps=0 w=15.47 l=1.93
X2 VDD2.t9 VN.t0 VTAIL.t2 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=2.55255 ps=15.8 w=15.47 l=1.93
X3 VTAIL.t16 VP.t1 VDD1.t8 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X4 VTAIL.t3 VN.t1 VDD2.t8 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X5 VDD1.t7 VP.t2 VTAIL.t18 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X6 VTAIL.t10 VP.t3 VDD1.t6 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X7 VDD1.t5 VP.t4 VTAIL.t14 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=6.0333 ps=31.72 w=15.47 l=1.93
X8 VDD2.t7 VN.t2 VTAIL.t0 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=6.0333 ps=31.72 w=15.47 l=1.93
X9 VTAIL.t7 VN.t3 VDD2.t6 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X10 VTAIL.t15 VP.t5 VDD1.t4 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X11 VDD2.t5 VN.t4 VTAIL.t4 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=2.55255 ps=15.8 w=15.47 l=1.93
X12 VDD1.t3 VP.t6 VTAIL.t19 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=6.0333 ps=31.72 w=15.47 l=1.93
X13 VDD2.t4 VN.t5 VTAIL.t5 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X14 VTAIL.t13 VP.t7 VDD1.t2 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X15 VDD1.t1 VP.t8 VTAIL.t11 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X16 VTAIL.t9 VN.t6 VDD2.t3 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X17 VDD1.t0 VP.t9 VTAIL.t12 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=2.55255 ps=15.8 w=15.47 l=1.93
X18 B.t8 B.t6 B.t7 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=0 ps=0 w=15.47 l=1.93
X19 VDD2.t2 VN.t7 VTAIL.t6 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=6.0333 ps=31.72 w=15.47 l=1.93
X20 B.t5 B.t3 B.t4 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=0 ps=0 w=15.47 l=1.93
X21 VDD2.t1 VN.t8 VTAIL.t1 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
X22 B.t2 B.t0 B.t1 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=6.0333 pd=31.72 as=0 ps=0 w=15.47 l=1.93
X23 VTAIL.t8 VN.t9 VDD2.t0 w_n3682_n4062# sky130_fd_pr__pfet_01v8 ad=2.55255 pd=15.8 as=2.55255 ps=15.8 w=15.47 l=1.93
R0 VP.n18 VP.t9 225.292
R1 VP.n60 VP.t2 193.175
R2 VP.n44 VP.t0 193.175
R3 VP.n7 VP.t1 193.175
R4 VP.n67 VP.t3 193.175
R5 VP.n75 VP.t6 193.175
R6 VP.n26 VP.t8 193.175
R7 VP.n41 VP.t4 193.175
R8 VP.n33 VP.t5 193.175
R9 VP.n17 VP.t7 193.175
R10 VP.n44 VP.n43 184.788
R11 VP.n76 VP.n75 184.788
R12 VP.n42 VP.n41 184.788
R13 VP.n20 VP.n19 161.3
R14 VP.n21 VP.n16 161.3
R15 VP.n23 VP.n22 161.3
R16 VP.n24 VP.n15 161.3
R17 VP.n26 VP.n25 161.3
R18 VP.n27 VP.n14 161.3
R19 VP.n29 VP.n28 161.3
R20 VP.n30 VP.n13 161.3
R21 VP.n32 VP.n31 161.3
R22 VP.n34 VP.n12 161.3
R23 VP.n36 VP.n35 161.3
R24 VP.n37 VP.n11 161.3
R25 VP.n39 VP.n38 161.3
R26 VP.n40 VP.n10 161.3
R27 VP.n74 VP.n0 161.3
R28 VP.n73 VP.n72 161.3
R29 VP.n71 VP.n1 161.3
R30 VP.n70 VP.n69 161.3
R31 VP.n68 VP.n2 161.3
R32 VP.n66 VP.n65 161.3
R33 VP.n64 VP.n3 161.3
R34 VP.n63 VP.n62 161.3
R35 VP.n61 VP.n4 161.3
R36 VP.n60 VP.n59 161.3
R37 VP.n58 VP.n5 161.3
R38 VP.n57 VP.n56 161.3
R39 VP.n55 VP.n6 161.3
R40 VP.n54 VP.n53 161.3
R41 VP.n52 VP.n51 161.3
R42 VP.n50 VP.n8 161.3
R43 VP.n49 VP.n48 161.3
R44 VP.n47 VP.n9 161.3
R45 VP.n46 VP.n45 161.3
R46 VP.n18 VP.n17 57.388
R47 VP.n56 VP.n55 53.1199
R48 VP.n62 VP.n3 53.1199
R49 VP.n28 VP.n13 53.1199
R50 VP.n22 VP.n21 53.1199
R51 VP.n43 VP.n42 51.9929
R52 VP.n50 VP.n49 51.1773
R53 VP.n69 VP.n1 51.1773
R54 VP.n35 VP.n11 51.1773
R55 VP.n49 VP.n9 29.8095
R56 VP.n73 VP.n1 29.8095
R57 VP.n39 VP.n11 29.8095
R58 VP.n56 VP.n5 27.8669
R59 VP.n62 VP.n61 27.8669
R60 VP.n28 VP.n27 27.8669
R61 VP.n22 VP.n15 27.8669
R62 VP.n45 VP.n9 24.4675
R63 VP.n51 VP.n50 24.4675
R64 VP.n55 VP.n54 24.4675
R65 VP.n60 VP.n5 24.4675
R66 VP.n61 VP.n60 24.4675
R67 VP.n66 VP.n3 24.4675
R68 VP.n69 VP.n68 24.4675
R69 VP.n74 VP.n73 24.4675
R70 VP.n40 VP.n39 24.4675
R71 VP.n32 VP.n13 24.4675
R72 VP.n35 VP.n34 24.4675
R73 VP.n26 VP.n15 24.4675
R74 VP.n27 VP.n26 24.4675
R75 VP.n21 VP.n20 24.4675
R76 VP.n54 VP.n7 12.7233
R77 VP.n67 VP.n66 12.7233
R78 VP.n33 VP.n32 12.7233
R79 VP.n20 VP.n17 12.7233
R80 VP.n19 VP.n18 12.5492
R81 VP.n51 VP.n7 11.7447
R82 VP.n68 VP.n67 11.7447
R83 VP.n34 VP.n33 11.7447
R84 VP.n45 VP.n44 0.97918
R85 VP.n75 VP.n74 0.97918
R86 VP.n41 VP.n40 0.97918
R87 VP.n19 VP.n16 0.189894
R88 VP.n23 VP.n16 0.189894
R89 VP.n24 VP.n23 0.189894
R90 VP.n25 VP.n24 0.189894
R91 VP.n25 VP.n14 0.189894
R92 VP.n29 VP.n14 0.189894
R93 VP.n30 VP.n29 0.189894
R94 VP.n31 VP.n30 0.189894
R95 VP.n31 VP.n12 0.189894
R96 VP.n36 VP.n12 0.189894
R97 VP.n37 VP.n36 0.189894
R98 VP.n38 VP.n37 0.189894
R99 VP.n38 VP.n10 0.189894
R100 VP.n42 VP.n10 0.189894
R101 VP.n46 VP.n43 0.189894
R102 VP.n47 VP.n46 0.189894
R103 VP.n48 VP.n47 0.189894
R104 VP.n48 VP.n8 0.189894
R105 VP.n52 VP.n8 0.189894
R106 VP.n53 VP.n52 0.189894
R107 VP.n53 VP.n6 0.189894
R108 VP.n57 VP.n6 0.189894
R109 VP.n58 VP.n57 0.189894
R110 VP.n59 VP.n58 0.189894
R111 VP.n59 VP.n4 0.189894
R112 VP.n63 VP.n4 0.189894
R113 VP.n64 VP.n63 0.189894
R114 VP.n65 VP.n64 0.189894
R115 VP.n65 VP.n2 0.189894
R116 VP.n70 VP.n2 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n72 VP.n71 0.189894
R119 VP.n72 VP.n0 0.189894
R120 VP.n76 VP.n0 0.189894
R121 VP VP.n76 0.0516364
R122 VTAIL.n352 VTAIL.n272 756.745
R123 VTAIL.n82 VTAIL.n2 756.745
R124 VTAIL.n266 VTAIL.n186 756.745
R125 VTAIL.n176 VTAIL.n96 756.745
R126 VTAIL.n301 VTAIL.n300 585
R127 VTAIL.n303 VTAIL.n302 585
R128 VTAIL.n296 VTAIL.n295 585
R129 VTAIL.n309 VTAIL.n308 585
R130 VTAIL.n311 VTAIL.n310 585
R131 VTAIL.n292 VTAIL.n291 585
R132 VTAIL.n317 VTAIL.n316 585
R133 VTAIL.n319 VTAIL.n318 585
R134 VTAIL.n288 VTAIL.n287 585
R135 VTAIL.n325 VTAIL.n324 585
R136 VTAIL.n327 VTAIL.n326 585
R137 VTAIL.n284 VTAIL.n283 585
R138 VTAIL.n333 VTAIL.n332 585
R139 VTAIL.n335 VTAIL.n334 585
R140 VTAIL.n280 VTAIL.n279 585
R141 VTAIL.n342 VTAIL.n341 585
R142 VTAIL.n343 VTAIL.n278 585
R143 VTAIL.n345 VTAIL.n344 585
R144 VTAIL.n276 VTAIL.n275 585
R145 VTAIL.n351 VTAIL.n350 585
R146 VTAIL.n353 VTAIL.n352 585
R147 VTAIL.n31 VTAIL.n30 585
R148 VTAIL.n33 VTAIL.n32 585
R149 VTAIL.n26 VTAIL.n25 585
R150 VTAIL.n39 VTAIL.n38 585
R151 VTAIL.n41 VTAIL.n40 585
R152 VTAIL.n22 VTAIL.n21 585
R153 VTAIL.n47 VTAIL.n46 585
R154 VTAIL.n49 VTAIL.n48 585
R155 VTAIL.n18 VTAIL.n17 585
R156 VTAIL.n55 VTAIL.n54 585
R157 VTAIL.n57 VTAIL.n56 585
R158 VTAIL.n14 VTAIL.n13 585
R159 VTAIL.n63 VTAIL.n62 585
R160 VTAIL.n65 VTAIL.n64 585
R161 VTAIL.n10 VTAIL.n9 585
R162 VTAIL.n72 VTAIL.n71 585
R163 VTAIL.n73 VTAIL.n8 585
R164 VTAIL.n75 VTAIL.n74 585
R165 VTAIL.n6 VTAIL.n5 585
R166 VTAIL.n81 VTAIL.n80 585
R167 VTAIL.n83 VTAIL.n82 585
R168 VTAIL.n267 VTAIL.n266 585
R169 VTAIL.n265 VTAIL.n264 585
R170 VTAIL.n190 VTAIL.n189 585
R171 VTAIL.n194 VTAIL.n192 585
R172 VTAIL.n259 VTAIL.n258 585
R173 VTAIL.n257 VTAIL.n256 585
R174 VTAIL.n196 VTAIL.n195 585
R175 VTAIL.n251 VTAIL.n250 585
R176 VTAIL.n249 VTAIL.n248 585
R177 VTAIL.n200 VTAIL.n199 585
R178 VTAIL.n243 VTAIL.n242 585
R179 VTAIL.n241 VTAIL.n240 585
R180 VTAIL.n204 VTAIL.n203 585
R181 VTAIL.n235 VTAIL.n234 585
R182 VTAIL.n233 VTAIL.n232 585
R183 VTAIL.n208 VTAIL.n207 585
R184 VTAIL.n227 VTAIL.n226 585
R185 VTAIL.n225 VTAIL.n224 585
R186 VTAIL.n212 VTAIL.n211 585
R187 VTAIL.n219 VTAIL.n218 585
R188 VTAIL.n217 VTAIL.n216 585
R189 VTAIL.n177 VTAIL.n176 585
R190 VTAIL.n175 VTAIL.n174 585
R191 VTAIL.n100 VTAIL.n99 585
R192 VTAIL.n104 VTAIL.n102 585
R193 VTAIL.n169 VTAIL.n168 585
R194 VTAIL.n167 VTAIL.n166 585
R195 VTAIL.n106 VTAIL.n105 585
R196 VTAIL.n161 VTAIL.n160 585
R197 VTAIL.n159 VTAIL.n158 585
R198 VTAIL.n110 VTAIL.n109 585
R199 VTAIL.n153 VTAIL.n152 585
R200 VTAIL.n151 VTAIL.n150 585
R201 VTAIL.n114 VTAIL.n113 585
R202 VTAIL.n145 VTAIL.n144 585
R203 VTAIL.n143 VTAIL.n142 585
R204 VTAIL.n118 VTAIL.n117 585
R205 VTAIL.n137 VTAIL.n136 585
R206 VTAIL.n135 VTAIL.n134 585
R207 VTAIL.n122 VTAIL.n121 585
R208 VTAIL.n129 VTAIL.n128 585
R209 VTAIL.n127 VTAIL.n126 585
R210 VTAIL.n299 VTAIL.t6 327.466
R211 VTAIL.n29 VTAIL.t19 327.466
R212 VTAIL.n215 VTAIL.t14 327.466
R213 VTAIL.n125 VTAIL.t0 327.466
R214 VTAIL.n302 VTAIL.n301 171.744
R215 VTAIL.n302 VTAIL.n295 171.744
R216 VTAIL.n309 VTAIL.n295 171.744
R217 VTAIL.n310 VTAIL.n309 171.744
R218 VTAIL.n310 VTAIL.n291 171.744
R219 VTAIL.n317 VTAIL.n291 171.744
R220 VTAIL.n318 VTAIL.n317 171.744
R221 VTAIL.n318 VTAIL.n287 171.744
R222 VTAIL.n325 VTAIL.n287 171.744
R223 VTAIL.n326 VTAIL.n325 171.744
R224 VTAIL.n326 VTAIL.n283 171.744
R225 VTAIL.n333 VTAIL.n283 171.744
R226 VTAIL.n334 VTAIL.n333 171.744
R227 VTAIL.n334 VTAIL.n279 171.744
R228 VTAIL.n342 VTAIL.n279 171.744
R229 VTAIL.n343 VTAIL.n342 171.744
R230 VTAIL.n344 VTAIL.n343 171.744
R231 VTAIL.n344 VTAIL.n275 171.744
R232 VTAIL.n351 VTAIL.n275 171.744
R233 VTAIL.n352 VTAIL.n351 171.744
R234 VTAIL.n32 VTAIL.n31 171.744
R235 VTAIL.n32 VTAIL.n25 171.744
R236 VTAIL.n39 VTAIL.n25 171.744
R237 VTAIL.n40 VTAIL.n39 171.744
R238 VTAIL.n40 VTAIL.n21 171.744
R239 VTAIL.n47 VTAIL.n21 171.744
R240 VTAIL.n48 VTAIL.n47 171.744
R241 VTAIL.n48 VTAIL.n17 171.744
R242 VTAIL.n55 VTAIL.n17 171.744
R243 VTAIL.n56 VTAIL.n55 171.744
R244 VTAIL.n56 VTAIL.n13 171.744
R245 VTAIL.n63 VTAIL.n13 171.744
R246 VTAIL.n64 VTAIL.n63 171.744
R247 VTAIL.n64 VTAIL.n9 171.744
R248 VTAIL.n72 VTAIL.n9 171.744
R249 VTAIL.n73 VTAIL.n72 171.744
R250 VTAIL.n74 VTAIL.n73 171.744
R251 VTAIL.n74 VTAIL.n5 171.744
R252 VTAIL.n81 VTAIL.n5 171.744
R253 VTAIL.n82 VTAIL.n81 171.744
R254 VTAIL.n266 VTAIL.n265 171.744
R255 VTAIL.n265 VTAIL.n189 171.744
R256 VTAIL.n194 VTAIL.n189 171.744
R257 VTAIL.n258 VTAIL.n194 171.744
R258 VTAIL.n258 VTAIL.n257 171.744
R259 VTAIL.n257 VTAIL.n195 171.744
R260 VTAIL.n250 VTAIL.n195 171.744
R261 VTAIL.n250 VTAIL.n249 171.744
R262 VTAIL.n249 VTAIL.n199 171.744
R263 VTAIL.n242 VTAIL.n199 171.744
R264 VTAIL.n242 VTAIL.n241 171.744
R265 VTAIL.n241 VTAIL.n203 171.744
R266 VTAIL.n234 VTAIL.n203 171.744
R267 VTAIL.n234 VTAIL.n233 171.744
R268 VTAIL.n233 VTAIL.n207 171.744
R269 VTAIL.n226 VTAIL.n207 171.744
R270 VTAIL.n226 VTAIL.n225 171.744
R271 VTAIL.n225 VTAIL.n211 171.744
R272 VTAIL.n218 VTAIL.n211 171.744
R273 VTAIL.n218 VTAIL.n217 171.744
R274 VTAIL.n176 VTAIL.n175 171.744
R275 VTAIL.n175 VTAIL.n99 171.744
R276 VTAIL.n104 VTAIL.n99 171.744
R277 VTAIL.n168 VTAIL.n104 171.744
R278 VTAIL.n168 VTAIL.n167 171.744
R279 VTAIL.n167 VTAIL.n105 171.744
R280 VTAIL.n160 VTAIL.n105 171.744
R281 VTAIL.n160 VTAIL.n159 171.744
R282 VTAIL.n159 VTAIL.n109 171.744
R283 VTAIL.n152 VTAIL.n109 171.744
R284 VTAIL.n152 VTAIL.n151 171.744
R285 VTAIL.n151 VTAIL.n113 171.744
R286 VTAIL.n144 VTAIL.n113 171.744
R287 VTAIL.n144 VTAIL.n143 171.744
R288 VTAIL.n143 VTAIL.n117 171.744
R289 VTAIL.n136 VTAIL.n117 171.744
R290 VTAIL.n136 VTAIL.n135 171.744
R291 VTAIL.n135 VTAIL.n121 171.744
R292 VTAIL.n128 VTAIL.n121 171.744
R293 VTAIL.n128 VTAIL.n127 171.744
R294 VTAIL.n301 VTAIL.t6 85.8723
R295 VTAIL.n31 VTAIL.t19 85.8723
R296 VTAIL.n217 VTAIL.t14 85.8723
R297 VTAIL.n127 VTAIL.t0 85.8723
R298 VTAIL.n185 VTAIL.n184 55.7127
R299 VTAIL.n183 VTAIL.n182 55.7127
R300 VTAIL.n95 VTAIL.n94 55.7127
R301 VTAIL.n93 VTAIL.n92 55.7127
R302 VTAIL.n359 VTAIL.n358 55.7125
R303 VTAIL.n1 VTAIL.n0 55.7125
R304 VTAIL.n89 VTAIL.n88 55.7125
R305 VTAIL.n91 VTAIL.n90 55.7125
R306 VTAIL.n357 VTAIL.n356 34.3187
R307 VTAIL.n87 VTAIL.n86 34.3187
R308 VTAIL.n271 VTAIL.n270 34.3187
R309 VTAIL.n181 VTAIL.n180 34.3187
R310 VTAIL.n93 VTAIL.n91 29.5996
R311 VTAIL.n357 VTAIL.n271 27.6514
R312 VTAIL.n300 VTAIL.n299 16.3895
R313 VTAIL.n30 VTAIL.n29 16.3895
R314 VTAIL.n216 VTAIL.n215 16.3895
R315 VTAIL.n126 VTAIL.n125 16.3895
R316 VTAIL.n345 VTAIL.n276 13.1884
R317 VTAIL.n75 VTAIL.n6 13.1884
R318 VTAIL.n192 VTAIL.n190 13.1884
R319 VTAIL.n102 VTAIL.n100 13.1884
R320 VTAIL.n303 VTAIL.n298 12.8005
R321 VTAIL.n346 VTAIL.n278 12.8005
R322 VTAIL.n350 VTAIL.n349 12.8005
R323 VTAIL.n33 VTAIL.n28 12.8005
R324 VTAIL.n76 VTAIL.n8 12.8005
R325 VTAIL.n80 VTAIL.n79 12.8005
R326 VTAIL.n264 VTAIL.n263 12.8005
R327 VTAIL.n260 VTAIL.n259 12.8005
R328 VTAIL.n219 VTAIL.n214 12.8005
R329 VTAIL.n174 VTAIL.n173 12.8005
R330 VTAIL.n170 VTAIL.n169 12.8005
R331 VTAIL.n129 VTAIL.n124 12.8005
R332 VTAIL.n304 VTAIL.n296 12.0247
R333 VTAIL.n341 VTAIL.n340 12.0247
R334 VTAIL.n353 VTAIL.n274 12.0247
R335 VTAIL.n34 VTAIL.n26 12.0247
R336 VTAIL.n71 VTAIL.n70 12.0247
R337 VTAIL.n83 VTAIL.n4 12.0247
R338 VTAIL.n267 VTAIL.n188 12.0247
R339 VTAIL.n256 VTAIL.n193 12.0247
R340 VTAIL.n220 VTAIL.n212 12.0247
R341 VTAIL.n177 VTAIL.n98 12.0247
R342 VTAIL.n166 VTAIL.n103 12.0247
R343 VTAIL.n130 VTAIL.n122 12.0247
R344 VTAIL.n308 VTAIL.n307 11.249
R345 VTAIL.n339 VTAIL.n280 11.249
R346 VTAIL.n354 VTAIL.n272 11.249
R347 VTAIL.n38 VTAIL.n37 11.249
R348 VTAIL.n69 VTAIL.n10 11.249
R349 VTAIL.n84 VTAIL.n2 11.249
R350 VTAIL.n268 VTAIL.n186 11.249
R351 VTAIL.n255 VTAIL.n196 11.249
R352 VTAIL.n224 VTAIL.n223 11.249
R353 VTAIL.n178 VTAIL.n96 11.249
R354 VTAIL.n165 VTAIL.n106 11.249
R355 VTAIL.n134 VTAIL.n133 11.249
R356 VTAIL.n311 VTAIL.n294 10.4732
R357 VTAIL.n336 VTAIL.n335 10.4732
R358 VTAIL.n41 VTAIL.n24 10.4732
R359 VTAIL.n66 VTAIL.n65 10.4732
R360 VTAIL.n252 VTAIL.n251 10.4732
R361 VTAIL.n227 VTAIL.n210 10.4732
R362 VTAIL.n162 VTAIL.n161 10.4732
R363 VTAIL.n137 VTAIL.n120 10.4732
R364 VTAIL.n312 VTAIL.n292 9.69747
R365 VTAIL.n332 VTAIL.n282 9.69747
R366 VTAIL.n42 VTAIL.n22 9.69747
R367 VTAIL.n62 VTAIL.n12 9.69747
R368 VTAIL.n248 VTAIL.n198 9.69747
R369 VTAIL.n228 VTAIL.n208 9.69747
R370 VTAIL.n158 VTAIL.n108 9.69747
R371 VTAIL.n138 VTAIL.n118 9.69747
R372 VTAIL.n356 VTAIL.n355 9.45567
R373 VTAIL.n86 VTAIL.n85 9.45567
R374 VTAIL.n270 VTAIL.n269 9.45567
R375 VTAIL.n180 VTAIL.n179 9.45567
R376 VTAIL.n355 VTAIL.n354 9.3005
R377 VTAIL.n274 VTAIL.n273 9.3005
R378 VTAIL.n349 VTAIL.n348 9.3005
R379 VTAIL.n321 VTAIL.n320 9.3005
R380 VTAIL.n290 VTAIL.n289 9.3005
R381 VTAIL.n315 VTAIL.n314 9.3005
R382 VTAIL.n313 VTAIL.n312 9.3005
R383 VTAIL.n294 VTAIL.n293 9.3005
R384 VTAIL.n307 VTAIL.n306 9.3005
R385 VTAIL.n305 VTAIL.n304 9.3005
R386 VTAIL.n298 VTAIL.n297 9.3005
R387 VTAIL.n323 VTAIL.n322 9.3005
R388 VTAIL.n286 VTAIL.n285 9.3005
R389 VTAIL.n329 VTAIL.n328 9.3005
R390 VTAIL.n331 VTAIL.n330 9.3005
R391 VTAIL.n282 VTAIL.n281 9.3005
R392 VTAIL.n337 VTAIL.n336 9.3005
R393 VTAIL.n339 VTAIL.n338 9.3005
R394 VTAIL.n340 VTAIL.n277 9.3005
R395 VTAIL.n347 VTAIL.n346 9.3005
R396 VTAIL.n85 VTAIL.n84 9.3005
R397 VTAIL.n4 VTAIL.n3 9.3005
R398 VTAIL.n79 VTAIL.n78 9.3005
R399 VTAIL.n51 VTAIL.n50 9.3005
R400 VTAIL.n20 VTAIL.n19 9.3005
R401 VTAIL.n45 VTAIL.n44 9.3005
R402 VTAIL.n43 VTAIL.n42 9.3005
R403 VTAIL.n24 VTAIL.n23 9.3005
R404 VTAIL.n37 VTAIL.n36 9.3005
R405 VTAIL.n35 VTAIL.n34 9.3005
R406 VTAIL.n28 VTAIL.n27 9.3005
R407 VTAIL.n53 VTAIL.n52 9.3005
R408 VTAIL.n16 VTAIL.n15 9.3005
R409 VTAIL.n59 VTAIL.n58 9.3005
R410 VTAIL.n61 VTAIL.n60 9.3005
R411 VTAIL.n12 VTAIL.n11 9.3005
R412 VTAIL.n67 VTAIL.n66 9.3005
R413 VTAIL.n69 VTAIL.n68 9.3005
R414 VTAIL.n70 VTAIL.n7 9.3005
R415 VTAIL.n77 VTAIL.n76 9.3005
R416 VTAIL.n202 VTAIL.n201 9.3005
R417 VTAIL.n245 VTAIL.n244 9.3005
R418 VTAIL.n247 VTAIL.n246 9.3005
R419 VTAIL.n198 VTAIL.n197 9.3005
R420 VTAIL.n253 VTAIL.n252 9.3005
R421 VTAIL.n255 VTAIL.n254 9.3005
R422 VTAIL.n193 VTAIL.n191 9.3005
R423 VTAIL.n261 VTAIL.n260 9.3005
R424 VTAIL.n269 VTAIL.n268 9.3005
R425 VTAIL.n188 VTAIL.n187 9.3005
R426 VTAIL.n263 VTAIL.n262 9.3005
R427 VTAIL.n239 VTAIL.n238 9.3005
R428 VTAIL.n237 VTAIL.n236 9.3005
R429 VTAIL.n206 VTAIL.n205 9.3005
R430 VTAIL.n231 VTAIL.n230 9.3005
R431 VTAIL.n229 VTAIL.n228 9.3005
R432 VTAIL.n210 VTAIL.n209 9.3005
R433 VTAIL.n223 VTAIL.n222 9.3005
R434 VTAIL.n221 VTAIL.n220 9.3005
R435 VTAIL.n214 VTAIL.n213 9.3005
R436 VTAIL.n112 VTAIL.n111 9.3005
R437 VTAIL.n155 VTAIL.n154 9.3005
R438 VTAIL.n157 VTAIL.n156 9.3005
R439 VTAIL.n108 VTAIL.n107 9.3005
R440 VTAIL.n163 VTAIL.n162 9.3005
R441 VTAIL.n165 VTAIL.n164 9.3005
R442 VTAIL.n103 VTAIL.n101 9.3005
R443 VTAIL.n171 VTAIL.n170 9.3005
R444 VTAIL.n179 VTAIL.n178 9.3005
R445 VTAIL.n98 VTAIL.n97 9.3005
R446 VTAIL.n173 VTAIL.n172 9.3005
R447 VTAIL.n149 VTAIL.n148 9.3005
R448 VTAIL.n147 VTAIL.n146 9.3005
R449 VTAIL.n116 VTAIL.n115 9.3005
R450 VTAIL.n141 VTAIL.n140 9.3005
R451 VTAIL.n139 VTAIL.n138 9.3005
R452 VTAIL.n120 VTAIL.n119 9.3005
R453 VTAIL.n133 VTAIL.n132 9.3005
R454 VTAIL.n131 VTAIL.n130 9.3005
R455 VTAIL.n124 VTAIL.n123 9.3005
R456 VTAIL.n316 VTAIL.n315 8.92171
R457 VTAIL.n331 VTAIL.n284 8.92171
R458 VTAIL.n46 VTAIL.n45 8.92171
R459 VTAIL.n61 VTAIL.n14 8.92171
R460 VTAIL.n247 VTAIL.n200 8.92171
R461 VTAIL.n232 VTAIL.n231 8.92171
R462 VTAIL.n157 VTAIL.n110 8.92171
R463 VTAIL.n142 VTAIL.n141 8.92171
R464 VTAIL.n319 VTAIL.n290 8.14595
R465 VTAIL.n328 VTAIL.n327 8.14595
R466 VTAIL.n49 VTAIL.n20 8.14595
R467 VTAIL.n58 VTAIL.n57 8.14595
R468 VTAIL.n244 VTAIL.n243 8.14595
R469 VTAIL.n235 VTAIL.n206 8.14595
R470 VTAIL.n154 VTAIL.n153 8.14595
R471 VTAIL.n145 VTAIL.n116 8.14595
R472 VTAIL.n320 VTAIL.n288 7.3702
R473 VTAIL.n324 VTAIL.n286 7.3702
R474 VTAIL.n50 VTAIL.n18 7.3702
R475 VTAIL.n54 VTAIL.n16 7.3702
R476 VTAIL.n240 VTAIL.n202 7.3702
R477 VTAIL.n236 VTAIL.n204 7.3702
R478 VTAIL.n150 VTAIL.n112 7.3702
R479 VTAIL.n146 VTAIL.n114 7.3702
R480 VTAIL.n323 VTAIL.n288 6.59444
R481 VTAIL.n324 VTAIL.n323 6.59444
R482 VTAIL.n53 VTAIL.n18 6.59444
R483 VTAIL.n54 VTAIL.n53 6.59444
R484 VTAIL.n240 VTAIL.n239 6.59444
R485 VTAIL.n239 VTAIL.n204 6.59444
R486 VTAIL.n150 VTAIL.n149 6.59444
R487 VTAIL.n149 VTAIL.n114 6.59444
R488 VTAIL.n320 VTAIL.n319 5.81868
R489 VTAIL.n327 VTAIL.n286 5.81868
R490 VTAIL.n50 VTAIL.n49 5.81868
R491 VTAIL.n57 VTAIL.n16 5.81868
R492 VTAIL.n243 VTAIL.n202 5.81868
R493 VTAIL.n236 VTAIL.n235 5.81868
R494 VTAIL.n153 VTAIL.n112 5.81868
R495 VTAIL.n146 VTAIL.n145 5.81868
R496 VTAIL.n316 VTAIL.n290 5.04292
R497 VTAIL.n328 VTAIL.n284 5.04292
R498 VTAIL.n46 VTAIL.n20 5.04292
R499 VTAIL.n58 VTAIL.n14 5.04292
R500 VTAIL.n244 VTAIL.n200 5.04292
R501 VTAIL.n232 VTAIL.n206 5.04292
R502 VTAIL.n154 VTAIL.n110 5.04292
R503 VTAIL.n142 VTAIL.n116 5.04292
R504 VTAIL.n315 VTAIL.n292 4.26717
R505 VTAIL.n332 VTAIL.n331 4.26717
R506 VTAIL.n45 VTAIL.n22 4.26717
R507 VTAIL.n62 VTAIL.n61 4.26717
R508 VTAIL.n248 VTAIL.n247 4.26717
R509 VTAIL.n231 VTAIL.n208 4.26717
R510 VTAIL.n158 VTAIL.n157 4.26717
R511 VTAIL.n141 VTAIL.n118 4.26717
R512 VTAIL.n299 VTAIL.n297 3.70982
R513 VTAIL.n29 VTAIL.n27 3.70982
R514 VTAIL.n215 VTAIL.n213 3.70982
R515 VTAIL.n125 VTAIL.n123 3.70982
R516 VTAIL.n312 VTAIL.n311 3.49141
R517 VTAIL.n335 VTAIL.n282 3.49141
R518 VTAIL.n42 VTAIL.n41 3.49141
R519 VTAIL.n65 VTAIL.n12 3.49141
R520 VTAIL.n251 VTAIL.n198 3.49141
R521 VTAIL.n228 VTAIL.n227 3.49141
R522 VTAIL.n161 VTAIL.n108 3.49141
R523 VTAIL.n138 VTAIL.n137 3.49141
R524 VTAIL.n308 VTAIL.n294 2.71565
R525 VTAIL.n336 VTAIL.n280 2.71565
R526 VTAIL.n356 VTAIL.n272 2.71565
R527 VTAIL.n38 VTAIL.n24 2.71565
R528 VTAIL.n66 VTAIL.n10 2.71565
R529 VTAIL.n86 VTAIL.n2 2.71565
R530 VTAIL.n270 VTAIL.n186 2.71565
R531 VTAIL.n252 VTAIL.n196 2.71565
R532 VTAIL.n224 VTAIL.n210 2.71565
R533 VTAIL.n180 VTAIL.n96 2.71565
R534 VTAIL.n162 VTAIL.n106 2.71565
R535 VTAIL.n134 VTAIL.n120 2.71565
R536 VTAIL.n358 VTAIL.t1 2.10166
R537 VTAIL.n358 VTAIL.t9 2.10166
R538 VTAIL.n0 VTAIL.t2 2.10166
R539 VTAIL.n0 VTAIL.t8 2.10166
R540 VTAIL.n88 VTAIL.t18 2.10166
R541 VTAIL.n88 VTAIL.t10 2.10166
R542 VTAIL.n90 VTAIL.t17 2.10166
R543 VTAIL.n90 VTAIL.t16 2.10166
R544 VTAIL.n184 VTAIL.t11 2.10166
R545 VTAIL.n184 VTAIL.t15 2.10166
R546 VTAIL.n182 VTAIL.t12 2.10166
R547 VTAIL.n182 VTAIL.t13 2.10166
R548 VTAIL.n94 VTAIL.t5 2.10166
R549 VTAIL.n94 VTAIL.t3 2.10166
R550 VTAIL.n92 VTAIL.t4 2.10166
R551 VTAIL.n92 VTAIL.t7 2.10166
R552 VTAIL.n95 VTAIL.n93 1.94878
R553 VTAIL.n181 VTAIL.n95 1.94878
R554 VTAIL.n185 VTAIL.n183 1.94878
R555 VTAIL.n271 VTAIL.n185 1.94878
R556 VTAIL.n91 VTAIL.n89 1.94878
R557 VTAIL.n89 VTAIL.n87 1.94878
R558 VTAIL.n359 VTAIL.n357 1.94878
R559 VTAIL.n307 VTAIL.n296 1.93989
R560 VTAIL.n341 VTAIL.n339 1.93989
R561 VTAIL.n354 VTAIL.n353 1.93989
R562 VTAIL.n37 VTAIL.n26 1.93989
R563 VTAIL.n71 VTAIL.n69 1.93989
R564 VTAIL.n84 VTAIL.n83 1.93989
R565 VTAIL.n268 VTAIL.n267 1.93989
R566 VTAIL.n256 VTAIL.n255 1.93989
R567 VTAIL.n223 VTAIL.n212 1.93989
R568 VTAIL.n178 VTAIL.n177 1.93989
R569 VTAIL.n166 VTAIL.n165 1.93989
R570 VTAIL.n133 VTAIL.n122 1.93989
R571 VTAIL VTAIL.n1 1.5199
R572 VTAIL.n183 VTAIL.n181 1.44447
R573 VTAIL.n87 VTAIL.n1 1.44447
R574 VTAIL.n304 VTAIL.n303 1.16414
R575 VTAIL.n340 VTAIL.n278 1.16414
R576 VTAIL.n350 VTAIL.n274 1.16414
R577 VTAIL.n34 VTAIL.n33 1.16414
R578 VTAIL.n70 VTAIL.n8 1.16414
R579 VTAIL.n80 VTAIL.n4 1.16414
R580 VTAIL.n264 VTAIL.n188 1.16414
R581 VTAIL.n259 VTAIL.n193 1.16414
R582 VTAIL.n220 VTAIL.n219 1.16414
R583 VTAIL.n174 VTAIL.n98 1.16414
R584 VTAIL.n169 VTAIL.n103 1.16414
R585 VTAIL.n130 VTAIL.n129 1.16414
R586 VTAIL VTAIL.n359 0.429379
R587 VTAIL.n300 VTAIL.n298 0.388379
R588 VTAIL.n346 VTAIL.n345 0.388379
R589 VTAIL.n349 VTAIL.n276 0.388379
R590 VTAIL.n30 VTAIL.n28 0.388379
R591 VTAIL.n76 VTAIL.n75 0.388379
R592 VTAIL.n79 VTAIL.n6 0.388379
R593 VTAIL.n263 VTAIL.n190 0.388379
R594 VTAIL.n260 VTAIL.n192 0.388379
R595 VTAIL.n216 VTAIL.n214 0.388379
R596 VTAIL.n173 VTAIL.n100 0.388379
R597 VTAIL.n170 VTAIL.n102 0.388379
R598 VTAIL.n126 VTAIL.n124 0.388379
R599 VTAIL.n305 VTAIL.n297 0.155672
R600 VTAIL.n306 VTAIL.n305 0.155672
R601 VTAIL.n306 VTAIL.n293 0.155672
R602 VTAIL.n313 VTAIL.n293 0.155672
R603 VTAIL.n314 VTAIL.n313 0.155672
R604 VTAIL.n314 VTAIL.n289 0.155672
R605 VTAIL.n321 VTAIL.n289 0.155672
R606 VTAIL.n322 VTAIL.n321 0.155672
R607 VTAIL.n322 VTAIL.n285 0.155672
R608 VTAIL.n329 VTAIL.n285 0.155672
R609 VTAIL.n330 VTAIL.n329 0.155672
R610 VTAIL.n330 VTAIL.n281 0.155672
R611 VTAIL.n337 VTAIL.n281 0.155672
R612 VTAIL.n338 VTAIL.n337 0.155672
R613 VTAIL.n338 VTAIL.n277 0.155672
R614 VTAIL.n347 VTAIL.n277 0.155672
R615 VTAIL.n348 VTAIL.n347 0.155672
R616 VTAIL.n348 VTAIL.n273 0.155672
R617 VTAIL.n355 VTAIL.n273 0.155672
R618 VTAIL.n35 VTAIL.n27 0.155672
R619 VTAIL.n36 VTAIL.n35 0.155672
R620 VTAIL.n36 VTAIL.n23 0.155672
R621 VTAIL.n43 VTAIL.n23 0.155672
R622 VTAIL.n44 VTAIL.n43 0.155672
R623 VTAIL.n44 VTAIL.n19 0.155672
R624 VTAIL.n51 VTAIL.n19 0.155672
R625 VTAIL.n52 VTAIL.n51 0.155672
R626 VTAIL.n52 VTAIL.n15 0.155672
R627 VTAIL.n59 VTAIL.n15 0.155672
R628 VTAIL.n60 VTAIL.n59 0.155672
R629 VTAIL.n60 VTAIL.n11 0.155672
R630 VTAIL.n67 VTAIL.n11 0.155672
R631 VTAIL.n68 VTAIL.n67 0.155672
R632 VTAIL.n68 VTAIL.n7 0.155672
R633 VTAIL.n77 VTAIL.n7 0.155672
R634 VTAIL.n78 VTAIL.n77 0.155672
R635 VTAIL.n78 VTAIL.n3 0.155672
R636 VTAIL.n85 VTAIL.n3 0.155672
R637 VTAIL.n269 VTAIL.n187 0.155672
R638 VTAIL.n262 VTAIL.n187 0.155672
R639 VTAIL.n262 VTAIL.n261 0.155672
R640 VTAIL.n261 VTAIL.n191 0.155672
R641 VTAIL.n254 VTAIL.n191 0.155672
R642 VTAIL.n254 VTAIL.n253 0.155672
R643 VTAIL.n253 VTAIL.n197 0.155672
R644 VTAIL.n246 VTAIL.n197 0.155672
R645 VTAIL.n246 VTAIL.n245 0.155672
R646 VTAIL.n245 VTAIL.n201 0.155672
R647 VTAIL.n238 VTAIL.n201 0.155672
R648 VTAIL.n238 VTAIL.n237 0.155672
R649 VTAIL.n237 VTAIL.n205 0.155672
R650 VTAIL.n230 VTAIL.n205 0.155672
R651 VTAIL.n230 VTAIL.n229 0.155672
R652 VTAIL.n229 VTAIL.n209 0.155672
R653 VTAIL.n222 VTAIL.n209 0.155672
R654 VTAIL.n222 VTAIL.n221 0.155672
R655 VTAIL.n221 VTAIL.n213 0.155672
R656 VTAIL.n179 VTAIL.n97 0.155672
R657 VTAIL.n172 VTAIL.n97 0.155672
R658 VTAIL.n172 VTAIL.n171 0.155672
R659 VTAIL.n171 VTAIL.n101 0.155672
R660 VTAIL.n164 VTAIL.n101 0.155672
R661 VTAIL.n164 VTAIL.n163 0.155672
R662 VTAIL.n163 VTAIL.n107 0.155672
R663 VTAIL.n156 VTAIL.n107 0.155672
R664 VTAIL.n156 VTAIL.n155 0.155672
R665 VTAIL.n155 VTAIL.n111 0.155672
R666 VTAIL.n148 VTAIL.n111 0.155672
R667 VTAIL.n148 VTAIL.n147 0.155672
R668 VTAIL.n147 VTAIL.n115 0.155672
R669 VTAIL.n140 VTAIL.n115 0.155672
R670 VTAIL.n140 VTAIL.n139 0.155672
R671 VTAIL.n139 VTAIL.n119 0.155672
R672 VTAIL.n132 VTAIL.n119 0.155672
R673 VTAIL.n132 VTAIL.n131 0.155672
R674 VTAIL.n131 VTAIL.n123 0.155672
R675 VDD1.n80 VDD1.n0 756.745
R676 VDD1.n167 VDD1.n87 756.745
R677 VDD1.n81 VDD1.n80 585
R678 VDD1.n79 VDD1.n78 585
R679 VDD1.n4 VDD1.n3 585
R680 VDD1.n8 VDD1.n6 585
R681 VDD1.n73 VDD1.n72 585
R682 VDD1.n71 VDD1.n70 585
R683 VDD1.n10 VDD1.n9 585
R684 VDD1.n65 VDD1.n64 585
R685 VDD1.n63 VDD1.n62 585
R686 VDD1.n14 VDD1.n13 585
R687 VDD1.n57 VDD1.n56 585
R688 VDD1.n55 VDD1.n54 585
R689 VDD1.n18 VDD1.n17 585
R690 VDD1.n49 VDD1.n48 585
R691 VDD1.n47 VDD1.n46 585
R692 VDD1.n22 VDD1.n21 585
R693 VDD1.n41 VDD1.n40 585
R694 VDD1.n39 VDD1.n38 585
R695 VDD1.n26 VDD1.n25 585
R696 VDD1.n33 VDD1.n32 585
R697 VDD1.n31 VDD1.n30 585
R698 VDD1.n116 VDD1.n115 585
R699 VDD1.n118 VDD1.n117 585
R700 VDD1.n111 VDD1.n110 585
R701 VDD1.n124 VDD1.n123 585
R702 VDD1.n126 VDD1.n125 585
R703 VDD1.n107 VDD1.n106 585
R704 VDD1.n132 VDD1.n131 585
R705 VDD1.n134 VDD1.n133 585
R706 VDD1.n103 VDD1.n102 585
R707 VDD1.n140 VDD1.n139 585
R708 VDD1.n142 VDD1.n141 585
R709 VDD1.n99 VDD1.n98 585
R710 VDD1.n148 VDD1.n147 585
R711 VDD1.n150 VDD1.n149 585
R712 VDD1.n95 VDD1.n94 585
R713 VDD1.n157 VDD1.n156 585
R714 VDD1.n158 VDD1.n93 585
R715 VDD1.n160 VDD1.n159 585
R716 VDD1.n91 VDD1.n90 585
R717 VDD1.n166 VDD1.n165 585
R718 VDD1.n168 VDD1.n167 585
R719 VDD1.n29 VDD1.t0 327.466
R720 VDD1.n114 VDD1.t9 327.466
R721 VDD1.n80 VDD1.n79 171.744
R722 VDD1.n79 VDD1.n3 171.744
R723 VDD1.n8 VDD1.n3 171.744
R724 VDD1.n72 VDD1.n8 171.744
R725 VDD1.n72 VDD1.n71 171.744
R726 VDD1.n71 VDD1.n9 171.744
R727 VDD1.n64 VDD1.n9 171.744
R728 VDD1.n64 VDD1.n63 171.744
R729 VDD1.n63 VDD1.n13 171.744
R730 VDD1.n56 VDD1.n13 171.744
R731 VDD1.n56 VDD1.n55 171.744
R732 VDD1.n55 VDD1.n17 171.744
R733 VDD1.n48 VDD1.n17 171.744
R734 VDD1.n48 VDD1.n47 171.744
R735 VDD1.n47 VDD1.n21 171.744
R736 VDD1.n40 VDD1.n21 171.744
R737 VDD1.n40 VDD1.n39 171.744
R738 VDD1.n39 VDD1.n25 171.744
R739 VDD1.n32 VDD1.n25 171.744
R740 VDD1.n32 VDD1.n31 171.744
R741 VDD1.n117 VDD1.n116 171.744
R742 VDD1.n117 VDD1.n110 171.744
R743 VDD1.n124 VDD1.n110 171.744
R744 VDD1.n125 VDD1.n124 171.744
R745 VDD1.n125 VDD1.n106 171.744
R746 VDD1.n132 VDD1.n106 171.744
R747 VDD1.n133 VDD1.n132 171.744
R748 VDD1.n133 VDD1.n102 171.744
R749 VDD1.n140 VDD1.n102 171.744
R750 VDD1.n141 VDD1.n140 171.744
R751 VDD1.n141 VDD1.n98 171.744
R752 VDD1.n148 VDD1.n98 171.744
R753 VDD1.n149 VDD1.n148 171.744
R754 VDD1.n149 VDD1.n94 171.744
R755 VDD1.n157 VDD1.n94 171.744
R756 VDD1.n158 VDD1.n157 171.744
R757 VDD1.n159 VDD1.n158 171.744
R758 VDD1.n159 VDD1.n90 171.744
R759 VDD1.n166 VDD1.n90 171.744
R760 VDD1.n167 VDD1.n166 171.744
R761 VDD1.n31 VDD1.t0 85.8723
R762 VDD1.n116 VDD1.t9 85.8723
R763 VDD1.n175 VDD1.n174 73.7972
R764 VDD1.n86 VDD1.n85 72.3915
R765 VDD1.n173 VDD1.n172 72.3913
R766 VDD1.n177 VDD1.n176 72.3913
R767 VDD1.n86 VDD1.n84 52.9457
R768 VDD1.n173 VDD1.n171 52.9457
R769 VDD1.n177 VDD1.n175 47.863
R770 VDD1.n30 VDD1.n29 16.3895
R771 VDD1.n115 VDD1.n114 16.3895
R772 VDD1.n6 VDD1.n4 13.1884
R773 VDD1.n160 VDD1.n91 13.1884
R774 VDD1.n78 VDD1.n77 12.8005
R775 VDD1.n74 VDD1.n73 12.8005
R776 VDD1.n33 VDD1.n28 12.8005
R777 VDD1.n118 VDD1.n113 12.8005
R778 VDD1.n161 VDD1.n93 12.8005
R779 VDD1.n165 VDD1.n164 12.8005
R780 VDD1.n81 VDD1.n2 12.0247
R781 VDD1.n70 VDD1.n7 12.0247
R782 VDD1.n34 VDD1.n26 12.0247
R783 VDD1.n119 VDD1.n111 12.0247
R784 VDD1.n156 VDD1.n155 12.0247
R785 VDD1.n168 VDD1.n89 12.0247
R786 VDD1.n82 VDD1.n0 11.249
R787 VDD1.n69 VDD1.n10 11.249
R788 VDD1.n38 VDD1.n37 11.249
R789 VDD1.n123 VDD1.n122 11.249
R790 VDD1.n154 VDD1.n95 11.249
R791 VDD1.n169 VDD1.n87 11.249
R792 VDD1.n66 VDD1.n65 10.4732
R793 VDD1.n41 VDD1.n24 10.4732
R794 VDD1.n126 VDD1.n109 10.4732
R795 VDD1.n151 VDD1.n150 10.4732
R796 VDD1.n62 VDD1.n12 9.69747
R797 VDD1.n42 VDD1.n22 9.69747
R798 VDD1.n127 VDD1.n107 9.69747
R799 VDD1.n147 VDD1.n97 9.69747
R800 VDD1.n84 VDD1.n83 9.45567
R801 VDD1.n171 VDD1.n170 9.45567
R802 VDD1.n16 VDD1.n15 9.3005
R803 VDD1.n59 VDD1.n58 9.3005
R804 VDD1.n61 VDD1.n60 9.3005
R805 VDD1.n12 VDD1.n11 9.3005
R806 VDD1.n67 VDD1.n66 9.3005
R807 VDD1.n69 VDD1.n68 9.3005
R808 VDD1.n7 VDD1.n5 9.3005
R809 VDD1.n75 VDD1.n74 9.3005
R810 VDD1.n83 VDD1.n82 9.3005
R811 VDD1.n2 VDD1.n1 9.3005
R812 VDD1.n77 VDD1.n76 9.3005
R813 VDD1.n53 VDD1.n52 9.3005
R814 VDD1.n51 VDD1.n50 9.3005
R815 VDD1.n20 VDD1.n19 9.3005
R816 VDD1.n45 VDD1.n44 9.3005
R817 VDD1.n43 VDD1.n42 9.3005
R818 VDD1.n24 VDD1.n23 9.3005
R819 VDD1.n37 VDD1.n36 9.3005
R820 VDD1.n35 VDD1.n34 9.3005
R821 VDD1.n28 VDD1.n27 9.3005
R822 VDD1.n170 VDD1.n169 9.3005
R823 VDD1.n89 VDD1.n88 9.3005
R824 VDD1.n164 VDD1.n163 9.3005
R825 VDD1.n136 VDD1.n135 9.3005
R826 VDD1.n105 VDD1.n104 9.3005
R827 VDD1.n130 VDD1.n129 9.3005
R828 VDD1.n128 VDD1.n127 9.3005
R829 VDD1.n109 VDD1.n108 9.3005
R830 VDD1.n122 VDD1.n121 9.3005
R831 VDD1.n120 VDD1.n119 9.3005
R832 VDD1.n113 VDD1.n112 9.3005
R833 VDD1.n138 VDD1.n137 9.3005
R834 VDD1.n101 VDD1.n100 9.3005
R835 VDD1.n144 VDD1.n143 9.3005
R836 VDD1.n146 VDD1.n145 9.3005
R837 VDD1.n97 VDD1.n96 9.3005
R838 VDD1.n152 VDD1.n151 9.3005
R839 VDD1.n154 VDD1.n153 9.3005
R840 VDD1.n155 VDD1.n92 9.3005
R841 VDD1.n162 VDD1.n161 9.3005
R842 VDD1.n61 VDD1.n14 8.92171
R843 VDD1.n46 VDD1.n45 8.92171
R844 VDD1.n131 VDD1.n130 8.92171
R845 VDD1.n146 VDD1.n99 8.92171
R846 VDD1.n58 VDD1.n57 8.14595
R847 VDD1.n49 VDD1.n20 8.14595
R848 VDD1.n134 VDD1.n105 8.14595
R849 VDD1.n143 VDD1.n142 8.14595
R850 VDD1.n54 VDD1.n16 7.3702
R851 VDD1.n50 VDD1.n18 7.3702
R852 VDD1.n135 VDD1.n103 7.3702
R853 VDD1.n139 VDD1.n101 7.3702
R854 VDD1.n54 VDD1.n53 6.59444
R855 VDD1.n53 VDD1.n18 6.59444
R856 VDD1.n138 VDD1.n103 6.59444
R857 VDD1.n139 VDD1.n138 6.59444
R858 VDD1.n57 VDD1.n16 5.81868
R859 VDD1.n50 VDD1.n49 5.81868
R860 VDD1.n135 VDD1.n134 5.81868
R861 VDD1.n142 VDD1.n101 5.81868
R862 VDD1.n58 VDD1.n14 5.04292
R863 VDD1.n46 VDD1.n20 5.04292
R864 VDD1.n131 VDD1.n105 5.04292
R865 VDD1.n143 VDD1.n99 5.04292
R866 VDD1.n62 VDD1.n61 4.26717
R867 VDD1.n45 VDD1.n22 4.26717
R868 VDD1.n130 VDD1.n107 4.26717
R869 VDD1.n147 VDD1.n146 4.26717
R870 VDD1.n29 VDD1.n27 3.70982
R871 VDD1.n114 VDD1.n112 3.70982
R872 VDD1.n65 VDD1.n12 3.49141
R873 VDD1.n42 VDD1.n41 3.49141
R874 VDD1.n127 VDD1.n126 3.49141
R875 VDD1.n150 VDD1.n97 3.49141
R876 VDD1.n84 VDD1.n0 2.71565
R877 VDD1.n66 VDD1.n10 2.71565
R878 VDD1.n38 VDD1.n24 2.71565
R879 VDD1.n123 VDD1.n109 2.71565
R880 VDD1.n151 VDD1.n95 2.71565
R881 VDD1.n171 VDD1.n87 2.71565
R882 VDD1.n176 VDD1.t4 2.10166
R883 VDD1.n176 VDD1.t5 2.10166
R884 VDD1.n85 VDD1.t2 2.10166
R885 VDD1.n85 VDD1.t1 2.10166
R886 VDD1.n174 VDD1.t6 2.10166
R887 VDD1.n174 VDD1.t3 2.10166
R888 VDD1.n172 VDD1.t8 2.10166
R889 VDD1.n172 VDD1.t7 2.10166
R890 VDD1.n82 VDD1.n81 1.93989
R891 VDD1.n70 VDD1.n69 1.93989
R892 VDD1.n37 VDD1.n26 1.93989
R893 VDD1.n122 VDD1.n111 1.93989
R894 VDD1.n156 VDD1.n154 1.93989
R895 VDD1.n169 VDD1.n168 1.93989
R896 VDD1 VDD1.n177 1.40352
R897 VDD1.n78 VDD1.n2 1.16414
R898 VDD1.n73 VDD1.n7 1.16414
R899 VDD1.n34 VDD1.n33 1.16414
R900 VDD1.n119 VDD1.n118 1.16414
R901 VDD1.n155 VDD1.n93 1.16414
R902 VDD1.n165 VDD1.n89 1.16414
R903 VDD1 VDD1.n86 0.545759
R904 VDD1.n175 VDD1.n173 0.432223
R905 VDD1.n77 VDD1.n4 0.388379
R906 VDD1.n74 VDD1.n6 0.388379
R907 VDD1.n30 VDD1.n28 0.388379
R908 VDD1.n115 VDD1.n113 0.388379
R909 VDD1.n161 VDD1.n160 0.388379
R910 VDD1.n164 VDD1.n91 0.388379
R911 VDD1.n83 VDD1.n1 0.155672
R912 VDD1.n76 VDD1.n1 0.155672
R913 VDD1.n76 VDD1.n75 0.155672
R914 VDD1.n75 VDD1.n5 0.155672
R915 VDD1.n68 VDD1.n5 0.155672
R916 VDD1.n68 VDD1.n67 0.155672
R917 VDD1.n67 VDD1.n11 0.155672
R918 VDD1.n60 VDD1.n11 0.155672
R919 VDD1.n60 VDD1.n59 0.155672
R920 VDD1.n59 VDD1.n15 0.155672
R921 VDD1.n52 VDD1.n15 0.155672
R922 VDD1.n52 VDD1.n51 0.155672
R923 VDD1.n51 VDD1.n19 0.155672
R924 VDD1.n44 VDD1.n19 0.155672
R925 VDD1.n44 VDD1.n43 0.155672
R926 VDD1.n43 VDD1.n23 0.155672
R927 VDD1.n36 VDD1.n23 0.155672
R928 VDD1.n36 VDD1.n35 0.155672
R929 VDD1.n35 VDD1.n27 0.155672
R930 VDD1.n120 VDD1.n112 0.155672
R931 VDD1.n121 VDD1.n120 0.155672
R932 VDD1.n121 VDD1.n108 0.155672
R933 VDD1.n128 VDD1.n108 0.155672
R934 VDD1.n129 VDD1.n128 0.155672
R935 VDD1.n129 VDD1.n104 0.155672
R936 VDD1.n136 VDD1.n104 0.155672
R937 VDD1.n137 VDD1.n136 0.155672
R938 VDD1.n137 VDD1.n100 0.155672
R939 VDD1.n144 VDD1.n100 0.155672
R940 VDD1.n145 VDD1.n144 0.155672
R941 VDD1.n145 VDD1.n96 0.155672
R942 VDD1.n152 VDD1.n96 0.155672
R943 VDD1.n153 VDD1.n152 0.155672
R944 VDD1.n153 VDD1.n92 0.155672
R945 VDD1.n162 VDD1.n92 0.155672
R946 VDD1.n163 VDD1.n162 0.155672
R947 VDD1.n163 VDD1.n88 0.155672
R948 VDD1.n170 VDD1.n88 0.155672
R949 B.n608 B.n607 585
R950 B.n609 B.n86 585
R951 B.n611 B.n610 585
R952 B.n612 B.n85 585
R953 B.n614 B.n613 585
R954 B.n615 B.n84 585
R955 B.n617 B.n616 585
R956 B.n618 B.n83 585
R957 B.n620 B.n619 585
R958 B.n621 B.n82 585
R959 B.n623 B.n622 585
R960 B.n624 B.n81 585
R961 B.n626 B.n625 585
R962 B.n627 B.n80 585
R963 B.n629 B.n628 585
R964 B.n630 B.n79 585
R965 B.n632 B.n631 585
R966 B.n633 B.n78 585
R967 B.n635 B.n634 585
R968 B.n636 B.n77 585
R969 B.n638 B.n637 585
R970 B.n639 B.n76 585
R971 B.n641 B.n640 585
R972 B.n642 B.n75 585
R973 B.n644 B.n643 585
R974 B.n645 B.n74 585
R975 B.n647 B.n646 585
R976 B.n648 B.n73 585
R977 B.n650 B.n649 585
R978 B.n651 B.n72 585
R979 B.n653 B.n652 585
R980 B.n654 B.n71 585
R981 B.n656 B.n655 585
R982 B.n657 B.n70 585
R983 B.n659 B.n658 585
R984 B.n660 B.n69 585
R985 B.n662 B.n661 585
R986 B.n663 B.n68 585
R987 B.n665 B.n664 585
R988 B.n666 B.n67 585
R989 B.n668 B.n667 585
R990 B.n669 B.n66 585
R991 B.n671 B.n670 585
R992 B.n672 B.n65 585
R993 B.n674 B.n673 585
R994 B.n675 B.n64 585
R995 B.n677 B.n676 585
R996 B.n678 B.n63 585
R997 B.n680 B.n679 585
R998 B.n681 B.n62 585
R999 B.n683 B.n682 585
R1000 B.n684 B.n59 585
R1001 B.n687 B.n686 585
R1002 B.n688 B.n58 585
R1003 B.n690 B.n689 585
R1004 B.n691 B.n57 585
R1005 B.n693 B.n692 585
R1006 B.n694 B.n56 585
R1007 B.n696 B.n695 585
R1008 B.n697 B.n55 585
R1009 B.n699 B.n698 585
R1010 B.n701 B.n700 585
R1011 B.n702 B.n51 585
R1012 B.n704 B.n703 585
R1013 B.n705 B.n50 585
R1014 B.n707 B.n706 585
R1015 B.n708 B.n49 585
R1016 B.n710 B.n709 585
R1017 B.n711 B.n48 585
R1018 B.n713 B.n712 585
R1019 B.n714 B.n47 585
R1020 B.n716 B.n715 585
R1021 B.n717 B.n46 585
R1022 B.n719 B.n718 585
R1023 B.n720 B.n45 585
R1024 B.n722 B.n721 585
R1025 B.n723 B.n44 585
R1026 B.n725 B.n724 585
R1027 B.n726 B.n43 585
R1028 B.n728 B.n727 585
R1029 B.n729 B.n42 585
R1030 B.n731 B.n730 585
R1031 B.n732 B.n41 585
R1032 B.n734 B.n733 585
R1033 B.n735 B.n40 585
R1034 B.n737 B.n736 585
R1035 B.n738 B.n39 585
R1036 B.n740 B.n739 585
R1037 B.n741 B.n38 585
R1038 B.n743 B.n742 585
R1039 B.n744 B.n37 585
R1040 B.n746 B.n745 585
R1041 B.n747 B.n36 585
R1042 B.n749 B.n748 585
R1043 B.n750 B.n35 585
R1044 B.n752 B.n751 585
R1045 B.n753 B.n34 585
R1046 B.n755 B.n754 585
R1047 B.n756 B.n33 585
R1048 B.n758 B.n757 585
R1049 B.n759 B.n32 585
R1050 B.n761 B.n760 585
R1051 B.n762 B.n31 585
R1052 B.n764 B.n763 585
R1053 B.n765 B.n30 585
R1054 B.n767 B.n766 585
R1055 B.n768 B.n29 585
R1056 B.n770 B.n769 585
R1057 B.n771 B.n28 585
R1058 B.n773 B.n772 585
R1059 B.n774 B.n27 585
R1060 B.n776 B.n775 585
R1061 B.n777 B.n26 585
R1062 B.n606 B.n87 585
R1063 B.n605 B.n604 585
R1064 B.n603 B.n88 585
R1065 B.n602 B.n601 585
R1066 B.n600 B.n89 585
R1067 B.n599 B.n598 585
R1068 B.n597 B.n90 585
R1069 B.n596 B.n595 585
R1070 B.n594 B.n91 585
R1071 B.n593 B.n592 585
R1072 B.n591 B.n92 585
R1073 B.n590 B.n589 585
R1074 B.n588 B.n93 585
R1075 B.n587 B.n586 585
R1076 B.n585 B.n94 585
R1077 B.n584 B.n583 585
R1078 B.n582 B.n95 585
R1079 B.n581 B.n580 585
R1080 B.n579 B.n96 585
R1081 B.n578 B.n577 585
R1082 B.n576 B.n97 585
R1083 B.n575 B.n574 585
R1084 B.n573 B.n98 585
R1085 B.n572 B.n571 585
R1086 B.n570 B.n99 585
R1087 B.n569 B.n568 585
R1088 B.n567 B.n100 585
R1089 B.n566 B.n565 585
R1090 B.n564 B.n101 585
R1091 B.n563 B.n562 585
R1092 B.n561 B.n102 585
R1093 B.n560 B.n559 585
R1094 B.n558 B.n103 585
R1095 B.n557 B.n556 585
R1096 B.n555 B.n104 585
R1097 B.n554 B.n553 585
R1098 B.n552 B.n105 585
R1099 B.n551 B.n550 585
R1100 B.n549 B.n106 585
R1101 B.n548 B.n547 585
R1102 B.n546 B.n107 585
R1103 B.n545 B.n544 585
R1104 B.n543 B.n108 585
R1105 B.n542 B.n541 585
R1106 B.n540 B.n109 585
R1107 B.n539 B.n538 585
R1108 B.n537 B.n110 585
R1109 B.n536 B.n535 585
R1110 B.n534 B.n111 585
R1111 B.n533 B.n532 585
R1112 B.n531 B.n112 585
R1113 B.n530 B.n529 585
R1114 B.n528 B.n113 585
R1115 B.n527 B.n526 585
R1116 B.n525 B.n114 585
R1117 B.n524 B.n523 585
R1118 B.n522 B.n115 585
R1119 B.n521 B.n520 585
R1120 B.n519 B.n116 585
R1121 B.n518 B.n517 585
R1122 B.n516 B.n117 585
R1123 B.n515 B.n514 585
R1124 B.n513 B.n118 585
R1125 B.n512 B.n511 585
R1126 B.n510 B.n119 585
R1127 B.n509 B.n508 585
R1128 B.n507 B.n120 585
R1129 B.n506 B.n505 585
R1130 B.n504 B.n121 585
R1131 B.n503 B.n502 585
R1132 B.n501 B.n122 585
R1133 B.n500 B.n499 585
R1134 B.n498 B.n123 585
R1135 B.n497 B.n496 585
R1136 B.n495 B.n124 585
R1137 B.n494 B.n493 585
R1138 B.n492 B.n125 585
R1139 B.n491 B.n490 585
R1140 B.n489 B.n126 585
R1141 B.n488 B.n487 585
R1142 B.n486 B.n127 585
R1143 B.n485 B.n484 585
R1144 B.n483 B.n128 585
R1145 B.n482 B.n481 585
R1146 B.n480 B.n129 585
R1147 B.n479 B.n478 585
R1148 B.n477 B.n130 585
R1149 B.n476 B.n475 585
R1150 B.n474 B.n131 585
R1151 B.n473 B.n472 585
R1152 B.n471 B.n132 585
R1153 B.n470 B.n469 585
R1154 B.n468 B.n133 585
R1155 B.n467 B.n466 585
R1156 B.n465 B.n134 585
R1157 B.n464 B.n463 585
R1158 B.n462 B.n135 585
R1159 B.n291 B.n196 585
R1160 B.n293 B.n292 585
R1161 B.n294 B.n195 585
R1162 B.n296 B.n295 585
R1163 B.n297 B.n194 585
R1164 B.n299 B.n298 585
R1165 B.n300 B.n193 585
R1166 B.n302 B.n301 585
R1167 B.n303 B.n192 585
R1168 B.n305 B.n304 585
R1169 B.n306 B.n191 585
R1170 B.n308 B.n307 585
R1171 B.n309 B.n190 585
R1172 B.n311 B.n310 585
R1173 B.n312 B.n189 585
R1174 B.n314 B.n313 585
R1175 B.n315 B.n188 585
R1176 B.n317 B.n316 585
R1177 B.n318 B.n187 585
R1178 B.n320 B.n319 585
R1179 B.n321 B.n186 585
R1180 B.n323 B.n322 585
R1181 B.n324 B.n185 585
R1182 B.n326 B.n325 585
R1183 B.n327 B.n184 585
R1184 B.n329 B.n328 585
R1185 B.n330 B.n183 585
R1186 B.n332 B.n331 585
R1187 B.n333 B.n182 585
R1188 B.n335 B.n334 585
R1189 B.n336 B.n181 585
R1190 B.n338 B.n337 585
R1191 B.n339 B.n180 585
R1192 B.n341 B.n340 585
R1193 B.n342 B.n179 585
R1194 B.n344 B.n343 585
R1195 B.n345 B.n178 585
R1196 B.n347 B.n346 585
R1197 B.n348 B.n177 585
R1198 B.n350 B.n349 585
R1199 B.n351 B.n176 585
R1200 B.n353 B.n352 585
R1201 B.n354 B.n175 585
R1202 B.n356 B.n355 585
R1203 B.n357 B.n174 585
R1204 B.n359 B.n358 585
R1205 B.n360 B.n173 585
R1206 B.n362 B.n361 585
R1207 B.n363 B.n172 585
R1208 B.n365 B.n364 585
R1209 B.n366 B.n171 585
R1210 B.n368 B.n367 585
R1211 B.n370 B.n369 585
R1212 B.n371 B.n167 585
R1213 B.n373 B.n372 585
R1214 B.n374 B.n166 585
R1215 B.n376 B.n375 585
R1216 B.n377 B.n165 585
R1217 B.n379 B.n378 585
R1218 B.n380 B.n164 585
R1219 B.n382 B.n381 585
R1220 B.n384 B.n161 585
R1221 B.n386 B.n385 585
R1222 B.n387 B.n160 585
R1223 B.n389 B.n388 585
R1224 B.n390 B.n159 585
R1225 B.n392 B.n391 585
R1226 B.n393 B.n158 585
R1227 B.n395 B.n394 585
R1228 B.n396 B.n157 585
R1229 B.n398 B.n397 585
R1230 B.n399 B.n156 585
R1231 B.n401 B.n400 585
R1232 B.n402 B.n155 585
R1233 B.n404 B.n403 585
R1234 B.n405 B.n154 585
R1235 B.n407 B.n406 585
R1236 B.n408 B.n153 585
R1237 B.n410 B.n409 585
R1238 B.n411 B.n152 585
R1239 B.n413 B.n412 585
R1240 B.n414 B.n151 585
R1241 B.n416 B.n415 585
R1242 B.n417 B.n150 585
R1243 B.n419 B.n418 585
R1244 B.n420 B.n149 585
R1245 B.n422 B.n421 585
R1246 B.n423 B.n148 585
R1247 B.n425 B.n424 585
R1248 B.n426 B.n147 585
R1249 B.n428 B.n427 585
R1250 B.n429 B.n146 585
R1251 B.n431 B.n430 585
R1252 B.n432 B.n145 585
R1253 B.n434 B.n433 585
R1254 B.n435 B.n144 585
R1255 B.n437 B.n436 585
R1256 B.n438 B.n143 585
R1257 B.n440 B.n439 585
R1258 B.n441 B.n142 585
R1259 B.n443 B.n442 585
R1260 B.n444 B.n141 585
R1261 B.n446 B.n445 585
R1262 B.n447 B.n140 585
R1263 B.n449 B.n448 585
R1264 B.n450 B.n139 585
R1265 B.n452 B.n451 585
R1266 B.n453 B.n138 585
R1267 B.n455 B.n454 585
R1268 B.n456 B.n137 585
R1269 B.n458 B.n457 585
R1270 B.n459 B.n136 585
R1271 B.n461 B.n460 585
R1272 B.n290 B.n289 585
R1273 B.n288 B.n197 585
R1274 B.n287 B.n286 585
R1275 B.n285 B.n198 585
R1276 B.n284 B.n283 585
R1277 B.n282 B.n199 585
R1278 B.n281 B.n280 585
R1279 B.n279 B.n200 585
R1280 B.n278 B.n277 585
R1281 B.n276 B.n201 585
R1282 B.n275 B.n274 585
R1283 B.n273 B.n202 585
R1284 B.n272 B.n271 585
R1285 B.n270 B.n203 585
R1286 B.n269 B.n268 585
R1287 B.n267 B.n204 585
R1288 B.n266 B.n265 585
R1289 B.n264 B.n205 585
R1290 B.n263 B.n262 585
R1291 B.n261 B.n206 585
R1292 B.n260 B.n259 585
R1293 B.n258 B.n207 585
R1294 B.n257 B.n256 585
R1295 B.n255 B.n208 585
R1296 B.n254 B.n253 585
R1297 B.n252 B.n209 585
R1298 B.n251 B.n250 585
R1299 B.n249 B.n210 585
R1300 B.n248 B.n247 585
R1301 B.n246 B.n211 585
R1302 B.n245 B.n244 585
R1303 B.n243 B.n212 585
R1304 B.n242 B.n241 585
R1305 B.n240 B.n213 585
R1306 B.n239 B.n238 585
R1307 B.n237 B.n214 585
R1308 B.n236 B.n235 585
R1309 B.n234 B.n215 585
R1310 B.n233 B.n232 585
R1311 B.n231 B.n216 585
R1312 B.n230 B.n229 585
R1313 B.n228 B.n217 585
R1314 B.n227 B.n226 585
R1315 B.n225 B.n218 585
R1316 B.n224 B.n223 585
R1317 B.n222 B.n219 585
R1318 B.n221 B.n220 585
R1319 B.n2 B.n0 585
R1320 B.n849 B.n1 585
R1321 B.n848 B.n847 585
R1322 B.n846 B.n3 585
R1323 B.n845 B.n844 585
R1324 B.n843 B.n4 585
R1325 B.n842 B.n841 585
R1326 B.n840 B.n5 585
R1327 B.n839 B.n838 585
R1328 B.n837 B.n6 585
R1329 B.n836 B.n835 585
R1330 B.n834 B.n7 585
R1331 B.n833 B.n832 585
R1332 B.n831 B.n8 585
R1333 B.n830 B.n829 585
R1334 B.n828 B.n9 585
R1335 B.n827 B.n826 585
R1336 B.n825 B.n10 585
R1337 B.n824 B.n823 585
R1338 B.n822 B.n11 585
R1339 B.n821 B.n820 585
R1340 B.n819 B.n12 585
R1341 B.n818 B.n817 585
R1342 B.n816 B.n13 585
R1343 B.n815 B.n814 585
R1344 B.n813 B.n14 585
R1345 B.n812 B.n811 585
R1346 B.n810 B.n15 585
R1347 B.n809 B.n808 585
R1348 B.n807 B.n16 585
R1349 B.n806 B.n805 585
R1350 B.n804 B.n17 585
R1351 B.n803 B.n802 585
R1352 B.n801 B.n18 585
R1353 B.n800 B.n799 585
R1354 B.n798 B.n19 585
R1355 B.n797 B.n796 585
R1356 B.n795 B.n20 585
R1357 B.n794 B.n793 585
R1358 B.n792 B.n21 585
R1359 B.n791 B.n790 585
R1360 B.n789 B.n22 585
R1361 B.n788 B.n787 585
R1362 B.n786 B.n23 585
R1363 B.n785 B.n784 585
R1364 B.n783 B.n24 585
R1365 B.n782 B.n781 585
R1366 B.n780 B.n25 585
R1367 B.n779 B.n778 585
R1368 B.n851 B.n850 585
R1369 B.n291 B.n290 516.524
R1370 B.n778 B.n777 516.524
R1371 B.n460 B.n135 516.524
R1372 B.n608 B.n87 516.524
R1373 B.n162 B.t11 481.957
R1374 B.n60 B.t7 481.957
R1375 B.n168 B.t2 481.957
R1376 B.n52 B.t4 481.957
R1377 B.n163 B.t10 438.125
R1378 B.n61 B.t8 438.125
R1379 B.n169 B.t1 438.125
R1380 B.n53 B.t5 438.125
R1381 B.n162 B.t9 399.923
R1382 B.n168 B.t0 399.923
R1383 B.n52 B.t3 399.923
R1384 B.n60 B.t6 399.923
R1385 B.n290 B.n197 163.367
R1386 B.n286 B.n197 163.367
R1387 B.n286 B.n285 163.367
R1388 B.n285 B.n284 163.367
R1389 B.n284 B.n199 163.367
R1390 B.n280 B.n199 163.367
R1391 B.n280 B.n279 163.367
R1392 B.n279 B.n278 163.367
R1393 B.n278 B.n201 163.367
R1394 B.n274 B.n201 163.367
R1395 B.n274 B.n273 163.367
R1396 B.n273 B.n272 163.367
R1397 B.n272 B.n203 163.367
R1398 B.n268 B.n203 163.367
R1399 B.n268 B.n267 163.367
R1400 B.n267 B.n266 163.367
R1401 B.n266 B.n205 163.367
R1402 B.n262 B.n205 163.367
R1403 B.n262 B.n261 163.367
R1404 B.n261 B.n260 163.367
R1405 B.n260 B.n207 163.367
R1406 B.n256 B.n207 163.367
R1407 B.n256 B.n255 163.367
R1408 B.n255 B.n254 163.367
R1409 B.n254 B.n209 163.367
R1410 B.n250 B.n209 163.367
R1411 B.n250 B.n249 163.367
R1412 B.n249 B.n248 163.367
R1413 B.n248 B.n211 163.367
R1414 B.n244 B.n211 163.367
R1415 B.n244 B.n243 163.367
R1416 B.n243 B.n242 163.367
R1417 B.n242 B.n213 163.367
R1418 B.n238 B.n213 163.367
R1419 B.n238 B.n237 163.367
R1420 B.n237 B.n236 163.367
R1421 B.n236 B.n215 163.367
R1422 B.n232 B.n215 163.367
R1423 B.n232 B.n231 163.367
R1424 B.n231 B.n230 163.367
R1425 B.n230 B.n217 163.367
R1426 B.n226 B.n217 163.367
R1427 B.n226 B.n225 163.367
R1428 B.n225 B.n224 163.367
R1429 B.n224 B.n219 163.367
R1430 B.n220 B.n219 163.367
R1431 B.n220 B.n2 163.367
R1432 B.n850 B.n2 163.367
R1433 B.n850 B.n849 163.367
R1434 B.n849 B.n848 163.367
R1435 B.n848 B.n3 163.367
R1436 B.n844 B.n3 163.367
R1437 B.n844 B.n843 163.367
R1438 B.n843 B.n842 163.367
R1439 B.n842 B.n5 163.367
R1440 B.n838 B.n5 163.367
R1441 B.n838 B.n837 163.367
R1442 B.n837 B.n836 163.367
R1443 B.n836 B.n7 163.367
R1444 B.n832 B.n7 163.367
R1445 B.n832 B.n831 163.367
R1446 B.n831 B.n830 163.367
R1447 B.n830 B.n9 163.367
R1448 B.n826 B.n9 163.367
R1449 B.n826 B.n825 163.367
R1450 B.n825 B.n824 163.367
R1451 B.n824 B.n11 163.367
R1452 B.n820 B.n11 163.367
R1453 B.n820 B.n819 163.367
R1454 B.n819 B.n818 163.367
R1455 B.n818 B.n13 163.367
R1456 B.n814 B.n13 163.367
R1457 B.n814 B.n813 163.367
R1458 B.n813 B.n812 163.367
R1459 B.n812 B.n15 163.367
R1460 B.n808 B.n15 163.367
R1461 B.n808 B.n807 163.367
R1462 B.n807 B.n806 163.367
R1463 B.n806 B.n17 163.367
R1464 B.n802 B.n17 163.367
R1465 B.n802 B.n801 163.367
R1466 B.n801 B.n800 163.367
R1467 B.n800 B.n19 163.367
R1468 B.n796 B.n19 163.367
R1469 B.n796 B.n795 163.367
R1470 B.n795 B.n794 163.367
R1471 B.n794 B.n21 163.367
R1472 B.n790 B.n21 163.367
R1473 B.n790 B.n789 163.367
R1474 B.n789 B.n788 163.367
R1475 B.n788 B.n23 163.367
R1476 B.n784 B.n23 163.367
R1477 B.n784 B.n783 163.367
R1478 B.n783 B.n782 163.367
R1479 B.n782 B.n25 163.367
R1480 B.n778 B.n25 163.367
R1481 B.n292 B.n291 163.367
R1482 B.n292 B.n195 163.367
R1483 B.n296 B.n195 163.367
R1484 B.n297 B.n296 163.367
R1485 B.n298 B.n297 163.367
R1486 B.n298 B.n193 163.367
R1487 B.n302 B.n193 163.367
R1488 B.n303 B.n302 163.367
R1489 B.n304 B.n303 163.367
R1490 B.n304 B.n191 163.367
R1491 B.n308 B.n191 163.367
R1492 B.n309 B.n308 163.367
R1493 B.n310 B.n309 163.367
R1494 B.n310 B.n189 163.367
R1495 B.n314 B.n189 163.367
R1496 B.n315 B.n314 163.367
R1497 B.n316 B.n315 163.367
R1498 B.n316 B.n187 163.367
R1499 B.n320 B.n187 163.367
R1500 B.n321 B.n320 163.367
R1501 B.n322 B.n321 163.367
R1502 B.n322 B.n185 163.367
R1503 B.n326 B.n185 163.367
R1504 B.n327 B.n326 163.367
R1505 B.n328 B.n327 163.367
R1506 B.n328 B.n183 163.367
R1507 B.n332 B.n183 163.367
R1508 B.n333 B.n332 163.367
R1509 B.n334 B.n333 163.367
R1510 B.n334 B.n181 163.367
R1511 B.n338 B.n181 163.367
R1512 B.n339 B.n338 163.367
R1513 B.n340 B.n339 163.367
R1514 B.n340 B.n179 163.367
R1515 B.n344 B.n179 163.367
R1516 B.n345 B.n344 163.367
R1517 B.n346 B.n345 163.367
R1518 B.n346 B.n177 163.367
R1519 B.n350 B.n177 163.367
R1520 B.n351 B.n350 163.367
R1521 B.n352 B.n351 163.367
R1522 B.n352 B.n175 163.367
R1523 B.n356 B.n175 163.367
R1524 B.n357 B.n356 163.367
R1525 B.n358 B.n357 163.367
R1526 B.n358 B.n173 163.367
R1527 B.n362 B.n173 163.367
R1528 B.n363 B.n362 163.367
R1529 B.n364 B.n363 163.367
R1530 B.n364 B.n171 163.367
R1531 B.n368 B.n171 163.367
R1532 B.n369 B.n368 163.367
R1533 B.n369 B.n167 163.367
R1534 B.n373 B.n167 163.367
R1535 B.n374 B.n373 163.367
R1536 B.n375 B.n374 163.367
R1537 B.n375 B.n165 163.367
R1538 B.n379 B.n165 163.367
R1539 B.n380 B.n379 163.367
R1540 B.n381 B.n380 163.367
R1541 B.n381 B.n161 163.367
R1542 B.n386 B.n161 163.367
R1543 B.n387 B.n386 163.367
R1544 B.n388 B.n387 163.367
R1545 B.n388 B.n159 163.367
R1546 B.n392 B.n159 163.367
R1547 B.n393 B.n392 163.367
R1548 B.n394 B.n393 163.367
R1549 B.n394 B.n157 163.367
R1550 B.n398 B.n157 163.367
R1551 B.n399 B.n398 163.367
R1552 B.n400 B.n399 163.367
R1553 B.n400 B.n155 163.367
R1554 B.n404 B.n155 163.367
R1555 B.n405 B.n404 163.367
R1556 B.n406 B.n405 163.367
R1557 B.n406 B.n153 163.367
R1558 B.n410 B.n153 163.367
R1559 B.n411 B.n410 163.367
R1560 B.n412 B.n411 163.367
R1561 B.n412 B.n151 163.367
R1562 B.n416 B.n151 163.367
R1563 B.n417 B.n416 163.367
R1564 B.n418 B.n417 163.367
R1565 B.n418 B.n149 163.367
R1566 B.n422 B.n149 163.367
R1567 B.n423 B.n422 163.367
R1568 B.n424 B.n423 163.367
R1569 B.n424 B.n147 163.367
R1570 B.n428 B.n147 163.367
R1571 B.n429 B.n428 163.367
R1572 B.n430 B.n429 163.367
R1573 B.n430 B.n145 163.367
R1574 B.n434 B.n145 163.367
R1575 B.n435 B.n434 163.367
R1576 B.n436 B.n435 163.367
R1577 B.n436 B.n143 163.367
R1578 B.n440 B.n143 163.367
R1579 B.n441 B.n440 163.367
R1580 B.n442 B.n441 163.367
R1581 B.n442 B.n141 163.367
R1582 B.n446 B.n141 163.367
R1583 B.n447 B.n446 163.367
R1584 B.n448 B.n447 163.367
R1585 B.n448 B.n139 163.367
R1586 B.n452 B.n139 163.367
R1587 B.n453 B.n452 163.367
R1588 B.n454 B.n453 163.367
R1589 B.n454 B.n137 163.367
R1590 B.n458 B.n137 163.367
R1591 B.n459 B.n458 163.367
R1592 B.n460 B.n459 163.367
R1593 B.n464 B.n135 163.367
R1594 B.n465 B.n464 163.367
R1595 B.n466 B.n465 163.367
R1596 B.n466 B.n133 163.367
R1597 B.n470 B.n133 163.367
R1598 B.n471 B.n470 163.367
R1599 B.n472 B.n471 163.367
R1600 B.n472 B.n131 163.367
R1601 B.n476 B.n131 163.367
R1602 B.n477 B.n476 163.367
R1603 B.n478 B.n477 163.367
R1604 B.n478 B.n129 163.367
R1605 B.n482 B.n129 163.367
R1606 B.n483 B.n482 163.367
R1607 B.n484 B.n483 163.367
R1608 B.n484 B.n127 163.367
R1609 B.n488 B.n127 163.367
R1610 B.n489 B.n488 163.367
R1611 B.n490 B.n489 163.367
R1612 B.n490 B.n125 163.367
R1613 B.n494 B.n125 163.367
R1614 B.n495 B.n494 163.367
R1615 B.n496 B.n495 163.367
R1616 B.n496 B.n123 163.367
R1617 B.n500 B.n123 163.367
R1618 B.n501 B.n500 163.367
R1619 B.n502 B.n501 163.367
R1620 B.n502 B.n121 163.367
R1621 B.n506 B.n121 163.367
R1622 B.n507 B.n506 163.367
R1623 B.n508 B.n507 163.367
R1624 B.n508 B.n119 163.367
R1625 B.n512 B.n119 163.367
R1626 B.n513 B.n512 163.367
R1627 B.n514 B.n513 163.367
R1628 B.n514 B.n117 163.367
R1629 B.n518 B.n117 163.367
R1630 B.n519 B.n518 163.367
R1631 B.n520 B.n519 163.367
R1632 B.n520 B.n115 163.367
R1633 B.n524 B.n115 163.367
R1634 B.n525 B.n524 163.367
R1635 B.n526 B.n525 163.367
R1636 B.n526 B.n113 163.367
R1637 B.n530 B.n113 163.367
R1638 B.n531 B.n530 163.367
R1639 B.n532 B.n531 163.367
R1640 B.n532 B.n111 163.367
R1641 B.n536 B.n111 163.367
R1642 B.n537 B.n536 163.367
R1643 B.n538 B.n537 163.367
R1644 B.n538 B.n109 163.367
R1645 B.n542 B.n109 163.367
R1646 B.n543 B.n542 163.367
R1647 B.n544 B.n543 163.367
R1648 B.n544 B.n107 163.367
R1649 B.n548 B.n107 163.367
R1650 B.n549 B.n548 163.367
R1651 B.n550 B.n549 163.367
R1652 B.n550 B.n105 163.367
R1653 B.n554 B.n105 163.367
R1654 B.n555 B.n554 163.367
R1655 B.n556 B.n555 163.367
R1656 B.n556 B.n103 163.367
R1657 B.n560 B.n103 163.367
R1658 B.n561 B.n560 163.367
R1659 B.n562 B.n561 163.367
R1660 B.n562 B.n101 163.367
R1661 B.n566 B.n101 163.367
R1662 B.n567 B.n566 163.367
R1663 B.n568 B.n567 163.367
R1664 B.n568 B.n99 163.367
R1665 B.n572 B.n99 163.367
R1666 B.n573 B.n572 163.367
R1667 B.n574 B.n573 163.367
R1668 B.n574 B.n97 163.367
R1669 B.n578 B.n97 163.367
R1670 B.n579 B.n578 163.367
R1671 B.n580 B.n579 163.367
R1672 B.n580 B.n95 163.367
R1673 B.n584 B.n95 163.367
R1674 B.n585 B.n584 163.367
R1675 B.n586 B.n585 163.367
R1676 B.n586 B.n93 163.367
R1677 B.n590 B.n93 163.367
R1678 B.n591 B.n590 163.367
R1679 B.n592 B.n591 163.367
R1680 B.n592 B.n91 163.367
R1681 B.n596 B.n91 163.367
R1682 B.n597 B.n596 163.367
R1683 B.n598 B.n597 163.367
R1684 B.n598 B.n89 163.367
R1685 B.n602 B.n89 163.367
R1686 B.n603 B.n602 163.367
R1687 B.n604 B.n603 163.367
R1688 B.n604 B.n87 163.367
R1689 B.n777 B.n776 163.367
R1690 B.n776 B.n27 163.367
R1691 B.n772 B.n27 163.367
R1692 B.n772 B.n771 163.367
R1693 B.n771 B.n770 163.367
R1694 B.n770 B.n29 163.367
R1695 B.n766 B.n29 163.367
R1696 B.n766 B.n765 163.367
R1697 B.n765 B.n764 163.367
R1698 B.n764 B.n31 163.367
R1699 B.n760 B.n31 163.367
R1700 B.n760 B.n759 163.367
R1701 B.n759 B.n758 163.367
R1702 B.n758 B.n33 163.367
R1703 B.n754 B.n33 163.367
R1704 B.n754 B.n753 163.367
R1705 B.n753 B.n752 163.367
R1706 B.n752 B.n35 163.367
R1707 B.n748 B.n35 163.367
R1708 B.n748 B.n747 163.367
R1709 B.n747 B.n746 163.367
R1710 B.n746 B.n37 163.367
R1711 B.n742 B.n37 163.367
R1712 B.n742 B.n741 163.367
R1713 B.n741 B.n740 163.367
R1714 B.n740 B.n39 163.367
R1715 B.n736 B.n39 163.367
R1716 B.n736 B.n735 163.367
R1717 B.n735 B.n734 163.367
R1718 B.n734 B.n41 163.367
R1719 B.n730 B.n41 163.367
R1720 B.n730 B.n729 163.367
R1721 B.n729 B.n728 163.367
R1722 B.n728 B.n43 163.367
R1723 B.n724 B.n43 163.367
R1724 B.n724 B.n723 163.367
R1725 B.n723 B.n722 163.367
R1726 B.n722 B.n45 163.367
R1727 B.n718 B.n45 163.367
R1728 B.n718 B.n717 163.367
R1729 B.n717 B.n716 163.367
R1730 B.n716 B.n47 163.367
R1731 B.n712 B.n47 163.367
R1732 B.n712 B.n711 163.367
R1733 B.n711 B.n710 163.367
R1734 B.n710 B.n49 163.367
R1735 B.n706 B.n49 163.367
R1736 B.n706 B.n705 163.367
R1737 B.n705 B.n704 163.367
R1738 B.n704 B.n51 163.367
R1739 B.n700 B.n51 163.367
R1740 B.n700 B.n699 163.367
R1741 B.n699 B.n55 163.367
R1742 B.n695 B.n55 163.367
R1743 B.n695 B.n694 163.367
R1744 B.n694 B.n693 163.367
R1745 B.n693 B.n57 163.367
R1746 B.n689 B.n57 163.367
R1747 B.n689 B.n688 163.367
R1748 B.n688 B.n687 163.367
R1749 B.n687 B.n59 163.367
R1750 B.n682 B.n59 163.367
R1751 B.n682 B.n681 163.367
R1752 B.n681 B.n680 163.367
R1753 B.n680 B.n63 163.367
R1754 B.n676 B.n63 163.367
R1755 B.n676 B.n675 163.367
R1756 B.n675 B.n674 163.367
R1757 B.n674 B.n65 163.367
R1758 B.n670 B.n65 163.367
R1759 B.n670 B.n669 163.367
R1760 B.n669 B.n668 163.367
R1761 B.n668 B.n67 163.367
R1762 B.n664 B.n67 163.367
R1763 B.n664 B.n663 163.367
R1764 B.n663 B.n662 163.367
R1765 B.n662 B.n69 163.367
R1766 B.n658 B.n69 163.367
R1767 B.n658 B.n657 163.367
R1768 B.n657 B.n656 163.367
R1769 B.n656 B.n71 163.367
R1770 B.n652 B.n71 163.367
R1771 B.n652 B.n651 163.367
R1772 B.n651 B.n650 163.367
R1773 B.n650 B.n73 163.367
R1774 B.n646 B.n73 163.367
R1775 B.n646 B.n645 163.367
R1776 B.n645 B.n644 163.367
R1777 B.n644 B.n75 163.367
R1778 B.n640 B.n75 163.367
R1779 B.n640 B.n639 163.367
R1780 B.n639 B.n638 163.367
R1781 B.n638 B.n77 163.367
R1782 B.n634 B.n77 163.367
R1783 B.n634 B.n633 163.367
R1784 B.n633 B.n632 163.367
R1785 B.n632 B.n79 163.367
R1786 B.n628 B.n79 163.367
R1787 B.n628 B.n627 163.367
R1788 B.n627 B.n626 163.367
R1789 B.n626 B.n81 163.367
R1790 B.n622 B.n81 163.367
R1791 B.n622 B.n621 163.367
R1792 B.n621 B.n620 163.367
R1793 B.n620 B.n83 163.367
R1794 B.n616 B.n83 163.367
R1795 B.n616 B.n615 163.367
R1796 B.n615 B.n614 163.367
R1797 B.n614 B.n85 163.367
R1798 B.n610 B.n85 163.367
R1799 B.n610 B.n609 163.367
R1800 B.n609 B.n608 163.367
R1801 B.n383 B.n163 59.5399
R1802 B.n170 B.n169 59.5399
R1803 B.n54 B.n53 59.5399
R1804 B.n685 B.n61 59.5399
R1805 B.n163 B.n162 43.8308
R1806 B.n169 B.n168 43.8308
R1807 B.n53 B.n52 43.8308
R1808 B.n61 B.n60 43.8308
R1809 B.n779 B.n26 33.5615
R1810 B.n607 B.n606 33.5615
R1811 B.n462 B.n461 33.5615
R1812 B.n289 B.n196 33.5615
R1813 B B.n851 18.0485
R1814 B.n775 B.n26 10.6151
R1815 B.n775 B.n774 10.6151
R1816 B.n774 B.n773 10.6151
R1817 B.n773 B.n28 10.6151
R1818 B.n769 B.n28 10.6151
R1819 B.n769 B.n768 10.6151
R1820 B.n768 B.n767 10.6151
R1821 B.n767 B.n30 10.6151
R1822 B.n763 B.n30 10.6151
R1823 B.n763 B.n762 10.6151
R1824 B.n762 B.n761 10.6151
R1825 B.n761 B.n32 10.6151
R1826 B.n757 B.n32 10.6151
R1827 B.n757 B.n756 10.6151
R1828 B.n756 B.n755 10.6151
R1829 B.n755 B.n34 10.6151
R1830 B.n751 B.n34 10.6151
R1831 B.n751 B.n750 10.6151
R1832 B.n750 B.n749 10.6151
R1833 B.n749 B.n36 10.6151
R1834 B.n745 B.n36 10.6151
R1835 B.n745 B.n744 10.6151
R1836 B.n744 B.n743 10.6151
R1837 B.n743 B.n38 10.6151
R1838 B.n739 B.n38 10.6151
R1839 B.n739 B.n738 10.6151
R1840 B.n738 B.n737 10.6151
R1841 B.n737 B.n40 10.6151
R1842 B.n733 B.n40 10.6151
R1843 B.n733 B.n732 10.6151
R1844 B.n732 B.n731 10.6151
R1845 B.n731 B.n42 10.6151
R1846 B.n727 B.n42 10.6151
R1847 B.n727 B.n726 10.6151
R1848 B.n726 B.n725 10.6151
R1849 B.n725 B.n44 10.6151
R1850 B.n721 B.n44 10.6151
R1851 B.n721 B.n720 10.6151
R1852 B.n720 B.n719 10.6151
R1853 B.n719 B.n46 10.6151
R1854 B.n715 B.n46 10.6151
R1855 B.n715 B.n714 10.6151
R1856 B.n714 B.n713 10.6151
R1857 B.n713 B.n48 10.6151
R1858 B.n709 B.n48 10.6151
R1859 B.n709 B.n708 10.6151
R1860 B.n708 B.n707 10.6151
R1861 B.n707 B.n50 10.6151
R1862 B.n703 B.n50 10.6151
R1863 B.n703 B.n702 10.6151
R1864 B.n702 B.n701 10.6151
R1865 B.n698 B.n697 10.6151
R1866 B.n697 B.n696 10.6151
R1867 B.n696 B.n56 10.6151
R1868 B.n692 B.n56 10.6151
R1869 B.n692 B.n691 10.6151
R1870 B.n691 B.n690 10.6151
R1871 B.n690 B.n58 10.6151
R1872 B.n686 B.n58 10.6151
R1873 B.n684 B.n683 10.6151
R1874 B.n683 B.n62 10.6151
R1875 B.n679 B.n62 10.6151
R1876 B.n679 B.n678 10.6151
R1877 B.n678 B.n677 10.6151
R1878 B.n677 B.n64 10.6151
R1879 B.n673 B.n64 10.6151
R1880 B.n673 B.n672 10.6151
R1881 B.n672 B.n671 10.6151
R1882 B.n671 B.n66 10.6151
R1883 B.n667 B.n66 10.6151
R1884 B.n667 B.n666 10.6151
R1885 B.n666 B.n665 10.6151
R1886 B.n665 B.n68 10.6151
R1887 B.n661 B.n68 10.6151
R1888 B.n661 B.n660 10.6151
R1889 B.n660 B.n659 10.6151
R1890 B.n659 B.n70 10.6151
R1891 B.n655 B.n70 10.6151
R1892 B.n655 B.n654 10.6151
R1893 B.n654 B.n653 10.6151
R1894 B.n653 B.n72 10.6151
R1895 B.n649 B.n72 10.6151
R1896 B.n649 B.n648 10.6151
R1897 B.n648 B.n647 10.6151
R1898 B.n647 B.n74 10.6151
R1899 B.n643 B.n74 10.6151
R1900 B.n643 B.n642 10.6151
R1901 B.n642 B.n641 10.6151
R1902 B.n641 B.n76 10.6151
R1903 B.n637 B.n76 10.6151
R1904 B.n637 B.n636 10.6151
R1905 B.n636 B.n635 10.6151
R1906 B.n635 B.n78 10.6151
R1907 B.n631 B.n78 10.6151
R1908 B.n631 B.n630 10.6151
R1909 B.n630 B.n629 10.6151
R1910 B.n629 B.n80 10.6151
R1911 B.n625 B.n80 10.6151
R1912 B.n625 B.n624 10.6151
R1913 B.n624 B.n623 10.6151
R1914 B.n623 B.n82 10.6151
R1915 B.n619 B.n82 10.6151
R1916 B.n619 B.n618 10.6151
R1917 B.n618 B.n617 10.6151
R1918 B.n617 B.n84 10.6151
R1919 B.n613 B.n84 10.6151
R1920 B.n613 B.n612 10.6151
R1921 B.n612 B.n611 10.6151
R1922 B.n611 B.n86 10.6151
R1923 B.n607 B.n86 10.6151
R1924 B.n463 B.n462 10.6151
R1925 B.n463 B.n134 10.6151
R1926 B.n467 B.n134 10.6151
R1927 B.n468 B.n467 10.6151
R1928 B.n469 B.n468 10.6151
R1929 B.n469 B.n132 10.6151
R1930 B.n473 B.n132 10.6151
R1931 B.n474 B.n473 10.6151
R1932 B.n475 B.n474 10.6151
R1933 B.n475 B.n130 10.6151
R1934 B.n479 B.n130 10.6151
R1935 B.n480 B.n479 10.6151
R1936 B.n481 B.n480 10.6151
R1937 B.n481 B.n128 10.6151
R1938 B.n485 B.n128 10.6151
R1939 B.n486 B.n485 10.6151
R1940 B.n487 B.n486 10.6151
R1941 B.n487 B.n126 10.6151
R1942 B.n491 B.n126 10.6151
R1943 B.n492 B.n491 10.6151
R1944 B.n493 B.n492 10.6151
R1945 B.n493 B.n124 10.6151
R1946 B.n497 B.n124 10.6151
R1947 B.n498 B.n497 10.6151
R1948 B.n499 B.n498 10.6151
R1949 B.n499 B.n122 10.6151
R1950 B.n503 B.n122 10.6151
R1951 B.n504 B.n503 10.6151
R1952 B.n505 B.n504 10.6151
R1953 B.n505 B.n120 10.6151
R1954 B.n509 B.n120 10.6151
R1955 B.n510 B.n509 10.6151
R1956 B.n511 B.n510 10.6151
R1957 B.n511 B.n118 10.6151
R1958 B.n515 B.n118 10.6151
R1959 B.n516 B.n515 10.6151
R1960 B.n517 B.n516 10.6151
R1961 B.n517 B.n116 10.6151
R1962 B.n521 B.n116 10.6151
R1963 B.n522 B.n521 10.6151
R1964 B.n523 B.n522 10.6151
R1965 B.n523 B.n114 10.6151
R1966 B.n527 B.n114 10.6151
R1967 B.n528 B.n527 10.6151
R1968 B.n529 B.n528 10.6151
R1969 B.n529 B.n112 10.6151
R1970 B.n533 B.n112 10.6151
R1971 B.n534 B.n533 10.6151
R1972 B.n535 B.n534 10.6151
R1973 B.n535 B.n110 10.6151
R1974 B.n539 B.n110 10.6151
R1975 B.n540 B.n539 10.6151
R1976 B.n541 B.n540 10.6151
R1977 B.n541 B.n108 10.6151
R1978 B.n545 B.n108 10.6151
R1979 B.n546 B.n545 10.6151
R1980 B.n547 B.n546 10.6151
R1981 B.n547 B.n106 10.6151
R1982 B.n551 B.n106 10.6151
R1983 B.n552 B.n551 10.6151
R1984 B.n553 B.n552 10.6151
R1985 B.n553 B.n104 10.6151
R1986 B.n557 B.n104 10.6151
R1987 B.n558 B.n557 10.6151
R1988 B.n559 B.n558 10.6151
R1989 B.n559 B.n102 10.6151
R1990 B.n563 B.n102 10.6151
R1991 B.n564 B.n563 10.6151
R1992 B.n565 B.n564 10.6151
R1993 B.n565 B.n100 10.6151
R1994 B.n569 B.n100 10.6151
R1995 B.n570 B.n569 10.6151
R1996 B.n571 B.n570 10.6151
R1997 B.n571 B.n98 10.6151
R1998 B.n575 B.n98 10.6151
R1999 B.n576 B.n575 10.6151
R2000 B.n577 B.n576 10.6151
R2001 B.n577 B.n96 10.6151
R2002 B.n581 B.n96 10.6151
R2003 B.n582 B.n581 10.6151
R2004 B.n583 B.n582 10.6151
R2005 B.n583 B.n94 10.6151
R2006 B.n587 B.n94 10.6151
R2007 B.n588 B.n587 10.6151
R2008 B.n589 B.n588 10.6151
R2009 B.n589 B.n92 10.6151
R2010 B.n593 B.n92 10.6151
R2011 B.n594 B.n593 10.6151
R2012 B.n595 B.n594 10.6151
R2013 B.n595 B.n90 10.6151
R2014 B.n599 B.n90 10.6151
R2015 B.n600 B.n599 10.6151
R2016 B.n601 B.n600 10.6151
R2017 B.n601 B.n88 10.6151
R2018 B.n605 B.n88 10.6151
R2019 B.n606 B.n605 10.6151
R2020 B.n293 B.n196 10.6151
R2021 B.n294 B.n293 10.6151
R2022 B.n295 B.n294 10.6151
R2023 B.n295 B.n194 10.6151
R2024 B.n299 B.n194 10.6151
R2025 B.n300 B.n299 10.6151
R2026 B.n301 B.n300 10.6151
R2027 B.n301 B.n192 10.6151
R2028 B.n305 B.n192 10.6151
R2029 B.n306 B.n305 10.6151
R2030 B.n307 B.n306 10.6151
R2031 B.n307 B.n190 10.6151
R2032 B.n311 B.n190 10.6151
R2033 B.n312 B.n311 10.6151
R2034 B.n313 B.n312 10.6151
R2035 B.n313 B.n188 10.6151
R2036 B.n317 B.n188 10.6151
R2037 B.n318 B.n317 10.6151
R2038 B.n319 B.n318 10.6151
R2039 B.n319 B.n186 10.6151
R2040 B.n323 B.n186 10.6151
R2041 B.n324 B.n323 10.6151
R2042 B.n325 B.n324 10.6151
R2043 B.n325 B.n184 10.6151
R2044 B.n329 B.n184 10.6151
R2045 B.n330 B.n329 10.6151
R2046 B.n331 B.n330 10.6151
R2047 B.n331 B.n182 10.6151
R2048 B.n335 B.n182 10.6151
R2049 B.n336 B.n335 10.6151
R2050 B.n337 B.n336 10.6151
R2051 B.n337 B.n180 10.6151
R2052 B.n341 B.n180 10.6151
R2053 B.n342 B.n341 10.6151
R2054 B.n343 B.n342 10.6151
R2055 B.n343 B.n178 10.6151
R2056 B.n347 B.n178 10.6151
R2057 B.n348 B.n347 10.6151
R2058 B.n349 B.n348 10.6151
R2059 B.n349 B.n176 10.6151
R2060 B.n353 B.n176 10.6151
R2061 B.n354 B.n353 10.6151
R2062 B.n355 B.n354 10.6151
R2063 B.n355 B.n174 10.6151
R2064 B.n359 B.n174 10.6151
R2065 B.n360 B.n359 10.6151
R2066 B.n361 B.n360 10.6151
R2067 B.n361 B.n172 10.6151
R2068 B.n365 B.n172 10.6151
R2069 B.n366 B.n365 10.6151
R2070 B.n367 B.n366 10.6151
R2071 B.n371 B.n370 10.6151
R2072 B.n372 B.n371 10.6151
R2073 B.n372 B.n166 10.6151
R2074 B.n376 B.n166 10.6151
R2075 B.n377 B.n376 10.6151
R2076 B.n378 B.n377 10.6151
R2077 B.n378 B.n164 10.6151
R2078 B.n382 B.n164 10.6151
R2079 B.n385 B.n384 10.6151
R2080 B.n385 B.n160 10.6151
R2081 B.n389 B.n160 10.6151
R2082 B.n390 B.n389 10.6151
R2083 B.n391 B.n390 10.6151
R2084 B.n391 B.n158 10.6151
R2085 B.n395 B.n158 10.6151
R2086 B.n396 B.n395 10.6151
R2087 B.n397 B.n396 10.6151
R2088 B.n397 B.n156 10.6151
R2089 B.n401 B.n156 10.6151
R2090 B.n402 B.n401 10.6151
R2091 B.n403 B.n402 10.6151
R2092 B.n403 B.n154 10.6151
R2093 B.n407 B.n154 10.6151
R2094 B.n408 B.n407 10.6151
R2095 B.n409 B.n408 10.6151
R2096 B.n409 B.n152 10.6151
R2097 B.n413 B.n152 10.6151
R2098 B.n414 B.n413 10.6151
R2099 B.n415 B.n414 10.6151
R2100 B.n415 B.n150 10.6151
R2101 B.n419 B.n150 10.6151
R2102 B.n420 B.n419 10.6151
R2103 B.n421 B.n420 10.6151
R2104 B.n421 B.n148 10.6151
R2105 B.n425 B.n148 10.6151
R2106 B.n426 B.n425 10.6151
R2107 B.n427 B.n426 10.6151
R2108 B.n427 B.n146 10.6151
R2109 B.n431 B.n146 10.6151
R2110 B.n432 B.n431 10.6151
R2111 B.n433 B.n432 10.6151
R2112 B.n433 B.n144 10.6151
R2113 B.n437 B.n144 10.6151
R2114 B.n438 B.n437 10.6151
R2115 B.n439 B.n438 10.6151
R2116 B.n439 B.n142 10.6151
R2117 B.n443 B.n142 10.6151
R2118 B.n444 B.n443 10.6151
R2119 B.n445 B.n444 10.6151
R2120 B.n445 B.n140 10.6151
R2121 B.n449 B.n140 10.6151
R2122 B.n450 B.n449 10.6151
R2123 B.n451 B.n450 10.6151
R2124 B.n451 B.n138 10.6151
R2125 B.n455 B.n138 10.6151
R2126 B.n456 B.n455 10.6151
R2127 B.n457 B.n456 10.6151
R2128 B.n457 B.n136 10.6151
R2129 B.n461 B.n136 10.6151
R2130 B.n289 B.n288 10.6151
R2131 B.n288 B.n287 10.6151
R2132 B.n287 B.n198 10.6151
R2133 B.n283 B.n198 10.6151
R2134 B.n283 B.n282 10.6151
R2135 B.n282 B.n281 10.6151
R2136 B.n281 B.n200 10.6151
R2137 B.n277 B.n200 10.6151
R2138 B.n277 B.n276 10.6151
R2139 B.n276 B.n275 10.6151
R2140 B.n275 B.n202 10.6151
R2141 B.n271 B.n202 10.6151
R2142 B.n271 B.n270 10.6151
R2143 B.n270 B.n269 10.6151
R2144 B.n269 B.n204 10.6151
R2145 B.n265 B.n204 10.6151
R2146 B.n265 B.n264 10.6151
R2147 B.n264 B.n263 10.6151
R2148 B.n263 B.n206 10.6151
R2149 B.n259 B.n206 10.6151
R2150 B.n259 B.n258 10.6151
R2151 B.n258 B.n257 10.6151
R2152 B.n257 B.n208 10.6151
R2153 B.n253 B.n208 10.6151
R2154 B.n253 B.n252 10.6151
R2155 B.n252 B.n251 10.6151
R2156 B.n251 B.n210 10.6151
R2157 B.n247 B.n210 10.6151
R2158 B.n247 B.n246 10.6151
R2159 B.n246 B.n245 10.6151
R2160 B.n245 B.n212 10.6151
R2161 B.n241 B.n212 10.6151
R2162 B.n241 B.n240 10.6151
R2163 B.n240 B.n239 10.6151
R2164 B.n239 B.n214 10.6151
R2165 B.n235 B.n214 10.6151
R2166 B.n235 B.n234 10.6151
R2167 B.n234 B.n233 10.6151
R2168 B.n233 B.n216 10.6151
R2169 B.n229 B.n216 10.6151
R2170 B.n229 B.n228 10.6151
R2171 B.n228 B.n227 10.6151
R2172 B.n227 B.n218 10.6151
R2173 B.n223 B.n218 10.6151
R2174 B.n223 B.n222 10.6151
R2175 B.n222 B.n221 10.6151
R2176 B.n221 B.n0 10.6151
R2177 B.n847 B.n1 10.6151
R2178 B.n847 B.n846 10.6151
R2179 B.n846 B.n845 10.6151
R2180 B.n845 B.n4 10.6151
R2181 B.n841 B.n4 10.6151
R2182 B.n841 B.n840 10.6151
R2183 B.n840 B.n839 10.6151
R2184 B.n839 B.n6 10.6151
R2185 B.n835 B.n6 10.6151
R2186 B.n835 B.n834 10.6151
R2187 B.n834 B.n833 10.6151
R2188 B.n833 B.n8 10.6151
R2189 B.n829 B.n8 10.6151
R2190 B.n829 B.n828 10.6151
R2191 B.n828 B.n827 10.6151
R2192 B.n827 B.n10 10.6151
R2193 B.n823 B.n10 10.6151
R2194 B.n823 B.n822 10.6151
R2195 B.n822 B.n821 10.6151
R2196 B.n821 B.n12 10.6151
R2197 B.n817 B.n12 10.6151
R2198 B.n817 B.n816 10.6151
R2199 B.n816 B.n815 10.6151
R2200 B.n815 B.n14 10.6151
R2201 B.n811 B.n14 10.6151
R2202 B.n811 B.n810 10.6151
R2203 B.n810 B.n809 10.6151
R2204 B.n809 B.n16 10.6151
R2205 B.n805 B.n16 10.6151
R2206 B.n805 B.n804 10.6151
R2207 B.n804 B.n803 10.6151
R2208 B.n803 B.n18 10.6151
R2209 B.n799 B.n18 10.6151
R2210 B.n799 B.n798 10.6151
R2211 B.n798 B.n797 10.6151
R2212 B.n797 B.n20 10.6151
R2213 B.n793 B.n20 10.6151
R2214 B.n793 B.n792 10.6151
R2215 B.n792 B.n791 10.6151
R2216 B.n791 B.n22 10.6151
R2217 B.n787 B.n22 10.6151
R2218 B.n787 B.n786 10.6151
R2219 B.n786 B.n785 10.6151
R2220 B.n785 B.n24 10.6151
R2221 B.n781 B.n24 10.6151
R2222 B.n781 B.n780 10.6151
R2223 B.n780 B.n779 10.6151
R2224 B.n698 B.n54 6.5566
R2225 B.n686 B.n685 6.5566
R2226 B.n370 B.n170 6.5566
R2227 B.n383 B.n382 6.5566
R2228 B.n701 B.n54 4.05904
R2229 B.n685 B.n684 4.05904
R2230 B.n367 B.n170 4.05904
R2231 B.n384 B.n383 4.05904
R2232 B.n851 B.n0 2.81026
R2233 B.n851 B.n1 2.81026
R2234 VN.n8 VN.t0 225.292
R2235 VN.n41 VN.t2 225.292
R2236 VN.n16 VN.t8 193.175
R2237 VN.n7 VN.t9 193.175
R2238 VN.n23 VN.t6 193.175
R2239 VN.n31 VN.t7 193.175
R2240 VN.n49 VN.t5 193.175
R2241 VN.n40 VN.t1 193.175
R2242 VN.n56 VN.t3 193.175
R2243 VN.n64 VN.t4 193.175
R2244 VN.n32 VN.n31 184.788
R2245 VN.n65 VN.n64 184.788
R2246 VN.n63 VN.n33 161.3
R2247 VN.n62 VN.n61 161.3
R2248 VN.n60 VN.n34 161.3
R2249 VN.n59 VN.n58 161.3
R2250 VN.n57 VN.n35 161.3
R2251 VN.n55 VN.n54 161.3
R2252 VN.n53 VN.n36 161.3
R2253 VN.n52 VN.n51 161.3
R2254 VN.n50 VN.n37 161.3
R2255 VN.n49 VN.n48 161.3
R2256 VN.n47 VN.n38 161.3
R2257 VN.n46 VN.n45 161.3
R2258 VN.n44 VN.n39 161.3
R2259 VN.n43 VN.n42 161.3
R2260 VN.n30 VN.n0 161.3
R2261 VN.n29 VN.n28 161.3
R2262 VN.n27 VN.n1 161.3
R2263 VN.n26 VN.n25 161.3
R2264 VN.n24 VN.n2 161.3
R2265 VN.n22 VN.n21 161.3
R2266 VN.n20 VN.n3 161.3
R2267 VN.n19 VN.n18 161.3
R2268 VN.n17 VN.n4 161.3
R2269 VN.n16 VN.n15 161.3
R2270 VN.n14 VN.n5 161.3
R2271 VN.n13 VN.n12 161.3
R2272 VN.n11 VN.n6 161.3
R2273 VN.n10 VN.n9 161.3
R2274 VN.n8 VN.n7 57.3879
R2275 VN.n41 VN.n40 57.3879
R2276 VN.n12 VN.n11 53.1199
R2277 VN.n18 VN.n3 53.1199
R2278 VN.n45 VN.n44 53.1199
R2279 VN.n51 VN.n36 53.1199
R2280 VN VN.n65 52.3736
R2281 VN.n25 VN.n1 51.1773
R2282 VN.n58 VN.n34 51.1773
R2283 VN.n29 VN.n1 29.8095
R2284 VN.n62 VN.n34 29.8095
R2285 VN.n12 VN.n5 27.8669
R2286 VN.n18 VN.n17 27.8669
R2287 VN.n45 VN.n38 27.8669
R2288 VN.n51 VN.n50 27.8669
R2289 VN.n11 VN.n10 24.4675
R2290 VN.n16 VN.n5 24.4675
R2291 VN.n17 VN.n16 24.4675
R2292 VN.n22 VN.n3 24.4675
R2293 VN.n25 VN.n24 24.4675
R2294 VN.n30 VN.n29 24.4675
R2295 VN.n44 VN.n43 24.4675
R2296 VN.n50 VN.n49 24.4675
R2297 VN.n49 VN.n38 24.4675
R2298 VN.n58 VN.n57 24.4675
R2299 VN.n55 VN.n36 24.4675
R2300 VN.n63 VN.n62 24.4675
R2301 VN.n10 VN.n7 12.7233
R2302 VN.n23 VN.n22 12.7233
R2303 VN.n43 VN.n40 12.7233
R2304 VN.n56 VN.n55 12.7233
R2305 VN.n42 VN.n41 12.5492
R2306 VN.n9 VN.n8 12.5492
R2307 VN.n24 VN.n23 11.7447
R2308 VN.n57 VN.n56 11.7447
R2309 VN.n31 VN.n30 0.97918
R2310 VN.n64 VN.n63 0.97918
R2311 VN.n65 VN.n33 0.189894
R2312 VN.n61 VN.n33 0.189894
R2313 VN.n61 VN.n60 0.189894
R2314 VN.n60 VN.n59 0.189894
R2315 VN.n59 VN.n35 0.189894
R2316 VN.n54 VN.n35 0.189894
R2317 VN.n54 VN.n53 0.189894
R2318 VN.n53 VN.n52 0.189894
R2319 VN.n52 VN.n37 0.189894
R2320 VN.n48 VN.n37 0.189894
R2321 VN.n48 VN.n47 0.189894
R2322 VN.n47 VN.n46 0.189894
R2323 VN.n46 VN.n39 0.189894
R2324 VN.n42 VN.n39 0.189894
R2325 VN.n9 VN.n6 0.189894
R2326 VN.n13 VN.n6 0.189894
R2327 VN.n14 VN.n13 0.189894
R2328 VN.n15 VN.n14 0.189894
R2329 VN.n15 VN.n4 0.189894
R2330 VN.n19 VN.n4 0.189894
R2331 VN.n20 VN.n19 0.189894
R2332 VN.n21 VN.n20 0.189894
R2333 VN.n21 VN.n2 0.189894
R2334 VN.n26 VN.n2 0.189894
R2335 VN.n27 VN.n26 0.189894
R2336 VN.n28 VN.n27 0.189894
R2337 VN.n28 VN.n0 0.189894
R2338 VN.n32 VN.n0 0.189894
R2339 VN VN.n32 0.0516364
R2340 VDD2.n169 VDD2.n89 756.745
R2341 VDD2.n80 VDD2.n0 756.745
R2342 VDD2.n170 VDD2.n169 585
R2343 VDD2.n168 VDD2.n167 585
R2344 VDD2.n93 VDD2.n92 585
R2345 VDD2.n97 VDD2.n95 585
R2346 VDD2.n162 VDD2.n161 585
R2347 VDD2.n160 VDD2.n159 585
R2348 VDD2.n99 VDD2.n98 585
R2349 VDD2.n154 VDD2.n153 585
R2350 VDD2.n152 VDD2.n151 585
R2351 VDD2.n103 VDD2.n102 585
R2352 VDD2.n146 VDD2.n145 585
R2353 VDD2.n144 VDD2.n143 585
R2354 VDD2.n107 VDD2.n106 585
R2355 VDD2.n138 VDD2.n137 585
R2356 VDD2.n136 VDD2.n135 585
R2357 VDD2.n111 VDD2.n110 585
R2358 VDD2.n130 VDD2.n129 585
R2359 VDD2.n128 VDD2.n127 585
R2360 VDD2.n115 VDD2.n114 585
R2361 VDD2.n122 VDD2.n121 585
R2362 VDD2.n120 VDD2.n119 585
R2363 VDD2.n29 VDD2.n28 585
R2364 VDD2.n31 VDD2.n30 585
R2365 VDD2.n24 VDD2.n23 585
R2366 VDD2.n37 VDD2.n36 585
R2367 VDD2.n39 VDD2.n38 585
R2368 VDD2.n20 VDD2.n19 585
R2369 VDD2.n45 VDD2.n44 585
R2370 VDD2.n47 VDD2.n46 585
R2371 VDD2.n16 VDD2.n15 585
R2372 VDD2.n53 VDD2.n52 585
R2373 VDD2.n55 VDD2.n54 585
R2374 VDD2.n12 VDD2.n11 585
R2375 VDD2.n61 VDD2.n60 585
R2376 VDD2.n63 VDD2.n62 585
R2377 VDD2.n8 VDD2.n7 585
R2378 VDD2.n70 VDD2.n69 585
R2379 VDD2.n71 VDD2.n6 585
R2380 VDD2.n73 VDD2.n72 585
R2381 VDD2.n4 VDD2.n3 585
R2382 VDD2.n79 VDD2.n78 585
R2383 VDD2.n81 VDD2.n80 585
R2384 VDD2.n118 VDD2.t5 327.466
R2385 VDD2.n27 VDD2.t9 327.466
R2386 VDD2.n169 VDD2.n168 171.744
R2387 VDD2.n168 VDD2.n92 171.744
R2388 VDD2.n97 VDD2.n92 171.744
R2389 VDD2.n161 VDD2.n97 171.744
R2390 VDD2.n161 VDD2.n160 171.744
R2391 VDD2.n160 VDD2.n98 171.744
R2392 VDD2.n153 VDD2.n98 171.744
R2393 VDD2.n153 VDD2.n152 171.744
R2394 VDD2.n152 VDD2.n102 171.744
R2395 VDD2.n145 VDD2.n102 171.744
R2396 VDD2.n145 VDD2.n144 171.744
R2397 VDD2.n144 VDD2.n106 171.744
R2398 VDD2.n137 VDD2.n106 171.744
R2399 VDD2.n137 VDD2.n136 171.744
R2400 VDD2.n136 VDD2.n110 171.744
R2401 VDD2.n129 VDD2.n110 171.744
R2402 VDD2.n129 VDD2.n128 171.744
R2403 VDD2.n128 VDD2.n114 171.744
R2404 VDD2.n121 VDD2.n114 171.744
R2405 VDD2.n121 VDD2.n120 171.744
R2406 VDD2.n30 VDD2.n29 171.744
R2407 VDD2.n30 VDD2.n23 171.744
R2408 VDD2.n37 VDD2.n23 171.744
R2409 VDD2.n38 VDD2.n37 171.744
R2410 VDD2.n38 VDD2.n19 171.744
R2411 VDD2.n45 VDD2.n19 171.744
R2412 VDD2.n46 VDD2.n45 171.744
R2413 VDD2.n46 VDD2.n15 171.744
R2414 VDD2.n53 VDD2.n15 171.744
R2415 VDD2.n54 VDD2.n53 171.744
R2416 VDD2.n54 VDD2.n11 171.744
R2417 VDD2.n61 VDD2.n11 171.744
R2418 VDD2.n62 VDD2.n61 171.744
R2419 VDD2.n62 VDD2.n7 171.744
R2420 VDD2.n70 VDD2.n7 171.744
R2421 VDD2.n71 VDD2.n70 171.744
R2422 VDD2.n72 VDD2.n71 171.744
R2423 VDD2.n72 VDD2.n3 171.744
R2424 VDD2.n79 VDD2.n3 171.744
R2425 VDD2.n80 VDD2.n79 171.744
R2426 VDD2.n120 VDD2.t5 85.8723
R2427 VDD2.n29 VDD2.t9 85.8723
R2428 VDD2.n88 VDD2.n87 73.7972
R2429 VDD2 VDD2.n177 73.7943
R2430 VDD2.n176 VDD2.n175 72.3915
R2431 VDD2.n86 VDD2.n85 72.3913
R2432 VDD2.n86 VDD2.n84 52.9457
R2433 VDD2.n174 VDD2.n173 50.9975
R2434 VDD2.n174 VDD2.n88 46.3058
R2435 VDD2.n119 VDD2.n118 16.3895
R2436 VDD2.n28 VDD2.n27 16.3895
R2437 VDD2.n95 VDD2.n93 13.1884
R2438 VDD2.n73 VDD2.n4 13.1884
R2439 VDD2.n167 VDD2.n166 12.8005
R2440 VDD2.n163 VDD2.n162 12.8005
R2441 VDD2.n122 VDD2.n117 12.8005
R2442 VDD2.n31 VDD2.n26 12.8005
R2443 VDD2.n74 VDD2.n6 12.8005
R2444 VDD2.n78 VDD2.n77 12.8005
R2445 VDD2.n170 VDD2.n91 12.0247
R2446 VDD2.n159 VDD2.n96 12.0247
R2447 VDD2.n123 VDD2.n115 12.0247
R2448 VDD2.n32 VDD2.n24 12.0247
R2449 VDD2.n69 VDD2.n68 12.0247
R2450 VDD2.n81 VDD2.n2 12.0247
R2451 VDD2.n171 VDD2.n89 11.249
R2452 VDD2.n158 VDD2.n99 11.249
R2453 VDD2.n127 VDD2.n126 11.249
R2454 VDD2.n36 VDD2.n35 11.249
R2455 VDD2.n67 VDD2.n8 11.249
R2456 VDD2.n82 VDD2.n0 11.249
R2457 VDD2.n155 VDD2.n154 10.4732
R2458 VDD2.n130 VDD2.n113 10.4732
R2459 VDD2.n39 VDD2.n22 10.4732
R2460 VDD2.n64 VDD2.n63 10.4732
R2461 VDD2.n151 VDD2.n101 9.69747
R2462 VDD2.n131 VDD2.n111 9.69747
R2463 VDD2.n40 VDD2.n20 9.69747
R2464 VDD2.n60 VDD2.n10 9.69747
R2465 VDD2.n173 VDD2.n172 9.45567
R2466 VDD2.n84 VDD2.n83 9.45567
R2467 VDD2.n105 VDD2.n104 9.3005
R2468 VDD2.n148 VDD2.n147 9.3005
R2469 VDD2.n150 VDD2.n149 9.3005
R2470 VDD2.n101 VDD2.n100 9.3005
R2471 VDD2.n156 VDD2.n155 9.3005
R2472 VDD2.n158 VDD2.n157 9.3005
R2473 VDD2.n96 VDD2.n94 9.3005
R2474 VDD2.n164 VDD2.n163 9.3005
R2475 VDD2.n172 VDD2.n171 9.3005
R2476 VDD2.n91 VDD2.n90 9.3005
R2477 VDD2.n166 VDD2.n165 9.3005
R2478 VDD2.n142 VDD2.n141 9.3005
R2479 VDD2.n140 VDD2.n139 9.3005
R2480 VDD2.n109 VDD2.n108 9.3005
R2481 VDD2.n134 VDD2.n133 9.3005
R2482 VDD2.n132 VDD2.n131 9.3005
R2483 VDD2.n113 VDD2.n112 9.3005
R2484 VDD2.n126 VDD2.n125 9.3005
R2485 VDD2.n124 VDD2.n123 9.3005
R2486 VDD2.n117 VDD2.n116 9.3005
R2487 VDD2.n83 VDD2.n82 9.3005
R2488 VDD2.n2 VDD2.n1 9.3005
R2489 VDD2.n77 VDD2.n76 9.3005
R2490 VDD2.n49 VDD2.n48 9.3005
R2491 VDD2.n18 VDD2.n17 9.3005
R2492 VDD2.n43 VDD2.n42 9.3005
R2493 VDD2.n41 VDD2.n40 9.3005
R2494 VDD2.n22 VDD2.n21 9.3005
R2495 VDD2.n35 VDD2.n34 9.3005
R2496 VDD2.n33 VDD2.n32 9.3005
R2497 VDD2.n26 VDD2.n25 9.3005
R2498 VDD2.n51 VDD2.n50 9.3005
R2499 VDD2.n14 VDD2.n13 9.3005
R2500 VDD2.n57 VDD2.n56 9.3005
R2501 VDD2.n59 VDD2.n58 9.3005
R2502 VDD2.n10 VDD2.n9 9.3005
R2503 VDD2.n65 VDD2.n64 9.3005
R2504 VDD2.n67 VDD2.n66 9.3005
R2505 VDD2.n68 VDD2.n5 9.3005
R2506 VDD2.n75 VDD2.n74 9.3005
R2507 VDD2.n150 VDD2.n103 8.92171
R2508 VDD2.n135 VDD2.n134 8.92171
R2509 VDD2.n44 VDD2.n43 8.92171
R2510 VDD2.n59 VDD2.n12 8.92171
R2511 VDD2.n147 VDD2.n146 8.14595
R2512 VDD2.n138 VDD2.n109 8.14595
R2513 VDD2.n47 VDD2.n18 8.14595
R2514 VDD2.n56 VDD2.n55 8.14595
R2515 VDD2.n143 VDD2.n105 7.3702
R2516 VDD2.n139 VDD2.n107 7.3702
R2517 VDD2.n48 VDD2.n16 7.3702
R2518 VDD2.n52 VDD2.n14 7.3702
R2519 VDD2.n143 VDD2.n142 6.59444
R2520 VDD2.n142 VDD2.n107 6.59444
R2521 VDD2.n51 VDD2.n16 6.59444
R2522 VDD2.n52 VDD2.n51 6.59444
R2523 VDD2.n146 VDD2.n105 5.81868
R2524 VDD2.n139 VDD2.n138 5.81868
R2525 VDD2.n48 VDD2.n47 5.81868
R2526 VDD2.n55 VDD2.n14 5.81868
R2527 VDD2.n147 VDD2.n103 5.04292
R2528 VDD2.n135 VDD2.n109 5.04292
R2529 VDD2.n44 VDD2.n18 5.04292
R2530 VDD2.n56 VDD2.n12 5.04292
R2531 VDD2.n151 VDD2.n150 4.26717
R2532 VDD2.n134 VDD2.n111 4.26717
R2533 VDD2.n43 VDD2.n20 4.26717
R2534 VDD2.n60 VDD2.n59 4.26717
R2535 VDD2.n118 VDD2.n116 3.70982
R2536 VDD2.n27 VDD2.n25 3.70982
R2537 VDD2.n154 VDD2.n101 3.49141
R2538 VDD2.n131 VDD2.n130 3.49141
R2539 VDD2.n40 VDD2.n39 3.49141
R2540 VDD2.n63 VDD2.n10 3.49141
R2541 VDD2.n173 VDD2.n89 2.71565
R2542 VDD2.n155 VDD2.n99 2.71565
R2543 VDD2.n127 VDD2.n113 2.71565
R2544 VDD2.n36 VDD2.n22 2.71565
R2545 VDD2.n64 VDD2.n8 2.71565
R2546 VDD2.n84 VDD2.n0 2.71565
R2547 VDD2.n177 VDD2.t8 2.10166
R2548 VDD2.n177 VDD2.t7 2.10166
R2549 VDD2.n175 VDD2.t6 2.10166
R2550 VDD2.n175 VDD2.t4 2.10166
R2551 VDD2.n87 VDD2.t3 2.10166
R2552 VDD2.n87 VDD2.t2 2.10166
R2553 VDD2.n85 VDD2.t0 2.10166
R2554 VDD2.n85 VDD2.t1 2.10166
R2555 VDD2.n176 VDD2.n174 1.94878
R2556 VDD2.n171 VDD2.n170 1.93989
R2557 VDD2.n159 VDD2.n158 1.93989
R2558 VDD2.n126 VDD2.n115 1.93989
R2559 VDD2.n35 VDD2.n24 1.93989
R2560 VDD2.n69 VDD2.n67 1.93989
R2561 VDD2.n82 VDD2.n81 1.93989
R2562 VDD2.n167 VDD2.n91 1.16414
R2563 VDD2.n162 VDD2.n96 1.16414
R2564 VDD2.n123 VDD2.n122 1.16414
R2565 VDD2.n32 VDD2.n31 1.16414
R2566 VDD2.n68 VDD2.n6 1.16414
R2567 VDD2.n78 VDD2.n2 1.16414
R2568 VDD2 VDD2.n176 0.545759
R2569 VDD2.n88 VDD2.n86 0.432223
R2570 VDD2.n166 VDD2.n93 0.388379
R2571 VDD2.n163 VDD2.n95 0.388379
R2572 VDD2.n119 VDD2.n117 0.388379
R2573 VDD2.n28 VDD2.n26 0.388379
R2574 VDD2.n74 VDD2.n73 0.388379
R2575 VDD2.n77 VDD2.n4 0.388379
R2576 VDD2.n172 VDD2.n90 0.155672
R2577 VDD2.n165 VDD2.n90 0.155672
R2578 VDD2.n165 VDD2.n164 0.155672
R2579 VDD2.n164 VDD2.n94 0.155672
R2580 VDD2.n157 VDD2.n94 0.155672
R2581 VDD2.n157 VDD2.n156 0.155672
R2582 VDD2.n156 VDD2.n100 0.155672
R2583 VDD2.n149 VDD2.n100 0.155672
R2584 VDD2.n149 VDD2.n148 0.155672
R2585 VDD2.n148 VDD2.n104 0.155672
R2586 VDD2.n141 VDD2.n104 0.155672
R2587 VDD2.n141 VDD2.n140 0.155672
R2588 VDD2.n140 VDD2.n108 0.155672
R2589 VDD2.n133 VDD2.n108 0.155672
R2590 VDD2.n133 VDD2.n132 0.155672
R2591 VDD2.n132 VDD2.n112 0.155672
R2592 VDD2.n125 VDD2.n112 0.155672
R2593 VDD2.n125 VDD2.n124 0.155672
R2594 VDD2.n124 VDD2.n116 0.155672
R2595 VDD2.n33 VDD2.n25 0.155672
R2596 VDD2.n34 VDD2.n33 0.155672
R2597 VDD2.n34 VDD2.n21 0.155672
R2598 VDD2.n41 VDD2.n21 0.155672
R2599 VDD2.n42 VDD2.n41 0.155672
R2600 VDD2.n42 VDD2.n17 0.155672
R2601 VDD2.n49 VDD2.n17 0.155672
R2602 VDD2.n50 VDD2.n49 0.155672
R2603 VDD2.n50 VDD2.n13 0.155672
R2604 VDD2.n57 VDD2.n13 0.155672
R2605 VDD2.n58 VDD2.n57 0.155672
R2606 VDD2.n58 VDD2.n9 0.155672
R2607 VDD2.n65 VDD2.n9 0.155672
R2608 VDD2.n66 VDD2.n65 0.155672
R2609 VDD2.n66 VDD2.n5 0.155672
R2610 VDD2.n75 VDD2.n5 0.155672
R2611 VDD2.n76 VDD2.n75 0.155672
R2612 VDD2.n76 VDD2.n1 0.155672
R2613 VDD2.n83 VDD2.n1 0.155672
C0 VTAIL VDD1 12.349401f
C1 w_n3682_n4062# VN 7.73309f
C2 VDD1 VN 0.151799f
C3 VTAIL VP 12.9342f
C4 VDD1 w_n3682_n4062# 2.77803f
C5 VP VN 8.05232f
C6 w_n3682_n4062# VP 8.210401f
C7 VTAIL B 4.16823f
C8 VDD1 VP 13.0429f
C9 VDD2 VTAIL 12.393901f
C10 B VN 1.1536f
C11 w_n3682_n4062# B 10.3931f
C12 VDD2 VN 12.700901f
C13 VDD1 B 2.48463f
C14 VDD2 w_n3682_n4062# 2.88685f
C15 VDD2 VDD1 1.73888f
C16 B VP 1.95253f
C17 VDD2 VP 0.498464f
C18 VDD2 B 2.57645f
C19 VTAIL VN 12.9198f
C20 VTAIL w_n3682_n4062# 3.62242f
C21 VDD2 VSUBS 1.963058f
C22 VDD1 VSUBS 1.773705f
C23 VTAIL VSUBS 1.262897f
C24 VN VSUBS 6.73984f
C25 VP VSUBS 3.496182f
C26 B VSUBS 4.827605f
C27 w_n3682_n4062# VSUBS 0.183319p
C28 VDD2.n0 VSUBS 0.028942f
C29 VDD2.n1 VSUBS 0.026962f
C30 VDD2.n2 VSUBS 0.014488f
C31 VDD2.n3 VSUBS 0.034245f
C32 VDD2.n4 VSUBS 0.014914f
C33 VDD2.n5 VSUBS 0.026962f
C34 VDD2.n6 VSUBS 0.015341f
C35 VDD2.n7 VSUBS 0.034245f
C36 VDD2.n8 VSUBS 0.015341f
C37 VDD2.n9 VSUBS 0.026962f
C38 VDD2.n10 VSUBS 0.014488f
C39 VDD2.n11 VSUBS 0.034245f
C40 VDD2.n12 VSUBS 0.015341f
C41 VDD2.n13 VSUBS 0.026962f
C42 VDD2.n14 VSUBS 0.014488f
C43 VDD2.n15 VSUBS 0.034245f
C44 VDD2.n16 VSUBS 0.015341f
C45 VDD2.n17 VSUBS 0.026962f
C46 VDD2.n18 VSUBS 0.014488f
C47 VDD2.n19 VSUBS 0.034245f
C48 VDD2.n20 VSUBS 0.015341f
C49 VDD2.n21 VSUBS 0.026962f
C50 VDD2.n22 VSUBS 0.014488f
C51 VDD2.n23 VSUBS 0.034245f
C52 VDD2.n24 VSUBS 0.015341f
C53 VDD2.n25 VSUBS 1.77913f
C54 VDD2.n26 VSUBS 0.014488f
C55 VDD2.t9 VSUBS 0.073344f
C56 VDD2.n27 VSUBS 0.193799f
C57 VDD2.n28 VSUBS 0.021785f
C58 VDD2.n29 VSUBS 0.025684f
C59 VDD2.n30 VSUBS 0.034245f
C60 VDD2.n31 VSUBS 0.015341f
C61 VDD2.n32 VSUBS 0.014488f
C62 VDD2.n33 VSUBS 0.026962f
C63 VDD2.n34 VSUBS 0.026962f
C64 VDD2.n35 VSUBS 0.014488f
C65 VDD2.n36 VSUBS 0.015341f
C66 VDD2.n37 VSUBS 0.034245f
C67 VDD2.n38 VSUBS 0.034245f
C68 VDD2.n39 VSUBS 0.015341f
C69 VDD2.n40 VSUBS 0.014488f
C70 VDD2.n41 VSUBS 0.026962f
C71 VDD2.n42 VSUBS 0.026962f
C72 VDD2.n43 VSUBS 0.014488f
C73 VDD2.n44 VSUBS 0.015341f
C74 VDD2.n45 VSUBS 0.034245f
C75 VDD2.n46 VSUBS 0.034245f
C76 VDD2.n47 VSUBS 0.015341f
C77 VDD2.n48 VSUBS 0.014488f
C78 VDD2.n49 VSUBS 0.026962f
C79 VDD2.n50 VSUBS 0.026962f
C80 VDD2.n51 VSUBS 0.014488f
C81 VDD2.n52 VSUBS 0.015341f
C82 VDD2.n53 VSUBS 0.034245f
C83 VDD2.n54 VSUBS 0.034245f
C84 VDD2.n55 VSUBS 0.015341f
C85 VDD2.n56 VSUBS 0.014488f
C86 VDD2.n57 VSUBS 0.026962f
C87 VDD2.n58 VSUBS 0.026962f
C88 VDD2.n59 VSUBS 0.014488f
C89 VDD2.n60 VSUBS 0.015341f
C90 VDD2.n61 VSUBS 0.034245f
C91 VDD2.n62 VSUBS 0.034245f
C92 VDD2.n63 VSUBS 0.015341f
C93 VDD2.n64 VSUBS 0.014488f
C94 VDD2.n65 VSUBS 0.026962f
C95 VDD2.n66 VSUBS 0.026962f
C96 VDD2.n67 VSUBS 0.014488f
C97 VDD2.n68 VSUBS 0.014488f
C98 VDD2.n69 VSUBS 0.015341f
C99 VDD2.n70 VSUBS 0.034245f
C100 VDD2.n71 VSUBS 0.034245f
C101 VDD2.n72 VSUBS 0.034245f
C102 VDD2.n73 VSUBS 0.014914f
C103 VDD2.n74 VSUBS 0.014488f
C104 VDD2.n75 VSUBS 0.026962f
C105 VDD2.n76 VSUBS 0.026962f
C106 VDD2.n77 VSUBS 0.014488f
C107 VDD2.n78 VSUBS 0.015341f
C108 VDD2.n79 VSUBS 0.034245f
C109 VDD2.n80 VSUBS 0.080573f
C110 VDD2.n81 VSUBS 0.015341f
C111 VDD2.n82 VSUBS 0.014488f
C112 VDD2.n83 VSUBS 0.066374f
C113 VDD2.n84 VSUBS 0.067349f
C114 VDD2.t0 VSUBS 0.329611f
C115 VDD2.t1 VSUBS 0.329611f
C116 VDD2.n85 VSUBS 2.69431f
C117 VDD2.n86 VSUBS 0.934089f
C118 VDD2.t3 VSUBS 0.329611f
C119 VDD2.t2 VSUBS 0.329611f
C120 VDD2.n87 VSUBS 2.70981f
C121 VDD2.n88 VSUBS 3.2718f
C122 VDD2.n89 VSUBS 0.028942f
C123 VDD2.n90 VSUBS 0.026962f
C124 VDD2.n91 VSUBS 0.014488f
C125 VDD2.n92 VSUBS 0.034245f
C126 VDD2.n93 VSUBS 0.014914f
C127 VDD2.n94 VSUBS 0.026962f
C128 VDD2.n95 VSUBS 0.014914f
C129 VDD2.n96 VSUBS 0.014488f
C130 VDD2.n97 VSUBS 0.034245f
C131 VDD2.n98 VSUBS 0.034245f
C132 VDD2.n99 VSUBS 0.015341f
C133 VDD2.n100 VSUBS 0.026962f
C134 VDD2.n101 VSUBS 0.014488f
C135 VDD2.n102 VSUBS 0.034245f
C136 VDD2.n103 VSUBS 0.015341f
C137 VDD2.n104 VSUBS 0.026962f
C138 VDD2.n105 VSUBS 0.014488f
C139 VDD2.n106 VSUBS 0.034245f
C140 VDD2.n107 VSUBS 0.015341f
C141 VDD2.n108 VSUBS 0.026962f
C142 VDD2.n109 VSUBS 0.014488f
C143 VDD2.n110 VSUBS 0.034245f
C144 VDD2.n111 VSUBS 0.015341f
C145 VDD2.n112 VSUBS 0.026962f
C146 VDD2.n113 VSUBS 0.014488f
C147 VDD2.n114 VSUBS 0.034245f
C148 VDD2.n115 VSUBS 0.015341f
C149 VDD2.n116 VSUBS 1.77913f
C150 VDD2.n117 VSUBS 0.014488f
C151 VDD2.t5 VSUBS 0.073344f
C152 VDD2.n118 VSUBS 0.193799f
C153 VDD2.n119 VSUBS 0.021785f
C154 VDD2.n120 VSUBS 0.025684f
C155 VDD2.n121 VSUBS 0.034245f
C156 VDD2.n122 VSUBS 0.015341f
C157 VDD2.n123 VSUBS 0.014488f
C158 VDD2.n124 VSUBS 0.026962f
C159 VDD2.n125 VSUBS 0.026962f
C160 VDD2.n126 VSUBS 0.014488f
C161 VDD2.n127 VSUBS 0.015341f
C162 VDD2.n128 VSUBS 0.034245f
C163 VDD2.n129 VSUBS 0.034245f
C164 VDD2.n130 VSUBS 0.015341f
C165 VDD2.n131 VSUBS 0.014488f
C166 VDD2.n132 VSUBS 0.026962f
C167 VDD2.n133 VSUBS 0.026962f
C168 VDD2.n134 VSUBS 0.014488f
C169 VDD2.n135 VSUBS 0.015341f
C170 VDD2.n136 VSUBS 0.034245f
C171 VDD2.n137 VSUBS 0.034245f
C172 VDD2.n138 VSUBS 0.015341f
C173 VDD2.n139 VSUBS 0.014488f
C174 VDD2.n140 VSUBS 0.026962f
C175 VDD2.n141 VSUBS 0.026962f
C176 VDD2.n142 VSUBS 0.014488f
C177 VDD2.n143 VSUBS 0.015341f
C178 VDD2.n144 VSUBS 0.034245f
C179 VDD2.n145 VSUBS 0.034245f
C180 VDD2.n146 VSUBS 0.015341f
C181 VDD2.n147 VSUBS 0.014488f
C182 VDD2.n148 VSUBS 0.026962f
C183 VDD2.n149 VSUBS 0.026962f
C184 VDD2.n150 VSUBS 0.014488f
C185 VDD2.n151 VSUBS 0.015341f
C186 VDD2.n152 VSUBS 0.034245f
C187 VDD2.n153 VSUBS 0.034245f
C188 VDD2.n154 VSUBS 0.015341f
C189 VDD2.n155 VSUBS 0.014488f
C190 VDD2.n156 VSUBS 0.026962f
C191 VDD2.n157 VSUBS 0.026962f
C192 VDD2.n158 VSUBS 0.014488f
C193 VDD2.n159 VSUBS 0.015341f
C194 VDD2.n160 VSUBS 0.034245f
C195 VDD2.n161 VSUBS 0.034245f
C196 VDD2.n162 VSUBS 0.015341f
C197 VDD2.n163 VSUBS 0.014488f
C198 VDD2.n164 VSUBS 0.026962f
C199 VDD2.n165 VSUBS 0.026962f
C200 VDD2.n166 VSUBS 0.014488f
C201 VDD2.n167 VSUBS 0.015341f
C202 VDD2.n168 VSUBS 0.034245f
C203 VDD2.n169 VSUBS 0.080573f
C204 VDD2.n170 VSUBS 0.015341f
C205 VDD2.n171 VSUBS 0.014488f
C206 VDD2.n172 VSUBS 0.066374f
C207 VDD2.n173 VSUBS 0.059124f
C208 VDD2.n174 VSUBS 3.12622f
C209 VDD2.t6 VSUBS 0.329611f
C210 VDD2.t4 VSUBS 0.329611f
C211 VDD2.n175 VSUBS 2.69432f
C212 VDD2.n176 VSUBS 0.727216f
C213 VDD2.t8 VSUBS 0.329611f
C214 VDD2.t7 VSUBS 0.329611f
C215 VDD2.n177 VSUBS 2.70976f
C216 VN.n0 VSUBS 0.031109f
C217 VN.t7 VSUBS 2.54689f
C218 VN.n1 VSUBS 0.030345f
C219 VN.n2 VSUBS 0.031109f
C220 VN.t6 VSUBS 2.54689f
C221 VN.n3 VSUBS 0.055197f
C222 VN.n4 VSUBS 0.031109f
C223 VN.t8 VSUBS 2.54689f
C224 VN.n5 VSUBS 0.06098f
C225 VN.n6 VSUBS 0.031109f
C226 VN.t9 VSUBS 2.54689f
C227 VN.n7 VSUBS 0.969482f
C228 VN.t0 VSUBS 2.69665f
C229 VN.n8 VSUBS 0.975077f
C230 VN.n9 VSUBS 0.231159f
C231 VN.n10 VSUBS 0.044239f
C232 VN.n11 VSUBS 0.055197f
C233 VN.n12 VSUBS 0.032628f
C234 VN.n13 VSUBS 0.031109f
C235 VN.n14 VSUBS 0.031109f
C236 VN.n15 VSUBS 0.031109f
C237 VN.n16 VSUBS 0.925637f
C238 VN.n17 VSUBS 0.06098f
C239 VN.n18 VSUBS 0.032628f
C240 VN.n19 VSUBS 0.031109f
C241 VN.n20 VSUBS 0.031109f
C242 VN.n21 VSUBS 0.031109f
C243 VN.n22 VSUBS 0.044239f
C244 VN.n23 VSUBS 0.896283f
C245 VN.n24 VSUBS 0.043094f
C246 VN.n25 VSUBS 0.056482f
C247 VN.n26 VSUBS 0.031109f
C248 VN.n27 VSUBS 0.031109f
C249 VN.n28 VSUBS 0.031109f
C250 VN.n29 VSUBS 0.061978f
C251 VN.n30 VSUBS 0.030499f
C252 VN.n31 VSUBS 0.969379f
C253 VN.n32 VSUBS 0.034752f
C254 VN.n33 VSUBS 0.031109f
C255 VN.t4 VSUBS 2.54689f
C256 VN.n34 VSUBS 0.030345f
C257 VN.n35 VSUBS 0.031109f
C258 VN.t3 VSUBS 2.54689f
C259 VN.n36 VSUBS 0.055197f
C260 VN.n37 VSUBS 0.031109f
C261 VN.t5 VSUBS 2.54689f
C262 VN.n38 VSUBS 0.06098f
C263 VN.n39 VSUBS 0.031109f
C264 VN.t1 VSUBS 2.54689f
C265 VN.n40 VSUBS 0.969482f
C266 VN.t2 VSUBS 2.69665f
C267 VN.n41 VSUBS 0.975077f
C268 VN.n42 VSUBS 0.231159f
C269 VN.n43 VSUBS 0.044239f
C270 VN.n44 VSUBS 0.055197f
C271 VN.n45 VSUBS 0.032628f
C272 VN.n46 VSUBS 0.031109f
C273 VN.n47 VSUBS 0.031109f
C274 VN.n48 VSUBS 0.031109f
C275 VN.n49 VSUBS 0.925637f
C276 VN.n50 VSUBS 0.06098f
C277 VN.n51 VSUBS 0.032628f
C278 VN.n52 VSUBS 0.031109f
C279 VN.n53 VSUBS 0.031109f
C280 VN.n54 VSUBS 0.031109f
C281 VN.n55 VSUBS 0.044239f
C282 VN.n56 VSUBS 0.896283f
C283 VN.n57 VSUBS 0.043094f
C284 VN.n58 VSUBS 0.056482f
C285 VN.n59 VSUBS 0.031109f
C286 VN.n60 VSUBS 0.031109f
C287 VN.n61 VSUBS 0.031109f
C288 VN.n62 VSUBS 0.061978f
C289 VN.n63 VSUBS 0.030499f
C290 VN.n64 VSUBS 0.969379f
C291 VN.n65 VSUBS 1.82345f
C292 B.n0 VSUBS 0.005179f
C293 B.n1 VSUBS 0.005179f
C294 B.n2 VSUBS 0.008191f
C295 B.n3 VSUBS 0.008191f
C296 B.n4 VSUBS 0.008191f
C297 B.n5 VSUBS 0.008191f
C298 B.n6 VSUBS 0.008191f
C299 B.n7 VSUBS 0.008191f
C300 B.n8 VSUBS 0.008191f
C301 B.n9 VSUBS 0.008191f
C302 B.n10 VSUBS 0.008191f
C303 B.n11 VSUBS 0.008191f
C304 B.n12 VSUBS 0.008191f
C305 B.n13 VSUBS 0.008191f
C306 B.n14 VSUBS 0.008191f
C307 B.n15 VSUBS 0.008191f
C308 B.n16 VSUBS 0.008191f
C309 B.n17 VSUBS 0.008191f
C310 B.n18 VSUBS 0.008191f
C311 B.n19 VSUBS 0.008191f
C312 B.n20 VSUBS 0.008191f
C313 B.n21 VSUBS 0.008191f
C314 B.n22 VSUBS 0.008191f
C315 B.n23 VSUBS 0.008191f
C316 B.n24 VSUBS 0.008191f
C317 B.n25 VSUBS 0.008191f
C318 B.n26 VSUBS 0.019869f
C319 B.n27 VSUBS 0.008191f
C320 B.n28 VSUBS 0.008191f
C321 B.n29 VSUBS 0.008191f
C322 B.n30 VSUBS 0.008191f
C323 B.n31 VSUBS 0.008191f
C324 B.n32 VSUBS 0.008191f
C325 B.n33 VSUBS 0.008191f
C326 B.n34 VSUBS 0.008191f
C327 B.n35 VSUBS 0.008191f
C328 B.n36 VSUBS 0.008191f
C329 B.n37 VSUBS 0.008191f
C330 B.n38 VSUBS 0.008191f
C331 B.n39 VSUBS 0.008191f
C332 B.n40 VSUBS 0.008191f
C333 B.n41 VSUBS 0.008191f
C334 B.n42 VSUBS 0.008191f
C335 B.n43 VSUBS 0.008191f
C336 B.n44 VSUBS 0.008191f
C337 B.n45 VSUBS 0.008191f
C338 B.n46 VSUBS 0.008191f
C339 B.n47 VSUBS 0.008191f
C340 B.n48 VSUBS 0.008191f
C341 B.n49 VSUBS 0.008191f
C342 B.n50 VSUBS 0.008191f
C343 B.n51 VSUBS 0.008191f
C344 B.t5 VSUBS 0.340084f
C345 B.t4 VSUBS 0.3704f
C346 B.t3 VSUBS 1.53091f
C347 B.n52 VSUBS 0.554709f
C348 B.n53 VSUBS 0.345042f
C349 B.n54 VSUBS 0.018977f
C350 B.n55 VSUBS 0.008191f
C351 B.n56 VSUBS 0.008191f
C352 B.n57 VSUBS 0.008191f
C353 B.n58 VSUBS 0.008191f
C354 B.n59 VSUBS 0.008191f
C355 B.t8 VSUBS 0.340088f
C356 B.t7 VSUBS 0.370404f
C357 B.t6 VSUBS 1.53091f
C358 B.n60 VSUBS 0.554705f
C359 B.n61 VSUBS 0.345039f
C360 B.n62 VSUBS 0.008191f
C361 B.n63 VSUBS 0.008191f
C362 B.n64 VSUBS 0.008191f
C363 B.n65 VSUBS 0.008191f
C364 B.n66 VSUBS 0.008191f
C365 B.n67 VSUBS 0.008191f
C366 B.n68 VSUBS 0.008191f
C367 B.n69 VSUBS 0.008191f
C368 B.n70 VSUBS 0.008191f
C369 B.n71 VSUBS 0.008191f
C370 B.n72 VSUBS 0.008191f
C371 B.n73 VSUBS 0.008191f
C372 B.n74 VSUBS 0.008191f
C373 B.n75 VSUBS 0.008191f
C374 B.n76 VSUBS 0.008191f
C375 B.n77 VSUBS 0.008191f
C376 B.n78 VSUBS 0.008191f
C377 B.n79 VSUBS 0.008191f
C378 B.n80 VSUBS 0.008191f
C379 B.n81 VSUBS 0.008191f
C380 B.n82 VSUBS 0.008191f
C381 B.n83 VSUBS 0.008191f
C382 B.n84 VSUBS 0.008191f
C383 B.n85 VSUBS 0.008191f
C384 B.n86 VSUBS 0.008191f
C385 B.n87 VSUBS 0.019157f
C386 B.n88 VSUBS 0.008191f
C387 B.n89 VSUBS 0.008191f
C388 B.n90 VSUBS 0.008191f
C389 B.n91 VSUBS 0.008191f
C390 B.n92 VSUBS 0.008191f
C391 B.n93 VSUBS 0.008191f
C392 B.n94 VSUBS 0.008191f
C393 B.n95 VSUBS 0.008191f
C394 B.n96 VSUBS 0.008191f
C395 B.n97 VSUBS 0.008191f
C396 B.n98 VSUBS 0.008191f
C397 B.n99 VSUBS 0.008191f
C398 B.n100 VSUBS 0.008191f
C399 B.n101 VSUBS 0.008191f
C400 B.n102 VSUBS 0.008191f
C401 B.n103 VSUBS 0.008191f
C402 B.n104 VSUBS 0.008191f
C403 B.n105 VSUBS 0.008191f
C404 B.n106 VSUBS 0.008191f
C405 B.n107 VSUBS 0.008191f
C406 B.n108 VSUBS 0.008191f
C407 B.n109 VSUBS 0.008191f
C408 B.n110 VSUBS 0.008191f
C409 B.n111 VSUBS 0.008191f
C410 B.n112 VSUBS 0.008191f
C411 B.n113 VSUBS 0.008191f
C412 B.n114 VSUBS 0.008191f
C413 B.n115 VSUBS 0.008191f
C414 B.n116 VSUBS 0.008191f
C415 B.n117 VSUBS 0.008191f
C416 B.n118 VSUBS 0.008191f
C417 B.n119 VSUBS 0.008191f
C418 B.n120 VSUBS 0.008191f
C419 B.n121 VSUBS 0.008191f
C420 B.n122 VSUBS 0.008191f
C421 B.n123 VSUBS 0.008191f
C422 B.n124 VSUBS 0.008191f
C423 B.n125 VSUBS 0.008191f
C424 B.n126 VSUBS 0.008191f
C425 B.n127 VSUBS 0.008191f
C426 B.n128 VSUBS 0.008191f
C427 B.n129 VSUBS 0.008191f
C428 B.n130 VSUBS 0.008191f
C429 B.n131 VSUBS 0.008191f
C430 B.n132 VSUBS 0.008191f
C431 B.n133 VSUBS 0.008191f
C432 B.n134 VSUBS 0.008191f
C433 B.n135 VSUBS 0.019157f
C434 B.n136 VSUBS 0.008191f
C435 B.n137 VSUBS 0.008191f
C436 B.n138 VSUBS 0.008191f
C437 B.n139 VSUBS 0.008191f
C438 B.n140 VSUBS 0.008191f
C439 B.n141 VSUBS 0.008191f
C440 B.n142 VSUBS 0.008191f
C441 B.n143 VSUBS 0.008191f
C442 B.n144 VSUBS 0.008191f
C443 B.n145 VSUBS 0.008191f
C444 B.n146 VSUBS 0.008191f
C445 B.n147 VSUBS 0.008191f
C446 B.n148 VSUBS 0.008191f
C447 B.n149 VSUBS 0.008191f
C448 B.n150 VSUBS 0.008191f
C449 B.n151 VSUBS 0.008191f
C450 B.n152 VSUBS 0.008191f
C451 B.n153 VSUBS 0.008191f
C452 B.n154 VSUBS 0.008191f
C453 B.n155 VSUBS 0.008191f
C454 B.n156 VSUBS 0.008191f
C455 B.n157 VSUBS 0.008191f
C456 B.n158 VSUBS 0.008191f
C457 B.n159 VSUBS 0.008191f
C458 B.n160 VSUBS 0.008191f
C459 B.n161 VSUBS 0.008191f
C460 B.t10 VSUBS 0.340088f
C461 B.t11 VSUBS 0.370404f
C462 B.t9 VSUBS 1.53091f
C463 B.n162 VSUBS 0.554705f
C464 B.n163 VSUBS 0.345039f
C465 B.n164 VSUBS 0.008191f
C466 B.n165 VSUBS 0.008191f
C467 B.n166 VSUBS 0.008191f
C468 B.n167 VSUBS 0.008191f
C469 B.t1 VSUBS 0.340084f
C470 B.t2 VSUBS 0.3704f
C471 B.t0 VSUBS 1.53091f
C472 B.n168 VSUBS 0.554709f
C473 B.n169 VSUBS 0.345042f
C474 B.n170 VSUBS 0.018977f
C475 B.n171 VSUBS 0.008191f
C476 B.n172 VSUBS 0.008191f
C477 B.n173 VSUBS 0.008191f
C478 B.n174 VSUBS 0.008191f
C479 B.n175 VSUBS 0.008191f
C480 B.n176 VSUBS 0.008191f
C481 B.n177 VSUBS 0.008191f
C482 B.n178 VSUBS 0.008191f
C483 B.n179 VSUBS 0.008191f
C484 B.n180 VSUBS 0.008191f
C485 B.n181 VSUBS 0.008191f
C486 B.n182 VSUBS 0.008191f
C487 B.n183 VSUBS 0.008191f
C488 B.n184 VSUBS 0.008191f
C489 B.n185 VSUBS 0.008191f
C490 B.n186 VSUBS 0.008191f
C491 B.n187 VSUBS 0.008191f
C492 B.n188 VSUBS 0.008191f
C493 B.n189 VSUBS 0.008191f
C494 B.n190 VSUBS 0.008191f
C495 B.n191 VSUBS 0.008191f
C496 B.n192 VSUBS 0.008191f
C497 B.n193 VSUBS 0.008191f
C498 B.n194 VSUBS 0.008191f
C499 B.n195 VSUBS 0.008191f
C500 B.n196 VSUBS 0.019869f
C501 B.n197 VSUBS 0.008191f
C502 B.n198 VSUBS 0.008191f
C503 B.n199 VSUBS 0.008191f
C504 B.n200 VSUBS 0.008191f
C505 B.n201 VSUBS 0.008191f
C506 B.n202 VSUBS 0.008191f
C507 B.n203 VSUBS 0.008191f
C508 B.n204 VSUBS 0.008191f
C509 B.n205 VSUBS 0.008191f
C510 B.n206 VSUBS 0.008191f
C511 B.n207 VSUBS 0.008191f
C512 B.n208 VSUBS 0.008191f
C513 B.n209 VSUBS 0.008191f
C514 B.n210 VSUBS 0.008191f
C515 B.n211 VSUBS 0.008191f
C516 B.n212 VSUBS 0.008191f
C517 B.n213 VSUBS 0.008191f
C518 B.n214 VSUBS 0.008191f
C519 B.n215 VSUBS 0.008191f
C520 B.n216 VSUBS 0.008191f
C521 B.n217 VSUBS 0.008191f
C522 B.n218 VSUBS 0.008191f
C523 B.n219 VSUBS 0.008191f
C524 B.n220 VSUBS 0.008191f
C525 B.n221 VSUBS 0.008191f
C526 B.n222 VSUBS 0.008191f
C527 B.n223 VSUBS 0.008191f
C528 B.n224 VSUBS 0.008191f
C529 B.n225 VSUBS 0.008191f
C530 B.n226 VSUBS 0.008191f
C531 B.n227 VSUBS 0.008191f
C532 B.n228 VSUBS 0.008191f
C533 B.n229 VSUBS 0.008191f
C534 B.n230 VSUBS 0.008191f
C535 B.n231 VSUBS 0.008191f
C536 B.n232 VSUBS 0.008191f
C537 B.n233 VSUBS 0.008191f
C538 B.n234 VSUBS 0.008191f
C539 B.n235 VSUBS 0.008191f
C540 B.n236 VSUBS 0.008191f
C541 B.n237 VSUBS 0.008191f
C542 B.n238 VSUBS 0.008191f
C543 B.n239 VSUBS 0.008191f
C544 B.n240 VSUBS 0.008191f
C545 B.n241 VSUBS 0.008191f
C546 B.n242 VSUBS 0.008191f
C547 B.n243 VSUBS 0.008191f
C548 B.n244 VSUBS 0.008191f
C549 B.n245 VSUBS 0.008191f
C550 B.n246 VSUBS 0.008191f
C551 B.n247 VSUBS 0.008191f
C552 B.n248 VSUBS 0.008191f
C553 B.n249 VSUBS 0.008191f
C554 B.n250 VSUBS 0.008191f
C555 B.n251 VSUBS 0.008191f
C556 B.n252 VSUBS 0.008191f
C557 B.n253 VSUBS 0.008191f
C558 B.n254 VSUBS 0.008191f
C559 B.n255 VSUBS 0.008191f
C560 B.n256 VSUBS 0.008191f
C561 B.n257 VSUBS 0.008191f
C562 B.n258 VSUBS 0.008191f
C563 B.n259 VSUBS 0.008191f
C564 B.n260 VSUBS 0.008191f
C565 B.n261 VSUBS 0.008191f
C566 B.n262 VSUBS 0.008191f
C567 B.n263 VSUBS 0.008191f
C568 B.n264 VSUBS 0.008191f
C569 B.n265 VSUBS 0.008191f
C570 B.n266 VSUBS 0.008191f
C571 B.n267 VSUBS 0.008191f
C572 B.n268 VSUBS 0.008191f
C573 B.n269 VSUBS 0.008191f
C574 B.n270 VSUBS 0.008191f
C575 B.n271 VSUBS 0.008191f
C576 B.n272 VSUBS 0.008191f
C577 B.n273 VSUBS 0.008191f
C578 B.n274 VSUBS 0.008191f
C579 B.n275 VSUBS 0.008191f
C580 B.n276 VSUBS 0.008191f
C581 B.n277 VSUBS 0.008191f
C582 B.n278 VSUBS 0.008191f
C583 B.n279 VSUBS 0.008191f
C584 B.n280 VSUBS 0.008191f
C585 B.n281 VSUBS 0.008191f
C586 B.n282 VSUBS 0.008191f
C587 B.n283 VSUBS 0.008191f
C588 B.n284 VSUBS 0.008191f
C589 B.n285 VSUBS 0.008191f
C590 B.n286 VSUBS 0.008191f
C591 B.n287 VSUBS 0.008191f
C592 B.n288 VSUBS 0.008191f
C593 B.n289 VSUBS 0.019157f
C594 B.n290 VSUBS 0.019157f
C595 B.n291 VSUBS 0.019869f
C596 B.n292 VSUBS 0.008191f
C597 B.n293 VSUBS 0.008191f
C598 B.n294 VSUBS 0.008191f
C599 B.n295 VSUBS 0.008191f
C600 B.n296 VSUBS 0.008191f
C601 B.n297 VSUBS 0.008191f
C602 B.n298 VSUBS 0.008191f
C603 B.n299 VSUBS 0.008191f
C604 B.n300 VSUBS 0.008191f
C605 B.n301 VSUBS 0.008191f
C606 B.n302 VSUBS 0.008191f
C607 B.n303 VSUBS 0.008191f
C608 B.n304 VSUBS 0.008191f
C609 B.n305 VSUBS 0.008191f
C610 B.n306 VSUBS 0.008191f
C611 B.n307 VSUBS 0.008191f
C612 B.n308 VSUBS 0.008191f
C613 B.n309 VSUBS 0.008191f
C614 B.n310 VSUBS 0.008191f
C615 B.n311 VSUBS 0.008191f
C616 B.n312 VSUBS 0.008191f
C617 B.n313 VSUBS 0.008191f
C618 B.n314 VSUBS 0.008191f
C619 B.n315 VSUBS 0.008191f
C620 B.n316 VSUBS 0.008191f
C621 B.n317 VSUBS 0.008191f
C622 B.n318 VSUBS 0.008191f
C623 B.n319 VSUBS 0.008191f
C624 B.n320 VSUBS 0.008191f
C625 B.n321 VSUBS 0.008191f
C626 B.n322 VSUBS 0.008191f
C627 B.n323 VSUBS 0.008191f
C628 B.n324 VSUBS 0.008191f
C629 B.n325 VSUBS 0.008191f
C630 B.n326 VSUBS 0.008191f
C631 B.n327 VSUBS 0.008191f
C632 B.n328 VSUBS 0.008191f
C633 B.n329 VSUBS 0.008191f
C634 B.n330 VSUBS 0.008191f
C635 B.n331 VSUBS 0.008191f
C636 B.n332 VSUBS 0.008191f
C637 B.n333 VSUBS 0.008191f
C638 B.n334 VSUBS 0.008191f
C639 B.n335 VSUBS 0.008191f
C640 B.n336 VSUBS 0.008191f
C641 B.n337 VSUBS 0.008191f
C642 B.n338 VSUBS 0.008191f
C643 B.n339 VSUBS 0.008191f
C644 B.n340 VSUBS 0.008191f
C645 B.n341 VSUBS 0.008191f
C646 B.n342 VSUBS 0.008191f
C647 B.n343 VSUBS 0.008191f
C648 B.n344 VSUBS 0.008191f
C649 B.n345 VSUBS 0.008191f
C650 B.n346 VSUBS 0.008191f
C651 B.n347 VSUBS 0.008191f
C652 B.n348 VSUBS 0.008191f
C653 B.n349 VSUBS 0.008191f
C654 B.n350 VSUBS 0.008191f
C655 B.n351 VSUBS 0.008191f
C656 B.n352 VSUBS 0.008191f
C657 B.n353 VSUBS 0.008191f
C658 B.n354 VSUBS 0.008191f
C659 B.n355 VSUBS 0.008191f
C660 B.n356 VSUBS 0.008191f
C661 B.n357 VSUBS 0.008191f
C662 B.n358 VSUBS 0.008191f
C663 B.n359 VSUBS 0.008191f
C664 B.n360 VSUBS 0.008191f
C665 B.n361 VSUBS 0.008191f
C666 B.n362 VSUBS 0.008191f
C667 B.n363 VSUBS 0.008191f
C668 B.n364 VSUBS 0.008191f
C669 B.n365 VSUBS 0.008191f
C670 B.n366 VSUBS 0.008191f
C671 B.n367 VSUBS 0.005661f
C672 B.n368 VSUBS 0.008191f
C673 B.n369 VSUBS 0.008191f
C674 B.n370 VSUBS 0.006625f
C675 B.n371 VSUBS 0.008191f
C676 B.n372 VSUBS 0.008191f
C677 B.n373 VSUBS 0.008191f
C678 B.n374 VSUBS 0.008191f
C679 B.n375 VSUBS 0.008191f
C680 B.n376 VSUBS 0.008191f
C681 B.n377 VSUBS 0.008191f
C682 B.n378 VSUBS 0.008191f
C683 B.n379 VSUBS 0.008191f
C684 B.n380 VSUBS 0.008191f
C685 B.n381 VSUBS 0.008191f
C686 B.n382 VSUBS 0.006625f
C687 B.n383 VSUBS 0.018977f
C688 B.n384 VSUBS 0.005661f
C689 B.n385 VSUBS 0.008191f
C690 B.n386 VSUBS 0.008191f
C691 B.n387 VSUBS 0.008191f
C692 B.n388 VSUBS 0.008191f
C693 B.n389 VSUBS 0.008191f
C694 B.n390 VSUBS 0.008191f
C695 B.n391 VSUBS 0.008191f
C696 B.n392 VSUBS 0.008191f
C697 B.n393 VSUBS 0.008191f
C698 B.n394 VSUBS 0.008191f
C699 B.n395 VSUBS 0.008191f
C700 B.n396 VSUBS 0.008191f
C701 B.n397 VSUBS 0.008191f
C702 B.n398 VSUBS 0.008191f
C703 B.n399 VSUBS 0.008191f
C704 B.n400 VSUBS 0.008191f
C705 B.n401 VSUBS 0.008191f
C706 B.n402 VSUBS 0.008191f
C707 B.n403 VSUBS 0.008191f
C708 B.n404 VSUBS 0.008191f
C709 B.n405 VSUBS 0.008191f
C710 B.n406 VSUBS 0.008191f
C711 B.n407 VSUBS 0.008191f
C712 B.n408 VSUBS 0.008191f
C713 B.n409 VSUBS 0.008191f
C714 B.n410 VSUBS 0.008191f
C715 B.n411 VSUBS 0.008191f
C716 B.n412 VSUBS 0.008191f
C717 B.n413 VSUBS 0.008191f
C718 B.n414 VSUBS 0.008191f
C719 B.n415 VSUBS 0.008191f
C720 B.n416 VSUBS 0.008191f
C721 B.n417 VSUBS 0.008191f
C722 B.n418 VSUBS 0.008191f
C723 B.n419 VSUBS 0.008191f
C724 B.n420 VSUBS 0.008191f
C725 B.n421 VSUBS 0.008191f
C726 B.n422 VSUBS 0.008191f
C727 B.n423 VSUBS 0.008191f
C728 B.n424 VSUBS 0.008191f
C729 B.n425 VSUBS 0.008191f
C730 B.n426 VSUBS 0.008191f
C731 B.n427 VSUBS 0.008191f
C732 B.n428 VSUBS 0.008191f
C733 B.n429 VSUBS 0.008191f
C734 B.n430 VSUBS 0.008191f
C735 B.n431 VSUBS 0.008191f
C736 B.n432 VSUBS 0.008191f
C737 B.n433 VSUBS 0.008191f
C738 B.n434 VSUBS 0.008191f
C739 B.n435 VSUBS 0.008191f
C740 B.n436 VSUBS 0.008191f
C741 B.n437 VSUBS 0.008191f
C742 B.n438 VSUBS 0.008191f
C743 B.n439 VSUBS 0.008191f
C744 B.n440 VSUBS 0.008191f
C745 B.n441 VSUBS 0.008191f
C746 B.n442 VSUBS 0.008191f
C747 B.n443 VSUBS 0.008191f
C748 B.n444 VSUBS 0.008191f
C749 B.n445 VSUBS 0.008191f
C750 B.n446 VSUBS 0.008191f
C751 B.n447 VSUBS 0.008191f
C752 B.n448 VSUBS 0.008191f
C753 B.n449 VSUBS 0.008191f
C754 B.n450 VSUBS 0.008191f
C755 B.n451 VSUBS 0.008191f
C756 B.n452 VSUBS 0.008191f
C757 B.n453 VSUBS 0.008191f
C758 B.n454 VSUBS 0.008191f
C759 B.n455 VSUBS 0.008191f
C760 B.n456 VSUBS 0.008191f
C761 B.n457 VSUBS 0.008191f
C762 B.n458 VSUBS 0.008191f
C763 B.n459 VSUBS 0.008191f
C764 B.n460 VSUBS 0.019869f
C765 B.n461 VSUBS 0.019869f
C766 B.n462 VSUBS 0.019157f
C767 B.n463 VSUBS 0.008191f
C768 B.n464 VSUBS 0.008191f
C769 B.n465 VSUBS 0.008191f
C770 B.n466 VSUBS 0.008191f
C771 B.n467 VSUBS 0.008191f
C772 B.n468 VSUBS 0.008191f
C773 B.n469 VSUBS 0.008191f
C774 B.n470 VSUBS 0.008191f
C775 B.n471 VSUBS 0.008191f
C776 B.n472 VSUBS 0.008191f
C777 B.n473 VSUBS 0.008191f
C778 B.n474 VSUBS 0.008191f
C779 B.n475 VSUBS 0.008191f
C780 B.n476 VSUBS 0.008191f
C781 B.n477 VSUBS 0.008191f
C782 B.n478 VSUBS 0.008191f
C783 B.n479 VSUBS 0.008191f
C784 B.n480 VSUBS 0.008191f
C785 B.n481 VSUBS 0.008191f
C786 B.n482 VSUBS 0.008191f
C787 B.n483 VSUBS 0.008191f
C788 B.n484 VSUBS 0.008191f
C789 B.n485 VSUBS 0.008191f
C790 B.n486 VSUBS 0.008191f
C791 B.n487 VSUBS 0.008191f
C792 B.n488 VSUBS 0.008191f
C793 B.n489 VSUBS 0.008191f
C794 B.n490 VSUBS 0.008191f
C795 B.n491 VSUBS 0.008191f
C796 B.n492 VSUBS 0.008191f
C797 B.n493 VSUBS 0.008191f
C798 B.n494 VSUBS 0.008191f
C799 B.n495 VSUBS 0.008191f
C800 B.n496 VSUBS 0.008191f
C801 B.n497 VSUBS 0.008191f
C802 B.n498 VSUBS 0.008191f
C803 B.n499 VSUBS 0.008191f
C804 B.n500 VSUBS 0.008191f
C805 B.n501 VSUBS 0.008191f
C806 B.n502 VSUBS 0.008191f
C807 B.n503 VSUBS 0.008191f
C808 B.n504 VSUBS 0.008191f
C809 B.n505 VSUBS 0.008191f
C810 B.n506 VSUBS 0.008191f
C811 B.n507 VSUBS 0.008191f
C812 B.n508 VSUBS 0.008191f
C813 B.n509 VSUBS 0.008191f
C814 B.n510 VSUBS 0.008191f
C815 B.n511 VSUBS 0.008191f
C816 B.n512 VSUBS 0.008191f
C817 B.n513 VSUBS 0.008191f
C818 B.n514 VSUBS 0.008191f
C819 B.n515 VSUBS 0.008191f
C820 B.n516 VSUBS 0.008191f
C821 B.n517 VSUBS 0.008191f
C822 B.n518 VSUBS 0.008191f
C823 B.n519 VSUBS 0.008191f
C824 B.n520 VSUBS 0.008191f
C825 B.n521 VSUBS 0.008191f
C826 B.n522 VSUBS 0.008191f
C827 B.n523 VSUBS 0.008191f
C828 B.n524 VSUBS 0.008191f
C829 B.n525 VSUBS 0.008191f
C830 B.n526 VSUBS 0.008191f
C831 B.n527 VSUBS 0.008191f
C832 B.n528 VSUBS 0.008191f
C833 B.n529 VSUBS 0.008191f
C834 B.n530 VSUBS 0.008191f
C835 B.n531 VSUBS 0.008191f
C836 B.n532 VSUBS 0.008191f
C837 B.n533 VSUBS 0.008191f
C838 B.n534 VSUBS 0.008191f
C839 B.n535 VSUBS 0.008191f
C840 B.n536 VSUBS 0.008191f
C841 B.n537 VSUBS 0.008191f
C842 B.n538 VSUBS 0.008191f
C843 B.n539 VSUBS 0.008191f
C844 B.n540 VSUBS 0.008191f
C845 B.n541 VSUBS 0.008191f
C846 B.n542 VSUBS 0.008191f
C847 B.n543 VSUBS 0.008191f
C848 B.n544 VSUBS 0.008191f
C849 B.n545 VSUBS 0.008191f
C850 B.n546 VSUBS 0.008191f
C851 B.n547 VSUBS 0.008191f
C852 B.n548 VSUBS 0.008191f
C853 B.n549 VSUBS 0.008191f
C854 B.n550 VSUBS 0.008191f
C855 B.n551 VSUBS 0.008191f
C856 B.n552 VSUBS 0.008191f
C857 B.n553 VSUBS 0.008191f
C858 B.n554 VSUBS 0.008191f
C859 B.n555 VSUBS 0.008191f
C860 B.n556 VSUBS 0.008191f
C861 B.n557 VSUBS 0.008191f
C862 B.n558 VSUBS 0.008191f
C863 B.n559 VSUBS 0.008191f
C864 B.n560 VSUBS 0.008191f
C865 B.n561 VSUBS 0.008191f
C866 B.n562 VSUBS 0.008191f
C867 B.n563 VSUBS 0.008191f
C868 B.n564 VSUBS 0.008191f
C869 B.n565 VSUBS 0.008191f
C870 B.n566 VSUBS 0.008191f
C871 B.n567 VSUBS 0.008191f
C872 B.n568 VSUBS 0.008191f
C873 B.n569 VSUBS 0.008191f
C874 B.n570 VSUBS 0.008191f
C875 B.n571 VSUBS 0.008191f
C876 B.n572 VSUBS 0.008191f
C877 B.n573 VSUBS 0.008191f
C878 B.n574 VSUBS 0.008191f
C879 B.n575 VSUBS 0.008191f
C880 B.n576 VSUBS 0.008191f
C881 B.n577 VSUBS 0.008191f
C882 B.n578 VSUBS 0.008191f
C883 B.n579 VSUBS 0.008191f
C884 B.n580 VSUBS 0.008191f
C885 B.n581 VSUBS 0.008191f
C886 B.n582 VSUBS 0.008191f
C887 B.n583 VSUBS 0.008191f
C888 B.n584 VSUBS 0.008191f
C889 B.n585 VSUBS 0.008191f
C890 B.n586 VSUBS 0.008191f
C891 B.n587 VSUBS 0.008191f
C892 B.n588 VSUBS 0.008191f
C893 B.n589 VSUBS 0.008191f
C894 B.n590 VSUBS 0.008191f
C895 B.n591 VSUBS 0.008191f
C896 B.n592 VSUBS 0.008191f
C897 B.n593 VSUBS 0.008191f
C898 B.n594 VSUBS 0.008191f
C899 B.n595 VSUBS 0.008191f
C900 B.n596 VSUBS 0.008191f
C901 B.n597 VSUBS 0.008191f
C902 B.n598 VSUBS 0.008191f
C903 B.n599 VSUBS 0.008191f
C904 B.n600 VSUBS 0.008191f
C905 B.n601 VSUBS 0.008191f
C906 B.n602 VSUBS 0.008191f
C907 B.n603 VSUBS 0.008191f
C908 B.n604 VSUBS 0.008191f
C909 B.n605 VSUBS 0.008191f
C910 B.n606 VSUBS 0.020098f
C911 B.n607 VSUBS 0.018927f
C912 B.n608 VSUBS 0.019869f
C913 B.n609 VSUBS 0.008191f
C914 B.n610 VSUBS 0.008191f
C915 B.n611 VSUBS 0.008191f
C916 B.n612 VSUBS 0.008191f
C917 B.n613 VSUBS 0.008191f
C918 B.n614 VSUBS 0.008191f
C919 B.n615 VSUBS 0.008191f
C920 B.n616 VSUBS 0.008191f
C921 B.n617 VSUBS 0.008191f
C922 B.n618 VSUBS 0.008191f
C923 B.n619 VSUBS 0.008191f
C924 B.n620 VSUBS 0.008191f
C925 B.n621 VSUBS 0.008191f
C926 B.n622 VSUBS 0.008191f
C927 B.n623 VSUBS 0.008191f
C928 B.n624 VSUBS 0.008191f
C929 B.n625 VSUBS 0.008191f
C930 B.n626 VSUBS 0.008191f
C931 B.n627 VSUBS 0.008191f
C932 B.n628 VSUBS 0.008191f
C933 B.n629 VSUBS 0.008191f
C934 B.n630 VSUBS 0.008191f
C935 B.n631 VSUBS 0.008191f
C936 B.n632 VSUBS 0.008191f
C937 B.n633 VSUBS 0.008191f
C938 B.n634 VSUBS 0.008191f
C939 B.n635 VSUBS 0.008191f
C940 B.n636 VSUBS 0.008191f
C941 B.n637 VSUBS 0.008191f
C942 B.n638 VSUBS 0.008191f
C943 B.n639 VSUBS 0.008191f
C944 B.n640 VSUBS 0.008191f
C945 B.n641 VSUBS 0.008191f
C946 B.n642 VSUBS 0.008191f
C947 B.n643 VSUBS 0.008191f
C948 B.n644 VSUBS 0.008191f
C949 B.n645 VSUBS 0.008191f
C950 B.n646 VSUBS 0.008191f
C951 B.n647 VSUBS 0.008191f
C952 B.n648 VSUBS 0.008191f
C953 B.n649 VSUBS 0.008191f
C954 B.n650 VSUBS 0.008191f
C955 B.n651 VSUBS 0.008191f
C956 B.n652 VSUBS 0.008191f
C957 B.n653 VSUBS 0.008191f
C958 B.n654 VSUBS 0.008191f
C959 B.n655 VSUBS 0.008191f
C960 B.n656 VSUBS 0.008191f
C961 B.n657 VSUBS 0.008191f
C962 B.n658 VSUBS 0.008191f
C963 B.n659 VSUBS 0.008191f
C964 B.n660 VSUBS 0.008191f
C965 B.n661 VSUBS 0.008191f
C966 B.n662 VSUBS 0.008191f
C967 B.n663 VSUBS 0.008191f
C968 B.n664 VSUBS 0.008191f
C969 B.n665 VSUBS 0.008191f
C970 B.n666 VSUBS 0.008191f
C971 B.n667 VSUBS 0.008191f
C972 B.n668 VSUBS 0.008191f
C973 B.n669 VSUBS 0.008191f
C974 B.n670 VSUBS 0.008191f
C975 B.n671 VSUBS 0.008191f
C976 B.n672 VSUBS 0.008191f
C977 B.n673 VSUBS 0.008191f
C978 B.n674 VSUBS 0.008191f
C979 B.n675 VSUBS 0.008191f
C980 B.n676 VSUBS 0.008191f
C981 B.n677 VSUBS 0.008191f
C982 B.n678 VSUBS 0.008191f
C983 B.n679 VSUBS 0.008191f
C984 B.n680 VSUBS 0.008191f
C985 B.n681 VSUBS 0.008191f
C986 B.n682 VSUBS 0.008191f
C987 B.n683 VSUBS 0.008191f
C988 B.n684 VSUBS 0.005661f
C989 B.n685 VSUBS 0.018977f
C990 B.n686 VSUBS 0.006625f
C991 B.n687 VSUBS 0.008191f
C992 B.n688 VSUBS 0.008191f
C993 B.n689 VSUBS 0.008191f
C994 B.n690 VSUBS 0.008191f
C995 B.n691 VSUBS 0.008191f
C996 B.n692 VSUBS 0.008191f
C997 B.n693 VSUBS 0.008191f
C998 B.n694 VSUBS 0.008191f
C999 B.n695 VSUBS 0.008191f
C1000 B.n696 VSUBS 0.008191f
C1001 B.n697 VSUBS 0.008191f
C1002 B.n698 VSUBS 0.006625f
C1003 B.n699 VSUBS 0.008191f
C1004 B.n700 VSUBS 0.008191f
C1005 B.n701 VSUBS 0.005661f
C1006 B.n702 VSUBS 0.008191f
C1007 B.n703 VSUBS 0.008191f
C1008 B.n704 VSUBS 0.008191f
C1009 B.n705 VSUBS 0.008191f
C1010 B.n706 VSUBS 0.008191f
C1011 B.n707 VSUBS 0.008191f
C1012 B.n708 VSUBS 0.008191f
C1013 B.n709 VSUBS 0.008191f
C1014 B.n710 VSUBS 0.008191f
C1015 B.n711 VSUBS 0.008191f
C1016 B.n712 VSUBS 0.008191f
C1017 B.n713 VSUBS 0.008191f
C1018 B.n714 VSUBS 0.008191f
C1019 B.n715 VSUBS 0.008191f
C1020 B.n716 VSUBS 0.008191f
C1021 B.n717 VSUBS 0.008191f
C1022 B.n718 VSUBS 0.008191f
C1023 B.n719 VSUBS 0.008191f
C1024 B.n720 VSUBS 0.008191f
C1025 B.n721 VSUBS 0.008191f
C1026 B.n722 VSUBS 0.008191f
C1027 B.n723 VSUBS 0.008191f
C1028 B.n724 VSUBS 0.008191f
C1029 B.n725 VSUBS 0.008191f
C1030 B.n726 VSUBS 0.008191f
C1031 B.n727 VSUBS 0.008191f
C1032 B.n728 VSUBS 0.008191f
C1033 B.n729 VSUBS 0.008191f
C1034 B.n730 VSUBS 0.008191f
C1035 B.n731 VSUBS 0.008191f
C1036 B.n732 VSUBS 0.008191f
C1037 B.n733 VSUBS 0.008191f
C1038 B.n734 VSUBS 0.008191f
C1039 B.n735 VSUBS 0.008191f
C1040 B.n736 VSUBS 0.008191f
C1041 B.n737 VSUBS 0.008191f
C1042 B.n738 VSUBS 0.008191f
C1043 B.n739 VSUBS 0.008191f
C1044 B.n740 VSUBS 0.008191f
C1045 B.n741 VSUBS 0.008191f
C1046 B.n742 VSUBS 0.008191f
C1047 B.n743 VSUBS 0.008191f
C1048 B.n744 VSUBS 0.008191f
C1049 B.n745 VSUBS 0.008191f
C1050 B.n746 VSUBS 0.008191f
C1051 B.n747 VSUBS 0.008191f
C1052 B.n748 VSUBS 0.008191f
C1053 B.n749 VSUBS 0.008191f
C1054 B.n750 VSUBS 0.008191f
C1055 B.n751 VSUBS 0.008191f
C1056 B.n752 VSUBS 0.008191f
C1057 B.n753 VSUBS 0.008191f
C1058 B.n754 VSUBS 0.008191f
C1059 B.n755 VSUBS 0.008191f
C1060 B.n756 VSUBS 0.008191f
C1061 B.n757 VSUBS 0.008191f
C1062 B.n758 VSUBS 0.008191f
C1063 B.n759 VSUBS 0.008191f
C1064 B.n760 VSUBS 0.008191f
C1065 B.n761 VSUBS 0.008191f
C1066 B.n762 VSUBS 0.008191f
C1067 B.n763 VSUBS 0.008191f
C1068 B.n764 VSUBS 0.008191f
C1069 B.n765 VSUBS 0.008191f
C1070 B.n766 VSUBS 0.008191f
C1071 B.n767 VSUBS 0.008191f
C1072 B.n768 VSUBS 0.008191f
C1073 B.n769 VSUBS 0.008191f
C1074 B.n770 VSUBS 0.008191f
C1075 B.n771 VSUBS 0.008191f
C1076 B.n772 VSUBS 0.008191f
C1077 B.n773 VSUBS 0.008191f
C1078 B.n774 VSUBS 0.008191f
C1079 B.n775 VSUBS 0.008191f
C1080 B.n776 VSUBS 0.008191f
C1081 B.n777 VSUBS 0.019869f
C1082 B.n778 VSUBS 0.019157f
C1083 B.n779 VSUBS 0.019157f
C1084 B.n780 VSUBS 0.008191f
C1085 B.n781 VSUBS 0.008191f
C1086 B.n782 VSUBS 0.008191f
C1087 B.n783 VSUBS 0.008191f
C1088 B.n784 VSUBS 0.008191f
C1089 B.n785 VSUBS 0.008191f
C1090 B.n786 VSUBS 0.008191f
C1091 B.n787 VSUBS 0.008191f
C1092 B.n788 VSUBS 0.008191f
C1093 B.n789 VSUBS 0.008191f
C1094 B.n790 VSUBS 0.008191f
C1095 B.n791 VSUBS 0.008191f
C1096 B.n792 VSUBS 0.008191f
C1097 B.n793 VSUBS 0.008191f
C1098 B.n794 VSUBS 0.008191f
C1099 B.n795 VSUBS 0.008191f
C1100 B.n796 VSUBS 0.008191f
C1101 B.n797 VSUBS 0.008191f
C1102 B.n798 VSUBS 0.008191f
C1103 B.n799 VSUBS 0.008191f
C1104 B.n800 VSUBS 0.008191f
C1105 B.n801 VSUBS 0.008191f
C1106 B.n802 VSUBS 0.008191f
C1107 B.n803 VSUBS 0.008191f
C1108 B.n804 VSUBS 0.008191f
C1109 B.n805 VSUBS 0.008191f
C1110 B.n806 VSUBS 0.008191f
C1111 B.n807 VSUBS 0.008191f
C1112 B.n808 VSUBS 0.008191f
C1113 B.n809 VSUBS 0.008191f
C1114 B.n810 VSUBS 0.008191f
C1115 B.n811 VSUBS 0.008191f
C1116 B.n812 VSUBS 0.008191f
C1117 B.n813 VSUBS 0.008191f
C1118 B.n814 VSUBS 0.008191f
C1119 B.n815 VSUBS 0.008191f
C1120 B.n816 VSUBS 0.008191f
C1121 B.n817 VSUBS 0.008191f
C1122 B.n818 VSUBS 0.008191f
C1123 B.n819 VSUBS 0.008191f
C1124 B.n820 VSUBS 0.008191f
C1125 B.n821 VSUBS 0.008191f
C1126 B.n822 VSUBS 0.008191f
C1127 B.n823 VSUBS 0.008191f
C1128 B.n824 VSUBS 0.008191f
C1129 B.n825 VSUBS 0.008191f
C1130 B.n826 VSUBS 0.008191f
C1131 B.n827 VSUBS 0.008191f
C1132 B.n828 VSUBS 0.008191f
C1133 B.n829 VSUBS 0.008191f
C1134 B.n830 VSUBS 0.008191f
C1135 B.n831 VSUBS 0.008191f
C1136 B.n832 VSUBS 0.008191f
C1137 B.n833 VSUBS 0.008191f
C1138 B.n834 VSUBS 0.008191f
C1139 B.n835 VSUBS 0.008191f
C1140 B.n836 VSUBS 0.008191f
C1141 B.n837 VSUBS 0.008191f
C1142 B.n838 VSUBS 0.008191f
C1143 B.n839 VSUBS 0.008191f
C1144 B.n840 VSUBS 0.008191f
C1145 B.n841 VSUBS 0.008191f
C1146 B.n842 VSUBS 0.008191f
C1147 B.n843 VSUBS 0.008191f
C1148 B.n844 VSUBS 0.008191f
C1149 B.n845 VSUBS 0.008191f
C1150 B.n846 VSUBS 0.008191f
C1151 B.n847 VSUBS 0.008191f
C1152 B.n848 VSUBS 0.008191f
C1153 B.n849 VSUBS 0.008191f
C1154 B.n850 VSUBS 0.008191f
C1155 B.n851 VSUBS 0.018546f
C1156 VDD1.n0 VSUBS 0.028848f
C1157 VDD1.n1 VSUBS 0.026875f
C1158 VDD1.n2 VSUBS 0.014441f
C1159 VDD1.n3 VSUBS 0.034134f
C1160 VDD1.n4 VSUBS 0.014866f
C1161 VDD1.n5 VSUBS 0.026875f
C1162 VDD1.n6 VSUBS 0.014866f
C1163 VDD1.n7 VSUBS 0.014441f
C1164 VDD1.n8 VSUBS 0.034134f
C1165 VDD1.n9 VSUBS 0.034134f
C1166 VDD1.n10 VSUBS 0.015291f
C1167 VDD1.n11 VSUBS 0.026875f
C1168 VDD1.n12 VSUBS 0.014441f
C1169 VDD1.n13 VSUBS 0.034134f
C1170 VDD1.n14 VSUBS 0.015291f
C1171 VDD1.n15 VSUBS 0.026875f
C1172 VDD1.n16 VSUBS 0.014441f
C1173 VDD1.n17 VSUBS 0.034134f
C1174 VDD1.n18 VSUBS 0.015291f
C1175 VDD1.n19 VSUBS 0.026875f
C1176 VDD1.n20 VSUBS 0.014441f
C1177 VDD1.n21 VSUBS 0.034134f
C1178 VDD1.n22 VSUBS 0.015291f
C1179 VDD1.n23 VSUBS 0.026875f
C1180 VDD1.n24 VSUBS 0.014441f
C1181 VDD1.n25 VSUBS 0.034134f
C1182 VDD1.n26 VSUBS 0.015291f
C1183 VDD1.n27 VSUBS 1.77336f
C1184 VDD1.n28 VSUBS 0.014441f
C1185 VDD1.t0 VSUBS 0.073106f
C1186 VDD1.n29 VSUBS 0.19317f
C1187 VDD1.n30 VSUBS 0.021715f
C1188 VDD1.n31 VSUBS 0.025601f
C1189 VDD1.n32 VSUBS 0.034134f
C1190 VDD1.n33 VSUBS 0.015291f
C1191 VDD1.n34 VSUBS 0.014441f
C1192 VDD1.n35 VSUBS 0.026875f
C1193 VDD1.n36 VSUBS 0.026875f
C1194 VDD1.n37 VSUBS 0.014441f
C1195 VDD1.n38 VSUBS 0.015291f
C1196 VDD1.n39 VSUBS 0.034134f
C1197 VDD1.n40 VSUBS 0.034134f
C1198 VDD1.n41 VSUBS 0.015291f
C1199 VDD1.n42 VSUBS 0.014441f
C1200 VDD1.n43 VSUBS 0.026875f
C1201 VDD1.n44 VSUBS 0.026875f
C1202 VDD1.n45 VSUBS 0.014441f
C1203 VDD1.n46 VSUBS 0.015291f
C1204 VDD1.n47 VSUBS 0.034134f
C1205 VDD1.n48 VSUBS 0.034134f
C1206 VDD1.n49 VSUBS 0.015291f
C1207 VDD1.n50 VSUBS 0.014441f
C1208 VDD1.n51 VSUBS 0.026875f
C1209 VDD1.n52 VSUBS 0.026875f
C1210 VDD1.n53 VSUBS 0.014441f
C1211 VDD1.n54 VSUBS 0.015291f
C1212 VDD1.n55 VSUBS 0.034134f
C1213 VDD1.n56 VSUBS 0.034134f
C1214 VDD1.n57 VSUBS 0.015291f
C1215 VDD1.n58 VSUBS 0.014441f
C1216 VDD1.n59 VSUBS 0.026875f
C1217 VDD1.n60 VSUBS 0.026875f
C1218 VDD1.n61 VSUBS 0.014441f
C1219 VDD1.n62 VSUBS 0.015291f
C1220 VDD1.n63 VSUBS 0.034134f
C1221 VDD1.n64 VSUBS 0.034134f
C1222 VDD1.n65 VSUBS 0.015291f
C1223 VDD1.n66 VSUBS 0.014441f
C1224 VDD1.n67 VSUBS 0.026875f
C1225 VDD1.n68 VSUBS 0.026875f
C1226 VDD1.n69 VSUBS 0.014441f
C1227 VDD1.n70 VSUBS 0.015291f
C1228 VDD1.n71 VSUBS 0.034134f
C1229 VDD1.n72 VSUBS 0.034134f
C1230 VDD1.n73 VSUBS 0.015291f
C1231 VDD1.n74 VSUBS 0.014441f
C1232 VDD1.n75 VSUBS 0.026875f
C1233 VDD1.n76 VSUBS 0.026875f
C1234 VDD1.n77 VSUBS 0.014441f
C1235 VDD1.n78 VSUBS 0.015291f
C1236 VDD1.n79 VSUBS 0.034134f
C1237 VDD1.n80 VSUBS 0.080312f
C1238 VDD1.n81 VSUBS 0.015291f
C1239 VDD1.n82 VSUBS 0.014441f
C1240 VDD1.n83 VSUBS 0.066159f
C1241 VDD1.n84 VSUBS 0.06713f
C1242 VDD1.t2 VSUBS 0.328542f
C1243 VDD1.t1 VSUBS 0.328542f
C1244 VDD1.n85 VSUBS 2.68558f
C1245 VDD1.n86 VSUBS 0.939435f
C1246 VDD1.n87 VSUBS 0.028848f
C1247 VDD1.n88 VSUBS 0.026875f
C1248 VDD1.n89 VSUBS 0.014441f
C1249 VDD1.n90 VSUBS 0.034134f
C1250 VDD1.n91 VSUBS 0.014866f
C1251 VDD1.n92 VSUBS 0.026875f
C1252 VDD1.n93 VSUBS 0.015291f
C1253 VDD1.n94 VSUBS 0.034134f
C1254 VDD1.n95 VSUBS 0.015291f
C1255 VDD1.n96 VSUBS 0.026875f
C1256 VDD1.n97 VSUBS 0.014441f
C1257 VDD1.n98 VSUBS 0.034134f
C1258 VDD1.n99 VSUBS 0.015291f
C1259 VDD1.n100 VSUBS 0.026875f
C1260 VDD1.n101 VSUBS 0.014441f
C1261 VDD1.n102 VSUBS 0.034134f
C1262 VDD1.n103 VSUBS 0.015291f
C1263 VDD1.n104 VSUBS 0.026875f
C1264 VDD1.n105 VSUBS 0.014441f
C1265 VDD1.n106 VSUBS 0.034134f
C1266 VDD1.n107 VSUBS 0.015291f
C1267 VDD1.n108 VSUBS 0.026875f
C1268 VDD1.n109 VSUBS 0.014441f
C1269 VDD1.n110 VSUBS 0.034134f
C1270 VDD1.n111 VSUBS 0.015291f
C1271 VDD1.n112 VSUBS 1.77336f
C1272 VDD1.n113 VSUBS 0.014441f
C1273 VDD1.t9 VSUBS 0.073106f
C1274 VDD1.n114 VSUBS 0.19317f
C1275 VDD1.n115 VSUBS 0.021715f
C1276 VDD1.n116 VSUBS 0.025601f
C1277 VDD1.n117 VSUBS 0.034134f
C1278 VDD1.n118 VSUBS 0.015291f
C1279 VDD1.n119 VSUBS 0.014441f
C1280 VDD1.n120 VSUBS 0.026875f
C1281 VDD1.n121 VSUBS 0.026875f
C1282 VDD1.n122 VSUBS 0.014441f
C1283 VDD1.n123 VSUBS 0.015291f
C1284 VDD1.n124 VSUBS 0.034134f
C1285 VDD1.n125 VSUBS 0.034134f
C1286 VDD1.n126 VSUBS 0.015291f
C1287 VDD1.n127 VSUBS 0.014441f
C1288 VDD1.n128 VSUBS 0.026875f
C1289 VDD1.n129 VSUBS 0.026875f
C1290 VDD1.n130 VSUBS 0.014441f
C1291 VDD1.n131 VSUBS 0.015291f
C1292 VDD1.n132 VSUBS 0.034134f
C1293 VDD1.n133 VSUBS 0.034134f
C1294 VDD1.n134 VSUBS 0.015291f
C1295 VDD1.n135 VSUBS 0.014441f
C1296 VDD1.n136 VSUBS 0.026875f
C1297 VDD1.n137 VSUBS 0.026875f
C1298 VDD1.n138 VSUBS 0.014441f
C1299 VDD1.n139 VSUBS 0.015291f
C1300 VDD1.n140 VSUBS 0.034134f
C1301 VDD1.n141 VSUBS 0.034134f
C1302 VDD1.n142 VSUBS 0.015291f
C1303 VDD1.n143 VSUBS 0.014441f
C1304 VDD1.n144 VSUBS 0.026875f
C1305 VDD1.n145 VSUBS 0.026875f
C1306 VDD1.n146 VSUBS 0.014441f
C1307 VDD1.n147 VSUBS 0.015291f
C1308 VDD1.n148 VSUBS 0.034134f
C1309 VDD1.n149 VSUBS 0.034134f
C1310 VDD1.n150 VSUBS 0.015291f
C1311 VDD1.n151 VSUBS 0.014441f
C1312 VDD1.n152 VSUBS 0.026875f
C1313 VDD1.n153 VSUBS 0.026875f
C1314 VDD1.n154 VSUBS 0.014441f
C1315 VDD1.n155 VSUBS 0.014441f
C1316 VDD1.n156 VSUBS 0.015291f
C1317 VDD1.n157 VSUBS 0.034134f
C1318 VDD1.n158 VSUBS 0.034134f
C1319 VDD1.n159 VSUBS 0.034134f
C1320 VDD1.n160 VSUBS 0.014866f
C1321 VDD1.n161 VSUBS 0.014441f
C1322 VDD1.n162 VSUBS 0.026875f
C1323 VDD1.n163 VSUBS 0.026875f
C1324 VDD1.n164 VSUBS 0.014441f
C1325 VDD1.n165 VSUBS 0.015291f
C1326 VDD1.n166 VSUBS 0.034134f
C1327 VDD1.n167 VSUBS 0.080312f
C1328 VDD1.n168 VSUBS 0.015291f
C1329 VDD1.n169 VSUBS 0.014441f
C1330 VDD1.n170 VSUBS 0.066159f
C1331 VDD1.n171 VSUBS 0.06713f
C1332 VDD1.t8 VSUBS 0.328542f
C1333 VDD1.t7 VSUBS 0.328542f
C1334 VDD1.n172 VSUBS 2.68557f
C1335 VDD1.n173 VSUBS 0.931059f
C1336 VDD1.t6 VSUBS 0.328542f
C1337 VDD1.t3 VSUBS 0.328542f
C1338 VDD1.n174 VSUBS 2.70102f
C1339 VDD1.n175 VSUBS 3.37865f
C1340 VDD1.t4 VSUBS 0.328542f
C1341 VDD1.t5 VSUBS 0.328542f
C1342 VDD1.n176 VSUBS 2.68557f
C1343 VDD1.n177 VSUBS 3.68508f
C1344 VTAIL.t2 VSUBS 0.335869f
C1345 VTAIL.t8 VSUBS 0.335869f
C1346 VTAIL.n0 VSUBS 2.59127f
C1347 VTAIL.n1 VSUBS 0.899479f
C1348 VTAIL.n2 VSUBS 0.029491f
C1349 VTAIL.n3 VSUBS 0.027474f
C1350 VTAIL.n4 VSUBS 0.014763f
C1351 VTAIL.n5 VSUBS 0.034896f
C1352 VTAIL.n6 VSUBS 0.015198f
C1353 VTAIL.n7 VSUBS 0.027474f
C1354 VTAIL.n8 VSUBS 0.015632f
C1355 VTAIL.n9 VSUBS 0.034896f
C1356 VTAIL.n10 VSUBS 0.015632f
C1357 VTAIL.n11 VSUBS 0.027474f
C1358 VTAIL.n12 VSUBS 0.014763f
C1359 VTAIL.n13 VSUBS 0.034896f
C1360 VTAIL.n14 VSUBS 0.015632f
C1361 VTAIL.n15 VSUBS 0.027474f
C1362 VTAIL.n16 VSUBS 0.014763f
C1363 VTAIL.n17 VSUBS 0.034896f
C1364 VTAIL.n18 VSUBS 0.015632f
C1365 VTAIL.n19 VSUBS 0.027474f
C1366 VTAIL.n20 VSUBS 0.014763f
C1367 VTAIL.n21 VSUBS 0.034896f
C1368 VTAIL.n22 VSUBS 0.015632f
C1369 VTAIL.n23 VSUBS 0.027474f
C1370 VTAIL.n24 VSUBS 0.014763f
C1371 VTAIL.n25 VSUBS 0.034896f
C1372 VTAIL.n26 VSUBS 0.015632f
C1373 VTAIL.n27 VSUBS 1.81291f
C1374 VTAIL.n28 VSUBS 0.014763f
C1375 VTAIL.t19 VSUBS 0.074736f
C1376 VTAIL.n29 VSUBS 0.197478f
C1377 VTAIL.n30 VSUBS 0.022199f
C1378 VTAIL.n31 VSUBS 0.026172f
C1379 VTAIL.n32 VSUBS 0.034896f
C1380 VTAIL.n33 VSUBS 0.015632f
C1381 VTAIL.n34 VSUBS 0.014763f
C1382 VTAIL.n35 VSUBS 0.027474f
C1383 VTAIL.n36 VSUBS 0.027474f
C1384 VTAIL.n37 VSUBS 0.014763f
C1385 VTAIL.n38 VSUBS 0.015632f
C1386 VTAIL.n39 VSUBS 0.034896f
C1387 VTAIL.n40 VSUBS 0.034896f
C1388 VTAIL.n41 VSUBS 0.015632f
C1389 VTAIL.n42 VSUBS 0.014763f
C1390 VTAIL.n43 VSUBS 0.027474f
C1391 VTAIL.n44 VSUBS 0.027474f
C1392 VTAIL.n45 VSUBS 0.014763f
C1393 VTAIL.n46 VSUBS 0.015632f
C1394 VTAIL.n47 VSUBS 0.034896f
C1395 VTAIL.n48 VSUBS 0.034896f
C1396 VTAIL.n49 VSUBS 0.015632f
C1397 VTAIL.n50 VSUBS 0.014763f
C1398 VTAIL.n51 VSUBS 0.027474f
C1399 VTAIL.n52 VSUBS 0.027474f
C1400 VTAIL.n53 VSUBS 0.014763f
C1401 VTAIL.n54 VSUBS 0.015632f
C1402 VTAIL.n55 VSUBS 0.034896f
C1403 VTAIL.n56 VSUBS 0.034896f
C1404 VTAIL.n57 VSUBS 0.015632f
C1405 VTAIL.n58 VSUBS 0.014763f
C1406 VTAIL.n59 VSUBS 0.027474f
C1407 VTAIL.n60 VSUBS 0.027474f
C1408 VTAIL.n61 VSUBS 0.014763f
C1409 VTAIL.n62 VSUBS 0.015632f
C1410 VTAIL.n63 VSUBS 0.034896f
C1411 VTAIL.n64 VSUBS 0.034896f
C1412 VTAIL.n65 VSUBS 0.015632f
C1413 VTAIL.n66 VSUBS 0.014763f
C1414 VTAIL.n67 VSUBS 0.027474f
C1415 VTAIL.n68 VSUBS 0.027474f
C1416 VTAIL.n69 VSUBS 0.014763f
C1417 VTAIL.n70 VSUBS 0.014763f
C1418 VTAIL.n71 VSUBS 0.015632f
C1419 VTAIL.n72 VSUBS 0.034896f
C1420 VTAIL.n73 VSUBS 0.034896f
C1421 VTAIL.n74 VSUBS 0.034896f
C1422 VTAIL.n75 VSUBS 0.015198f
C1423 VTAIL.n76 VSUBS 0.014763f
C1424 VTAIL.n77 VSUBS 0.027474f
C1425 VTAIL.n78 VSUBS 0.027474f
C1426 VTAIL.n79 VSUBS 0.014763f
C1427 VTAIL.n80 VSUBS 0.015632f
C1428 VTAIL.n81 VSUBS 0.034896f
C1429 VTAIL.n82 VSUBS 0.082103f
C1430 VTAIL.n83 VSUBS 0.015632f
C1431 VTAIL.n84 VSUBS 0.014763f
C1432 VTAIL.n85 VSUBS 0.067634f
C1433 VTAIL.n86 VSUBS 0.041307f
C1434 VTAIL.n87 VSUBS 0.326108f
C1435 VTAIL.t18 VSUBS 0.335869f
C1436 VTAIL.t10 VSUBS 0.335869f
C1437 VTAIL.n88 VSUBS 2.59127f
C1438 VTAIL.n89 VSUBS 0.982093f
C1439 VTAIL.t17 VSUBS 0.335869f
C1440 VTAIL.t16 VSUBS 0.335869f
C1441 VTAIL.n90 VSUBS 2.59127f
C1442 VTAIL.n91 VSUBS 2.7084f
C1443 VTAIL.t4 VSUBS 0.335869f
C1444 VTAIL.t7 VSUBS 0.335869f
C1445 VTAIL.n92 VSUBS 2.59129f
C1446 VTAIL.n93 VSUBS 2.70839f
C1447 VTAIL.t5 VSUBS 0.335869f
C1448 VTAIL.t3 VSUBS 0.335869f
C1449 VTAIL.n94 VSUBS 2.59129f
C1450 VTAIL.n95 VSUBS 0.982077f
C1451 VTAIL.n96 VSUBS 0.029491f
C1452 VTAIL.n97 VSUBS 0.027474f
C1453 VTAIL.n98 VSUBS 0.014763f
C1454 VTAIL.n99 VSUBS 0.034896f
C1455 VTAIL.n100 VSUBS 0.015198f
C1456 VTAIL.n101 VSUBS 0.027474f
C1457 VTAIL.n102 VSUBS 0.015198f
C1458 VTAIL.n103 VSUBS 0.014763f
C1459 VTAIL.n104 VSUBS 0.034896f
C1460 VTAIL.n105 VSUBS 0.034896f
C1461 VTAIL.n106 VSUBS 0.015632f
C1462 VTAIL.n107 VSUBS 0.027474f
C1463 VTAIL.n108 VSUBS 0.014763f
C1464 VTAIL.n109 VSUBS 0.034896f
C1465 VTAIL.n110 VSUBS 0.015632f
C1466 VTAIL.n111 VSUBS 0.027474f
C1467 VTAIL.n112 VSUBS 0.014763f
C1468 VTAIL.n113 VSUBS 0.034896f
C1469 VTAIL.n114 VSUBS 0.015632f
C1470 VTAIL.n115 VSUBS 0.027474f
C1471 VTAIL.n116 VSUBS 0.014763f
C1472 VTAIL.n117 VSUBS 0.034896f
C1473 VTAIL.n118 VSUBS 0.015632f
C1474 VTAIL.n119 VSUBS 0.027474f
C1475 VTAIL.n120 VSUBS 0.014763f
C1476 VTAIL.n121 VSUBS 0.034896f
C1477 VTAIL.n122 VSUBS 0.015632f
C1478 VTAIL.n123 VSUBS 1.81291f
C1479 VTAIL.n124 VSUBS 0.014763f
C1480 VTAIL.t0 VSUBS 0.074736f
C1481 VTAIL.n125 VSUBS 0.197478f
C1482 VTAIL.n126 VSUBS 0.022199f
C1483 VTAIL.n127 VSUBS 0.026172f
C1484 VTAIL.n128 VSUBS 0.034896f
C1485 VTAIL.n129 VSUBS 0.015632f
C1486 VTAIL.n130 VSUBS 0.014763f
C1487 VTAIL.n131 VSUBS 0.027474f
C1488 VTAIL.n132 VSUBS 0.027474f
C1489 VTAIL.n133 VSUBS 0.014763f
C1490 VTAIL.n134 VSUBS 0.015632f
C1491 VTAIL.n135 VSUBS 0.034896f
C1492 VTAIL.n136 VSUBS 0.034896f
C1493 VTAIL.n137 VSUBS 0.015632f
C1494 VTAIL.n138 VSUBS 0.014763f
C1495 VTAIL.n139 VSUBS 0.027474f
C1496 VTAIL.n140 VSUBS 0.027474f
C1497 VTAIL.n141 VSUBS 0.014763f
C1498 VTAIL.n142 VSUBS 0.015632f
C1499 VTAIL.n143 VSUBS 0.034896f
C1500 VTAIL.n144 VSUBS 0.034896f
C1501 VTAIL.n145 VSUBS 0.015632f
C1502 VTAIL.n146 VSUBS 0.014763f
C1503 VTAIL.n147 VSUBS 0.027474f
C1504 VTAIL.n148 VSUBS 0.027474f
C1505 VTAIL.n149 VSUBS 0.014763f
C1506 VTAIL.n150 VSUBS 0.015632f
C1507 VTAIL.n151 VSUBS 0.034896f
C1508 VTAIL.n152 VSUBS 0.034896f
C1509 VTAIL.n153 VSUBS 0.015632f
C1510 VTAIL.n154 VSUBS 0.014763f
C1511 VTAIL.n155 VSUBS 0.027474f
C1512 VTAIL.n156 VSUBS 0.027474f
C1513 VTAIL.n157 VSUBS 0.014763f
C1514 VTAIL.n158 VSUBS 0.015632f
C1515 VTAIL.n159 VSUBS 0.034896f
C1516 VTAIL.n160 VSUBS 0.034896f
C1517 VTAIL.n161 VSUBS 0.015632f
C1518 VTAIL.n162 VSUBS 0.014763f
C1519 VTAIL.n163 VSUBS 0.027474f
C1520 VTAIL.n164 VSUBS 0.027474f
C1521 VTAIL.n165 VSUBS 0.014763f
C1522 VTAIL.n166 VSUBS 0.015632f
C1523 VTAIL.n167 VSUBS 0.034896f
C1524 VTAIL.n168 VSUBS 0.034896f
C1525 VTAIL.n169 VSUBS 0.015632f
C1526 VTAIL.n170 VSUBS 0.014763f
C1527 VTAIL.n171 VSUBS 0.027474f
C1528 VTAIL.n172 VSUBS 0.027474f
C1529 VTAIL.n173 VSUBS 0.014763f
C1530 VTAIL.n174 VSUBS 0.015632f
C1531 VTAIL.n175 VSUBS 0.034896f
C1532 VTAIL.n176 VSUBS 0.082103f
C1533 VTAIL.n177 VSUBS 0.015632f
C1534 VTAIL.n178 VSUBS 0.014763f
C1535 VTAIL.n179 VSUBS 0.067634f
C1536 VTAIL.n180 VSUBS 0.041307f
C1537 VTAIL.n181 VSUBS 0.326108f
C1538 VTAIL.t12 VSUBS 0.335869f
C1539 VTAIL.t13 VSUBS 0.335869f
C1540 VTAIL.n182 VSUBS 2.59129f
C1541 VTAIL.n183 VSUBS 0.937431f
C1542 VTAIL.t11 VSUBS 0.335869f
C1543 VTAIL.t15 VSUBS 0.335869f
C1544 VTAIL.n184 VSUBS 2.59129f
C1545 VTAIL.n185 VSUBS 0.982077f
C1546 VTAIL.n186 VSUBS 0.029491f
C1547 VTAIL.n187 VSUBS 0.027474f
C1548 VTAIL.n188 VSUBS 0.014763f
C1549 VTAIL.n189 VSUBS 0.034896f
C1550 VTAIL.n190 VSUBS 0.015198f
C1551 VTAIL.n191 VSUBS 0.027474f
C1552 VTAIL.n192 VSUBS 0.015198f
C1553 VTAIL.n193 VSUBS 0.014763f
C1554 VTAIL.n194 VSUBS 0.034896f
C1555 VTAIL.n195 VSUBS 0.034896f
C1556 VTAIL.n196 VSUBS 0.015632f
C1557 VTAIL.n197 VSUBS 0.027474f
C1558 VTAIL.n198 VSUBS 0.014763f
C1559 VTAIL.n199 VSUBS 0.034896f
C1560 VTAIL.n200 VSUBS 0.015632f
C1561 VTAIL.n201 VSUBS 0.027474f
C1562 VTAIL.n202 VSUBS 0.014763f
C1563 VTAIL.n203 VSUBS 0.034896f
C1564 VTAIL.n204 VSUBS 0.015632f
C1565 VTAIL.n205 VSUBS 0.027474f
C1566 VTAIL.n206 VSUBS 0.014763f
C1567 VTAIL.n207 VSUBS 0.034896f
C1568 VTAIL.n208 VSUBS 0.015632f
C1569 VTAIL.n209 VSUBS 0.027474f
C1570 VTAIL.n210 VSUBS 0.014763f
C1571 VTAIL.n211 VSUBS 0.034896f
C1572 VTAIL.n212 VSUBS 0.015632f
C1573 VTAIL.n213 VSUBS 1.81291f
C1574 VTAIL.n214 VSUBS 0.014763f
C1575 VTAIL.t14 VSUBS 0.074736f
C1576 VTAIL.n215 VSUBS 0.197478f
C1577 VTAIL.n216 VSUBS 0.022199f
C1578 VTAIL.n217 VSUBS 0.026172f
C1579 VTAIL.n218 VSUBS 0.034896f
C1580 VTAIL.n219 VSUBS 0.015632f
C1581 VTAIL.n220 VSUBS 0.014763f
C1582 VTAIL.n221 VSUBS 0.027474f
C1583 VTAIL.n222 VSUBS 0.027474f
C1584 VTAIL.n223 VSUBS 0.014763f
C1585 VTAIL.n224 VSUBS 0.015632f
C1586 VTAIL.n225 VSUBS 0.034896f
C1587 VTAIL.n226 VSUBS 0.034896f
C1588 VTAIL.n227 VSUBS 0.015632f
C1589 VTAIL.n228 VSUBS 0.014763f
C1590 VTAIL.n229 VSUBS 0.027474f
C1591 VTAIL.n230 VSUBS 0.027474f
C1592 VTAIL.n231 VSUBS 0.014763f
C1593 VTAIL.n232 VSUBS 0.015632f
C1594 VTAIL.n233 VSUBS 0.034896f
C1595 VTAIL.n234 VSUBS 0.034896f
C1596 VTAIL.n235 VSUBS 0.015632f
C1597 VTAIL.n236 VSUBS 0.014763f
C1598 VTAIL.n237 VSUBS 0.027474f
C1599 VTAIL.n238 VSUBS 0.027474f
C1600 VTAIL.n239 VSUBS 0.014763f
C1601 VTAIL.n240 VSUBS 0.015632f
C1602 VTAIL.n241 VSUBS 0.034896f
C1603 VTAIL.n242 VSUBS 0.034896f
C1604 VTAIL.n243 VSUBS 0.015632f
C1605 VTAIL.n244 VSUBS 0.014763f
C1606 VTAIL.n245 VSUBS 0.027474f
C1607 VTAIL.n246 VSUBS 0.027474f
C1608 VTAIL.n247 VSUBS 0.014763f
C1609 VTAIL.n248 VSUBS 0.015632f
C1610 VTAIL.n249 VSUBS 0.034896f
C1611 VTAIL.n250 VSUBS 0.034896f
C1612 VTAIL.n251 VSUBS 0.015632f
C1613 VTAIL.n252 VSUBS 0.014763f
C1614 VTAIL.n253 VSUBS 0.027474f
C1615 VTAIL.n254 VSUBS 0.027474f
C1616 VTAIL.n255 VSUBS 0.014763f
C1617 VTAIL.n256 VSUBS 0.015632f
C1618 VTAIL.n257 VSUBS 0.034896f
C1619 VTAIL.n258 VSUBS 0.034896f
C1620 VTAIL.n259 VSUBS 0.015632f
C1621 VTAIL.n260 VSUBS 0.014763f
C1622 VTAIL.n261 VSUBS 0.027474f
C1623 VTAIL.n262 VSUBS 0.027474f
C1624 VTAIL.n263 VSUBS 0.014763f
C1625 VTAIL.n264 VSUBS 0.015632f
C1626 VTAIL.n265 VSUBS 0.034896f
C1627 VTAIL.n266 VSUBS 0.082103f
C1628 VTAIL.n267 VSUBS 0.015632f
C1629 VTAIL.n268 VSUBS 0.014763f
C1630 VTAIL.n269 VSUBS 0.067634f
C1631 VTAIL.n270 VSUBS 0.041307f
C1632 VTAIL.n271 VSUBS 1.92459f
C1633 VTAIL.n272 VSUBS 0.029491f
C1634 VTAIL.n273 VSUBS 0.027474f
C1635 VTAIL.n274 VSUBS 0.014763f
C1636 VTAIL.n275 VSUBS 0.034896f
C1637 VTAIL.n276 VSUBS 0.015198f
C1638 VTAIL.n277 VSUBS 0.027474f
C1639 VTAIL.n278 VSUBS 0.015632f
C1640 VTAIL.n279 VSUBS 0.034896f
C1641 VTAIL.n280 VSUBS 0.015632f
C1642 VTAIL.n281 VSUBS 0.027474f
C1643 VTAIL.n282 VSUBS 0.014763f
C1644 VTAIL.n283 VSUBS 0.034896f
C1645 VTAIL.n284 VSUBS 0.015632f
C1646 VTAIL.n285 VSUBS 0.027474f
C1647 VTAIL.n286 VSUBS 0.014763f
C1648 VTAIL.n287 VSUBS 0.034896f
C1649 VTAIL.n288 VSUBS 0.015632f
C1650 VTAIL.n289 VSUBS 0.027474f
C1651 VTAIL.n290 VSUBS 0.014763f
C1652 VTAIL.n291 VSUBS 0.034896f
C1653 VTAIL.n292 VSUBS 0.015632f
C1654 VTAIL.n293 VSUBS 0.027474f
C1655 VTAIL.n294 VSUBS 0.014763f
C1656 VTAIL.n295 VSUBS 0.034896f
C1657 VTAIL.n296 VSUBS 0.015632f
C1658 VTAIL.n297 VSUBS 1.81291f
C1659 VTAIL.n298 VSUBS 0.014763f
C1660 VTAIL.t6 VSUBS 0.074736f
C1661 VTAIL.n299 VSUBS 0.197478f
C1662 VTAIL.n300 VSUBS 0.022199f
C1663 VTAIL.n301 VSUBS 0.026172f
C1664 VTAIL.n302 VSUBS 0.034896f
C1665 VTAIL.n303 VSUBS 0.015632f
C1666 VTAIL.n304 VSUBS 0.014763f
C1667 VTAIL.n305 VSUBS 0.027474f
C1668 VTAIL.n306 VSUBS 0.027474f
C1669 VTAIL.n307 VSUBS 0.014763f
C1670 VTAIL.n308 VSUBS 0.015632f
C1671 VTAIL.n309 VSUBS 0.034896f
C1672 VTAIL.n310 VSUBS 0.034896f
C1673 VTAIL.n311 VSUBS 0.015632f
C1674 VTAIL.n312 VSUBS 0.014763f
C1675 VTAIL.n313 VSUBS 0.027474f
C1676 VTAIL.n314 VSUBS 0.027474f
C1677 VTAIL.n315 VSUBS 0.014763f
C1678 VTAIL.n316 VSUBS 0.015632f
C1679 VTAIL.n317 VSUBS 0.034896f
C1680 VTAIL.n318 VSUBS 0.034896f
C1681 VTAIL.n319 VSUBS 0.015632f
C1682 VTAIL.n320 VSUBS 0.014763f
C1683 VTAIL.n321 VSUBS 0.027474f
C1684 VTAIL.n322 VSUBS 0.027474f
C1685 VTAIL.n323 VSUBS 0.014763f
C1686 VTAIL.n324 VSUBS 0.015632f
C1687 VTAIL.n325 VSUBS 0.034896f
C1688 VTAIL.n326 VSUBS 0.034896f
C1689 VTAIL.n327 VSUBS 0.015632f
C1690 VTAIL.n328 VSUBS 0.014763f
C1691 VTAIL.n329 VSUBS 0.027474f
C1692 VTAIL.n330 VSUBS 0.027474f
C1693 VTAIL.n331 VSUBS 0.014763f
C1694 VTAIL.n332 VSUBS 0.015632f
C1695 VTAIL.n333 VSUBS 0.034896f
C1696 VTAIL.n334 VSUBS 0.034896f
C1697 VTAIL.n335 VSUBS 0.015632f
C1698 VTAIL.n336 VSUBS 0.014763f
C1699 VTAIL.n337 VSUBS 0.027474f
C1700 VTAIL.n338 VSUBS 0.027474f
C1701 VTAIL.n339 VSUBS 0.014763f
C1702 VTAIL.n340 VSUBS 0.014763f
C1703 VTAIL.n341 VSUBS 0.015632f
C1704 VTAIL.n342 VSUBS 0.034896f
C1705 VTAIL.n343 VSUBS 0.034896f
C1706 VTAIL.n344 VSUBS 0.034896f
C1707 VTAIL.n345 VSUBS 0.015198f
C1708 VTAIL.n346 VSUBS 0.014763f
C1709 VTAIL.n347 VSUBS 0.027474f
C1710 VTAIL.n348 VSUBS 0.027474f
C1711 VTAIL.n349 VSUBS 0.014763f
C1712 VTAIL.n350 VSUBS 0.015632f
C1713 VTAIL.n351 VSUBS 0.034896f
C1714 VTAIL.n352 VSUBS 0.082103f
C1715 VTAIL.n353 VSUBS 0.015632f
C1716 VTAIL.n354 VSUBS 0.014763f
C1717 VTAIL.n355 VSUBS 0.067634f
C1718 VTAIL.n356 VSUBS 0.041307f
C1719 VTAIL.n357 VSUBS 1.92459f
C1720 VTAIL.t1 VSUBS 0.335869f
C1721 VTAIL.t9 VSUBS 0.335869f
C1722 VTAIL.n358 VSUBS 2.59127f
C1723 VTAIL.n359 VSUBS 0.847583f
C1724 VP.n0 VSUBS 0.031743f
C1725 VP.t6 VSUBS 2.59885f
C1726 VP.n1 VSUBS 0.030964f
C1727 VP.n2 VSUBS 0.031743f
C1728 VP.t3 VSUBS 2.59885f
C1729 VP.n3 VSUBS 0.056323f
C1730 VP.n4 VSUBS 0.031743f
C1731 VP.t2 VSUBS 2.59885f
C1732 VP.n5 VSUBS 0.062224f
C1733 VP.n6 VSUBS 0.031743f
C1734 VP.t1 VSUBS 2.59885f
C1735 VP.n7 VSUBS 0.914568f
C1736 VP.n8 VSUBS 0.031743f
C1737 VP.n9 VSUBS 0.063242f
C1738 VP.n10 VSUBS 0.031743f
C1739 VP.t4 VSUBS 2.59885f
C1740 VP.n11 VSUBS 0.030964f
C1741 VP.n12 VSUBS 0.031743f
C1742 VP.t5 VSUBS 2.59885f
C1743 VP.n13 VSUBS 0.056323f
C1744 VP.n14 VSUBS 0.031743f
C1745 VP.t8 VSUBS 2.59885f
C1746 VP.n15 VSUBS 0.062224f
C1747 VP.n16 VSUBS 0.031743f
C1748 VP.t7 VSUBS 2.59885f
C1749 VP.n17 VSUBS 0.989261f
C1750 VP.t9 VSUBS 2.75166f
C1751 VP.n18 VSUBS 0.99497f
C1752 VP.n19 VSUBS 0.235875f
C1753 VP.n20 VSUBS 0.045142f
C1754 VP.n21 VSUBS 0.056323f
C1755 VP.n22 VSUBS 0.033294f
C1756 VP.n23 VSUBS 0.031743f
C1757 VP.n24 VSUBS 0.031743f
C1758 VP.n25 VSUBS 0.031743f
C1759 VP.n26 VSUBS 0.944521f
C1760 VP.n27 VSUBS 0.062224f
C1761 VP.n28 VSUBS 0.033294f
C1762 VP.n29 VSUBS 0.031743f
C1763 VP.n30 VSUBS 0.031743f
C1764 VP.n31 VSUBS 0.031743f
C1765 VP.n32 VSUBS 0.045142f
C1766 VP.n33 VSUBS 0.914568f
C1767 VP.n34 VSUBS 0.043973f
C1768 VP.n35 VSUBS 0.057634f
C1769 VP.n36 VSUBS 0.031743f
C1770 VP.n37 VSUBS 0.031743f
C1771 VP.n38 VSUBS 0.031743f
C1772 VP.n39 VSUBS 0.063242f
C1773 VP.n40 VSUBS 0.031121f
C1774 VP.n41 VSUBS 0.989156f
C1775 VP.n42 VSUBS 1.84005f
C1776 VP.n43 VSUBS 1.862f
C1777 VP.t0 VSUBS 2.59885f
C1778 VP.n44 VSUBS 0.989156f
C1779 VP.n45 VSUBS 0.031121f
C1780 VP.n46 VSUBS 0.031743f
C1781 VP.n47 VSUBS 0.031743f
C1782 VP.n48 VSUBS 0.031743f
C1783 VP.n49 VSUBS 0.030964f
C1784 VP.n50 VSUBS 0.057634f
C1785 VP.n51 VSUBS 0.043973f
C1786 VP.n52 VSUBS 0.031743f
C1787 VP.n53 VSUBS 0.031743f
C1788 VP.n54 VSUBS 0.045142f
C1789 VP.n55 VSUBS 0.056323f
C1790 VP.n56 VSUBS 0.033294f
C1791 VP.n57 VSUBS 0.031743f
C1792 VP.n58 VSUBS 0.031743f
C1793 VP.n59 VSUBS 0.031743f
C1794 VP.n60 VSUBS 0.944521f
C1795 VP.n61 VSUBS 0.062224f
C1796 VP.n62 VSUBS 0.033294f
C1797 VP.n63 VSUBS 0.031743f
C1798 VP.n64 VSUBS 0.031743f
C1799 VP.n65 VSUBS 0.031743f
C1800 VP.n66 VSUBS 0.045142f
C1801 VP.n67 VSUBS 0.914568f
C1802 VP.n68 VSUBS 0.043973f
C1803 VP.n69 VSUBS 0.057634f
C1804 VP.n70 VSUBS 0.031743f
C1805 VP.n71 VSUBS 0.031743f
C1806 VP.n72 VSUBS 0.031743f
C1807 VP.n73 VSUBS 0.063242f
C1808 VP.n74 VSUBS 0.031121f
C1809 VP.n75 VSUBS 0.989156f
C1810 VP.n76 VSUBS 0.035461f
.ends

