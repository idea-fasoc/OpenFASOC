* NGSPICE file created from diff_pair_sample_1725.ext - technology: sky130A

.subckt diff_pair_sample_1725 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=0 ps=0 w=16.44 l=3.25
X1 VTAIL.t7 VN.t0 VDD2.t0 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=2.7126 ps=16.77 w=16.44 l=3.25
X2 VDD1.t3 VP.t0 VTAIL.t1 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=2.7126 pd=16.77 as=6.4116 ps=33.66 w=16.44 l=3.25
X3 VTAIL.t6 VN.t1 VDD2.t3 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=2.7126 ps=16.77 w=16.44 l=3.25
X4 VTAIL.t3 VP.t1 VDD1.t2 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=2.7126 ps=16.77 w=16.44 l=3.25
X5 VDD2.t1 VN.t2 VTAIL.t5 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=2.7126 pd=16.77 as=6.4116 ps=33.66 w=16.44 l=3.25
X6 B.t8 B.t6 B.t7 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=0 ps=0 w=16.44 l=3.25
X7 VDD1.t1 VP.t2 VTAIL.t0 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=2.7126 pd=16.77 as=6.4116 ps=33.66 w=16.44 l=3.25
X8 B.t5 B.t3 B.t4 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=0 ps=0 w=16.44 l=3.25
X9 B.t2 B.t0 B.t1 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=0 ps=0 w=16.44 l=3.25
X10 VDD2.t2 VN.t3 VTAIL.t4 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=2.7126 pd=16.77 as=6.4116 ps=33.66 w=16.44 l=3.25
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n3118_n4256# sky130_fd_pr__pfet_01v8 ad=6.4116 pd=33.66 as=2.7126 ps=16.77 w=16.44 l=3.25
R0 B.n444 B.n125 585
R1 B.n443 B.n442 585
R2 B.n441 B.n126 585
R3 B.n440 B.n439 585
R4 B.n438 B.n127 585
R5 B.n437 B.n436 585
R6 B.n435 B.n128 585
R7 B.n434 B.n433 585
R8 B.n432 B.n129 585
R9 B.n431 B.n430 585
R10 B.n429 B.n130 585
R11 B.n428 B.n427 585
R12 B.n426 B.n131 585
R13 B.n425 B.n424 585
R14 B.n423 B.n132 585
R15 B.n422 B.n421 585
R16 B.n420 B.n133 585
R17 B.n419 B.n418 585
R18 B.n417 B.n134 585
R19 B.n416 B.n415 585
R20 B.n414 B.n135 585
R21 B.n413 B.n412 585
R22 B.n411 B.n136 585
R23 B.n410 B.n409 585
R24 B.n408 B.n137 585
R25 B.n407 B.n406 585
R26 B.n405 B.n138 585
R27 B.n404 B.n403 585
R28 B.n402 B.n139 585
R29 B.n401 B.n400 585
R30 B.n399 B.n140 585
R31 B.n398 B.n397 585
R32 B.n396 B.n141 585
R33 B.n395 B.n394 585
R34 B.n393 B.n142 585
R35 B.n392 B.n391 585
R36 B.n390 B.n143 585
R37 B.n389 B.n388 585
R38 B.n387 B.n144 585
R39 B.n386 B.n385 585
R40 B.n384 B.n145 585
R41 B.n383 B.n382 585
R42 B.n381 B.n146 585
R43 B.n380 B.n379 585
R44 B.n378 B.n147 585
R45 B.n377 B.n376 585
R46 B.n375 B.n148 585
R47 B.n374 B.n373 585
R48 B.n372 B.n149 585
R49 B.n371 B.n370 585
R50 B.n369 B.n150 585
R51 B.n368 B.n367 585
R52 B.n366 B.n151 585
R53 B.n365 B.n364 585
R54 B.n363 B.n152 585
R55 B.n362 B.n361 585
R56 B.n357 B.n153 585
R57 B.n356 B.n355 585
R58 B.n354 B.n154 585
R59 B.n353 B.n352 585
R60 B.n351 B.n155 585
R61 B.n350 B.n349 585
R62 B.n348 B.n156 585
R63 B.n347 B.n346 585
R64 B.n344 B.n157 585
R65 B.n343 B.n342 585
R66 B.n341 B.n160 585
R67 B.n340 B.n339 585
R68 B.n338 B.n161 585
R69 B.n337 B.n336 585
R70 B.n335 B.n162 585
R71 B.n334 B.n333 585
R72 B.n332 B.n163 585
R73 B.n331 B.n330 585
R74 B.n329 B.n164 585
R75 B.n328 B.n327 585
R76 B.n326 B.n165 585
R77 B.n325 B.n324 585
R78 B.n323 B.n166 585
R79 B.n322 B.n321 585
R80 B.n320 B.n167 585
R81 B.n319 B.n318 585
R82 B.n317 B.n168 585
R83 B.n316 B.n315 585
R84 B.n314 B.n169 585
R85 B.n313 B.n312 585
R86 B.n311 B.n170 585
R87 B.n310 B.n309 585
R88 B.n308 B.n171 585
R89 B.n307 B.n306 585
R90 B.n305 B.n172 585
R91 B.n304 B.n303 585
R92 B.n302 B.n173 585
R93 B.n301 B.n300 585
R94 B.n299 B.n174 585
R95 B.n298 B.n297 585
R96 B.n296 B.n175 585
R97 B.n295 B.n294 585
R98 B.n293 B.n176 585
R99 B.n292 B.n291 585
R100 B.n290 B.n177 585
R101 B.n289 B.n288 585
R102 B.n287 B.n178 585
R103 B.n286 B.n285 585
R104 B.n284 B.n179 585
R105 B.n283 B.n282 585
R106 B.n281 B.n180 585
R107 B.n280 B.n279 585
R108 B.n278 B.n181 585
R109 B.n277 B.n276 585
R110 B.n275 B.n182 585
R111 B.n274 B.n273 585
R112 B.n272 B.n183 585
R113 B.n271 B.n270 585
R114 B.n269 B.n184 585
R115 B.n268 B.n267 585
R116 B.n266 B.n185 585
R117 B.n265 B.n264 585
R118 B.n263 B.n186 585
R119 B.n446 B.n445 585
R120 B.n447 B.n124 585
R121 B.n449 B.n448 585
R122 B.n450 B.n123 585
R123 B.n452 B.n451 585
R124 B.n453 B.n122 585
R125 B.n455 B.n454 585
R126 B.n456 B.n121 585
R127 B.n458 B.n457 585
R128 B.n459 B.n120 585
R129 B.n461 B.n460 585
R130 B.n462 B.n119 585
R131 B.n464 B.n463 585
R132 B.n465 B.n118 585
R133 B.n467 B.n466 585
R134 B.n468 B.n117 585
R135 B.n470 B.n469 585
R136 B.n471 B.n116 585
R137 B.n473 B.n472 585
R138 B.n474 B.n115 585
R139 B.n476 B.n475 585
R140 B.n477 B.n114 585
R141 B.n479 B.n478 585
R142 B.n480 B.n113 585
R143 B.n482 B.n481 585
R144 B.n483 B.n112 585
R145 B.n485 B.n484 585
R146 B.n486 B.n111 585
R147 B.n488 B.n487 585
R148 B.n489 B.n110 585
R149 B.n491 B.n490 585
R150 B.n492 B.n109 585
R151 B.n494 B.n493 585
R152 B.n495 B.n108 585
R153 B.n497 B.n496 585
R154 B.n498 B.n107 585
R155 B.n500 B.n499 585
R156 B.n501 B.n106 585
R157 B.n503 B.n502 585
R158 B.n504 B.n105 585
R159 B.n506 B.n505 585
R160 B.n507 B.n104 585
R161 B.n509 B.n508 585
R162 B.n510 B.n103 585
R163 B.n512 B.n511 585
R164 B.n513 B.n102 585
R165 B.n515 B.n514 585
R166 B.n516 B.n101 585
R167 B.n518 B.n517 585
R168 B.n519 B.n100 585
R169 B.n521 B.n520 585
R170 B.n522 B.n99 585
R171 B.n524 B.n523 585
R172 B.n525 B.n98 585
R173 B.n527 B.n526 585
R174 B.n528 B.n97 585
R175 B.n530 B.n529 585
R176 B.n531 B.n96 585
R177 B.n533 B.n532 585
R178 B.n534 B.n95 585
R179 B.n536 B.n535 585
R180 B.n537 B.n94 585
R181 B.n539 B.n538 585
R182 B.n540 B.n93 585
R183 B.n542 B.n541 585
R184 B.n543 B.n92 585
R185 B.n545 B.n544 585
R186 B.n546 B.n91 585
R187 B.n548 B.n547 585
R188 B.n549 B.n90 585
R189 B.n551 B.n550 585
R190 B.n552 B.n89 585
R191 B.n554 B.n553 585
R192 B.n555 B.n88 585
R193 B.n557 B.n556 585
R194 B.n558 B.n87 585
R195 B.n560 B.n559 585
R196 B.n561 B.n86 585
R197 B.n563 B.n562 585
R198 B.n564 B.n85 585
R199 B.n745 B.n744 585
R200 B.n743 B.n22 585
R201 B.n742 B.n741 585
R202 B.n740 B.n23 585
R203 B.n739 B.n738 585
R204 B.n737 B.n24 585
R205 B.n736 B.n735 585
R206 B.n734 B.n25 585
R207 B.n733 B.n732 585
R208 B.n731 B.n26 585
R209 B.n730 B.n729 585
R210 B.n728 B.n27 585
R211 B.n727 B.n726 585
R212 B.n725 B.n28 585
R213 B.n724 B.n723 585
R214 B.n722 B.n29 585
R215 B.n721 B.n720 585
R216 B.n719 B.n30 585
R217 B.n718 B.n717 585
R218 B.n716 B.n31 585
R219 B.n715 B.n714 585
R220 B.n713 B.n32 585
R221 B.n712 B.n711 585
R222 B.n710 B.n33 585
R223 B.n709 B.n708 585
R224 B.n707 B.n34 585
R225 B.n706 B.n705 585
R226 B.n704 B.n35 585
R227 B.n703 B.n702 585
R228 B.n701 B.n36 585
R229 B.n700 B.n699 585
R230 B.n698 B.n37 585
R231 B.n697 B.n696 585
R232 B.n695 B.n38 585
R233 B.n694 B.n693 585
R234 B.n692 B.n39 585
R235 B.n691 B.n690 585
R236 B.n689 B.n40 585
R237 B.n688 B.n687 585
R238 B.n686 B.n41 585
R239 B.n685 B.n684 585
R240 B.n683 B.n42 585
R241 B.n682 B.n681 585
R242 B.n680 B.n43 585
R243 B.n679 B.n678 585
R244 B.n677 B.n44 585
R245 B.n676 B.n675 585
R246 B.n674 B.n45 585
R247 B.n673 B.n672 585
R248 B.n671 B.n46 585
R249 B.n670 B.n669 585
R250 B.n668 B.n47 585
R251 B.n667 B.n666 585
R252 B.n665 B.n48 585
R253 B.n664 B.n663 585
R254 B.n661 B.n49 585
R255 B.n660 B.n659 585
R256 B.n658 B.n52 585
R257 B.n657 B.n656 585
R258 B.n655 B.n53 585
R259 B.n654 B.n653 585
R260 B.n652 B.n54 585
R261 B.n651 B.n650 585
R262 B.n649 B.n55 585
R263 B.n647 B.n646 585
R264 B.n645 B.n58 585
R265 B.n644 B.n643 585
R266 B.n642 B.n59 585
R267 B.n641 B.n640 585
R268 B.n639 B.n60 585
R269 B.n638 B.n637 585
R270 B.n636 B.n61 585
R271 B.n635 B.n634 585
R272 B.n633 B.n62 585
R273 B.n632 B.n631 585
R274 B.n630 B.n63 585
R275 B.n629 B.n628 585
R276 B.n627 B.n64 585
R277 B.n626 B.n625 585
R278 B.n624 B.n65 585
R279 B.n623 B.n622 585
R280 B.n621 B.n66 585
R281 B.n620 B.n619 585
R282 B.n618 B.n67 585
R283 B.n617 B.n616 585
R284 B.n615 B.n68 585
R285 B.n614 B.n613 585
R286 B.n612 B.n69 585
R287 B.n611 B.n610 585
R288 B.n609 B.n70 585
R289 B.n608 B.n607 585
R290 B.n606 B.n71 585
R291 B.n605 B.n604 585
R292 B.n603 B.n72 585
R293 B.n602 B.n601 585
R294 B.n600 B.n73 585
R295 B.n599 B.n598 585
R296 B.n597 B.n74 585
R297 B.n596 B.n595 585
R298 B.n594 B.n75 585
R299 B.n593 B.n592 585
R300 B.n591 B.n76 585
R301 B.n590 B.n589 585
R302 B.n588 B.n77 585
R303 B.n587 B.n586 585
R304 B.n585 B.n78 585
R305 B.n584 B.n583 585
R306 B.n582 B.n79 585
R307 B.n581 B.n580 585
R308 B.n579 B.n80 585
R309 B.n578 B.n577 585
R310 B.n576 B.n81 585
R311 B.n575 B.n574 585
R312 B.n573 B.n82 585
R313 B.n572 B.n571 585
R314 B.n570 B.n83 585
R315 B.n569 B.n568 585
R316 B.n567 B.n84 585
R317 B.n566 B.n565 585
R318 B.n746 B.n21 585
R319 B.n748 B.n747 585
R320 B.n749 B.n20 585
R321 B.n751 B.n750 585
R322 B.n752 B.n19 585
R323 B.n754 B.n753 585
R324 B.n755 B.n18 585
R325 B.n757 B.n756 585
R326 B.n758 B.n17 585
R327 B.n760 B.n759 585
R328 B.n761 B.n16 585
R329 B.n763 B.n762 585
R330 B.n764 B.n15 585
R331 B.n766 B.n765 585
R332 B.n767 B.n14 585
R333 B.n769 B.n768 585
R334 B.n770 B.n13 585
R335 B.n772 B.n771 585
R336 B.n773 B.n12 585
R337 B.n775 B.n774 585
R338 B.n776 B.n11 585
R339 B.n778 B.n777 585
R340 B.n779 B.n10 585
R341 B.n781 B.n780 585
R342 B.n782 B.n9 585
R343 B.n784 B.n783 585
R344 B.n785 B.n8 585
R345 B.n787 B.n786 585
R346 B.n788 B.n7 585
R347 B.n790 B.n789 585
R348 B.n791 B.n6 585
R349 B.n793 B.n792 585
R350 B.n794 B.n5 585
R351 B.n796 B.n795 585
R352 B.n797 B.n4 585
R353 B.n799 B.n798 585
R354 B.n800 B.n3 585
R355 B.n802 B.n801 585
R356 B.n803 B.n0 585
R357 B.n2 B.n1 585
R358 B.n206 B.n205 585
R359 B.n208 B.n207 585
R360 B.n209 B.n204 585
R361 B.n211 B.n210 585
R362 B.n212 B.n203 585
R363 B.n214 B.n213 585
R364 B.n215 B.n202 585
R365 B.n217 B.n216 585
R366 B.n218 B.n201 585
R367 B.n220 B.n219 585
R368 B.n221 B.n200 585
R369 B.n223 B.n222 585
R370 B.n224 B.n199 585
R371 B.n226 B.n225 585
R372 B.n227 B.n198 585
R373 B.n229 B.n228 585
R374 B.n230 B.n197 585
R375 B.n232 B.n231 585
R376 B.n233 B.n196 585
R377 B.n235 B.n234 585
R378 B.n236 B.n195 585
R379 B.n238 B.n237 585
R380 B.n239 B.n194 585
R381 B.n241 B.n240 585
R382 B.n242 B.n193 585
R383 B.n244 B.n243 585
R384 B.n245 B.n192 585
R385 B.n247 B.n246 585
R386 B.n248 B.n191 585
R387 B.n250 B.n249 585
R388 B.n251 B.n190 585
R389 B.n253 B.n252 585
R390 B.n254 B.n189 585
R391 B.n256 B.n255 585
R392 B.n257 B.n188 585
R393 B.n259 B.n258 585
R394 B.n260 B.n187 585
R395 B.n262 B.n261 585
R396 B.n263 B.n262 526.135
R397 B.n446 B.n125 526.135
R398 B.n566 B.n85 526.135
R399 B.n744 B.n21 526.135
R400 B.n158 B.t9 330.764
R401 B.n358 B.t3 330.764
R402 B.n56 B.t0 330.764
R403 B.n50 B.t6 330.764
R404 B.n805 B.n804 256.663
R405 B.n804 B.n803 235.042
R406 B.n804 B.n2 235.042
R407 B.n358 B.t4 178.131
R408 B.n56 B.t2 178.131
R409 B.n158 B.t10 178.109
R410 B.n50 B.t8 178.109
R411 B.n264 B.n263 163.367
R412 B.n264 B.n185 163.367
R413 B.n268 B.n185 163.367
R414 B.n269 B.n268 163.367
R415 B.n270 B.n269 163.367
R416 B.n270 B.n183 163.367
R417 B.n274 B.n183 163.367
R418 B.n275 B.n274 163.367
R419 B.n276 B.n275 163.367
R420 B.n276 B.n181 163.367
R421 B.n280 B.n181 163.367
R422 B.n281 B.n280 163.367
R423 B.n282 B.n281 163.367
R424 B.n282 B.n179 163.367
R425 B.n286 B.n179 163.367
R426 B.n287 B.n286 163.367
R427 B.n288 B.n287 163.367
R428 B.n288 B.n177 163.367
R429 B.n292 B.n177 163.367
R430 B.n293 B.n292 163.367
R431 B.n294 B.n293 163.367
R432 B.n294 B.n175 163.367
R433 B.n298 B.n175 163.367
R434 B.n299 B.n298 163.367
R435 B.n300 B.n299 163.367
R436 B.n300 B.n173 163.367
R437 B.n304 B.n173 163.367
R438 B.n305 B.n304 163.367
R439 B.n306 B.n305 163.367
R440 B.n306 B.n171 163.367
R441 B.n310 B.n171 163.367
R442 B.n311 B.n310 163.367
R443 B.n312 B.n311 163.367
R444 B.n312 B.n169 163.367
R445 B.n316 B.n169 163.367
R446 B.n317 B.n316 163.367
R447 B.n318 B.n317 163.367
R448 B.n318 B.n167 163.367
R449 B.n322 B.n167 163.367
R450 B.n323 B.n322 163.367
R451 B.n324 B.n323 163.367
R452 B.n324 B.n165 163.367
R453 B.n328 B.n165 163.367
R454 B.n329 B.n328 163.367
R455 B.n330 B.n329 163.367
R456 B.n330 B.n163 163.367
R457 B.n334 B.n163 163.367
R458 B.n335 B.n334 163.367
R459 B.n336 B.n335 163.367
R460 B.n336 B.n161 163.367
R461 B.n340 B.n161 163.367
R462 B.n341 B.n340 163.367
R463 B.n342 B.n341 163.367
R464 B.n342 B.n157 163.367
R465 B.n347 B.n157 163.367
R466 B.n348 B.n347 163.367
R467 B.n349 B.n348 163.367
R468 B.n349 B.n155 163.367
R469 B.n353 B.n155 163.367
R470 B.n354 B.n353 163.367
R471 B.n355 B.n354 163.367
R472 B.n355 B.n153 163.367
R473 B.n362 B.n153 163.367
R474 B.n363 B.n362 163.367
R475 B.n364 B.n363 163.367
R476 B.n364 B.n151 163.367
R477 B.n368 B.n151 163.367
R478 B.n369 B.n368 163.367
R479 B.n370 B.n369 163.367
R480 B.n370 B.n149 163.367
R481 B.n374 B.n149 163.367
R482 B.n375 B.n374 163.367
R483 B.n376 B.n375 163.367
R484 B.n376 B.n147 163.367
R485 B.n380 B.n147 163.367
R486 B.n381 B.n380 163.367
R487 B.n382 B.n381 163.367
R488 B.n382 B.n145 163.367
R489 B.n386 B.n145 163.367
R490 B.n387 B.n386 163.367
R491 B.n388 B.n387 163.367
R492 B.n388 B.n143 163.367
R493 B.n392 B.n143 163.367
R494 B.n393 B.n392 163.367
R495 B.n394 B.n393 163.367
R496 B.n394 B.n141 163.367
R497 B.n398 B.n141 163.367
R498 B.n399 B.n398 163.367
R499 B.n400 B.n399 163.367
R500 B.n400 B.n139 163.367
R501 B.n404 B.n139 163.367
R502 B.n405 B.n404 163.367
R503 B.n406 B.n405 163.367
R504 B.n406 B.n137 163.367
R505 B.n410 B.n137 163.367
R506 B.n411 B.n410 163.367
R507 B.n412 B.n411 163.367
R508 B.n412 B.n135 163.367
R509 B.n416 B.n135 163.367
R510 B.n417 B.n416 163.367
R511 B.n418 B.n417 163.367
R512 B.n418 B.n133 163.367
R513 B.n422 B.n133 163.367
R514 B.n423 B.n422 163.367
R515 B.n424 B.n423 163.367
R516 B.n424 B.n131 163.367
R517 B.n428 B.n131 163.367
R518 B.n429 B.n428 163.367
R519 B.n430 B.n429 163.367
R520 B.n430 B.n129 163.367
R521 B.n434 B.n129 163.367
R522 B.n435 B.n434 163.367
R523 B.n436 B.n435 163.367
R524 B.n436 B.n127 163.367
R525 B.n440 B.n127 163.367
R526 B.n441 B.n440 163.367
R527 B.n442 B.n441 163.367
R528 B.n442 B.n125 163.367
R529 B.n562 B.n85 163.367
R530 B.n562 B.n561 163.367
R531 B.n561 B.n560 163.367
R532 B.n560 B.n87 163.367
R533 B.n556 B.n87 163.367
R534 B.n556 B.n555 163.367
R535 B.n555 B.n554 163.367
R536 B.n554 B.n89 163.367
R537 B.n550 B.n89 163.367
R538 B.n550 B.n549 163.367
R539 B.n549 B.n548 163.367
R540 B.n548 B.n91 163.367
R541 B.n544 B.n91 163.367
R542 B.n544 B.n543 163.367
R543 B.n543 B.n542 163.367
R544 B.n542 B.n93 163.367
R545 B.n538 B.n93 163.367
R546 B.n538 B.n537 163.367
R547 B.n537 B.n536 163.367
R548 B.n536 B.n95 163.367
R549 B.n532 B.n95 163.367
R550 B.n532 B.n531 163.367
R551 B.n531 B.n530 163.367
R552 B.n530 B.n97 163.367
R553 B.n526 B.n97 163.367
R554 B.n526 B.n525 163.367
R555 B.n525 B.n524 163.367
R556 B.n524 B.n99 163.367
R557 B.n520 B.n99 163.367
R558 B.n520 B.n519 163.367
R559 B.n519 B.n518 163.367
R560 B.n518 B.n101 163.367
R561 B.n514 B.n101 163.367
R562 B.n514 B.n513 163.367
R563 B.n513 B.n512 163.367
R564 B.n512 B.n103 163.367
R565 B.n508 B.n103 163.367
R566 B.n508 B.n507 163.367
R567 B.n507 B.n506 163.367
R568 B.n506 B.n105 163.367
R569 B.n502 B.n105 163.367
R570 B.n502 B.n501 163.367
R571 B.n501 B.n500 163.367
R572 B.n500 B.n107 163.367
R573 B.n496 B.n107 163.367
R574 B.n496 B.n495 163.367
R575 B.n495 B.n494 163.367
R576 B.n494 B.n109 163.367
R577 B.n490 B.n109 163.367
R578 B.n490 B.n489 163.367
R579 B.n489 B.n488 163.367
R580 B.n488 B.n111 163.367
R581 B.n484 B.n111 163.367
R582 B.n484 B.n483 163.367
R583 B.n483 B.n482 163.367
R584 B.n482 B.n113 163.367
R585 B.n478 B.n113 163.367
R586 B.n478 B.n477 163.367
R587 B.n477 B.n476 163.367
R588 B.n476 B.n115 163.367
R589 B.n472 B.n115 163.367
R590 B.n472 B.n471 163.367
R591 B.n471 B.n470 163.367
R592 B.n470 B.n117 163.367
R593 B.n466 B.n117 163.367
R594 B.n466 B.n465 163.367
R595 B.n465 B.n464 163.367
R596 B.n464 B.n119 163.367
R597 B.n460 B.n119 163.367
R598 B.n460 B.n459 163.367
R599 B.n459 B.n458 163.367
R600 B.n458 B.n121 163.367
R601 B.n454 B.n121 163.367
R602 B.n454 B.n453 163.367
R603 B.n453 B.n452 163.367
R604 B.n452 B.n123 163.367
R605 B.n448 B.n123 163.367
R606 B.n448 B.n447 163.367
R607 B.n447 B.n446 163.367
R608 B.n744 B.n743 163.367
R609 B.n743 B.n742 163.367
R610 B.n742 B.n23 163.367
R611 B.n738 B.n23 163.367
R612 B.n738 B.n737 163.367
R613 B.n737 B.n736 163.367
R614 B.n736 B.n25 163.367
R615 B.n732 B.n25 163.367
R616 B.n732 B.n731 163.367
R617 B.n731 B.n730 163.367
R618 B.n730 B.n27 163.367
R619 B.n726 B.n27 163.367
R620 B.n726 B.n725 163.367
R621 B.n725 B.n724 163.367
R622 B.n724 B.n29 163.367
R623 B.n720 B.n29 163.367
R624 B.n720 B.n719 163.367
R625 B.n719 B.n718 163.367
R626 B.n718 B.n31 163.367
R627 B.n714 B.n31 163.367
R628 B.n714 B.n713 163.367
R629 B.n713 B.n712 163.367
R630 B.n712 B.n33 163.367
R631 B.n708 B.n33 163.367
R632 B.n708 B.n707 163.367
R633 B.n707 B.n706 163.367
R634 B.n706 B.n35 163.367
R635 B.n702 B.n35 163.367
R636 B.n702 B.n701 163.367
R637 B.n701 B.n700 163.367
R638 B.n700 B.n37 163.367
R639 B.n696 B.n37 163.367
R640 B.n696 B.n695 163.367
R641 B.n695 B.n694 163.367
R642 B.n694 B.n39 163.367
R643 B.n690 B.n39 163.367
R644 B.n690 B.n689 163.367
R645 B.n689 B.n688 163.367
R646 B.n688 B.n41 163.367
R647 B.n684 B.n41 163.367
R648 B.n684 B.n683 163.367
R649 B.n683 B.n682 163.367
R650 B.n682 B.n43 163.367
R651 B.n678 B.n43 163.367
R652 B.n678 B.n677 163.367
R653 B.n677 B.n676 163.367
R654 B.n676 B.n45 163.367
R655 B.n672 B.n45 163.367
R656 B.n672 B.n671 163.367
R657 B.n671 B.n670 163.367
R658 B.n670 B.n47 163.367
R659 B.n666 B.n47 163.367
R660 B.n666 B.n665 163.367
R661 B.n665 B.n664 163.367
R662 B.n664 B.n49 163.367
R663 B.n659 B.n49 163.367
R664 B.n659 B.n658 163.367
R665 B.n658 B.n657 163.367
R666 B.n657 B.n53 163.367
R667 B.n653 B.n53 163.367
R668 B.n653 B.n652 163.367
R669 B.n652 B.n651 163.367
R670 B.n651 B.n55 163.367
R671 B.n646 B.n55 163.367
R672 B.n646 B.n645 163.367
R673 B.n645 B.n644 163.367
R674 B.n644 B.n59 163.367
R675 B.n640 B.n59 163.367
R676 B.n640 B.n639 163.367
R677 B.n639 B.n638 163.367
R678 B.n638 B.n61 163.367
R679 B.n634 B.n61 163.367
R680 B.n634 B.n633 163.367
R681 B.n633 B.n632 163.367
R682 B.n632 B.n63 163.367
R683 B.n628 B.n63 163.367
R684 B.n628 B.n627 163.367
R685 B.n627 B.n626 163.367
R686 B.n626 B.n65 163.367
R687 B.n622 B.n65 163.367
R688 B.n622 B.n621 163.367
R689 B.n621 B.n620 163.367
R690 B.n620 B.n67 163.367
R691 B.n616 B.n67 163.367
R692 B.n616 B.n615 163.367
R693 B.n615 B.n614 163.367
R694 B.n614 B.n69 163.367
R695 B.n610 B.n69 163.367
R696 B.n610 B.n609 163.367
R697 B.n609 B.n608 163.367
R698 B.n608 B.n71 163.367
R699 B.n604 B.n71 163.367
R700 B.n604 B.n603 163.367
R701 B.n603 B.n602 163.367
R702 B.n602 B.n73 163.367
R703 B.n598 B.n73 163.367
R704 B.n598 B.n597 163.367
R705 B.n597 B.n596 163.367
R706 B.n596 B.n75 163.367
R707 B.n592 B.n75 163.367
R708 B.n592 B.n591 163.367
R709 B.n591 B.n590 163.367
R710 B.n590 B.n77 163.367
R711 B.n586 B.n77 163.367
R712 B.n586 B.n585 163.367
R713 B.n585 B.n584 163.367
R714 B.n584 B.n79 163.367
R715 B.n580 B.n79 163.367
R716 B.n580 B.n579 163.367
R717 B.n579 B.n578 163.367
R718 B.n578 B.n81 163.367
R719 B.n574 B.n81 163.367
R720 B.n574 B.n573 163.367
R721 B.n573 B.n572 163.367
R722 B.n572 B.n83 163.367
R723 B.n568 B.n83 163.367
R724 B.n568 B.n567 163.367
R725 B.n567 B.n566 163.367
R726 B.n748 B.n21 163.367
R727 B.n749 B.n748 163.367
R728 B.n750 B.n749 163.367
R729 B.n750 B.n19 163.367
R730 B.n754 B.n19 163.367
R731 B.n755 B.n754 163.367
R732 B.n756 B.n755 163.367
R733 B.n756 B.n17 163.367
R734 B.n760 B.n17 163.367
R735 B.n761 B.n760 163.367
R736 B.n762 B.n761 163.367
R737 B.n762 B.n15 163.367
R738 B.n766 B.n15 163.367
R739 B.n767 B.n766 163.367
R740 B.n768 B.n767 163.367
R741 B.n768 B.n13 163.367
R742 B.n772 B.n13 163.367
R743 B.n773 B.n772 163.367
R744 B.n774 B.n773 163.367
R745 B.n774 B.n11 163.367
R746 B.n778 B.n11 163.367
R747 B.n779 B.n778 163.367
R748 B.n780 B.n779 163.367
R749 B.n780 B.n9 163.367
R750 B.n784 B.n9 163.367
R751 B.n785 B.n784 163.367
R752 B.n786 B.n785 163.367
R753 B.n786 B.n7 163.367
R754 B.n790 B.n7 163.367
R755 B.n791 B.n790 163.367
R756 B.n792 B.n791 163.367
R757 B.n792 B.n5 163.367
R758 B.n796 B.n5 163.367
R759 B.n797 B.n796 163.367
R760 B.n798 B.n797 163.367
R761 B.n798 B.n3 163.367
R762 B.n802 B.n3 163.367
R763 B.n803 B.n802 163.367
R764 B.n205 B.n2 163.367
R765 B.n208 B.n205 163.367
R766 B.n209 B.n208 163.367
R767 B.n210 B.n209 163.367
R768 B.n210 B.n203 163.367
R769 B.n214 B.n203 163.367
R770 B.n215 B.n214 163.367
R771 B.n216 B.n215 163.367
R772 B.n216 B.n201 163.367
R773 B.n220 B.n201 163.367
R774 B.n221 B.n220 163.367
R775 B.n222 B.n221 163.367
R776 B.n222 B.n199 163.367
R777 B.n226 B.n199 163.367
R778 B.n227 B.n226 163.367
R779 B.n228 B.n227 163.367
R780 B.n228 B.n197 163.367
R781 B.n232 B.n197 163.367
R782 B.n233 B.n232 163.367
R783 B.n234 B.n233 163.367
R784 B.n234 B.n195 163.367
R785 B.n238 B.n195 163.367
R786 B.n239 B.n238 163.367
R787 B.n240 B.n239 163.367
R788 B.n240 B.n193 163.367
R789 B.n244 B.n193 163.367
R790 B.n245 B.n244 163.367
R791 B.n246 B.n245 163.367
R792 B.n246 B.n191 163.367
R793 B.n250 B.n191 163.367
R794 B.n251 B.n250 163.367
R795 B.n252 B.n251 163.367
R796 B.n252 B.n189 163.367
R797 B.n256 B.n189 163.367
R798 B.n257 B.n256 163.367
R799 B.n258 B.n257 163.367
R800 B.n258 B.n187 163.367
R801 B.n262 B.n187 163.367
R802 B.n359 B.t5 108.701
R803 B.n57 B.t1 108.701
R804 B.n159 B.t11 108.68
R805 B.n51 B.t7 108.68
R806 B.n159 B.n158 69.4308
R807 B.n359 B.n358 69.4308
R808 B.n57 B.n56 69.4308
R809 B.n51 B.n50 69.4308
R810 B.n345 B.n159 59.5399
R811 B.n360 B.n359 59.5399
R812 B.n648 B.n57 59.5399
R813 B.n662 B.n51 59.5399
R814 B.n746 B.n745 34.1859
R815 B.n565 B.n564 34.1859
R816 B.n445 B.n444 34.1859
R817 B.n261 B.n186 34.1859
R818 B B.n805 18.0485
R819 B.n747 B.n746 10.6151
R820 B.n747 B.n20 10.6151
R821 B.n751 B.n20 10.6151
R822 B.n752 B.n751 10.6151
R823 B.n753 B.n752 10.6151
R824 B.n753 B.n18 10.6151
R825 B.n757 B.n18 10.6151
R826 B.n758 B.n757 10.6151
R827 B.n759 B.n758 10.6151
R828 B.n759 B.n16 10.6151
R829 B.n763 B.n16 10.6151
R830 B.n764 B.n763 10.6151
R831 B.n765 B.n764 10.6151
R832 B.n765 B.n14 10.6151
R833 B.n769 B.n14 10.6151
R834 B.n770 B.n769 10.6151
R835 B.n771 B.n770 10.6151
R836 B.n771 B.n12 10.6151
R837 B.n775 B.n12 10.6151
R838 B.n776 B.n775 10.6151
R839 B.n777 B.n776 10.6151
R840 B.n777 B.n10 10.6151
R841 B.n781 B.n10 10.6151
R842 B.n782 B.n781 10.6151
R843 B.n783 B.n782 10.6151
R844 B.n783 B.n8 10.6151
R845 B.n787 B.n8 10.6151
R846 B.n788 B.n787 10.6151
R847 B.n789 B.n788 10.6151
R848 B.n789 B.n6 10.6151
R849 B.n793 B.n6 10.6151
R850 B.n794 B.n793 10.6151
R851 B.n795 B.n794 10.6151
R852 B.n795 B.n4 10.6151
R853 B.n799 B.n4 10.6151
R854 B.n800 B.n799 10.6151
R855 B.n801 B.n800 10.6151
R856 B.n801 B.n0 10.6151
R857 B.n745 B.n22 10.6151
R858 B.n741 B.n22 10.6151
R859 B.n741 B.n740 10.6151
R860 B.n740 B.n739 10.6151
R861 B.n739 B.n24 10.6151
R862 B.n735 B.n24 10.6151
R863 B.n735 B.n734 10.6151
R864 B.n734 B.n733 10.6151
R865 B.n733 B.n26 10.6151
R866 B.n729 B.n26 10.6151
R867 B.n729 B.n728 10.6151
R868 B.n728 B.n727 10.6151
R869 B.n727 B.n28 10.6151
R870 B.n723 B.n28 10.6151
R871 B.n723 B.n722 10.6151
R872 B.n722 B.n721 10.6151
R873 B.n721 B.n30 10.6151
R874 B.n717 B.n30 10.6151
R875 B.n717 B.n716 10.6151
R876 B.n716 B.n715 10.6151
R877 B.n715 B.n32 10.6151
R878 B.n711 B.n32 10.6151
R879 B.n711 B.n710 10.6151
R880 B.n710 B.n709 10.6151
R881 B.n709 B.n34 10.6151
R882 B.n705 B.n34 10.6151
R883 B.n705 B.n704 10.6151
R884 B.n704 B.n703 10.6151
R885 B.n703 B.n36 10.6151
R886 B.n699 B.n36 10.6151
R887 B.n699 B.n698 10.6151
R888 B.n698 B.n697 10.6151
R889 B.n697 B.n38 10.6151
R890 B.n693 B.n38 10.6151
R891 B.n693 B.n692 10.6151
R892 B.n692 B.n691 10.6151
R893 B.n691 B.n40 10.6151
R894 B.n687 B.n40 10.6151
R895 B.n687 B.n686 10.6151
R896 B.n686 B.n685 10.6151
R897 B.n685 B.n42 10.6151
R898 B.n681 B.n42 10.6151
R899 B.n681 B.n680 10.6151
R900 B.n680 B.n679 10.6151
R901 B.n679 B.n44 10.6151
R902 B.n675 B.n44 10.6151
R903 B.n675 B.n674 10.6151
R904 B.n674 B.n673 10.6151
R905 B.n673 B.n46 10.6151
R906 B.n669 B.n46 10.6151
R907 B.n669 B.n668 10.6151
R908 B.n668 B.n667 10.6151
R909 B.n667 B.n48 10.6151
R910 B.n663 B.n48 10.6151
R911 B.n661 B.n660 10.6151
R912 B.n660 B.n52 10.6151
R913 B.n656 B.n52 10.6151
R914 B.n656 B.n655 10.6151
R915 B.n655 B.n654 10.6151
R916 B.n654 B.n54 10.6151
R917 B.n650 B.n54 10.6151
R918 B.n650 B.n649 10.6151
R919 B.n647 B.n58 10.6151
R920 B.n643 B.n58 10.6151
R921 B.n643 B.n642 10.6151
R922 B.n642 B.n641 10.6151
R923 B.n641 B.n60 10.6151
R924 B.n637 B.n60 10.6151
R925 B.n637 B.n636 10.6151
R926 B.n636 B.n635 10.6151
R927 B.n635 B.n62 10.6151
R928 B.n631 B.n62 10.6151
R929 B.n631 B.n630 10.6151
R930 B.n630 B.n629 10.6151
R931 B.n629 B.n64 10.6151
R932 B.n625 B.n64 10.6151
R933 B.n625 B.n624 10.6151
R934 B.n624 B.n623 10.6151
R935 B.n623 B.n66 10.6151
R936 B.n619 B.n66 10.6151
R937 B.n619 B.n618 10.6151
R938 B.n618 B.n617 10.6151
R939 B.n617 B.n68 10.6151
R940 B.n613 B.n68 10.6151
R941 B.n613 B.n612 10.6151
R942 B.n612 B.n611 10.6151
R943 B.n611 B.n70 10.6151
R944 B.n607 B.n70 10.6151
R945 B.n607 B.n606 10.6151
R946 B.n606 B.n605 10.6151
R947 B.n605 B.n72 10.6151
R948 B.n601 B.n72 10.6151
R949 B.n601 B.n600 10.6151
R950 B.n600 B.n599 10.6151
R951 B.n599 B.n74 10.6151
R952 B.n595 B.n74 10.6151
R953 B.n595 B.n594 10.6151
R954 B.n594 B.n593 10.6151
R955 B.n593 B.n76 10.6151
R956 B.n589 B.n76 10.6151
R957 B.n589 B.n588 10.6151
R958 B.n588 B.n587 10.6151
R959 B.n587 B.n78 10.6151
R960 B.n583 B.n78 10.6151
R961 B.n583 B.n582 10.6151
R962 B.n582 B.n581 10.6151
R963 B.n581 B.n80 10.6151
R964 B.n577 B.n80 10.6151
R965 B.n577 B.n576 10.6151
R966 B.n576 B.n575 10.6151
R967 B.n575 B.n82 10.6151
R968 B.n571 B.n82 10.6151
R969 B.n571 B.n570 10.6151
R970 B.n570 B.n569 10.6151
R971 B.n569 B.n84 10.6151
R972 B.n565 B.n84 10.6151
R973 B.n564 B.n563 10.6151
R974 B.n563 B.n86 10.6151
R975 B.n559 B.n86 10.6151
R976 B.n559 B.n558 10.6151
R977 B.n558 B.n557 10.6151
R978 B.n557 B.n88 10.6151
R979 B.n553 B.n88 10.6151
R980 B.n553 B.n552 10.6151
R981 B.n552 B.n551 10.6151
R982 B.n551 B.n90 10.6151
R983 B.n547 B.n90 10.6151
R984 B.n547 B.n546 10.6151
R985 B.n546 B.n545 10.6151
R986 B.n545 B.n92 10.6151
R987 B.n541 B.n92 10.6151
R988 B.n541 B.n540 10.6151
R989 B.n540 B.n539 10.6151
R990 B.n539 B.n94 10.6151
R991 B.n535 B.n94 10.6151
R992 B.n535 B.n534 10.6151
R993 B.n534 B.n533 10.6151
R994 B.n533 B.n96 10.6151
R995 B.n529 B.n96 10.6151
R996 B.n529 B.n528 10.6151
R997 B.n528 B.n527 10.6151
R998 B.n527 B.n98 10.6151
R999 B.n523 B.n98 10.6151
R1000 B.n523 B.n522 10.6151
R1001 B.n522 B.n521 10.6151
R1002 B.n521 B.n100 10.6151
R1003 B.n517 B.n100 10.6151
R1004 B.n517 B.n516 10.6151
R1005 B.n516 B.n515 10.6151
R1006 B.n515 B.n102 10.6151
R1007 B.n511 B.n102 10.6151
R1008 B.n511 B.n510 10.6151
R1009 B.n510 B.n509 10.6151
R1010 B.n509 B.n104 10.6151
R1011 B.n505 B.n104 10.6151
R1012 B.n505 B.n504 10.6151
R1013 B.n504 B.n503 10.6151
R1014 B.n503 B.n106 10.6151
R1015 B.n499 B.n106 10.6151
R1016 B.n499 B.n498 10.6151
R1017 B.n498 B.n497 10.6151
R1018 B.n497 B.n108 10.6151
R1019 B.n493 B.n108 10.6151
R1020 B.n493 B.n492 10.6151
R1021 B.n492 B.n491 10.6151
R1022 B.n491 B.n110 10.6151
R1023 B.n487 B.n110 10.6151
R1024 B.n487 B.n486 10.6151
R1025 B.n486 B.n485 10.6151
R1026 B.n485 B.n112 10.6151
R1027 B.n481 B.n112 10.6151
R1028 B.n481 B.n480 10.6151
R1029 B.n480 B.n479 10.6151
R1030 B.n479 B.n114 10.6151
R1031 B.n475 B.n114 10.6151
R1032 B.n475 B.n474 10.6151
R1033 B.n474 B.n473 10.6151
R1034 B.n473 B.n116 10.6151
R1035 B.n469 B.n116 10.6151
R1036 B.n469 B.n468 10.6151
R1037 B.n468 B.n467 10.6151
R1038 B.n467 B.n118 10.6151
R1039 B.n463 B.n118 10.6151
R1040 B.n463 B.n462 10.6151
R1041 B.n462 B.n461 10.6151
R1042 B.n461 B.n120 10.6151
R1043 B.n457 B.n120 10.6151
R1044 B.n457 B.n456 10.6151
R1045 B.n456 B.n455 10.6151
R1046 B.n455 B.n122 10.6151
R1047 B.n451 B.n122 10.6151
R1048 B.n451 B.n450 10.6151
R1049 B.n450 B.n449 10.6151
R1050 B.n449 B.n124 10.6151
R1051 B.n445 B.n124 10.6151
R1052 B.n206 B.n1 10.6151
R1053 B.n207 B.n206 10.6151
R1054 B.n207 B.n204 10.6151
R1055 B.n211 B.n204 10.6151
R1056 B.n212 B.n211 10.6151
R1057 B.n213 B.n212 10.6151
R1058 B.n213 B.n202 10.6151
R1059 B.n217 B.n202 10.6151
R1060 B.n218 B.n217 10.6151
R1061 B.n219 B.n218 10.6151
R1062 B.n219 B.n200 10.6151
R1063 B.n223 B.n200 10.6151
R1064 B.n224 B.n223 10.6151
R1065 B.n225 B.n224 10.6151
R1066 B.n225 B.n198 10.6151
R1067 B.n229 B.n198 10.6151
R1068 B.n230 B.n229 10.6151
R1069 B.n231 B.n230 10.6151
R1070 B.n231 B.n196 10.6151
R1071 B.n235 B.n196 10.6151
R1072 B.n236 B.n235 10.6151
R1073 B.n237 B.n236 10.6151
R1074 B.n237 B.n194 10.6151
R1075 B.n241 B.n194 10.6151
R1076 B.n242 B.n241 10.6151
R1077 B.n243 B.n242 10.6151
R1078 B.n243 B.n192 10.6151
R1079 B.n247 B.n192 10.6151
R1080 B.n248 B.n247 10.6151
R1081 B.n249 B.n248 10.6151
R1082 B.n249 B.n190 10.6151
R1083 B.n253 B.n190 10.6151
R1084 B.n254 B.n253 10.6151
R1085 B.n255 B.n254 10.6151
R1086 B.n255 B.n188 10.6151
R1087 B.n259 B.n188 10.6151
R1088 B.n260 B.n259 10.6151
R1089 B.n261 B.n260 10.6151
R1090 B.n265 B.n186 10.6151
R1091 B.n266 B.n265 10.6151
R1092 B.n267 B.n266 10.6151
R1093 B.n267 B.n184 10.6151
R1094 B.n271 B.n184 10.6151
R1095 B.n272 B.n271 10.6151
R1096 B.n273 B.n272 10.6151
R1097 B.n273 B.n182 10.6151
R1098 B.n277 B.n182 10.6151
R1099 B.n278 B.n277 10.6151
R1100 B.n279 B.n278 10.6151
R1101 B.n279 B.n180 10.6151
R1102 B.n283 B.n180 10.6151
R1103 B.n284 B.n283 10.6151
R1104 B.n285 B.n284 10.6151
R1105 B.n285 B.n178 10.6151
R1106 B.n289 B.n178 10.6151
R1107 B.n290 B.n289 10.6151
R1108 B.n291 B.n290 10.6151
R1109 B.n291 B.n176 10.6151
R1110 B.n295 B.n176 10.6151
R1111 B.n296 B.n295 10.6151
R1112 B.n297 B.n296 10.6151
R1113 B.n297 B.n174 10.6151
R1114 B.n301 B.n174 10.6151
R1115 B.n302 B.n301 10.6151
R1116 B.n303 B.n302 10.6151
R1117 B.n303 B.n172 10.6151
R1118 B.n307 B.n172 10.6151
R1119 B.n308 B.n307 10.6151
R1120 B.n309 B.n308 10.6151
R1121 B.n309 B.n170 10.6151
R1122 B.n313 B.n170 10.6151
R1123 B.n314 B.n313 10.6151
R1124 B.n315 B.n314 10.6151
R1125 B.n315 B.n168 10.6151
R1126 B.n319 B.n168 10.6151
R1127 B.n320 B.n319 10.6151
R1128 B.n321 B.n320 10.6151
R1129 B.n321 B.n166 10.6151
R1130 B.n325 B.n166 10.6151
R1131 B.n326 B.n325 10.6151
R1132 B.n327 B.n326 10.6151
R1133 B.n327 B.n164 10.6151
R1134 B.n331 B.n164 10.6151
R1135 B.n332 B.n331 10.6151
R1136 B.n333 B.n332 10.6151
R1137 B.n333 B.n162 10.6151
R1138 B.n337 B.n162 10.6151
R1139 B.n338 B.n337 10.6151
R1140 B.n339 B.n338 10.6151
R1141 B.n339 B.n160 10.6151
R1142 B.n343 B.n160 10.6151
R1143 B.n344 B.n343 10.6151
R1144 B.n346 B.n156 10.6151
R1145 B.n350 B.n156 10.6151
R1146 B.n351 B.n350 10.6151
R1147 B.n352 B.n351 10.6151
R1148 B.n352 B.n154 10.6151
R1149 B.n356 B.n154 10.6151
R1150 B.n357 B.n356 10.6151
R1151 B.n361 B.n357 10.6151
R1152 B.n365 B.n152 10.6151
R1153 B.n366 B.n365 10.6151
R1154 B.n367 B.n366 10.6151
R1155 B.n367 B.n150 10.6151
R1156 B.n371 B.n150 10.6151
R1157 B.n372 B.n371 10.6151
R1158 B.n373 B.n372 10.6151
R1159 B.n373 B.n148 10.6151
R1160 B.n377 B.n148 10.6151
R1161 B.n378 B.n377 10.6151
R1162 B.n379 B.n378 10.6151
R1163 B.n379 B.n146 10.6151
R1164 B.n383 B.n146 10.6151
R1165 B.n384 B.n383 10.6151
R1166 B.n385 B.n384 10.6151
R1167 B.n385 B.n144 10.6151
R1168 B.n389 B.n144 10.6151
R1169 B.n390 B.n389 10.6151
R1170 B.n391 B.n390 10.6151
R1171 B.n391 B.n142 10.6151
R1172 B.n395 B.n142 10.6151
R1173 B.n396 B.n395 10.6151
R1174 B.n397 B.n396 10.6151
R1175 B.n397 B.n140 10.6151
R1176 B.n401 B.n140 10.6151
R1177 B.n402 B.n401 10.6151
R1178 B.n403 B.n402 10.6151
R1179 B.n403 B.n138 10.6151
R1180 B.n407 B.n138 10.6151
R1181 B.n408 B.n407 10.6151
R1182 B.n409 B.n408 10.6151
R1183 B.n409 B.n136 10.6151
R1184 B.n413 B.n136 10.6151
R1185 B.n414 B.n413 10.6151
R1186 B.n415 B.n414 10.6151
R1187 B.n415 B.n134 10.6151
R1188 B.n419 B.n134 10.6151
R1189 B.n420 B.n419 10.6151
R1190 B.n421 B.n420 10.6151
R1191 B.n421 B.n132 10.6151
R1192 B.n425 B.n132 10.6151
R1193 B.n426 B.n425 10.6151
R1194 B.n427 B.n426 10.6151
R1195 B.n427 B.n130 10.6151
R1196 B.n431 B.n130 10.6151
R1197 B.n432 B.n431 10.6151
R1198 B.n433 B.n432 10.6151
R1199 B.n433 B.n128 10.6151
R1200 B.n437 B.n128 10.6151
R1201 B.n438 B.n437 10.6151
R1202 B.n439 B.n438 10.6151
R1203 B.n439 B.n126 10.6151
R1204 B.n443 B.n126 10.6151
R1205 B.n444 B.n443 10.6151
R1206 B.n805 B.n0 8.11757
R1207 B.n805 B.n1 8.11757
R1208 B.n662 B.n661 6.5566
R1209 B.n649 B.n648 6.5566
R1210 B.n346 B.n345 6.5566
R1211 B.n361 B.n360 6.5566
R1212 B.n663 B.n662 4.05904
R1213 B.n648 B.n647 4.05904
R1214 B.n345 B.n344 4.05904
R1215 B.n360 B.n152 4.05904
R1216 VN.n1 VN.t2 156.633
R1217 VN.n0 VN.t0 156.633
R1218 VN.n0 VN.t3 155.528
R1219 VN.n1 VN.t1 155.528
R1220 VN VN.n1 54.4298
R1221 VN VN.n0 2.56238
R1222 VDD2.n2 VDD2.n0 116.737
R1223 VDD2.n2 VDD2.n1 69.5913
R1224 VDD2.n1 VDD2.t3 1.97769
R1225 VDD2.n1 VDD2.t1 1.97769
R1226 VDD2.n0 VDD2.t0 1.97769
R1227 VDD2.n0 VDD2.t2 1.97769
R1228 VDD2 VDD2.n2 0.0586897
R1229 VTAIL.n5 VTAIL.t3 54.8899
R1230 VTAIL.n4 VTAIL.t5 54.8899
R1231 VTAIL.n3 VTAIL.t6 54.8899
R1232 VTAIL.n7 VTAIL.t4 54.8896
R1233 VTAIL.n0 VTAIL.t7 54.8896
R1234 VTAIL.n1 VTAIL.t0 54.8896
R1235 VTAIL.n2 VTAIL.t2 54.8896
R1236 VTAIL.n6 VTAIL.t1 54.8896
R1237 VTAIL.n7 VTAIL.n6 29.6255
R1238 VTAIL.n3 VTAIL.n2 29.6255
R1239 VTAIL.n4 VTAIL.n3 3.08671
R1240 VTAIL.n6 VTAIL.n5 3.08671
R1241 VTAIL.n2 VTAIL.n1 3.08671
R1242 VTAIL VTAIL.n0 1.60179
R1243 VTAIL VTAIL.n7 1.48541
R1244 VTAIL.n5 VTAIL.n4 0.470328
R1245 VTAIL.n1 VTAIL.n0 0.470328
R1246 VP.n17 VP.n16 161.3
R1247 VP.n15 VP.n1 161.3
R1248 VP.n14 VP.n13 161.3
R1249 VP.n12 VP.n2 161.3
R1250 VP.n11 VP.n10 161.3
R1251 VP.n9 VP.n3 161.3
R1252 VP.n8 VP.n7 161.3
R1253 VP.n5 VP.t1 156.633
R1254 VP.n5 VP.t0 155.528
R1255 VP.n4 VP.t3 121.909
R1256 VP.n0 VP.t2 121.909
R1257 VP.n6 VP.n4 75.7718
R1258 VP.n18 VP.n0 75.7718
R1259 VP.n6 VP.n5 54.2643
R1260 VP.n10 VP.n2 40.4106
R1261 VP.n14 VP.n2 40.4106
R1262 VP.n9 VP.n8 24.3439
R1263 VP.n10 VP.n9 24.3439
R1264 VP.n15 VP.n14 24.3439
R1265 VP.n16 VP.n15 24.3439
R1266 VP.n8 VP.n4 14.1197
R1267 VP.n16 VP.n0 14.1197
R1268 VP.n7 VP.n6 0.355081
R1269 VP.n18 VP.n17 0.355081
R1270 VP VP.n18 0.26685
R1271 VP.n7 VP.n3 0.189894
R1272 VP.n11 VP.n3 0.189894
R1273 VP.n12 VP.n11 0.189894
R1274 VP.n13 VP.n12 0.189894
R1275 VP.n13 VP.n1 0.189894
R1276 VP.n17 VP.n1 0.189894
R1277 VDD1 VDD1.n1 117.261
R1278 VDD1 VDD1.n0 69.6495
R1279 VDD1.n0 VDD1.t2 1.97769
R1280 VDD1.n0 VDD1.t3 1.97769
R1281 VDD1.n1 VDD1.t0 1.97769
R1282 VDD1.n1 VDD1.t1 1.97769
C0 VDD2 VDD1 1.18571f
C1 VTAIL VDD1 6.53302f
C2 VN VP 7.48816f
C3 VDD1 w_n3118_n4256# 1.69245f
C4 VP B 1.95087f
C5 VP VDD2 0.435177f
C6 VTAIL VP 6.44554f
C7 VN B 1.27995f
C8 VP w_n3118_n4256# 5.89879f
C9 VN VDD2 6.63369f
C10 B VDD2 1.55905f
C11 VTAIL VN 6.43144f
C12 VTAIL B 6.7263f
C13 VN w_n3118_n4256# 5.49631f
C14 B w_n3118_n4256# 11.2895f
C15 VTAIL VDD2 6.59158f
C16 VDD2 w_n3118_n4256# 1.76295f
C17 VTAIL w_n3118_n4256# 4.97332f
C18 VP VDD1 6.91886f
C19 VN VDD1 0.149098f
C20 B VDD1 1.49612f
C21 VDD2 VSUBS 1.150583f
C22 VDD1 VSUBS 6.6263f
C23 VTAIL VSUBS 1.496716f
C24 VN VSUBS 5.94108f
C25 VP VSUBS 2.792252f
C26 B VSUBS 5.210573f
C27 w_n3118_n4256# VSUBS 0.162498p
C28 VDD1.t2 VSUBS 0.349083f
C29 VDD1.t3 VSUBS 0.349083f
C30 VDD1.n0 VSUBS 2.86721f
C31 VDD1.t0 VSUBS 0.349083f
C32 VDD1.t1 VSUBS 0.349083f
C33 VDD1.n1 VSUBS 3.83242f
C34 VP.t2 VSUBS 4.01802f
C35 VP.n0 VSUBS 1.49855f
C36 VP.n1 VSUBS 0.027389f
C37 VP.n2 VSUBS 0.022164f
C38 VP.n3 VSUBS 0.027389f
C39 VP.t3 VSUBS 4.01802f
C40 VP.n4 VSUBS 1.49855f
C41 VP.t1 VSUBS 4.37221f
C42 VP.t0 VSUBS 4.36129f
C43 VP.n5 VSUBS 4.52485f
C44 VP.n6 VSUBS 1.74689f
C45 VP.n7 VSUBS 0.044213f
C46 VP.n8 VSUBS 0.040664f
C47 VP.n9 VSUBS 0.051303f
C48 VP.n10 VSUBS 0.054727f
C49 VP.n11 VSUBS 0.027389f
C50 VP.n12 VSUBS 0.027389f
C51 VP.n13 VSUBS 0.027389f
C52 VP.n14 VSUBS 0.054727f
C53 VP.n15 VSUBS 0.051303f
C54 VP.n16 VSUBS 0.040664f
C55 VP.n17 VSUBS 0.044213f
C56 VP.n18 VSUBS 0.066303f
C57 VTAIL.t7 VSUBS 3.00937f
C58 VTAIL.n0 VSUBS 0.807355f
C59 VTAIL.t0 VSUBS 3.00937f
C60 VTAIL.n1 VSUBS 0.916771f
C61 VTAIL.t2 VSUBS 3.00937f
C62 VTAIL.n2 VSUBS 2.46448f
C63 VTAIL.t6 VSUBS 3.00938f
C64 VTAIL.n3 VSUBS 2.46447f
C65 VTAIL.t5 VSUBS 3.00938f
C66 VTAIL.n4 VSUBS 0.916766f
C67 VTAIL.t3 VSUBS 3.00938f
C68 VTAIL.n5 VSUBS 0.916766f
C69 VTAIL.t1 VSUBS 3.00937f
C70 VTAIL.n6 VSUBS 2.46448f
C71 VTAIL.t4 VSUBS 3.00937f
C72 VTAIL.n7 VSUBS 2.34649f
C73 VDD2.t0 VSUBS 0.346439f
C74 VDD2.t2 VSUBS 0.346439f
C75 VDD2.n0 VSUBS 3.77598f
C76 VDD2.t3 VSUBS 0.346439f
C77 VDD2.t1 VSUBS 0.346439f
C78 VDD2.n1 VSUBS 2.84482f
C79 VDD2.n2 VSUBS 4.92252f
C80 VN.t3 VSUBS 4.24084f
C81 VN.t0 VSUBS 4.25145f
C82 VN.n0 VSUBS 2.62691f
C83 VN.t1 VSUBS 4.24084f
C84 VN.t2 VSUBS 4.25145f
C85 VN.n1 VSUBS 4.41042f
C86 B.n0 VSUBS 0.005139f
C87 B.n1 VSUBS 0.005139f
C88 B.n2 VSUBS 0.0076f
C89 B.n3 VSUBS 0.005824f
C90 B.n4 VSUBS 0.005824f
C91 B.n5 VSUBS 0.005824f
C92 B.n6 VSUBS 0.005824f
C93 B.n7 VSUBS 0.005824f
C94 B.n8 VSUBS 0.005824f
C95 B.n9 VSUBS 0.005824f
C96 B.n10 VSUBS 0.005824f
C97 B.n11 VSUBS 0.005824f
C98 B.n12 VSUBS 0.005824f
C99 B.n13 VSUBS 0.005824f
C100 B.n14 VSUBS 0.005824f
C101 B.n15 VSUBS 0.005824f
C102 B.n16 VSUBS 0.005824f
C103 B.n17 VSUBS 0.005824f
C104 B.n18 VSUBS 0.005824f
C105 B.n19 VSUBS 0.005824f
C106 B.n20 VSUBS 0.005824f
C107 B.n21 VSUBS 0.013605f
C108 B.n22 VSUBS 0.005824f
C109 B.n23 VSUBS 0.005824f
C110 B.n24 VSUBS 0.005824f
C111 B.n25 VSUBS 0.005824f
C112 B.n26 VSUBS 0.005824f
C113 B.n27 VSUBS 0.005824f
C114 B.n28 VSUBS 0.005824f
C115 B.n29 VSUBS 0.005824f
C116 B.n30 VSUBS 0.005824f
C117 B.n31 VSUBS 0.005824f
C118 B.n32 VSUBS 0.005824f
C119 B.n33 VSUBS 0.005824f
C120 B.n34 VSUBS 0.005824f
C121 B.n35 VSUBS 0.005824f
C122 B.n36 VSUBS 0.005824f
C123 B.n37 VSUBS 0.005824f
C124 B.n38 VSUBS 0.005824f
C125 B.n39 VSUBS 0.005824f
C126 B.n40 VSUBS 0.005824f
C127 B.n41 VSUBS 0.005824f
C128 B.n42 VSUBS 0.005824f
C129 B.n43 VSUBS 0.005824f
C130 B.n44 VSUBS 0.005824f
C131 B.n45 VSUBS 0.005824f
C132 B.n46 VSUBS 0.005824f
C133 B.n47 VSUBS 0.005824f
C134 B.n48 VSUBS 0.005824f
C135 B.n49 VSUBS 0.005824f
C136 B.t7 VSUBS 0.458706f
C137 B.t8 VSUBS 0.47971f
C138 B.t6 VSUBS 2.01572f
C139 B.n50 VSUBS 0.278622f
C140 B.n51 VSUBS 0.062188f
C141 B.n52 VSUBS 0.005824f
C142 B.n53 VSUBS 0.005824f
C143 B.n54 VSUBS 0.005824f
C144 B.n55 VSUBS 0.005824f
C145 B.t1 VSUBS 0.458692f
C146 B.t2 VSUBS 0.479699f
C147 B.t0 VSUBS 2.01572f
C148 B.n56 VSUBS 0.278634f
C149 B.n57 VSUBS 0.062203f
C150 B.n58 VSUBS 0.005824f
C151 B.n59 VSUBS 0.005824f
C152 B.n60 VSUBS 0.005824f
C153 B.n61 VSUBS 0.005824f
C154 B.n62 VSUBS 0.005824f
C155 B.n63 VSUBS 0.005824f
C156 B.n64 VSUBS 0.005824f
C157 B.n65 VSUBS 0.005824f
C158 B.n66 VSUBS 0.005824f
C159 B.n67 VSUBS 0.005824f
C160 B.n68 VSUBS 0.005824f
C161 B.n69 VSUBS 0.005824f
C162 B.n70 VSUBS 0.005824f
C163 B.n71 VSUBS 0.005824f
C164 B.n72 VSUBS 0.005824f
C165 B.n73 VSUBS 0.005824f
C166 B.n74 VSUBS 0.005824f
C167 B.n75 VSUBS 0.005824f
C168 B.n76 VSUBS 0.005824f
C169 B.n77 VSUBS 0.005824f
C170 B.n78 VSUBS 0.005824f
C171 B.n79 VSUBS 0.005824f
C172 B.n80 VSUBS 0.005824f
C173 B.n81 VSUBS 0.005824f
C174 B.n82 VSUBS 0.005824f
C175 B.n83 VSUBS 0.005824f
C176 B.n84 VSUBS 0.005824f
C177 B.n85 VSUBS 0.013605f
C178 B.n86 VSUBS 0.005824f
C179 B.n87 VSUBS 0.005824f
C180 B.n88 VSUBS 0.005824f
C181 B.n89 VSUBS 0.005824f
C182 B.n90 VSUBS 0.005824f
C183 B.n91 VSUBS 0.005824f
C184 B.n92 VSUBS 0.005824f
C185 B.n93 VSUBS 0.005824f
C186 B.n94 VSUBS 0.005824f
C187 B.n95 VSUBS 0.005824f
C188 B.n96 VSUBS 0.005824f
C189 B.n97 VSUBS 0.005824f
C190 B.n98 VSUBS 0.005824f
C191 B.n99 VSUBS 0.005824f
C192 B.n100 VSUBS 0.005824f
C193 B.n101 VSUBS 0.005824f
C194 B.n102 VSUBS 0.005824f
C195 B.n103 VSUBS 0.005824f
C196 B.n104 VSUBS 0.005824f
C197 B.n105 VSUBS 0.005824f
C198 B.n106 VSUBS 0.005824f
C199 B.n107 VSUBS 0.005824f
C200 B.n108 VSUBS 0.005824f
C201 B.n109 VSUBS 0.005824f
C202 B.n110 VSUBS 0.005824f
C203 B.n111 VSUBS 0.005824f
C204 B.n112 VSUBS 0.005824f
C205 B.n113 VSUBS 0.005824f
C206 B.n114 VSUBS 0.005824f
C207 B.n115 VSUBS 0.005824f
C208 B.n116 VSUBS 0.005824f
C209 B.n117 VSUBS 0.005824f
C210 B.n118 VSUBS 0.005824f
C211 B.n119 VSUBS 0.005824f
C212 B.n120 VSUBS 0.005824f
C213 B.n121 VSUBS 0.005824f
C214 B.n122 VSUBS 0.005824f
C215 B.n123 VSUBS 0.005824f
C216 B.n124 VSUBS 0.005824f
C217 B.n125 VSUBS 0.014487f
C218 B.n126 VSUBS 0.005824f
C219 B.n127 VSUBS 0.005824f
C220 B.n128 VSUBS 0.005824f
C221 B.n129 VSUBS 0.005824f
C222 B.n130 VSUBS 0.005824f
C223 B.n131 VSUBS 0.005824f
C224 B.n132 VSUBS 0.005824f
C225 B.n133 VSUBS 0.005824f
C226 B.n134 VSUBS 0.005824f
C227 B.n135 VSUBS 0.005824f
C228 B.n136 VSUBS 0.005824f
C229 B.n137 VSUBS 0.005824f
C230 B.n138 VSUBS 0.005824f
C231 B.n139 VSUBS 0.005824f
C232 B.n140 VSUBS 0.005824f
C233 B.n141 VSUBS 0.005824f
C234 B.n142 VSUBS 0.005824f
C235 B.n143 VSUBS 0.005824f
C236 B.n144 VSUBS 0.005824f
C237 B.n145 VSUBS 0.005824f
C238 B.n146 VSUBS 0.005824f
C239 B.n147 VSUBS 0.005824f
C240 B.n148 VSUBS 0.005824f
C241 B.n149 VSUBS 0.005824f
C242 B.n150 VSUBS 0.005824f
C243 B.n151 VSUBS 0.005824f
C244 B.n152 VSUBS 0.004025f
C245 B.n153 VSUBS 0.005824f
C246 B.n154 VSUBS 0.005824f
C247 B.n155 VSUBS 0.005824f
C248 B.n156 VSUBS 0.005824f
C249 B.n157 VSUBS 0.005824f
C250 B.t11 VSUBS 0.458706f
C251 B.t10 VSUBS 0.47971f
C252 B.t9 VSUBS 2.01572f
C253 B.n158 VSUBS 0.278622f
C254 B.n159 VSUBS 0.062188f
C255 B.n160 VSUBS 0.005824f
C256 B.n161 VSUBS 0.005824f
C257 B.n162 VSUBS 0.005824f
C258 B.n163 VSUBS 0.005824f
C259 B.n164 VSUBS 0.005824f
C260 B.n165 VSUBS 0.005824f
C261 B.n166 VSUBS 0.005824f
C262 B.n167 VSUBS 0.005824f
C263 B.n168 VSUBS 0.005824f
C264 B.n169 VSUBS 0.005824f
C265 B.n170 VSUBS 0.005824f
C266 B.n171 VSUBS 0.005824f
C267 B.n172 VSUBS 0.005824f
C268 B.n173 VSUBS 0.005824f
C269 B.n174 VSUBS 0.005824f
C270 B.n175 VSUBS 0.005824f
C271 B.n176 VSUBS 0.005824f
C272 B.n177 VSUBS 0.005824f
C273 B.n178 VSUBS 0.005824f
C274 B.n179 VSUBS 0.005824f
C275 B.n180 VSUBS 0.005824f
C276 B.n181 VSUBS 0.005824f
C277 B.n182 VSUBS 0.005824f
C278 B.n183 VSUBS 0.005824f
C279 B.n184 VSUBS 0.005824f
C280 B.n185 VSUBS 0.005824f
C281 B.n186 VSUBS 0.014487f
C282 B.n187 VSUBS 0.005824f
C283 B.n188 VSUBS 0.005824f
C284 B.n189 VSUBS 0.005824f
C285 B.n190 VSUBS 0.005824f
C286 B.n191 VSUBS 0.005824f
C287 B.n192 VSUBS 0.005824f
C288 B.n193 VSUBS 0.005824f
C289 B.n194 VSUBS 0.005824f
C290 B.n195 VSUBS 0.005824f
C291 B.n196 VSUBS 0.005824f
C292 B.n197 VSUBS 0.005824f
C293 B.n198 VSUBS 0.005824f
C294 B.n199 VSUBS 0.005824f
C295 B.n200 VSUBS 0.005824f
C296 B.n201 VSUBS 0.005824f
C297 B.n202 VSUBS 0.005824f
C298 B.n203 VSUBS 0.005824f
C299 B.n204 VSUBS 0.005824f
C300 B.n205 VSUBS 0.005824f
C301 B.n206 VSUBS 0.005824f
C302 B.n207 VSUBS 0.005824f
C303 B.n208 VSUBS 0.005824f
C304 B.n209 VSUBS 0.005824f
C305 B.n210 VSUBS 0.005824f
C306 B.n211 VSUBS 0.005824f
C307 B.n212 VSUBS 0.005824f
C308 B.n213 VSUBS 0.005824f
C309 B.n214 VSUBS 0.005824f
C310 B.n215 VSUBS 0.005824f
C311 B.n216 VSUBS 0.005824f
C312 B.n217 VSUBS 0.005824f
C313 B.n218 VSUBS 0.005824f
C314 B.n219 VSUBS 0.005824f
C315 B.n220 VSUBS 0.005824f
C316 B.n221 VSUBS 0.005824f
C317 B.n222 VSUBS 0.005824f
C318 B.n223 VSUBS 0.005824f
C319 B.n224 VSUBS 0.005824f
C320 B.n225 VSUBS 0.005824f
C321 B.n226 VSUBS 0.005824f
C322 B.n227 VSUBS 0.005824f
C323 B.n228 VSUBS 0.005824f
C324 B.n229 VSUBS 0.005824f
C325 B.n230 VSUBS 0.005824f
C326 B.n231 VSUBS 0.005824f
C327 B.n232 VSUBS 0.005824f
C328 B.n233 VSUBS 0.005824f
C329 B.n234 VSUBS 0.005824f
C330 B.n235 VSUBS 0.005824f
C331 B.n236 VSUBS 0.005824f
C332 B.n237 VSUBS 0.005824f
C333 B.n238 VSUBS 0.005824f
C334 B.n239 VSUBS 0.005824f
C335 B.n240 VSUBS 0.005824f
C336 B.n241 VSUBS 0.005824f
C337 B.n242 VSUBS 0.005824f
C338 B.n243 VSUBS 0.005824f
C339 B.n244 VSUBS 0.005824f
C340 B.n245 VSUBS 0.005824f
C341 B.n246 VSUBS 0.005824f
C342 B.n247 VSUBS 0.005824f
C343 B.n248 VSUBS 0.005824f
C344 B.n249 VSUBS 0.005824f
C345 B.n250 VSUBS 0.005824f
C346 B.n251 VSUBS 0.005824f
C347 B.n252 VSUBS 0.005824f
C348 B.n253 VSUBS 0.005824f
C349 B.n254 VSUBS 0.005824f
C350 B.n255 VSUBS 0.005824f
C351 B.n256 VSUBS 0.005824f
C352 B.n257 VSUBS 0.005824f
C353 B.n258 VSUBS 0.005824f
C354 B.n259 VSUBS 0.005824f
C355 B.n260 VSUBS 0.005824f
C356 B.n261 VSUBS 0.013605f
C357 B.n262 VSUBS 0.013605f
C358 B.n263 VSUBS 0.014487f
C359 B.n264 VSUBS 0.005824f
C360 B.n265 VSUBS 0.005824f
C361 B.n266 VSUBS 0.005824f
C362 B.n267 VSUBS 0.005824f
C363 B.n268 VSUBS 0.005824f
C364 B.n269 VSUBS 0.005824f
C365 B.n270 VSUBS 0.005824f
C366 B.n271 VSUBS 0.005824f
C367 B.n272 VSUBS 0.005824f
C368 B.n273 VSUBS 0.005824f
C369 B.n274 VSUBS 0.005824f
C370 B.n275 VSUBS 0.005824f
C371 B.n276 VSUBS 0.005824f
C372 B.n277 VSUBS 0.005824f
C373 B.n278 VSUBS 0.005824f
C374 B.n279 VSUBS 0.005824f
C375 B.n280 VSUBS 0.005824f
C376 B.n281 VSUBS 0.005824f
C377 B.n282 VSUBS 0.005824f
C378 B.n283 VSUBS 0.005824f
C379 B.n284 VSUBS 0.005824f
C380 B.n285 VSUBS 0.005824f
C381 B.n286 VSUBS 0.005824f
C382 B.n287 VSUBS 0.005824f
C383 B.n288 VSUBS 0.005824f
C384 B.n289 VSUBS 0.005824f
C385 B.n290 VSUBS 0.005824f
C386 B.n291 VSUBS 0.005824f
C387 B.n292 VSUBS 0.005824f
C388 B.n293 VSUBS 0.005824f
C389 B.n294 VSUBS 0.005824f
C390 B.n295 VSUBS 0.005824f
C391 B.n296 VSUBS 0.005824f
C392 B.n297 VSUBS 0.005824f
C393 B.n298 VSUBS 0.005824f
C394 B.n299 VSUBS 0.005824f
C395 B.n300 VSUBS 0.005824f
C396 B.n301 VSUBS 0.005824f
C397 B.n302 VSUBS 0.005824f
C398 B.n303 VSUBS 0.005824f
C399 B.n304 VSUBS 0.005824f
C400 B.n305 VSUBS 0.005824f
C401 B.n306 VSUBS 0.005824f
C402 B.n307 VSUBS 0.005824f
C403 B.n308 VSUBS 0.005824f
C404 B.n309 VSUBS 0.005824f
C405 B.n310 VSUBS 0.005824f
C406 B.n311 VSUBS 0.005824f
C407 B.n312 VSUBS 0.005824f
C408 B.n313 VSUBS 0.005824f
C409 B.n314 VSUBS 0.005824f
C410 B.n315 VSUBS 0.005824f
C411 B.n316 VSUBS 0.005824f
C412 B.n317 VSUBS 0.005824f
C413 B.n318 VSUBS 0.005824f
C414 B.n319 VSUBS 0.005824f
C415 B.n320 VSUBS 0.005824f
C416 B.n321 VSUBS 0.005824f
C417 B.n322 VSUBS 0.005824f
C418 B.n323 VSUBS 0.005824f
C419 B.n324 VSUBS 0.005824f
C420 B.n325 VSUBS 0.005824f
C421 B.n326 VSUBS 0.005824f
C422 B.n327 VSUBS 0.005824f
C423 B.n328 VSUBS 0.005824f
C424 B.n329 VSUBS 0.005824f
C425 B.n330 VSUBS 0.005824f
C426 B.n331 VSUBS 0.005824f
C427 B.n332 VSUBS 0.005824f
C428 B.n333 VSUBS 0.005824f
C429 B.n334 VSUBS 0.005824f
C430 B.n335 VSUBS 0.005824f
C431 B.n336 VSUBS 0.005824f
C432 B.n337 VSUBS 0.005824f
C433 B.n338 VSUBS 0.005824f
C434 B.n339 VSUBS 0.005824f
C435 B.n340 VSUBS 0.005824f
C436 B.n341 VSUBS 0.005824f
C437 B.n342 VSUBS 0.005824f
C438 B.n343 VSUBS 0.005824f
C439 B.n344 VSUBS 0.004025f
C440 B.n345 VSUBS 0.013493f
C441 B.n346 VSUBS 0.004711f
C442 B.n347 VSUBS 0.005824f
C443 B.n348 VSUBS 0.005824f
C444 B.n349 VSUBS 0.005824f
C445 B.n350 VSUBS 0.005824f
C446 B.n351 VSUBS 0.005824f
C447 B.n352 VSUBS 0.005824f
C448 B.n353 VSUBS 0.005824f
C449 B.n354 VSUBS 0.005824f
C450 B.n355 VSUBS 0.005824f
C451 B.n356 VSUBS 0.005824f
C452 B.n357 VSUBS 0.005824f
C453 B.t5 VSUBS 0.458692f
C454 B.t4 VSUBS 0.479699f
C455 B.t3 VSUBS 2.01572f
C456 B.n358 VSUBS 0.278634f
C457 B.n359 VSUBS 0.062203f
C458 B.n360 VSUBS 0.013493f
C459 B.n361 VSUBS 0.004711f
C460 B.n362 VSUBS 0.005824f
C461 B.n363 VSUBS 0.005824f
C462 B.n364 VSUBS 0.005824f
C463 B.n365 VSUBS 0.005824f
C464 B.n366 VSUBS 0.005824f
C465 B.n367 VSUBS 0.005824f
C466 B.n368 VSUBS 0.005824f
C467 B.n369 VSUBS 0.005824f
C468 B.n370 VSUBS 0.005824f
C469 B.n371 VSUBS 0.005824f
C470 B.n372 VSUBS 0.005824f
C471 B.n373 VSUBS 0.005824f
C472 B.n374 VSUBS 0.005824f
C473 B.n375 VSUBS 0.005824f
C474 B.n376 VSUBS 0.005824f
C475 B.n377 VSUBS 0.005824f
C476 B.n378 VSUBS 0.005824f
C477 B.n379 VSUBS 0.005824f
C478 B.n380 VSUBS 0.005824f
C479 B.n381 VSUBS 0.005824f
C480 B.n382 VSUBS 0.005824f
C481 B.n383 VSUBS 0.005824f
C482 B.n384 VSUBS 0.005824f
C483 B.n385 VSUBS 0.005824f
C484 B.n386 VSUBS 0.005824f
C485 B.n387 VSUBS 0.005824f
C486 B.n388 VSUBS 0.005824f
C487 B.n389 VSUBS 0.005824f
C488 B.n390 VSUBS 0.005824f
C489 B.n391 VSUBS 0.005824f
C490 B.n392 VSUBS 0.005824f
C491 B.n393 VSUBS 0.005824f
C492 B.n394 VSUBS 0.005824f
C493 B.n395 VSUBS 0.005824f
C494 B.n396 VSUBS 0.005824f
C495 B.n397 VSUBS 0.005824f
C496 B.n398 VSUBS 0.005824f
C497 B.n399 VSUBS 0.005824f
C498 B.n400 VSUBS 0.005824f
C499 B.n401 VSUBS 0.005824f
C500 B.n402 VSUBS 0.005824f
C501 B.n403 VSUBS 0.005824f
C502 B.n404 VSUBS 0.005824f
C503 B.n405 VSUBS 0.005824f
C504 B.n406 VSUBS 0.005824f
C505 B.n407 VSUBS 0.005824f
C506 B.n408 VSUBS 0.005824f
C507 B.n409 VSUBS 0.005824f
C508 B.n410 VSUBS 0.005824f
C509 B.n411 VSUBS 0.005824f
C510 B.n412 VSUBS 0.005824f
C511 B.n413 VSUBS 0.005824f
C512 B.n414 VSUBS 0.005824f
C513 B.n415 VSUBS 0.005824f
C514 B.n416 VSUBS 0.005824f
C515 B.n417 VSUBS 0.005824f
C516 B.n418 VSUBS 0.005824f
C517 B.n419 VSUBS 0.005824f
C518 B.n420 VSUBS 0.005824f
C519 B.n421 VSUBS 0.005824f
C520 B.n422 VSUBS 0.005824f
C521 B.n423 VSUBS 0.005824f
C522 B.n424 VSUBS 0.005824f
C523 B.n425 VSUBS 0.005824f
C524 B.n426 VSUBS 0.005824f
C525 B.n427 VSUBS 0.005824f
C526 B.n428 VSUBS 0.005824f
C527 B.n429 VSUBS 0.005824f
C528 B.n430 VSUBS 0.005824f
C529 B.n431 VSUBS 0.005824f
C530 B.n432 VSUBS 0.005824f
C531 B.n433 VSUBS 0.005824f
C532 B.n434 VSUBS 0.005824f
C533 B.n435 VSUBS 0.005824f
C534 B.n436 VSUBS 0.005824f
C535 B.n437 VSUBS 0.005824f
C536 B.n438 VSUBS 0.005824f
C537 B.n439 VSUBS 0.005824f
C538 B.n440 VSUBS 0.005824f
C539 B.n441 VSUBS 0.005824f
C540 B.n442 VSUBS 0.005824f
C541 B.n443 VSUBS 0.005824f
C542 B.n444 VSUBS 0.01383f
C543 B.n445 VSUBS 0.014262f
C544 B.n446 VSUBS 0.013605f
C545 B.n447 VSUBS 0.005824f
C546 B.n448 VSUBS 0.005824f
C547 B.n449 VSUBS 0.005824f
C548 B.n450 VSUBS 0.005824f
C549 B.n451 VSUBS 0.005824f
C550 B.n452 VSUBS 0.005824f
C551 B.n453 VSUBS 0.005824f
C552 B.n454 VSUBS 0.005824f
C553 B.n455 VSUBS 0.005824f
C554 B.n456 VSUBS 0.005824f
C555 B.n457 VSUBS 0.005824f
C556 B.n458 VSUBS 0.005824f
C557 B.n459 VSUBS 0.005824f
C558 B.n460 VSUBS 0.005824f
C559 B.n461 VSUBS 0.005824f
C560 B.n462 VSUBS 0.005824f
C561 B.n463 VSUBS 0.005824f
C562 B.n464 VSUBS 0.005824f
C563 B.n465 VSUBS 0.005824f
C564 B.n466 VSUBS 0.005824f
C565 B.n467 VSUBS 0.005824f
C566 B.n468 VSUBS 0.005824f
C567 B.n469 VSUBS 0.005824f
C568 B.n470 VSUBS 0.005824f
C569 B.n471 VSUBS 0.005824f
C570 B.n472 VSUBS 0.005824f
C571 B.n473 VSUBS 0.005824f
C572 B.n474 VSUBS 0.005824f
C573 B.n475 VSUBS 0.005824f
C574 B.n476 VSUBS 0.005824f
C575 B.n477 VSUBS 0.005824f
C576 B.n478 VSUBS 0.005824f
C577 B.n479 VSUBS 0.005824f
C578 B.n480 VSUBS 0.005824f
C579 B.n481 VSUBS 0.005824f
C580 B.n482 VSUBS 0.005824f
C581 B.n483 VSUBS 0.005824f
C582 B.n484 VSUBS 0.005824f
C583 B.n485 VSUBS 0.005824f
C584 B.n486 VSUBS 0.005824f
C585 B.n487 VSUBS 0.005824f
C586 B.n488 VSUBS 0.005824f
C587 B.n489 VSUBS 0.005824f
C588 B.n490 VSUBS 0.005824f
C589 B.n491 VSUBS 0.005824f
C590 B.n492 VSUBS 0.005824f
C591 B.n493 VSUBS 0.005824f
C592 B.n494 VSUBS 0.005824f
C593 B.n495 VSUBS 0.005824f
C594 B.n496 VSUBS 0.005824f
C595 B.n497 VSUBS 0.005824f
C596 B.n498 VSUBS 0.005824f
C597 B.n499 VSUBS 0.005824f
C598 B.n500 VSUBS 0.005824f
C599 B.n501 VSUBS 0.005824f
C600 B.n502 VSUBS 0.005824f
C601 B.n503 VSUBS 0.005824f
C602 B.n504 VSUBS 0.005824f
C603 B.n505 VSUBS 0.005824f
C604 B.n506 VSUBS 0.005824f
C605 B.n507 VSUBS 0.005824f
C606 B.n508 VSUBS 0.005824f
C607 B.n509 VSUBS 0.005824f
C608 B.n510 VSUBS 0.005824f
C609 B.n511 VSUBS 0.005824f
C610 B.n512 VSUBS 0.005824f
C611 B.n513 VSUBS 0.005824f
C612 B.n514 VSUBS 0.005824f
C613 B.n515 VSUBS 0.005824f
C614 B.n516 VSUBS 0.005824f
C615 B.n517 VSUBS 0.005824f
C616 B.n518 VSUBS 0.005824f
C617 B.n519 VSUBS 0.005824f
C618 B.n520 VSUBS 0.005824f
C619 B.n521 VSUBS 0.005824f
C620 B.n522 VSUBS 0.005824f
C621 B.n523 VSUBS 0.005824f
C622 B.n524 VSUBS 0.005824f
C623 B.n525 VSUBS 0.005824f
C624 B.n526 VSUBS 0.005824f
C625 B.n527 VSUBS 0.005824f
C626 B.n528 VSUBS 0.005824f
C627 B.n529 VSUBS 0.005824f
C628 B.n530 VSUBS 0.005824f
C629 B.n531 VSUBS 0.005824f
C630 B.n532 VSUBS 0.005824f
C631 B.n533 VSUBS 0.005824f
C632 B.n534 VSUBS 0.005824f
C633 B.n535 VSUBS 0.005824f
C634 B.n536 VSUBS 0.005824f
C635 B.n537 VSUBS 0.005824f
C636 B.n538 VSUBS 0.005824f
C637 B.n539 VSUBS 0.005824f
C638 B.n540 VSUBS 0.005824f
C639 B.n541 VSUBS 0.005824f
C640 B.n542 VSUBS 0.005824f
C641 B.n543 VSUBS 0.005824f
C642 B.n544 VSUBS 0.005824f
C643 B.n545 VSUBS 0.005824f
C644 B.n546 VSUBS 0.005824f
C645 B.n547 VSUBS 0.005824f
C646 B.n548 VSUBS 0.005824f
C647 B.n549 VSUBS 0.005824f
C648 B.n550 VSUBS 0.005824f
C649 B.n551 VSUBS 0.005824f
C650 B.n552 VSUBS 0.005824f
C651 B.n553 VSUBS 0.005824f
C652 B.n554 VSUBS 0.005824f
C653 B.n555 VSUBS 0.005824f
C654 B.n556 VSUBS 0.005824f
C655 B.n557 VSUBS 0.005824f
C656 B.n558 VSUBS 0.005824f
C657 B.n559 VSUBS 0.005824f
C658 B.n560 VSUBS 0.005824f
C659 B.n561 VSUBS 0.005824f
C660 B.n562 VSUBS 0.005824f
C661 B.n563 VSUBS 0.005824f
C662 B.n564 VSUBS 0.013605f
C663 B.n565 VSUBS 0.014487f
C664 B.n566 VSUBS 0.014487f
C665 B.n567 VSUBS 0.005824f
C666 B.n568 VSUBS 0.005824f
C667 B.n569 VSUBS 0.005824f
C668 B.n570 VSUBS 0.005824f
C669 B.n571 VSUBS 0.005824f
C670 B.n572 VSUBS 0.005824f
C671 B.n573 VSUBS 0.005824f
C672 B.n574 VSUBS 0.005824f
C673 B.n575 VSUBS 0.005824f
C674 B.n576 VSUBS 0.005824f
C675 B.n577 VSUBS 0.005824f
C676 B.n578 VSUBS 0.005824f
C677 B.n579 VSUBS 0.005824f
C678 B.n580 VSUBS 0.005824f
C679 B.n581 VSUBS 0.005824f
C680 B.n582 VSUBS 0.005824f
C681 B.n583 VSUBS 0.005824f
C682 B.n584 VSUBS 0.005824f
C683 B.n585 VSUBS 0.005824f
C684 B.n586 VSUBS 0.005824f
C685 B.n587 VSUBS 0.005824f
C686 B.n588 VSUBS 0.005824f
C687 B.n589 VSUBS 0.005824f
C688 B.n590 VSUBS 0.005824f
C689 B.n591 VSUBS 0.005824f
C690 B.n592 VSUBS 0.005824f
C691 B.n593 VSUBS 0.005824f
C692 B.n594 VSUBS 0.005824f
C693 B.n595 VSUBS 0.005824f
C694 B.n596 VSUBS 0.005824f
C695 B.n597 VSUBS 0.005824f
C696 B.n598 VSUBS 0.005824f
C697 B.n599 VSUBS 0.005824f
C698 B.n600 VSUBS 0.005824f
C699 B.n601 VSUBS 0.005824f
C700 B.n602 VSUBS 0.005824f
C701 B.n603 VSUBS 0.005824f
C702 B.n604 VSUBS 0.005824f
C703 B.n605 VSUBS 0.005824f
C704 B.n606 VSUBS 0.005824f
C705 B.n607 VSUBS 0.005824f
C706 B.n608 VSUBS 0.005824f
C707 B.n609 VSUBS 0.005824f
C708 B.n610 VSUBS 0.005824f
C709 B.n611 VSUBS 0.005824f
C710 B.n612 VSUBS 0.005824f
C711 B.n613 VSUBS 0.005824f
C712 B.n614 VSUBS 0.005824f
C713 B.n615 VSUBS 0.005824f
C714 B.n616 VSUBS 0.005824f
C715 B.n617 VSUBS 0.005824f
C716 B.n618 VSUBS 0.005824f
C717 B.n619 VSUBS 0.005824f
C718 B.n620 VSUBS 0.005824f
C719 B.n621 VSUBS 0.005824f
C720 B.n622 VSUBS 0.005824f
C721 B.n623 VSUBS 0.005824f
C722 B.n624 VSUBS 0.005824f
C723 B.n625 VSUBS 0.005824f
C724 B.n626 VSUBS 0.005824f
C725 B.n627 VSUBS 0.005824f
C726 B.n628 VSUBS 0.005824f
C727 B.n629 VSUBS 0.005824f
C728 B.n630 VSUBS 0.005824f
C729 B.n631 VSUBS 0.005824f
C730 B.n632 VSUBS 0.005824f
C731 B.n633 VSUBS 0.005824f
C732 B.n634 VSUBS 0.005824f
C733 B.n635 VSUBS 0.005824f
C734 B.n636 VSUBS 0.005824f
C735 B.n637 VSUBS 0.005824f
C736 B.n638 VSUBS 0.005824f
C737 B.n639 VSUBS 0.005824f
C738 B.n640 VSUBS 0.005824f
C739 B.n641 VSUBS 0.005824f
C740 B.n642 VSUBS 0.005824f
C741 B.n643 VSUBS 0.005824f
C742 B.n644 VSUBS 0.005824f
C743 B.n645 VSUBS 0.005824f
C744 B.n646 VSUBS 0.005824f
C745 B.n647 VSUBS 0.004025f
C746 B.n648 VSUBS 0.013493f
C747 B.n649 VSUBS 0.004711f
C748 B.n650 VSUBS 0.005824f
C749 B.n651 VSUBS 0.005824f
C750 B.n652 VSUBS 0.005824f
C751 B.n653 VSUBS 0.005824f
C752 B.n654 VSUBS 0.005824f
C753 B.n655 VSUBS 0.005824f
C754 B.n656 VSUBS 0.005824f
C755 B.n657 VSUBS 0.005824f
C756 B.n658 VSUBS 0.005824f
C757 B.n659 VSUBS 0.005824f
C758 B.n660 VSUBS 0.005824f
C759 B.n661 VSUBS 0.004711f
C760 B.n662 VSUBS 0.013493f
C761 B.n663 VSUBS 0.004025f
C762 B.n664 VSUBS 0.005824f
C763 B.n665 VSUBS 0.005824f
C764 B.n666 VSUBS 0.005824f
C765 B.n667 VSUBS 0.005824f
C766 B.n668 VSUBS 0.005824f
C767 B.n669 VSUBS 0.005824f
C768 B.n670 VSUBS 0.005824f
C769 B.n671 VSUBS 0.005824f
C770 B.n672 VSUBS 0.005824f
C771 B.n673 VSUBS 0.005824f
C772 B.n674 VSUBS 0.005824f
C773 B.n675 VSUBS 0.005824f
C774 B.n676 VSUBS 0.005824f
C775 B.n677 VSUBS 0.005824f
C776 B.n678 VSUBS 0.005824f
C777 B.n679 VSUBS 0.005824f
C778 B.n680 VSUBS 0.005824f
C779 B.n681 VSUBS 0.005824f
C780 B.n682 VSUBS 0.005824f
C781 B.n683 VSUBS 0.005824f
C782 B.n684 VSUBS 0.005824f
C783 B.n685 VSUBS 0.005824f
C784 B.n686 VSUBS 0.005824f
C785 B.n687 VSUBS 0.005824f
C786 B.n688 VSUBS 0.005824f
C787 B.n689 VSUBS 0.005824f
C788 B.n690 VSUBS 0.005824f
C789 B.n691 VSUBS 0.005824f
C790 B.n692 VSUBS 0.005824f
C791 B.n693 VSUBS 0.005824f
C792 B.n694 VSUBS 0.005824f
C793 B.n695 VSUBS 0.005824f
C794 B.n696 VSUBS 0.005824f
C795 B.n697 VSUBS 0.005824f
C796 B.n698 VSUBS 0.005824f
C797 B.n699 VSUBS 0.005824f
C798 B.n700 VSUBS 0.005824f
C799 B.n701 VSUBS 0.005824f
C800 B.n702 VSUBS 0.005824f
C801 B.n703 VSUBS 0.005824f
C802 B.n704 VSUBS 0.005824f
C803 B.n705 VSUBS 0.005824f
C804 B.n706 VSUBS 0.005824f
C805 B.n707 VSUBS 0.005824f
C806 B.n708 VSUBS 0.005824f
C807 B.n709 VSUBS 0.005824f
C808 B.n710 VSUBS 0.005824f
C809 B.n711 VSUBS 0.005824f
C810 B.n712 VSUBS 0.005824f
C811 B.n713 VSUBS 0.005824f
C812 B.n714 VSUBS 0.005824f
C813 B.n715 VSUBS 0.005824f
C814 B.n716 VSUBS 0.005824f
C815 B.n717 VSUBS 0.005824f
C816 B.n718 VSUBS 0.005824f
C817 B.n719 VSUBS 0.005824f
C818 B.n720 VSUBS 0.005824f
C819 B.n721 VSUBS 0.005824f
C820 B.n722 VSUBS 0.005824f
C821 B.n723 VSUBS 0.005824f
C822 B.n724 VSUBS 0.005824f
C823 B.n725 VSUBS 0.005824f
C824 B.n726 VSUBS 0.005824f
C825 B.n727 VSUBS 0.005824f
C826 B.n728 VSUBS 0.005824f
C827 B.n729 VSUBS 0.005824f
C828 B.n730 VSUBS 0.005824f
C829 B.n731 VSUBS 0.005824f
C830 B.n732 VSUBS 0.005824f
C831 B.n733 VSUBS 0.005824f
C832 B.n734 VSUBS 0.005824f
C833 B.n735 VSUBS 0.005824f
C834 B.n736 VSUBS 0.005824f
C835 B.n737 VSUBS 0.005824f
C836 B.n738 VSUBS 0.005824f
C837 B.n739 VSUBS 0.005824f
C838 B.n740 VSUBS 0.005824f
C839 B.n741 VSUBS 0.005824f
C840 B.n742 VSUBS 0.005824f
C841 B.n743 VSUBS 0.005824f
C842 B.n744 VSUBS 0.014487f
C843 B.n745 VSUBS 0.014487f
C844 B.n746 VSUBS 0.013605f
C845 B.n747 VSUBS 0.005824f
C846 B.n748 VSUBS 0.005824f
C847 B.n749 VSUBS 0.005824f
C848 B.n750 VSUBS 0.005824f
C849 B.n751 VSUBS 0.005824f
C850 B.n752 VSUBS 0.005824f
C851 B.n753 VSUBS 0.005824f
C852 B.n754 VSUBS 0.005824f
C853 B.n755 VSUBS 0.005824f
C854 B.n756 VSUBS 0.005824f
C855 B.n757 VSUBS 0.005824f
C856 B.n758 VSUBS 0.005824f
C857 B.n759 VSUBS 0.005824f
C858 B.n760 VSUBS 0.005824f
C859 B.n761 VSUBS 0.005824f
C860 B.n762 VSUBS 0.005824f
C861 B.n763 VSUBS 0.005824f
C862 B.n764 VSUBS 0.005824f
C863 B.n765 VSUBS 0.005824f
C864 B.n766 VSUBS 0.005824f
C865 B.n767 VSUBS 0.005824f
C866 B.n768 VSUBS 0.005824f
C867 B.n769 VSUBS 0.005824f
C868 B.n770 VSUBS 0.005824f
C869 B.n771 VSUBS 0.005824f
C870 B.n772 VSUBS 0.005824f
C871 B.n773 VSUBS 0.005824f
C872 B.n774 VSUBS 0.005824f
C873 B.n775 VSUBS 0.005824f
C874 B.n776 VSUBS 0.005824f
C875 B.n777 VSUBS 0.005824f
C876 B.n778 VSUBS 0.005824f
C877 B.n779 VSUBS 0.005824f
C878 B.n780 VSUBS 0.005824f
C879 B.n781 VSUBS 0.005824f
C880 B.n782 VSUBS 0.005824f
C881 B.n783 VSUBS 0.005824f
C882 B.n784 VSUBS 0.005824f
C883 B.n785 VSUBS 0.005824f
C884 B.n786 VSUBS 0.005824f
C885 B.n787 VSUBS 0.005824f
C886 B.n788 VSUBS 0.005824f
C887 B.n789 VSUBS 0.005824f
C888 B.n790 VSUBS 0.005824f
C889 B.n791 VSUBS 0.005824f
C890 B.n792 VSUBS 0.005824f
C891 B.n793 VSUBS 0.005824f
C892 B.n794 VSUBS 0.005824f
C893 B.n795 VSUBS 0.005824f
C894 B.n796 VSUBS 0.005824f
C895 B.n797 VSUBS 0.005824f
C896 B.n798 VSUBS 0.005824f
C897 B.n799 VSUBS 0.005824f
C898 B.n800 VSUBS 0.005824f
C899 B.n801 VSUBS 0.005824f
C900 B.n802 VSUBS 0.005824f
C901 B.n803 VSUBS 0.0076f
C902 B.n804 VSUBS 0.008096f
C903 B.n805 VSUBS 0.0161f
.ends

