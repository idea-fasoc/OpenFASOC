* NGSPICE file created from diff_pair_sample_0043.ext - technology: sky130A

.subckt diff_pair_sample_0043 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=0 ps=0 w=9.69 l=1.06
X1 VDD1.t1 VP.t0 VTAIL.t2 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=3.7791 ps=20.16 w=9.69 l=1.06
X2 VDD1.t0 VP.t1 VTAIL.t3 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=3.7791 ps=20.16 w=9.69 l=1.06
X3 B.t8 B.t6 B.t7 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=0 ps=0 w=9.69 l=1.06
X4 B.t5 B.t3 B.t4 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=0 ps=0 w=9.69 l=1.06
X5 B.t2 B.t0 B.t1 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=0 ps=0 w=9.69 l=1.06
X6 VDD2.t1 VN.t0 VTAIL.t1 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=3.7791 ps=20.16 w=9.69 l=1.06
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1526_n2910# sky130_fd_pr__pfet_01v8 ad=3.7791 pd=20.16 as=3.7791 ps=20.16 w=9.69 l=1.06
R0 B.n264 B.n71 585
R1 B.n263 B.n262 585
R2 B.n261 B.n72 585
R3 B.n260 B.n259 585
R4 B.n258 B.n73 585
R5 B.n257 B.n256 585
R6 B.n255 B.n74 585
R7 B.n254 B.n253 585
R8 B.n252 B.n75 585
R9 B.n251 B.n250 585
R10 B.n249 B.n76 585
R11 B.n248 B.n247 585
R12 B.n246 B.n77 585
R13 B.n245 B.n244 585
R14 B.n243 B.n78 585
R15 B.n242 B.n241 585
R16 B.n240 B.n79 585
R17 B.n239 B.n238 585
R18 B.n237 B.n80 585
R19 B.n236 B.n235 585
R20 B.n234 B.n81 585
R21 B.n233 B.n232 585
R22 B.n231 B.n82 585
R23 B.n230 B.n229 585
R24 B.n228 B.n83 585
R25 B.n227 B.n226 585
R26 B.n225 B.n84 585
R27 B.n224 B.n223 585
R28 B.n222 B.n85 585
R29 B.n221 B.n220 585
R30 B.n219 B.n86 585
R31 B.n218 B.n217 585
R32 B.n216 B.n87 585
R33 B.n215 B.n214 585
R34 B.n213 B.n88 585
R35 B.n212 B.n211 585
R36 B.n207 B.n89 585
R37 B.n206 B.n205 585
R38 B.n204 B.n90 585
R39 B.n203 B.n202 585
R40 B.n201 B.n91 585
R41 B.n200 B.n199 585
R42 B.n198 B.n92 585
R43 B.n197 B.n196 585
R44 B.n194 B.n93 585
R45 B.n193 B.n192 585
R46 B.n191 B.n96 585
R47 B.n190 B.n189 585
R48 B.n188 B.n97 585
R49 B.n187 B.n186 585
R50 B.n185 B.n98 585
R51 B.n184 B.n183 585
R52 B.n182 B.n99 585
R53 B.n181 B.n180 585
R54 B.n179 B.n100 585
R55 B.n178 B.n177 585
R56 B.n176 B.n101 585
R57 B.n175 B.n174 585
R58 B.n173 B.n102 585
R59 B.n172 B.n171 585
R60 B.n170 B.n103 585
R61 B.n169 B.n168 585
R62 B.n167 B.n104 585
R63 B.n166 B.n165 585
R64 B.n164 B.n105 585
R65 B.n163 B.n162 585
R66 B.n161 B.n106 585
R67 B.n160 B.n159 585
R68 B.n158 B.n107 585
R69 B.n157 B.n156 585
R70 B.n155 B.n108 585
R71 B.n154 B.n153 585
R72 B.n152 B.n109 585
R73 B.n151 B.n150 585
R74 B.n149 B.n110 585
R75 B.n148 B.n147 585
R76 B.n146 B.n111 585
R77 B.n145 B.n144 585
R78 B.n143 B.n112 585
R79 B.n266 B.n265 585
R80 B.n267 B.n70 585
R81 B.n269 B.n268 585
R82 B.n270 B.n69 585
R83 B.n272 B.n271 585
R84 B.n273 B.n68 585
R85 B.n275 B.n274 585
R86 B.n276 B.n67 585
R87 B.n278 B.n277 585
R88 B.n279 B.n66 585
R89 B.n281 B.n280 585
R90 B.n282 B.n65 585
R91 B.n284 B.n283 585
R92 B.n285 B.n64 585
R93 B.n287 B.n286 585
R94 B.n288 B.n63 585
R95 B.n290 B.n289 585
R96 B.n291 B.n62 585
R97 B.n293 B.n292 585
R98 B.n294 B.n61 585
R99 B.n296 B.n295 585
R100 B.n297 B.n60 585
R101 B.n299 B.n298 585
R102 B.n300 B.n59 585
R103 B.n302 B.n301 585
R104 B.n303 B.n58 585
R105 B.n305 B.n304 585
R106 B.n306 B.n57 585
R107 B.n308 B.n307 585
R108 B.n309 B.n56 585
R109 B.n311 B.n310 585
R110 B.n312 B.n55 585
R111 B.n314 B.n313 585
R112 B.n315 B.n54 585
R113 B.n435 B.n10 585
R114 B.n434 B.n433 585
R115 B.n432 B.n11 585
R116 B.n431 B.n430 585
R117 B.n429 B.n12 585
R118 B.n428 B.n427 585
R119 B.n426 B.n13 585
R120 B.n425 B.n424 585
R121 B.n423 B.n14 585
R122 B.n422 B.n421 585
R123 B.n420 B.n15 585
R124 B.n419 B.n418 585
R125 B.n417 B.n16 585
R126 B.n416 B.n415 585
R127 B.n414 B.n17 585
R128 B.n413 B.n412 585
R129 B.n411 B.n18 585
R130 B.n410 B.n409 585
R131 B.n408 B.n19 585
R132 B.n407 B.n406 585
R133 B.n405 B.n20 585
R134 B.n404 B.n403 585
R135 B.n402 B.n21 585
R136 B.n401 B.n400 585
R137 B.n399 B.n22 585
R138 B.n398 B.n397 585
R139 B.n396 B.n23 585
R140 B.n395 B.n394 585
R141 B.n393 B.n24 585
R142 B.n392 B.n391 585
R143 B.n390 B.n25 585
R144 B.n389 B.n388 585
R145 B.n387 B.n26 585
R146 B.n386 B.n385 585
R147 B.n384 B.n27 585
R148 B.n382 B.n381 585
R149 B.n380 B.n30 585
R150 B.n379 B.n378 585
R151 B.n377 B.n31 585
R152 B.n376 B.n375 585
R153 B.n374 B.n32 585
R154 B.n373 B.n372 585
R155 B.n371 B.n33 585
R156 B.n370 B.n369 585
R157 B.n368 B.n367 585
R158 B.n366 B.n37 585
R159 B.n365 B.n364 585
R160 B.n363 B.n38 585
R161 B.n362 B.n361 585
R162 B.n360 B.n39 585
R163 B.n359 B.n358 585
R164 B.n357 B.n40 585
R165 B.n356 B.n355 585
R166 B.n354 B.n41 585
R167 B.n353 B.n352 585
R168 B.n351 B.n42 585
R169 B.n350 B.n349 585
R170 B.n348 B.n43 585
R171 B.n347 B.n346 585
R172 B.n345 B.n44 585
R173 B.n344 B.n343 585
R174 B.n342 B.n45 585
R175 B.n341 B.n340 585
R176 B.n339 B.n46 585
R177 B.n338 B.n337 585
R178 B.n336 B.n47 585
R179 B.n335 B.n334 585
R180 B.n333 B.n48 585
R181 B.n332 B.n331 585
R182 B.n330 B.n49 585
R183 B.n329 B.n328 585
R184 B.n327 B.n50 585
R185 B.n326 B.n325 585
R186 B.n324 B.n51 585
R187 B.n323 B.n322 585
R188 B.n321 B.n52 585
R189 B.n320 B.n319 585
R190 B.n318 B.n53 585
R191 B.n317 B.n316 585
R192 B.n437 B.n436 585
R193 B.n438 B.n9 585
R194 B.n440 B.n439 585
R195 B.n441 B.n8 585
R196 B.n443 B.n442 585
R197 B.n444 B.n7 585
R198 B.n446 B.n445 585
R199 B.n447 B.n6 585
R200 B.n449 B.n448 585
R201 B.n450 B.n5 585
R202 B.n452 B.n451 585
R203 B.n453 B.n4 585
R204 B.n455 B.n454 585
R205 B.n456 B.n3 585
R206 B.n458 B.n457 585
R207 B.n459 B.n0 585
R208 B.n2 B.n1 585
R209 B.n121 B.n120 585
R210 B.n122 B.n119 585
R211 B.n124 B.n123 585
R212 B.n125 B.n118 585
R213 B.n127 B.n126 585
R214 B.n128 B.n117 585
R215 B.n130 B.n129 585
R216 B.n131 B.n116 585
R217 B.n133 B.n132 585
R218 B.n134 B.n115 585
R219 B.n136 B.n135 585
R220 B.n137 B.n114 585
R221 B.n139 B.n138 585
R222 B.n140 B.n113 585
R223 B.n142 B.n141 585
R224 B.n143 B.n142 492.5
R225 B.n266 B.n71 492.5
R226 B.n316 B.n315 492.5
R227 B.n436 B.n435 492.5
R228 B.n94 B.t9 423.627
R229 B.n208 B.t0 423.627
R230 B.n34 B.t6 423.627
R231 B.n28 B.t3 423.627
R232 B.n461 B.n460 256.663
R233 B.n460 B.n459 235.042
R234 B.n460 B.n2 235.042
R235 B.n144 B.n143 163.367
R236 B.n144 B.n111 163.367
R237 B.n148 B.n111 163.367
R238 B.n149 B.n148 163.367
R239 B.n150 B.n149 163.367
R240 B.n150 B.n109 163.367
R241 B.n154 B.n109 163.367
R242 B.n155 B.n154 163.367
R243 B.n156 B.n155 163.367
R244 B.n156 B.n107 163.367
R245 B.n160 B.n107 163.367
R246 B.n161 B.n160 163.367
R247 B.n162 B.n161 163.367
R248 B.n162 B.n105 163.367
R249 B.n166 B.n105 163.367
R250 B.n167 B.n166 163.367
R251 B.n168 B.n167 163.367
R252 B.n168 B.n103 163.367
R253 B.n172 B.n103 163.367
R254 B.n173 B.n172 163.367
R255 B.n174 B.n173 163.367
R256 B.n174 B.n101 163.367
R257 B.n178 B.n101 163.367
R258 B.n179 B.n178 163.367
R259 B.n180 B.n179 163.367
R260 B.n180 B.n99 163.367
R261 B.n184 B.n99 163.367
R262 B.n185 B.n184 163.367
R263 B.n186 B.n185 163.367
R264 B.n186 B.n97 163.367
R265 B.n190 B.n97 163.367
R266 B.n191 B.n190 163.367
R267 B.n192 B.n191 163.367
R268 B.n192 B.n93 163.367
R269 B.n197 B.n93 163.367
R270 B.n198 B.n197 163.367
R271 B.n199 B.n198 163.367
R272 B.n199 B.n91 163.367
R273 B.n203 B.n91 163.367
R274 B.n204 B.n203 163.367
R275 B.n205 B.n204 163.367
R276 B.n205 B.n89 163.367
R277 B.n212 B.n89 163.367
R278 B.n213 B.n212 163.367
R279 B.n214 B.n213 163.367
R280 B.n214 B.n87 163.367
R281 B.n218 B.n87 163.367
R282 B.n219 B.n218 163.367
R283 B.n220 B.n219 163.367
R284 B.n220 B.n85 163.367
R285 B.n224 B.n85 163.367
R286 B.n225 B.n224 163.367
R287 B.n226 B.n225 163.367
R288 B.n226 B.n83 163.367
R289 B.n230 B.n83 163.367
R290 B.n231 B.n230 163.367
R291 B.n232 B.n231 163.367
R292 B.n232 B.n81 163.367
R293 B.n236 B.n81 163.367
R294 B.n237 B.n236 163.367
R295 B.n238 B.n237 163.367
R296 B.n238 B.n79 163.367
R297 B.n242 B.n79 163.367
R298 B.n243 B.n242 163.367
R299 B.n244 B.n243 163.367
R300 B.n244 B.n77 163.367
R301 B.n248 B.n77 163.367
R302 B.n249 B.n248 163.367
R303 B.n250 B.n249 163.367
R304 B.n250 B.n75 163.367
R305 B.n254 B.n75 163.367
R306 B.n255 B.n254 163.367
R307 B.n256 B.n255 163.367
R308 B.n256 B.n73 163.367
R309 B.n260 B.n73 163.367
R310 B.n261 B.n260 163.367
R311 B.n262 B.n261 163.367
R312 B.n262 B.n71 163.367
R313 B.n315 B.n314 163.367
R314 B.n314 B.n55 163.367
R315 B.n310 B.n55 163.367
R316 B.n310 B.n309 163.367
R317 B.n309 B.n308 163.367
R318 B.n308 B.n57 163.367
R319 B.n304 B.n57 163.367
R320 B.n304 B.n303 163.367
R321 B.n303 B.n302 163.367
R322 B.n302 B.n59 163.367
R323 B.n298 B.n59 163.367
R324 B.n298 B.n297 163.367
R325 B.n297 B.n296 163.367
R326 B.n296 B.n61 163.367
R327 B.n292 B.n61 163.367
R328 B.n292 B.n291 163.367
R329 B.n291 B.n290 163.367
R330 B.n290 B.n63 163.367
R331 B.n286 B.n63 163.367
R332 B.n286 B.n285 163.367
R333 B.n285 B.n284 163.367
R334 B.n284 B.n65 163.367
R335 B.n280 B.n65 163.367
R336 B.n280 B.n279 163.367
R337 B.n279 B.n278 163.367
R338 B.n278 B.n67 163.367
R339 B.n274 B.n67 163.367
R340 B.n274 B.n273 163.367
R341 B.n273 B.n272 163.367
R342 B.n272 B.n69 163.367
R343 B.n268 B.n69 163.367
R344 B.n268 B.n267 163.367
R345 B.n267 B.n266 163.367
R346 B.n435 B.n434 163.367
R347 B.n434 B.n11 163.367
R348 B.n430 B.n11 163.367
R349 B.n430 B.n429 163.367
R350 B.n429 B.n428 163.367
R351 B.n428 B.n13 163.367
R352 B.n424 B.n13 163.367
R353 B.n424 B.n423 163.367
R354 B.n423 B.n422 163.367
R355 B.n422 B.n15 163.367
R356 B.n418 B.n15 163.367
R357 B.n418 B.n417 163.367
R358 B.n417 B.n416 163.367
R359 B.n416 B.n17 163.367
R360 B.n412 B.n17 163.367
R361 B.n412 B.n411 163.367
R362 B.n411 B.n410 163.367
R363 B.n410 B.n19 163.367
R364 B.n406 B.n19 163.367
R365 B.n406 B.n405 163.367
R366 B.n405 B.n404 163.367
R367 B.n404 B.n21 163.367
R368 B.n400 B.n21 163.367
R369 B.n400 B.n399 163.367
R370 B.n399 B.n398 163.367
R371 B.n398 B.n23 163.367
R372 B.n394 B.n23 163.367
R373 B.n394 B.n393 163.367
R374 B.n393 B.n392 163.367
R375 B.n392 B.n25 163.367
R376 B.n388 B.n25 163.367
R377 B.n388 B.n387 163.367
R378 B.n387 B.n386 163.367
R379 B.n386 B.n27 163.367
R380 B.n381 B.n27 163.367
R381 B.n381 B.n380 163.367
R382 B.n380 B.n379 163.367
R383 B.n379 B.n31 163.367
R384 B.n375 B.n31 163.367
R385 B.n375 B.n374 163.367
R386 B.n374 B.n373 163.367
R387 B.n373 B.n33 163.367
R388 B.n369 B.n33 163.367
R389 B.n369 B.n368 163.367
R390 B.n368 B.n37 163.367
R391 B.n364 B.n37 163.367
R392 B.n364 B.n363 163.367
R393 B.n363 B.n362 163.367
R394 B.n362 B.n39 163.367
R395 B.n358 B.n39 163.367
R396 B.n358 B.n357 163.367
R397 B.n357 B.n356 163.367
R398 B.n356 B.n41 163.367
R399 B.n352 B.n41 163.367
R400 B.n352 B.n351 163.367
R401 B.n351 B.n350 163.367
R402 B.n350 B.n43 163.367
R403 B.n346 B.n43 163.367
R404 B.n346 B.n345 163.367
R405 B.n345 B.n344 163.367
R406 B.n344 B.n45 163.367
R407 B.n340 B.n45 163.367
R408 B.n340 B.n339 163.367
R409 B.n339 B.n338 163.367
R410 B.n338 B.n47 163.367
R411 B.n334 B.n47 163.367
R412 B.n334 B.n333 163.367
R413 B.n333 B.n332 163.367
R414 B.n332 B.n49 163.367
R415 B.n328 B.n49 163.367
R416 B.n328 B.n327 163.367
R417 B.n327 B.n326 163.367
R418 B.n326 B.n51 163.367
R419 B.n322 B.n51 163.367
R420 B.n322 B.n321 163.367
R421 B.n321 B.n320 163.367
R422 B.n320 B.n53 163.367
R423 B.n316 B.n53 163.367
R424 B.n436 B.n9 163.367
R425 B.n440 B.n9 163.367
R426 B.n441 B.n440 163.367
R427 B.n442 B.n441 163.367
R428 B.n442 B.n7 163.367
R429 B.n446 B.n7 163.367
R430 B.n447 B.n446 163.367
R431 B.n448 B.n447 163.367
R432 B.n448 B.n5 163.367
R433 B.n452 B.n5 163.367
R434 B.n453 B.n452 163.367
R435 B.n454 B.n453 163.367
R436 B.n454 B.n3 163.367
R437 B.n458 B.n3 163.367
R438 B.n459 B.n458 163.367
R439 B.n120 B.n2 163.367
R440 B.n120 B.n119 163.367
R441 B.n124 B.n119 163.367
R442 B.n125 B.n124 163.367
R443 B.n126 B.n125 163.367
R444 B.n126 B.n117 163.367
R445 B.n130 B.n117 163.367
R446 B.n131 B.n130 163.367
R447 B.n132 B.n131 163.367
R448 B.n132 B.n115 163.367
R449 B.n136 B.n115 163.367
R450 B.n137 B.n136 163.367
R451 B.n138 B.n137 163.367
R452 B.n138 B.n113 163.367
R453 B.n142 B.n113 163.367
R454 B.n208 B.t1 138.048
R455 B.n34 B.t8 138.048
R456 B.n94 B.t10 138.037
R457 B.n28 B.t5 138.037
R458 B.n209 B.t2 111.091
R459 B.n35 B.t7 111.091
R460 B.n95 B.t11 111.079
R461 B.n29 B.t4 111.079
R462 B.n195 B.n95 59.5399
R463 B.n210 B.n209 59.5399
R464 B.n36 B.n35 59.5399
R465 B.n383 B.n29 59.5399
R466 B.n437 B.n10 32.0005
R467 B.n317 B.n54 32.0005
R468 B.n265 B.n264 32.0005
R469 B.n141 B.n112 32.0005
R470 B.n95 B.n94 26.9581
R471 B.n209 B.n208 26.9581
R472 B.n35 B.n34 26.9581
R473 B.n29 B.n28 26.9581
R474 B B.n461 18.0485
R475 B.n438 B.n437 10.6151
R476 B.n439 B.n438 10.6151
R477 B.n439 B.n8 10.6151
R478 B.n443 B.n8 10.6151
R479 B.n444 B.n443 10.6151
R480 B.n445 B.n444 10.6151
R481 B.n445 B.n6 10.6151
R482 B.n449 B.n6 10.6151
R483 B.n450 B.n449 10.6151
R484 B.n451 B.n450 10.6151
R485 B.n451 B.n4 10.6151
R486 B.n455 B.n4 10.6151
R487 B.n456 B.n455 10.6151
R488 B.n457 B.n456 10.6151
R489 B.n457 B.n0 10.6151
R490 B.n433 B.n10 10.6151
R491 B.n433 B.n432 10.6151
R492 B.n432 B.n431 10.6151
R493 B.n431 B.n12 10.6151
R494 B.n427 B.n12 10.6151
R495 B.n427 B.n426 10.6151
R496 B.n426 B.n425 10.6151
R497 B.n425 B.n14 10.6151
R498 B.n421 B.n14 10.6151
R499 B.n421 B.n420 10.6151
R500 B.n420 B.n419 10.6151
R501 B.n419 B.n16 10.6151
R502 B.n415 B.n16 10.6151
R503 B.n415 B.n414 10.6151
R504 B.n414 B.n413 10.6151
R505 B.n413 B.n18 10.6151
R506 B.n409 B.n18 10.6151
R507 B.n409 B.n408 10.6151
R508 B.n408 B.n407 10.6151
R509 B.n407 B.n20 10.6151
R510 B.n403 B.n20 10.6151
R511 B.n403 B.n402 10.6151
R512 B.n402 B.n401 10.6151
R513 B.n401 B.n22 10.6151
R514 B.n397 B.n22 10.6151
R515 B.n397 B.n396 10.6151
R516 B.n396 B.n395 10.6151
R517 B.n395 B.n24 10.6151
R518 B.n391 B.n24 10.6151
R519 B.n391 B.n390 10.6151
R520 B.n390 B.n389 10.6151
R521 B.n389 B.n26 10.6151
R522 B.n385 B.n26 10.6151
R523 B.n385 B.n384 10.6151
R524 B.n382 B.n30 10.6151
R525 B.n378 B.n30 10.6151
R526 B.n378 B.n377 10.6151
R527 B.n377 B.n376 10.6151
R528 B.n376 B.n32 10.6151
R529 B.n372 B.n32 10.6151
R530 B.n372 B.n371 10.6151
R531 B.n371 B.n370 10.6151
R532 B.n367 B.n366 10.6151
R533 B.n366 B.n365 10.6151
R534 B.n365 B.n38 10.6151
R535 B.n361 B.n38 10.6151
R536 B.n361 B.n360 10.6151
R537 B.n360 B.n359 10.6151
R538 B.n359 B.n40 10.6151
R539 B.n355 B.n40 10.6151
R540 B.n355 B.n354 10.6151
R541 B.n354 B.n353 10.6151
R542 B.n353 B.n42 10.6151
R543 B.n349 B.n42 10.6151
R544 B.n349 B.n348 10.6151
R545 B.n348 B.n347 10.6151
R546 B.n347 B.n44 10.6151
R547 B.n343 B.n44 10.6151
R548 B.n343 B.n342 10.6151
R549 B.n342 B.n341 10.6151
R550 B.n341 B.n46 10.6151
R551 B.n337 B.n46 10.6151
R552 B.n337 B.n336 10.6151
R553 B.n336 B.n335 10.6151
R554 B.n335 B.n48 10.6151
R555 B.n331 B.n48 10.6151
R556 B.n331 B.n330 10.6151
R557 B.n330 B.n329 10.6151
R558 B.n329 B.n50 10.6151
R559 B.n325 B.n50 10.6151
R560 B.n325 B.n324 10.6151
R561 B.n324 B.n323 10.6151
R562 B.n323 B.n52 10.6151
R563 B.n319 B.n52 10.6151
R564 B.n319 B.n318 10.6151
R565 B.n318 B.n317 10.6151
R566 B.n313 B.n54 10.6151
R567 B.n313 B.n312 10.6151
R568 B.n312 B.n311 10.6151
R569 B.n311 B.n56 10.6151
R570 B.n307 B.n56 10.6151
R571 B.n307 B.n306 10.6151
R572 B.n306 B.n305 10.6151
R573 B.n305 B.n58 10.6151
R574 B.n301 B.n58 10.6151
R575 B.n301 B.n300 10.6151
R576 B.n300 B.n299 10.6151
R577 B.n299 B.n60 10.6151
R578 B.n295 B.n60 10.6151
R579 B.n295 B.n294 10.6151
R580 B.n294 B.n293 10.6151
R581 B.n293 B.n62 10.6151
R582 B.n289 B.n62 10.6151
R583 B.n289 B.n288 10.6151
R584 B.n288 B.n287 10.6151
R585 B.n287 B.n64 10.6151
R586 B.n283 B.n64 10.6151
R587 B.n283 B.n282 10.6151
R588 B.n282 B.n281 10.6151
R589 B.n281 B.n66 10.6151
R590 B.n277 B.n66 10.6151
R591 B.n277 B.n276 10.6151
R592 B.n276 B.n275 10.6151
R593 B.n275 B.n68 10.6151
R594 B.n271 B.n68 10.6151
R595 B.n271 B.n270 10.6151
R596 B.n270 B.n269 10.6151
R597 B.n269 B.n70 10.6151
R598 B.n265 B.n70 10.6151
R599 B.n121 B.n1 10.6151
R600 B.n122 B.n121 10.6151
R601 B.n123 B.n122 10.6151
R602 B.n123 B.n118 10.6151
R603 B.n127 B.n118 10.6151
R604 B.n128 B.n127 10.6151
R605 B.n129 B.n128 10.6151
R606 B.n129 B.n116 10.6151
R607 B.n133 B.n116 10.6151
R608 B.n134 B.n133 10.6151
R609 B.n135 B.n134 10.6151
R610 B.n135 B.n114 10.6151
R611 B.n139 B.n114 10.6151
R612 B.n140 B.n139 10.6151
R613 B.n141 B.n140 10.6151
R614 B.n145 B.n112 10.6151
R615 B.n146 B.n145 10.6151
R616 B.n147 B.n146 10.6151
R617 B.n147 B.n110 10.6151
R618 B.n151 B.n110 10.6151
R619 B.n152 B.n151 10.6151
R620 B.n153 B.n152 10.6151
R621 B.n153 B.n108 10.6151
R622 B.n157 B.n108 10.6151
R623 B.n158 B.n157 10.6151
R624 B.n159 B.n158 10.6151
R625 B.n159 B.n106 10.6151
R626 B.n163 B.n106 10.6151
R627 B.n164 B.n163 10.6151
R628 B.n165 B.n164 10.6151
R629 B.n165 B.n104 10.6151
R630 B.n169 B.n104 10.6151
R631 B.n170 B.n169 10.6151
R632 B.n171 B.n170 10.6151
R633 B.n171 B.n102 10.6151
R634 B.n175 B.n102 10.6151
R635 B.n176 B.n175 10.6151
R636 B.n177 B.n176 10.6151
R637 B.n177 B.n100 10.6151
R638 B.n181 B.n100 10.6151
R639 B.n182 B.n181 10.6151
R640 B.n183 B.n182 10.6151
R641 B.n183 B.n98 10.6151
R642 B.n187 B.n98 10.6151
R643 B.n188 B.n187 10.6151
R644 B.n189 B.n188 10.6151
R645 B.n189 B.n96 10.6151
R646 B.n193 B.n96 10.6151
R647 B.n194 B.n193 10.6151
R648 B.n196 B.n92 10.6151
R649 B.n200 B.n92 10.6151
R650 B.n201 B.n200 10.6151
R651 B.n202 B.n201 10.6151
R652 B.n202 B.n90 10.6151
R653 B.n206 B.n90 10.6151
R654 B.n207 B.n206 10.6151
R655 B.n211 B.n207 10.6151
R656 B.n215 B.n88 10.6151
R657 B.n216 B.n215 10.6151
R658 B.n217 B.n216 10.6151
R659 B.n217 B.n86 10.6151
R660 B.n221 B.n86 10.6151
R661 B.n222 B.n221 10.6151
R662 B.n223 B.n222 10.6151
R663 B.n223 B.n84 10.6151
R664 B.n227 B.n84 10.6151
R665 B.n228 B.n227 10.6151
R666 B.n229 B.n228 10.6151
R667 B.n229 B.n82 10.6151
R668 B.n233 B.n82 10.6151
R669 B.n234 B.n233 10.6151
R670 B.n235 B.n234 10.6151
R671 B.n235 B.n80 10.6151
R672 B.n239 B.n80 10.6151
R673 B.n240 B.n239 10.6151
R674 B.n241 B.n240 10.6151
R675 B.n241 B.n78 10.6151
R676 B.n245 B.n78 10.6151
R677 B.n246 B.n245 10.6151
R678 B.n247 B.n246 10.6151
R679 B.n247 B.n76 10.6151
R680 B.n251 B.n76 10.6151
R681 B.n252 B.n251 10.6151
R682 B.n253 B.n252 10.6151
R683 B.n253 B.n74 10.6151
R684 B.n257 B.n74 10.6151
R685 B.n258 B.n257 10.6151
R686 B.n259 B.n258 10.6151
R687 B.n259 B.n72 10.6151
R688 B.n263 B.n72 10.6151
R689 B.n264 B.n263 10.6151
R690 B.n461 B.n0 8.11757
R691 B.n461 B.n1 8.11757
R692 B.n383 B.n382 7.18099
R693 B.n370 B.n36 7.18099
R694 B.n196 B.n195 7.18099
R695 B.n211 B.n210 7.18099
R696 B.n384 B.n383 3.43465
R697 B.n367 B.n36 3.43465
R698 B.n195 B.n194 3.43465
R699 B.n210 B.n88 3.43465
R700 VP.n0 VP.t0 457.735
R701 VP.n0 VP.t1 418.897
R702 VP VP.n0 0.0516364
R703 VTAIL.n1 VTAIL.t0 66.2415
R704 VTAIL.n3 VTAIL.t1 66.2414
R705 VTAIL.n0 VTAIL.t3 66.2414
R706 VTAIL.n2 VTAIL.t2 66.2414
R707 VTAIL.n1 VTAIL.n0 23.1341
R708 VTAIL.n3 VTAIL.n2 21.9358
R709 VTAIL.n2 VTAIL.n1 1.06947
R710 VTAIL VTAIL.n0 0.828086
R711 VTAIL VTAIL.n3 0.241879
R712 VDD1 VDD1.t0 118.171
R713 VDD1 VDD1.t1 83.2779
R714 VN VN.t1 458.115
R715 VN VN.t0 418.949
R716 VDD2.n0 VDD2.t1 117.347
R717 VDD2.n0 VDD2.t0 82.9201
R718 VDD2 VDD2.n0 0.358259
C0 VP VN 4.29653f
C1 VDD2 w_n1526_n2910# 1.45125f
C2 VDD1 VP 2.00081f
C3 VTAIL VN 1.52863f
C4 VDD1 VTAIL 4.5059f
C5 VDD1 VN 0.148753f
C6 VDD2 B 1.3232f
C7 w_n1526_n2910# B 6.50203f
C8 VDD2 VP 0.269664f
C9 VDD2 VTAIL 4.54445f
C10 VP w_n1526_n2910# 2.11328f
C11 VDD2 VN 1.88303f
C12 w_n1526_n2910# VTAIL 2.4958f
C13 VDD1 VDD2 0.497833f
C14 w_n1526_n2910# VN 1.92222f
C15 VDD1 w_n1526_n2910# 1.44297f
C16 VP B 1.07011f
C17 VTAIL B 2.4768f
C18 VN B 0.762169f
C19 VDD1 B 1.30611f
C20 VP VTAIL 1.54306f
C21 VDD2 VSUBS 0.677589f
C22 VDD1 VSUBS 3.7622f
C23 VTAIL VSUBS 0.715689f
C24 VN VSUBS 4.04261f
C25 VP VSUBS 1.128873f
C26 B VSUBS 2.565328f
C27 w_n1526_n2910# VSUBS 54.8811f
C28 VDD2.t1 VSUBS 1.37388f
C29 VDD2.t0 VSUBS 1.08735f
C30 VDD2.n0 VSUBS 1.99407f
C31 VN.t0 VSUBS 0.926266f
C32 VN.t1 VSUBS 1.02981f
C33 VDD1.t1 VSUBS 1.55426f
C34 VDD1.t0 VSUBS 1.98437f
C35 VTAIL.t3 VSUBS 1.70566f
C36 VTAIL.n0 VSUBS 1.82222f
C37 VTAIL.t0 VSUBS 1.70567f
C38 VTAIL.n1 VSUBS 1.84102f
C39 VTAIL.t2 VSUBS 1.70566f
C40 VTAIL.n2 VSUBS 1.74765f
C41 VTAIL.t1 VSUBS 1.70566f
C42 VTAIL.n3 VSUBS 1.68316f
C43 VP.t0 VSUBS 2.02498f
C44 VP.t1 VSUBS 1.82565f
C45 VP.n0 VSUBS 4.51875f
C46 B.n0 VSUBS 0.006579f
C47 B.n1 VSUBS 0.006579f
C48 B.n2 VSUBS 0.009731f
C49 B.n3 VSUBS 0.007457f
C50 B.n4 VSUBS 0.007457f
C51 B.n5 VSUBS 0.007457f
C52 B.n6 VSUBS 0.007457f
C53 B.n7 VSUBS 0.007457f
C54 B.n8 VSUBS 0.007457f
C55 B.n9 VSUBS 0.007457f
C56 B.n10 VSUBS 0.017359f
C57 B.n11 VSUBS 0.007457f
C58 B.n12 VSUBS 0.007457f
C59 B.n13 VSUBS 0.007457f
C60 B.n14 VSUBS 0.007457f
C61 B.n15 VSUBS 0.007457f
C62 B.n16 VSUBS 0.007457f
C63 B.n17 VSUBS 0.007457f
C64 B.n18 VSUBS 0.007457f
C65 B.n19 VSUBS 0.007457f
C66 B.n20 VSUBS 0.007457f
C67 B.n21 VSUBS 0.007457f
C68 B.n22 VSUBS 0.007457f
C69 B.n23 VSUBS 0.007457f
C70 B.n24 VSUBS 0.007457f
C71 B.n25 VSUBS 0.007457f
C72 B.n26 VSUBS 0.007457f
C73 B.n27 VSUBS 0.007457f
C74 B.t4 VSUBS 0.327817f
C75 B.t5 VSUBS 0.339308f
C76 B.t3 VSUBS 0.472626f
C77 B.n28 VSUBS 0.142244f
C78 B.n29 VSUBS 0.069475f
C79 B.n30 VSUBS 0.007457f
C80 B.n31 VSUBS 0.007457f
C81 B.n32 VSUBS 0.007457f
C82 B.n33 VSUBS 0.007457f
C83 B.t7 VSUBS 0.327813f
C84 B.t8 VSUBS 0.339303f
C85 B.t6 VSUBS 0.472626f
C86 B.n34 VSUBS 0.142248f
C87 B.n35 VSUBS 0.069479f
C88 B.n36 VSUBS 0.017276f
C89 B.n37 VSUBS 0.007457f
C90 B.n38 VSUBS 0.007457f
C91 B.n39 VSUBS 0.007457f
C92 B.n40 VSUBS 0.007457f
C93 B.n41 VSUBS 0.007457f
C94 B.n42 VSUBS 0.007457f
C95 B.n43 VSUBS 0.007457f
C96 B.n44 VSUBS 0.007457f
C97 B.n45 VSUBS 0.007457f
C98 B.n46 VSUBS 0.007457f
C99 B.n47 VSUBS 0.007457f
C100 B.n48 VSUBS 0.007457f
C101 B.n49 VSUBS 0.007457f
C102 B.n50 VSUBS 0.007457f
C103 B.n51 VSUBS 0.007457f
C104 B.n52 VSUBS 0.007457f
C105 B.n53 VSUBS 0.007457f
C106 B.n54 VSUBS 0.017073f
C107 B.n55 VSUBS 0.007457f
C108 B.n56 VSUBS 0.007457f
C109 B.n57 VSUBS 0.007457f
C110 B.n58 VSUBS 0.007457f
C111 B.n59 VSUBS 0.007457f
C112 B.n60 VSUBS 0.007457f
C113 B.n61 VSUBS 0.007457f
C114 B.n62 VSUBS 0.007457f
C115 B.n63 VSUBS 0.007457f
C116 B.n64 VSUBS 0.007457f
C117 B.n65 VSUBS 0.007457f
C118 B.n66 VSUBS 0.007457f
C119 B.n67 VSUBS 0.007457f
C120 B.n68 VSUBS 0.007457f
C121 B.n69 VSUBS 0.007457f
C122 B.n70 VSUBS 0.007457f
C123 B.n71 VSUBS 0.017359f
C124 B.n72 VSUBS 0.007457f
C125 B.n73 VSUBS 0.007457f
C126 B.n74 VSUBS 0.007457f
C127 B.n75 VSUBS 0.007457f
C128 B.n76 VSUBS 0.007457f
C129 B.n77 VSUBS 0.007457f
C130 B.n78 VSUBS 0.007457f
C131 B.n79 VSUBS 0.007457f
C132 B.n80 VSUBS 0.007457f
C133 B.n81 VSUBS 0.007457f
C134 B.n82 VSUBS 0.007457f
C135 B.n83 VSUBS 0.007457f
C136 B.n84 VSUBS 0.007457f
C137 B.n85 VSUBS 0.007457f
C138 B.n86 VSUBS 0.007457f
C139 B.n87 VSUBS 0.007457f
C140 B.n88 VSUBS 0.004935f
C141 B.n89 VSUBS 0.007457f
C142 B.n90 VSUBS 0.007457f
C143 B.n91 VSUBS 0.007457f
C144 B.n92 VSUBS 0.007457f
C145 B.n93 VSUBS 0.007457f
C146 B.t11 VSUBS 0.327817f
C147 B.t10 VSUBS 0.339308f
C148 B.t9 VSUBS 0.472626f
C149 B.n94 VSUBS 0.142244f
C150 B.n95 VSUBS 0.069475f
C151 B.n96 VSUBS 0.007457f
C152 B.n97 VSUBS 0.007457f
C153 B.n98 VSUBS 0.007457f
C154 B.n99 VSUBS 0.007457f
C155 B.n100 VSUBS 0.007457f
C156 B.n101 VSUBS 0.007457f
C157 B.n102 VSUBS 0.007457f
C158 B.n103 VSUBS 0.007457f
C159 B.n104 VSUBS 0.007457f
C160 B.n105 VSUBS 0.007457f
C161 B.n106 VSUBS 0.007457f
C162 B.n107 VSUBS 0.007457f
C163 B.n108 VSUBS 0.007457f
C164 B.n109 VSUBS 0.007457f
C165 B.n110 VSUBS 0.007457f
C166 B.n111 VSUBS 0.007457f
C167 B.n112 VSUBS 0.017359f
C168 B.n113 VSUBS 0.007457f
C169 B.n114 VSUBS 0.007457f
C170 B.n115 VSUBS 0.007457f
C171 B.n116 VSUBS 0.007457f
C172 B.n117 VSUBS 0.007457f
C173 B.n118 VSUBS 0.007457f
C174 B.n119 VSUBS 0.007457f
C175 B.n120 VSUBS 0.007457f
C176 B.n121 VSUBS 0.007457f
C177 B.n122 VSUBS 0.007457f
C178 B.n123 VSUBS 0.007457f
C179 B.n124 VSUBS 0.007457f
C180 B.n125 VSUBS 0.007457f
C181 B.n126 VSUBS 0.007457f
C182 B.n127 VSUBS 0.007457f
C183 B.n128 VSUBS 0.007457f
C184 B.n129 VSUBS 0.007457f
C185 B.n130 VSUBS 0.007457f
C186 B.n131 VSUBS 0.007457f
C187 B.n132 VSUBS 0.007457f
C188 B.n133 VSUBS 0.007457f
C189 B.n134 VSUBS 0.007457f
C190 B.n135 VSUBS 0.007457f
C191 B.n136 VSUBS 0.007457f
C192 B.n137 VSUBS 0.007457f
C193 B.n138 VSUBS 0.007457f
C194 B.n139 VSUBS 0.007457f
C195 B.n140 VSUBS 0.007457f
C196 B.n141 VSUBS 0.017073f
C197 B.n142 VSUBS 0.017073f
C198 B.n143 VSUBS 0.017359f
C199 B.n144 VSUBS 0.007457f
C200 B.n145 VSUBS 0.007457f
C201 B.n146 VSUBS 0.007457f
C202 B.n147 VSUBS 0.007457f
C203 B.n148 VSUBS 0.007457f
C204 B.n149 VSUBS 0.007457f
C205 B.n150 VSUBS 0.007457f
C206 B.n151 VSUBS 0.007457f
C207 B.n152 VSUBS 0.007457f
C208 B.n153 VSUBS 0.007457f
C209 B.n154 VSUBS 0.007457f
C210 B.n155 VSUBS 0.007457f
C211 B.n156 VSUBS 0.007457f
C212 B.n157 VSUBS 0.007457f
C213 B.n158 VSUBS 0.007457f
C214 B.n159 VSUBS 0.007457f
C215 B.n160 VSUBS 0.007457f
C216 B.n161 VSUBS 0.007457f
C217 B.n162 VSUBS 0.007457f
C218 B.n163 VSUBS 0.007457f
C219 B.n164 VSUBS 0.007457f
C220 B.n165 VSUBS 0.007457f
C221 B.n166 VSUBS 0.007457f
C222 B.n167 VSUBS 0.007457f
C223 B.n168 VSUBS 0.007457f
C224 B.n169 VSUBS 0.007457f
C225 B.n170 VSUBS 0.007457f
C226 B.n171 VSUBS 0.007457f
C227 B.n172 VSUBS 0.007457f
C228 B.n173 VSUBS 0.007457f
C229 B.n174 VSUBS 0.007457f
C230 B.n175 VSUBS 0.007457f
C231 B.n176 VSUBS 0.007457f
C232 B.n177 VSUBS 0.007457f
C233 B.n178 VSUBS 0.007457f
C234 B.n179 VSUBS 0.007457f
C235 B.n180 VSUBS 0.007457f
C236 B.n181 VSUBS 0.007457f
C237 B.n182 VSUBS 0.007457f
C238 B.n183 VSUBS 0.007457f
C239 B.n184 VSUBS 0.007457f
C240 B.n185 VSUBS 0.007457f
C241 B.n186 VSUBS 0.007457f
C242 B.n187 VSUBS 0.007457f
C243 B.n188 VSUBS 0.007457f
C244 B.n189 VSUBS 0.007457f
C245 B.n190 VSUBS 0.007457f
C246 B.n191 VSUBS 0.007457f
C247 B.n192 VSUBS 0.007457f
C248 B.n193 VSUBS 0.007457f
C249 B.n194 VSUBS 0.004935f
C250 B.n195 VSUBS 0.017276f
C251 B.n196 VSUBS 0.00625f
C252 B.n197 VSUBS 0.007457f
C253 B.n198 VSUBS 0.007457f
C254 B.n199 VSUBS 0.007457f
C255 B.n200 VSUBS 0.007457f
C256 B.n201 VSUBS 0.007457f
C257 B.n202 VSUBS 0.007457f
C258 B.n203 VSUBS 0.007457f
C259 B.n204 VSUBS 0.007457f
C260 B.n205 VSUBS 0.007457f
C261 B.n206 VSUBS 0.007457f
C262 B.n207 VSUBS 0.007457f
C263 B.t2 VSUBS 0.327813f
C264 B.t1 VSUBS 0.339303f
C265 B.t0 VSUBS 0.472626f
C266 B.n208 VSUBS 0.142248f
C267 B.n209 VSUBS 0.069479f
C268 B.n210 VSUBS 0.017276f
C269 B.n211 VSUBS 0.00625f
C270 B.n212 VSUBS 0.007457f
C271 B.n213 VSUBS 0.007457f
C272 B.n214 VSUBS 0.007457f
C273 B.n215 VSUBS 0.007457f
C274 B.n216 VSUBS 0.007457f
C275 B.n217 VSUBS 0.007457f
C276 B.n218 VSUBS 0.007457f
C277 B.n219 VSUBS 0.007457f
C278 B.n220 VSUBS 0.007457f
C279 B.n221 VSUBS 0.007457f
C280 B.n222 VSUBS 0.007457f
C281 B.n223 VSUBS 0.007457f
C282 B.n224 VSUBS 0.007457f
C283 B.n225 VSUBS 0.007457f
C284 B.n226 VSUBS 0.007457f
C285 B.n227 VSUBS 0.007457f
C286 B.n228 VSUBS 0.007457f
C287 B.n229 VSUBS 0.007457f
C288 B.n230 VSUBS 0.007457f
C289 B.n231 VSUBS 0.007457f
C290 B.n232 VSUBS 0.007457f
C291 B.n233 VSUBS 0.007457f
C292 B.n234 VSUBS 0.007457f
C293 B.n235 VSUBS 0.007457f
C294 B.n236 VSUBS 0.007457f
C295 B.n237 VSUBS 0.007457f
C296 B.n238 VSUBS 0.007457f
C297 B.n239 VSUBS 0.007457f
C298 B.n240 VSUBS 0.007457f
C299 B.n241 VSUBS 0.007457f
C300 B.n242 VSUBS 0.007457f
C301 B.n243 VSUBS 0.007457f
C302 B.n244 VSUBS 0.007457f
C303 B.n245 VSUBS 0.007457f
C304 B.n246 VSUBS 0.007457f
C305 B.n247 VSUBS 0.007457f
C306 B.n248 VSUBS 0.007457f
C307 B.n249 VSUBS 0.007457f
C308 B.n250 VSUBS 0.007457f
C309 B.n251 VSUBS 0.007457f
C310 B.n252 VSUBS 0.007457f
C311 B.n253 VSUBS 0.007457f
C312 B.n254 VSUBS 0.007457f
C313 B.n255 VSUBS 0.007457f
C314 B.n256 VSUBS 0.007457f
C315 B.n257 VSUBS 0.007457f
C316 B.n258 VSUBS 0.007457f
C317 B.n259 VSUBS 0.007457f
C318 B.n260 VSUBS 0.007457f
C319 B.n261 VSUBS 0.007457f
C320 B.n262 VSUBS 0.007457f
C321 B.n263 VSUBS 0.007457f
C322 B.n264 VSUBS 0.01646f
C323 B.n265 VSUBS 0.017973f
C324 B.n266 VSUBS 0.017073f
C325 B.n267 VSUBS 0.007457f
C326 B.n268 VSUBS 0.007457f
C327 B.n269 VSUBS 0.007457f
C328 B.n270 VSUBS 0.007457f
C329 B.n271 VSUBS 0.007457f
C330 B.n272 VSUBS 0.007457f
C331 B.n273 VSUBS 0.007457f
C332 B.n274 VSUBS 0.007457f
C333 B.n275 VSUBS 0.007457f
C334 B.n276 VSUBS 0.007457f
C335 B.n277 VSUBS 0.007457f
C336 B.n278 VSUBS 0.007457f
C337 B.n279 VSUBS 0.007457f
C338 B.n280 VSUBS 0.007457f
C339 B.n281 VSUBS 0.007457f
C340 B.n282 VSUBS 0.007457f
C341 B.n283 VSUBS 0.007457f
C342 B.n284 VSUBS 0.007457f
C343 B.n285 VSUBS 0.007457f
C344 B.n286 VSUBS 0.007457f
C345 B.n287 VSUBS 0.007457f
C346 B.n288 VSUBS 0.007457f
C347 B.n289 VSUBS 0.007457f
C348 B.n290 VSUBS 0.007457f
C349 B.n291 VSUBS 0.007457f
C350 B.n292 VSUBS 0.007457f
C351 B.n293 VSUBS 0.007457f
C352 B.n294 VSUBS 0.007457f
C353 B.n295 VSUBS 0.007457f
C354 B.n296 VSUBS 0.007457f
C355 B.n297 VSUBS 0.007457f
C356 B.n298 VSUBS 0.007457f
C357 B.n299 VSUBS 0.007457f
C358 B.n300 VSUBS 0.007457f
C359 B.n301 VSUBS 0.007457f
C360 B.n302 VSUBS 0.007457f
C361 B.n303 VSUBS 0.007457f
C362 B.n304 VSUBS 0.007457f
C363 B.n305 VSUBS 0.007457f
C364 B.n306 VSUBS 0.007457f
C365 B.n307 VSUBS 0.007457f
C366 B.n308 VSUBS 0.007457f
C367 B.n309 VSUBS 0.007457f
C368 B.n310 VSUBS 0.007457f
C369 B.n311 VSUBS 0.007457f
C370 B.n312 VSUBS 0.007457f
C371 B.n313 VSUBS 0.007457f
C372 B.n314 VSUBS 0.007457f
C373 B.n315 VSUBS 0.017073f
C374 B.n316 VSUBS 0.017359f
C375 B.n317 VSUBS 0.017359f
C376 B.n318 VSUBS 0.007457f
C377 B.n319 VSUBS 0.007457f
C378 B.n320 VSUBS 0.007457f
C379 B.n321 VSUBS 0.007457f
C380 B.n322 VSUBS 0.007457f
C381 B.n323 VSUBS 0.007457f
C382 B.n324 VSUBS 0.007457f
C383 B.n325 VSUBS 0.007457f
C384 B.n326 VSUBS 0.007457f
C385 B.n327 VSUBS 0.007457f
C386 B.n328 VSUBS 0.007457f
C387 B.n329 VSUBS 0.007457f
C388 B.n330 VSUBS 0.007457f
C389 B.n331 VSUBS 0.007457f
C390 B.n332 VSUBS 0.007457f
C391 B.n333 VSUBS 0.007457f
C392 B.n334 VSUBS 0.007457f
C393 B.n335 VSUBS 0.007457f
C394 B.n336 VSUBS 0.007457f
C395 B.n337 VSUBS 0.007457f
C396 B.n338 VSUBS 0.007457f
C397 B.n339 VSUBS 0.007457f
C398 B.n340 VSUBS 0.007457f
C399 B.n341 VSUBS 0.007457f
C400 B.n342 VSUBS 0.007457f
C401 B.n343 VSUBS 0.007457f
C402 B.n344 VSUBS 0.007457f
C403 B.n345 VSUBS 0.007457f
C404 B.n346 VSUBS 0.007457f
C405 B.n347 VSUBS 0.007457f
C406 B.n348 VSUBS 0.007457f
C407 B.n349 VSUBS 0.007457f
C408 B.n350 VSUBS 0.007457f
C409 B.n351 VSUBS 0.007457f
C410 B.n352 VSUBS 0.007457f
C411 B.n353 VSUBS 0.007457f
C412 B.n354 VSUBS 0.007457f
C413 B.n355 VSUBS 0.007457f
C414 B.n356 VSUBS 0.007457f
C415 B.n357 VSUBS 0.007457f
C416 B.n358 VSUBS 0.007457f
C417 B.n359 VSUBS 0.007457f
C418 B.n360 VSUBS 0.007457f
C419 B.n361 VSUBS 0.007457f
C420 B.n362 VSUBS 0.007457f
C421 B.n363 VSUBS 0.007457f
C422 B.n364 VSUBS 0.007457f
C423 B.n365 VSUBS 0.007457f
C424 B.n366 VSUBS 0.007457f
C425 B.n367 VSUBS 0.004935f
C426 B.n368 VSUBS 0.007457f
C427 B.n369 VSUBS 0.007457f
C428 B.n370 VSUBS 0.00625f
C429 B.n371 VSUBS 0.007457f
C430 B.n372 VSUBS 0.007457f
C431 B.n373 VSUBS 0.007457f
C432 B.n374 VSUBS 0.007457f
C433 B.n375 VSUBS 0.007457f
C434 B.n376 VSUBS 0.007457f
C435 B.n377 VSUBS 0.007457f
C436 B.n378 VSUBS 0.007457f
C437 B.n379 VSUBS 0.007457f
C438 B.n380 VSUBS 0.007457f
C439 B.n381 VSUBS 0.007457f
C440 B.n382 VSUBS 0.00625f
C441 B.n383 VSUBS 0.017276f
C442 B.n384 VSUBS 0.004935f
C443 B.n385 VSUBS 0.007457f
C444 B.n386 VSUBS 0.007457f
C445 B.n387 VSUBS 0.007457f
C446 B.n388 VSUBS 0.007457f
C447 B.n389 VSUBS 0.007457f
C448 B.n390 VSUBS 0.007457f
C449 B.n391 VSUBS 0.007457f
C450 B.n392 VSUBS 0.007457f
C451 B.n393 VSUBS 0.007457f
C452 B.n394 VSUBS 0.007457f
C453 B.n395 VSUBS 0.007457f
C454 B.n396 VSUBS 0.007457f
C455 B.n397 VSUBS 0.007457f
C456 B.n398 VSUBS 0.007457f
C457 B.n399 VSUBS 0.007457f
C458 B.n400 VSUBS 0.007457f
C459 B.n401 VSUBS 0.007457f
C460 B.n402 VSUBS 0.007457f
C461 B.n403 VSUBS 0.007457f
C462 B.n404 VSUBS 0.007457f
C463 B.n405 VSUBS 0.007457f
C464 B.n406 VSUBS 0.007457f
C465 B.n407 VSUBS 0.007457f
C466 B.n408 VSUBS 0.007457f
C467 B.n409 VSUBS 0.007457f
C468 B.n410 VSUBS 0.007457f
C469 B.n411 VSUBS 0.007457f
C470 B.n412 VSUBS 0.007457f
C471 B.n413 VSUBS 0.007457f
C472 B.n414 VSUBS 0.007457f
C473 B.n415 VSUBS 0.007457f
C474 B.n416 VSUBS 0.007457f
C475 B.n417 VSUBS 0.007457f
C476 B.n418 VSUBS 0.007457f
C477 B.n419 VSUBS 0.007457f
C478 B.n420 VSUBS 0.007457f
C479 B.n421 VSUBS 0.007457f
C480 B.n422 VSUBS 0.007457f
C481 B.n423 VSUBS 0.007457f
C482 B.n424 VSUBS 0.007457f
C483 B.n425 VSUBS 0.007457f
C484 B.n426 VSUBS 0.007457f
C485 B.n427 VSUBS 0.007457f
C486 B.n428 VSUBS 0.007457f
C487 B.n429 VSUBS 0.007457f
C488 B.n430 VSUBS 0.007457f
C489 B.n431 VSUBS 0.007457f
C490 B.n432 VSUBS 0.007457f
C491 B.n433 VSUBS 0.007457f
C492 B.n434 VSUBS 0.007457f
C493 B.n435 VSUBS 0.017359f
C494 B.n436 VSUBS 0.017073f
C495 B.n437 VSUBS 0.017073f
C496 B.n438 VSUBS 0.007457f
C497 B.n439 VSUBS 0.007457f
C498 B.n440 VSUBS 0.007457f
C499 B.n441 VSUBS 0.007457f
C500 B.n442 VSUBS 0.007457f
C501 B.n443 VSUBS 0.007457f
C502 B.n444 VSUBS 0.007457f
C503 B.n445 VSUBS 0.007457f
C504 B.n446 VSUBS 0.007457f
C505 B.n447 VSUBS 0.007457f
C506 B.n448 VSUBS 0.007457f
C507 B.n449 VSUBS 0.007457f
C508 B.n450 VSUBS 0.007457f
C509 B.n451 VSUBS 0.007457f
C510 B.n452 VSUBS 0.007457f
C511 B.n453 VSUBS 0.007457f
C512 B.n454 VSUBS 0.007457f
C513 B.n455 VSUBS 0.007457f
C514 B.n456 VSUBS 0.007457f
C515 B.n457 VSUBS 0.007457f
C516 B.n458 VSUBS 0.007457f
C517 B.n459 VSUBS 0.009731f
C518 B.n460 VSUBS 0.010366f
C519 B.n461 VSUBS 0.020613f
.ends

