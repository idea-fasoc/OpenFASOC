* NGSPICE file created from diff_pair_sample_0927.ext - technology: sky130A

.subckt diff_pair_sample_0927 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t14 B.t6 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X1 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=0 ps=0 w=8.47 l=1.41
X2 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=0 ps=0 w=8.47 l=1.41
X3 VDD1.t7 VP.t0 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=3.3033 ps=17.72 w=8.47 l=1.41
X4 VTAIL.t15 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X5 VTAIL.t2 VP.t1 VDD1.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X6 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=0 ps=0 w=8.47 l=1.41
X7 VTAIL.t9 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=1.39755 ps=8.8 w=8.47 l=1.41
X8 VTAIL.t7 VP.t2 VDD1.t5 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=1.39755 ps=8.8 w=8.47 l=1.41
X9 VTAIL.t5 VP.t3 VDD1.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X10 VDD2.t4 VN.t3 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=3.3033 ps=17.72 w=8.47 l=1.41
X11 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=0 ps=0 w=8.47 l=1.41
X12 VTAIL.t10 VN.t4 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X13 VTAIL.t1 VP.t4 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=1.39755 ps=8.8 w=8.47 l=1.41
X14 VDD2.t2 VN.t5 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=3.3033 ps=17.72 w=8.47 l=1.41
X15 VDD1.t2 VP.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X16 VDD2.t1 VN.t6 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X17 VTAIL.t8 VN.t7 VDD2.t0 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3033 pd=17.72 as=1.39755 ps=8.8 w=8.47 l=1.41
X18 VDD1.t1 VP.t6 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=1.39755 ps=8.8 w=8.47 l=1.41
X19 VDD1.t0 VP.t7 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.39755 pd=8.8 as=3.3033 ps=17.72 w=8.47 l=1.41
R0 VN.n18 VN.n17 180.385
R1 VN.n37 VN.n36 180.385
R2 VN.n5 VN.t7 176.014
R3 VN.n24 VN.t3 176.014
R4 VN.n35 VN.n19 161.3
R5 VN.n34 VN.n33 161.3
R6 VN.n32 VN.n20 161.3
R7 VN.n31 VN.n30 161.3
R8 VN.n28 VN.n21 161.3
R9 VN.n27 VN.n26 161.3
R10 VN.n25 VN.n22 161.3
R11 VN.n16 VN.n0 161.3
R12 VN.n15 VN.n14 161.3
R13 VN.n13 VN.n1 161.3
R14 VN.n12 VN.n11 161.3
R15 VN.n9 VN.n2 161.3
R16 VN.n8 VN.n7 161.3
R17 VN.n6 VN.n3 161.3
R18 VN.n4 VN.t0 144.772
R19 VN.n10 VN.t4 144.772
R20 VN.n17 VN.t5 144.772
R21 VN.n23 VN.t1 144.772
R22 VN.n29 VN.t6 144.772
R23 VN.n36 VN.t2 144.772
R24 VN.n15 VN.n1 56.5193
R25 VN.n34 VN.n20 56.5193
R26 VN.n5 VN.n4 47.8106
R27 VN.n24 VN.n23 47.8106
R28 VN VN.n37 42.866
R29 VN.n8 VN.n3 40.4934
R30 VN.n9 VN.n8 40.4934
R31 VN.n27 VN.n22 40.4934
R32 VN.n28 VN.n27 40.4934
R33 VN.n11 VN.n1 24.4675
R34 VN.n16 VN.n15 24.4675
R35 VN.n30 VN.n20 24.4675
R36 VN.n35 VN.n34 24.4675
R37 VN.n25 VN.n24 18.2406
R38 VN.n6 VN.n5 18.2406
R39 VN.n4 VN.n3 18.1061
R40 VN.n10 VN.n9 18.1061
R41 VN.n23 VN.n22 18.1061
R42 VN.n29 VN.n28 18.1061
R43 VN.n11 VN.n10 6.36192
R44 VN.n30 VN.n29 6.36192
R45 VN.n17 VN.n16 5.38324
R46 VN.n36 VN.n35 5.38324
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n26 VN.n21 0.189894
R53 VN.n26 VN.n25 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VTAIL.n11 VTAIL.t7 48.8952
R63 VTAIL.n10 VTAIL.t12 48.8952
R64 VTAIL.n7 VTAIL.t9 48.8952
R65 VTAIL.n14 VTAIL.t4 48.8952
R66 VTAIL.n15 VTAIL.t13 48.895
R67 VTAIL.n2 VTAIL.t8 48.895
R68 VTAIL.n3 VTAIL.t0 48.895
R69 VTAIL.n6 VTAIL.t1 48.895
R70 VTAIL.n13 VTAIL.n12 46.5576
R71 VTAIL.n9 VTAIL.n8 46.5576
R72 VTAIL.n1 VTAIL.n0 46.5575
R73 VTAIL.n5 VTAIL.n4 46.5575
R74 VTAIL.n15 VTAIL.n14 21.1686
R75 VTAIL.n7 VTAIL.n6 21.1686
R76 VTAIL.n0 VTAIL.t14 2.33816
R77 VTAIL.n0 VTAIL.t10 2.33816
R78 VTAIL.n4 VTAIL.t3 2.33816
R79 VTAIL.n4 VTAIL.t2 2.33816
R80 VTAIL.n12 VTAIL.t6 2.33816
R81 VTAIL.n12 VTAIL.t5 2.33816
R82 VTAIL.n8 VTAIL.t11 2.33816
R83 VTAIL.n8 VTAIL.t15 2.33816
R84 VTAIL.n9 VTAIL.n7 1.5005
R85 VTAIL.n10 VTAIL.n9 1.5005
R86 VTAIL.n13 VTAIL.n11 1.5005
R87 VTAIL.n14 VTAIL.n13 1.5005
R88 VTAIL.n6 VTAIL.n5 1.5005
R89 VTAIL.n5 VTAIL.n3 1.5005
R90 VTAIL.n2 VTAIL.n1 1.5005
R91 VTAIL VTAIL.n15 1.44231
R92 VTAIL.n11 VTAIL.n10 0.470328
R93 VTAIL.n3 VTAIL.n2 0.470328
R94 VTAIL VTAIL.n1 0.0586897
R95 VDD2.n2 VDD2.n1 63.931
R96 VDD2.n2 VDD2.n0 63.931
R97 VDD2 VDD2.n5 63.9282
R98 VDD2.n4 VDD2.n3 63.2364
R99 VDD2.n4 VDD2.n2 37.767
R100 VDD2.n5 VDD2.t6 2.33816
R101 VDD2.n5 VDD2.t4 2.33816
R102 VDD2.n3 VDD2.t5 2.33816
R103 VDD2.n3 VDD2.t1 2.33816
R104 VDD2.n1 VDD2.t3 2.33816
R105 VDD2.n1 VDD2.t2 2.33816
R106 VDD2.n0 VDD2.t0 2.33816
R107 VDD2.n0 VDD2.t7 2.33816
R108 VDD2 VDD2.n4 0.80869
R109 B.n640 B.n639 585
R110 B.n245 B.n98 585
R111 B.n244 B.n243 585
R112 B.n242 B.n241 585
R113 B.n240 B.n239 585
R114 B.n238 B.n237 585
R115 B.n236 B.n235 585
R116 B.n234 B.n233 585
R117 B.n232 B.n231 585
R118 B.n230 B.n229 585
R119 B.n228 B.n227 585
R120 B.n226 B.n225 585
R121 B.n224 B.n223 585
R122 B.n222 B.n221 585
R123 B.n220 B.n219 585
R124 B.n218 B.n217 585
R125 B.n216 B.n215 585
R126 B.n214 B.n213 585
R127 B.n212 B.n211 585
R128 B.n210 B.n209 585
R129 B.n208 B.n207 585
R130 B.n206 B.n205 585
R131 B.n204 B.n203 585
R132 B.n202 B.n201 585
R133 B.n200 B.n199 585
R134 B.n198 B.n197 585
R135 B.n196 B.n195 585
R136 B.n194 B.n193 585
R137 B.n192 B.n191 585
R138 B.n190 B.n189 585
R139 B.n188 B.n187 585
R140 B.n185 B.n184 585
R141 B.n183 B.n182 585
R142 B.n181 B.n180 585
R143 B.n179 B.n178 585
R144 B.n177 B.n176 585
R145 B.n175 B.n174 585
R146 B.n173 B.n172 585
R147 B.n171 B.n170 585
R148 B.n169 B.n168 585
R149 B.n167 B.n166 585
R150 B.n164 B.n163 585
R151 B.n162 B.n161 585
R152 B.n160 B.n159 585
R153 B.n158 B.n157 585
R154 B.n156 B.n155 585
R155 B.n154 B.n153 585
R156 B.n152 B.n151 585
R157 B.n150 B.n149 585
R158 B.n148 B.n147 585
R159 B.n146 B.n145 585
R160 B.n144 B.n143 585
R161 B.n142 B.n141 585
R162 B.n140 B.n139 585
R163 B.n138 B.n137 585
R164 B.n136 B.n135 585
R165 B.n134 B.n133 585
R166 B.n132 B.n131 585
R167 B.n130 B.n129 585
R168 B.n128 B.n127 585
R169 B.n126 B.n125 585
R170 B.n124 B.n123 585
R171 B.n122 B.n121 585
R172 B.n120 B.n119 585
R173 B.n118 B.n117 585
R174 B.n116 B.n115 585
R175 B.n114 B.n113 585
R176 B.n112 B.n111 585
R177 B.n110 B.n109 585
R178 B.n108 B.n107 585
R179 B.n106 B.n105 585
R180 B.n104 B.n103 585
R181 B.n638 B.n62 585
R182 B.n643 B.n62 585
R183 B.n637 B.n61 585
R184 B.n644 B.n61 585
R185 B.n636 B.n635 585
R186 B.n635 B.n57 585
R187 B.n634 B.n56 585
R188 B.n650 B.n56 585
R189 B.n633 B.n55 585
R190 B.n651 B.n55 585
R191 B.n632 B.n54 585
R192 B.n652 B.n54 585
R193 B.n631 B.n630 585
R194 B.n630 B.n50 585
R195 B.n629 B.n49 585
R196 B.n658 B.n49 585
R197 B.n628 B.n48 585
R198 B.n659 B.n48 585
R199 B.n627 B.n47 585
R200 B.n660 B.n47 585
R201 B.n626 B.n625 585
R202 B.n625 B.n43 585
R203 B.n624 B.n42 585
R204 B.n666 B.n42 585
R205 B.n623 B.n41 585
R206 B.n667 B.n41 585
R207 B.n622 B.n40 585
R208 B.n668 B.n40 585
R209 B.n621 B.n620 585
R210 B.n620 B.n36 585
R211 B.n619 B.n35 585
R212 B.n674 B.n35 585
R213 B.n618 B.n34 585
R214 B.n675 B.n34 585
R215 B.n617 B.n33 585
R216 B.n676 B.n33 585
R217 B.n616 B.n615 585
R218 B.n615 B.n29 585
R219 B.n614 B.n28 585
R220 B.n682 B.n28 585
R221 B.n613 B.n27 585
R222 B.n683 B.n27 585
R223 B.n612 B.n26 585
R224 B.n684 B.n26 585
R225 B.n611 B.n610 585
R226 B.n610 B.n22 585
R227 B.n609 B.n21 585
R228 B.n690 B.n21 585
R229 B.n608 B.n20 585
R230 B.n691 B.n20 585
R231 B.n607 B.n19 585
R232 B.n692 B.n19 585
R233 B.n606 B.n605 585
R234 B.n605 B.n15 585
R235 B.n604 B.n14 585
R236 B.n698 B.n14 585
R237 B.n603 B.n13 585
R238 B.n699 B.n13 585
R239 B.n602 B.n12 585
R240 B.n700 B.n12 585
R241 B.n601 B.n600 585
R242 B.n600 B.n599 585
R243 B.n598 B.n597 585
R244 B.n598 B.n8 585
R245 B.n596 B.n7 585
R246 B.n707 B.n7 585
R247 B.n595 B.n6 585
R248 B.n708 B.n6 585
R249 B.n594 B.n5 585
R250 B.n709 B.n5 585
R251 B.n593 B.n592 585
R252 B.n592 B.n4 585
R253 B.n591 B.n246 585
R254 B.n591 B.n590 585
R255 B.n581 B.n247 585
R256 B.n248 B.n247 585
R257 B.n583 B.n582 585
R258 B.n584 B.n583 585
R259 B.n580 B.n253 585
R260 B.n253 B.n252 585
R261 B.n579 B.n578 585
R262 B.n578 B.n577 585
R263 B.n255 B.n254 585
R264 B.n256 B.n255 585
R265 B.n570 B.n569 585
R266 B.n571 B.n570 585
R267 B.n568 B.n260 585
R268 B.n264 B.n260 585
R269 B.n567 B.n566 585
R270 B.n566 B.n565 585
R271 B.n262 B.n261 585
R272 B.n263 B.n262 585
R273 B.n558 B.n557 585
R274 B.n559 B.n558 585
R275 B.n556 B.n269 585
R276 B.n269 B.n268 585
R277 B.n555 B.n554 585
R278 B.n554 B.n553 585
R279 B.n271 B.n270 585
R280 B.n272 B.n271 585
R281 B.n546 B.n545 585
R282 B.n547 B.n546 585
R283 B.n544 B.n277 585
R284 B.n277 B.n276 585
R285 B.n543 B.n542 585
R286 B.n542 B.n541 585
R287 B.n279 B.n278 585
R288 B.n280 B.n279 585
R289 B.n534 B.n533 585
R290 B.n535 B.n534 585
R291 B.n532 B.n285 585
R292 B.n285 B.n284 585
R293 B.n531 B.n530 585
R294 B.n530 B.n529 585
R295 B.n287 B.n286 585
R296 B.n288 B.n287 585
R297 B.n522 B.n521 585
R298 B.n523 B.n522 585
R299 B.n520 B.n293 585
R300 B.n293 B.n292 585
R301 B.n519 B.n518 585
R302 B.n518 B.n517 585
R303 B.n295 B.n294 585
R304 B.n296 B.n295 585
R305 B.n510 B.n509 585
R306 B.n511 B.n510 585
R307 B.n508 B.n301 585
R308 B.n301 B.n300 585
R309 B.n507 B.n506 585
R310 B.n506 B.n505 585
R311 B.n303 B.n302 585
R312 B.n304 B.n303 585
R313 B.n498 B.n497 585
R314 B.n499 B.n498 585
R315 B.n496 B.n309 585
R316 B.n309 B.n308 585
R317 B.n491 B.n490 585
R318 B.n489 B.n347 585
R319 B.n488 B.n346 585
R320 B.n493 B.n346 585
R321 B.n487 B.n486 585
R322 B.n485 B.n484 585
R323 B.n483 B.n482 585
R324 B.n481 B.n480 585
R325 B.n479 B.n478 585
R326 B.n477 B.n476 585
R327 B.n475 B.n474 585
R328 B.n473 B.n472 585
R329 B.n471 B.n470 585
R330 B.n469 B.n468 585
R331 B.n467 B.n466 585
R332 B.n465 B.n464 585
R333 B.n463 B.n462 585
R334 B.n461 B.n460 585
R335 B.n459 B.n458 585
R336 B.n457 B.n456 585
R337 B.n455 B.n454 585
R338 B.n453 B.n452 585
R339 B.n451 B.n450 585
R340 B.n449 B.n448 585
R341 B.n447 B.n446 585
R342 B.n445 B.n444 585
R343 B.n443 B.n442 585
R344 B.n441 B.n440 585
R345 B.n439 B.n438 585
R346 B.n437 B.n436 585
R347 B.n435 B.n434 585
R348 B.n433 B.n432 585
R349 B.n431 B.n430 585
R350 B.n429 B.n428 585
R351 B.n427 B.n426 585
R352 B.n425 B.n424 585
R353 B.n423 B.n422 585
R354 B.n421 B.n420 585
R355 B.n419 B.n418 585
R356 B.n417 B.n416 585
R357 B.n415 B.n414 585
R358 B.n413 B.n412 585
R359 B.n411 B.n410 585
R360 B.n409 B.n408 585
R361 B.n407 B.n406 585
R362 B.n405 B.n404 585
R363 B.n403 B.n402 585
R364 B.n401 B.n400 585
R365 B.n399 B.n398 585
R366 B.n397 B.n396 585
R367 B.n395 B.n394 585
R368 B.n393 B.n392 585
R369 B.n391 B.n390 585
R370 B.n389 B.n388 585
R371 B.n387 B.n386 585
R372 B.n385 B.n384 585
R373 B.n383 B.n382 585
R374 B.n381 B.n380 585
R375 B.n379 B.n378 585
R376 B.n377 B.n376 585
R377 B.n375 B.n374 585
R378 B.n373 B.n372 585
R379 B.n371 B.n370 585
R380 B.n369 B.n368 585
R381 B.n367 B.n366 585
R382 B.n365 B.n364 585
R383 B.n363 B.n362 585
R384 B.n361 B.n360 585
R385 B.n359 B.n358 585
R386 B.n357 B.n356 585
R387 B.n355 B.n354 585
R388 B.n311 B.n310 585
R389 B.n495 B.n494 585
R390 B.n494 B.n493 585
R391 B.n307 B.n306 585
R392 B.n308 B.n307 585
R393 B.n501 B.n500 585
R394 B.n500 B.n499 585
R395 B.n502 B.n305 585
R396 B.n305 B.n304 585
R397 B.n504 B.n503 585
R398 B.n505 B.n504 585
R399 B.n299 B.n298 585
R400 B.n300 B.n299 585
R401 B.n513 B.n512 585
R402 B.n512 B.n511 585
R403 B.n514 B.n297 585
R404 B.n297 B.n296 585
R405 B.n516 B.n515 585
R406 B.n517 B.n516 585
R407 B.n291 B.n290 585
R408 B.n292 B.n291 585
R409 B.n525 B.n524 585
R410 B.n524 B.n523 585
R411 B.n526 B.n289 585
R412 B.n289 B.n288 585
R413 B.n528 B.n527 585
R414 B.n529 B.n528 585
R415 B.n283 B.n282 585
R416 B.n284 B.n283 585
R417 B.n537 B.n536 585
R418 B.n536 B.n535 585
R419 B.n538 B.n281 585
R420 B.n281 B.n280 585
R421 B.n540 B.n539 585
R422 B.n541 B.n540 585
R423 B.n275 B.n274 585
R424 B.n276 B.n275 585
R425 B.n549 B.n548 585
R426 B.n548 B.n547 585
R427 B.n550 B.n273 585
R428 B.n273 B.n272 585
R429 B.n552 B.n551 585
R430 B.n553 B.n552 585
R431 B.n267 B.n266 585
R432 B.n268 B.n267 585
R433 B.n561 B.n560 585
R434 B.n560 B.n559 585
R435 B.n562 B.n265 585
R436 B.n265 B.n263 585
R437 B.n564 B.n563 585
R438 B.n565 B.n564 585
R439 B.n259 B.n258 585
R440 B.n264 B.n259 585
R441 B.n573 B.n572 585
R442 B.n572 B.n571 585
R443 B.n574 B.n257 585
R444 B.n257 B.n256 585
R445 B.n576 B.n575 585
R446 B.n577 B.n576 585
R447 B.n251 B.n250 585
R448 B.n252 B.n251 585
R449 B.n586 B.n585 585
R450 B.n585 B.n584 585
R451 B.n587 B.n249 585
R452 B.n249 B.n248 585
R453 B.n589 B.n588 585
R454 B.n590 B.n589 585
R455 B.n3 B.n0 585
R456 B.n4 B.n3 585
R457 B.n706 B.n1 585
R458 B.n707 B.n706 585
R459 B.n705 B.n704 585
R460 B.n705 B.n8 585
R461 B.n703 B.n9 585
R462 B.n599 B.n9 585
R463 B.n702 B.n701 585
R464 B.n701 B.n700 585
R465 B.n11 B.n10 585
R466 B.n699 B.n11 585
R467 B.n697 B.n696 585
R468 B.n698 B.n697 585
R469 B.n695 B.n16 585
R470 B.n16 B.n15 585
R471 B.n694 B.n693 585
R472 B.n693 B.n692 585
R473 B.n18 B.n17 585
R474 B.n691 B.n18 585
R475 B.n689 B.n688 585
R476 B.n690 B.n689 585
R477 B.n687 B.n23 585
R478 B.n23 B.n22 585
R479 B.n686 B.n685 585
R480 B.n685 B.n684 585
R481 B.n25 B.n24 585
R482 B.n683 B.n25 585
R483 B.n681 B.n680 585
R484 B.n682 B.n681 585
R485 B.n679 B.n30 585
R486 B.n30 B.n29 585
R487 B.n678 B.n677 585
R488 B.n677 B.n676 585
R489 B.n32 B.n31 585
R490 B.n675 B.n32 585
R491 B.n673 B.n672 585
R492 B.n674 B.n673 585
R493 B.n671 B.n37 585
R494 B.n37 B.n36 585
R495 B.n670 B.n669 585
R496 B.n669 B.n668 585
R497 B.n39 B.n38 585
R498 B.n667 B.n39 585
R499 B.n665 B.n664 585
R500 B.n666 B.n665 585
R501 B.n663 B.n44 585
R502 B.n44 B.n43 585
R503 B.n662 B.n661 585
R504 B.n661 B.n660 585
R505 B.n46 B.n45 585
R506 B.n659 B.n46 585
R507 B.n657 B.n656 585
R508 B.n658 B.n657 585
R509 B.n655 B.n51 585
R510 B.n51 B.n50 585
R511 B.n654 B.n653 585
R512 B.n653 B.n652 585
R513 B.n53 B.n52 585
R514 B.n651 B.n53 585
R515 B.n649 B.n648 585
R516 B.n650 B.n649 585
R517 B.n647 B.n58 585
R518 B.n58 B.n57 585
R519 B.n646 B.n645 585
R520 B.n645 B.n644 585
R521 B.n60 B.n59 585
R522 B.n643 B.n60 585
R523 B.n710 B.n709 585
R524 B.n708 B.n2 585
R525 B.n103 B.n60 535.745
R526 B.n640 B.n62 535.745
R527 B.n494 B.n309 535.745
R528 B.n491 B.n307 535.745
R529 B.n101 B.t15 349.86
R530 B.n99 B.t19 349.86
R531 B.n351 B.t12 349.86
R532 B.n348 B.t8 349.86
R533 B.n642 B.n641 256.663
R534 B.n642 B.n97 256.663
R535 B.n642 B.n96 256.663
R536 B.n642 B.n95 256.663
R537 B.n642 B.n94 256.663
R538 B.n642 B.n93 256.663
R539 B.n642 B.n92 256.663
R540 B.n642 B.n91 256.663
R541 B.n642 B.n90 256.663
R542 B.n642 B.n89 256.663
R543 B.n642 B.n88 256.663
R544 B.n642 B.n87 256.663
R545 B.n642 B.n86 256.663
R546 B.n642 B.n85 256.663
R547 B.n642 B.n84 256.663
R548 B.n642 B.n83 256.663
R549 B.n642 B.n82 256.663
R550 B.n642 B.n81 256.663
R551 B.n642 B.n80 256.663
R552 B.n642 B.n79 256.663
R553 B.n642 B.n78 256.663
R554 B.n642 B.n77 256.663
R555 B.n642 B.n76 256.663
R556 B.n642 B.n75 256.663
R557 B.n642 B.n74 256.663
R558 B.n642 B.n73 256.663
R559 B.n642 B.n72 256.663
R560 B.n642 B.n71 256.663
R561 B.n642 B.n70 256.663
R562 B.n642 B.n69 256.663
R563 B.n642 B.n68 256.663
R564 B.n642 B.n67 256.663
R565 B.n642 B.n66 256.663
R566 B.n642 B.n65 256.663
R567 B.n642 B.n64 256.663
R568 B.n642 B.n63 256.663
R569 B.n493 B.n492 256.663
R570 B.n493 B.n312 256.663
R571 B.n493 B.n313 256.663
R572 B.n493 B.n314 256.663
R573 B.n493 B.n315 256.663
R574 B.n493 B.n316 256.663
R575 B.n493 B.n317 256.663
R576 B.n493 B.n318 256.663
R577 B.n493 B.n319 256.663
R578 B.n493 B.n320 256.663
R579 B.n493 B.n321 256.663
R580 B.n493 B.n322 256.663
R581 B.n493 B.n323 256.663
R582 B.n493 B.n324 256.663
R583 B.n493 B.n325 256.663
R584 B.n493 B.n326 256.663
R585 B.n493 B.n327 256.663
R586 B.n493 B.n328 256.663
R587 B.n493 B.n329 256.663
R588 B.n493 B.n330 256.663
R589 B.n493 B.n331 256.663
R590 B.n493 B.n332 256.663
R591 B.n493 B.n333 256.663
R592 B.n493 B.n334 256.663
R593 B.n493 B.n335 256.663
R594 B.n493 B.n336 256.663
R595 B.n493 B.n337 256.663
R596 B.n493 B.n338 256.663
R597 B.n493 B.n339 256.663
R598 B.n493 B.n340 256.663
R599 B.n493 B.n341 256.663
R600 B.n493 B.n342 256.663
R601 B.n493 B.n343 256.663
R602 B.n493 B.n344 256.663
R603 B.n493 B.n345 256.663
R604 B.n712 B.n711 256.663
R605 B.n107 B.n106 163.367
R606 B.n111 B.n110 163.367
R607 B.n115 B.n114 163.367
R608 B.n119 B.n118 163.367
R609 B.n123 B.n122 163.367
R610 B.n127 B.n126 163.367
R611 B.n131 B.n130 163.367
R612 B.n135 B.n134 163.367
R613 B.n139 B.n138 163.367
R614 B.n143 B.n142 163.367
R615 B.n147 B.n146 163.367
R616 B.n151 B.n150 163.367
R617 B.n155 B.n154 163.367
R618 B.n159 B.n158 163.367
R619 B.n163 B.n162 163.367
R620 B.n168 B.n167 163.367
R621 B.n172 B.n171 163.367
R622 B.n176 B.n175 163.367
R623 B.n180 B.n179 163.367
R624 B.n184 B.n183 163.367
R625 B.n189 B.n188 163.367
R626 B.n193 B.n192 163.367
R627 B.n197 B.n196 163.367
R628 B.n201 B.n200 163.367
R629 B.n205 B.n204 163.367
R630 B.n209 B.n208 163.367
R631 B.n213 B.n212 163.367
R632 B.n217 B.n216 163.367
R633 B.n221 B.n220 163.367
R634 B.n225 B.n224 163.367
R635 B.n229 B.n228 163.367
R636 B.n233 B.n232 163.367
R637 B.n237 B.n236 163.367
R638 B.n241 B.n240 163.367
R639 B.n243 B.n98 163.367
R640 B.n498 B.n309 163.367
R641 B.n498 B.n303 163.367
R642 B.n506 B.n303 163.367
R643 B.n506 B.n301 163.367
R644 B.n510 B.n301 163.367
R645 B.n510 B.n295 163.367
R646 B.n518 B.n295 163.367
R647 B.n518 B.n293 163.367
R648 B.n522 B.n293 163.367
R649 B.n522 B.n287 163.367
R650 B.n530 B.n287 163.367
R651 B.n530 B.n285 163.367
R652 B.n534 B.n285 163.367
R653 B.n534 B.n279 163.367
R654 B.n542 B.n279 163.367
R655 B.n542 B.n277 163.367
R656 B.n546 B.n277 163.367
R657 B.n546 B.n271 163.367
R658 B.n554 B.n271 163.367
R659 B.n554 B.n269 163.367
R660 B.n558 B.n269 163.367
R661 B.n558 B.n262 163.367
R662 B.n566 B.n262 163.367
R663 B.n566 B.n260 163.367
R664 B.n570 B.n260 163.367
R665 B.n570 B.n255 163.367
R666 B.n578 B.n255 163.367
R667 B.n578 B.n253 163.367
R668 B.n583 B.n253 163.367
R669 B.n583 B.n247 163.367
R670 B.n591 B.n247 163.367
R671 B.n592 B.n591 163.367
R672 B.n592 B.n5 163.367
R673 B.n6 B.n5 163.367
R674 B.n7 B.n6 163.367
R675 B.n598 B.n7 163.367
R676 B.n600 B.n598 163.367
R677 B.n600 B.n12 163.367
R678 B.n13 B.n12 163.367
R679 B.n14 B.n13 163.367
R680 B.n605 B.n14 163.367
R681 B.n605 B.n19 163.367
R682 B.n20 B.n19 163.367
R683 B.n21 B.n20 163.367
R684 B.n610 B.n21 163.367
R685 B.n610 B.n26 163.367
R686 B.n27 B.n26 163.367
R687 B.n28 B.n27 163.367
R688 B.n615 B.n28 163.367
R689 B.n615 B.n33 163.367
R690 B.n34 B.n33 163.367
R691 B.n35 B.n34 163.367
R692 B.n620 B.n35 163.367
R693 B.n620 B.n40 163.367
R694 B.n41 B.n40 163.367
R695 B.n42 B.n41 163.367
R696 B.n625 B.n42 163.367
R697 B.n625 B.n47 163.367
R698 B.n48 B.n47 163.367
R699 B.n49 B.n48 163.367
R700 B.n630 B.n49 163.367
R701 B.n630 B.n54 163.367
R702 B.n55 B.n54 163.367
R703 B.n56 B.n55 163.367
R704 B.n635 B.n56 163.367
R705 B.n635 B.n61 163.367
R706 B.n62 B.n61 163.367
R707 B.n347 B.n346 163.367
R708 B.n486 B.n346 163.367
R709 B.n484 B.n483 163.367
R710 B.n480 B.n479 163.367
R711 B.n476 B.n475 163.367
R712 B.n472 B.n471 163.367
R713 B.n468 B.n467 163.367
R714 B.n464 B.n463 163.367
R715 B.n460 B.n459 163.367
R716 B.n456 B.n455 163.367
R717 B.n452 B.n451 163.367
R718 B.n448 B.n447 163.367
R719 B.n444 B.n443 163.367
R720 B.n440 B.n439 163.367
R721 B.n436 B.n435 163.367
R722 B.n432 B.n431 163.367
R723 B.n428 B.n427 163.367
R724 B.n424 B.n423 163.367
R725 B.n420 B.n419 163.367
R726 B.n416 B.n415 163.367
R727 B.n412 B.n411 163.367
R728 B.n408 B.n407 163.367
R729 B.n404 B.n403 163.367
R730 B.n400 B.n399 163.367
R731 B.n396 B.n395 163.367
R732 B.n392 B.n391 163.367
R733 B.n388 B.n387 163.367
R734 B.n384 B.n383 163.367
R735 B.n380 B.n379 163.367
R736 B.n376 B.n375 163.367
R737 B.n372 B.n371 163.367
R738 B.n368 B.n367 163.367
R739 B.n364 B.n363 163.367
R740 B.n360 B.n359 163.367
R741 B.n356 B.n355 163.367
R742 B.n494 B.n311 163.367
R743 B.n500 B.n307 163.367
R744 B.n500 B.n305 163.367
R745 B.n504 B.n305 163.367
R746 B.n504 B.n299 163.367
R747 B.n512 B.n299 163.367
R748 B.n512 B.n297 163.367
R749 B.n516 B.n297 163.367
R750 B.n516 B.n291 163.367
R751 B.n524 B.n291 163.367
R752 B.n524 B.n289 163.367
R753 B.n528 B.n289 163.367
R754 B.n528 B.n283 163.367
R755 B.n536 B.n283 163.367
R756 B.n536 B.n281 163.367
R757 B.n540 B.n281 163.367
R758 B.n540 B.n275 163.367
R759 B.n548 B.n275 163.367
R760 B.n548 B.n273 163.367
R761 B.n552 B.n273 163.367
R762 B.n552 B.n267 163.367
R763 B.n560 B.n267 163.367
R764 B.n560 B.n265 163.367
R765 B.n564 B.n265 163.367
R766 B.n564 B.n259 163.367
R767 B.n572 B.n259 163.367
R768 B.n572 B.n257 163.367
R769 B.n576 B.n257 163.367
R770 B.n576 B.n251 163.367
R771 B.n585 B.n251 163.367
R772 B.n585 B.n249 163.367
R773 B.n589 B.n249 163.367
R774 B.n589 B.n3 163.367
R775 B.n710 B.n3 163.367
R776 B.n706 B.n2 163.367
R777 B.n706 B.n705 163.367
R778 B.n705 B.n9 163.367
R779 B.n701 B.n9 163.367
R780 B.n701 B.n11 163.367
R781 B.n697 B.n11 163.367
R782 B.n697 B.n16 163.367
R783 B.n693 B.n16 163.367
R784 B.n693 B.n18 163.367
R785 B.n689 B.n18 163.367
R786 B.n689 B.n23 163.367
R787 B.n685 B.n23 163.367
R788 B.n685 B.n25 163.367
R789 B.n681 B.n25 163.367
R790 B.n681 B.n30 163.367
R791 B.n677 B.n30 163.367
R792 B.n677 B.n32 163.367
R793 B.n673 B.n32 163.367
R794 B.n673 B.n37 163.367
R795 B.n669 B.n37 163.367
R796 B.n669 B.n39 163.367
R797 B.n665 B.n39 163.367
R798 B.n665 B.n44 163.367
R799 B.n661 B.n44 163.367
R800 B.n661 B.n46 163.367
R801 B.n657 B.n46 163.367
R802 B.n657 B.n51 163.367
R803 B.n653 B.n51 163.367
R804 B.n653 B.n53 163.367
R805 B.n649 B.n53 163.367
R806 B.n649 B.n58 163.367
R807 B.n645 B.n58 163.367
R808 B.n645 B.n60 163.367
R809 B.n493 B.n308 109.641
R810 B.n643 B.n642 109.641
R811 B.n99 B.t20 108.231
R812 B.n351 B.t14 108.231
R813 B.n101 B.t17 108.221
R814 B.n348 B.t11 108.221
R815 B.n100 B.t21 74.4847
R816 B.n352 B.t13 74.4847
R817 B.n102 B.t18 74.4749
R818 B.n349 B.t10 74.4749
R819 B.n103 B.n63 71.676
R820 B.n107 B.n64 71.676
R821 B.n111 B.n65 71.676
R822 B.n115 B.n66 71.676
R823 B.n119 B.n67 71.676
R824 B.n123 B.n68 71.676
R825 B.n127 B.n69 71.676
R826 B.n131 B.n70 71.676
R827 B.n135 B.n71 71.676
R828 B.n139 B.n72 71.676
R829 B.n143 B.n73 71.676
R830 B.n147 B.n74 71.676
R831 B.n151 B.n75 71.676
R832 B.n155 B.n76 71.676
R833 B.n159 B.n77 71.676
R834 B.n163 B.n78 71.676
R835 B.n168 B.n79 71.676
R836 B.n172 B.n80 71.676
R837 B.n176 B.n81 71.676
R838 B.n180 B.n82 71.676
R839 B.n184 B.n83 71.676
R840 B.n189 B.n84 71.676
R841 B.n193 B.n85 71.676
R842 B.n197 B.n86 71.676
R843 B.n201 B.n87 71.676
R844 B.n205 B.n88 71.676
R845 B.n209 B.n89 71.676
R846 B.n213 B.n90 71.676
R847 B.n217 B.n91 71.676
R848 B.n221 B.n92 71.676
R849 B.n225 B.n93 71.676
R850 B.n229 B.n94 71.676
R851 B.n233 B.n95 71.676
R852 B.n237 B.n96 71.676
R853 B.n241 B.n97 71.676
R854 B.n641 B.n98 71.676
R855 B.n641 B.n640 71.676
R856 B.n243 B.n97 71.676
R857 B.n240 B.n96 71.676
R858 B.n236 B.n95 71.676
R859 B.n232 B.n94 71.676
R860 B.n228 B.n93 71.676
R861 B.n224 B.n92 71.676
R862 B.n220 B.n91 71.676
R863 B.n216 B.n90 71.676
R864 B.n212 B.n89 71.676
R865 B.n208 B.n88 71.676
R866 B.n204 B.n87 71.676
R867 B.n200 B.n86 71.676
R868 B.n196 B.n85 71.676
R869 B.n192 B.n84 71.676
R870 B.n188 B.n83 71.676
R871 B.n183 B.n82 71.676
R872 B.n179 B.n81 71.676
R873 B.n175 B.n80 71.676
R874 B.n171 B.n79 71.676
R875 B.n167 B.n78 71.676
R876 B.n162 B.n77 71.676
R877 B.n158 B.n76 71.676
R878 B.n154 B.n75 71.676
R879 B.n150 B.n74 71.676
R880 B.n146 B.n73 71.676
R881 B.n142 B.n72 71.676
R882 B.n138 B.n71 71.676
R883 B.n134 B.n70 71.676
R884 B.n130 B.n69 71.676
R885 B.n126 B.n68 71.676
R886 B.n122 B.n67 71.676
R887 B.n118 B.n66 71.676
R888 B.n114 B.n65 71.676
R889 B.n110 B.n64 71.676
R890 B.n106 B.n63 71.676
R891 B.n492 B.n491 71.676
R892 B.n486 B.n312 71.676
R893 B.n483 B.n313 71.676
R894 B.n479 B.n314 71.676
R895 B.n475 B.n315 71.676
R896 B.n471 B.n316 71.676
R897 B.n467 B.n317 71.676
R898 B.n463 B.n318 71.676
R899 B.n459 B.n319 71.676
R900 B.n455 B.n320 71.676
R901 B.n451 B.n321 71.676
R902 B.n447 B.n322 71.676
R903 B.n443 B.n323 71.676
R904 B.n439 B.n324 71.676
R905 B.n435 B.n325 71.676
R906 B.n431 B.n326 71.676
R907 B.n427 B.n327 71.676
R908 B.n423 B.n328 71.676
R909 B.n419 B.n329 71.676
R910 B.n415 B.n330 71.676
R911 B.n411 B.n331 71.676
R912 B.n407 B.n332 71.676
R913 B.n403 B.n333 71.676
R914 B.n399 B.n334 71.676
R915 B.n395 B.n335 71.676
R916 B.n391 B.n336 71.676
R917 B.n387 B.n337 71.676
R918 B.n383 B.n338 71.676
R919 B.n379 B.n339 71.676
R920 B.n375 B.n340 71.676
R921 B.n371 B.n341 71.676
R922 B.n367 B.n342 71.676
R923 B.n363 B.n343 71.676
R924 B.n359 B.n344 71.676
R925 B.n355 B.n345 71.676
R926 B.n492 B.n347 71.676
R927 B.n484 B.n312 71.676
R928 B.n480 B.n313 71.676
R929 B.n476 B.n314 71.676
R930 B.n472 B.n315 71.676
R931 B.n468 B.n316 71.676
R932 B.n464 B.n317 71.676
R933 B.n460 B.n318 71.676
R934 B.n456 B.n319 71.676
R935 B.n452 B.n320 71.676
R936 B.n448 B.n321 71.676
R937 B.n444 B.n322 71.676
R938 B.n440 B.n323 71.676
R939 B.n436 B.n324 71.676
R940 B.n432 B.n325 71.676
R941 B.n428 B.n326 71.676
R942 B.n424 B.n327 71.676
R943 B.n420 B.n328 71.676
R944 B.n416 B.n329 71.676
R945 B.n412 B.n330 71.676
R946 B.n408 B.n331 71.676
R947 B.n404 B.n332 71.676
R948 B.n400 B.n333 71.676
R949 B.n396 B.n334 71.676
R950 B.n392 B.n335 71.676
R951 B.n388 B.n336 71.676
R952 B.n384 B.n337 71.676
R953 B.n380 B.n338 71.676
R954 B.n376 B.n339 71.676
R955 B.n372 B.n340 71.676
R956 B.n368 B.n341 71.676
R957 B.n364 B.n342 71.676
R958 B.n360 B.n343 71.676
R959 B.n356 B.n344 71.676
R960 B.n345 B.n311 71.676
R961 B.n711 B.n710 71.676
R962 B.n711 B.n2 71.676
R963 B.n165 B.n102 59.5399
R964 B.n186 B.n100 59.5399
R965 B.n353 B.n352 59.5399
R966 B.n350 B.n349 59.5399
R967 B.n499 B.n308 54.4203
R968 B.n499 B.n304 54.4203
R969 B.n505 B.n304 54.4203
R970 B.n505 B.n300 54.4203
R971 B.n511 B.n300 54.4203
R972 B.n517 B.n296 54.4203
R973 B.n517 B.n292 54.4203
R974 B.n523 B.n292 54.4203
R975 B.n523 B.n288 54.4203
R976 B.n529 B.n288 54.4203
R977 B.n529 B.n284 54.4203
R978 B.n535 B.n284 54.4203
R979 B.n541 B.n280 54.4203
R980 B.n541 B.n276 54.4203
R981 B.n547 B.n276 54.4203
R982 B.n547 B.n272 54.4203
R983 B.n553 B.n272 54.4203
R984 B.n559 B.n268 54.4203
R985 B.n559 B.n263 54.4203
R986 B.n565 B.n263 54.4203
R987 B.n565 B.n264 54.4203
R988 B.n571 B.n256 54.4203
R989 B.n577 B.n256 54.4203
R990 B.n577 B.n252 54.4203
R991 B.n584 B.n252 54.4203
R992 B.n590 B.n248 54.4203
R993 B.n590 B.n4 54.4203
R994 B.n709 B.n4 54.4203
R995 B.n709 B.n708 54.4203
R996 B.n708 B.n707 54.4203
R997 B.n707 B.n8 54.4203
R998 B.n599 B.n8 54.4203
R999 B.n700 B.n699 54.4203
R1000 B.n699 B.n698 54.4203
R1001 B.n698 B.n15 54.4203
R1002 B.n692 B.n15 54.4203
R1003 B.n691 B.n690 54.4203
R1004 B.n690 B.n22 54.4203
R1005 B.n684 B.n22 54.4203
R1006 B.n684 B.n683 54.4203
R1007 B.n682 B.n29 54.4203
R1008 B.n676 B.n29 54.4203
R1009 B.n676 B.n675 54.4203
R1010 B.n675 B.n674 54.4203
R1011 B.n674 B.n36 54.4203
R1012 B.n668 B.n667 54.4203
R1013 B.n667 B.n666 54.4203
R1014 B.n666 B.n43 54.4203
R1015 B.n660 B.n43 54.4203
R1016 B.n660 B.n659 54.4203
R1017 B.n659 B.n658 54.4203
R1018 B.n658 B.n50 54.4203
R1019 B.n652 B.n651 54.4203
R1020 B.n651 B.n650 54.4203
R1021 B.n650 B.n57 54.4203
R1022 B.n644 B.n57 54.4203
R1023 B.n644 B.n643 54.4203
R1024 B.n535 B.t1 53.62
R1025 B.n668 B.t4 53.62
R1026 B.t3 B.n268 48.8182
R1027 B.n683 B.t5 48.8182
R1028 B.n571 B.t2 42.4159
R1029 B.n692 B.t6 42.4159
R1030 B.n511 B.t9 36.0136
R1031 B.t0 B.n248 36.0136
R1032 B.n599 B.t7 36.0136
R1033 B.n652 B.t16 36.0136
R1034 B.n490 B.n306 34.8103
R1035 B.n496 B.n495 34.8103
R1036 B.n639 B.n638 34.8103
R1037 B.n104 B.n59 34.8103
R1038 B.n102 B.n101 33.746
R1039 B.n100 B.n99 33.746
R1040 B.n352 B.n351 33.746
R1041 B.n349 B.n348 33.746
R1042 B.t9 B.n296 18.4072
R1043 B.n584 B.t0 18.4072
R1044 B.n700 B.t7 18.4072
R1045 B.t16 B.n50 18.4072
R1046 B B.n712 18.0485
R1047 B.n264 B.t2 12.0049
R1048 B.t6 B.n691 12.0049
R1049 B.n501 B.n306 10.6151
R1050 B.n502 B.n501 10.6151
R1051 B.n503 B.n502 10.6151
R1052 B.n503 B.n298 10.6151
R1053 B.n513 B.n298 10.6151
R1054 B.n514 B.n513 10.6151
R1055 B.n515 B.n514 10.6151
R1056 B.n515 B.n290 10.6151
R1057 B.n525 B.n290 10.6151
R1058 B.n526 B.n525 10.6151
R1059 B.n527 B.n526 10.6151
R1060 B.n527 B.n282 10.6151
R1061 B.n537 B.n282 10.6151
R1062 B.n538 B.n537 10.6151
R1063 B.n539 B.n538 10.6151
R1064 B.n539 B.n274 10.6151
R1065 B.n549 B.n274 10.6151
R1066 B.n550 B.n549 10.6151
R1067 B.n551 B.n550 10.6151
R1068 B.n551 B.n266 10.6151
R1069 B.n561 B.n266 10.6151
R1070 B.n562 B.n561 10.6151
R1071 B.n563 B.n562 10.6151
R1072 B.n563 B.n258 10.6151
R1073 B.n573 B.n258 10.6151
R1074 B.n574 B.n573 10.6151
R1075 B.n575 B.n574 10.6151
R1076 B.n575 B.n250 10.6151
R1077 B.n586 B.n250 10.6151
R1078 B.n587 B.n586 10.6151
R1079 B.n588 B.n587 10.6151
R1080 B.n588 B.n0 10.6151
R1081 B.n490 B.n489 10.6151
R1082 B.n489 B.n488 10.6151
R1083 B.n488 B.n487 10.6151
R1084 B.n487 B.n485 10.6151
R1085 B.n485 B.n482 10.6151
R1086 B.n482 B.n481 10.6151
R1087 B.n481 B.n478 10.6151
R1088 B.n478 B.n477 10.6151
R1089 B.n477 B.n474 10.6151
R1090 B.n474 B.n473 10.6151
R1091 B.n473 B.n470 10.6151
R1092 B.n470 B.n469 10.6151
R1093 B.n469 B.n466 10.6151
R1094 B.n466 B.n465 10.6151
R1095 B.n465 B.n462 10.6151
R1096 B.n462 B.n461 10.6151
R1097 B.n461 B.n458 10.6151
R1098 B.n458 B.n457 10.6151
R1099 B.n457 B.n454 10.6151
R1100 B.n454 B.n453 10.6151
R1101 B.n453 B.n450 10.6151
R1102 B.n450 B.n449 10.6151
R1103 B.n449 B.n446 10.6151
R1104 B.n446 B.n445 10.6151
R1105 B.n445 B.n442 10.6151
R1106 B.n442 B.n441 10.6151
R1107 B.n441 B.n438 10.6151
R1108 B.n438 B.n437 10.6151
R1109 B.n437 B.n434 10.6151
R1110 B.n434 B.n433 10.6151
R1111 B.n430 B.n429 10.6151
R1112 B.n429 B.n426 10.6151
R1113 B.n426 B.n425 10.6151
R1114 B.n425 B.n422 10.6151
R1115 B.n422 B.n421 10.6151
R1116 B.n421 B.n418 10.6151
R1117 B.n418 B.n417 10.6151
R1118 B.n417 B.n414 10.6151
R1119 B.n414 B.n413 10.6151
R1120 B.n410 B.n409 10.6151
R1121 B.n409 B.n406 10.6151
R1122 B.n406 B.n405 10.6151
R1123 B.n405 B.n402 10.6151
R1124 B.n402 B.n401 10.6151
R1125 B.n401 B.n398 10.6151
R1126 B.n398 B.n397 10.6151
R1127 B.n397 B.n394 10.6151
R1128 B.n394 B.n393 10.6151
R1129 B.n393 B.n390 10.6151
R1130 B.n390 B.n389 10.6151
R1131 B.n389 B.n386 10.6151
R1132 B.n386 B.n385 10.6151
R1133 B.n385 B.n382 10.6151
R1134 B.n382 B.n381 10.6151
R1135 B.n381 B.n378 10.6151
R1136 B.n378 B.n377 10.6151
R1137 B.n377 B.n374 10.6151
R1138 B.n374 B.n373 10.6151
R1139 B.n373 B.n370 10.6151
R1140 B.n370 B.n369 10.6151
R1141 B.n369 B.n366 10.6151
R1142 B.n366 B.n365 10.6151
R1143 B.n365 B.n362 10.6151
R1144 B.n362 B.n361 10.6151
R1145 B.n361 B.n358 10.6151
R1146 B.n358 B.n357 10.6151
R1147 B.n357 B.n354 10.6151
R1148 B.n354 B.n310 10.6151
R1149 B.n495 B.n310 10.6151
R1150 B.n497 B.n496 10.6151
R1151 B.n497 B.n302 10.6151
R1152 B.n507 B.n302 10.6151
R1153 B.n508 B.n507 10.6151
R1154 B.n509 B.n508 10.6151
R1155 B.n509 B.n294 10.6151
R1156 B.n519 B.n294 10.6151
R1157 B.n520 B.n519 10.6151
R1158 B.n521 B.n520 10.6151
R1159 B.n521 B.n286 10.6151
R1160 B.n531 B.n286 10.6151
R1161 B.n532 B.n531 10.6151
R1162 B.n533 B.n532 10.6151
R1163 B.n533 B.n278 10.6151
R1164 B.n543 B.n278 10.6151
R1165 B.n544 B.n543 10.6151
R1166 B.n545 B.n544 10.6151
R1167 B.n545 B.n270 10.6151
R1168 B.n555 B.n270 10.6151
R1169 B.n556 B.n555 10.6151
R1170 B.n557 B.n556 10.6151
R1171 B.n557 B.n261 10.6151
R1172 B.n567 B.n261 10.6151
R1173 B.n568 B.n567 10.6151
R1174 B.n569 B.n568 10.6151
R1175 B.n569 B.n254 10.6151
R1176 B.n579 B.n254 10.6151
R1177 B.n580 B.n579 10.6151
R1178 B.n582 B.n580 10.6151
R1179 B.n582 B.n581 10.6151
R1180 B.n581 B.n246 10.6151
R1181 B.n593 B.n246 10.6151
R1182 B.n594 B.n593 10.6151
R1183 B.n595 B.n594 10.6151
R1184 B.n596 B.n595 10.6151
R1185 B.n597 B.n596 10.6151
R1186 B.n601 B.n597 10.6151
R1187 B.n602 B.n601 10.6151
R1188 B.n603 B.n602 10.6151
R1189 B.n604 B.n603 10.6151
R1190 B.n606 B.n604 10.6151
R1191 B.n607 B.n606 10.6151
R1192 B.n608 B.n607 10.6151
R1193 B.n609 B.n608 10.6151
R1194 B.n611 B.n609 10.6151
R1195 B.n612 B.n611 10.6151
R1196 B.n613 B.n612 10.6151
R1197 B.n614 B.n613 10.6151
R1198 B.n616 B.n614 10.6151
R1199 B.n617 B.n616 10.6151
R1200 B.n618 B.n617 10.6151
R1201 B.n619 B.n618 10.6151
R1202 B.n621 B.n619 10.6151
R1203 B.n622 B.n621 10.6151
R1204 B.n623 B.n622 10.6151
R1205 B.n624 B.n623 10.6151
R1206 B.n626 B.n624 10.6151
R1207 B.n627 B.n626 10.6151
R1208 B.n628 B.n627 10.6151
R1209 B.n629 B.n628 10.6151
R1210 B.n631 B.n629 10.6151
R1211 B.n632 B.n631 10.6151
R1212 B.n633 B.n632 10.6151
R1213 B.n634 B.n633 10.6151
R1214 B.n636 B.n634 10.6151
R1215 B.n637 B.n636 10.6151
R1216 B.n638 B.n637 10.6151
R1217 B.n704 B.n1 10.6151
R1218 B.n704 B.n703 10.6151
R1219 B.n703 B.n702 10.6151
R1220 B.n702 B.n10 10.6151
R1221 B.n696 B.n10 10.6151
R1222 B.n696 B.n695 10.6151
R1223 B.n695 B.n694 10.6151
R1224 B.n694 B.n17 10.6151
R1225 B.n688 B.n17 10.6151
R1226 B.n688 B.n687 10.6151
R1227 B.n687 B.n686 10.6151
R1228 B.n686 B.n24 10.6151
R1229 B.n680 B.n24 10.6151
R1230 B.n680 B.n679 10.6151
R1231 B.n679 B.n678 10.6151
R1232 B.n678 B.n31 10.6151
R1233 B.n672 B.n31 10.6151
R1234 B.n672 B.n671 10.6151
R1235 B.n671 B.n670 10.6151
R1236 B.n670 B.n38 10.6151
R1237 B.n664 B.n38 10.6151
R1238 B.n664 B.n663 10.6151
R1239 B.n663 B.n662 10.6151
R1240 B.n662 B.n45 10.6151
R1241 B.n656 B.n45 10.6151
R1242 B.n656 B.n655 10.6151
R1243 B.n655 B.n654 10.6151
R1244 B.n654 B.n52 10.6151
R1245 B.n648 B.n52 10.6151
R1246 B.n648 B.n647 10.6151
R1247 B.n647 B.n646 10.6151
R1248 B.n646 B.n59 10.6151
R1249 B.n105 B.n104 10.6151
R1250 B.n108 B.n105 10.6151
R1251 B.n109 B.n108 10.6151
R1252 B.n112 B.n109 10.6151
R1253 B.n113 B.n112 10.6151
R1254 B.n116 B.n113 10.6151
R1255 B.n117 B.n116 10.6151
R1256 B.n120 B.n117 10.6151
R1257 B.n121 B.n120 10.6151
R1258 B.n124 B.n121 10.6151
R1259 B.n125 B.n124 10.6151
R1260 B.n128 B.n125 10.6151
R1261 B.n129 B.n128 10.6151
R1262 B.n132 B.n129 10.6151
R1263 B.n133 B.n132 10.6151
R1264 B.n136 B.n133 10.6151
R1265 B.n137 B.n136 10.6151
R1266 B.n140 B.n137 10.6151
R1267 B.n141 B.n140 10.6151
R1268 B.n144 B.n141 10.6151
R1269 B.n145 B.n144 10.6151
R1270 B.n148 B.n145 10.6151
R1271 B.n149 B.n148 10.6151
R1272 B.n152 B.n149 10.6151
R1273 B.n153 B.n152 10.6151
R1274 B.n156 B.n153 10.6151
R1275 B.n157 B.n156 10.6151
R1276 B.n160 B.n157 10.6151
R1277 B.n161 B.n160 10.6151
R1278 B.n164 B.n161 10.6151
R1279 B.n169 B.n166 10.6151
R1280 B.n170 B.n169 10.6151
R1281 B.n173 B.n170 10.6151
R1282 B.n174 B.n173 10.6151
R1283 B.n177 B.n174 10.6151
R1284 B.n178 B.n177 10.6151
R1285 B.n181 B.n178 10.6151
R1286 B.n182 B.n181 10.6151
R1287 B.n185 B.n182 10.6151
R1288 B.n190 B.n187 10.6151
R1289 B.n191 B.n190 10.6151
R1290 B.n194 B.n191 10.6151
R1291 B.n195 B.n194 10.6151
R1292 B.n198 B.n195 10.6151
R1293 B.n199 B.n198 10.6151
R1294 B.n202 B.n199 10.6151
R1295 B.n203 B.n202 10.6151
R1296 B.n206 B.n203 10.6151
R1297 B.n207 B.n206 10.6151
R1298 B.n210 B.n207 10.6151
R1299 B.n211 B.n210 10.6151
R1300 B.n214 B.n211 10.6151
R1301 B.n215 B.n214 10.6151
R1302 B.n218 B.n215 10.6151
R1303 B.n219 B.n218 10.6151
R1304 B.n222 B.n219 10.6151
R1305 B.n223 B.n222 10.6151
R1306 B.n226 B.n223 10.6151
R1307 B.n227 B.n226 10.6151
R1308 B.n230 B.n227 10.6151
R1309 B.n231 B.n230 10.6151
R1310 B.n234 B.n231 10.6151
R1311 B.n235 B.n234 10.6151
R1312 B.n238 B.n235 10.6151
R1313 B.n239 B.n238 10.6151
R1314 B.n242 B.n239 10.6151
R1315 B.n244 B.n242 10.6151
R1316 B.n245 B.n244 10.6151
R1317 B.n639 B.n245 10.6151
R1318 B.n433 B.n350 9.36635
R1319 B.n410 B.n353 9.36635
R1320 B.n165 B.n164 9.36635
R1321 B.n187 B.n186 9.36635
R1322 B.n712 B.n0 8.11757
R1323 B.n712 B.n1 8.11757
R1324 B.n553 B.t3 5.60254
R1325 B.t5 B.n682 5.60254
R1326 B.n430 B.n350 1.24928
R1327 B.n413 B.n353 1.24928
R1328 B.n166 B.n165 1.24928
R1329 B.n186 B.n185 1.24928
R1330 B.t1 B.n280 0.800791
R1331 B.t4 B.n36 0.800791
R1332 VP.n26 VP.n25 180.385
R1333 VP.n46 VP.n45 180.385
R1334 VP.n24 VP.n23 180.385
R1335 VP.n11 VP.t2 176.014
R1336 VP.n12 VP.n9 161.3
R1337 VP.n14 VP.n13 161.3
R1338 VP.n15 VP.n8 161.3
R1339 VP.n18 VP.n17 161.3
R1340 VP.n19 VP.n7 161.3
R1341 VP.n21 VP.n20 161.3
R1342 VP.n22 VP.n6 161.3
R1343 VP.n44 VP.n0 161.3
R1344 VP.n43 VP.n42 161.3
R1345 VP.n41 VP.n1 161.3
R1346 VP.n40 VP.n39 161.3
R1347 VP.n37 VP.n2 161.3
R1348 VP.n36 VP.n35 161.3
R1349 VP.n34 VP.n3 161.3
R1350 VP.n33 VP.n32 161.3
R1351 VP.n30 VP.n4 161.3
R1352 VP.n29 VP.n28 161.3
R1353 VP.n27 VP.n5 161.3
R1354 VP.n25 VP.t4 144.772
R1355 VP.n31 VP.t5 144.772
R1356 VP.n38 VP.t1 144.772
R1357 VP.n45 VP.t7 144.772
R1358 VP.n23 VP.t0 144.772
R1359 VP.n16 VP.t3 144.772
R1360 VP.n10 VP.t6 144.772
R1361 VP.n30 VP.n29 56.5193
R1362 VP.n43 VP.n1 56.5193
R1363 VP.n21 VP.n7 56.5193
R1364 VP.n11 VP.n10 47.8106
R1365 VP.n26 VP.n24 42.4853
R1366 VP.n36 VP.n3 40.4934
R1367 VP.n37 VP.n36 40.4934
R1368 VP.n15 VP.n14 40.4934
R1369 VP.n14 VP.n9 40.4934
R1370 VP.n29 VP.n5 24.4675
R1371 VP.n32 VP.n30 24.4675
R1372 VP.n39 VP.n1 24.4675
R1373 VP.n44 VP.n43 24.4675
R1374 VP.n22 VP.n21 24.4675
R1375 VP.n17 VP.n7 24.4675
R1376 VP.n12 VP.n11 18.2406
R1377 VP.n31 VP.n3 18.1061
R1378 VP.n38 VP.n37 18.1061
R1379 VP.n16 VP.n15 18.1061
R1380 VP.n10 VP.n9 18.1061
R1381 VP.n32 VP.n31 6.36192
R1382 VP.n39 VP.n38 6.36192
R1383 VP.n17 VP.n16 6.36192
R1384 VP.n25 VP.n5 5.38324
R1385 VP.n45 VP.n44 5.38324
R1386 VP.n23 VP.n22 5.38324
R1387 VP.n13 VP.n12 0.189894
R1388 VP.n13 VP.n8 0.189894
R1389 VP.n18 VP.n8 0.189894
R1390 VP.n19 VP.n18 0.189894
R1391 VP.n20 VP.n19 0.189894
R1392 VP.n20 VP.n6 0.189894
R1393 VP.n24 VP.n6 0.189894
R1394 VP.n27 VP.n26 0.189894
R1395 VP.n28 VP.n27 0.189894
R1396 VP.n28 VP.n4 0.189894
R1397 VP.n33 VP.n4 0.189894
R1398 VP.n34 VP.n33 0.189894
R1399 VP.n35 VP.n34 0.189894
R1400 VP.n35 VP.n2 0.189894
R1401 VP.n40 VP.n2 0.189894
R1402 VP.n41 VP.n40 0.189894
R1403 VP.n42 VP.n41 0.189894
R1404 VP.n42 VP.n0 0.189894
R1405 VP.n46 VP.n0 0.189894
R1406 VP VP.n46 0.0516364
R1407 VDD1 VDD1.n0 64.0446
R1408 VDD1.n3 VDD1.n2 63.931
R1409 VDD1.n3 VDD1.n1 63.931
R1410 VDD1.n5 VDD1.n4 63.2364
R1411 VDD1.n5 VDD1.n3 38.35
R1412 VDD1.n4 VDD1.t4 2.33816
R1413 VDD1.n4 VDD1.t7 2.33816
R1414 VDD1.n0 VDD1.t5 2.33816
R1415 VDD1.n0 VDD1.t1 2.33816
R1416 VDD1.n2 VDD1.t6 2.33816
R1417 VDD1.n2 VDD1.t0 2.33816
R1418 VDD1.n1 VDD1.t3 2.33816
R1419 VDD1.n1 VDD1.t2 2.33816
R1420 VDD1 VDD1.n5 0.69231
C0 VP VTAIL 5.52528f
C1 VDD1 VDD2 1.18364f
C2 VDD1 VP 5.59166f
C3 VDD1 VTAIL 6.89801f
C4 VN VDD2 5.34899f
C5 VN VP 5.55774f
C6 VN VTAIL 5.51117f
C7 VP VDD2 0.393108f
C8 VDD1 VN 0.149642f
C9 VTAIL VDD2 6.94445f
C10 VDD2 B 3.904134f
C11 VDD1 B 4.218867f
C12 VTAIL B 7.519164f
C13 VN B 10.71106f
C14 VP B 9.179649f
C15 VDD1.t5 B 0.168873f
C16 VDD1.t1 B 0.168873f
C17 VDD1.n0 B 1.46452f
C18 VDD1.t3 B 0.168873f
C19 VDD1.t2 B 0.168873f
C20 VDD1.n1 B 1.4637f
C21 VDD1.t6 B 0.168873f
C22 VDD1.t0 B 0.168873f
C23 VDD1.n2 B 1.4637f
C24 VDD1.n3 B 2.45402f
C25 VDD1.t4 B 0.168873f
C26 VDD1.t7 B 0.168873f
C27 VDD1.n4 B 1.45935f
C28 VDD1.n5 B 2.31742f
C29 VP.n0 B 0.033388f
C30 VP.t7 B 1.07348f
C31 VP.n1 B 0.04781f
C32 VP.n2 B 0.033388f
C33 VP.t1 B 1.07348f
C34 VP.n3 B 0.05837f
C35 VP.n4 B 0.033388f
C36 VP.n5 B 0.038264f
C37 VP.n6 B 0.033388f
C38 VP.t0 B 1.07348f
C39 VP.n7 B 0.04781f
C40 VP.n8 B 0.033388f
C41 VP.t3 B 1.07348f
C42 VP.n9 B 0.05837f
C43 VP.t2 B 1.16652f
C44 VP.t6 B 1.07348f
C45 VP.n10 B 0.46983f
C46 VP.n11 B 0.478907f
C47 VP.n12 B 0.206329f
C48 VP.n13 B 0.033388f
C49 VP.n14 B 0.026991f
C50 VP.n15 B 0.05837f
C51 VP.n16 B 0.403207f
C52 VP.n17 B 0.039492f
C53 VP.n18 B 0.033388f
C54 VP.n19 B 0.033388f
C55 VP.n20 B 0.033388f
C56 VP.n21 B 0.049671f
C57 VP.n22 B 0.038264f
C58 VP.n23 B 0.459949f
C59 VP.n24 B 1.4114f
C60 VP.t4 B 1.07348f
C61 VP.n25 B 0.459949f
C62 VP.n26 B 1.43965f
C63 VP.n27 B 0.033388f
C64 VP.n28 B 0.033388f
C65 VP.n29 B 0.049671f
C66 VP.n30 B 0.04781f
C67 VP.t5 B 1.07348f
C68 VP.n31 B 0.403207f
C69 VP.n32 B 0.039492f
C70 VP.n33 B 0.033388f
C71 VP.n34 B 0.033388f
C72 VP.n35 B 0.033388f
C73 VP.n36 B 0.026991f
C74 VP.n37 B 0.05837f
C75 VP.n38 B 0.403207f
C76 VP.n39 B 0.039492f
C77 VP.n40 B 0.033388f
C78 VP.n41 B 0.033388f
C79 VP.n42 B 0.033388f
C80 VP.n43 B 0.049671f
C81 VP.n44 B 0.038264f
C82 VP.n45 B 0.459949f
C83 VP.n46 B 0.032588f
C84 VDD2.t0 B 0.166058f
C85 VDD2.t7 B 0.166058f
C86 VDD2.n0 B 1.43931f
C87 VDD2.t3 B 0.166058f
C88 VDD2.t2 B 0.166058f
C89 VDD2.n1 B 1.43931f
C90 VDD2.n2 B 2.36056f
C91 VDD2.t5 B 0.166058f
C92 VDD2.t1 B 0.166058f
C93 VDD2.n3 B 1.43502f
C94 VDD2.n4 B 2.24902f
C95 VDD2.t6 B 0.166058f
C96 VDD2.t4 B 0.166058f
C97 VDD2.n5 B 1.43928f
C98 VTAIL.t14 B 0.135039f
C99 VTAIL.t10 B 0.135039f
C100 VTAIL.n0 B 1.10769f
C101 VTAIL.n1 B 0.302437f
C102 VTAIL.t8 B 1.41186f
C103 VTAIL.n2 B 0.393311f
C104 VTAIL.t0 B 1.41186f
C105 VTAIL.n3 B 0.393311f
C106 VTAIL.t3 B 0.135039f
C107 VTAIL.t2 B 0.135039f
C108 VTAIL.n4 B 1.10769f
C109 VTAIL.n5 B 0.396168f
C110 VTAIL.t1 B 1.41186f
C111 VTAIL.n6 B 1.20902f
C112 VTAIL.t9 B 1.41187f
C113 VTAIL.n7 B 1.20902f
C114 VTAIL.t11 B 0.135039f
C115 VTAIL.t15 B 0.135039f
C116 VTAIL.n8 B 1.10769f
C117 VTAIL.n9 B 0.396166f
C118 VTAIL.t12 B 1.41187f
C119 VTAIL.n10 B 0.393305f
C120 VTAIL.t7 B 1.41187f
C121 VTAIL.n11 B 0.393305f
C122 VTAIL.t6 B 0.135039f
C123 VTAIL.t5 B 0.135039f
C124 VTAIL.n12 B 1.10769f
C125 VTAIL.n13 B 0.396166f
C126 VTAIL.t4 B 1.41187f
C127 VTAIL.n14 B 1.20902f
C128 VTAIL.t13 B 1.41186f
C129 VTAIL.n15 B 1.20524f
C130 VN.n0 B 0.032696f
C131 VN.t5 B 1.05124f
C132 VN.n1 B 0.046819f
C133 VN.n2 B 0.032696f
C134 VN.t4 B 1.05124f
C135 VN.n3 B 0.057161f
C136 VN.t7 B 1.14236f
C137 VN.t0 B 1.05124f
C138 VN.n4 B 0.460097f
C139 VN.n5 B 0.468986f
C140 VN.n6 B 0.202054f
C141 VN.n7 B 0.032696f
C142 VN.n8 B 0.026432f
C143 VN.n9 B 0.057161f
C144 VN.n10 B 0.394854f
C145 VN.n11 B 0.038674f
C146 VN.n12 B 0.032696f
C147 VN.n13 B 0.032696f
C148 VN.n14 B 0.032696f
C149 VN.n15 B 0.048641f
C150 VN.n16 B 0.037471f
C151 VN.n17 B 0.450421f
C152 VN.n18 B 0.031913f
C153 VN.n19 B 0.032696f
C154 VN.t2 B 1.05124f
C155 VN.n20 B 0.046819f
C156 VN.n21 B 0.032696f
C157 VN.t6 B 1.05124f
C158 VN.n22 B 0.057161f
C159 VN.t3 B 1.14236f
C160 VN.t1 B 1.05124f
C161 VN.n23 B 0.460097f
C162 VN.n24 B 0.468986f
C163 VN.n25 B 0.202054f
C164 VN.n26 B 0.032696f
C165 VN.n27 B 0.026432f
C166 VN.n28 B 0.057161f
C167 VN.n29 B 0.394854f
C168 VN.n30 B 0.038674f
C169 VN.n31 B 0.032696f
C170 VN.n32 B 0.032696f
C171 VN.n33 B 0.032696f
C172 VN.n34 B 0.048641f
C173 VN.n35 B 0.037471f
C174 VN.n36 B 0.450421f
C175 VN.n37 B 1.40361f
.ends

