* NGSPICE file created from diff_pair_sample_0360.ext - technology: sky130A

.subckt diff_pair_sample_0360 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t12 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=7.2423 ps=37.92 w=18.57 l=3.41
X1 VDD1.t9 VP.t0 VTAIL.t18 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=3.06405 ps=18.9 w=18.57 l=3.41
X2 VTAIL.t8 VN.t1 VDD2.t8 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X3 VDD1.t8 VP.t1 VTAIL.t16 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=7.2423 ps=37.92 w=18.57 l=3.41
X4 B.t11 B.t9 B.t10 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=0 ps=0 w=18.57 l=3.41
X5 VTAIL.t4 VP.t2 VDD1.t7 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X6 VDD2.t7 VN.t2 VTAIL.t10 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X7 VDD2.t6 VN.t3 VTAIL.t7 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X8 VDD1.t6 VP.t3 VTAIL.t3 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=3.06405 ps=18.9 w=18.57 l=3.41
X9 VTAIL.t9 VN.t4 VDD2.t5 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X10 VTAIL.t15 VP.t4 VDD1.t5 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X11 VDD2.t4 VN.t5 VTAIL.t13 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=7.2423 ps=37.92 w=18.57 l=3.41
X12 VDD2.t3 VN.t6 VTAIL.t11 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=3.06405 ps=18.9 w=18.57 l=3.41
X13 B.t8 B.t6 B.t7 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=0 ps=0 w=18.57 l=3.41
X14 VDD1.t4 VP.t5 VTAIL.t19 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X15 VTAIL.t17 VP.t6 VDD1.t3 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X16 VTAIL.t2 VP.t7 VDD1.t2 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X17 VDD2.t2 VN.t7 VTAIL.t14 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=3.06405 ps=18.9 w=18.57 l=3.41
X18 B.t5 B.t3 B.t4 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=0 ps=0 w=18.57 l=3.41
X19 B.t2 B.t0 B.t1 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=7.2423 pd=37.92 as=0 ps=0 w=18.57 l=3.41
X20 VTAIL.t6 VN.t8 VDD2.t1 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X21 VDD1.t1 VP.t8 VTAIL.t1 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
X22 VDD1.t0 VP.t9 VTAIL.t0 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=7.2423 ps=37.92 w=18.57 l=3.41
X23 VTAIL.t5 VN.t9 VDD2.t0 w_n5458_n4682# sky130_fd_pr__pfet_01v8 ad=3.06405 pd=18.9 as=3.06405 ps=18.9 w=18.57 l=3.41
R0 VN.n64 VN.t5 164.869
R1 VN.n13 VN.t6 164.869
R2 VN.n98 VN.n97 161.3
R3 VN.n96 VN.n51 161.3
R4 VN.n95 VN.n94 161.3
R5 VN.n93 VN.n52 161.3
R6 VN.n92 VN.n91 161.3
R7 VN.n90 VN.n53 161.3
R8 VN.n89 VN.n88 161.3
R9 VN.n87 VN.n54 161.3
R10 VN.n86 VN.n85 161.3
R11 VN.n84 VN.n55 161.3
R12 VN.n83 VN.n82 161.3
R13 VN.n81 VN.n57 161.3
R14 VN.n80 VN.n79 161.3
R15 VN.n78 VN.n58 161.3
R16 VN.n77 VN.n76 161.3
R17 VN.n75 VN.n74 161.3
R18 VN.n73 VN.n60 161.3
R19 VN.n72 VN.n71 161.3
R20 VN.n70 VN.n61 161.3
R21 VN.n69 VN.n68 161.3
R22 VN.n67 VN.n62 161.3
R23 VN.n66 VN.n65 161.3
R24 VN.n48 VN.n47 161.3
R25 VN.n46 VN.n1 161.3
R26 VN.n45 VN.n44 161.3
R27 VN.n43 VN.n2 161.3
R28 VN.n42 VN.n41 161.3
R29 VN.n40 VN.n3 161.3
R30 VN.n39 VN.n38 161.3
R31 VN.n37 VN.n4 161.3
R32 VN.n36 VN.n35 161.3
R33 VN.n33 VN.n5 161.3
R34 VN.n32 VN.n31 161.3
R35 VN.n30 VN.n6 161.3
R36 VN.n29 VN.n28 161.3
R37 VN.n27 VN.n7 161.3
R38 VN.n26 VN.n25 161.3
R39 VN.n24 VN.n23 161.3
R40 VN.n22 VN.n9 161.3
R41 VN.n21 VN.n20 161.3
R42 VN.n19 VN.n10 161.3
R43 VN.n18 VN.n17 161.3
R44 VN.n16 VN.n11 161.3
R45 VN.n15 VN.n14 161.3
R46 VN.n12 VN.t1 131.244
R47 VN.n8 VN.t3 131.244
R48 VN.n34 VN.t9 131.244
R49 VN.n0 VN.t0 131.244
R50 VN.n63 VN.t8 131.244
R51 VN.n59 VN.t2 131.244
R52 VN.n56 VN.t4 131.244
R53 VN.n50 VN.t7 131.244
R54 VN.n49 VN.n0 78.8126
R55 VN.n99 VN.n50 78.8126
R56 VN VN.n99 62.748
R57 VN.n41 VN.n2 54.0911
R58 VN.n91 VN.n52 54.0911
R59 VN.n17 VN.n10 52.1486
R60 VN.n32 VN.n6 52.1486
R61 VN.n68 VN.n61 52.1486
R62 VN.n83 VN.n57 52.1486
R63 VN.n13 VN.n12 50.6338
R64 VN.n64 VN.n63 50.6338
R65 VN.n21 VN.n10 28.8382
R66 VN.n28 VN.n6 28.8382
R67 VN.n72 VN.n61 28.8382
R68 VN.n79 VN.n57 28.8382
R69 VN.n45 VN.n2 26.8957
R70 VN.n95 VN.n52 26.8957
R71 VN.n16 VN.n15 24.4675
R72 VN.n17 VN.n16 24.4675
R73 VN.n22 VN.n21 24.4675
R74 VN.n23 VN.n22 24.4675
R75 VN.n27 VN.n26 24.4675
R76 VN.n28 VN.n27 24.4675
R77 VN.n33 VN.n32 24.4675
R78 VN.n35 VN.n33 24.4675
R79 VN.n39 VN.n4 24.4675
R80 VN.n40 VN.n39 24.4675
R81 VN.n41 VN.n40 24.4675
R82 VN.n46 VN.n45 24.4675
R83 VN.n47 VN.n46 24.4675
R84 VN.n68 VN.n67 24.4675
R85 VN.n67 VN.n66 24.4675
R86 VN.n79 VN.n78 24.4675
R87 VN.n78 VN.n77 24.4675
R88 VN.n74 VN.n73 24.4675
R89 VN.n73 VN.n72 24.4675
R90 VN.n91 VN.n90 24.4675
R91 VN.n90 VN.n89 24.4675
R92 VN.n89 VN.n54 24.4675
R93 VN.n85 VN.n84 24.4675
R94 VN.n84 VN.n83 24.4675
R95 VN.n97 VN.n96 24.4675
R96 VN.n96 VN.n95 24.4675
R97 VN.n15 VN.n12 23.9782
R98 VN.n35 VN.n34 23.9782
R99 VN.n66 VN.n63 23.9782
R100 VN.n85 VN.n56 23.9782
R101 VN.n23 VN.n8 12.234
R102 VN.n26 VN.n8 12.234
R103 VN.n77 VN.n59 12.234
R104 VN.n74 VN.n59 12.234
R105 VN.n47 VN.n0 11.2553
R106 VN.n97 VN.n50 11.2553
R107 VN.n65 VN.n64 3.11119
R108 VN.n14 VN.n13 3.11119
R109 VN.n34 VN.n4 0.48984
R110 VN.n56 VN.n54 0.48984
R111 VN.n99 VN.n98 0.354971
R112 VN.n49 VN.n48 0.354971
R113 VN VN.n49 0.26696
R114 VN.n98 VN.n51 0.189894
R115 VN.n94 VN.n51 0.189894
R116 VN.n94 VN.n93 0.189894
R117 VN.n93 VN.n92 0.189894
R118 VN.n92 VN.n53 0.189894
R119 VN.n88 VN.n53 0.189894
R120 VN.n88 VN.n87 0.189894
R121 VN.n87 VN.n86 0.189894
R122 VN.n86 VN.n55 0.189894
R123 VN.n82 VN.n55 0.189894
R124 VN.n82 VN.n81 0.189894
R125 VN.n81 VN.n80 0.189894
R126 VN.n80 VN.n58 0.189894
R127 VN.n76 VN.n58 0.189894
R128 VN.n76 VN.n75 0.189894
R129 VN.n75 VN.n60 0.189894
R130 VN.n71 VN.n60 0.189894
R131 VN.n71 VN.n70 0.189894
R132 VN.n70 VN.n69 0.189894
R133 VN.n69 VN.n62 0.189894
R134 VN.n65 VN.n62 0.189894
R135 VN.n14 VN.n11 0.189894
R136 VN.n18 VN.n11 0.189894
R137 VN.n19 VN.n18 0.189894
R138 VN.n20 VN.n19 0.189894
R139 VN.n20 VN.n9 0.189894
R140 VN.n24 VN.n9 0.189894
R141 VN.n25 VN.n24 0.189894
R142 VN.n25 VN.n7 0.189894
R143 VN.n29 VN.n7 0.189894
R144 VN.n30 VN.n29 0.189894
R145 VN.n31 VN.n30 0.189894
R146 VN.n31 VN.n5 0.189894
R147 VN.n36 VN.n5 0.189894
R148 VN.n37 VN.n36 0.189894
R149 VN.n38 VN.n37 0.189894
R150 VN.n38 VN.n3 0.189894
R151 VN.n42 VN.n3 0.189894
R152 VN.n43 VN.n42 0.189894
R153 VN.n44 VN.n43 0.189894
R154 VN.n44 VN.n1 0.189894
R155 VN.n48 VN.n1 0.189894
R156 VTAIL.n11 VTAIL.t13 53.0223
R157 VTAIL.n17 VTAIL.t12 53.0221
R158 VTAIL.n2 VTAIL.t0 53.0221
R159 VTAIL.n16 VTAIL.t16 53.0221
R160 VTAIL.n15 VTAIL.n14 51.2719
R161 VTAIL.n13 VTAIL.n12 51.2719
R162 VTAIL.n10 VTAIL.n9 51.2719
R163 VTAIL.n8 VTAIL.n7 51.2719
R164 VTAIL.n19 VTAIL.n18 51.2717
R165 VTAIL.n1 VTAIL.n0 51.2717
R166 VTAIL.n4 VTAIL.n3 51.2717
R167 VTAIL.n6 VTAIL.n5 51.2717
R168 VTAIL.n8 VTAIL.n6 34.8238
R169 VTAIL.n17 VTAIL.n16 31.5996
R170 VTAIL.n10 VTAIL.n8 3.22464
R171 VTAIL.n11 VTAIL.n10 3.22464
R172 VTAIL.n15 VTAIL.n13 3.22464
R173 VTAIL.n16 VTAIL.n15 3.22464
R174 VTAIL.n6 VTAIL.n4 3.22464
R175 VTAIL.n4 VTAIL.n2 3.22464
R176 VTAIL.n19 VTAIL.n17 3.22464
R177 VTAIL VTAIL.n1 2.47679
R178 VTAIL.n13 VTAIL.n11 2.0824
R179 VTAIL.n2 VTAIL.n1 2.0824
R180 VTAIL.n18 VTAIL.t7 1.7509
R181 VTAIL.n18 VTAIL.t5 1.7509
R182 VTAIL.n0 VTAIL.t11 1.7509
R183 VTAIL.n0 VTAIL.t8 1.7509
R184 VTAIL.n3 VTAIL.t1 1.7509
R185 VTAIL.n3 VTAIL.t17 1.7509
R186 VTAIL.n5 VTAIL.t3 1.7509
R187 VTAIL.n5 VTAIL.t15 1.7509
R188 VTAIL.n14 VTAIL.t19 1.7509
R189 VTAIL.n14 VTAIL.t2 1.7509
R190 VTAIL.n12 VTAIL.t18 1.7509
R191 VTAIL.n12 VTAIL.t4 1.7509
R192 VTAIL.n9 VTAIL.t10 1.7509
R193 VTAIL.n9 VTAIL.t6 1.7509
R194 VTAIL.n7 VTAIL.t14 1.7509
R195 VTAIL.n7 VTAIL.t9 1.7509
R196 VTAIL VTAIL.n19 0.748345
R197 VDD2.n1 VDD2.t3 72.9251
R198 VDD2.n3 VDD2.n2 70.3132
R199 VDD2 VDD2.n7 70.3104
R200 VDD2.n4 VDD2.t2 69.7011
R201 VDD2.n6 VDD2.n5 67.9507
R202 VDD2.n1 VDD2.n0 67.9505
R203 VDD2.n4 VDD2.n3 55.0386
R204 VDD2.n6 VDD2.n4 3.22464
R205 VDD2.n7 VDD2.t1 1.7509
R206 VDD2.n7 VDD2.t4 1.7509
R207 VDD2.n5 VDD2.t5 1.7509
R208 VDD2.n5 VDD2.t7 1.7509
R209 VDD2.n2 VDD2.t0 1.7509
R210 VDD2.n2 VDD2.t9 1.7509
R211 VDD2.n0 VDD2.t8 1.7509
R212 VDD2.n0 VDD2.t6 1.7509
R213 VDD2 VDD2.n6 0.864724
R214 VDD2.n3 VDD2.n1 0.751188
R215 VP.n30 VP.t0 164.869
R216 VP.n32 VP.n31 161.3
R217 VP.n33 VP.n28 161.3
R218 VP.n35 VP.n34 161.3
R219 VP.n36 VP.n27 161.3
R220 VP.n38 VP.n37 161.3
R221 VP.n39 VP.n26 161.3
R222 VP.n41 VP.n40 161.3
R223 VP.n43 VP.n42 161.3
R224 VP.n44 VP.n24 161.3
R225 VP.n46 VP.n45 161.3
R226 VP.n47 VP.n23 161.3
R227 VP.n49 VP.n48 161.3
R228 VP.n50 VP.n22 161.3
R229 VP.n53 VP.n52 161.3
R230 VP.n54 VP.n21 161.3
R231 VP.n56 VP.n55 161.3
R232 VP.n57 VP.n20 161.3
R233 VP.n59 VP.n58 161.3
R234 VP.n60 VP.n19 161.3
R235 VP.n62 VP.n61 161.3
R236 VP.n63 VP.n18 161.3
R237 VP.n65 VP.n64 161.3
R238 VP.n115 VP.n114 161.3
R239 VP.n113 VP.n1 161.3
R240 VP.n112 VP.n111 161.3
R241 VP.n110 VP.n2 161.3
R242 VP.n109 VP.n108 161.3
R243 VP.n107 VP.n3 161.3
R244 VP.n106 VP.n105 161.3
R245 VP.n104 VP.n4 161.3
R246 VP.n103 VP.n102 161.3
R247 VP.n100 VP.n5 161.3
R248 VP.n99 VP.n98 161.3
R249 VP.n97 VP.n6 161.3
R250 VP.n96 VP.n95 161.3
R251 VP.n94 VP.n7 161.3
R252 VP.n93 VP.n92 161.3
R253 VP.n91 VP.n90 161.3
R254 VP.n89 VP.n9 161.3
R255 VP.n88 VP.n87 161.3
R256 VP.n86 VP.n10 161.3
R257 VP.n85 VP.n84 161.3
R258 VP.n83 VP.n11 161.3
R259 VP.n82 VP.n81 161.3
R260 VP.n80 VP.n79 161.3
R261 VP.n78 VP.n13 161.3
R262 VP.n77 VP.n76 161.3
R263 VP.n75 VP.n14 161.3
R264 VP.n74 VP.n73 161.3
R265 VP.n72 VP.n15 161.3
R266 VP.n71 VP.n70 161.3
R267 VP.n69 VP.n16 161.3
R268 VP.n67 VP.t3 131.244
R269 VP.n12 VP.t4 131.244
R270 VP.n8 VP.t8 131.244
R271 VP.n101 VP.t6 131.244
R272 VP.n0 VP.t9 131.244
R273 VP.n17 VP.t1 131.244
R274 VP.n51 VP.t7 131.244
R275 VP.n25 VP.t5 131.244
R276 VP.n29 VP.t2 131.244
R277 VP.n68 VP.n67 78.8126
R278 VP.n116 VP.n0 78.8126
R279 VP.n66 VP.n17 78.8126
R280 VP.n68 VP.n66 62.5827
R281 VP.n73 VP.n14 54.0911
R282 VP.n108 VP.n2 54.0911
R283 VP.n58 VP.n19 54.0911
R284 VP.n84 VP.n10 52.1486
R285 VP.n99 VP.n6 52.1486
R286 VP.n49 VP.n23 52.1486
R287 VP.n34 VP.n27 52.1486
R288 VP.n30 VP.n29 50.6338
R289 VP.n88 VP.n10 28.8382
R290 VP.n95 VP.n6 28.8382
R291 VP.n45 VP.n23 28.8382
R292 VP.n38 VP.n27 28.8382
R293 VP.n73 VP.n72 26.8957
R294 VP.n112 VP.n2 26.8957
R295 VP.n62 VP.n19 26.8957
R296 VP.n71 VP.n16 24.4675
R297 VP.n72 VP.n71 24.4675
R298 VP.n77 VP.n14 24.4675
R299 VP.n78 VP.n77 24.4675
R300 VP.n79 VP.n78 24.4675
R301 VP.n83 VP.n82 24.4675
R302 VP.n84 VP.n83 24.4675
R303 VP.n89 VP.n88 24.4675
R304 VP.n90 VP.n89 24.4675
R305 VP.n94 VP.n93 24.4675
R306 VP.n95 VP.n94 24.4675
R307 VP.n100 VP.n99 24.4675
R308 VP.n102 VP.n100 24.4675
R309 VP.n106 VP.n4 24.4675
R310 VP.n107 VP.n106 24.4675
R311 VP.n108 VP.n107 24.4675
R312 VP.n113 VP.n112 24.4675
R313 VP.n114 VP.n113 24.4675
R314 VP.n63 VP.n62 24.4675
R315 VP.n64 VP.n63 24.4675
R316 VP.n50 VP.n49 24.4675
R317 VP.n52 VP.n50 24.4675
R318 VP.n56 VP.n21 24.4675
R319 VP.n57 VP.n56 24.4675
R320 VP.n58 VP.n57 24.4675
R321 VP.n39 VP.n38 24.4675
R322 VP.n40 VP.n39 24.4675
R323 VP.n44 VP.n43 24.4675
R324 VP.n45 VP.n44 24.4675
R325 VP.n33 VP.n32 24.4675
R326 VP.n34 VP.n33 24.4675
R327 VP.n82 VP.n12 23.9782
R328 VP.n102 VP.n101 23.9782
R329 VP.n52 VP.n51 23.9782
R330 VP.n32 VP.n29 23.9782
R331 VP.n90 VP.n8 12.234
R332 VP.n93 VP.n8 12.234
R333 VP.n40 VP.n25 12.234
R334 VP.n43 VP.n25 12.234
R335 VP.n67 VP.n16 11.2553
R336 VP.n114 VP.n0 11.2553
R337 VP.n64 VP.n17 11.2553
R338 VP.n31 VP.n30 3.11118
R339 VP.n79 VP.n12 0.48984
R340 VP.n101 VP.n4 0.48984
R341 VP.n51 VP.n21 0.48984
R342 VP.n66 VP.n65 0.354971
R343 VP.n69 VP.n68 0.354971
R344 VP.n116 VP.n115 0.354971
R345 VP VP.n116 0.26696
R346 VP.n31 VP.n28 0.189894
R347 VP.n35 VP.n28 0.189894
R348 VP.n36 VP.n35 0.189894
R349 VP.n37 VP.n36 0.189894
R350 VP.n37 VP.n26 0.189894
R351 VP.n41 VP.n26 0.189894
R352 VP.n42 VP.n41 0.189894
R353 VP.n42 VP.n24 0.189894
R354 VP.n46 VP.n24 0.189894
R355 VP.n47 VP.n46 0.189894
R356 VP.n48 VP.n47 0.189894
R357 VP.n48 VP.n22 0.189894
R358 VP.n53 VP.n22 0.189894
R359 VP.n54 VP.n53 0.189894
R360 VP.n55 VP.n54 0.189894
R361 VP.n55 VP.n20 0.189894
R362 VP.n59 VP.n20 0.189894
R363 VP.n60 VP.n59 0.189894
R364 VP.n61 VP.n60 0.189894
R365 VP.n61 VP.n18 0.189894
R366 VP.n65 VP.n18 0.189894
R367 VP.n70 VP.n69 0.189894
R368 VP.n70 VP.n15 0.189894
R369 VP.n74 VP.n15 0.189894
R370 VP.n75 VP.n74 0.189894
R371 VP.n76 VP.n75 0.189894
R372 VP.n76 VP.n13 0.189894
R373 VP.n80 VP.n13 0.189894
R374 VP.n81 VP.n80 0.189894
R375 VP.n81 VP.n11 0.189894
R376 VP.n85 VP.n11 0.189894
R377 VP.n86 VP.n85 0.189894
R378 VP.n87 VP.n86 0.189894
R379 VP.n87 VP.n9 0.189894
R380 VP.n91 VP.n9 0.189894
R381 VP.n92 VP.n91 0.189894
R382 VP.n92 VP.n7 0.189894
R383 VP.n96 VP.n7 0.189894
R384 VP.n97 VP.n96 0.189894
R385 VP.n98 VP.n97 0.189894
R386 VP.n98 VP.n5 0.189894
R387 VP.n103 VP.n5 0.189894
R388 VP.n104 VP.n103 0.189894
R389 VP.n105 VP.n104 0.189894
R390 VP.n105 VP.n3 0.189894
R391 VP.n109 VP.n3 0.189894
R392 VP.n110 VP.n109 0.189894
R393 VP.n111 VP.n110 0.189894
R394 VP.n111 VP.n1 0.189894
R395 VP.n115 VP.n1 0.189894
R396 VDD1.n1 VDD1.t9 72.9252
R397 VDD1.n3 VDD1.t6 72.9251
R398 VDD1.n5 VDD1.n4 70.3132
R399 VDD1.n1 VDD1.n0 67.9507
R400 VDD1.n7 VDD1.n6 67.9505
R401 VDD1.n3 VDD1.n2 67.9505
R402 VDD1.n7 VDD1.n5 57.2337
R403 VDD1 VDD1.n7 2.36041
R404 VDD1.n6 VDD1.t2 1.7509
R405 VDD1.n6 VDD1.t8 1.7509
R406 VDD1.n0 VDD1.t7 1.7509
R407 VDD1.n0 VDD1.t4 1.7509
R408 VDD1.n4 VDD1.t3 1.7509
R409 VDD1.n4 VDD1.t0 1.7509
R410 VDD1.n2 VDD1.t5 1.7509
R411 VDD1.n2 VDD1.t1 1.7509
R412 VDD1 VDD1.n1 0.864724
R413 VDD1.n5 VDD1.n3 0.751188
R414 B.n822 B.n821 585
R415 B.n823 B.n108 585
R416 B.n825 B.n824 585
R417 B.n826 B.n107 585
R418 B.n828 B.n827 585
R419 B.n829 B.n106 585
R420 B.n831 B.n830 585
R421 B.n832 B.n105 585
R422 B.n834 B.n833 585
R423 B.n835 B.n104 585
R424 B.n837 B.n836 585
R425 B.n838 B.n103 585
R426 B.n840 B.n839 585
R427 B.n841 B.n102 585
R428 B.n843 B.n842 585
R429 B.n844 B.n101 585
R430 B.n846 B.n845 585
R431 B.n847 B.n100 585
R432 B.n849 B.n848 585
R433 B.n850 B.n99 585
R434 B.n852 B.n851 585
R435 B.n853 B.n98 585
R436 B.n855 B.n854 585
R437 B.n856 B.n97 585
R438 B.n858 B.n857 585
R439 B.n859 B.n96 585
R440 B.n861 B.n860 585
R441 B.n862 B.n95 585
R442 B.n864 B.n863 585
R443 B.n865 B.n94 585
R444 B.n867 B.n866 585
R445 B.n868 B.n93 585
R446 B.n870 B.n869 585
R447 B.n871 B.n92 585
R448 B.n873 B.n872 585
R449 B.n874 B.n91 585
R450 B.n876 B.n875 585
R451 B.n877 B.n90 585
R452 B.n879 B.n878 585
R453 B.n880 B.n89 585
R454 B.n882 B.n881 585
R455 B.n883 B.n88 585
R456 B.n885 B.n884 585
R457 B.n886 B.n87 585
R458 B.n888 B.n887 585
R459 B.n889 B.n86 585
R460 B.n891 B.n890 585
R461 B.n892 B.n85 585
R462 B.n894 B.n893 585
R463 B.n895 B.n84 585
R464 B.n897 B.n896 585
R465 B.n898 B.n83 585
R466 B.n900 B.n899 585
R467 B.n901 B.n82 585
R468 B.n903 B.n902 585
R469 B.n904 B.n81 585
R470 B.n906 B.n905 585
R471 B.n907 B.n80 585
R472 B.n909 B.n908 585
R473 B.n910 B.n79 585
R474 B.n912 B.n911 585
R475 B.n914 B.n913 585
R476 B.n915 B.n75 585
R477 B.n917 B.n916 585
R478 B.n918 B.n74 585
R479 B.n920 B.n919 585
R480 B.n921 B.n73 585
R481 B.n923 B.n922 585
R482 B.n924 B.n72 585
R483 B.n926 B.n925 585
R484 B.n928 B.n69 585
R485 B.n930 B.n929 585
R486 B.n931 B.n68 585
R487 B.n933 B.n932 585
R488 B.n934 B.n67 585
R489 B.n936 B.n935 585
R490 B.n937 B.n66 585
R491 B.n939 B.n938 585
R492 B.n940 B.n65 585
R493 B.n942 B.n941 585
R494 B.n943 B.n64 585
R495 B.n945 B.n944 585
R496 B.n946 B.n63 585
R497 B.n948 B.n947 585
R498 B.n949 B.n62 585
R499 B.n951 B.n950 585
R500 B.n952 B.n61 585
R501 B.n954 B.n953 585
R502 B.n955 B.n60 585
R503 B.n957 B.n956 585
R504 B.n958 B.n59 585
R505 B.n960 B.n959 585
R506 B.n961 B.n58 585
R507 B.n963 B.n962 585
R508 B.n964 B.n57 585
R509 B.n966 B.n965 585
R510 B.n967 B.n56 585
R511 B.n969 B.n968 585
R512 B.n970 B.n55 585
R513 B.n972 B.n971 585
R514 B.n973 B.n54 585
R515 B.n975 B.n974 585
R516 B.n976 B.n53 585
R517 B.n978 B.n977 585
R518 B.n979 B.n52 585
R519 B.n981 B.n980 585
R520 B.n982 B.n51 585
R521 B.n984 B.n983 585
R522 B.n985 B.n50 585
R523 B.n987 B.n986 585
R524 B.n988 B.n49 585
R525 B.n990 B.n989 585
R526 B.n991 B.n48 585
R527 B.n993 B.n992 585
R528 B.n994 B.n47 585
R529 B.n996 B.n995 585
R530 B.n997 B.n46 585
R531 B.n999 B.n998 585
R532 B.n1000 B.n45 585
R533 B.n1002 B.n1001 585
R534 B.n1003 B.n44 585
R535 B.n1005 B.n1004 585
R536 B.n1006 B.n43 585
R537 B.n1008 B.n1007 585
R538 B.n1009 B.n42 585
R539 B.n1011 B.n1010 585
R540 B.n1012 B.n41 585
R541 B.n1014 B.n1013 585
R542 B.n1015 B.n40 585
R543 B.n1017 B.n1016 585
R544 B.n1018 B.n39 585
R545 B.n820 B.n109 585
R546 B.n819 B.n818 585
R547 B.n817 B.n110 585
R548 B.n816 B.n815 585
R549 B.n814 B.n111 585
R550 B.n813 B.n812 585
R551 B.n811 B.n112 585
R552 B.n810 B.n809 585
R553 B.n808 B.n113 585
R554 B.n807 B.n806 585
R555 B.n805 B.n114 585
R556 B.n804 B.n803 585
R557 B.n802 B.n115 585
R558 B.n801 B.n800 585
R559 B.n799 B.n116 585
R560 B.n798 B.n797 585
R561 B.n796 B.n117 585
R562 B.n795 B.n794 585
R563 B.n793 B.n118 585
R564 B.n792 B.n791 585
R565 B.n790 B.n119 585
R566 B.n789 B.n788 585
R567 B.n787 B.n120 585
R568 B.n786 B.n785 585
R569 B.n784 B.n121 585
R570 B.n783 B.n782 585
R571 B.n781 B.n122 585
R572 B.n780 B.n779 585
R573 B.n778 B.n123 585
R574 B.n777 B.n776 585
R575 B.n775 B.n124 585
R576 B.n774 B.n773 585
R577 B.n772 B.n125 585
R578 B.n771 B.n770 585
R579 B.n769 B.n126 585
R580 B.n768 B.n767 585
R581 B.n766 B.n127 585
R582 B.n765 B.n764 585
R583 B.n763 B.n128 585
R584 B.n762 B.n761 585
R585 B.n760 B.n129 585
R586 B.n759 B.n758 585
R587 B.n757 B.n130 585
R588 B.n756 B.n755 585
R589 B.n754 B.n131 585
R590 B.n753 B.n752 585
R591 B.n751 B.n132 585
R592 B.n750 B.n749 585
R593 B.n748 B.n133 585
R594 B.n747 B.n746 585
R595 B.n745 B.n134 585
R596 B.n744 B.n743 585
R597 B.n742 B.n135 585
R598 B.n741 B.n740 585
R599 B.n739 B.n136 585
R600 B.n738 B.n737 585
R601 B.n736 B.n137 585
R602 B.n735 B.n734 585
R603 B.n733 B.n138 585
R604 B.n732 B.n731 585
R605 B.n730 B.n139 585
R606 B.n729 B.n728 585
R607 B.n727 B.n140 585
R608 B.n726 B.n725 585
R609 B.n724 B.n141 585
R610 B.n723 B.n722 585
R611 B.n721 B.n142 585
R612 B.n720 B.n719 585
R613 B.n718 B.n143 585
R614 B.n717 B.n716 585
R615 B.n715 B.n144 585
R616 B.n714 B.n713 585
R617 B.n712 B.n145 585
R618 B.n711 B.n710 585
R619 B.n709 B.n146 585
R620 B.n708 B.n707 585
R621 B.n706 B.n147 585
R622 B.n705 B.n704 585
R623 B.n703 B.n148 585
R624 B.n702 B.n701 585
R625 B.n700 B.n149 585
R626 B.n699 B.n698 585
R627 B.n697 B.n150 585
R628 B.n696 B.n695 585
R629 B.n694 B.n151 585
R630 B.n693 B.n692 585
R631 B.n691 B.n152 585
R632 B.n690 B.n689 585
R633 B.n688 B.n153 585
R634 B.n687 B.n686 585
R635 B.n685 B.n154 585
R636 B.n684 B.n683 585
R637 B.n682 B.n155 585
R638 B.n681 B.n680 585
R639 B.n679 B.n156 585
R640 B.n678 B.n677 585
R641 B.n676 B.n157 585
R642 B.n675 B.n674 585
R643 B.n673 B.n158 585
R644 B.n672 B.n671 585
R645 B.n670 B.n159 585
R646 B.n669 B.n668 585
R647 B.n667 B.n160 585
R648 B.n666 B.n665 585
R649 B.n664 B.n161 585
R650 B.n663 B.n662 585
R651 B.n661 B.n162 585
R652 B.n660 B.n659 585
R653 B.n658 B.n163 585
R654 B.n657 B.n656 585
R655 B.n655 B.n164 585
R656 B.n654 B.n653 585
R657 B.n652 B.n165 585
R658 B.n651 B.n650 585
R659 B.n649 B.n166 585
R660 B.n648 B.n647 585
R661 B.n646 B.n167 585
R662 B.n645 B.n644 585
R663 B.n643 B.n168 585
R664 B.n642 B.n641 585
R665 B.n640 B.n169 585
R666 B.n639 B.n638 585
R667 B.n637 B.n170 585
R668 B.n636 B.n635 585
R669 B.n634 B.n171 585
R670 B.n633 B.n632 585
R671 B.n631 B.n172 585
R672 B.n630 B.n629 585
R673 B.n628 B.n173 585
R674 B.n627 B.n626 585
R675 B.n625 B.n174 585
R676 B.n624 B.n623 585
R677 B.n622 B.n175 585
R678 B.n621 B.n620 585
R679 B.n619 B.n176 585
R680 B.n618 B.n617 585
R681 B.n616 B.n177 585
R682 B.n615 B.n614 585
R683 B.n613 B.n178 585
R684 B.n612 B.n611 585
R685 B.n610 B.n179 585
R686 B.n609 B.n608 585
R687 B.n607 B.n180 585
R688 B.n606 B.n605 585
R689 B.n604 B.n181 585
R690 B.n603 B.n602 585
R691 B.n601 B.n182 585
R692 B.n600 B.n599 585
R693 B.n598 B.n183 585
R694 B.n400 B.n253 585
R695 B.n402 B.n401 585
R696 B.n403 B.n252 585
R697 B.n405 B.n404 585
R698 B.n406 B.n251 585
R699 B.n408 B.n407 585
R700 B.n409 B.n250 585
R701 B.n411 B.n410 585
R702 B.n412 B.n249 585
R703 B.n414 B.n413 585
R704 B.n415 B.n248 585
R705 B.n417 B.n416 585
R706 B.n418 B.n247 585
R707 B.n420 B.n419 585
R708 B.n421 B.n246 585
R709 B.n423 B.n422 585
R710 B.n424 B.n245 585
R711 B.n426 B.n425 585
R712 B.n427 B.n244 585
R713 B.n429 B.n428 585
R714 B.n430 B.n243 585
R715 B.n432 B.n431 585
R716 B.n433 B.n242 585
R717 B.n435 B.n434 585
R718 B.n436 B.n241 585
R719 B.n438 B.n437 585
R720 B.n439 B.n240 585
R721 B.n441 B.n440 585
R722 B.n442 B.n239 585
R723 B.n444 B.n443 585
R724 B.n445 B.n238 585
R725 B.n447 B.n446 585
R726 B.n448 B.n237 585
R727 B.n450 B.n449 585
R728 B.n451 B.n236 585
R729 B.n453 B.n452 585
R730 B.n454 B.n235 585
R731 B.n456 B.n455 585
R732 B.n457 B.n234 585
R733 B.n459 B.n458 585
R734 B.n460 B.n233 585
R735 B.n462 B.n461 585
R736 B.n463 B.n232 585
R737 B.n465 B.n464 585
R738 B.n466 B.n231 585
R739 B.n468 B.n467 585
R740 B.n469 B.n230 585
R741 B.n471 B.n470 585
R742 B.n472 B.n229 585
R743 B.n474 B.n473 585
R744 B.n475 B.n228 585
R745 B.n477 B.n476 585
R746 B.n478 B.n227 585
R747 B.n480 B.n479 585
R748 B.n481 B.n226 585
R749 B.n483 B.n482 585
R750 B.n484 B.n225 585
R751 B.n486 B.n485 585
R752 B.n487 B.n224 585
R753 B.n489 B.n488 585
R754 B.n490 B.n221 585
R755 B.n493 B.n492 585
R756 B.n494 B.n220 585
R757 B.n496 B.n495 585
R758 B.n497 B.n219 585
R759 B.n499 B.n498 585
R760 B.n500 B.n218 585
R761 B.n502 B.n501 585
R762 B.n503 B.n217 585
R763 B.n505 B.n504 585
R764 B.n507 B.n506 585
R765 B.n508 B.n213 585
R766 B.n510 B.n509 585
R767 B.n511 B.n212 585
R768 B.n513 B.n512 585
R769 B.n514 B.n211 585
R770 B.n516 B.n515 585
R771 B.n517 B.n210 585
R772 B.n519 B.n518 585
R773 B.n520 B.n209 585
R774 B.n522 B.n521 585
R775 B.n523 B.n208 585
R776 B.n525 B.n524 585
R777 B.n526 B.n207 585
R778 B.n528 B.n527 585
R779 B.n529 B.n206 585
R780 B.n531 B.n530 585
R781 B.n532 B.n205 585
R782 B.n534 B.n533 585
R783 B.n535 B.n204 585
R784 B.n537 B.n536 585
R785 B.n538 B.n203 585
R786 B.n540 B.n539 585
R787 B.n541 B.n202 585
R788 B.n543 B.n542 585
R789 B.n544 B.n201 585
R790 B.n546 B.n545 585
R791 B.n547 B.n200 585
R792 B.n549 B.n548 585
R793 B.n550 B.n199 585
R794 B.n552 B.n551 585
R795 B.n553 B.n198 585
R796 B.n555 B.n554 585
R797 B.n556 B.n197 585
R798 B.n558 B.n557 585
R799 B.n559 B.n196 585
R800 B.n561 B.n560 585
R801 B.n562 B.n195 585
R802 B.n564 B.n563 585
R803 B.n565 B.n194 585
R804 B.n567 B.n566 585
R805 B.n568 B.n193 585
R806 B.n570 B.n569 585
R807 B.n571 B.n192 585
R808 B.n573 B.n572 585
R809 B.n574 B.n191 585
R810 B.n576 B.n575 585
R811 B.n577 B.n190 585
R812 B.n579 B.n578 585
R813 B.n580 B.n189 585
R814 B.n582 B.n581 585
R815 B.n583 B.n188 585
R816 B.n585 B.n584 585
R817 B.n586 B.n187 585
R818 B.n588 B.n587 585
R819 B.n589 B.n186 585
R820 B.n591 B.n590 585
R821 B.n592 B.n185 585
R822 B.n594 B.n593 585
R823 B.n595 B.n184 585
R824 B.n597 B.n596 585
R825 B.n399 B.n398 585
R826 B.n397 B.n254 585
R827 B.n396 B.n395 585
R828 B.n394 B.n255 585
R829 B.n393 B.n392 585
R830 B.n391 B.n256 585
R831 B.n390 B.n389 585
R832 B.n388 B.n257 585
R833 B.n387 B.n386 585
R834 B.n385 B.n258 585
R835 B.n384 B.n383 585
R836 B.n382 B.n259 585
R837 B.n381 B.n380 585
R838 B.n379 B.n260 585
R839 B.n378 B.n377 585
R840 B.n376 B.n261 585
R841 B.n375 B.n374 585
R842 B.n373 B.n262 585
R843 B.n372 B.n371 585
R844 B.n370 B.n263 585
R845 B.n369 B.n368 585
R846 B.n367 B.n264 585
R847 B.n366 B.n365 585
R848 B.n364 B.n265 585
R849 B.n363 B.n362 585
R850 B.n361 B.n266 585
R851 B.n360 B.n359 585
R852 B.n358 B.n267 585
R853 B.n357 B.n356 585
R854 B.n355 B.n268 585
R855 B.n354 B.n353 585
R856 B.n352 B.n269 585
R857 B.n351 B.n350 585
R858 B.n349 B.n270 585
R859 B.n348 B.n347 585
R860 B.n346 B.n271 585
R861 B.n345 B.n344 585
R862 B.n343 B.n272 585
R863 B.n342 B.n341 585
R864 B.n340 B.n273 585
R865 B.n339 B.n338 585
R866 B.n337 B.n274 585
R867 B.n336 B.n335 585
R868 B.n334 B.n275 585
R869 B.n333 B.n332 585
R870 B.n331 B.n276 585
R871 B.n330 B.n329 585
R872 B.n328 B.n277 585
R873 B.n327 B.n326 585
R874 B.n325 B.n278 585
R875 B.n324 B.n323 585
R876 B.n322 B.n279 585
R877 B.n321 B.n320 585
R878 B.n319 B.n280 585
R879 B.n318 B.n317 585
R880 B.n316 B.n281 585
R881 B.n315 B.n314 585
R882 B.n313 B.n282 585
R883 B.n312 B.n311 585
R884 B.n310 B.n283 585
R885 B.n309 B.n308 585
R886 B.n307 B.n284 585
R887 B.n306 B.n305 585
R888 B.n304 B.n285 585
R889 B.n303 B.n302 585
R890 B.n301 B.n286 585
R891 B.n300 B.n299 585
R892 B.n298 B.n287 585
R893 B.n297 B.n296 585
R894 B.n295 B.n288 585
R895 B.n294 B.n293 585
R896 B.n292 B.n289 585
R897 B.n291 B.n290 585
R898 B.n2 B.n0 585
R899 B.n1129 B.n1 585
R900 B.n1128 B.n1127 585
R901 B.n1126 B.n3 585
R902 B.n1125 B.n1124 585
R903 B.n1123 B.n4 585
R904 B.n1122 B.n1121 585
R905 B.n1120 B.n5 585
R906 B.n1119 B.n1118 585
R907 B.n1117 B.n6 585
R908 B.n1116 B.n1115 585
R909 B.n1114 B.n7 585
R910 B.n1113 B.n1112 585
R911 B.n1111 B.n8 585
R912 B.n1110 B.n1109 585
R913 B.n1108 B.n9 585
R914 B.n1107 B.n1106 585
R915 B.n1105 B.n10 585
R916 B.n1104 B.n1103 585
R917 B.n1102 B.n11 585
R918 B.n1101 B.n1100 585
R919 B.n1099 B.n12 585
R920 B.n1098 B.n1097 585
R921 B.n1096 B.n13 585
R922 B.n1095 B.n1094 585
R923 B.n1093 B.n14 585
R924 B.n1092 B.n1091 585
R925 B.n1090 B.n15 585
R926 B.n1089 B.n1088 585
R927 B.n1087 B.n16 585
R928 B.n1086 B.n1085 585
R929 B.n1084 B.n17 585
R930 B.n1083 B.n1082 585
R931 B.n1081 B.n18 585
R932 B.n1080 B.n1079 585
R933 B.n1078 B.n19 585
R934 B.n1077 B.n1076 585
R935 B.n1075 B.n20 585
R936 B.n1074 B.n1073 585
R937 B.n1072 B.n21 585
R938 B.n1071 B.n1070 585
R939 B.n1069 B.n22 585
R940 B.n1068 B.n1067 585
R941 B.n1066 B.n23 585
R942 B.n1065 B.n1064 585
R943 B.n1063 B.n24 585
R944 B.n1062 B.n1061 585
R945 B.n1060 B.n25 585
R946 B.n1059 B.n1058 585
R947 B.n1057 B.n26 585
R948 B.n1056 B.n1055 585
R949 B.n1054 B.n27 585
R950 B.n1053 B.n1052 585
R951 B.n1051 B.n28 585
R952 B.n1050 B.n1049 585
R953 B.n1048 B.n29 585
R954 B.n1047 B.n1046 585
R955 B.n1045 B.n30 585
R956 B.n1044 B.n1043 585
R957 B.n1042 B.n31 585
R958 B.n1041 B.n1040 585
R959 B.n1039 B.n32 585
R960 B.n1038 B.n1037 585
R961 B.n1036 B.n33 585
R962 B.n1035 B.n1034 585
R963 B.n1033 B.n34 585
R964 B.n1032 B.n1031 585
R965 B.n1030 B.n35 585
R966 B.n1029 B.n1028 585
R967 B.n1027 B.n36 585
R968 B.n1026 B.n1025 585
R969 B.n1024 B.n37 585
R970 B.n1023 B.n1022 585
R971 B.n1021 B.n38 585
R972 B.n1020 B.n1019 585
R973 B.n1131 B.n1130 585
R974 B.n398 B.n253 554.963
R975 B.n1020 B.n39 554.963
R976 B.n596 B.n183 554.963
R977 B.n822 B.n109 554.963
R978 B.n214 B.t9 340.253
R979 B.n222 B.t6 340.253
R980 B.n70 B.t0 340.253
R981 B.n76 B.t3 340.253
R982 B.n214 B.t11 182.756
R983 B.n76 B.t4 182.756
R984 B.n222 B.t8 182.732
R985 B.n70 B.t1 182.732
R986 B.n398 B.n397 163.367
R987 B.n397 B.n396 163.367
R988 B.n396 B.n255 163.367
R989 B.n392 B.n255 163.367
R990 B.n392 B.n391 163.367
R991 B.n391 B.n390 163.367
R992 B.n390 B.n257 163.367
R993 B.n386 B.n257 163.367
R994 B.n386 B.n385 163.367
R995 B.n385 B.n384 163.367
R996 B.n384 B.n259 163.367
R997 B.n380 B.n259 163.367
R998 B.n380 B.n379 163.367
R999 B.n379 B.n378 163.367
R1000 B.n378 B.n261 163.367
R1001 B.n374 B.n261 163.367
R1002 B.n374 B.n373 163.367
R1003 B.n373 B.n372 163.367
R1004 B.n372 B.n263 163.367
R1005 B.n368 B.n263 163.367
R1006 B.n368 B.n367 163.367
R1007 B.n367 B.n366 163.367
R1008 B.n366 B.n265 163.367
R1009 B.n362 B.n265 163.367
R1010 B.n362 B.n361 163.367
R1011 B.n361 B.n360 163.367
R1012 B.n360 B.n267 163.367
R1013 B.n356 B.n267 163.367
R1014 B.n356 B.n355 163.367
R1015 B.n355 B.n354 163.367
R1016 B.n354 B.n269 163.367
R1017 B.n350 B.n269 163.367
R1018 B.n350 B.n349 163.367
R1019 B.n349 B.n348 163.367
R1020 B.n348 B.n271 163.367
R1021 B.n344 B.n271 163.367
R1022 B.n344 B.n343 163.367
R1023 B.n343 B.n342 163.367
R1024 B.n342 B.n273 163.367
R1025 B.n338 B.n273 163.367
R1026 B.n338 B.n337 163.367
R1027 B.n337 B.n336 163.367
R1028 B.n336 B.n275 163.367
R1029 B.n332 B.n275 163.367
R1030 B.n332 B.n331 163.367
R1031 B.n331 B.n330 163.367
R1032 B.n330 B.n277 163.367
R1033 B.n326 B.n277 163.367
R1034 B.n326 B.n325 163.367
R1035 B.n325 B.n324 163.367
R1036 B.n324 B.n279 163.367
R1037 B.n320 B.n279 163.367
R1038 B.n320 B.n319 163.367
R1039 B.n319 B.n318 163.367
R1040 B.n318 B.n281 163.367
R1041 B.n314 B.n281 163.367
R1042 B.n314 B.n313 163.367
R1043 B.n313 B.n312 163.367
R1044 B.n312 B.n283 163.367
R1045 B.n308 B.n283 163.367
R1046 B.n308 B.n307 163.367
R1047 B.n307 B.n306 163.367
R1048 B.n306 B.n285 163.367
R1049 B.n302 B.n285 163.367
R1050 B.n302 B.n301 163.367
R1051 B.n301 B.n300 163.367
R1052 B.n300 B.n287 163.367
R1053 B.n296 B.n287 163.367
R1054 B.n296 B.n295 163.367
R1055 B.n295 B.n294 163.367
R1056 B.n294 B.n289 163.367
R1057 B.n290 B.n289 163.367
R1058 B.n290 B.n2 163.367
R1059 B.n1130 B.n2 163.367
R1060 B.n1130 B.n1129 163.367
R1061 B.n1129 B.n1128 163.367
R1062 B.n1128 B.n3 163.367
R1063 B.n1124 B.n3 163.367
R1064 B.n1124 B.n1123 163.367
R1065 B.n1123 B.n1122 163.367
R1066 B.n1122 B.n5 163.367
R1067 B.n1118 B.n5 163.367
R1068 B.n1118 B.n1117 163.367
R1069 B.n1117 B.n1116 163.367
R1070 B.n1116 B.n7 163.367
R1071 B.n1112 B.n7 163.367
R1072 B.n1112 B.n1111 163.367
R1073 B.n1111 B.n1110 163.367
R1074 B.n1110 B.n9 163.367
R1075 B.n1106 B.n9 163.367
R1076 B.n1106 B.n1105 163.367
R1077 B.n1105 B.n1104 163.367
R1078 B.n1104 B.n11 163.367
R1079 B.n1100 B.n11 163.367
R1080 B.n1100 B.n1099 163.367
R1081 B.n1099 B.n1098 163.367
R1082 B.n1098 B.n13 163.367
R1083 B.n1094 B.n13 163.367
R1084 B.n1094 B.n1093 163.367
R1085 B.n1093 B.n1092 163.367
R1086 B.n1092 B.n15 163.367
R1087 B.n1088 B.n15 163.367
R1088 B.n1088 B.n1087 163.367
R1089 B.n1087 B.n1086 163.367
R1090 B.n1086 B.n17 163.367
R1091 B.n1082 B.n17 163.367
R1092 B.n1082 B.n1081 163.367
R1093 B.n1081 B.n1080 163.367
R1094 B.n1080 B.n19 163.367
R1095 B.n1076 B.n19 163.367
R1096 B.n1076 B.n1075 163.367
R1097 B.n1075 B.n1074 163.367
R1098 B.n1074 B.n21 163.367
R1099 B.n1070 B.n21 163.367
R1100 B.n1070 B.n1069 163.367
R1101 B.n1069 B.n1068 163.367
R1102 B.n1068 B.n23 163.367
R1103 B.n1064 B.n23 163.367
R1104 B.n1064 B.n1063 163.367
R1105 B.n1063 B.n1062 163.367
R1106 B.n1062 B.n25 163.367
R1107 B.n1058 B.n25 163.367
R1108 B.n1058 B.n1057 163.367
R1109 B.n1057 B.n1056 163.367
R1110 B.n1056 B.n27 163.367
R1111 B.n1052 B.n27 163.367
R1112 B.n1052 B.n1051 163.367
R1113 B.n1051 B.n1050 163.367
R1114 B.n1050 B.n29 163.367
R1115 B.n1046 B.n29 163.367
R1116 B.n1046 B.n1045 163.367
R1117 B.n1045 B.n1044 163.367
R1118 B.n1044 B.n31 163.367
R1119 B.n1040 B.n31 163.367
R1120 B.n1040 B.n1039 163.367
R1121 B.n1039 B.n1038 163.367
R1122 B.n1038 B.n33 163.367
R1123 B.n1034 B.n33 163.367
R1124 B.n1034 B.n1033 163.367
R1125 B.n1033 B.n1032 163.367
R1126 B.n1032 B.n35 163.367
R1127 B.n1028 B.n35 163.367
R1128 B.n1028 B.n1027 163.367
R1129 B.n1027 B.n1026 163.367
R1130 B.n1026 B.n37 163.367
R1131 B.n1022 B.n37 163.367
R1132 B.n1022 B.n1021 163.367
R1133 B.n1021 B.n1020 163.367
R1134 B.n402 B.n253 163.367
R1135 B.n403 B.n402 163.367
R1136 B.n404 B.n403 163.367
R1137 B.n404 B.n251 163.367
R1138 B.n408 B.n251 163.367
R1139 B.n409 B.n408 163.367
R1140 B.n410 B.n409 163.367
R1141 B.n410 B.n249 163.367
R1142 B.n414 B.n249 163.367
R1143 B.n415 B.n414 163.367
R1144 B.n416 B.n415 163.367
R1145 B.n416 B.n247 163.367
R1146 B.n420 B.n247 163.367
R1147 B.n421 B.n420 163.367
R1148 B.n422 B.n421 163.367
R1149 B.n422 B.n245 163.367
R1150 B.n426 B.n245 163.367
R1151 B.n427 B.n426 163.367
R1152 B.n428 B.n427 163.367
R1153 B.n428 B.n243 163.367
R1154 B.n432 B.n243 163.367
R1155 B.n433 B.n432 163.367
R1156 B.n434 B.n433 163.367
R1157 B.n434 B.n241 163.367
R1158 B.n438 B.n241 163.367
R1159 B.n439 B.n438 163.367
R1160 B.n440 B.n439 163.367
R1161 B.n440 B.n239 163.367
R1162 B.n444 B.n239 163.367
R1163 B.n445 B.n444 163.367
R1164 B.n446 B.n445 163.367
R1165 B.n446 B.n237 163.367
R1166 B.n450 B.n237 163.367
R1167 B.n451 B.n450 163.367
R1168 B.n452 B.n451 163.367
R1169 B.n452 B.n235 163.367
R1170 B.n456 B.n235 163.367
R1171 B.n457 B.n456 163.367
R1172 B.n458 B.n457 163.367
R1173 B.n458 B.n233 163.367
R1174 B.n462 B.n233 163.367
R1175 B.n463 B.n462 163.367
R1176 B.n464 B.n463 163.367
R1177 B.n464 B.n231 163.367
R1178 B.n468 B.n231 163.367
R1179 B.n469 B.n468 163.367
R1180 B.n470 B.n469 163.367
R1181 B.n470 B.n229 163.367
R1182 B.n474 B.n229 163.367
R1183 B.n475 B.n474 163.367
R1184 B.n476 B.n475 163.367
R1185 B.n476 B.n227 163.367
R1186 B.n480 B.n227 163.367
R1187 B.n481 B.n480 163.367
R1188 B.n482 B.n481 163.367
R1189 B.n482 B.n225 163.367
R1190 B.n486 B.n225 163.367
R1191 B.n487 B.n486 163.367
R1192 B.n488 B.n487 163.367
R1193 B.n488 B.n221 163.367
R1194 B.n493 B.n221 163.367
R1195 B.n494 B.n493 163.367
R1196 B.n495 B.n494 163.367
R1197 B.n495 B.n219 163.367
R1198 B.n499 B.n219 163.367
R1199 B.n500 B.n499 163.367
R1200 B.n501 B.n500 163.367
R1201 B.n501 B.n217 163.367
R1202 B.n505 B.n217 163.367
R1203 B.n506 B.n505 163.367
R1204 B.n506 B.n213 163.367
R1205 B.n510 B.n213 163.367
R1206 B.n511 B.n510 163.367
R1207 B.n512 B.n511 163.367
R1208 B.n512 B.n211 163.367
R1209 B.n516 B.n211 163.367
R1210 B.n517 B.n516 163.367
R1211 B.n518 B.n517 163.367
R1212 B.n518 B.n209 163.367
R1213 B.n522 B.n209 163.367
R1214 B.n523 B.n522 163.367
R1215 B.n524 B.n523 163.367
R1216 B.n524 B.n207 163.367
R1217 B.n528 B.n207 163.367
R1218 B.n529 B.n528 163.367
R1219 B.n530 B.n529 163.367
R1220 B.n530 B.n205 163.367
R1221 B.n534 B.n205 163.367
R1222 B.n535 B.n534 163.367
R1223 B.n536 B.n535 163.367
R1224 B.n536 B.n203 163.367
R1225 B.n540 B.n203 163.367
R1226 B.n541 B.n540 163.367
R1227 B.n542 B.n541 163.367
R1228 B.n542 B.n201 163.367
R1229 B.n546 B.n201 163.367
R1230 B.n547 B.n546 163.367
R1231 B.n548 B.n547 163.367
R1232 B.n548 B.n199 163.367
R1233 B.n552 B.n199 163.367
R1234 B.n553 B.n552 163.367
R1235 B.n554 B.n553 163.367
R1236 B.n554 B.n197 163.367
R1237 B.n558 B.n197 163.367
R1238 B.n559 B.n558 163.367
R1239 B.n560 B.n559 163.367
R1240 B.n560 B.n195 163.367
R1241 B.n564 B.n195 163.367
R1242 B.n565 B.n564 163.367
R1243 B.n566 B.n565 163.367
R1244 B.n566 B.n193 163.367
R1245 B.n570 B.n193 163.367
R1246 B.n571 B.n570 163.367
R1247 B.n572 B.n571 163.367
R1248 B.n572 B.n191 163.367
R1249 B.n576 B.n191 163.367
R1250 B.n577 B.n576 163.367
R1251 B.n578 B.n577 163.367
R1252 B.n578 B.n189 163.367
R1253 B.n582 B.n189 163.367
R1254 B.n583 B.n582 163.367
R1255 B.n584 B.n583 163.367
R1256 B.n584 B.n187 163.367
R1257 B.n588 B.n187 163.367
R1258 B.n589 B.n588 163.367
R1259 B.n590 B.n589 163.367
R1260 B.n590 B.n185 163.367
R1261 B.n594 B.n185 163.367
R1262 B.n595 B.n594 163.367
R1263 B.n596 B.n595 163.367
R1264 B.n600 B.n183 163.367
R1265 B.n601 B.n600 163.367
R1266 B.n602 B.n601 163.367
R1267 B.n602 B.n181 163.367
R1268 B.n606 B.n181 163.367
R1269 B.n607 B.n606 163.367
R1270 B.n608 B.n607 163.367
R1271 B.n608 B.n179 163.367
R1272 B.n612 B.n179 163.367
R1273 B.n613 B.n612 163.367
R1274 B.n614 B.n613 163.367
R1275 B.n614 B.n177 163.367
R1276 B.n618 B.n177 163.367
R1277 B.n619 B.n618 163.367
R1278 B.n620 B.n619 163.367
R1279 B.n620 B.n175 163.367
R1280 B.n624 B.n175 163.367
R1281 B.n625 B.n624 163.367
R1282 B.n626 B.n625 163.367
R1283 B.n626 B.n173 163.367
R1284 B.n630 B.n173 163.367
R1285 B.n631 B.n630 163.367
R1286 B.n632 B.n631 163.367
R1287 B.n632 B.n171 163.367
R1288 B.n636 B.n171 163.367
R1289 B.n637 B.n636 163.367
R1290 B.n638 B.n637 163.367
R1291 B.n638 B.n169 163.367
R1292 B.n642 B.n169 163.367
R1293 B.n643 B.n642 163.367
R1294 B.n644 B.n643 163.367
R1295 B.n644 B.n167 163.367
R1296 B.n648 B.n167 163.367
R1297 B.n649 B.n648 163.367
R1298 B.n650 B.n649 163.367
R1299 B.n650 B.n165 163.367
R1300 B.n654 B.n165 163.367
R1301 B.n655 B.n654 163.367
R1302 B.n656 B.n655 163.367
R1303 B.n656 B.n163 163.367
R1304 B.n660 B.n163 163.367
R1305 B.n661 B.n660 163.367
R1306 B.n662 B.n661 163.367
R1307 B.n662 B.n161 163.367
R1308 B.n666 B.n161 163.367
R1309 B.n667 B.n666 163.367
R1310 B.n668 B.n667 163.367
R1311 B.n668 B.n159 163.367
R1312 B.n672 B.n159 163.367
R1313 B.n673 B.n672 163.367
R1314 B.n674 B.n673 163.367
R1315 B.n674 B.n157 163.367
R1316 B.n678 B.n157 163.367
R1317 B.n679 B.n678 163.367
R1318 B.n680 B.n679 163.367
R1319 B.n680 B.n155 163.367
R1320 B.n684 B.n155 163.367
R1321 B.n685 B.n684 163.367
R1322 B.n686 B.n685 163.367
R1323 B.n686 B.n153 163.367
R1324 B.n690 B.n153 163.367
R1325 B.n691 B.n690 163.367
R1326 B.n692 B.n691 163.367
R1327 B.n692 B.n151 163.367
R1328 B.n696 B.n151 163.367
R1329 B.n697 B.n696 163.367
R1330 B.n698 B.n697 163.367
R1331 B.n698 B.n149 163.367
R1332 B.n702 B.n149 163.367
R1333 B.n703 B.n702 163.367
R1334 B.n704 B.n703 163.367
R1335 B.n704 B.n147 163.367
R1336 B.n708 B.n147 163.367
R1337 B.n709 B.n708 163.367
R1338 B.n710 B.n709 163.367
R1339 B.n710 B.n145 163.367
R1340 B.n714 B.n145 163.367
R1341 B.n715 B.n714 163.367
R1342 B.n716 B.n715 163.367
R1343 B.n716 B.n143 163.367
R1344 B.n720 B.n143 163.367
R1345 B.n721 B.n720 163.367
R1346 B.n722 B.n721 163.367
R1347 B.n722 B.n141 163.367
R1348 B.n726 B.n141 163.367
R1349 B.n727 B.n726 163.367
R1350 B.n728 B.n727 163.367
R1351 B.n728 B.n139 163.367
R1352 B.n732 B.n139 163.367
R1353 B.n733 B.n732 163.367
R1354 B.n734 B.n733 163.367
R1355 B.n734 B.n137 163.367
R1356 B.n738 B.n137 163.367
R1357 B.n739 B.n738 163.367
R1358 B.n740 B.n739 163.367
R1359 B.n740 B.n135 163.367
R1360 B.n744 B.n135 163.367
R1361 B.n745 B.n744 163.367
R1362 B.n746 B.n745 163.367
R1363 B.n746 B.n133 163.367
R1364 B.n750 B.n133 163.367
R1365 B.n751 B.n750 163.367
R1366 B.n752 B.n751 163.367
R1367 B.n752 B.n131 163.367
R1368 B.n756 B.n131 163.367
R1369 B.n757 B.n756 163.367
R1370 B.n758 B.n757 163.367
R1371 B.n758 B.n129 163.367
R1372 B.n762 B.n129 163.367
R1373 B.n763 B.n762 163.367
R1374 B.n764 B.n763 163.367
R1375 B.n764 B.n127 163.367
R1376 B.n768 B.n127 163.367
R1377 B.n769 B.n768 163.367
R1378 B.n770 B.n769 163.367
R1379 B.n770 B.n125 163.367
R1380 B.n774 B.n125 163.367
R1381 B.n775 B.n774 163.367
R1382 B.n776 B.n775 163.367
R1383 B.n776 B.n123 163.367
R1384 B.n780 B.n123 163.367
R1385 B.n781 B.n780 163.367
R1386 B.n782 B.n781 163.367
R1387 B.n782 B.n121 163.367
R1388 B.n786 B.n121 163.367
R1389 B.n787 B.n786 163.367
R1390 B.n788 B.n787 163.367
R1391 B.n788 B.n119 163.367
R1392 B.n792 B.n119 163.367
R1393 B.n793 B.n792 163.367
R1394 B.n794 B.n793 163.367
R1395 B.n794 B.n117 163.367
R1396 B.n798 B.n117 163.367
R1397 B.n799 B.n798 163.367
R1398 B.n800 B.n799 163.367
R1399 B.n800 B.n115 163.367
R1400 B.n804 B.n115 163.367
R1401 B.n805 B.n804 163.367
R1402 B.n806 B.n805 163.367
R1403 B.n806 B.n113 163.367
R1404 B.n810 B.n113 163.367
R1405 B.n811 B.n810 163.367
R1406 B.n812 B.n811 163.367
R1407 B.n812 B.n111 163.367
R1408 B.n816 B.n111 163.367
R1409 B.n817 B.n816 163.367
R1410 B.n818 B.n817 163.367
R1411 B.n818 B.n109 163.367
R1412 B.n1016 B.n39 163.367
R1413 B.n1016 B.n1015 163.367
R1414 B.n1015 B.n1014 163.367
R1415 B.n1014 B.n41 163.367
R1416 B.n1010 B.n41 163.367
R1417 B.n1010 B.n1009 163.367
R1418 B.n1009 B.n1008 163.367
R1419 B.n1008 B.n43 163.367
R1420 B.n1004 B.n43 163.367
R1421 B.n1004 B.n1003 163.367
R1422 B.n1003 B.n1002 163.367
R1423 B.n1002 B.n45 163.367
R1424 B.n998 B.n45 163.367
R1425 B.n998 B.n997 163.367
R1426 B.n997 B.n996 163.367
R1427 B.n996 B.n47 163.367
R1428 B.n992 B.n47 163.367
R1429 B.n992 B.n991 163.367
R1430 B.n991 B.n990 163.367
R1431 B.n990 B.n49 163.367
R1432 B.n986 B.n49 163.367
R1433 B.n986 B.n985 163.367
R1434 B.n985 B.n984 163.367
R1435 B.n984 B.n51 163.367
R1436 B.n980 B.n51 163.367
R1437 B.n980 B.n979 163.367
R1438 B.n979 B.n978 163.367
R1439 B.n978 B.n53 163.367
R1440 B.n974 B.n53 163.367
R1441 B.n974 B.n973 163.367
R1442 B.n973 B.n972 163.367
R1443 B.n972 B.n55 163.367
R1444 B.n968 B.n55 163.367
R1445 B.n968 B.n967 163.367
R1446 B.n967 B.n966 163.367
R1447 B.n966 B.n57 163.367
R1448 B.n962 B.n57 163.367
R1449 B.n962 B.n961 163.367
R1450 B.n961 B.n960 163.367
R1451 B.n960 B.n59 163.367
R1452 B.n956 B.n59 163.367
R1453 B.n956 B.n955 163.367
R1454 B.n955 B.n954 163.367
R1455 B.n954 B.n61 163.367
R1456 B.n950 B.n61 163.367
R1457 B.n950 B.n949 163.367
R1458 B.n949 B.n948 163.367
R1459 B.n948 B.n63 163.367
R1460 B.n944 B.n63 163.367
R1461 B.n944 B.n943 163.367
R1462 B.n943 B.n942 163.367
R1463 B.n942 B.n65 163.367
R1464 B.n938 B.n65 163.367
R1465 B.n938 B.n937 163.367
R1466 B.n937 B.n936 163.367
R1467 B.n936 B.n67 163.367
R1468 B.n932 B.n67 163.367
R1469 B.n932 B.n931 163.367
R1470 B.n931 B.n930 163.367
R1471 B.n930 B.n69 163.367
R1472 B.n925 B.n69 163.367
R1473 B.n925 B.n924 163.367
R1474 B.n924 B.n923 163.367
R1475 B.n923 B.n73 163.367
R1476 B.n919 B.n73 163.367
R1477 B.n919 B.n918 163.367
R1478 B.n918 B.n917 163.367
R1479 B.n917 B.n75 163.367
R1480 B.n913 B.n75 163.367
R1481 B.n913 B.n912 163.367
R1482 B.n912 B.n79 163.367
R1483 B.n908 B.n79 163.367
R1484 B.n908 B.n907 163.367
R1485 B.n907 B.n906 163.367
R1486 B.n906 B.n81 163.367
R1487 B.n902 B.n81 163.367
R1488 B.n902 B.n901 163.367
R1489 B.n901 B.n900 163.367
R1490 B.n900 B.n83 163.367
R1491 B.n896 B.n83 163.367
R1492 B.n896 B.n895 163.367
R1493 B.n895 B.n894 163.367
R1494 B.n894 B.n85 163.367
R1495 B.n890 B.n85 163.367
R1496 B.n890 B.n889 163.367
R1497 B.n889 B.n888 163.367
R1498 B.n888 B.n87 163.367
R1499 B.n884 B.n87 163.367
R1500 B.n884 B.n883 163.367
R1501 B.n883 B.n882 163.367
R1502 B.n882 B.n89 163.367
R1503 B.n878 B.n89 163.367
R1504 B.n878 B.n877 163.367
R1505 B.n877 B.n876 163.367
R1506 B.n876 B.n91 163.367
R1507 B.n872 B.n91 163.367
R1508 B.n872 B.n871 163.367
R1509 B.n871 B.n870 163.367
R1510 B.n870 B.n93 163.367
R1511 B.n866 B.n93 163.367
R1512 B.n866 B.n865 163.367
R1513 B.n865 B.n864 163.367
R1514 B.n864 B.n95 163.367
R1515 B.n860 B.n95 163.367
R1516 B.n860 B.n859 163.367
R1517 B.n859 B.n858 163.367
R1518 B.n858 B.n97 163.367
R1519 B.n854 B.n97 163.367
R1520 B.n854 B.n853 163.367
R1521 B.n853 B.n852 163.367
R1522 B.n852 B.n99 163.367
R1523 B.n848 B.n99 163.367
R1524 B.n848 B.n847 163.367
R1525 B.n847 B.n846 163.367
R1526 B.n846 B.n101 163.367
R1527 B.n842 B.n101 163.367
R1528 B.n842 B.n841 163.367
R1529 B.n841 B.n840 163.367
R1530 B.n840 B.n103 163.367
R1531 B.n836 B.n103 163.367
R1532 B.n836 B.n835 163.367
R1533 B.n835 B.n834 163.367
R1534 B.n834 B.n105 163.367
R1535 B.n830 B.n105 163.367
R1536 B.n830 B.n829 163.367
R1537 B.n829 B.n828 163.367
R1538 B.n828 B.n107 163.367
R1539 B.n824 B.n107 163.367
R1540 B.n824 B.n823 163.367
R1541 B.n823 B.n822 163.367
R1542 B.n215 B.t10 110.222
R1543 B.n77 B.t5 110.222
R1544 B.n223 B.t7 110.198
R1545 B.n71 B.t2 110.198
R1546 B.n215 B.n214 72.5338
R1547 B.n223 B.n222 72.5338
R1548 B.n71 B.n70 72.5338
R1549 B.n77 B.n76 72.5338
R1550 B.n216 B.n215 59.5399
R1551 B.n491 B.n223 59.5399
R1552 B.n927 B.n71 59.5399
R1553 B.n78 B.n77 59.5399
R1554 B.n1019 B.n1018 36.059
R1555 B.n598 B.n597 36.059
R1556 B.n400 B.n399 36.059
R1557 B.n821 B.n820 36.059
R1558 B B.n1131 18.0485
R1559 B.n1018 B.n1017 10.6151
R1560 B.n1017 B.n40 10.6151
R1561 B.n1013 B.n40 10.6151
R1562 B.n1013 B.n1012 10.6151
R1563 B.n1012 B.n1011 10.6151
R1564 B.n1011 B.n42 10.6151
R1565 B.n1007 B.n42 10.6151
R1566 B.n1007 B.n1006 10.6151
R1567 B.n1006 B.n1005 10.6151
R1568 B.n1005 B.n44 10.6151
R1569 B.n1001 B.n44 10.6151
R1570 B.n1001 B.n1000 10.6151
R1571 B.n1000 B.n999 10.6151
R1572 B.n999 B.n46 10.6151
R1573 B.n995 B.n46 10.6151
R1574 B.n995 B.n994 10.6151
R1575 B.n994 B.n993 10.6151
R1576 B.n993 B.n48 10.6151
R1577 B.n989 B.n48 10.6151
R1578 B.n989 B.n988 10.6151
R1579 B.n988 B.n987 10.6151
R1580 B.n987 B.n50 10.6151
R1581 B.n983 B.n50 10.6151
R1582 B.n983 B.n982 10.6151
R1583 B.n982 B.n981 10.6151
R1584 B.n981 B.n52 10.6151
R1585 B.n977 B.n52 10.6151
R1586 B.n977 B.n976 10.6151
R1587 B.n976 B.n975 10.6151
R1588 B.n975 B.n54 10.6151
R1589 B.n971 B.n54 10.6151
R1590 B.n971 B.n970 10.6151
R1591 B.n970 B.n969 10.6151
R1592 B.n969 B.n56 10.6151
R1593 B.n965 B.n56 10.6151
R1594 B.n965 B.n964 10.6151
R1595 B.n964 B.n963 10.6151
R1596 B.n963 B.n58 10.6151
R1597 B.n959 B.n58 10.6151
R1598 B.n959 B.n958 10.6151
R1599 B.n958 B.n957 10.6151
R1600 B.n957 B.n60 10.6151
R1601 B.n953 B.n60 10.6151
R1602 B.n953 B.n952 10.6151
R1603 B.n952 B.n951 10.6151
R1604 B.n951 B.n62 10.6151
R1605 B.n947 B.n62 10.6151
R1606 B.n947 B.n946 10.6151
R1607 B.n946 B.n945 10.6151
R1608 B.n945 B.n64 10.6151
R1609 B.n941 B.n64 10.6151
R1610 B.n941 B.n940 10.6151
R1611 B.n940 B.n939 10.6151
R1612 B.n939 B.n66 10.6151
R1613 B.n935 B.n66 10.6151
R1614 B.n935 B.n934 10.6151
R1615 B.n934 B.n933 10.6151
R1616 B.n933 B.n68 10.6151
R1617 B.n929 B.n68 10.6151
R1618 B.n929 B.n928 10.6151
R1619 B.n926 B.n72 10.6151
R1620 B.n922 B.n72 10.6151
R1621 B.n922 B.n921 10.6151
R1622 B.n921 B.n920 10.6151
R1623 B.n920 B.n74 10.6151
R1624 B.n916 B.n74 10.6151
R1625 B.n916 B.n915 10.6151
R1626 B.n915 B.n914 10.6151
R1627 B.n911 B.n910 10.6151
R1628 B.n910 B.n909 10.6151
R1629 B.n909 B.n80 10.6151
R1630 B.n905 B.n80 10.6151
R1631 B.n905 B.n904 10.6151
R1632 B.n904 B.n903 10.6151
R1633 B.n903 B.n82 10.6151
R1634 B.n899 B.n82 10.6151
R1635 B.n899 B.n898 10.6151
R1636 B.n898 B.n897 10.6151
R1637 B.n897 B.n84 10.6151
R1638 B.n893 B.n84 10.6151
R1639 B.n893 B.n892 10.6151
R1640 B.n892 B.n891 10.6151
R1641 B.n891 B.n86 10.6151
R1642 B.n887 B.n86 10.6151
R1643 B.n887 B.n886 10.6151
R1644 B.n886 B.n885 10.6151
R1645 B.n885 B.n88 10.6151
R1646 B.n881 B.n88 10.6151
R1647 B.n881 B.n880 10.6151
R1648 B.n880 B.n879 10.6151
R1649 B.n879 B.n90 10.6151
R1650 B.n875 B.n90 10.6151
R1651 B.n875 B.n874 10.6151
R1652 B.n874 B.n873 10.6151
R1653 B.n873 B.n92 10.6151
R1654 B.n869 B.n92 10.6151
R1655 B.n869 B.n868 10.6151
R1656 B.n868 B.n867 10.6151
R1657 B.n867 B.n94 10.6151
R1658 B.n863 B.n94 10.6151
R1659 B.n863 B.n862 10.6151
R1660 B.n862 B.n861 10.6151
R1661 B.n861 B.n96 10.6151
R1662 B.n857 B.n96 10.6151
R1663 B.n857 B.n856 10.6151
R1664 B.n856 B.n855 10.6151
R1665 B.n855 B.n98 10.6151
R1666 B.n851 B.n98 10.6151
R1667 B.n851 B.n850 10.6151
R1668 B.n850 B.n849 10.6151
R1669 B.n849 B.n100 10.6151
R1670 B.n845 B.n100 10.6151
R1671 B.n845 B.n844 10.6151
R1672 B.n844 B.n843 10.6151
R1673 B.n843 B.n102 10.6151
R1674 B.n839 B.n102 10.6151
R1675 B.n839 B.n838 10.6151
R1676 B.n838 B.n837 10.6151
R1677 B.n837 B.n104 10.6151
R1678 B.n833 B.n104 10.6151
R1679 B.n833 B.n832 10.6151
R1680 B.n832 B.n831 10.6151
R1681 B.n831 B.n106 10.6151
R1682 B.n827 B.n106 10.6151
R1683 B.n827 B.n826 10.6151
R1684 B.n826 B.n825 10.6151
R1685 B.n825 B.n108 10.6151
R1686 B.n821 B.n108 10.6151
R1687 B.n599 B.n598 10.6151
R1688 B.n599 B.n182 10.6151
R1689 B.n603 B.n182 10.6151
R1690 B.n604 B.n603 10.6151
R1691 B.n605 B.n604 10.6151
R1692 B.n605 B.n180 10.6151
R1693 B.n609 B.n180 10.6151
R1694 B.n610 B.n609 10.6151
R1695 B.n611 B.n610 10.6151
R1696 B.n611 B.n178 10.6151
R1697 B.n615 B.n178 10.6151
R1698 B.n616 B.n615 10.6151
R1699 B.n617 B.n616 10.6151
R1700 B.n617 B.n176 10.6151
R1701 B.n621 B.n176 10.6151
R1702 B.n622 B.n621 10.6151
R1703 B.n623 B.n622 10.6151
R1704 B.n623 B.n174 10.6151
R1705 B.n627 B.n174 10.6151
R1706 B.n628 B.n627 10.6151
R1707 B.n629 B.n628 10.6151
R1708 B.n629 B.n172 10.6151
R1709 B.n633 B.n172 10.6151
R1710 B.n634 B.n633 10.6151
R1711 B.n635 B.n634 10.6151
R1712 B.n635 B.n170 10.6151
R1713 B.n639 B.n170 10.6151
R1714 B.n640 B.n639 10.6151
R1715 B.n641 B.n640 10.6151
R1716 B.n641 B.n168 10.6151
R1717 B.n645 B.n168 10.6151
R1718 B.n646 B.n645 10.6151
R1719 B.n647 B.n646 10.6151
R1720 B.n647 B.n166 10.6151
R1721 B.n651 B.n166 10.6151
R1722 B.n652 B.n651 10.6151
R1723 B.n653 B.n652 10.6151
R1724 B.n653 B.n164 10.6151
R1725 B.n657 B.n164 10.6151
R1726 B.n658 B.n657 10.6151
R1727 B.n659 B.n658 10.6151
R1728 B.n659 B.n162 10.6151
R1729 B.n663 B.n162 10.6151
R1730 B.n664 B.n663 10.6151
R1731 B.n665 B.n664 10.6151
R1732 B.n665 B.n160 10.6151
R1733 B.n669 B.n160 10.6151
R1734 B.n670 B.n669 10.6151
R1735 B.n671 B.n670 10.6151
R1736 B.n671 B.n158 10.6151
R1737 B.n675 B.n158 10.6151
R1738 B.n676 B.n675 10.6151
R1739 B.n677 B.n676 10.6151
R1740 B.n677 B.n156 10.6151
R1741 B.n681 B.n156 10.6151
R1742 B.n682 B.n681 10.6151
R1743 B.n683 B.n682 10.6151
R1744 B.n683 B.n154 10.6151
R1745 B.n687 B.n154 10.6151
R1746 B.n688 B.n687 10.6151
R1747 B.n689 B.n688 10.6151
R1748 B.n689 B.n152 10.6151
R1749 B.n693 B.n152 10.6151
R1750 B.n694 B.n693 10.6151
R1751 B.n695 B.n694 10.6151
R1752 B.n695 B.n150 10.6151
R1753 B.n699 B.n150 10.6151
R1754 B.n700 B.n699 10.6151
R1755 B.n701 B.n700 10.6151
R1756 B.n701 B.n148 10.6151
R1757 B.n705 B.n148 10.6151
R1758 B.n706 B.n705 10.6151
R1759 B.n707 B.n706 10.6151
R1760 B.n707 B.n146 10.6151
R1761 B.n711 B.n146 10.6151
R1762 B.n712 B.n711 10.6151
R1763 B.n713 B.n712 10.6151
R1764 B.n713 B.n144 10.6151
R1765 B.n717 B.n144 10.6151
R1766 B.n718 B.n717 10.6151
R1767 B.n719 B.n718 10.6151
R1768 B.n719 B.n142 10.6151
R1769 B.n723 B.n142 10.6151
R1770 B.n724 B.n723 10.6151
R1771 B.n725 B.n724 10.6151
R1772 B.n725 B.n140 10.6151
R1773 B.n729 B.n140 10.6151
R1774 B.n730 B.n729 10.6151
R1775 B.n731 B.n730 10.6151
R1776 B.n731 B.n138 10.6151
R1777 B.n735 B.n138 10.6151
R1778 B.n736 B.n735 10.6151
R1779 B.n737 B.n736 10.6151
R1780 B.n737 B.n136 10.6151
R1781 B.n741 B.n136 10.6151
R1782 B.n742 B.n741 10.6151
R1783 B.n743 B.n742 10.6151
R1784 B.n743 B.n134 10.6151
R1785 B.n747 B.n134 10.6151
R1786 B.n748 B.n747 10.6151
R1787 B.n749 B.n748 10.6151
R1788 B.n749 B.n132 10.6151
R1789 B.n753 B.n132 10.6151
R1790 B.n754 B.n753 10.6151
R1791 B.n755 B.n754 10.6151
R1792 B.n755 B.n130 10.6151
R1793 B.n759 B.n130 10.6151
R1794 B.n760 B.n759 10.6151
R1795 B.n761 B.n760 10.6151
R1796 B.n761 B.n128 10.6151
R1797 B.n765 B.n128 10.6151
R1798 B.n766 B.n765 10.6151
R1799 B.n767 B.n766 10.6151
R1800 B.n767 B.n126 10.6151
R1801 B.n771 B.n126 10.6151
R1802 B.n772 B.n771 10.6151
R1803 B.n773 B.n772 10.6151
R1804 B.n773 B.n124 10.6151
R1805 B.n777 B.n124 10.6151
R1806 B.n778 B.n777 10.6151
R1807 B.n779 B.n778 10.6151
R1808 B.n779 B.n122 10.6151
R1809 B.n783 B.n122 10.6151
R1810 B.n784 B.n783 10.6151
R1811 B.n785 B.n784 10.6151
R1812 B.n785 B.n120 10.6151
R1813 B.n789 B.n120 10.6151
R1814 B.n790 B.n789 10.6151
R1815 B.n791 B.n790 10.6151
R1816 B.n791 B.n118 10.6151
R1817 B.n795 B.n118 10.6151
R1818 B.n796 B.n795 10.6151
R1819 B.n797 B.n796 10.6151
R1820 B.n797 B.n116 10.6151
R1821 B.n801 B.n116 10.6151
R1822 B.n802 B.n801 10.6151
R1823 B.n803 B.n802 10.6151
R1824 B.n803 B.n114 10.6151
R1825 B.n807 B.n114 10.6151
R1826 B.n808 B.n807 10.6151
R1827 B.n809 B.n808 10.6151
R1828 B.n809 B.n112 10.6151
R1829 B.n813 B.n112 10.6151
R1830 B.n814 B.n813 10.6151
R1831 B.n815 B.n814 10.6151
R1832 B.n815 B.n110 10.6151
R1833 B.n819 B.n110 10.6151
R1834 B.n820 B.n819 10.6151
R1835 B.n401 B.n400 10.6151
R1836 B.n401 B.n252 10.6151
R1837 B.n405 B.n252 10.6151
R1838 B.n406 B.n405 10.6151
R1839 B.n407 B.n406 10.6151
R1840 B.n407 B.n250 10.6151
R1841 B.n411 B.n250 10.6151
R1842 B.n412 B.n411 10.6151
R1843 B.n413 B.n412 10.6151
R1844 B.n413 B.n248 10.6151
R1845 B.n417 B.n248 10.6151
R1846 B.n418 B.n417 10.6151
R1847 B.n419 B.n418 10.6151
R1848 B.n419 B.n246 10.6151
R1849 B.n423 B.n246 10.6151
R1850 B.n424 B.n423 10.6151
R1851 B.n425 B.n424 10.6151
R1852 B.n425 B.n244 10.6151
R1853 B.n429 B.n244 10.6151
R1854 B.n430 B.n429 10.6151
R1855 B.n431 B.n430 10.6151
R1856 B.n431 B.n242 10.6151
R1857 B.n435 B.n242 10.6151
R1858 B.n436 B.n435 10.6151
R1859 B.n437 B.n436 10.6151
R1860 B.n437 B.n240 10.6151
R1861 B.n441 B.n240 10.6151
R1862 B.n442 B.n441 10.6151
R1863 B.n443 B.n442 10.6151
R1864 B.n443 B.n238 10.6151
R1865 B.n447 B.n238 10.6151
R1866 B.n448 B.n447 10.6151
R1867 B.n449 B.n448 10.6151
R1868 B.n449 B.n236 10.6151
R1869 B.n453 B.n236 10.6151
R1870 B.n454 B.n453 10.6151
R1871 B.n455 B.n454 10.6151
R1872 B.n455 B.n234 10.6151
R1873 B.n459 B.n234 10.6151
R1874 B.n460 B.n459 10.6151
R1875 B.n461 B.n460 10.6151
R1876 B.n461 B.n232 10.6151
R1877 B.n465 B.n232 10.6151
R1878 B.n466 B.n465 10.6151
R1879 B.n467 B.n466 10.6151
R1880 B.n467 B.n230 10.6151
R1881 B.n471 B.n230 10.6151
R1882 B.n472 B.n471 10.6151
R1883 B.n473 B.n472 10.6151
R1884 B.n473 B.n228 10.6151
R1885 B.n477 B.n228 10.6151
R1886 B.n478 B.n477 10.6151
R1887 B.n479 B.n478 10.6151
R1888 B.n479 B.n226 10.6151
R1889 B.n483 B.n226 10.6151
R1890 B.n484 B.n483 10.6151
R1891 B.n485 B.n484 10.6151
R1892 B.n485 B.n224 10.6151
R1893 B.n489 B.n224 10.6151
R1894 B.n490 B.n489 10.6151
R1895 B.n492 B.n220 10.6151
R1896 B.n496 B.n220 10.6151
R1897 B.n497 B.n496 10.6151
R1898 B.n498 B.n497 10.6151
R1899 B.n498 B.n218 10.6151
R1900 B.n502 B.n218 10.6151
R1901 B.n503 B.n502 10.6151
R1902 B.n504 B.n503 10.6151
R1903 B.n508 B.n507 10.6151
R1904 B.n509 B.n508 10.6151
R1905 B.n509 B.n212 10.6151
R1906 B.n513 B.n212 10.6151
R1907 B.n514 B.n513 10.6151
R1908 B.n515 B.n514 10.6151
R1909 B.n515 B.n210 10.6151
R1910 B.n519 B.n210 10.6151
R1911 B.n520 B.n519 10.6151
R1912 B.n521 B.n520 10.6151
R1913 B.n521 B.n208 10.6151
R1914 B.n525 B.n208 10.6151
R1915 B.n526 B.n525 10.6151
R1916 B.n527 B.n526 10.6151
R1917 B.n527 B.n206 10.6151
R1918 B.n531 B.n206 10.6151
R1919 B.n532 B.n531 10.6151
R1920 B.n533 B.n532 10.6151
R1921 B.n533 B.n204 10.6151
R1922 B.n537 B.n204 10.6151
R1923 B.n538 B.n537 10.6151
R1924 B.n539 B.n538 10.6151
R1925 B.n539 B.n202 10.6151
R1926 B.n543 B.n202 10.6151
R1927 B.n544 B.n543 10.6151
R1928 B.n545 B.n544 10.6151
R1929 B.n545 B.n200 10.6151
R1930 B.n549 B.n200 10.6151
R1931 B.n550 B.n549 10.6151
R1932 B.n551 B.n550 10.6151
R1933 B.n551 B.n198 10.6151
R1934 B.n555 B.n198 10.6151
R1935 B.n556 B.n555 10.6151
R1936 B.n557 B.n556 10.6151
R1937 B.n557 B.n196 10.6151
R1938 B.n561 B.n196 10.6151
R1939 B.n562 B.n561 10.6151
R1940 B.n563 B.n562 10.6151
R1941 B.n563 B.n194 10.6151
R1942 B.n567 B.n194 10.6151
R1943 B.n568 B.n567 10.6151
R1944 B.n569 B.n568 10.6151
R1945 B.n569 B.n192 10.6151
R1946 B.n573 B.n192 10.6151
R1947 B.n574 B.n573 10.6151
R1948 B.n575 B.n574 10.6151
R1949 B.n575 B.n190 10.6151
R1950 B.n579 B.n190 10.6151
R1951 B.n580 B.n579 10.6151
R1952 B.n581 B.n580 10.6151
R1953 B.n581 B.n188 10.6151
R1954 B.n585 B.n188 10.6151
R1955 B.n586 B.n585 10.6151
R1956 B.n587 B.n586 10.6151
R1957 B.n587 B.n186 10.6151
R1958 B.n591 B.n186 10.6151
R1959 B.n592 B.n591 10.6151
R1960 B.n593 B.n592 10.6151
R1961 B.n593 B.n184 10.6151
R1962 B.n597 B.n184 10.6151
R1963 B.n399 B.n254 10.6151
R1964 B.n395 B.n254 10.6151
R1965 B.n395 B.n394 10.6151
R1966 B.n394 B.n393 10.6151
R1967 B.n393 B.n256 10.6151
R1968 B.n389 B.n256 10.6151
R1969 B.n389 B.n388 10.6151
R1970 B.n388 B.n387 10.6151
R1971 B.n387 B.n258 10.6151
R1972 B.n383 B.n258 10.6151
R1973 B.n383 B.n382 10.6151
R1974 B.n382 B.n381 10.6151
R1975 B.n381 B.n260 10.6151
R1976 B.n377 B.n260 10.6151
R1977 B.n377 B.n376 10.6151
R1978 B.n376 B.n375 10.6151
R1979 B.n375 B.n262 10.6151
R1980 B.n371 B.n262 10.6151
R1981 B.n371 B.n370 10.6151
R1982 B.n370 B.n369 10.6151
R1983 B.n369 B.n264 10.6151
R1984 B.n365 B.n264 10.6151
R1985 B.n365 B.n364 10.6151
R1986 B.n364 B.n363 10.6151
R1987 B.n363 B.n266 10.6151
R1988 B.n359 B.n266 10.6151
R1989 B.n359 B.n358 10.6151
R1990 B.n358 B.n357 10.6151
R1991 B.n357 B.n268 10.6151
R1992 B.n353 B.n268 10.6151
R1993 B.n353 B.n352 10.6151
R1994 B.n352 B.n351 10.6151
R1995 B.n351 B.n270 10.6151
R1996 B.n347 B.n270 10.6151
R1997 B.n347 B.n346 10.6151
R1998 B.n346 B.n345 10.6151
R1999 B.n345 B.n272 10.6151
R2000 B.n341 B.n272 10.6151
R2001 B.n341 B.n340 10.6151
R2002 B.n340 B.n339 10.6151
R2003 B.n339 B.n274 10.6151
R2004 B.n335 B.n274 10.6151
R2005 B.n335 B.n334 10.6151
R2006 B.n334 B.n333 10.6151
R2007 B.n333 B.n276 10.6151
R2008 B.n329 B.n276 10.6151
R2009 B.n329 B.n328 10.6151
R2010 B.n328 B.n327 10.6151
R2011 B.n327 B.n278 10.6151
R2012 B.n323 B.n278 10.6151
R2013 B.n323 B.n322 10.6151
R2014 B.n322 B.n321 10.6151
R2015 B.n321 B.n280 10.6151
R2016 B.n317 B.n280 10.6151
R2017 B.n317 B.n316 10.6151
R2018 B.n316 B.n315 10.6151
R2019 B.n315 B.n282 10.6151
R2020 B.n311 B.n282 10.6151
R2021 B.n311 B.n310 10.6151
R2022 B.n310 B.n309 10.6151
R2023 B.n309 B.n284 10.6151
R2024 B.n305 B.n284 10.6151
R2025 B.n305 B.n304 10.6151
R2026 B.n304 B.n303 10.6151
R2027 B.n303 B.n286 10.6151
R2028 B.n299 B.n286 10.6151
R2029 B.n299 B.n298 10.6151
R2030 B.n298 B.n297 10.6151
R2031 B.n297 B.n288 10.6151
R2032 B.n293 B.n288 10.6151
R2033 B.n293 B.n292 10.6151
R2034 B.n292 B.n291 10.6151
R2035 B.n291 B.n0 10.6151
R2036 B.n1127 B.n1 10.6151
R2037 B.n1127 B.n1126 10.6151
R2038 B.n1126 B.n1125 10.6151
R2039 B.n1125 B.n4 10.6151
R2040 B.n1121 B.n4 10.6151
R2041 B.n1121 B.n1120 10.6151
R2042 B.n1120 B.n1119 10.6151
R2043 B.n1119 B.n6 10.6151
R2044 B.n1115 B.n6 10.6151
R2045 B.n1115 B.n1114 10.6151
R2046 B.n1114 B.n1113 10.6151
R2047 B.n1113 B.n8 10.6151
R2048 B.n1109 B.n8 10.6151
R2049 B.n1109 B.n1108 10.6151
R2050 B.n1108 B.n1107 10.6151
R2051 B.n1107 B.n10 10.6151
R2052 B.n1103 B.n10 10.6151
R2053 B.n1103 B.n1102 10.6151
R2054 B.n1102 B.n1101 10.6151
R2055 B.n1101 B.n12 10.6151
R2056 B.n1097 B.n12 10.6151
R2057 B.n1097 B.n1096 10.6151
R2058 B.n1096 B.n1095 10.6151
R2059 B.n1095 B.n14 10.6151
R2060 B.n1091 B.n14 10.6151
R2061 B.n1091 B.n1090 10.6151
R2062 B.n1090 B.n1089 10.6151
R2063 B.n1089 B.n16 10.6151
R2064 B.n1085 B.n16 10.6151
R2065 B.n1085 B.n1084 10.6151
R2066 B.n1084 B.n1083 10.6151
R2067 B.n1083 B.n18 10.6151
R2068 B.n1079 B.n18 10.6151
R2069 B.n1079 B.n1078 10.6151
R2070 B.n1078 B.n1077 10.6151
R2071 B.n1077 B.n20 10.6151
R2072 B.n1073 B.n20 10.6151
R2073 B.n1073 B.n1072 10.6151
R2074 B.n1072 B.n1071 10.6151
R2075 B.n1071 B.n22 10.6151
R2076 B.n1067 B.n22 10.6151
R2077 B.n1067 B.n1066 10.6151
R2078 B.n1066 B.n1065 10.6151
R2079 B.n1065 B.n24 10.6151
R2080 B.n1061 B.n24 10.6151
R2081 B.n1061 B.n1060 10.6151
R2082 B.n1060 B.n1059 10.6151
R2083 B.n1059 B.n26 10.6151
R2084 B.n1055 B.n26 10.6151
R2085 B.n1055 B.n1054 10.6151
R2086 B.n1054 B.n1053 10.6151
R2087 B.n1053 B.n28 10.6151
R2088 B.n1049 B.n28 10.6151
R2089 B.n1049 B.n1048 10.6151
R2090 B.n1048 B.n1047 10.6151
R2091 B.n1047 B.n30 10.6151
R2092 B.n1043 B.n30 10.6151
R2093 B.n1043 B.n1042 10.6151
R2094 B.n1042 B.n1041 10.6151
R2095 B.n1041 B.n32 10.6151
R2096 B.n1037 B.n32 10.6151
R2097 B.n1037 B.n1036 10.6151
R2098 B.n1036 B.n1035 10.6151
R2099 B.n1035 B.n34 10.6151
R2100 B.n1031 B.n34 10.6151
R2101 B.n1031 B.n1030 10.6151
R2102 B.n1030 B.n1029 10.6151
R2103 B.n1029 B.n36 10.6151
R2104 B.n1025 B.n36 10.6151
R2105 B.n1025 B.n1024 10.6151
R2106 B.n1024 B.n1023 10.6151
R2107 B.n1023 B.n38 10.6151
R2108 B.n1019 B.n38 10.6151
R2109 B.n927 B.n926 6.5566
R2110 B.n914 B.n78 6.5566
R2111 B.n492 B.n491 6.5566
R2112 B.n504 B.n216 6.5566
R2113 B.n928 B.n927 4.05904
R2114 B.n911 B.n78 4.05904
R2115 B.n491 B.n490 4.05904
R2116 B.n507 B.n216 4.05904
R2117 B.n1131 B.n0 2.81026
R2118 B.n1131 B.n1 2.81026
C0 VP B 2.77017f
C1 VP w_n5458_n4682# 12.757299f
C2 VP VTAIL 17.7205f
C3 VN VP 10.8109f
C4 w_n5458_n4682# B 13.7505f
C5 VDD1 VP 17.5519f
C6 VP VDD2 0.68738f
C7 VTAIL B 5.58692f
C8 VN B 1.56658f
C9 w_n5458_n4682# VTAIL 4.22228f
C10 VN w_n5458_n4682# 12.0442f
C11 VN VTAIL 17.7062f
C12 VDD1 B 3.32338f
C13 VDD2 B 3.47284f
C14 VDD1 w_n5458_n4682# 3.54735f
C15 w_n5458_n4682# VDD2 3.733f
C16 VDD1 VTAIL 13.411901f
C17 VDD2 VTAIL 13.4678f
C18 VDD1 VN 0.155244f
C19 VN VDD2 17.0246f
C20 VDD1 VDD2 2.70283f
C21 VDD2 VSUBS 2.59294f
C22 VDD1 VSUBS 2.459325f
C23 VTAIL VSUBS 1.717581f
C24 VN VSUBS 9.24902f
C25 VP VSUBS 5.511901f
C26 B VSUBS 6.925285f
C27 w_n5458_n4682# VSUBS 0.31235p
C28 B.n0 VSUBS 0.004839f
C29 B.n1 VSUBS 0.004839f
C30 B.n2 VSUBS 0.007653f
C31 B.n3 VSUBS 0.007653f
C32 B.n4 VSUBS 0.007653f
C33 B.n5 VSUBS 0.007653f
C34 B.n6 VSUBS 0.007653f
C35 B.n7 VSUBS 0.007653f
C36 B.n8 VSUBS 0.007653f
C37 B.n9 VSUBS 0.007653f
C38 B.n10 VSUBS 0.007653f
C39 B.n11 VSUBS 0.007653f
C40 B.n12 VSUBS 0.007653f
C41 B.n13 VSUBS 0.007653f
C42 B.n14 VSUBS 0.007653f
C43 B.n15 VSUBS 0.007653f
C44 B.n16 VSUBS 0.007653f
C45 B.n17 VSUBS 0.007653f
C46 B.n18 VSUBS 0.007653f
C47 B.n19 VSUBS 0.007653f
C48 B.n20 VSUBS 0.007653f
C49 B.n21 VSUBS 0.007653f
C50 B.n22 VSUBS 0.007653f
C51 B.n23 VSUBS 0.007653f
C52 B.n24 VSUBS 0.007653f
C53 B.n25 VSUBS 0.007653f
C54 B.n26 VSUBS 0.007653f
C55 B.n27 VSUBS 0.007653f
C56 B.n28 VSUBS 0.007653f
C57 B.n29 VSUBS 0.007653f
C58 B.n30 VSUBS 0.007653f
C59 B.n31 VSUBS 0.007653f
C60 B.n32 VSUBS 0.007653f
C61 B.n33 VSUBS 0.007653f
C62 B.n34 VSUBS 0.007653f
C63 B.n35 VSUBS 0.007653f
C64 B.n36 VSUBS 0.007653f
C65 B.n37 VSUBS 0.007653f
C66 B.n38 VSUBS 0.007653f
C67 B.n39 VSUBS 0.019441f
C68 B.n40 VSUBS 0.007653f
C69 B.n41 VSUBS 0.007653f
C70 B.n42 VSUBS 0.007653f
C71 B.n43 VSUBS 0.007653f
C72 B.n44 VSUBS 0.007653f
C73 B.n45 VSUBS 0.007653f
C74 B.n46 VSUBS 0.007653f
C75 B.n47 VSUBS 0.007653f
C76 B.n48 VSUBS 0.007653f
C77 B.n49 VSUBS 0.007653f
C78 B.n50 VSUBS 0.007653f
C79 B.n51 VSUBS 0.007653f
C80 B.n52 VSUBS 0.007653f
C81 B.n53 VSUBS 0.007653f
C82 B.n54 VSUBS 0.007653f
C83 B.n55 VSUBS 0.007653f
C84 B.n56 VSUBS 0.007653f
C85 B.n57 VSUBS 0.007653f
C86 B.n58 VSUBS 0.007653f
C87 B.n59 VSUBS 0.007653f
C88 B.n60 VSUBS 0.007653f
C89 B.n61 VSUBS 0.007653f
C90 B.n62 VSUBS 0.007653f
C91 B.n63 VSUBS 0.007653f
C92 B.n64 VSUBS 0.007653f
C93 B.n65 VSUBS 0.007653f
C94 B.n66 VSUBS 0.007653f
C95 B.n67 VSUBS 0.007653f
C96 B.n68 VSUBS 0.007653f
C97 B.n69 VSUBS 0.007653f
C98 B.t2 VSUBS 0.68686f
C99 B.t1 VSUBS 0.71528f
C100 B.t0 VSUBS 3.12515f
C101 B.n70 VSUBS 0.434191f
C102 B.n71 VSUBS 0.082512f
C103 B.n72 VSUBS 0.007653f
C104 B.n73 VSUBS 0.007653f
C105 B.n74 VSUBS 0.007653f
C106 B.n75 VSUBS 0.007653f
C107 B.t5 VSUBS 0.686833f
C108 B.t4 VSUBS 0.71526f
C109 B.t3 VSUBS 3.12515f
C110 B.n76 VSUBS 0.43421f
C111 B.n77 VSUBS 0.082539f
C112 B.n78 VSUBS 0.01773f
C113 B.n79 VSUBS 0.007653f
C114 B.n80 VSUBS 0.007653f
C115 B.n81 VSUBS 0.007653f
C116 B.n82 VSUBS 0.007653f
C117 B.n83 VSUBS 0.007653f
C118 B.n84 VSUBS 0.007653f
C119 B.n85 VSUBS 0.007653f
C120 B.n86 VSUBS 0.007653f
C121 B.n87 VSUBS 0.007653f
C122 B.n88 VSUBS 0.007653f
C123 B.n89 VSUBS 0.007653f
C124 B.n90 VSUBS 0.007653f
C125 B.n91 VSUBS 0.007653f
C126 B.n92 VSUBS 0.007653f
C127 B.n93 VSUBS 0.007653f
C128 B.n94 VSUBS 0.007653f
C129 B.n95 VSUBS 0.007653f
C130 B.n96 VSUBS 0.007653f
C131 B.n97 VSUBS 0.007653f
C132 B.n98 VSUBS 0.007653f
C133 B.n99 VSUBS 0.007653f
C134 B.n100 VSUBS 0.007653f
C135 B.n101 VSUBS 0.007653f
C136 B.n102 VSUBS 0.007653f
C137 B.n103 VSUBS 0.007653f
C138 B.n104 VSUBS 0.007653f
C139 B.n105 VSUBS 0.007653f
C140 B.n106 VSUBS 0.007653f
C141 B.n107 VSUBS 0.007653f
C142 B.n108 VSUBS 0.007653f
C143 B.n109 VSUBS 0.018822f
C144 B.n110 VSUBS 0.007653f
C145 B.n111 VSUBS 0.007653f
C146 B.n112 VSUBS 0.007653f
C147 B.n113 VSUBS 0.007653f
C148 B.n114 VSUBS 0.007653f
C149 B.n115 VSUBS 0.007653f
C150 B.n116 VSUBS 0.007653f
C151 B.n117 VSUBS 0.007653f
C152 B.n118 VSUBS 0.007653f
C153 B.n119 VSUBS 0.007653f
C154 B.n120 VSUBS 0.007653f
C155 B.n121 VSUBS 0.007653f
C156 B.n122 VSUBS 0.007653f
C157 B.n123 VSUBS 0.007653f
C158 B.n124 VSUBS 0.007653f
C159 B.n125 VSUBS 0.007653f
C160 B.n126 VSUBS 0.007653f
C161 B.n127 VSUBS 0.007653f
C162 B.n128 VSUBS 0.007653f
C163 B.n129 VSUBS 0.007653f
C164 B.n130 VSUBS 0.007653f
C165 B.n131 VSUBS 0.007653f
C166 B.n132 VSUBS 0.007653f
C167 B.n133 VSUBS 0.007653f
C168 B.n134 VSUBS 0.007653f
C169 B.n135 VSUBS 0.007653f
C170 B.n136 VSUBS 0.007653f
C171 B.n137 VSUBS 0.007653f
C172 B.n138 VSUBS 0.007653f
C173 B.n139 VSUBS 0.007653f
C174 B.n140 VSUBS 0.007653f
C175 B.n141 VSUBS 0.007653f
C176 B.n142 VSUBS 0.007653f
C177 B.n143 VSUBS 0.007653f
C178 B.n144 VSUBS 0.007653f
C179 B.n145 VSUBS 0.007653f
C180 B.n146 VSUBS 0.007653f
C181 B.n147 VSUBS 0.007653f
C182 B.n148 VSUBS 0.007653f
C183 B.n149 VSUBS 0.007653f
C184 B.n150 VSUBS 0.007653f
C185 B.n151 VSUBS 0.007653f
C186 B.n152 VSUBS 0.007653f
C187 B.n153 VSUBS 0.007653f
C188 B.n154 VSUBS 0.007653f
C189 B.n155 VSUBS 0.007653f
C190 B.n156 VSUBS 0.007653f
C191 B.n157 VSUBS 0.007653f
C192 B.n158 VSUBS 0.007653f
C193 B.n159 VSUBS 0.007653f
C194 B.n160 VSUBS 0.007653f
C195 B.n161 VSUBS 0.007653f
C196 B.n162 VSUBS 0.007653f
C197 B.n163 VSUBS 0.007653f
C198 B.n164 VSUBS 0.007653f
C199 B.n165 VSUBS 0.007653f
C200 B.n166 VSUBS 0.007653f
C201 B.n167 VSUBS 0.007653f
C202 B.n168 VSUBS 0.007653f
C203 B.n169 VSUBS 0.007653f
C204 B.n170 VSUBS 0.007653f
C205 B.n171 VSUBS 0.007653f
C206 B.n172 VSUBS 0.007653f
C207 B.n173 VSUBS 0.007653f
C208 B.n174 VSUBS 0.007653f
C209 B.n175 VSUBS 0.007653f
C210 B.n176 VSUBS 0.007653f
C211 B.n177 VSUBS 0.007653f
C212 B.n178 VSUBS 0.007653f
C213 B.n179 VSUBS 0.007653f
C214 B.n180 VSUBS 0.007653f
C215 B.n181 VSUBS 0.007653f
C216 B.n182 VSUBS 0.007653f
C217 B.n183 VSUBS 0.018822f
C218 B.n184 VSUBS 0.007653f
C219 B.n185 VSUBS 0.007653f
C220 B.n186 VSUBS 0.007653f
C221 B.n187 VSUBS 0.007653f
C222 B.n188 VSUBS 0.007653f
C223 B.n189 VSUBS 0.007653f
C224 B.n190 VSUBS 0.007653f
C225 B.n191 VSUBS 0.007653f
C226 B.n192 VSUBS 0.007653f
C227 B.n193 VSUBS 0.007653f
C228 B.n194 VSUBS 0.007653f
C229 B.n195 VSUBS 0.007653f
C230 B.n196 VSUBS 0.007653f
C231 B.n197 VSUBS 0.007653f
C232 B.n198 VSUBS 0.007653f
C233 B.n199 VSUBS 0.007653f
C234 B.n200 VSUBS 0.007653f
C235 B.n201 VSUBS 0.007653f
C236 B.n202 VSUBS 0.007653f
C237 B.n203 VSUBS 0.007653f
C238 B.n204 VSUBS 0.007653f
C239 B.n205 VSUBS 0.007653f
C240 B.n206 VSUBS 0.007653f
C241 B.n207 VSUBS 0.007653f
C242 B.n208 VSUBS 0.007653f
C243 B.n209 VSUBS 0.007653f
C244 B.n210 VSUBS 0.007653f
C245 B.n211 VSUBS 0.007653f
C246 B.n212 VSUBS 0.007653f
C247 B.n213 VSUBS 0.007653f
C248 B.t10 VSUBS 0.686833f
C249 B.t11 VSUBS 0.71526f
C250 B.t9 VSUBS 3.12515f
C251 B.n214 VSUBS 0.43421f
C252 B.n215 VSUBS 0.082539f
C253 B.n216 VSUBS 0.01773f
C254 B.n217 VSUBS 0.007653f
C255 B.n218 VSUBS 0.007653f
C256 B.n219 VSUBS 0.007653f
C257 B.n220 VSUBS 0.007653f
C258 B.n221 VSUBS 0.007653f
C259 B.t7 VSUBS 0.68686f
C260 B.t8 VSUBS 0.71528f
C261 B.t6 VSUBS 3.12515f
C262 B.n222 VSUBS 0.434191f
C263 B.n223 VSUBS 0.082512f
C264 B.n224 VSUBS 0.007653f
C265 B.n225 VSUBS 0.007653f
C266 B.n226 VSUBS 0.007653f
C267 B.n227 VSUBS 0.007653f
C268 B.n228 VSUBS 0.007653f
C269 B.n229 VSUBS 0.007653f
C270 B.n230 VSUBS 0.007653f
C271 B.n231 VSUBS 0.007653f
C272 B.n232 VSUBS 0.007653f
C273 B.n233 VSUBS 0.007653f
C274 B.n234 VSUBS 0.007653f
C275 B.n235 VSUBS 0.007653f
C276 B.n236 VSUBS 0.007653f
C277 B.n237 VSUBS 0.007653f
C278 B.n238 VSUBS 0.007653f
C279 B.n239 VSUBS 0.007653f
C280 B.n240 VSUBS 0.007653f
C281 B.n241 VSUBS 0.007653f
C282 B.n242 VSUBS 0.007653f
C283 B.n243 VSUBS 0.007653f
C284 B.n244 VSUBS 0.007653f
C285 B.n245 VSUBS 0.007653f
C286 B.n246 VSUBS 0.007653f
C287 B.n247 VSUBS 0.007653f
C288 B.n248 VSUBS 0.007653f
C289 B.n249 VSUBS 0.007653f
C290 B.n250 VSUBS 0.007653f
C291 B.n251 VSUBS 0.007653f
C292 B.n252 VSUBS 0.007653f
C293 B.n253 VSUBS 0.019441f
C294 B.n254 VSUBS 0.007653f
C295 B.n255 VSUBS 0.007653f
C296 B.n256 VSUBS 0.007653f
C297 B.n257 VSUBS 0.007653f
C298 B.n258 VSUBS 0.007653f
C299 B.n259 VSUBS 0.007653f
C300 B.n260 VSUBS 0.007653f
C301 B.n261 VSUBS 0.007653f
C302 B.n262 VSUBS 0.007653f
C303 B.n263 VSUBS 0.007653f
C304 B.n264 VSUBS 0.007653f
C305 B.n265 VSUBS 0.007653f
C306 B.n266 VSUBS 0.007653f
C307 B.n267 VSUBS 0.007653f
C308 B.n268 VSUBS 0.007653f
C309 B.n269 VSUBS 0.007653f
C310 B.n270 VSUBS 0.007653f
C311 B.n271 VSUBS 0.007653f
C312 B.n272 VSUBS 0.007653f
C313 B.n273 VSUBS 0.007653f
C314 B.n274 VSUBS 0.007653f
C315 B.n275 VSUBS 0.007653f
C316 B.n276 VSUBS 0.007653f
C317 B.n277 VSUBS 0.007653f
C318 B.n278 VSUBS 0.007653f
C319 B.n279 VSUBS 0.007653f
C320 B.n280 VSUBS 0.007653f
C321 B.n281 VSUBS 0.007653f
C322 B.n282 VSUBS 0.007653f
C323 B.n283 VSUBS 0.007653f
C324 B.n284 VSUBS 0.007653f
C325 B.n285 VSUBS 0.007653f
C326 B.n286 VSUBS 0.007653f
C327 B.n287 VSUBS 0.007653f
C328 B.n288 VSUBS 0.007653f
C329 B.n289 VSUBS 0.007653f
C330 B.n290 VSUBS 0.007653f
C331 B.n291 VSUBS 0.007653f
C332 B.n292 VSUBS 0.007653f
C333 B.n293 VSUBS 0.007653f
C334 B.n294 VSUBS 0.007653f
C335 B.n295 VSUBS 0.007653f
C336 B.n296 VSUBS 0.007653f
C337 B.n297 VSUBS 0.007653f
C338 B.n298 VSUBS 0.007653f
C339 B.n299 VSUBS 0.007653f
C340 B.n300 VSUBS 0.007653f
C341 B.n301 VSUBS 0.007653f
C342 B.n302 VSUBS 0.007653f
C343 B.n303 VSUBS 0.007653f
C344 B.n304 VSUBS 0.007653f
C345 B.n305 VSUBS 0.007653f
C346 B.n306 VSUBS 0.007653f
C347 B.n307 VSUBS 0.007653f
C348 B.n308 VSUBS 0.007653f
C349 B.n309 VSUBS 0.007653f
C350 B.n310 VSUBS 0.007653f
C351 B.n311 VSUBS 0.007653f
C352 B.n312 VSUBS 0.007653f
C353 B.n313 VSUBS 0.007653f
C354 B.n314 VSUBS 0.007653f
C355 B.n315 VSUBS 0.007653f
C356 B.n316 VSUBS 0.007653f
C357 B.n317 VSUBS 0.007653f
C358 B.n318 VSUBS 0.007653f
C359 B.n319 VSUBS 0.007653f
C360 B.n320 VSUBS 0.007653f
C361 B.n321 VSUBS 0.007653f
C362 B.n322 VSUBS 0.007653f
C363 B.n323 VSUBS 0.007653f
C364 B.n324 VSUBS 0.007653f
C365 B.n325 VSUBS 0.007653f
C366 B.n326 VSUBS 0.007653f
C367 B.n327 VSUBS 0.007653f
C368 B.n328 VSUBS 0.007653f
C369 B.n329 VSUBS 0.007653f
C370 B.n330 VSUBS 0.007653f
C371 B.n331 VSUBS 0.007653f
C372 B.n332 VSUBS 0.007653f
C373 B.n333 VSUBS 0.007653f
C374 B.n334 VSUBS 0.007653f
C375 B.n335 VSUBS 0.007653f
C376 B.n336 VSUBS 0.007653f
C377 B.n337 VSUBS 0.007653f
C378 B.n338 VSUBS 0.007653f
C379 B.n339 VSUBS 0.007653f
C380 B.n340 VSUBS 0.007653f
C381 B.n341 VSUBS 0.007653f
C382 B.n342 VSUBS 0.007653f
C383 B.n343 VSUBS 0.007653f
C384 B.n344 VSUBS 0.007653f
C385 B.n345 VSUBS 0.007653f
C386 B.n346 VSUBS 0.007653f
C387 B.n347 VSUBS 0.007653f
C388 B.n348 VSUBS 0.007653f
C389 B.n349 VSUBS 0.007653f
C390 B.n350 VSUBS 0.007653f
C391 B.n351 VSUBS 0.007653f
C392 B.n352 VSUBS 0.007653f
C393 B.n353 VSUBS 0.007653f
C394 B.n354 VSUBS 0.007653f
C395 B.n355 VSUBS 0.007653f
C396 B.n356 VSUBS 0.007653f
C397 B.n357 VSUBS 0.007653f
C398 B.n358 VSUBS 0.007653f
C399 B.n359 VSUBS 0.007653f
C400 B.n360 VSUBS 0.007653f
C401 B.n361 VSUBS 0.007653f
C402 B.n362 VSUBS 0.007653f
C403 B.n363 VSUBS 0.007653f
C404 B.n364 VSUBS 0.007653f
C405 B.n365 VSUBS 0.007653f
C406 B.n366 VSUBS 0.007653f
C407 B.n367 VSUBS 0.007653f
C408 B.n368 VSUBS 0.007653f
C409 B.n369 VSUBS 0.007653f
C410 B.n370 VSUBS 0.007653f
C411 B.n371 VSUBS 0.007653f
C412 B.n372 VSUBS 0.007653f
C413 B.n373 VSUBS 0.007653f
C414 B.n374 VSUBS 0.007653f
C415 B.n375 VSUBS 0.007653f
C416 B.n376 VSUBS 0.007653f
C417 B.n377 VSUBS 0.007653f
C418 B.n378 VSUBS 0.007653f
C419 B.n379 VSUBS 0.007653f
C420 B.n380 VSUBS 0.007653f
C421 B.n381 VSUBS 0.007653f
C422 B.n382 VSUBS 0.007653f
C423 B.n383 VSUBS 0.007653f
C424 B.n384 VSUBS 0.007653f
C425 B.n385 VSUBS 0.007653f
C426 B.n386 VSUBS 0.007653f
C427 B.n387 VSUBS 0.007653f
C428 B.n388 VSUBS 0.007653f
C429 B.n389 VSUBS 0.007653f
C430 B.n390 VSUBS 0.007653f
C431 B.n391 VSUBS 0.007653f
C432 B.n392 VSUBS 0.007653f
C433 B.n393 VSUBS 0.007653f
C434 B.n394 VSUBS 0.007653f
C435 B.n395 VSUBS 0.007653f
C436 B.n396 VSUBS 0.007653f
C437 B.n397 VSUBS 0.007653f
C438 B.n398 VSUBS 0.018822f
C439 B.n399 VSUBS 0.018822f
C440 B.n400 VSUBS 0.019441f
C441 B.n401 VSUBS 0.007653f
C442 B.n402 VSUBS 0.007653f
C443 B.n403 VSUBS 0.007653f
C444 B.n404 VSUBS 0.007653f
C445 B.n405 VSUBS 0.007653f
C446 B.n406 VSUBS 0.007653f
C447 B.n407 VSUBS 0.007653f
C448 B.n408 VSUBS 0.007653f
C449 B.n409 VSUBS 0.007653f
C450 B.n410 VSUBS 0.007653f
C451 B.n411 VSUBS 0.007653f
C452 B.n412 VSUBS 0.007653f
C453 B.n413 VSUBS 0.007653f
C454 B.n414 VSUBS 0.007653f
C455 B.n415 VSUBS 0.007653f
C456 B.n416 VSUBS 0.007653f
C457 B.n417 VSUBS 0.007653f
C458 B.n418 VSUBS 0.007653f
C459 B.n419 VSUBS 0.007653f
C460 B.n420 VSUBS 0.007653f
C461 B.n421 VSUBS 0.007653f
C462 B.n422 VSUBS 0.007653f
C463 B.n423 VSUBS 0.007653f
C464 B.n424 VSUBS 0.007653f
C465 B.n425 VSUBS 0.007653f
C466 B.n426 VSUBS 0.007653f
C467 B.n427 VSUBS 0.007653f
C468 B.n428 VSUBS 0.007653f
C469 B.n429 VSUBS 0.007653f
C470 B.n430 VSUBS 0.007653f
C471 B.n431 VSUBS 0.007653f
C472 B.n432 VSUBS 0.007653f
C473 B.n433 VSUBS 0.007653f
C474 B.n434 VSUBS 0.007653f
C475 B.n435 VSUBS 0.007653f
C476 B.n436 VSUBS 0.007653f
C477 B.n437 VSUBS 0.007653f
C478 B.n438 VSUBS 0.007653f
C479 B.n439 VSUBS 0.007653f
C480 B.n440 VSUBS 0.007653f
C481 B.n441 VSUBS 0.007653f
C482 B.n442 VSUBS 0.007653f
C483 B.n443 VSUBS 0.007653f
C484 B.n444 VSUBS 0.007653f
C485 B.n445 VSUBS 0.007653f
C486 B.n446 VSUBS 0.007653f
C487 B.n447 VSUBS 0.007653f
C488 B.n448 VSUBS 0.007653f
C489 B.n449 VSUBS 0.007653f
C490 B.n450 VSUBS 0.007653f
C491 B.n451 VSUBS 0.007653f
C492 B.n452 VSUBS 0.007653f
C493 B.n453 VSUBS 0.007653f
C494 B.n454 VSUBS 0.007653f
C495 B.n455 VSUBS 0.007653f
C496 B.n456 VSUBS 0.007653f
C497 B.n457 VSUBS 0.007653f
C498 B.n458 VSUBS 0.007653f
C499 B.n459 VSUBS 0.007653f
C500 B.n460 VSUBS 0.007653f
C501 B.n461 VSUBS 0.007653f
C502 B.n462 VSUBS 0.007653f
C503 B.n463 VSUBS 0.007653f
C504 B.n464 VSUBS 0.007653f
C505 B.n465 VSUBS 0.007653f
C506 B.n466 VSUBS 0.007653f
C507 B.n467 VSUBS 0.007653f
C508 B.n468 VSUBS 0.007653f
C509 B.n469 VSUBS 0.007653f
C510 B.n470 VSUBS 0.007653f
C511 B.n471 VSUBS 0.007653f
C512 B.n472 VSUBS 0.007653f
C513 B.n473 VSUBS 0.007653f
C514 B.n474 VSUBS 0.007653f
C515 B.n475 VSUBS 0.007653f
C516 B.n476 VSUBS 0.007653f
C517 B.n477 VSUBS 0.007653f
C518 B.n478 VSUBS 0.007653f
C519 B.n479 VSUBS 0.007653f
C520 B.n480 VSUBS 0.007653f
C521 B.n481 VSUBS 0.007653f
C522 B.n482 VSUBS 0.007653f
C523 B.n483 VSUBS 0.007653f
C524 B.n484 VSUBS 0.007653f
C525 B.n485 VSUBS 0.007653f
C526 B.n486 VSUBS 0.007653f
C527 B.n487 VSUBS 0.007653f
C528 B.n488 VSUBS 0.007653f
C529 B.n489 VSUBS 0.007653f
C530 B.n490 VSUBS 0.005289f
C531 B.n491 VSUBS 0.01773f
C532 B.n492 VSUBS 0.00619f
C533 B.n493 VSUBS 0.007653f
C534 B.n494 VSUBS 0.007653f
C535 B.n495 VSUBS 0.007653f
C536 B.n496 VSUBS 0.007653f
C537 B.n497 VSUBS 0.007653f
C538 B.n498 VSUBS 0.007653f
C539 B.n499 VSUBS 0.007653f
C540 B.n500 VSUBS 0.007653f
C541 B.n501 VSUBS 0.007653f
C542 B.n502 VSUBS 0.007653f
C543 B.n503 VSUBS 0.007653f
C544 B.n504 VSUBS 0.00619f
C545 B.n505 VSUBS 0.007653f
C546 B.n506 VSUBS 0.007653f
C547 B.n507 VSUBS 0.005289f
C548 B.n508 VSUBS 0.007653f
C549 B.n509 VSUBS 0.007653f
C550 B.n510 VSUBS 0.007653f
C551 B.n511 VSUBS 0.007653f
C552 B.n512 VSUBS 0.007653f
C553 B.n513 VSUBS 0.007653f
C554 B.n514 VSUBS 0.007653f
C555 B.n515 VSUBS 0.007653f
C556 B.n516 VSUBS 0.007653f
C557 B.n517 VSUBS 0.007653f
C558 B.n518 VSUBS 0.007653f
C559 B.n519 VSUBS 0.007653f
C560 B.n520 VSUBS 0.007653f
C561 B.n521 VSUBS 0.007653f
C562 B.n522 VSUBS 0.007653f
C563 B.n523 VSUBS 0.007653f
C564 B.n524 VSUBS 0.007653f
C565 B.n525 VSUBS 0.007653f
C566 B.n526 VSUBS 0.007653f
C567 B.n527 VSUBS 0.007653f
C568 B.n528 VSUBS 0.007653f
C569 B.n529 VSUBS 0.007653f
C570 B.n530 VSUBS 0.007653f
C571 B.n531 VSUBS 0.007653f
C572 B.n532 VSUBS 0.007653f
C573 B.n533 VSUBS 0.007653f
C574 B.n534 VSUBS 0.007653f
C575 B.n535 VSUBS 0.007653f
C576 B.n536 VSUBS 0.007653f
C577 B.n537 VSUBS 0.007653f
C578 B.n538 VSUBS 0.007653f
C579 B.n539 VSUBS 0.007653f
C580 B.n540 VSUBS 0.007653f
C581 B.n541 VSUBS 0.007653f
C582 B.n542 VSUBS 0.007653f
C583 B.n543 VSUBS 0.007653f
C584 B.n544 VSUBS 0.007653f
C585 B.n545 VSUBS 0.007653f
C586 B.n546 VSUBS 0.007653f
C587 B.n547 VSUBS 0.007653f
C588 B.n548 VSUBS 0.007653f
C589 B.n549 VSUBS 0.007653f
C590 B.n550 VSUBS 0.007653f
C591 B.n551 VSUBS 0.007653f
C592 B.n552 VSUBS 0.007653f
C593 B.n553 VSUBS 0.007653f
C594 B.n554 VSUBS 0.007653f
C595 B.n555 VSUBS 0.007653f
C596 B.n556 VSUBS 0.007653f
C597 B.n557 VSUBS 0.007653f
C598 B.n558 VSUBS 0.007653f
C599 B.n559 VSUBS 0.007653f
C600 B.n560 VSUBS 0.007653f
C601 B.n561 VSUBS 0.007653f
C602 B.n562 VSUBS 0.007653f
C603 B.n563 VSUBS 0.007653f
C604 B.n564 VSUBS 0.007653f
C605 B.n565 VSUBS 0.007653f
C606 B.n566 VSUBS 0.007653f
C607 B.n567 VSUBS 0.007653f
C608 B.n568 VSUBS 0.007653f
C609 B.n569 VSUBS 0.007653f
C610 B.n570 VSUBS 0.007653f
C611 B.n571 VSUBS 0.007653f
C612 B.n572 VSUBS 0.007653f
C613 B.n573 VSUBS 0.007653f
C614 B.n574 VSUBS 0.007653f
C615 B.n575 VSUBS 0.007653f
C616 B.n576 VSUBS 0.007653f
C617 B.n577 VSUBS 0.007653f
C618 B.n578 VSUBS 0.007653f
C619 B.n579 VSUBS 0.007653f
C620 B.n580 VSUBS 0.007653f
C621 B.n581 VSUBS 0.007653f
C622 B.n582 VSUBS 0.007653f
C623 B.n583 VSUBS 0.007653f
C624 B.n584 VSUBS 0.007653f
C625 B.n585 VSUBS 0.007653f
C626 B.n586 VSUBS 0.007653f
C627 B.n587 VSUBS 0.007653f
C628 B.n588 VSUBS 0.007653f
C629 B.n589 VSUBS 0.007653f
C630 B.n590 VSUBS 0.007653f
C631 B.n591 VSUBS 0.007653f
C632 B.n592 VSUBS 0.007653f
C633 B.n593 VSUBS 0.007653f
C634 B.n594 VSUBS 0.007653f
C635 B.n595 VSUBS 0.007653f
C636 B.n596 VSUBS 0.019441f
C637 B.n597 VSUBS 0.019441f
C638 B.n598 VSUBS 0.018822f
C639 B.n599 VSUBS 0.007653f
C640 B.n600 VSUBS 0.007653f
C641 B.n601 VSUBS 0.007653f
C642 B.n602 VSUBS 0.007653f
C643 B.n603 VSUBS 0.007653f
C644 B.n604 VSUBS 0.007653f
C645 B.n605 VSUBS 0.007653f
C646 B.n606 VSUBS 0.007653f
C647 B.n607 VSUBS 0.007653f
C648 B.n608 VSUBS 0.007653f
C649 B.n609 VSUBS 0.007653f
C650 B.n610 VSUBS 0.007653f
C651 B.n611 VSUBS 0.007653f
C652 B.n612 VSUBS 0.007653f
C653 B.n613 VSUBS 0.007653f
C654 B.n614 VSUBS 0.007653f
C655 B.n615 VSUBS 0.007653f
C656 B.n616 VSUBS 0.007653f
C657 B.n617 VSUBS 0.007653f
C658 B.n618 VSUBS 0.007653f
C659 B.n619 VSUBS 0.007653f
C660 B.n620 VSUBS 0.007653f
C661 B.n621 VSUBS 0.007653f
C662 B.n622 VSUBS 0.007653f
C663 B.n623 VSUBS 0.007653f
C664 B.n624 VSUBS 0.007653f
C665 B.n625 VSUBS 0.007653f
C666 B.n626 VSUBS 0.007653f
C667 B.n627 VSUBS 0.007653f
C668 B.n628 VSUBS 0.007653f
C669 B.n629 VSUBS 0.007653f
C670 B.n630 VSUBS 0.007653f
C671 B.n631 VSUBS 0.007653f
C672 B.n632 VSUBS 0.007653f
C673 B.n633 VSUBS 0.007653f
C674 B.n634 VSUBS 0.007653f
C675 B.n635 VSUBS 0.007653f
C676 B.n636 VSUBS 0.007653f
C677 B.n637 VSUBS 0.007653f
C678 B.n638 VSUBS 0.007653f
C679 B.n639 VSUBS 0.007653f
C680 B.n640 VSUBS 0.007653f
C681 B.n641 VSUBS 0.007653f
C682 B.n642 VSUBS 0.007653f
C683 B.n643 VSUBS 0.007653f
C684 B.n644 VSUBS 0.007653f
C685 B.n645 VSUBS 0.007653f
C686 B.n646 VSUBS 0.007653f
C687 B.n647 VSUBS 0.007653f
C688 B.n648 VSUBS 0.007653f
C689 B.n649 VSUBS 0.007653f
C690 B.n650 VSUBS 0.007653f
C691 B.n651 VSUBS 0.007653f
C692 B.n652 VSUBS 0.007653f
C693 B.n653 VSUBS 0.007653f
C694 B.n654 VSUBS 0.007653f
C695 B.n655 VSUBS 0.007653f
C696 B.n656 VSUBS 0.007653f
C697 B.n657 VSUBS 0.007653f
C698 B.n658 VSUBS 0.007653f
C699 B.n659 VSUBS 0.007653f
C700 B.n660 VSUBS 0.007653f
C701 B.n661 VSUBS 0.007653f
C702 B.n662 VSUBS 0.007653f
C703 B.n663 VSUBS 0.007653f
C704 B.n664 VSUBS 0.007653f
C705 B.n665 VSUBS 0.007653f
C706 B.n666 VSUBS 0.007653f
C707 B.n667 VSUBS 0.007653f
C708 B.n668 VSUBS 0.007653f
C709 B.n669 VSUBS 0.007653f
C710 B.n670 VSUBS 0.007653f
C711 B.n671 VSUBS 0.007653f
C712 B.n672 VSUBS 0.007653f
C713 B.n673 VSUBS 0.007653f
C714 B.n674 VSUBS 0.007653f
C715 B.n675 VSUBS 0.007653f
C716 B.n676 VSUBS 0.007653f
C717 B.n677 VSUBS 0.007653f
C718 B.n678 VSUBS 0.007653f
C719 B.n679 VSUBS 0.007653f
C720 B.n680 VSUBS 0.007653f
C721 B.n681 VSUBS 0.007653f
C722 B.n682 VSUBS 0.007653f
C723 B.n683 VSUBS 0.007653f
C724 B.n684 VSUBS 0.007653f
C725 B.n685 VSUBS 0.007653f
C726 B.n686 VSUBS 0.007653f
C727 B.n687 VSUBS 0.007653f
C728 B.n688 VSUBS 0.007653f
C729 B.n689 VSUBS 0.007653f
C730 B.n690 VSUBS 0.007653f
C731 B.n691 VSUBS 0.007653f
C732 B.n692 VSUBS 0.007653f
C733 B.n693 VSUBS 0.007653f
C734 B.n694 VSUBS 0.007653f
C735 B.n695 VSUBS 0.007653f
C736 B.n696 VSUBS 0.007653f
C737 B.n697 VSUBS 0.007653f
C738 B.n698 VSUBS 0.007653f
C739 B.n699 VSUBS 0.007653f
C740 B.n700 VSUBS 0.007653f
C741 B.n701 VSUBS 0.007653f
C742 B.n702 VSUBS 0.007653f
C743 B.n703 VSUBS 0.007653f
C744 B.n704 VSUBS 0.007653f
C745 B.n705 VSUBS 0.007653f
C746 B.n706 VSUBS 0.007653f
C747 B.n707 VSUBS 0.007653f
C748 B.n708 VSUBS 0.007653f
C749 B.n709 VSUBS 0.007653f
C750 B.n710 VSUBS 0.007653f
C751 B.n711 VSUBS 0.007653f
C752 B.n712 VSUBS 0.007653f
C753 B.n713 VSUBS 0.007653f
C754 B.n714 VSUBS 0.007653f
C755 B.n715 VSUBS 0.007653f
C756 B.n716 VSUBS 0.007653f
C757 B.n717 VSUBS 0.007653f
C758 B.n718 VSUBS 0.007653f
C759 B.n719 VSUBS 0.007653f
C760 B.n720 VSUBS 0.007653f
C761 B.n721 VSUBS 0.007653f
C762 B.n722 VSUBS 0.007653f
C763 B.n723 VSUBS 0.007653f
C764 B.n724 VSUBS 0.007653f
C765 B.n725 VSUBS 0.007653f
C766 B.n726 VSUBS 0.007653f
C767 B.n727 VSUBS 0.007653f
C768 B.n728 VSUBS 0.007653f
C769 B.n729 VSUBS 0.007653f
C770 B.n730 VSUBS 0.007653f
C771 B.n731 VSUBS 0.007653f
C772 B.n732 VSUBS 0.007653f
C773 B.n733 VSUBS 0.007653f
C774 B.n734 VSUBS 0.007653f
C775 B.n735 VSUBS 0.007653f
C776 B.n736 VSUBS 0.007653f
C777 B.n737 VSUBS 0.007653f
C778 B.n738 VSUBS 0.007653f
C779 B.n739 VSUBS 0.007653f
C780 B.n740 VSUBS 0.007653f
C781 B.n741 VSUBS 0.007653f
C782 B.n742 VSUBS 0.007653f
C783 B.n743 VSUBS 0.007653f
C784 B.n744 VSUBS 0.007653f
C785 B.n745 VSUBS 0.007653f
C786 B.n746 VSUBS 0.007653f
C787 B.n747 VSUBS 0.007653f
C788 B.n748 VSUBS 0.007653f
C789 B.n749 VSUBS 0.007653f
C790 B.n750 VSUBS 0.007653f
C791 B.n751 VSUBS 0.007653f
C792 B.n752 VSUBS 0.007653f
C793 B.n753 VSUBS 0.007653f
C794 B.n754 VSUBS 0.007653f
C795 B.n755 VSUBS 0.007653f
C796 B.n756 VSUBS 0.007653f
C797 B.n757 VSUBS 0.007653f
C798 B.n758 VSUBS 0.007653f
C799 B.n759 VSUBS 0.007653f
C800 B.n760 VSUBS 0.007653f
C801 B.n761 VSUBS 0.007653f
C802 B.n762 VSUBS 0.007653f
C803 B.n763 VSUBS 0.007653f
C804 B.n764 VSUBS 0.007653f
C805 B.n765 VSUBS 0.007653f
C806 B.n766 VSUBS 0.007653f
C807 B.n767 VSUBS 0.007653f
C808 B.n768 VSUBS 0.007653f
C809 B.n769 VSUBS 0.007653f
C810 B.n770 VSUBS 0.007653f
C811 B.n771 VSUBS 0.007653f
C812 B.n772 VSUBS 0.007653f
C813 B.n773 VSUBS 0.007653f
C814 B.n774 VSUBS 0.007653f
C815 B.n775 VSUBS 0.007653f
C816 B.n776 VSUBS 0.007653f
C817 B.n777 VSUBS 0.007653f
C818 B.n778 VSUBS 0.007653f
C819 B.n779 VSUBS 0.007653f
C820 B.n780 VSUBS 0.007653f
C821 B.n781 VSUBS 0.007653f
C822 B.n782 VSUBS 0.007653f
C823 B.n783 VSUBS 0.007653f
C824 B.n784 VSUBS 0.007653f
C825 B.n785 VSUBS 0.007653f
C826 B.n786 VSUBS 0.007653f
C827 B.n787 VSUBS 0.007653f
C828 B.n788 VSUBS 0.007653f
C829 B.n789 VSUBS 0.007653f
C830 B.n790 VSUBS 0.007653f
C831 B.n791 VSUBS 0.007653f
C832 B.n792 VSUBS 0.007653f
C833 B.n793 VSUBS 0.007653f
C834 B.n794 VSUBS 0.007653f
C835 B.n795 VSUBS 0.007653f
C836 B.n796 VSUBS 0.007653f
C837 B.n797 VSUBS 0.007653f
C838 B.n798 VSUBS 0.007653f
C839 B.n799 VSUBS 0.007653f
C840 B.n800 VSUBS 0.007653f
C841 B.n801 VSUBS 0.007653f
C842 B.n802 VSUBS 0.007653f
C843 B.n803 VSUBS 0.007653f
C844 B.n804 VSUBS 0.007653f
C845 B.n805 VSUBS 0.007653f
C846 B.n806 VSUBS 0.007653f
C847 B.n807 VSUBS 0.007653f
C848 B.n808 VSUBS 0.007653f
C849 B.n809 VSUBS 0.007653f
C850 B.n810 VSUBS 0.007653f
C851 B.n811 VSUBS 0.007653f
C852 B.n812 VSUBS 0.007653f
C853 B.n813 VSUBS 0.007653f
C854 B.n814 VSUBS 0.007653f
C855 B.n815 VSUBS 0.007653f
C856 B.n816 VSUBS 0.007653f
C857 B.n817 VSUBS 0.007653f
C858 B.n818 VSUBS 0.007653f
C859 B.n819 VSUBS 0.007653f
C860 B.n820 VSUBS 0.019641f
C861 B.n821 VSUBS 0.018622f
C862 B.n822 VSUBS 0.019441f
C863 B.n823 VSUBS 0.007653f
C864 B.n824 VSUBS 0.007653f
C865 B.n825 VSUBS 0.007653f
C866 B.n826 VSUBS 0.007653f
C867 B.n827 VSUBS 0.007653f
C868 B.n828 VSUBS 0.007653f
C869 B.n829 VSUBS 0.007653f
C870 B.n830 VSUBS 0.007653f
C871 B.n831 VSUBS 0.007653f
C872 B.n832 VSUBS 0.007653f
C873 B.n833 VSUBS 0.007653f
C874 B.n834 VSUBS 0.007653f
C875 B.n835 VSUBS 0.007653f
C876 B.n836 VSUBS 0.007653f
C877 B.n837 VSUBS 0.007653f
C878 B.n838 VSUBS 0.007653f
C879 B.n839 VSUBS 0.007653f
C880 B.n840 VSUBS 0.007653f
C881 B.n841 VSUBS 0.007653f
C882 B.n842 VSUBS 0.007653f
C883 B.n843 VSUBS 0.007653f
C884 B.n844 VSUBS 0.007653f
C885 B.n845 VSUBS 0.007653f
C886 B.n846 VSUBS 0.007653f
C887 B.n847 VSUBS 0.007653f
C888 B.n848 VSUBS 0.007653f
C889 B.n849 VSUBS 0.007653f
C890 B.n850 VSUBS 0.007653f
C891 B.n851 VSUBS 0.007653f
C892 B.n852 VSUBS 0.007653f
C893 B.n853 VSUBS 0.007653f
C894 B.n854 VSUBS 0.007653f
C895 B.n855 VSUBS 0.007653f
C896 B.n856 VSUBS 0.007653f
C897 B.n857 VSUBS 0.007653f
C898 B.n858 VSUBS 0.007653f
C899 B.n859 VSUBS 0.007653f
C900 B.n860 VSUBS 0.007653f
C901 B.n861 VSUBS 0.007653f
C902 B.n862 VSUBS 0.007653f
C903 B.n863 VSUBS 0.007653f
C904 B.n864 VSUBS 0.007653f
C905 B.n865 VSUBS 0.007653f
C906 B.n866 VSUBS 0.007653f
C907 B.n867 VSUBS 0.007653f
C908 B.n868 VSUBS 0.007653f
C909 B.n869 VSUBS 0.007653f
C910 B.n870 VSUBS 0.007653f
C911 B.n871 VSUBS 0.007653f
C912 B.n872 VSUBS 0.007653f
C913 B.n873 VSUBS 0.007653f
C914 B.n874 VSUBS 0.007653f
C915 B.n875 VSUBS 0.007653f
C916 B.n876 VSUBS 0.007653f
C917 B.n877 VSUBS 0.007653f
C918 B.n878 VSUBS 0.007653f
C919 B.n879 VSUBS 0.007653f
C920 B.n880 VSUBS 0.007653f
C921 B.n881 VSUBS 0.007653f
C922 B.n882 VSUBS 0.007653f
C923 B.n883 VSUBS 0.007653f
C924 B.n884 VSUBS 0.007653f
C925 B.n885 VSUBS 0.007653f
C926 B.n886 VSUBS 0.007653f
C927 B.n887 VSUBS 0.007653f
C928 B.n888 VSUBS 0.007653f
C929 B.n889 VSUBS 0.007653f
C930 B.n890 VSUBS 0.007653f
C931 B.n891 VSUBS 0.007653f
C932 B.n892 VSUBS 0.007653f
C933 B.n893 VSUBS 0.007653f
C934 B.n894 VSUBS 0.007653f
C935 B.n895 VSUBS 0.007653f
C936 B.n896 VSUBS 0.007653f
C937 B.n897 VSUBS 0.007653f
C938 B.n898 VSUBS 0.007653f
C939 B.n899 VSUBS 0.007653f
C940 B.n900 VSUBS 0.007653f
C941 B.n901 VSUBS 0.007653f
C942 B.n902 VSUBS 0.007653f
C943 B.n903 VSUBS 0.007653f
C944 B.n904 VSUBS 0.007653f
C945 B.n905 VSUBS 0.007653f
C946 B.n906 VSUBS 0.007653f
C947 B.n907 VSUBS 0.007653f
C948 B.n908 VSUBS 0.007653f
C949 B.n909 VSUBS 0.007653f
C950 B.n910 VSUBS 0.007653f
C951 B.n911 VSUBS 0.005289f
C952 B.n912 VSUBS 0.007653f
C953 B.n913 VSUBS 0.007653f
C954 B.n914 VSUBS 0.00619f
C955 B.n915 VSUBS 0.007653f
C956 B.n916 VSUBS 0.007653f
C957 B.n917 VSUBS 0.007653f
C958 B.n918 VSUBS 0.007653f
C959 B.n919 VSUBS 0.007653f
C960 B.n920 VSUBS 0.007653f
C961 B.n921 VSUBS 0.007653f
C962 B.n922 VSUBS 0.007653f
C963 B.n923 VSUBS 0.007653f
C964 B.n924 VSUBS 0.007653f
C965 B.n925 VSUBS 0.007653f
C966 B.n926 VSUBS 0.00619f
C967 B.n927 VSUBS 0.01773f
C968 B.n928 VSUBS 0.005289f
C969 B.n929 VSUBS 0.007653f
C970 B.n930 VSUBS 0.007653f
C971 B.n931 VSUBS 0.007653f
C972 B.n932 VSUBS 0.007653f
C973 B.n933 VSUBS 0.007653f
C974 B.n934 VSUBS 0.007653f
C975 B.n935 VSUBS 0.007653f
C976 B.n936 VSUBS 0.007653f
C977 B.n937 VSUBS 0.007653f
C978 B.n938 VSUBS 0.007653f
C979 B.n939 VSUBS 0.007653f
C980 B.n940 VSUBS 0.007653f
C981 B.n941 VSUBS 0.007653f
C982 B.n942 VSUBS 0.007653f
C983 B.n943 VSUBS 0.007653f
C984 B.n944 VSUBS 0.007653f
C985 B.n945 VSUBS 0.007653f
C986 B.n946 VSUBS 0.007653f
C987 B.n947 VSUBS 0.007653f
C988 B.n948 VSUBS 0.007653f
C989 B.n949 VSUBS 0.007653f
C990 B.n950 VSUBS 0.007653f
C991 B.n951 VSUBS 0.007653f
C992 B.n952 VSUBS 0.007653f
C993 B.n953 VSUBS 0.007653f
C994 B.n954 VSUBS 0.007653f
C995 B.n955 VSUBS 0.007653f
C996 B.n956 VSUBS 0.007653f
C997 B.n957 VSUBS 0.007653f
C998 B.n958 VSUBS 0.007653f
C999 B.n959 VSUBS 0.007653f
C1000 B.n960 VSUBS 0.007653f
C1001 B.n961 VSUBS 0.007653f
C1002 B.n962 VSUBS 0.007653f
C1003 B.n963 VSUBS 0.007653f
C1004 B.n964 VSUBS 0.007653f
C1005 B.n965 VSUBS 0.007653f
C1006 B.n966 VSUBS 0.007653f
C1007 B.n967 VSUBS 0.007653f
C1008 B.n968 VSUBS 0.007653f
C1009 B.n969 VSUBS 0.007653f
C1010 B.n970 VSUBS 0.007653f
C1011 B.n971 VSUBS 0.007653f
C1012 B.n972 VSUBS 0.007653f
C1013 B.n973 VSUBS 0.007653f
C1014 B.n974 VSUBS 0.007653f
C1015 B.n975 VSUBS 0.007653f
C1016 B.n976 VSUBS 0.007653f
C1017 B.n977 VSUBS 0.007653f
C1018 B.n978 VSUBS 0.007653f
C1019 B.n979 VSUBS 0.007653f
C1020 B.n980 VSUBS 0.007653f
C1021 B.n981 VSUBS 0.007653f
C1022 B.n982 VSUBS 0.007653f
C1023 B.n983 VSUBS 0.007653f
C1024 B.n984 VSUBS 0.007653f
C1025 B.n985 VSUBS 0.007653f
C1026 B.n986 VSUBS 0.007653f
C1027 B.n987 VSUBS 0.007653f
C1028 B.n988 VSUBS 0.007653f
C1029 B.n989 VSUBS 0.007653f
C1030 B.n990 VSUBS 0.007653f
C1031 B.n991 VSUBS 0.007653f
C1032 B.n992 VSUBS 0.007653f
C1033 B.n993 VSUBS 0.007653f
C1034 B.n994 VSUBS 0.007653f
C1035 B.n995 VSUBS 0.007653f
C1036 B.n996 VSUBS 0.007653f
C1037 B.n997 VSUBS 0.007653f
C1038 B.n998 VSUBS 0.007653f
C1039 B.n999 VSUBS 0.007653f
C1040 B.n1000 VSUBS 0.007653f
C1041 B.n1001 VSUBS 0.007653f
C1042 B.n1002 VSUBS 0.007653f
C1043 B.n1003 VSUBS 0.007653f
C1044 B.n1004 VSUBS 0.007653f
C1045 B.n1005 VSUBS 0.007653f
C1046 B.n1006 VSUBS 0.007653f
C1047 B.n1007 VSUBS 0.007653f
C1048 B.n1008 VSUBS 0.007653f
C1049 B.n1009 VSUBS 0.007653f
C1050 B.n1010 VSUBS 0.007653f
C1051 B.n1011 VSUBS 0.007653f
C1052 B.n1012 VSUBS 0.007653f
C1053 B.n1013 VSUBS 0.007653f
C1054 B.n1014 VSUBS 0.007653f
C1055 B.n1015 VSUBS 0.007653f
C1056 B.n1016 VSUBS 0.007653f
C1057 B.n1017 VSUBS 0.007653f
C1058 B.n1018 VSUBS 0.019441f
C1059 B.n1019 VSUBS 0.018822f
C1060 B.n1020 VSUBS 0.018822f
C1061 B.n1021 VSUBS 0.007653f
C1062 B.n1022 VSUBS 0.007653f
C1063 B.n1023 VSUBS 0.007653f
C1064 B.n1024 VSUBS 0.007653f
C1065 B.n1025 VSUBS 0.007653f
C1066 B.n1026 VSUBS 0.007653f
C1067 B.n1027 VSUBS 0.007653f
C1068 B.n1028 VSUBS 0.007653f
C1069 B.n1029 VSUBS 0.007653f
C1070 B.n1030 VSUBS 0.007653f
C1071 B.n1031 VSUBS 0.007653f
C1072 B.n1032 VSUBS 0.007653f
C1073 B.n1033 VSUBS 0.007653f
C1074 B.n1034 VSUBS 0.007653f
C1075 B.n1035 VSUBS 0.007653f
C1076 B.n1036 VSUBS 0.007653f
C1077 B.n1037 VSUBS 0.007653f
C1078 B.n1038 VSUBS 0.007653f
C1079 B.n1039 VSUBS 0.007653f
C1080 B.n1040 VSUBS 0.007653f
C1081 B.n1041 VSUBS 0.007653f
C1082 B.n1042 VSUBS 0.007653f
C1083 B.n1043 VSUBS 0.007653f
C1084 B.n1044 VSUBS 0.007653f
C1085 B.n1045 VSUBS 0.007653f
C1086 B.n1046 VSUBS 0.007653f
C1087 B.n1047 VSUBS 0.007653f
C1088 B.n1048 VSUBS 0.007653f
C1089 B.n1049 VSUBS 0.007653f
C1090 B.n1050 VSUBS 0.007653f
C1091 B.n1051 VSUBS 0.007653f
C1092 B.n1052 VSUBS 0.007653f
C1093 B.n1053 VSUBS 0.007653f
C1094 B.n1054 VSUBS 0.007653f
C1095 B.n1055 VSUBS 0.007653f
C1096 B.n1056 VSUBS 0.007653f
C1097 B.n1057 VSUBS 0.007653f
C1098 B.n1058 VSUBS 0.007653f
C1099 B.n1059 VSUBS 0.007653f
C1100 B.n1060 VSUBS 0.007653f
C1101 B.n1061 VSUBS 0.007653f
C1102 B.n1062 VSUBS 0.007653f
C1103 B.n1063 VSUBS 0.007653f
C1104 B.n1064 VSUBS 0.007653f
C1105 B.n1065 VSUBS 0.007653f
C1106 B.n1066 VSUBS 0.007653f
C1107 B.n1067 VSUBS 0.007653f
C1108 B.n1068 VSUBS 0.007653f
C1109 B.n1069 VSUBS 0.007653f
C1110 B.n1070 VSUBS 0.007653f
C1111 B.n1071 VSUBS 0.007653f
C1112 B.n1072 VSUBS 0.007653f
C1113 B.n1073 VSUBS 0.007653f
C1114 B.n1074 VSUBS 0.007653f
C1115 B.n1075 VSUBS 0.007653f
C1116 B.n1076 VSUBS 0.007653f
C1117 B.n1077 VSUBS 0.007653f
C1118 B.n1078 VSUBS 0.007653f
C1119 B.n1079 VSUBS 0.007653f
C1120 B.n1080 VSUBS 0.007653f
C1121 B.n1081 VSUBS 0.007653f
C1122 B.n1082 VSUBS 0.007653f
C1123 B.n1083 VSUBS 0.007653f
C1124 B.n1084 VSUBS 0.007653f
C1125 B.n1085 VSUBS 0.007653f
C1126 B.n1086 VSUBS 0.007653f
C1127 B.n1087 VSUBS 0.007653f
C1128 B.n1088 VSUBS 0.007653f
C1129 B.n1089 VSUBS 0.007653f
C1130 B.n1090 VSUBS 0.007653f
C1131 B.n1091 VSUBS 0.007653f
C1132 B.n1092 VSUBS 0.007653f
C1133 B.n1093 VSUBS 0.007653f
C1134 B.n1094 VSUBS 0.007653f
C1135 B.n1095 VSUBS 0.007653f
C1136 B.n1096 VSUBS 0.007653f
C1137 B.n1097 VSUBS 0.007653f
C1138 B.n1098 VSUBS 0.007653f
C1139 B.n1099 VSUBS 0.007653f
C1140 B.n1100 VSUBS 0.007653f
C1141 B.n1101 VSUBS 0.007653f
C1142 B.n1102 VSUBS 0.007653f
C1143 B.n1103 VSUBS 0.007653f
C1144 B.n1104 VSUBS 0.007653f
C1145 B.n1105 VSUBS 0.007653f
C1146 B.n1106 VSUBS 0.007653f
C1147 B.n1107 VSUBS 0.007653f
C1148 B.n1108 VSUBS 0.007653f
C1149 B.n1109 VSUBS 0.007653f
C1150 B.n1110 VSUBS 0.007653f
C1151 B.n1111 VSUBS 0.007653f
C1152 B.n1112 VSUBS 0.007653f
C1153 B.n1113 VSUBS 0.007653f
C1154 B.n1114 VSUBS 0.007653f
C1155 B.n1115 VSUBS 0.007653f
C1156 B.n1116 VSUBS 0.007653f
C1157 B.n1117 VSUBS 0.007653f
C1158 B.n1118 VSUBS 0.007653f
C1159 B.n1119 VSUBS 0.007653f
C1160 B.n1120 VSUBS 0.007653f
C1161 B.n1121 VSUBS 0.007653f
C1162 B.n1122 VSUBS 0.007653f
C1163 B.n1123 VSUBS 0.007653f
C1164 B.n1124 VSUBS 0.007653f
C1165 B.n1125 VSUBS 0.007653f
C1166 B.n1126 VSUBS 0.007653f
C1167 B.n1127 VSUBS 0.007653f
C1168 B.n1128 VSUBS 0.007653f
C1169 B.n1129 VSUBS 0.007653f
C1170 B.n1130 VSUBS 0.007653f
C1171 B.n1131 VSUBS 0.017328f
C1172 VDD1.t9 VSUBS 4.60128f
C1173 VDD1.t7 VSUBS 0.421858f
C1174 VDD1.t4 VSUBS 0.421858f
C1175 VDD1.n0 VSUBS 3.51349f
C1176 VDD1.n1 VSUBS 1.89909f
C1177 VDD1.t6 VSUBS 4.60125f
C1178 VDD1.t5 VSUBS 0.421858f
C1179 VDD1.t1 VSUBS 0.421858f
C1180 VDD1.n2 VSUBS 3.51348f
C1181 VDD1.n3 VSUBS 1.88949f
C1182 VDD1.t3 VSUBS 0.421858f
C1183 VDD1.t0 VSUBS 0.421858f
C1184 VDD1.n4 VSUBS 3.55055f
C1185 VDD1.n5 VSUBS 4.80392f
C1186 VDD1.t2 VSUBS 0.421858f
C1187 VDD1.t8 VSUBS 0.421858f
C1188 VDD1.n6 VSUBS 3.51347f
C1189 VDD1.n7 VSUBS 4.94044f
C1190 VP.t9 VSUBS 4.00595f
C1191 VP.n0 VSUBS 1.46915f
C1192 VP.n1 VSUBS 0.022986f
C1193 VP.n2 VSUBS 0.025104f
C1194 VP.n3 VSUBS 0.022986f
C1195 VP.n4 VSUBS 0.022113f
C1196 VP.n5 VSUBS 0.022986f
C1197 VP.n6 VSUBS 0.023217f
C1198 VP.n7 VSUBS 0.022986f
C1199 VP.t8 VSUBS 4.00595f
C1200 VP.n8 VSUBS 1.38087f
C1201 VP.n9 VSUBS 0.022986f
C1202 VP.n10 VSUBS 0.023217f
C1203 VP.n11 VSUBS 0.022986f
C1204 VP.t4 VSUBS 4.00595f
C1205 VP.n12 VSUBS 1.38087f
C1206 VP.n13 VSUBS 0.022986f
C1207 VP.n14 VSUBS 0.04029f
C1208 VP.n15 VSUBS 0.022986f
C1209 VP.n16 VSUBS 0.031419f
C1210 VP.t1 VSUBS 4.00595f
C1211 VP.n17 VSUBS 1.46915f
C1212 VP.n18 VSUBS 0.022986f
C1213 VP.n19 VSUBS 0.025104f
C1214 VP.n20 VSUBS 0.022986f
C1215 VP.n21 VSUBS 0.022113f
C1216 VP.n22 VSUBS 0.022986f
C1217 VP.n23 VSUBS 0.023217f
C1218 VP.n24 VSUBS 0.022986f
C1219 VP.t5 VSUBS 4.00595f
C1220 VP.n25 VSUBS 1.38087f
C1221 VP.n26 VSUBS 0.022986f
C1222 VP.n27 VSUBS 0.023217f
C1223 VP.n28 VSUBS 0.022986f
C1224 VP.t2 VSUBS 4.00595f
C1225 VP.n29 VSUBS 1.47116f
C1226 VP.t0 VSUBS 4.32236f
C1227 VP.n30 VSUBS 1.40072f
C1228 VP.n31 VSUBS 0.280976f
C1229 VP.n32 VSUBS 0.042417f
C1230 VP.n33 VSUBS 0.04284f
C1231 VP.n34 VSUBS 0.041267f
C1232 VP.n35 VSUBS 0.022986f
C1233 VP.n36 VSUBS 0.022986f
C1234 VP.n37 VSUBS 0.022986f
C1235 VP.n38 VSUBS 0.045468f
C1236 VP.n39 VSUBS 0.04284f
C1237 VP.n40 VSUBS 0.032265f
C1238 VP.n41 VSUBS 0.022986f
C1239 VP.n42 VSUBS 0.022986f
C1240 VP.n43 VSUBS 0.032265f
C1241 VP.n44 VSUBS 0.04284f
C1242 VP.n45 VSUBS 0.045468f
C1243 VP.n46 VSUBS 0.022986f
C1244 VP.n47 VSUBS 0.022986f
C1245 VP.n48 VSUBS 0.022986f
C1246 VP.n49 VSUBS 0.041267f
C1247 VP.n50 VSUBS 0.04284f
C1248 VP.t7 VSUBS 4.00595f
C1249 VP.n51 VSUBS 1.38087f
C1250 VP.n52 VSUBS 0.042417f
C1251 VP.n53 VSUBS 0.022986f
C1252 VP.n54 VSUBS 0.022986f
C1253 VP.n55 VSUBS 0.022986f
C1254 VP.n56 VSUBS 0.04284f
C1255 VP.n57 VSUBS 0.04284f
C1256 VP.n58 VSUBS 0.04029f
C1257 VP.n59 VSUBS 0.022986f
C1258 VP.n60 VSUBS 0.022986f
C1259 VP.n61 VSUBS 0.022986f
C1260 VP.n62 VSUBS 0.044558f
C1261 VP.n63 VSUBS 0.04284f
C1262 VP.n64 VSUBS 0.031419f
C1263 VP.n65 VSUBS 0.037099f
C1264 VP.n66 VSUBS 1.78402f
C1265 VP.t3 VSUBS 4.00595f
C1266 VP.n67 VSUBS 1.46915f
C1267 VP.n68 VSUBS 1.79722f
C1268 VP.n69 VSUBS 0.037099f
C1269 VP.n70 VSUBS 0.022986f
C1270 VP.n71 VSUBS 0.04284f
C1271 VP.n72 VSUBS 0.044558f
C1272 VP.n73 VSUBS 0.025104f
C1273 VP.n74 VSUBS 0.022986f
C1274 VP.n75 VSUBS 0.022986f
C1275 VP.n76 VSUBS 0.022986f
C1276 VP.n77 VSUBS 0.04284f
C1277 VP.n78 VSUBS 0.04284f
C1278 VP.n79 VSUBS 0.022113f
C1279 VP.n80 VSUBS 0.022986f
C1280 VP.n81 VSUBS 0.022986f
C1281 VP.n82 VSUBS 0.042417f
C1282 VP.n83 VSUBS 0.04284f
C1283 VP.n84 VSUBS 0.041267f
C1284 VP.n85 VSUBS 0.022986f
C1285 VP.n86 VSUBS 0.022986f
C1286 VP.n87 VSUBS 0.022986f
C1287 VP.n88 VSUBS 0.045468f
C1288 VP.n89 VSUBS 0.04284f
C1289 VP.n90 VSUBS 0.032265f
C1290 VP.n91 VSUBS 0.022986f
C1291 VP.n92 VSUBS 0.022986f
C1292 VP.n93 VSUBS 0.032265f
C1293 VP.n94 VSUBS 0.04284f
C1294 VP.n95 VSUBS 0.045468f
C1295 VP.n96 VSUBS 0.022986f
C1296 VP.n97 VSUBS 0.022986f
C1297 VP.n98 VSUBS 0.022986f
C1298 VP.n99 VSUBS 0.041267f
C1299 VP.n100 VSUBS 0.04284f
C1300 VP.t6 VSUBS 4.00595f
C1301 VP.n101 VSUBS 1.38087f
C1302 VP.n102 VSUBS 0.042417f
C1303 VP.n103 VSUBS 0.022986f
C1304 VP.n104 VSUBS 0.022986f
C1305 VP.n105 VSUBS 0.022986f
C1306 VP.n106 VSUBS 0.04284f
C1307 VP.n107 VSUBS 0.04284f
C1308 VP.n108 VSUBS 0.04029f
C1309 VP.n109 VSUBS 0.022986f
C1310 VP.n110 VSUBS 0.022986f
C1311 VP.n111 VSUBS 0.022986f
C1312 VP.n112 VSUBS 0.044558f
C1313 VP.n113 VSUBS 0.04284f
C1314 VP.n114 VSUBS 0.031419f
C1315 VP.n115 VSUBS 0.037099f
C1316 VP.n116 VSUBS 0.059734f
C1317 VDD2.t3 VSUBS 4.60196f
C1318 VDD2.t8 VSUBS 0.421923f
C1319 VDD2.t6 VSUBS 0.421923f
C1320 VDD2.n0 VSUBS 3.51402f
C1321 VDD2.n1 VSUBS 1.88978f
C1322 VDD2.t0 VSUBS 0.421923f
C1323 VDD2.t9 VSUBS 0.421923f
C1324 VDD2.n2 VSUBS 3.55109f
C1325 VDD2.n3 VSUBS 4.63025f
C1326 VDD2.t2 VSUBS 4.55819f
C1327 VDD2.n4 VSUBS 4.8973f
C1328 VDD2.t5 VSUBS 0.421923f
C1329 VDD2.t7 VSUBS 0.421923f
C1330 VDD2.n5 VSUBS 3.51403f
C1331 VDD2.n6 VSUBS 0.952561f
C1332 VDD2.t1 VSUBS 0.421923f
C1333 VDD2.t4 VSUBS 0.421923f
C1334 VDD2.n7 VSUBS 3.55102f
C1335 VTAIL.t11 VSUBS 0.406823f
C1336 VTAIL.t8 VSUBS 0.406823f
C1337 VTAIL.n0 VSUBS 3.21f
C1338 VTAIL.n1 VSUBS 1.10103f
C1339 VTAIL.t0 VSUBS 4.19033f
C1340 VTAIL.n2 VSUBS 1.29701f
C1341 VTAIL.t1 VSUBS 0.406823f
C1342 VTAIL.t17 VSUBS 0.406823f
C1343 VTAIL.n3 VSUBS 3.21f
C1344 VTAIL.n4 VSUBS 1.26987f
C1345 VTAIL.t3 VSUBS 0.406823f
C1346 VTAIL.t15 VSUBS 0.406823f
C1347 VTAIL.n5 VSUBS 3.21f
C1348 VTAIL.n6 VSUBS 3.36451f
C1349 VTAIL.t14 VSUBS 0.406823f
C1350 VTAIL.t9 VSUBS 0.406823f
C1351 VTAIL.n7 VSUBS 3.21f
C1352 VTAIL.n8 VSUBS 3.3645f
C1353 VTAIL.t10 VSUBS 0.406823f
C1354 VTAIL.t6 VSUBS 0.406823f
C1355 VTAIL.n9 VSUBS 3.21f
C1356 VTAIL.n10 VSUBS 1.26986f
C1357 VTAIL.t13 VSUBS 4.19037f
C1358 VTAIL.n11 VSUBS 1.29698f
C1359 VTAIL.t18 VSUBS 0.406823f
C1360 VTAIL.t4 VSUBS 0.406823f
C1361 VTAIL.n12 VSUBS 3.21f
C1362 VTAIL.n13 VSUBS 1.16782f
C1363 VTAIL.t19 VSUBS 0.406823f
C1364 VTAIL.t2 VSUBS 0.406823f
C1365 VTAIL.n14 VSUBS 3.21f
C1366 VTAIL.n15 VSUBS 1.26986f
C1367 VTAIL.t16 VSUBS 4.19033f
C1368 VTAIL.n16 VSUBS 3.20568f
C1369 VTAIL.t12 VSUBS 4.19033f
C1370 VTAIL.n17 VSUBS 3.20568f
C1371 VTAIL.t7 VSUBS 0.406823f
C1372 VTAIL.t5 VSUBS 0.406823f
C1373 VTAIL.n18 VSUBS 3.21f
C1374 VTAIL.n19 VSUBS 1.04866f
C1375 VN.t0 VSUBS 3.73131f
C1376 VN.n0 VSUBS 1.36843f
C1377 VN.n1 VSUBS 0.02141f
C1378 VN.n2 VSUBS 0.023383f
C1379 VN.n3 VSUBS 0.02141f
C1380 VN.n4 VSUBS 0.020597f
C1381 VN.n5 VSUBS 0.02141f
C1382 VN.n6 VSUBS 0.021625f
C1383 VN.n7 VSUBS 0.02141f
C1384 VN.t3 VSUBS 3.73131f
C1385 VN.n8 VSUBS 1.2862f
C1386 VN.n9 VSUBS 0.02141f
C1387 VN.n10 VSUBS 0.021625f
C1388 VN.n11 VSUBS 0.02141f
C1389 VN.t1 VSUBS 3.73131f
C1390 VN.n12 VSUBS 1.3703f
C1391 VN.t6 VSUBS 4.02603f
C1392 VN.n13 VSUBS 1.30469f
C1393 VN.n14 VSUBS 0.261712f
C1394 VN.n15 VSUBS 0.039509f
C1395 VN.n16 VSUBS 0.039903f
C1396 VN.n17 VSUBS 0.038437f
C1397 VN.n18 VSUBS 0.02141f
C1398 VN.n19 VSUBS 0.02141f
C1399 VN.n20 VSUBS 0.02141f
C1400 VN.n21 VSUBS 0.04235f
C1401 VN.n22 VSUBS 0.039903f
C1402 VN.n23 VSUBS 0.030053f
C1403 VN.n24 VSUBS 0.02141f
C1404 VN.n25 VSUBS 0.02141f
C1405 VN.n26 VSUBS 0.030053f
C1406 VN.n27 VSUBS 0.039903f
C1407 VN.n28 VSUBS 0.04235f
C1408 VN.n29 VSUBS 0.02141f
C1409 VN.n30 VSUBS 0.02141f
C1410 VN.n31 VSUBS 0.02141f
C1411 VN.n32 VSUBS 0.038437f
C1412 VN.n33 VSUBS 0.039903f
C1413 VN.t9 VSUBS 3.73131f
C1414 VN.n34 VSUBS 1.2862f
C1415 VN.n35 VSUBS 0.039509f
C1416 VN.n36 VSUBS 0.02141f
C1417 VN.n37 VSUBS 0.02141f
C1418 VN.n38 VSUBS 0.02141f
C1419 VN.n39 VSUBS 0.039903f
C1420 VN.n40 VSUBS 0.039903f
C1421 VN.n41 VSUBS 0.037528f
C1422 VN.n42 VSUBS 0.02141f
C1423 VN.n43 VSUBS 0.02141f
C1424 VN.n44 VSUBS 0.02141f
C1425 VN.n45 VSUBS 0.041503f
C1426 VN.n46 VSUBS 0.039903f
C1427 VN.n47 VSUBS 0.029265f
C1428 VN.n48 VSUBS 0.034556f
C1429 VN.n49 VSUBS 0.055639f
C1430 VN.t7 VSUBS 3.73131f
C1431 VN.n50 VSUBS 1.36843f
C1432 VN.n51 VSUBS 0.02141f
C1433 VN.n52 VSUBS 0.023383f
C1434 VN.n53 VSUBS 0.02141f
C1435 VN.n54 VSUBS 0.020597f
C1436 VN.n55 VSUBS 0.02141f
C1437 VN.t4 VSUBS 3.73131f
C1438 VN.n56 VSUBS 1.2862f
C1439 VN.n57 VSUBS 0.021625f
C1440 VN.n58 VSUBS 0.02141f
C1441 VN.t2 VSUBS 3.73131f
C1442 VN.n59 VSUBS 1.2862f
C1443 VN.n60 VSUBS 0.02141f
C1444 VN.n61 VSUBS 0.021625f
C1445 VN.n62 VSUBS 0.02141f
C1446 VN.t8 VSUBS 3.73131f
C1447 VN.n63 VSUBS 1.3703f
C1448 VN.t5 VSUBS 4.02603f
C1449 VN.n64 VSUBS 1.30469f
C1450 VN.n65 VSUBS 0.261712f
C1451 VN.n66 VSUBS 0.039509f
C1452 VN.n67 VSUBS 0.039903f
C1453 VN.n68 VSUBS 0.038437f
C1454 VN.n69 VSUBS 0.02141f
C1455 VN.n70 VSUBS 0.02141f
C1456 VN.n71 VSUBS 0.02141f
C1457 VN.n72 VSUBS 0.04235f
C1458 VN.n73 VSUBS 0.039903f
C1459 VN.n74 VSUBS 0.030053f
C1460 VN.n75 VSUBS 0.02141f
C1461 VN.n76 VSUBS 0.02141f
C1462 VN.n77 VSUBS 0.030053f
C1463 VN.n78 VSUBS 0.039903f
C1464 VN.n79 VSUBS 0.04235f
C1465 VN.n80 VSUBS 0.02141f
C1466 VN.n81 VSUBS 0.02141f
C1467 VN.n82 VSUBS 0.02141f
C1468 VN.n83 VSUBS 0.038437f
C1469 VN.n84 VSUBS 0.039903f
C1470 VN.n85 VSUBS 0.039509f
C1471 VN.n86 VSUBS 0.02141f
C1472 VN.n87 VSUBS 0.02141f
C1473 VN.n88 VSUBS 0.02141f
C1474 VN.n89 VSUBS 0.039903f
C1475 VN.n90 VSUBS 0.039903f
C1476 VN.n91 VSUBS 0.037528f
C1477 VN.n92 VSUBS 0.02141f
C1478 VN.n93 VSUBS 0.02141f
C1479 VN.n94 VSUBS 0.02141f
C1480 VN.n95 VSUBS 0.041503f
C1481 VN.n96 VSUBS 0.039903f
C1482 VN.n97 VSUBS 0.029265f
C1483 VN.n98 VSUBS 0.034556f
C1484 VN.n99 VSUBS 1.66986f
.ends

