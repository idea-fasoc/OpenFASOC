* NGSPICE file created from diff_pair_sample_1230.ext - technology: sky130A

.subckt diff_pair_sample_1230 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=0 ps=0 w=10.74 l=0.65
X1 VDD1.t7 VP.t0 VTAIL.t11 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=4.1886 ps=22.26 w=10.74 l=0.65
X2 VTAIL.t0 VN.t0 VDD2.t7 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
X3 VDD2.t6 VN.t1 VTAIL.t15 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=4.1886 ps=22.26 w=10.74 l=0.65
X4 VTAIL.t8 VP.t1 VDD1.t6 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=1.7721 ps=11.07 w=10.74 l=0.65
X5 VDD1.t5 VP.t2 VTAIL.t12 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=4.1886 ps=22.26 w=10.74 l=0.65
X6 VDD2.t5 VN.t2 VTAIL.t1 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=4.1886 ps=22.26 w=10.74 l=0.65
X7 VTAIL.t13 VP.t3 VDD1.t4 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
X8 VDD1.t3 VP.t4 VTAIL.t9 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
X9 VTAIL.t7 VP.t5 VDD1.t2 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=1.7721 ps=11.07 w=10.74 l=0.65
X10 B.t8 B.t6 B.t7 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=0 ps=0 w=10.74 l=0.65
X11 B.t5 B.t3 B.t4 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=0 ps=0 w=10.74 l=0.65
X12 VTAIL.t2 VN.t3 VDD2.t4 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=1.7721 ps=11.07 w=10.74 l=0.65
X13 VTAIL.t6 VN.t4 VDD2.t3 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=1.7721 ps=11.07 w=10.74 l=0.65
X14 VTAIL.t10 VP.t6 VDD1.t1 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
X15 VDD2.t2 VN.t5 VTAIL.t5 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
X16 B.t2 B.t0 B.t1 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=4.1886 pd=22.26 as=0 ps=0 w=10.74 l=0.65
X17 VTAIL.t3 VN.t6 VDD2.t1 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
X18 VDD2.t0 VN.t7 VTAIL.t4 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
X19 VDD1.t0 VP.t7 VTAIL.t14 w_n1950_n3116# sky130_fd_pr__pfet_01v8 ad=1.7721 pd=11.07 as=1.7721 ps=11.07 w=10.74 l=0.65
R0 B.n110 B.t3 601.833
R1 B.n102 B.t9 601.833
R2 B.n40 B.t6 601.833
R3 B.n32 B.t0 601.833
R4 B.n300 B.n83 585
R5 B.n299 B.n298 585
R6 B.n297 B.n84 585
R7 B.n296 B.n295 585
R8 B.n294 B.n85 585
R9 B.n293 B.n292 585
R10 B.n291 B.n86 585
R11 B.n290 B.n289 585
R12 B.n288 B.n87 585
R13 B.n287 B.n286 585
R14 B.n285 B.n88 585
R15 B.n284 B.n283 585
R16 B.n282 B.n89 585
R17 B.n281 B.n280 585
R18 B.n279 B.n90 585
R19 B.n278 B.n277 585
R20 B.n276 B.n91 585
R21 B.n275 B.n274 585
R22 B.n273 B.n92 585
R23 B.n272 B.n271 585
R24 B.n270 B.n93 585
R25 B.n269 B.n268 585
R26 B.n267 B.n94 585
R27 B.n266 B.n265 585
R28 B.n264 B.n95 585
R29 B.n263 B.n262 585
R30 B.n261 B.n96 585
R31 B.n260 B.n259 585
R32 B.n258 B.n97 585
R33 B.n257 B.n256 585
R34 B.n255 B.n98 585
R35 B.n254 B.n253 585
R36 B.n252 B.n99 585
R37 B.n251 B.n250 585
R38 B.n249 B.n100 585
R39 B.n248 B.n247 585
R40 B.n246 B.n101 585
R41 B.n245 B.n244 585
R42 B.n243 B.n242 585
R43 B.n241 B.n105 585
R44 B.n240 B.n239 585
R45 B.n238 B.n106 585
R46 B.n237 B.n236 585
R47 B.n235 B.n107 585
R48 B.n234 B.n233 585
R49 B.n232 B.n108 585
R50 B.n231 B.n230 585
R51 B.n228 B.n109 585
R52 B.n227 B.n226 585
R53 B.n225 B.n112 585
R54 B.n224 B.n223 585
R55 B.n222 B.n113 585
R56 B.n221 B.n220 585
R57 B.n219 B.n114 585
R58 B.n218 B.n217 585
R59 B.n216 B.n115 585
R60 B.n215 B.n214 585
R61 B.n213 B.n116 585
R62 B.n212 B.n211 585
R63 B.n210 B.n117 585
R64 B.n209 B.n208 585
R65 B.n207 B.n118 585
R66 B.n206 B.n205 585
R67 B.n204 B.n119 585
R68 B.n203 B.n202 585
R69 B.n201 B.n120 585
R70 B.n200 B.n199 585
R71 B.n198 B.n121 585
R72 B.n197 B.n196 585
R73 B.n195 B.n122 585
R74 B.n194 B.n193 585
R75 B.n192 B.n123 585
R76 B.n191 B.n190 585
R77 B.n189 B.n124 585
R78 B.n188 B.n187 585
R79 B.n186 B.n125 585
R80 B.n185 B.n184 585
R81 B.n183 B.n126 585
R82 B.n182 B.n181 585
R83 B.n180 B.n127 585
R84 B.n179 B.n178 585
R85 B.n177 B.n128 585
R86 B.n176 B.n175 585
R87 B.n174 B.n129 585
R88 B.n173 B.n172 585
R89 B.n302 B.n301 585
R90 B.n303 B.n82 585
R91 B.n305 B.n304 585
R92 B.n306 B.n81 585
R93 B.n308 B.n307 585
R94 B.n309 B.n80 585
R95 B.n311 B.n310 585
R96 B.n312 B.n79 585
R97 B.n314 B.n313 585
R98 B.n315 B.n78 585
R99 B.n317 B.n316 585
R100 B.n318 B.n77 585
R101 B.n320 B.n319 585
R102 B.n321 B.n76 585
R103 B.n323 B.n322 585
R104 B.n324 B.n75 585
R105 B.n326 B.n325 585
R106 B.n327 B.n74 585
R107 B.n329 B.n328 585
R108 B.n330 B.n73 585
R109 B.n332 B.n331 585
R110 B.n333 B.n72 585
R111 B.n335 B.n334 585
R112 B.n336 B.n71 585
R113 B.n338 B.n337 585
R114 B.n339 B.n70 585
R115 B.n341 B.n340 585
R116 B.n342 B.n69 585
R117 B.n344 B.n343 585
R118 B.n345 B.n68 585
R119 B.n347 B.n346 585
R120 B.n348 B.n67 585
R121 B.n350 B.n349 585
R122 B.n351 B.n66 585
R123 B.n353 B.n352 585
R124 B.n354 B.n65 585
R125 B.n356 B.n355 585
R126 B.n357 B.n64 585
R127 B.n359 B.n358 585
R128 B.n360 B.n63 585
R129 B.n362 B.n361 585
R130 B.n363 B.n62 585
R131 B.n365 B.n364 585
R132 B.n366 B.n61 585
R133 B.n368 B.n367 585
R134 B.n369 B.n60 585
R135 B.n498 B.n13 585
R136 B.n497 B.n496 585
R137 B.n495 B.n14 585
R138 B.n494 B.n493 585
R139 B.n492 B.n15 585
R140 B.n491 B.n490 585
R141 B.n489 B.n16 585
R142 B.n488 B.n487 585
R143 B.n486 B.n17 585
R144 B.n485 B.n484 585
R145 B.n483 B.n18 585
R146 B.n482 B.n481 585
R147 B.n480 B.n19 585
R148 B.n479 B.n478 585
R149 B.n477 B.n20 585
R150 B.n476 B.n475 585
R151 B.n474 B.n21 585
R152 B.n473 B.n472 585
R153 B.n471 B.n22 585
R154 B.n470 B.n469 585
R155 B.n468 B.n23 585
R156 B.n467 B.n466 585
R157 B.n465 B.n24 585
R158 B.n464 B.n463 585
R159 B.n462 B.n25 585
R160 B.n461 B.n460 585
R161 B.n459 B.n26 585
R162 B.n458 B.n457 585
R163 B.n456 B.n27 585
R164 B.n455 B.n454 585
R165 B.n453 B.n28 585
R166 B.n452 B.n451 585
R167 B.n450 B.n29 585
R168 B.n449 B.n448 585
R169 B.n447 B.n30 585
R170 B.n446 B.n445 585
R171 B.n444 B.n31 585
R172 B.n443 B.n442 585
R173 B.n441 B.n440 585
R174 B.n439 B.n35 585
R175 B.n438 B.n437 585
R176 B.n436 B.n36 585
R177 B.n435 B.n434 585
R178 B.n433 B.n37 585
R179 B.n432 B.n431 585
R180 B.n430 B.n38 585
R181 B.n429 B.n428 585
R182 B.n426 B.n39 585
R183 B.n425 B.n424 585
R184 B.n423 B.n42 585
R185 B.n422 B.n421 585
R186 B.n420 B.n43 585
R187 B.n419 B.n418 585
R188 B.n417 B.n44 585
R189 B.n416 B.n415 585
R190 B.n414 B.n45 585
R191 B.n413 B.n412 585
R192 B.n411 B.n46 585
R193 B.n410 B.n409 585
R194 B.n408 B.n47 585
R195 B.n407 B.n406 585
R196 B.n405 B.n48 585
R197 B.n404 B.n403 585
R198 B.n402 B.n49 585
R199 B.n401 B.n400 585
R200 B.n399 B.n50 585
R201 B.n398 B.n397 585
R202 B.n396 B.n51 585
R203 B.n395 B.n394 585
R204 B.n393 B.n52 585
R205 B.n392 B.n391 585
R206 B.n390 B.n53 585
R207 B.n389 B.n388 585
R208 B.n387 B.n54 585
R209 B.n386 B.n385 585
R210 B.n384 B.n55 585
R211 B.n383 B.n382 585
R212 B.n381 B.n56 585
R213 B.n380 B.n379 585
R214 B.n378 B.n57 585
R215 B.n377 B.n376 585
R216 B.n375 B.n58 585
R217 B.n374 B.n373 585
R218 B.n372 B.n59 585
R219 B.n371 B.n370 585
R220 B.n500 B.n499 585
R221 B.n501 B.n12 585
R222 B.n503 B.n502 585
R223 B.n504 B.n11 585
R224 B.n506 B.n505 585
R225 B.n507 B.n10 585
R226 B.n509 B.n508 585
R227 B.n510 B.n9 585
R228 B.n512 B.n511 585
R229 B.n513 B.n8 585
R230 B.n515 B.n514 585
R231 B.n516 B.n7 585
R232 B.n518 B.n517 585
R233 B.n519 B.n6 585
R234 B.n521 B.n520 585
R235 B.n522 B.n5 585
R236 B.n524 B.n523 585
R237 B.n525 B.n4 585
R238 B.n527 B.n526 585
R239 B.n528 B.n3 585
R240 B.n530 B.n529 585
R241 B.n531 B.n0 585
R242 B.n2 B.n1 585
R243 B.n141 B.n140 585
R244 B.n143 B.n142 585
R245 B.n144 B.n139 585
R246 B.n146 B.n145 585
R247 B.n147 B.n138 585
R248 B.n149 B.n148 585
R249 B.n150 B.n137 585
R250 B.n152 B.n151 585
R251 B.n153 B.n136 585
R252 B.n155 B.n154 585
R253 B.n156 B.n135 585
R254 B.n158 B.n157 585
R255 B.n159 B.n134 585
R256 B.n161 B.n160 585
R257 B.n162 B.n133 585
R258 B.n164 B.n163 585
R259 B.n165 B.n132 585
R260 B.n167 B.n166 585
R261 B.n168 B.n131 585
R262 B.n170 B.n169 585
R263 B.n171 B.n130 585
R264 B.n172 B.n171 535.745
R265 B.n302 B.n83 535.745
R266 B.n370 B.n369 535.745
R267 B.n500 B.n13 535.745
R268 B.n102 B.t10 371.986
R269 B.n40 B.t8 371.986
R270 B.n110 B.t4 371.986
R271 B.n32 B.t2 371.986
R272 B.n103 B.t11 352.981
R273 B.n41 B.t7 352.981
R274 B.n111 B.t5 352.979
R275 B.n33 B.t1 352.979
R276 B.n533 B.n532 256.663
R277 B.n532 B.n531 235.042
R278 B.n532 B.n2 235.042
R279 B.n172 B.n129 163.367
R280 B.n176 B.n129 163.367
R281 B.n177 B.n176 163.367
R282 B.n178 B.n177 163.367
R283 B.n178 B.n127 163.367
R284 B.n182 B.n127 163.367
R285 B.n183 B.n182 163.367
R286 B.n184 B.n183 163.367
R287 B.n184 B.n125 163.367
R288 B.n188 B.n125 163.367
R289 B.n189 B.n188 163.367
R290 B.n190 B.n189 163.367
R291 B.n190 B.n123 163.367
R292 B.n194 B.n123 163.367
R293 B.n195 B.n194 163.367
R294 B.n196 B.n195 163.367
R295 B.n196 B.n121 163.367
R296 B.n200 B.n121 163.367
R297 B.n201 B.n200 163.367
R298 B.n202 B.n201 163.367
R299 B.n202 B.n119 163.367
R300 B.n206 B.n119 163.367
R301 B.n207 B.n206 163.367
R302 B.n208 B.n207 163.367
R303 B.n208 B.n117 163.367
R304 B.n212 B.n117 163.367
R305 B.n213 B.n212 163.367
R306 B.n214 B.n213 163.367
R307 B.n214 B.n115 163.367
R308 B.n218 B.n115 163.367
R309 B.n219 B.n218 163.367
R310 B.n220 B.n219 163.367
R311 B.n220 B.n113 163.367
R312 B.n224 B.n113 163.367
R313 B.n225 B.n224 163.367
R314 B.n226 B.n225 163.367
R315 B.n226 B.n109 163.367
R316 B.n231 B.n109 163.367
R317 B.n232 B.n231 163.367
R318 B.n233 B.n232 163.367
R319 B.n233 B.n107 163.367
R320 B.n237 B.n107 163.367
R321 B.n238 B.n237 163.367
R322 B.n239 B.n238 163.367
R323 B.n239 B.n105 163.367
R324 B.n243 B.n105 163.367
R325 B.n244 B.n243 163.367
R326 B.n244 B.n101 163.367
R327 B.n248 B.n101 163.367
R328 B.n249 B.n248 163.367
R329 B.n250 B.n249 163.367
R330 B.n250 B.n99 163.367
R331 B.n254 B.n99 163.367
R332 B.n255 B.n254 163.367
R333 B.n256 B.n255 163.367
R334 B.n256 B.n97 163.367
R335 B.n260 B.n97 163.367
R336 B.n261 B.n260 163.367
R337 B.n262 B.n261 163.367
R338 B.n262 B.n95 163.367
R339 B.n266 B.n95 163.367
R340 B.n267 B.n266 163.367
R341 B.n268 B.n267 163.367
R342 B.n268 B.n93 163.367
R343 B.n272 B.n93 163.367
R344 B.n273 B.n272 163.367
R345 B.n274 B.n273 163.367
R346 B.n274 B.n91 163.367
R347 B.n278 B.n91 163.367
R348 B.n279 B.n278 163.367
R349 B.n280 B.n279 163.367
R350 B.n280 B.n89 163.367
R351 B.n284 B.n89 163.367
R352 B.n285 B.n284 163.367
R353 B.n286 B.n285 163.367
R354 B.n286 B.n87 163.367
R355 B.n290 B.n87 163.367
R356 B.n291 B.n290 163.367
R357 B.n292 B.n291 163.367
R358 B.n292 B.n85 163.367
R359 B.n296 B.n85 163.367
R360 B.n297 B.n296 163.367
R361 B.n298 B.n297 163.367
R362 B.n298 B.n83 163.367
R363 B.n369 B.n368 163.367
R364 B.n368 B.n61 163.367
R365 B.n364 B.n61 163.367
R366 B.n364 B.n363 163.367
R367 B.n363 B.n362 163.367
R368 B.n362 B.n63 163.367
R369 B.n358 B.n63 163.367
R370 B.n358 B.n357 163.367
R371 B.n357 B.n356 163.367
R372 B.n356 B.n65 163.367
R373 B.n352 B.n65 163.367
R374 B.n352 B.n351 163.367
R375 B.n351 B.n350 163.367
R376 B.n350 B.n67 163.367
R377 B.n346 B.n67 163.367
R378 B.n346 B.n345 163.367
R379 B.n345 B.n344 163.367
R380 B.n344 B.n69 163.367
R381 B.n340 B.n69 163.367
R382 B.n340 B.n339 163.367
R383 B.n339 B.n338 163.367
R384 B.n338 B.n71 163.367
R385 B.n334 B.n71 163.367
R386 B.n334 B.n333 163.367
R387 B.n333 B.n332 163.367
R388 B.n332 B.n73 163.367
R389 B.n328 B.n73 163.367
R390 B.n328 B.n327 163.367
R391 B.n327 B.n326 163.367
R392 B.n326 B.n75 163.367
R393 B.n322 B.n75 163.367
R394 B.n322 B.n321 163.367
R395 B.n321 B.n320 163.367
R396 B.n320 B.n77 163.367
R397 B.n316 B.n77 163.367
R398 B.n316 B.n315 163.367
R399 B.n315 B.n314 163.367
R400 B.n314 B.n79 163.367
R401 B.n310 B.n79 163.367
R402 B.n310 B.n309 163.367
R403 B.n309 B.n308 163.367
R404 B.n308 B.n81 163.367
R405 B.n304 B.n81 163.367
R406 B.n304 B.n303 163.367
R407 B.n303 B.n302 163.367
R408 B.n496 B.n13 163.367
R409 B.n496 B.n495 163.367
R410 B.n495 B.n494 163.367
R411 B.n494 B.n15 163.367
R412 B.n490 B.n15 163.367
R413 B.n490 B.n489 163.367
R414 B.n489 B.n488 163.367
R415 B.n488 B.n17 163.367
R416 B.n484 B.n17 163.367
R417 B.n484 B.n483 163.367
R418 B.n483 B.n482 163.367
R419 B.n482 B.n19 163.367
R420 B.n478 B.n19 163.367
R421 B.n478 B.n477 163.367
R422 B.n477 B.n476 163.367
R423 B.n476 B.n21 163.367
R424 B.n472 B.n21 163.367
R425 B.n472 B.n471 163.367
R426 B.n471 B.n470 163.367
R427 B.n470 B.n23 163.367
R428 B.n466 B.n23 163.367
R429 B.n466 B.n465 163.367
R430 B.n465 B.n464 163.367
R431 B.n464 B.n25 163.367
R432 B.n460 B.n25 163.367
R433 B.n460 B.n459 163.367
R434 B.n459 B.n458 163.367
R435 B.n458 B.n27 163.367
R436 B.n454 B.n27 163.367
R437 B.n454 B.n453 163.367
R438 B.n453 B.n452 163.367
R439 B.n452 B.n29 163.367
R440 B.n448 B.n29 163.367
R441 B.n448 B.n447 163.367
R442 B.n447 B.n446 163.367
R443 B.n446 B.n31 163.367
R444 B.n442 B.n31 163.367
R445 B.n442 B.n441 163.367
R446 B.n441 B.n35 163.367
R447 B.n437 B.n35 163.367
R448 B.n437 B.n436 163.367
R449 B.n436 B.n435 163.367
R450 B.n435 B.n37 163.367
R451 B.n431 B.n37 163.367
R452 B.n431 B.n430 163.367
R453 B.n430 B.n429 163.367
R454 B.n429 B.n39 163.367
R455 B.n424 B.n39 163.367
R456 B.n424 B.n423 163.367
R457 B.n423 B.n422 163.367
R458 B.n422 B.n43 163.367
R459 B.n418 B.n43 163.367
R460 B.n418 B.n417 163.367
R461 B.n417 B.n416 163.367
R462 B.n416 B.n45 163.367
R463 B.n412 B.n45 163.367
R464 B.n412 B.n411 163.367
R465 B.n411 B.n410 163.367
R466 B.n410 B.n47 163.367
R467 B.n406 B.n47 163.367
R468 B.n406 B.n405 163.367
R469 B.n405 B.n404 163.367
R470 B.n404 B.n49 163.367
R471 B.n400 B.n49 163.367
R472 B.n400 B.n399 163.367
R473 B.n399 B.n398 163.367
R474 B.n398 B.n51 163.367
R475 B.n394 B.n51 163.367
R476 B.n394 B.n393 163.367
R477 B.n393 B.n392 163.367
R478 B.n392 B.n53 163.367
R479 B.n388 B.n53 163.367
R480 B.n388 B.n387 163.367
R481 B.n387 B.n386 163.367
R482 B.n386 B.n55 163.367
R483 B.n382 B.n55 163.367
R484 B.n382 B.n381 163.367
R485 B.n381 B.n380 163.367
R486 B.n380 B.n57 163.367
R487 B.n376 B.n57 163.367
R488 B.n376 B.n375 163.367
R489 B.n375 B.n374 163.367
R490 B.n374 B.n59 163.367
R491 B.n370 B.n59 163.367
R492 B.n501 B.n500 163.367
R493 B.n502 B.n501 163.367
R494 B.n502 B.n11 163.367
R495 B.n506 B.n11 163.367
R496 B.n507 B.n506 163.367
R497 B.n508 B.n507 163.367
R498 B.n508 B.n9 163.367
R499 B.n512 B.n9 163.367
R500 B.n513 B.n512 163.367
R501 B.n514 B.n513 163.367
R502 B.n514 B.n7 163.367
R503 B.n518 B.n7 163.367
R504 B.n519 B.n518 163.367
R505 B.n520 B.n519 163.367
R506 B.n520 B.n5 163.367
R507 B.n524 B.n5 163.367
R508 B.n525 B.n524 163.367
R509 B.n526 B.n525 163.367
R510 B.n526 B.n3 163.367
R511 B.n530 B.n3 163.367
R512 B.n531 B.n530 163.367
R513 B.n141 B.n2 163.367
R514 B.n142 B.n141 163.367
R515 B.n142 B.n139 163.367
R516 B.n146 B.n139 163.367
R517 B.n147 B.n146 163.367
R518 B.n148 B.n147 163.367
R519 B.n148 B.n137 163.367
R520 B.n152 B.n137 163.367
R521 B.n153 B.n152 163.367
R522 B.n154 B.n153 163.367
R523 B.n154 B.n135 163.367
R524 B.n158 B.n135 163.367
R525 B.n159 B.n158 163.367
R526 B.n160 B.n159 163.367
R527 B.n160 B.n133 163.367
R528 B.n164 B.n133 163.367
R529 B.n165 B.n164 163.367
R530 B.n166 B.n165 163.367
R531 B.n166 B.n131 163.367
R532 B.n170 B.n131 163.367
R533 B.n171 B.n170 163.367
R534 B.n229 B.n111 59.5399
R535 B.n104 B.n103 59.5399
R536 B.n427 B.n41 59.5399
R537 B.n34 B.n33 59.5399
R538 B.n499 B.n498 34.8103
R539 B.n371 B.n60 34.8103
R540 B.n301 B.n300 34.8103
R541 B.n173 B.n130 34.8103
R542 B.n111 B.n110 19.0066
R543 B.n103 B.n102 19.0066
R544 B.n41 B.n40 19.0066
R545 B.n33 B.n32 19.0066
R546 B B.n533 18.0485
R547 B.n499 B.n12 10.6151
R548 B.n503 B.n12 10.6151
R549 B.n504 B.n503 10.6151
R550 B.n505 B.n504 10.6151
R551 B.n505 B.n10 10.6151
R552 B.n509 B.n10 10.6151
R553 B.n510 B.n509 10.6151
R554 B.n511 B.n510 10.6151
R555 B.n511 B.n8 10.6151
R556 B.n515 B.n8 10.6151
R557 B.n516 B.n515 10.6151
R558 B.n517 B.n516 10.6151
R559 B.n517 B.n6 10.6151
R560 B.n521 B.n6 10.6151
R561 B.n522 B.n521 10.6151
R562 B.n523 B.n522 10.6151
R563 B.n523 B.n4 10.6151
R564 B.n527 B.n4 10.6151
R565 B.n528 B.n527 10.6151
R566 B.n529 B.n528 10.6151
R567 B.n529 B.n0 10.6151
R568 B.n498 B.n497 10.6151
R569 B.n497 B.n14 10.6151
R570 B.n493 B.n14 10.6151
R571 B.n493 B.n492 10.6151
R572 B.n492 B.n491 10.6151
R573 B.n491 B.n16 10.6151
R574 B.n487 B.n16 10.6151
R575 B.n487 B.n486 10.6151
R576 B.n486 B.n485 10.6151
R577 B.n485 B.n18 10.6151
R578 B.n481 B.n18 10.6151
R579 B.n481 B.n480 10.6151
R580 B.n480 B.n479 10.6151
R581 B.n479 B.n20 10.6151
R582 B.n475 B.n20 10.6151
R583 B.n475 B.n474 10.6151
R584 B.n474 B.n473 10.6151
R585 B.n473 B.n22 10.6151
R586 B.n469 B.n22 10.6151
R587 B.n469 B.n468 10.6151
R588 B.n468 B.n467 10.6151
R589 B.n467 B.n24 10.6151
R590 B.n463 B.n24 10.6151
R591 B.n463 B.n462 10.6151
R592 B.n462 B.n461 10.6151
R593 B.n461 B.n26 10.6151
R594 B.n457 B.n26 10.6151
R595 B.n457 B.n456 10.6151
R596 B.n456 B.n455 10.6151
R597 B.n455 B.n28 10.6151
R598 B.n451 B.n28 10.6151
R599 B.n451 B.n450 10.6151
R600 B.n450 B.n449 10.6151
R601 B.n449 B.n30 10.6151
R602 B.n445 B.n30 10.6151
R603 B.n445 B.n444 10.6151
R604 B.n444 B.n443 10.6151
R605 B.n440 B.n439 10.6151
R606 B.n439 B.n438 10.6151
R607 B.n438 B.n36 10.6151
R608 B.n434 B.n36 10.6151
R609 B.n434 B.n433 10.6151
R610 B.n433 B.n432 10.6151
R611 B.n432 B.n38 10.6151
R612 B.n428 B.n38 10.6151
R613 B.n426 B.n425 10.6151
R614 B.n425 B.n42 10.6151
R615 B.n421 B.n42 10.6151
R616 B.n421 B.n420 10.6151
R617 B.n420 B.n419 10.6151
R618 B.n419 B.n44 10.6151
R619 B.n415 B.n44 10.6151
R620 B.n415 B.n414 10.6151
R621 B.n414 B.n413 10.6151
R622 B.n413 B.n46 10.6151
R623 B.n409 B.n46 10.6151
R624 B.n409 B.n408 10.6151
R625 B.n408 B.n407 10.6151
R626 B.n407 B.n48 10.6151
R627 B.n403 B.n48 10.6151
R628 B.n403 B.n402 10.6151
R629 B.n402 B.n401 10.6151
R630 B.n401 B.n50 10.6151
R631 B.n397 B.n50 10.6151
R632 B.n397 B.n396 10.6151
R633 B.n396 B.n395 10.6151
R634 B.n395 B.n52 10.6151
R635 B.n391 B.n52 10.6151
R636 B.n391 B.n390 10.6151
R637 B.n390 B.n389 10.6151
R638 B.n389 B.n54 10.6151
R639 B.n385 B.n54 10.6151
R640 B.n385 B.n384 10.6151
R641 B.n384 B.n383 10.6151
R642 B.n383 B.n56 10.6151
R643 B.n379 B.n56 10.6151
R644 B.n379 B.n378 10.6151
R645 B.n378 B.n377 10.6151
R646 B.n377 B.n58 10.6151
R647 B.n373 B.n58 10.6151
R648 B.n373 B.n372 10.6151
R649 B.n372 B.n371 10.6151
R650 B.n367 B.n60 10.6151
R651 B.n367 B.n366 10.6151
R652 B.n366 B.n365 10.6151
R653 B.n365 B.n62 10.6151
R654 B.n361 B.n62 10.6151
R655 B.n361 B.n360 10.6151
R656 B.n360 B.n359 10.6151
R657 B.n359 B.n64 10.6151
R658 B.n355 B.n64 10.6151
R659 B.n355 B.n354 10.6151
R660 B.n354 B.n353 10.6151
R661 B.n353 B.n66 10.6151
R662 B.n349 B.n66 10.6151
R663 B.n349 B.n348 10.6151
R664 B.n348 B.n347 10.6151
R665 B.n347 B.n68 10.6151
R666 B.n343 B.n68 10.6151
R667 B.n343 B.n342 10.6151
R668 B.n342 B.n341 10.6151
R669 B.n341 B.n70 10.6151
R670 B.n337 B.n70 10.6151
R671 B.n337 B.n336 10.6151
R672 B.n336 B.n335 10.6151
R673 B.n335 B.n72 10.6151
R674 B.n331 B.n72 10.6151
R675 B.n331 B.n330 10.6151
R676 B.n330 B.n329 10.6151
R677 B.n329 B.n74 10.6151
R678 B.n325 B.n74 10.6151
R679 B.n325 B.n324 10.6151
R680 B.n324 B.n323 10.6151
R681 B.n323 B.n76 10.6151
R682 B.n319 B.n76 10.6151
R683 B.n319 B.n318 10.6151
R684 B.n318 B.n317 10.6151
R685 B.n317 B.n78 10.6151
R686 B.n313 B.n78 10.6151
R687 B.n313 B.n312 10.6151
R688 B.n312 B.n311 10.6151
R689 B.n311 B.n80 10.6151
R690 B.n307 B.n80 10.6151
R691 B.n307 B.n306 10.6151
R692 B.n306 B.n305 10.6151
R693 B.n305 B.n82 10.6151
R694 B.n301 B.n82 10.6151
R695 B.n140 B.n1 10.6151
R696 B.n143 B.n140 10.6151
R697 B.n144 B.n143 10.6151
R698 B.n145 B.n144 10.6151
R699 B.n145 B.n138 10.6151
R700 B.n149 B.n138 10.6151
R701 B.n150 B.n149 10.6151
R702 B.n151 B.n150 10.6151
R703 B.n151 B.n136 10.6151
R704 B.n155 B.n136 10.6151
R705 B.n156 B.n155 10.6151
R706 B.n157 B.n156 10.6151
R707 B.n157 B.n134 10.6151
R708 B.n161 B.n134 10.6151
R709 B.n162 B.n161 10.6151
R710 B.n163 B.n162 10.6151
R711 B.n163 B.n132 10.6151
R712 B.n167 B.n132 10.6151
R713 B.n168 B.n167 10.6151
R714 B.n169 B.n168 10.6151
R715 B.n169 B.n130 10.6151
R716 B.n174 B.n173 10.6151
R717 B.n175 B.n174 10.6151
R718 B.n175 B.n128 10.6151
R719 B.n179 B.n128 10.6151
R720 B.n180 B.n179 10.6151
R721 B.n181 B.n180 10.6151
R722 B.n181 B.n126 10.6151
R723 B.n185 B.n126 10.6151
R724 B.n186 B.n185 10.6151
R725 B.n187 B.n186 10.6151
R726 B.n187 B.n124 10.6151
R727 B.n191 B.n124 10.6151
R728 B.n192 B.n191 10.6151
R729 B.n193 B.n192 10.6151
R730 B.n193 B.n122 10.6151
R731 B.n197 B.n122 10.6151
R732 B.n198 B.n197 10.6151
R733 B.n199 B.n198 10.6151
R734 B.n199 B.n120 10.6151
R735 B.n203 B.n120 10.6151
R736 B.n204 B.n203 10.6151
R737 B.n205 B.n204 10.6151
R738 B.n205 B.n118 10.6151
R739 B.n209 B.n118 10.6151
R740 B.n210 B.n209 10.6151
R741 B.n211 B.n210 10.6151
R742 B.n211 B.n116 10.6151
R743 B.n215 B.n116 10.6151
R744 B.n216 B.n215 10.6151
R745 B.n217 B.n216 10.6151
R746 B.n217 B.n114 10.6151
R747 B.n221 B.n114 10.6151
R748 B.n222 B.n221 10.6151
R749 B.n223 B.n222 10.6151
R750 B.n223 B.n112 10.6151
R751 B.n227 B.n112 10.6151
R752 B.n228 B.n227 10.6151
R753 B.n230 B.n108 10.6151
R754 B.n234 B.n108 10.6151
R755 B.n235 B.n234 10.6151
R756 B.n236 B.n235 10.6151
R757 B.n236 B.n106 10.6151
R758 B.n240 B.n106 10.6151
R759 B.n241 B.n240 10.6151
R760 B.n242 B.n241 10.6151
R761 B.n246 B.n245 10.6151
R762 B.n247 B.n246 10.6151
R763 B.n247 B.n100 10.6151
R764 B.n251 B.n100 10.6151
R765 B.n252 B.n251 10.6151
R766 B.n253 B.n252 10.6151
R767 B.n253 B.n98 10.6151
R768 B.n257 B.n98 10.6151
R769 B.n258 B.n257 10.6151
R770 B.n259 B.n258 10.6151
R771 B.n259 B.n96 10.6151
R772 B.n263 B.n96 10.6151
R773 B.n264 B.n263 10.6151
R774 B.n265 B.n264 10.6151
R775 B.n265 B.n94 10.6151
R776 B.n269 B.n94 10.6151
R777 B.n270 B.n269 10.6151
R778 B.n271 B.n270 10.6151
R779 B.n271 B.n92 10.6151
R780 B.n275 B.n92 10.6151
R781 B.n276 B.n275 10.6151
R782 B.n277 B.n276 10.6151
R783 B.n277 B.n90 10.6151
R784 B.n281 B.n90 10.6151
R785 B.n282 B.n281 10.6151
R786 B.n283 B.n282 10.6151
R787 B.n283 B.n88 10.6151
R788 B.n287 B.n88 10.6151
R789 B.n288 B.n287 10.6151
R790 B.n289 B.n288 10.6151
R791 B.n289 B.n86 10.6151
R792 B.n293 B.n86 10.6151
R793 B.n294 B.n293 10.6151
R794 B.n295 B.n294 10.6151
R795 B.n295 B.n84 10.6151
R796 B.n299 B.n84 10.6151
R797 B.n300 B.n299 10.6151
R798 B.n533 B.n0 8.11757
R799 B.n533 B.n1 8.11757
R800 B.n440 B.n34 6.5566
R801 B.n428 B.n427 6.5566
R802 B.n230 B.n229 6.5566
R803 B.n242 B.n104 6.5566
R804 B.n443 B.n34 4.05904
R805 B.n427 B.n426 4.05904
R806 B.n229 B.n228 4.05904
R807 B.n245 B.n104 4.05904
R808 VP.n3 VP.t1 486.204
R809 VP.n1 VP.t5 459.384
R810 VP.n10 VP.t4 459.384
R811 VP.n11 VP.t3 459.384
R812 VP.n12 VP.t0 459.384
R813 VP.n6 VP.t2 459.384
R814 VP.n5 VP.t6 459.384
R815 VP.n4 VP.t7 459.384
R816 VP.n13 VP.n12 161.3
R817 VP.n7 VP.n6 161.3
R818 VP.n8 VP.n1 161.3
R819 VP.n5 VP.n2 80.6037
R820 VP.n11 VP.n0 80.6037
R821 VP.n10 VP.n9 80.6037
R822 VP.n10 VP.n1 48.2005
R823 VP.n11 VP.n10 48.2005
R824 VP.n12 VP.n11 48.2005
R825 VP.n6 VP.n5 48.2005
R826 VP.n5 VP.n4 48.2005
R827 VP.n3 VP.n2 45.2318
R828 VP.n8 VP.n7 40.9247
R829 VP.n4 VP.n3 13.3799
R830 VP.n9 VP.n0 0.380177
R831 VP.n7 VP.n2 0.285035
R832 VP.n9 VP.n8 0.285035
R833 VP.n13 VP.n0 0.285035
R834 VP VP.n13 0.0516364
R835 VTAIL.n466 VTAIL.n414 756.745
R836 VTAIL.n54 VTAIL.n2 756.745
R837 VTAIL.n112 VTAIL.n60 756.745
R838 VTAIL.n172 VTAIL.n120 756.745
R839 VTAIL.n408 VTAIL.n356 756.745
R840 VTAIL.n348 VTAIL.n296 756.745
R841 VTAIL.n290 VTAIL.n238 756.745
R842 VTAIL.n230 VTAIL.n178 756.745
R843 VTAIL.n433 VTAIL.n432 585
R844 VTAIL.n430 VTAIL.n429 585
R845 VTAIL.n439 VTAIL.n438 585
R846 VTAIL.n441 VTAIL.n440 585
R847 VTAIL.n426 VTAIL.n425 585
R848 VTAIL.n447 VTAIL.n446 585
R849 VTAIL.n450 VTAIL.n449 585
R850 VTAIL.n448 VTAIL.n422 585
R851 VTAIL.n455 VTAIL.n421 585
R852 VTAIL.n457 VTAIL.n456 585
R853 VTAIL.n459 VTAIL.n458 585
R854 VTAIL.n418 VTAIL.n417 585
R855 VTAIL.n465 VTAIL.n464 585
R856 VTAIL.n467 VTAIL.n466 585
R857 VTAIL.n21 VTAIL.n20 585
R858 VTAIL.n18 VTAIL.n17 585
R859 VTAIL.n27 VTAIL.n26 585
R860 VTAIL.n29 VTAIL.n28 585
R861 VTAIL.n14 VTAIL.n13 585
R862 VTAIL.n35 VTAIL.n34 585
R863 VTAIL.n38 VTAIL.n37 585
R864 VTAIL.n36 VTAIL.n10 585
R865 VTAIL.n43 VTAIL.n9 585
R866 VTAIL.n45 VTAIL.n44 585
R867 VTAIL.n47 VTAIL.n46 585
R868 VTAIL.n6 VTAIL.n5 585
R869 VTAIL.n53 VTAIL.n52 585
R870 VTAIL.n55 VTAIL.n54 585
R871 VTAIL.n79 VTAIL.n78 585
R872 VTAIL.n76 VTAIL.n75 585
R873 VTAIL.n85 VTAIL.n84 585
R874 VTAIL.n87 VTAIL.n86 585
R875 VTAIL.n72 VTAIL.n71 585
R876 VTAIL.n93 VTAIL.n92 585
R877 VTAIL.n96 VTAIL.n95 585
R878 VTAIL.n94 VTAIL.n68 585
R879 VTAIL.n101 VTAIL.n67 585
R880 VTAIL.n103 VTAIL.n102 585
R881 VTAIL.n105 VTAIL.n104 585
R882 VTAIL.n64 VTAIL.n63 585
R883 VTAIL.n111 VTAIL.n110 585
R884 VTAIL.n113 VTAIL.n112 585
R885 VTAIL.n139 VTAIL.n138 585
R886 VTAIL.n136 VTAIL.n135 585
R887 VTAIL.n145 VTAIL.n144 585
R888 VTAIL.n147 VTAIL.n146 585
R889 VTAIL.n132 VTAIL.n131 585
R890 VTAIL.n153 VTAIL.n152 585
R891 VTAIL.n156 VTAIL.n155 585
R892 VTAIL.n154 VTAIL.n128 585
R893 VTAIL.n161 VTAIL.n127 585
R894 VTAIL.n163 VTAIL.n162 585
R895 VTAIL.n165 VTAIL.n164 585
R896 VTAIL.n124 VTAIL.n123 585
R897 VTAIL.n171 VTAIL.n170 585
R898 VTAIL.n173 VTAIL.n172 585
R899 VTAIL.n409 VTAIL.n408 585
R900 VTAIL.n407 VTAIL.n406 585
R901 VTAIL.n360 VTAIL.n359 585
R902 VTAIL.n401 VTAIL.n400 585
R903 VTAIL.n399 VTAIL.n398 585
R904 VTAIL.n397 VTAIL.n363 585
R905 VTAIL.n367 VTAIL.n364 585
R906 VTAIL.n392 VTAIL.n391 585
R907 VTAIL.n390 VTAIL.n389 585
R908 VTAIL.n369 VTAIL.n368 585
R909 VTAIL.n384 VTAIL.n383 585
R910 VTAIL.n382 VTAIL.n381 585
R911 VTAIL.n373 VTAIL.n372 585
R912 VTAIL.n376 VTAIL.n375 585
R913 VTAIL.n349 VTAIL.n348 585
R914 VTAIL.n347 VTAIL.n346 585
R915 VTAIL.n300 VTAIL.n299 585
R916 VTAIL.n341 VTAIL.n340 585
R917 VTAIL.n339 VTAIL.n338 585
R918 VTAIL.n337 VTAIL.n303 585
R919 VTAIL.n307 VTAIL.n304 585
R920 VTAIL.n332 VTAIL.n331 585
R921 VTAIL.n330 VTAIL.n329 585
R922 VTAIL.n309 VTAIL.n308 585
R923 VTAIL.n324 VTAIL.n323 585
R924 VTAIL.n322 VTAIL.n321 585
R925 VTAIL.n313 VTAIL.n312 585
R926 VTAIL.n316 VTAIL.n315 585
R927 VTAIL.n291 VTAIL.n290 585
R928 VTAIL.n289 VTAIL.n288 585
R929 VTAIL.n242 VTAIL.n241 585
R930 VTAIL.n283 VTAIL.n282 585
R931 VTAIL.n281 VTAIL.n280 585
R932 VTAIL.n279 VTAIL.n245 585
R933 VTAIL.n249 VTAIL.n246 585
R934 VTAIL.n274 VTAIL.n273 585
R935 VTAIL.n272 VTAIL.n271 585
R936 VTAIL.n251 VTAIL.n250 585
R937 VTAIL.n266 VTAIL.n265 585
R938 VTAIL.n264 VTAIL.n263 585
R939 VTAIL.n255 VTAIL.n254 585
R940 VTAIL.n258 VTAIL.n257 585
R941 VTAIL.n231 VTAIL.n230 585
R942 VTAIL.n229 VTAIL.n228 585
R943 VTAIL.n182 VTAIL.n181 585
R944 VTAIL.n223 VTAIL.n222 585
R945 VTAIL.n221 VTAIL.n220 585
R946 VTAIL.n219 VTAIL.n185 585
R947 VTAIL.n189 VTAIL.n186 585
R948 VTAIL.n214 VTAIL.n213 585
R949 VTAIL.n212 VTAIL.n211 585
R950 VTAIL.n191 VTAIL.n190 585
R951 VTAIL.n206 VTAIL.n205 585
R952 VTAIL.n204 VTAIL.n203 585
R953 VTAIL.n195 VTAIL.n194 585
R954 VTAIL.n198 VTAIL.n197 585
R955 VTAIL.t12 VTAIL.n374 329.038
R956 VTAIL.t8 VTAIL.n314 329.038
R957 VTAIL.t1 VTAIL.n256 329.038
R958 VTAIL.t2 VTAIL.n196 329.038
R959 VTAIL.t15 VTAIL.n431 329.038
R960 VTAIL.t6 VTAIL.n19 329.038
R961 VTAIL.t11 VTAIL.n77 329.038
R962 VTAIL.t7 VTAIL.n137 329.038
R963 VTAIL.n432 VTAIL.n429 171.744
R964 VTAIL.n439 VTAIL.n429 171.744
R965 VTAIL.n440 VTAIL.n439 171.744
R966 VTAIL.n440 VTAIL.n425 171.744
R967 VTAIL.n447 VTAIL.n425 171.744
R968 VTAIL.n449 VTAIL.n447 171.744
R969 VTAIL.n449 VTAIL.n448 171.744
R970 VTAIL.n448 VTAIL.n421 171.744
R971 VTAIL.n457 VTAIL.n421 171.744
R972 VTAIL.n458 VTAIL.n457 171.744
R973 VTAIL.n458 VTAIL.n417 171.744
R974 VTAIL.n465 VTAIL.n417 171.744
R975 VTAIL.n466 VTAIL.n465 171.744
R976 VTAIL.n20 VTAIL.n17 171.744
R977 VTAIL.n27 VTAIL.n17 171.744
R978 VTAIL.n28 VTAIL.n27 171.744
R979 VTAIL.n28 VTAIL.n13 171.744
R980 VTAIL.n35 VTAIL.n13 171.744
R981 VTAIL.n37 VTAIL.n35 171.744
R982 VTAIL.n37 VTAIL.n36 171.744
R983 VTAIL.n36 VTAIL.n9 171.744
R984 VTAIL.n45 VTAIL.n9 171.744
R985 VTAIL.n46 VTAIL.n45 171.744
R986 VTAIL.n46 VTAIL.n5 171.744
R987 VTAIL.n53 VTAIL.n5 171.744
R988 VTAIL.n54 VTAIL.n53 171.744
R989 VTAIL.n78 VTAIL.n75 171.744
R990 VTAIL.n85 VTAIL.n75 171.744
R991 VTAIL.n86 VTAIL.n85 171.744
R992 VTAIL.n86 VTAIL.n71 171.744
R993 VTAIL.n93 VTAIL.n71 171.744
R994 VTAIL.n95 VTAIL.n93 171.744
R995 VTAIL.n95 VTAIL.n94 171.744
R996 VTAIL.n94 VTAIL.n67 171.744
R997 VTAIL.n103 VTAIL.n67 171.744
R998 VTAIL.n104 VTAIL.n103 171.744
R999 VTAIL.n104 VTAIL.n63 171.744
R1000 VTAIL.n111 VTAIL.n63 171.744
R1001 VTAIL.n112 VTAIL.n111 171.744
R1002 VTAIL.n138 VTAIL.n135 171.744
R1003 VTAIL.n145 VTAIL.n135 171.744
R1004 VTAIL.n146 VTAIL.n145 171.744
R1005 VTAIL.n146 VTAIL.n131 171.744
R1006 VTAIL.n153 VTAIL.n131 171.744
R1007 VTAIL.n155 VTAIL.n153 171.744
R1008 VTAIL.n155 VTAIL.n154 171.744
R1009 VTAIL.n154 VTAIL.n127 171.744
R1010 VTAIL.n163 VTAIL.n127 171.744
R1011 VTAIL.n164 VTAIL.n163 171.744
R1012 VTAIL.n164 VTAIL.n123 171.744
R1013 VTAIL.n171 VTAIL.n123 171.744
R1014 VTAIL.n172 VTAIL.n171 171.744
R1015 VTAIL.n408 VTAIL.n407 171.744
R1016 VTAIL.n407 VTAIL.n359 171.744
R1017 VTAIL.n400 VTAIL.n359 171.744
R1018 VTAIL.n400 VTAIL.n399 171.744
R1019 VTAIL.n399 VTAIL.n363 171.744
R1020 VTAIL.n367 VTAIL.n363 171.744
R1021 VTAIL.n391 VTAIL.n367 171.744
R1022 VTAIL.n391 VTAIL.n390 171.744
R1023 VTAIL.n390 VTAIL.n368 171.744
R1024 VTAIL.n383 VTAIL.n368 171.744
R1025 VTAIL.n383 VTAIL.n382 171.744
R1026 VTAIL.n382 VTAIL.n372 171.744
R1027 VTAIL.n375 VTAIL.n372 171.744
R1028 VTAIL.n348 VTAIL.n347 171.744
R1029 VTAIL.n347 VTAIL.n299 171.744
R1030 VTAIL.n340 VTAIL.n299 171.744
R1031 VTAIL.n340 VTAIL.n339 171.744
R1032 VTAIL.n339 VTAIL.n303 171.744
R1033 VTAIL.n307 VTAIL.n303 171.744
R1034 VTAIL.n331 VTAIL.n307 171.744
R1035 VTAIL.n331 VTAIL.n330 171.744
R1036 VTAIL.n330 VTAIL.n308 171.744
R1037 VTAIL.n323 VTAIL.n308 171.744
R1038 VTAIL.n323 VTAIL.n322 171.744
R1039 VTAIL.n322 VTAIL.n312 171.744
R1040 VTAIL.n315 VTAIL.n312 171.744
R1041 VTAIL.n290 VTAIL.n289 171.744
R1042 VTAIL.n289 VTAIL.n241 171.744
R1043 VTAIL.n282 VTAIL.n241 171.744
R1044 VTAIL.n282 VTAIL.n281 171.744
R1045 VTAIL.n281 VTAIL.n245 171.744
R1046 VTAIL.n249 VTAIL.n245 171.744
R1047 VTAIL.n273 VTAIL.n249 171.744
R1048 VTAIL.n273 VTAIL.n272 171.744
R1049 VTAIL.n272 VTAIL.n250 171.744
R1050 VTAIL.n265 VTAIL.n250 171.744
R1051 VTAIL.n265 VTAIL.n264 171.744
R1052 VTAIL.n264 VTAIL.n254 171.744
R1053 VTAIL.n257 VTAIL.n254 171.744
R1054 VTAIL.n230 VTAIL.n229 171.744
R1055 VTAIL.n229 VTAIL.n181 171.744
R1056 VTAIL.n222 VTAIL.n181 171.744
R1057 VTAIL.n222 VTAIL.n221 171.744
R1058 VTAIL.n221 VTAIL.n185 171.744
R1059 VTAIL.n189 VTAIL.n185 171.744
R1060 VTAIL.n213 VTAIL.n189 171.744
R1061 VTAIL.n213 VTAIL.n212 171.744
R1062 VTAIL.n212 VTAIL.n190 171.744
R1063 VTAIL.n205 VTAIL.n190 171.744
R1064 VTAIL.n205 VTAIL.n204 171.744
R1065 VTAIL.n204 VTAIL.n194 171.744
R1066 VTAIL.n197 VTAIL.n194 171.744
R1067 VTAIL.n432 VTAIL.t15 85.8723
R1068 VTAIL.n20 VTAIL.t6 85.8723
R1069 VTAIL.n78 VTAIL.t11 85.8723
R1070 VTAIL.n138 VTAIL.t7 85.8723
R1071 VTAIL.n375 VTAIL.t12 85.8723
R1072 VTAIL.n315 VTAIL.t8 85.8723
R1073 VTAIL.n257 VTAIL.t1 85.8723
R1074 VTAIL.n197 VTAIL.t2 85.8723
R1075 VTAIL.n355 VTAIL.n354 60.351
R1076 VTAIL.n237 VTAIL.n236 60.351
R1077 VTAIL.n1 VTAIL.n0 60.3508
R1078 VTAIL.n119 VTAIL.n118 60.3508
R1079 VTAIL.n471 VTAIL.n470 33.349
R1080 VTAIL.n59 VTAIL.n58 33.349
R1081 VTAIL.n117 VTAIL.n116 33.349
R1082 VTAIL.n177 VTAIL.n176 33.349
R1083 VTAIL.n413 VTAIL.n412 33.349
R1084 VTAIL.n353 VTAIL.n352 33.349
R1085 VTAIL.n295 VTAIL.n294 33.349
R1086 VTAIL.n235 VTAIL.n234 33.349
R1087 VTAIL.n471 VTAIL.n413 22.4703
R1088 VTAIL.n235 VTAIL.n177 22.4703
R1089 VTAIL.n456 VTAIL.n455 13.1884
R1090 VTAIL.n44 VTAIL.n43 13.1884
R1091 VTAIL.n102 VTAIL.n101 13.1884
R1092 VTAIL.n162 VTAIL.n161 13.1884
R1093 VTAIL.n398 VTAIL.n397 13.1884
R1094 VTAIL.n338 VTAIL.n337 13.1884
R1095 VTAIL.n280 VTAIL.n279 13.1884
R1096 VTAIL.n220 VTAIL.n219 13.1884
R1097 VTAIL.n454 VTAIL.n422 12.8005
R1098 VTAIL.n459 VTAIL.n420 12.8005
R1099 VTAIL.n42 VTAIL.n10 12.8005
R1100 VTAIL.n47 VTAIL.n8 12.8005
R1101 VTAIL.n100 VTAIL.n68 12.8005
R1102 VTAIL.n105 VTAIL.n66 12.8005
R1103 VTAIL.n160 VTAIL.n128 12.8005
R1104 VTAIL.n165 VTAIL.n126 12.8005
R1105 VTAIL.n401 VTAIL.n362 12.8005
R1106 VTAIL.n396 VTAIL.n364 12.8005
R1107 VTAIL.n341 VTAIL.n302 12.8005
R1108 VTAIL.n336 VTAIL.n304 12.8005
R1109 VTAIL.n283 VTAIL.n244 12.8005
R1110 VTAIL.n278 VTAIL.n246 12.8005
R1111 VTAIL.n223 VTAIL.n184 12.8005
R1112 VTAIL.n218 VTAIL.n186 12.8005
R1113 VTAIL.n451 VTAIL.n450 12.0247
R1114 VTAIL.n460 VTAIL.n418 12.0247
R1115 VTAIL.n39 VTAIL.n38 12.0247
R1116 VTAIL.n48 VTAIL.n6 12.0247
R1117 VTAIL.n97 VTAIL.n96 12.0247
R1118 VTAIL.n106 VTAIL.n64 12.0247
R1119 VTAIL.n157 VTAIL.n156 12.0247
R1120 VTAIL.n166 VTAIL.n124 12.0247
R1121 VTAIL.n402 VTAIL.n360 12.0247
R1122 VTAIL.n393 VTAIL.n392 12.0247
R1123 VTAIL.n342 VTAIL.n300 12.0247
R1124 VTAIL.n333 VTAIL.n332 12.0247
R1125 VTAIL.n284 VTAIL.n242 12.0247
R1126 VTAIL.n275 VTAIL.n274 12.0247
R1127 VTAIL.n224 VTAIL.n182 12.0247
R1128 VTAIL.n215 VTAIL.n214 12.0247
R1129 VTAIL.n446 VTAIL.n424 11.249
R1130 VTAIL.n464 VTAIL.n463 11.249
R1131 VTAIL.n34 VTAIL.n12 11.249
R1132 VTAIL.n52 VTAIL.n51 11.249
R1133 VTAIL.n92 VTAIL.n70 11.249
R1134 VTAIL.n110 VTAIL.n109 11.249
R1135 VTAIL.n152 VTAIL.n130 11.249
R1136 VTAIL.n170 VTAIL.n169 11.249
R1137 VTAIL.n406 VTAIL.n405 11.249
R1138 VTAIL.n389 VTAIL.n366 11.249
R1139 VTAIL.n346 VTAIL.n345 11.249
R1140 VTAIL.n329 VTAIL.n306 11.249
R1141 VTAIL.n288 VTAIL.n287 11.249
R1142 VTAIL.n271 VTAIL.n248 11.249
R1143 VTAIL.n228 VTAIL.n227 11.249
R1144 VTAIL.n211 VTAIL.n188 11.249
R1145 VTAIL.n433 VTAIL.n431 10.7239
R1146 VTAIL.n21 VTAIL.n19 10.7239
R1147 VTAIL.n79 VTAIL.n77 10.7239
R1148 VTAIL.n139 VTAIL.n137 10.7239
R1149 VTAIL.n376 VTAIL.n374 10.7239
R1150 VTAIL.n316 VTAIL.n314 10.7239
R1151 VTAIL.n258 VTAIL.n256 10.7239
R1152 VTAIL.n198 VTAIL.n196 10.7239
R1153 VTAIL.n445 VTAIL.n426 10.4732
R1154 VTAIL.n467 VTAIL.n416 10.4732
R1155 VTAIL.n33 VTAIL.n14 10.4732
R1156 VTAIL.n55 VTAIL.n4 10.4732
R1157 VTAIL.n91 VTAIL.n72 10.4732
R1158 VTAIL.n113 VTAIL.n62 10.4732
R1159 VTAIL.n151 VTAIL.n132 10.4732
R1160 VTAIL.n173 VTAIL.n122 10.4732
R1161 VTAIL.n409 VTAIL.n358 10.4732
R1162 VTAIL.n388 VTAIL.n369 10.4732
R1163 VTAIL.n349 VTAIL.n298 10.4732
R1164 VTAIL.n328 VTAIL.n309 10.4732
R1165 VTAIL.n291 VTAIL.n240 10.4732
R1166 VTAIL.n270 VTAIL.n251 10.4732
R1167 VTAIL.n231 VTAIL.n180 10.4732
R1168 VTAIL.n210 VTAIL.n191 10.4732
R1169 VTAIL.n442 VTAIL.n441 9.69747
R1170 VTAIL.n468 VTAIL.n414 9.69747
R1171 VTAIL.n30 VTAIL.n29 9.69747
R1172 VTAIL.n56 VTAIL.n2 9.69747
R1173 VTAIL.n88 VTAIL.n87 9.69747
R1174 VTAIL.n114 VTAIL.n60 9.69747
R1175 VTAIL.n148 VTAIL.n147 9.69747
R1176 VTAIL.n174 VTAIL.n120 9.69747
R1177 VTAIL.n410 VTAIL.n356 9.69747
R1178 VTAIL.n385 VTAIL.n384 9.69747
R1179 VTAIL.n350 VTAIL.n296 9.69747
R1180 VTAIL.n325 VTAIL.n324 9.69747
R1181 VTAIL.n292 VTAIL.n238 9.69747
R1182 VTAIL.n267 VTAIL.n266 9.69747
R1183 VTAIL.n232 VTAIL.n178 9.69747
R1184 VTAIL.n207 VTAIL.n206 9.69747
R1185 VTAIL.n470 VTAIL.n469 9.45567
R1186 VTAIL.n58 VTAIL.n57 9.45567
R1187 VTAIL.n116 VTAIL.n115 9.45567
R1188 VTAIL.n176 VTAIL.n175 9.45567
R1189 VTAIL.n412 VTAIL.n411 9.45567
R1190 VTAIL.n352 VTAIL.n351 9.45567
R1191 VTAIL.n294 VTAIL.n293 9.45567
R1192 VTAIL.n234 VTAIL.n233 9.45567
R1193 VTAIL.n469 VTAIL.n468 9.3005
R1194 VTAIL.n416 VTAIL.n415 9.3005
R1195 VTAIL.n463 VTAIL.n462 9.3005
R1196 VTAIL.n461 VTAIL.n460 9.3005
R1197 VTAIL.n420 VTAIL.n419 9.3005
R1198 VTAIL.n435 VTAIL.n434 9.3005
R1199 VTAIL.n437 VTAIL.n436 9.3005
R1200 VTAIL.n428 VTAIL.n427 9.3005
R1201 VTAIL.n443 VTAIL.n442 9.3005
R1202 VTAIL.n445 VTAIL.n444 9.3005
R1203 VTAIL.n424 VTAIL.n423 9.3005
R1204 VTAIL.n452 VTAIL.n451 9.3005
R1205 VTAIL.n454 VTAIL.n453 9.3005
R1206 VTAIL.n57 VTAIL.n56 9.3005
R1207 VTAIL.n4 VTAIL.n3 9.3005
R1208 VTAIL.n51 VTAIL.n50 9.3005
R1209 VTAIL.n49 VTAIL.n48 9.3005
R1210 VTAIL.n8 VTAIL.n7 9.3005
R1211 VTAIL.n23 VTAIL.n22 9.3005
R1212 VTAIL.n25 VTAIL.n24 9.3005
R1213 VTAIL.n16 VTAIL.n15 9.3005
R1214 VTAIL.n31 VTAIL.n30 9.3005
R1215 VTAIL.n33 VTAIL.n32 9.3005
R1216 VTAIL.n12 VTAIL.n11 9.3005
R1217 VTAIL.n40 VTAIL.n39 9.3005
R1218 VTAIL.n42 VTAIL.n41 9.3005
R1219 VTAIL.n115 VTAIL.n114 9.3005
R1220 VTAIL.n62 VTAIL.n61 9.3005
R1221 VTAIL.n109 VTAIL.n108 9.3005
R1222 VTAIL.n107 VTAIL.n106 9.3005
R1223 VTAIL.n66 VTAIL.n65 9.3005
R1224 VTAIL.n81 VTAIL.n80 9.3005
R1225 VTAIL.n83 VTAIL.n82 9.3005
R1226 VTAIL.n74 VTAIL.n73 9.3005
R1227 VTAIL.n89 VTAIL.n88 9.3005
R1228 VTAIL.n91 VTAIL.n90 9.3005
R1229 VTAIL.n70 VTAIL.n69 9.3005
R1230 VTAIL.n98 VTAIL.n97 9.3005
R1231 VTAIL.n100 VTAIL.n99 9.3005
R1232 VTAIL.n175 VTAIL.n174 9.3005
R1233 VTAIL.n122 VTAIL.n121 9.3005
R1234 VTAIL.n169 VTAIL.n168 9.3005
R1235 VTAIL.n167 VTAIL.n166 9.3005
R1236 VTAIL.n126 VTAIL.n125 9.3005
R1237 VTAIL.n141 VTAIL.n140 9.3005
R1238 VTAIL.n143 VTAIL.n142 9.3005
R1239 VTAIL.n134 VTAIL.n133 9.3005
R1240 VTAIL.n149 VTAIL.n148 9.3005
R1241 VTAIL.n151 VTAIL.n150 9.3005
R1242 VTAIL.n130 VTAIL.n129 9.3005
R1243 VTAIL.n158 VTAIL.n157 9.3005
R1244 VTAIL.n160 VTAIL.n159 9.3005
R1245 VTAIL.n378 VTAIL.n377 9.3005
R1246 VTAIL.n380 VTAIL.n379 9.3005
R1247 VTAIL.n371 VTAIL.n370 9.3005
R1248 VTAIL.n386 VTAIL.n385 9.3005
R1249 VTAIL.n388 VTAIL.n387 9.3005
R1250 VTAIL.n366 VTAIL.n365 9.3005
R1251 VTAIL.n394 VTAIL.n393 9.3005
R1252 VTAIL.n396 VTAIL.n395 9.3005
R1253 VTAIL.n411 VTAIL.n410 9.3005
R1254 VTAIL.n358 VTAIL.n357 9.3005
R1255 VTAIL.n405 VTAIL.n404 9.3005
R1256 VTAIL.n403 VTAIL.n402 9.3005
R1257 VTAIL.n362 VTAIL.n361 9.3005
R1258 VTAIL.n318 VTAIL.n317 9.3005
R1259 VTAIL.n320 VTAIL.n319 9.3005
R1260 VTAIL.n311 VTAIL.n310 9.3005
R1261 VTAIL.n326 VTAIL.n325 9.3005
R1262 VTAIL.n328 VTAIL.n327 9.3005
R1263 VTAIL.n306 VTAIL.n305 9.3005
R1264 VTAIL.n334 VTAIL.n333 9.3005
R1265 VTAIL.n336 VTAIL.n335 9.3005
R1266 VTAIL.n351 VTAIL.n350 9.3005
R1267 VTAIL.n298 VTAIL.n297 9.3005
R1268 VTAIL.n345 VTAIL.n344 9.3005
R1269 VTAIL.n343 VTAIL.n342 9.3005
R1270 VTAIL.n302 VTAIL.n301 9.3005
R1271 VTAIL.n260 VTAIL.n259 9.3005
R1272 VTAIL.n262 VTAIL.n261 9.3005
R1273 VTAIL.n253 VTAIL.n252 9.3005
R1274 VTAIL.n268 VTAIL.n267 9.3005
R1275 VTAIL.n270 VTAIL.n269 9.3005
R1276 VTAIL.n248 VTAIL.n247 9.3005
R1277 VTAIL.n276 VTAIL.n275 9.3005
R1278 VTAIL.n278 VTAIL.n277 9.3005
R1279 VTAIL.n293 VTAIL.n292 9.3005
R1280 VTAIL.n240 VTAIL.n239 9.3005
R1281 VTAIL.n287 VTAIL.n286 9.3005
R1282 VTAIL.n285 VTAIL.n284 9.3005
R1283 VTAIL.n244 VTAIL.n243 9.3005
R1284 VTAIL.n200 VTAIL.n199 9.3005
R1285 VTAIL.n202 VTAIL.n201 9.3005
R1286 VTAIL.n193 VTAIL.n192 9.3005
R1287 VTAIL.n208 VTAIL.n207 9.3005
R1288 VTAIL.n210 VTAIL.n209 9.3005
R1289 VTAIL.n188 VTAIL.n187 9.3005
R1290 VTAIL.n216 VTAIL.n215 9.3005
R1291 VTAIL.n218 VTAIL.n217 9.3005
R1292 VTAIL.n233 VTAIL.n232 9.3005
R1293 VTAIL.n180 VTAIL.n179 9.3005
R1294 VTAIL.n227 VTAIL.n226 9.3005
R1295 VTAIL.n225 VTAIL.n224 9.3005
R1296 VTAIL.n184 VTAIL.n183 9.3005
R1297 VTAIL.n438 VTAIL.n428 8.92171
R1298 VTAIL.n26 VTAIL.n16 8.92171
R1299 VTAIL.n84 VTAIL.n74 8.92171
R1300 VTAIL.n144 VTAIL.n134 8.92171
R1301 VTAIL.n381 VTAIL.n371 8.92171
R1302 VTAIL.n321 VTAIL.n311 8.92171
R1303 VTAIL.n263 VTAIL.n253 8.92171
R1304 VTAIL.n203 VTAIL.n193 8.92171
R1305 VTAIL.n437 VTAIL.n430 8.14595
R1306 VTAIL.n25 VTAIL.n18 8.14595
R1307 VTAIL.n83 VTAIL.n76 8.14595
R1308 VTAIL.n143 VTAIL.n136 8.14595
R1309 VTAIL.n380 VTAIL.n373 8.14595
R1310 VTAIL.n320 VTAIL.n313 8.14595
R1311 VTAIL.n262 VTAIL.n255 8.14595
R1312 VTAIL.n202 VTAIL.n195 8.14595
R1313 VTAIL.n434 VTAIL.n433 7.3702
R1314 VTAIL.n22 VTAIL.n21 7.3702
R1315 VTAIL.n80 VTAIL.n79 7.3702
R1316 VTAIL.n140 VTAIL.n139 7.3702
R1317 VTAIL.n377 VTAIL.n376 7.3702
R1318 VTAIL.n317 VTAIL.n316 7.3702
R1319 VTAIL.n259 VTAIL.n258 7.3702
R1320 VTAIL.n199 VTAIL.n198 7.3702
R1321 VTAIL.n434 VTAIL.n430 5.81868
R1322 VTAIL.n22 VTAIL.n18 5.81868
R1323 VTAIL.n80 VTAIL.n76 5.81868
R1324 VTAIL.n140 VTAIL.n136 5.81868
R1325 VTAIL.n377 VTAIL.n373 5.81868
R1326 VTAIL.n317 VTAIL.n313 5.81868
R1327 VTAIL.n259 VTAIL.n255 5.81868
R1328 VTAIL.n199 VTAIL.n195 5.81868
R1329 VTAIL.n438 VTAIL.n437 5.04292
R1330 VTAIL.n26 VTAIL.n25 5.04292
R1331 VTAIL.n84 VTAIL.n83 5.04292
R1332 VTAIL.n144 VTAIL.n143 5.04292
R1333 VTAIL.n381 VTAIL.n380 5.04292
R1334 VTAIL.n321 VTAIL.n320 5.04292
R1335 VTAIL.n263 VTAIL.n262 5.04292
R1336 VTAIL.n203 VTAIL.n202 5.04292
R1337 VTAIL.n441 VTAIL.n428 4.26717
R1338 VTAIL.n470 VTAIL.n414 4.26717
R1339 VTAIL.n29 VTAIL.n16 4.26717
R1340 VTAIL.n58 VTAIL.n2 4.26717
R1341 VTAIL.n87 VTAIL.n74 4.26717
R1342 VTAIL.n116 VTAIL.n60 4.26717
R1343 VTAIL.n147 VTAIL.n134 4.26717
R1344 VTAIL.n176 VTAIL.n120 4.26717
R1345 VTAIL.n412 VTAIL.n356 4.26717
R1346 VTAIL.n384 VTAIL.n371 4.26717
R1347 VTAIL.n352 VTAIL.n296 4.26717
R1348 VTAIL.n324 VTAIL.n311 4.26717
R1349 VTAIL.n294 VTAIL.n238 4.26717
R1350 VTAIL.n266 VTAIL.n253 4.26717
R1351 VTAIL.n234 VTAIL.n178 4.26717
R1352 VTAIL.n206 VTAIL.n193 4.26717
R1353 VTAIL.n442 VTAIL.n426 3.49141
R1354 VTAIL.n468 VTAIL.n467 3.49141
R1355 VTAIL.n30 VTAIL.n14 3.49141
R1356 VTAIL.n56 VTAIL.n55 3.49141
R1357 VTAIL.n88 VTAIL.n72 3.49141
R1358 VTAIL.n114 VTAIL.n113 3.49141
R1359 VTAIL.n148 VTAIL.n132 3.49141
R1360 VTAIL.n174 VTAIL.n173 3.49141
R1361 VTAIL.n410 VTAIL.n409 3.49141
R1362 VTAIL.n385 VTAIL.n369 3.49141
R1363 VTAIL.n350 VTAIL.n349 3.49141
R1364 VTAIL.n325 VTAIL.n309 3.49141
R1365 VTAIL.n292 VTAIL.n291 3.49141
R1366 VTAIL.n267 VTAIL.n251 3.49141
R1367 VTAIL.n232 VTAIL.n231 3.49141
R1368 VTAIL.n207 VTAIL.n191 3.49141
R1369 VTAIL.n0 VTAIL.t4 3.02704
R1370 VTAIL.n0 VTAIL.t3 3.02704
R1371 VTAIL.n118 VTAIL.t9 3.02704
R1372 VTAIL.n118 VTAIL.t13 3.02704
R1373 VTAIL.n354 VTAIL.t14 3.02704
R1374 VTAIL.n354 VTAIL.t10 3.02704
R1375 VTAIL.n236 VTAIL.t5 3.02704
R1376 VTAIL.n236 VTAIL.t0 3.02704
R1377 VTAIL.n446 VTAIL.n445 2.71565
R1378 VTAIL.n464 VTAIL.n416 2.71565
R1379 VTAIL.n34 VTAIL.n33 2.71565
R1380 VTAIL.n52 VTAIL.n4 2.71565
R1381 VTAIL.n92 VTAIL.n91 2.71565
R1382 VTAIL.n110 VTAIL.n62 2.71565
R1383 VTAIL.n152 VTAIL.n151 2.71565
R1384 VTAIL.n170 VTAIL.n122 2.71565
R1385 VTAIL.n406 VTAIL.n358 2.71565
R1386 VTAIL.n389 VTAIL.n388 2.71565
R1387 VTAIL.n346 VTAIL.n298 2.71565
R1388 VTAIL.n329 VTAIL.n328 2.71565
R1389 VTAIL.n288 VTAIL.n240 2.71565
R1390 VTAIL.n271 VTAIL.n270 2.71565
R1391 VTAIL.n228 VTAIL.n180 2.71565
R1392 VTAIL.n211 VTAIL.n210 2.71565
R1393 VTAIL.n435 VTAIL.n431 2.41282
R1394 VTAIL.n23 VTAIL.n19 2.41282
R1395 VTAIL.n81 VTAIL.n77 2.41282
R1396 VTAIL.n141 VTAIL.n137 2.41282
R1397 VTAIL.n378 VTAIL.n374 2.41282
R1398 VTAIL.n318 VTAIL.n314 2.41282
R1399 VTAIL.n260 VTAIL.n256 2.41282
R1400 VTAIL.n200 VTAIL.n196 2.41282
R1401 VTAIL.n450 VTAIL.n424 1.93989
R1402 VTAIL.n463 VTAIL.n418 1.93989
R1403 VTAIL.n38 VTAIL.n12 1.93989
R1404 VTAIL.n51 VTAIL.n6 1.93989
R1405 VTAIL.n96 VTAIL.n70 1.93989
R1406 VTAIL.n109 VTAIL.n64 1.93989
R1407 VTAIL.n156 VTAIL.n130 1.93989
R1408 VTAIL.n169 VTAIL.n124 1.93989
R1409 VTAIL.n405 VTAIL.n360 1.93989
R1410 VTAIL.n392 VTAIL.n366 1.93989
R1411 VTAIL.n345 VTAIL.n300 1.93989
R1412 VTAIL.n332 VTAIL.n306 1.93989
R1413 VTAIL.n287 VTAIL.n242 1.93989
R1414 VTAIL.n274 VTAIL.n248 1.93989
R1415 VTAIL.n227 VTAIL.n182 1.93989
R1416 VTAIL.n214 VTAIL.n188 1.93989
R1417 VTAIL.n451 VTAIL.n422 1.16414
R1418 VTAIL.n460 VTAIL.n459 1.16414
R1419 VTAIL.n39 VTAIL.n10 1.16414
R1420 VTAIL.n48 VTAIL.n47 1.16414
R1421 VTAIL.n97 VTAIL.n68 1.16414
R1422 VTAIL.n106 VTAIL.n105 1.16414
R1423 VTAIL.n157 VTAIL.n128 1.16414
R1424 VTAIL.n166 VTAIL.n165 1.16414
R1425 VTAIL.n402 VTAIL.n401 1.16414
R1426 VTAIL.n393 VTAIL.n364 1.16414
R1427 VTAIL.n342 VTAIL.n341 1.16414
R1428 VTAIL.n333 VTAIL.n304 1.16414
R1429 VTAIL.n284 VTAIL.n283 1.16414
R1430 VTAIL.n275 VTAIL.n246 1.16414
R1431 VTAIL.n224 VTAIL.n223 1.16414
R1432 VTAIL.n215 VTAIL.n186 1.16414
R1433 VTAIL.n237 VTAIL.n235 0.845328
R1434 VTAIL.n295 VTAIL.n237 0.845328
R1435 VTAIL.n355 VTAIL.n353 0.845328
R1436 VTAIL.n413 VTAIL.n355 0.845328
R1437 VTAIL.n177 VTAIL.n119 0.845328
R1438 VTAIL.n119 VTAIL.n117 0.845328
R1439 VTAIL.n59 VTAIL.n1 0.845328
R1440 VTAIL VTAIL.n471 0.787138
R1441 VTAIL.n353 VTAIL.n295 0.470328
R1442 VTAIL.n117 VTAIL.n59 0.470328
R1443 VTAIL.n455 VTAIL.n454 0.388379
R1444 VTAIL.n456 VTAIL.n420 0.388379
R1445 VTAIL.n43 VTAIL.n42 0.388379
R1446 VTAIL.n44 VTAIL.n8 0.388379
R1447 VTAIL.n101 VTAIL.n100 0.388379
R1448 VTAIL.n102 VTAIL.n66 0.388379
R1449 VTAIL.n161 VTAIL.n160 0.388379
R1450 VTAIL.n162 VTAIL.n126 0.388379
R1451 VTAIL.n398 VTAIL.n362 0.388379
R1452 VTAIL.n397 VTAIL.n396 0.388379
R1453 VTAIL.n338 VTAIL.n302 0.388379
R1454 VTAIL.n337 VTAIL.n336 0.388379
R1455 VTAIL.n280 VTAIL.n244 0.388379
R1456 VTAIL.n279 VTAIL.n278 0.388379
R1457 VTAIL.n220 VTAIL.n184 0.388379
R1458 VTAIL.n219 VTAIL.n218 0.388379
R1459 VTAIL.n436 VTAIL.n435 0.155672
R1460 VTAIL.n436 VTAIL.n427 0.155672
R1461 VTAIL.n443 VTAIL.n427 0.155672
R1462 VTAIL.n444 VTAIL.n443 0.155672
R1463 VTAIL.n444 VTAIL.n423 0.155672
R1464 VTAIL.n452 VTAIL.n423 0.155672
R1465 VTAIL.n453 VTAIL.n452 0.155672
R1466 VTAIL.n453 VTAIL.n419 0.155672
R1467 VTAIL.n461 VTAIL.n419 0.155672
R1468 VTAIL.n462 VTAIL.n461 0.155672
R1469 VTAIL.n462 VTAIL.n415 0.155672
R1470 VTAIL.n469 VTAIL.n415 0.155672
R1471 VTAIL.n24 VTAIL.n23 0.155672
R1472 VTAIL.n24 VTAIL.n15 0.155672
R1473 VTAIL.n31 VTAIL.n15 0.155672
R1474 VTAIL.n32 VTAIL.n31 0.155672
R1475 VTAIL.n32 VTAIL.n11 0.155672
R1476 VTAIL.n40 VTAIL.n11 0.155672
R1477 VTAIL.n41 VTAIL.n40 0.155672
R1478 VTAIL.n41 VTAIL.n7 0.155672
R1479 VTAIL.n49 VTAIL.n7 0.155672
R1480 VTAIL.n50 VTAIL.n49 0.155672
R1481 VTAIL.n50 VTAIL.n3 0.155672
R1482 VTAIL.n57 VTAIL.n3 0.155672
R1483 VTAIL.n82 VTAIL.n81 0.155672
R1484 VTAIL.n82 VTAIL.n73 0.155672
R1485 VTAIL.n89 VTAIL.n73 0.155672
R1486 VTAIL.n90 VTAIL.n89 0.155672
R1487 VTAIL.n90 VTAIL.n69 0.155672
R1488 VTAIL.n98 VTAIL.n69 0.155672
R1489 VTAIL.n99 VTAIL.n98 0.155672
R1490 VTAIL.n99 VTAIL.n65 0.155672
R1491 VTAIL.n107 VTAIL.n65 0.155672
R1492 VTAIL.n108 VTAIL.n107 0.155672
R1493 VTAIL.n108 VTAIL.n61 0.155672
R1494 VTAIL.n115 VTAIL.n61 0.155672
R1495 VTAIL.n142 VTAIL.n141 0.155672
R1496 VTAIL.n142 VTAIL.n133 0.155672
R1497 VTAIL.n149 VTAIL.n133 0.155672
R1498 VTAIL.n150 VTAIL.n149 0.155672
R1499 VTAIL.n150 VTAIL.n129 0.155672
R1500 VTAIL.n158 VTAIL.n129 0.155672
R1501 VTAIL.n159 VTAIL.n158 0.155672
R1502 VTAIL.n159 VTAIL.n125 0.155672
R1503 VTAIL.n167 VTAIL.n125 0.155672
R1504 VTAIL.n168 VTAIL.n167 0.155672
R1505 VTAIL.n168 VTAIL.n121 0.155672
R1506 VTAIL.n175 VTAIL.n121 0.155672
R1507 VTAIL.n411 VTAIL.n357 0.155672
R1508 VTAIL.n404 VTAIL.n357 0.155672
R1509 VTAIL.n404 VTAIL.n403 0.155672
R1510 VTAIL.n403 VTAIL.n361 0.155672
R1511 VTAIL.n395 VTAIL.n361 0.155672
R1512 VTAIL.n395 VTAIL.n394 0.155672
R1513 VTAIL.n394 VTAIL.n365 0.155672
R1514 VTAIL.n387 VTAIL.n365 0.155672
R1515 VTAIL.n387 VTAIL.n386 0.155672
R1516 VTAIL.n386 VTAIL.n370 0.155672
R1517 VTAIL.n379 VTAIL.n370 0.155672
R1518 VTAIL.n379 VTAIL.n378 0.155672
R1519 VTAIL.n351 VTAIL.n297 0.155672
R1520 VTAIL.n344 VTAIL.n297 0.155672
R1521 VTAIL.n344 VTAIL.n343 0.155672
R1522 VTAIL.n343 VTAIL.n301 0.155672
R1523 VTAIL.n335 VTAIL.n301 0.155672
R1524 VTAIL.n335 VTAIL.n334 0.155672
R1525 VTAIL.n334 VTAIL.n305 0.155672
R1526 VTAIL.n327 VTAIL.n305 0.155672
R1527 VTAIL.n327 VTAIL.n326 0.155672
R1528 VTAIL.n326 VTAIL.n310 0.155672
R1529 VTAIL.n319 VTAIL.n310 0.155672
R1530 VTAIL.n319 VTAIL.n318 0.155672
R1531 VTAIL.n293 VTAIL.n239 0.155672
R1532 VTAIL.n286 VTAIL.n239 0.155672
R1533 VTAIL.n286 VTAIL.n285 0.155672
R1534 VTAIL.n285 VTAIL.n243 0.155672
R1535 VTAIL.n277 VTAIL.n243 0.155672
R1536 VTAIL.n277 VTAIL.n276 0.155672
R1537 VTAIL.n276 VTAIL.n247 0.155672
R1538 VTAIL.n269 VTAIL.n247 0.155672
R1539 VTAIL.n269 VTAIL.n268 0.155672
R1540 VTAIL.n268 VTAIL.n252 0.155672
R1541 VTAIL.n261 VTAIL.n252 0.155672
R1542 VTAIL.n261 VTAIL.n260 0.155672
R1543 VTAIL.n233 VTAIL.n179 0.155672
R1544 VTAIL.n226 VTAIL.n179 0.155672
R1545 VTAIL.n226 VTAIL.n225 0.155672
R1546 VTAIL.n225 VTAIL.n183 0.155672
R1547 VTAIL.n217 VTAIL.n183 0.155672
R1548 VTAIL.n217 VTAIL.n216 0.155672
R1549 VTAIL.n216 VTAIL.n187 0.155672
R1550 VTAIL.n209 VTAIL.n187 0.155672
R1551 VTAIL.n209 VTAIL.n208 0.155672
R1552 VTAIL.n208 VTAIL.n192 0.155672
R1553 VTAIL.n201 VTAIL.n192 0.155672
R1554 VTAIL.n201 VTAIL.n200 0.155672
R1555 VTAIL VTAIL.n1 0.0586897
R1556 VDD1 VDD1.n0 77.5104
R1557 VDD1.n3 VDD1.n2 77.3967
R1558 VDD1.n3 VDD1.n1 77.3967
R1559 VDD1.n5 VDD1.n4 77.0296
R1560 VDD1.n5 VDD1.n3 37.3586
R1561 VDD1.n4 VDD1.t1 3.02704
R1562 VDD1.n4 VDD1.t5 3.02704
R1563 VDD1.n0 VDD1.t6 3.02704
R1564 VDD1.n0 VDD1.t0 3.02704
R1565 VDD1.n2 VDD1.t4 3.02704
R1566 VDD1.n2 VDD1.t7 3.02704
R1567 VDD1.n1 VDD1.t2 3.02704
R1568 VDD1.n1 VDD1.t3 3.02704
R1569 VDD1 VDD1.n5 0.364724
R1570 VN.n1 VN.t4 486.204
R1571 VN.n7 VN.t2 486.204
R1572 VN.n2 VN.t7 459.384
R1573 VN.n3 VN.t6 459.384
R1574 VN.n4 VN.t1 459.384
R1575 VN.n8 VN.t0 459.384
R1576 VN.n9 VN.t5 459.384
R1577 VN.n10 VN.t3 459.384
R1578 VN.n5 VN.n4 161.3
R1579 VN.n11 VN.n10 161.3
R1580 VN.n9 VN.n6 80.6037
R1581 VN.n3 VN.n0 80.6037
R1582 VN.n3 VN.n2 48.2005
R1583 VN.n4 VN.n3 48.2005
R1584 VN.n9 VN.n8 48.2005
R1585 VN.n10 VN.n9 48.2005
R1586 VN.n7 VN.n6 45.2318
R1587 VN.n1 VN.n0 45.2318
R1588 VN VN.n11 41.3054
R1589 VN.n8 VN.n7 13.3799
R1590 VN.n2 VN.n1 13.3799
R1591 VN.n11 VN.n6 0.285035
R1592 VN.n5 VN.n0 0.285035
R1593 VN VN.n5 0.0516364
R1594 VDD2.n2 VDD2.n1 77.3967
R1595 VDD2.n2 VDD2.n0 77.3967
R1596 VDD2 VDD2.n5 77.3938
R1597 VDD2.n4 VDD2.n3 77.0298
R1598 VDD2.n4 VDD2.n2 36.7756
R1599 VDD2.n5 VDD2.t7 3.02704
R1600 VDD2.n5 VDD2.t5 3.02704
R1601 VDD2.n3 VDD2.t4 3.02704
R1602 VDD2.n3 VDD2.t2 3.02704
R1603 VDD2.n1 VDD2.t1 3.02704
R1604 VDD2.n1 VDD2.t6 3.02704
R1605 VDD2.n0 VDD2.t3 3.02704
R1606 VDD2.n0 VDD2.t0 3.02704
R1607 VDD2 VDD2.n4 0.481103
C0 VP B 1.15689f
C1 VDD1 VN 0.147912f
C2 VTAIL B 3.46222f
C3 VDD2 B 1.05591f
C4 VDD1 w_n1950_n3116# 1.24835f
C5 VN w_n1950_n3116# 3.3903f
C6 VDD1 B 1.02079f
C7 B VN 0.752557f
C8 VP VTAIL 4.57665f
C9 VDD2 VP 0.31188f
C10 VDD2 VTAIL 10.5099f
C11 B w_n1950_n3116# 6.77882f
C12 VP VDD1 4.94033f
C13 VTAIL VDD1 10.4685f
C14 VDD2 VDD1 0.801833f
C15 VP VN 5.04358f
C16 VTAIL VN 4.56254f
C17 VDD2 VN 4.77677f
C18 VP w_n1950_n3116# 3.6377f
C19 VTAIL w_n1950_n3116# 3.90302f
C20 VDD2 w_n1950_n3116# 1.28112f
C21 VDD2 VSUBS 1.289471f
C22 VDD1 VSUBS 1.585937f
C23 VTAIL VSUBS 0.822149f
C24 VN VSUBS 4.55056f
C25 VP VSUBS 1.556731f
C26 B VSUBS 2.716571f
C27 w_n1950_n3116# VSUBS 74.9502f
C28 VDD2.t3 VSUBS 0.234729f
C29 VDD2.t0 VSUBS 0.234729f
C30 VDD2.n0 VSUBS 1.80289f
C31 VDD2.t1 VSUBS 0.234729f
C32 VDD2.t6 VSUBS 0.234729f
C33 VDD2.n1 VSUBS 1.80289f
C34 VDD2.n2 VSUBS 2.83636f
C35 VDD2.t4 VSUBS 0.234729f
C36 VDD2.t2 VSUBS 0.234729f
C37 VDD2.n3 VSUBS 1.79993f
C38 VDD2.n4 VSUBS 2.68206f
C39 VDD2.t7 VSUBS 0.234729f
C40 VDD2.t5 VSUBS 0.234729f
C41 VDD2.n5 VSUBS 1.80286f
C42 VN.n0 VSUBS 0.279925f
C43 VN.t4 VSUBS 1.14298f
C44 VN.n1 VSUBS 0.43305f
C45 VN.t7 VSUBS 1.11779f
C46 VN.n2 VSUBS 0.469202f
C47 VN.t6 VSUBS 1.11779f
C48 VN.n3 VSUBS 0.469202f
C49 VN.t1 VSUBS 1.11779f
C50 VN.n4 VSUBS 0.456493f
C51 VN.n5 VSUBS 0.062129f
C52 VN.n6 VSUBS 0.279925f
C53 VN.t0 VSUBS 1.11779f
C54 VN.t2 VSUBS 1.14298f
C55 VN.n7 VSUBS 0.43305f
C56 VN.n8 VSUBS 0.469202f
C57 VN.t5 VSUBS 1.11779f
C58 VN.n9 VSUBS 0.469202f
C59 VN.t3 VSUBS 1.11779f
C60 VN.n10 VSUBS 0.456493f
C61 VN.n11 VSUBS 2.2687f
C62 VDD1.t6 VSUBS 0.234697f
C63 VDD1.t0 VSUBS 0.234697f
C64 VDD1.n0 VSUBS 1.80361f
C65 VDD1.t2 VSUBS 0.234697f
C66 VDD1.t3 VSUBS 0.234697f
C67 VDD1.n1 VSUBS 1.80264f
C68 VDD1.t4 VSUBS 0.234697f
C69 VDD1.t7 VSUBS 0.234697f
C70 VDD1.n2 VSUBS 1.80264f
C71 VDD1.n3 VSUBS 2.89509f
C72 VDD1.t1 VSUBS 0.234697f
C73 VDD1.t5 VSUBS 0.234697f
C74 VDD1.n4 VSUBS 1.79967f
C75 VDD1.n5 VSUBS 2.71433f
C76 VTAIL.t4 VSUBS 0.217006f
C77 VTAIL.t3 VSUBS 0.217006f
C78 VTAIL.n0 VSUBS 1.53661f
C79 VTAIL.n1 VSUBS 0.632942f
C80 VTAIL.n2 VSUBS 0.027771f
C81 VTAIL.n3 VSUBS 0.025569f
C82 VTAIL.n4 VSUBS 0.01374f
C83 VTAIL.n5 VSUBS 0.032476f
C84 VTAIL.n6 VSUBS 0.014548f
C85 VTAIL.n7 VSUBS 0.025569f
C86 VTAIL.n8 VSUBS 0.01374f
C87 VTAIL.n9 VSUBS 0.032476f
C88 VTAIL.n10 VSUBS 0.014548f
C89 VTAIL.n11 VSUBS 0.025569f
C90 VTAIL.n12 VSUBS 0.01374f
C91 VTAIL.n13 VSUBS 0.032476f
C92 VTAIL.n14 VSUBS 0.014548f
C93 VTAIL.n15 VSUBS 0.025569f
C94 VTAIL.n16 VSUBS 0.01374f
C95 VTAIL.n17 VSUBS 0.032476f
C96 VTAIL.n18 VSUBS 0.014548f
C97 VTAIL.n19 VSUBS 0.186813f
C98 VTAIL.t6 VSUBS 0.069883f
C99 VTAIL.n20 VSUBS 0.024357f
C100 VTAIL.n21 VSUBS 0.02443f
C101 VTAIL.n22 VSUBS 0.01374f
C102 VTAIL.n23 VSUBS 1.1151f
C103 VTAIL.n24 VSUBS 0.025569f
C104 VTAIL.n25 VSUBS 0.01374f
C105 VTAIL.n26 VSUBS 0.014548f
C106 VTAIL.n27 VSUBS 0.032476f
C107 VTAIL.n28 VSUBS 0.032476f
C108 VTAIL.n29 VSUBS 0.014548f
C109 VTAIL.n30 VSUBS 0.01374f
C110 VTAIL.n31 VSUBS 0.025569f
C111 VTAIL.n32 VSUBS 0.025569f
C112 VTAIL.n33 VSUBS 0.01374f
C113 VTAIL.n34 VSUBS 0.014548f
C114 VTAIL.n35 VSUBS 0.032476f
C115 VTAIL.n36 VSUBS 0.032476f
C116 VTAIL.n37 VSUBS 0.032476f
C117 VTAIL.n38 VSUBS 0.014548f
C118 VTAIL.n39 VSUBS 0.01374f
C119 VTAIL.n40 VSUBS 0.025569f
C120 VTAIL.n41 VSUBS 0.025569f
C121 VTAIL.n42 VSUBS 0.01374f
C122 VTAIL.n43 VSUBS 0.014144f
C123 VTAIL.n44 VSUBS 0.014144f
C124 VTAIL.n45 VSUBS 0.032476f
C125 VTAIL.n46 VSUBS 0.032476f
C126 VTAIL.n47 VSUBS 0.014548f
C127 VTAIL.n48 VSUBS 0.01374f
C128 VTAIL.n49 VSUBS 0.025569f
C129 VTAIL.n50 VSUBS 0.025569f
C130 VTAIL.n51 VSUBS 0.01374f
C131 VTAIL.n52 VSUBS 0.014548f
C132 VTAIL.n53 VSUBS 0.032476f
C133 VTAIL.n54 VSUBS 0.077517f
C134 VTAIL.n55 VSUBS 0.014548f
C135 VTAIL.n56 VSUBS 0.01374f
C136 VTAIL.n57 VSUBS 0.061197f
C137 VTAIL.n58 VSUBS 0.038997f
C138 VTAIL.n59 VSUBS 0.131335f
C139 VTAIL.n60 VSUBS 0.027771f
C140 VTAIL.n61 VSUBS 0.025569f
C141 VTAIL.n62 VSUBS 0.01374f
C142 VTAIL.n63 VSUBS 0.032476f
C143 VTAIL.n64 VSUBS 0.014548f
C144 VTAIL.n65 VSUBS 0.025569f
C145 VTAIL.n66 VSUBS 0.01374f
C146 VTAIL.n67 VSUBS 0.032476f
C147 VTAIL.n68 VSUBS 0.014548f
C148 VTAIL.n69 VSUBS 0.025569f
C149 VTAIL.n70 VSUBS 0.01374f
C150 VTAIL.n71 VSUBS 0.032476f
C151 VTAIL.n72 VSUBS 0.014548f
C152 VTAIL.n73 VSUBS 0.025569f
C153 VTAIL.n74 VSUBS 0.01374f
C154 VTAIL.n75 VSUBS 0.032476f
C155 VTAIL.n76 VSUBS 0.014548f
C156 VTAIL.n77 VSUBS 0.186813f
C157 VTAIL.t11 VSUBS 0.069883f
C158 VTAIL.n78 VSUBS 0.024357f
C159 VTAIL.n79 VSUBS 0.02443f
C160 VTAIL.n80 VSUBS 0.01374f
C161 VTAIL.n81 VSUBS 1.1151f
C162 VTAIL.n82 VSUBS 0.025569f
C163 VTAIL.n83 VSUBS 0.01374f
C164 VTAIL.n84 VSUBS 0.014548f
C165 VTAIL.n85 VSUBS 0.032476f
C166 VTAIL.n86 VSUBS 0.032476f
C167 VTAIL.n87 VSUBS 0.014548f
C168 VTAIL.n88 VSUBS 0.01374f
C169 VTAIL.n89 VSUBS 0.025569f
C170 VTAIL.n90 VSUBS 0.025569f
C171 VTAIL.n91 VSUBS 0.01374f
C172 VTAIL.n92 VSUBS 0.014548f
C173 VTAIL.n93 VSUBS 0.032476f
C174 VTAIL.n94 VSUBS 0.032476f
C175 VTAIL.n95 VSUBS 0.032476f
C176 VTAIL.n96 VSUBS 0.014548f
C177 VTAIL.n97 VSUBS 0.01374f
C178 VTAIL.n98 VSUBS 0.025569f
C179 VTAIL.n99 VSUBS 0.025569f
C180 VTAIL.n100 VSUBS 0.01374f
C181 VTAIL.n101 VSUBS 0.014144f
C182 VTAIL.n102 VSUBS 0.014144f
C183 VTAIL.n103 VSUBS 0.032476f
C184 VTAIL.n104 VSUBS 0.032476f
C185 VTAIL.n105 VSUBS 0.014548f
C186 VTAIL.n106 VSUBS 0.01374f
C187 VTAIL.n107 VSUBS 0.025569f
C188 VTAIL.n108 VSUBS 0.025569f
C189 VTAIL.n109 VSUBS 0.01374f
C190 VTAIL.n110 VSUBS 0.014548f
C191 VTAIL.n111 VSUBS 0.032476f
C192 VTAIL.n112 VSUBS 0.077517f
C193 VTAIL.n113 VSUBS 0.014548f
C194 VTAIL.n114 VSUBS 0.01374f
C195 VTAIL.n115 VSUBS 0.061197f
C196 VTAIL.n116 VSUBS 0.038997f
C197 VTAIL.n117 VSUBS 0.131335f
C198 VTAIL.t9 VSUBS 0.217006f
C199 VTAIL.t13 VSUBS 0.217006f
C200 VTAIL.n118 VSUBS 1.53661f
C201 VTAIL.n119 VSUBS 0.697753f
C202 VTAIL.n120 VSUBS 0.027771f
C203 VTAIL.n121 VSUBS 0.025569f
C204 VTAIL.n122 VSUBS 0.01374f
C205 VTAIL.n123 VSUBS 0.032476f
C206 VTAIL.n124 VSUBS 0.014548f
C207 VTAIL.n125 VSUBS 0.025569f
C208 VTAIL.n126 VSUBS 0.01374f
C209 VTAIL.n127 VSUBS 0.032476f
C210 VTAIL.n128 VSUBS 0.014548f
C211 VTAIL.n129 VSUBS 0.025569f
C212 VTAIL.n130 VSUBS 0.01374f
C213 VTAIL.n131 VSUBS 0.032476f
C214 VTAIL.n132 VSUBS 0.014548f
C215 VTAIL.n133 VSUBS 0.025569f
C216 VTAIL.n134 VSUBS 0.01374f
C217 VTAIL.n135 VSUBS 0.032476f
C218 VTAIL.n136 VSUBS 0.014548f
C219 VTAIL.n137 VSUBS 0.186813f
C220 VTAIL.t7 VSUBS 0.069883f
C221 VTAIL.n138 VSUBS 0.024357f
C222 VTAIL.n139 VSUBS 0.02443f
C223 VTAIL.n140 VSUBS 0.01374f
C224 VTAIL.n141 VSUBS 1.1151f
C225 VTAIL.n142 VSUBS 0.025569f
C226 VTAIL.n143 VSUBS 0.01374f
C227 VTAIL.n144 VSUBS 0.014548f
C228 VTAIL.n145 VSUBS 0.032476f
C229 VTAIL.n146 VSUBS 0.032476f
C230 VTAIL.n147 VSUBS 0.014548f
C231 VTAIL.n148 VSUBS 0.01374f
C232 VTAIL.n149 VSUBS 0.025569f
C233 VTAIL.n150 VSUBS 0.025569f
C234 VTAIL.n151 VSUBS 0.01374f
C235 VTAIL.n152 VSUBS 0.014548f
C236 VTAIL.n153 VSUBS 0.032476f
C237 VTAIL.n154 VSUBS 0.032476f
C238 VTAIL.n155 VSUBS 0.032476f
C239 VTAIL.n156 VSUBS 0.014548f
C240 VTAIL.n157 VSUBS 0.01374f
C241 VTAIL.n158 VSUBS 0.025569f
C242 VTAIL.n159 VSUBS 0.025569f
C243 VTAIL.n160 VSUBS 0.01374f
C244 VTAIL.n161 VSUBS 0.014144f
C245 VTAIL.n162 VSUBS 0.014144f
C246 VTAIL.n163 VSUBS 0.032476f
C247 VTAIL.n164 VSUBS 0.032476f
C248 VTAIL.n165 VSUBS 0.014548f
C249 VTAIL.n166 VSUBS 0.01374f
C250 VTAIL.n167 VSUBS 0.025569f
C251 VTAIL.n168 VSUBS 0.025569f
C252 VTAIL.n169 VSUBS 0.01374f
C253 VTAIL.n170 VSUBS 0.014548f
C254 VTAIL.n171 VSUBS 0.032476f
C255 VTAIL.n172 VSUBS 0.077517f
C256 VTAIL.n173 VSUBS 0.014548f
C257 VTAIL.n174 VSUBS 0.01374f
C258 VTAIL.n175 VSUBS 0.061197f
C259 VTAIL.n176 VSUBS 0.038997f
C260 VTAIL.n177 VSUBS 1.27236f
C261 VTAIL.n178 VSUBS 0.027771f
C262 VTAIL.n179 VSUBS 0.025569f
C263 VTAIL.n180 VSUBS 0.01374f
C264 VTAIL.n181 VSUBS 0.032476f
C265 VTAIL.n182 VSUBS 0.014548f
C266 VTAIL.n183 VSUBS 0.025569f
C267 VTAIL.n184 VSUBS 0.01374f
C268 VTAIL.n185 VSUBS 0.032476f
C269 VTAIL.n186 VSUBS 0.014548f
C270 VTAIL.n187 VSUBS 0.025569f
C271 VTAIL.n188 VSUBS 0.01374f
C272 VTAIL.n189 VSUBS 0.032476f
C273 VTAIL.n190 VSUBS 0.032476f
C274 VTAIL.n191 VSUBS 0.014548f
C275 VTAIL.n192 VSUBS 0.025569f
C276 VTAIL.n193 VSUBS 0.01374f
C277 VTAIL.n194 VSUBS 0.032476f
C278 VTAIL.n195 VSUBS 0.014548f
C279 VTAIL.n196 VSUBS 0.186813f
C280 VTAIL.t2 VSUBS 0.069883f
C281 VTAIL.n197 VSUBS 0.024357f
C282 VTAIL.n198 VSUBS 0.02443f
C283 VTAIL.n199 VSUBS 0.01374f
C284 VTAIL.n200 VSUBS 1.1151f
C285 VTAIL.n201 VSUBS 0.025569f
C286 VTAIL.n202 VSUBS 0.01374f
C287 VTAIL.n203 VSUBS 0.014548f
C288 VTAIL.n204 VSUBS 0.032476f
C289 VTAIL.n205 VSUBS 0.032476f
C290 VTAIL.n206 VSUBS 0.014548f
C291 VTAIL.n207 VSUBS 0.01374f
C292 VTAIL.n208 VSUBS 0.025569f
C293 VTAIL.n209 VSUBS 0.025569f
C294 VTAIL.n210 VSUBS 0.01374f
C295 VTAIL.n211 VSUBS 0.014548f
C296 VTAIL.n212 VSUBS 0.032476f
C297 VTAIL.n213 VSUBS 0.032476f
C298 VTAIL.n214 VSUBS 0.014548f
C299 VTAIL.n215 VSUBS 0.01374f
C300 VTAIL.n216 VSUBS 0.025569f
C301 VTAIL.n217 VSUBS 0.025569f
C302 VTAIL.n218 VSUBS 0.01374f
C303 VTAIL.n219 VSUBS 0.014144f
C304 VTAIL.n220 VSUBS 0.014144f
C305 VTAIL.n221 VSUBS 0.032476f
C306 VTAIL.n222 VSUBS 0.032476f
C307 VTAIL.n223 VSUBS 0.014548f
C308 VTAIL.n224 VSUBS 0.01374f
C309 VTAIL.n225 VSUBS 0.025569f
C310 VTAIL.n226 VSUBS 0.025569f
C311 VTAIL.n227 VSUBS 0.01374f
C312 VTAIL.n228 VSUBS 0.014548f
C313 VTAIL.n229 VSUBS 0.032476f
C314 VTAIL.n230 VSUBS 0.077517f
C315 VTAIL.n231 VSUBS 0.014548f
C316 VTAIL.n232 VSUBS 0.01374f
C317 VTAIL.n233 VSUBS 0.061197f
C318 VTAIL.n234 VSUBS 0.038997f
C319 VTAIL.n235 VSUBS 1.27236f
C320 VTAIL.t5 VSUBS 0.217006f
C321 VTAIL.t0 VSUBS 0.217006f
C322 VTAIL.n236 VSUBS 1.53662f
C323 VTAIL.n237 VSUBS 0.697742f
C324 VTAIL.n238 VSUBS 0.027771f
C325 VTAIL.n239 VSUBS 0.025569f
C326 VTAIL.n240 VSUBS 0.01374f
C327 VTAIL.n241 VSUBS 0.032476f
C328 VTAIL.n242 VSUBS 0.014548f
C329 VTAIL.n243 VSUBS 0.025569f
C330 VTAIL.n244 VSUBS 0.01374f
C331 VTAIL.n245 VSUBS 0.032476f
C332 VTAIL.n246 VSUBS 0.014548f
C333 VTAIL.n247 VSUBS 0.025569f
C334 VTAIL.n248 VSUBS 0.01374f
C335 VTAIL.n249 VSUBS 0.032476f
C336 VTAIL.n250 VSUBS 0.032476f
C337 VTAIL.n251 VSUBS 0.014548f
C338 VTAIL.n252 VSUBS 0.025569f
C339 VTAIL.n253 VSUBS 0.01374f
C340 VTAIL.n254 VSUBS 0.032476f
C341 VTAIL.n255 VSUBS 0.014548f
C342 VTAIL.n256 VSUBS 0.186813f
C343 VTAIL.t1 VSUBS 0.069883f
C344 VTAIL.n257 VSUBS 0.024357f
C345 VTAIL.n258 VSUBS 0.02443f
C346 VTAIL.n259 VSUBS 0.01374f
C347 VTAIL.n260 VSUBS 1.1151f
C348 VTAIL.n261 VSUBS 0.025569f
C349 VTAIL.n262 VSUBS 0.01374f
C350 VTAIL.n263 VSUBS 0.014548f
C351 VTAIL.n264 VSUBS 0.032476f
C352 VTAIL.n265 VSUBS 0.032476f
C353 VTAIL.n266 VSUBS 0.014548f
C354 VTAIL.n267 VSUBS 0.01374f
C355 VTAIL.n268 VSUBS 0.025569f
C356 VTAIL.n269 VSUBS 0.025569f
C357 VTAIL.n270 VSUBS 0.01374f
C358 VTAIL.n271 VSUBS 0.014548f
C359 VTAIL.n272 VSUBS 0.032476f
C360 VTAIL.n273 VSUBS 0.032476f
C361 VTAIL.n274 VSUBS 0.014548f
C362 VTAIL.n275 VSUBS 0.01374f
C363 VTAIL.n276 VSUBS 0.025569f
C364 VTAIL.n277 VSUBS 0.025569f
C365 VTAIL.n278 VSUBS 0.01374f
C366 VTAIL.n279 VSUBS 0.014144f
C367 VTAIL.n280 VSUBS 0.014144f
C368 VTAIL.n281 VSUBS 0.032476f
C369 VTAIL.n282 VSUBS 0.032476f
C370 VTAIL.n283 VSUBS 0.014548f
C371 VTAIL.n284 VSUBS 0.01374f
C372 VTAIL.n285 VSUBS 0.025569f
C373 VTAIL.n286 VSUBS 0.025569f
C374 VTAIL.n287 VSUBS 0.01374f
C375 VTAIL.n288 VSUBS 0.014548f
C376 VTAIL.n289 VSUBS 0.032476f
C377 VTAIL.n290 VSUBS 0.077517f
C378 VTAIL.n291 VSUBS 0.014548f
C379 VTAIL.n292 VSUBS 0.01374f
C380 VTAIL.n293 VSUBS 0.061197f
C381 VTAIL.n294 VSUBS 0.038997f
C382 VTAIL.n295 VSUBS 0.131335f
C383 VTAIL.n296 VSUBS 0.027771f
C384 VTAIL.n297 VSUBS 0.025569f
C385 VTAIL.n298 VSUBS 0.01374f
C386 VTAIL.n299 VSUBS 0.032476f
C387 VTAIL.n300 VSUBS 0.014548f
C388 VTAIL.n301 VSUBS 0.025569f
C389 VTAIL.n302 VSUBS 0.01374f
C390 VTAIL.n303 VSUBS 0.032476f
C391 VTAIL.n304 VSUBS 0.014548f
C392 VTAIL.n305 VSUBS 0.025569f
C393 VTAIL.n306 VSUBS 0.01374f
C394 VTAIL.n307 VSUBS 0.032476f
C395 VTAIL.n308 VSUBS 0.032476f
C396 VTAIL.n309 VSUBS 0.014548f
C397 VTAIL.n310 VSUBS 0.025569f
C398 VTAIL.n311 VSUBS 0.01374f
C399 VTAIL.n312 VSUBS 0.032476f
C400 VTAIL.n313 VSUBS 0.014548f
C401 VTAIL.n314 VSUBS 0.186813f
C402 VTAIL.t8 VSUBS 0.069883f
C403 VTAIL.n315 VSUBS 0.024357f
C404 VTAIL.n316 VSUBS 0.02443f
C405 VTAIL.n317 VSUBS 0.01374f
C406 VTAIL.n318 VSUBS 1.1151f
C407 VTAIL.n319 VSUBS 0.025569f
C408 VTAIL.n320 VSUBS 0.01374f
C409 VTAIL.n321 VSUBS 0.014548f
C410 VTAIL.n322 VSUBS 0.032476f
C411 VTAIL.n323 VSUBS 0.032476f
C412 VTAIL.n324 VSUBS 0.014548f
C413 VTAIL.n325 VSUBS 0.01374f
C414 VTAIL.n326 VSUBS 0.025569f
C415 VTAIL.n327 VSUBS 0.025569f
C416 VTAIL.n328 VSUBS 0.01374f
C417 VTAIL.n329 VSUBS 0.014548f
C418 VTAIL.n330 VSUBS 0.032476f
C419 VTAIL.n331 VSUBS 0.032476f
C420 VTAIL.n332 VSUBS 0.014548f
C421 VTAIL.n333 VSUBS 0.01374f
C422 VTAIL.n334 VSUBS 0.025569f
C423 VTAIL.n335 VSUBS 0.025569f
C424 VTAIL.n336 VSUBS 0.01374f
C425 VTAIL.n337 VSUBS 0.014144f
C426 VTAIL.n338 VSUBS 0.014144f
C427 VTAIL.n339 VSUBS 0.032476f
C428 VTAIL.n340 VSUBS 0.032476f
C429 VTAIL.n341 VSUBS 0.014548f
C430 VTAIL.n342 VSUBS 0.01374f
C431 VTAIL.n343 VSUBS 0.025569f
C432 VTAIL.n344 VSUBS 0.025569f
C433 VTAIL.n345 VSUBS 0.01374f
C434 VTAIL.n346 VSUBS 0.014548f
C435 VTAIL.n347 VSUBS 0.032476f
C436 VTAIL.n348 VSUBS 0.077517f
C437 VTAIL.n349 VSUBS 0.014548f
C438 VTAIL.n350 VSUBS 0.01374f
C439 VTAIL.n351 VSUBS 0.061197f
C440 VTAIL.n352 VSUBS 0.038997f
C441 VTAIL.n353 VSUBS 0.131335f
C442 VTAIL.t14 VSUBS 0.217006f
C443 VTAIL.t10 VSUBS 0.217006f
C444 VTAIL.n354 VSUBS 1.53662f
C445 VTAIL.n355 VSUBS 0.697742f
C446 VTAIL.n356 VSUBS 0.027771f
C447 VTAIL.n357 VSUBS 0.025569f
C448 VTAIL.n358 VSUBS 0.01374f
C449 VTAIL.n359 VSUBS 0.032476f
C450 VTAIL.n360 VSUBS 0.014548f
C451 VTAIL.n361 VSUBS 0.025569f
C452 VTAIL.n362 VSUBS 0.01374f
C453 VTAIL.n363 VSUBS 0.032476f
C454 VTAIL.n364 VSUBS 0.014548f
C455 VTAIL.n365 VSUBS 0.025569f
C456 VTAIL.n366 VSUBS 0.01374f
C457 VTAIL.n367 VSUBS 0.032476f
C458 VTAIL.n368 VSUBS 0.032476f
C459 VTAIL.n369 VSUBS 0.014548f
C460 VTAIL.n370 VSUBS 0.025569f
C461 VTAIL.n371 VSUBS 0.01374f
C462 VTAIL.n372 VSUBS 0.032476f
C463 VTAIL.n373 VSUBS 0.014548f
C464 VTAIL.n374 VSUBS 0.186813f
C465 VTAIL.t12 VSUBS 0.069883f
C466 VTAIL.n375 VSUBS 0.024357f
C467 VTAIL.n376 VSUBS 0.02443f
C468 VTAIL.n377 VSUBS 0.01374f
C469 VTAIL.n378 VSUBS 1.1151f
C470 VTAIL.n379 VSUBS 0.025569f
C471 VTAIL.n380 VSUBS 0.01374f
C472 VTAIL.n381 VSUBS 0.014548f
C473 VTAIL.n382 VSUBS 0.032476f
C474 VTAIL.n383 VSUBS 0.032476f
C475 VTAIL.n384 VSUBS 0.014548f
C476 VTAIL.n385 VSUBS 0.01374f
C477 VTAIL.n386 VSUBS 0.025569f
C478 VTAIL.n387 VSUBS 0.025569f
C479 VTAIL.n388 VSUBS 0.01374f
C480 VTAIL.n389 VSUBS 0.014548f
C481 VTAIL.n390 VSUBS 0.032476f
C482 VTAIL.n391 VSUBS 0.032476f
C483 VTAIL.n392 VSUBS 0.014548f
C484 VTAIL.n393 VSUBS 0.01374f
C485 VTAIL.n394 VSUBS 0.025569f
C486 VTAIL.n395 VSUBS 0.025569f
C487 VTAIL.n396 VSUBS 0.01374f
C488 VTAIL.n397 VSUBS 0.014144f
C489 VTAIL.n398 VSUBS 0.014144f
C490 VTAIL.n399 VSUBS 0.032476f
C491 VTAIL.n400 VSUBS 0.032476f
C492 VTAIL.n401 VSUBS 0.014548f
C493 VTAIL.n402 VSUBS 0.01374f
C494 VTAIL.n403 VSUBS 0.025569f
C495 VTAIL.n404 VSUBS 0.025569f
C496 VTAIL.n405 VSUBS 0.01374f
C497 VTAIL.n406 VSUBS 0.014548f
C498 VTAIL.n407 VSUBS 0.032476f
C499 VTAIL.n408 VSUBS 0.077517f
C500 VTAIL.n409 VSUBS 0.014548f
C501 VTAIL.n410 VSUBS 0.01374f
C502 VTAIL.n411 VSUBS 0.061197f
C503 VTAIL.n412 VSUBS 0.038997f
C504 VTAIL.n413 VSUBS 1.27236f
C505 VTAIL.n414 VSUBS 0.027771f
C506 VTAIL.n415 VSUBS 0.025569f
C507 VTAIL.n416 VSUBS 0.01374f
C508 VTAIL.n417 VSUBS 0.032476f
C509 VTAIL.n418 VSUBS 0.014548f
C510 VTAIL.n419 VSUBS 0.025569f
C511 VTAIL.n420 VSUBS 0.01374f
C512 VTAIL.n421 VSUBS 0.032476f
C513 VTAIL.n422 VSUBS 0.014548f
C514 VTAIL.n423 VSUBS 0.025569f
C515 VTAIL.n424 VSUBS 0.01374f
C516 VTAIL.n425 VSUBS 0.032476f
C517 VTAIL.n426 VSUBS 0.014548f
C518 VTAIL.n427 VSUBS 0.025569f
C519 VTAIL.n428 VSUBS 0.01374f
C520 VTAIL.n429 VSUBS 0.032476f
C521 VTAIL.n430 VSUBS 0.014548f
C522 VTAIL.n431 VSUBS 0.186813f
C523 VTAIL.t15 VSUBS 0.069883f
C524 VTAIL.n432 VSUBS 0.024357f
C525 VTAIL.n433 VSUBS 0.02443f
C526 VTAIL.n434 VSUBS 0.01374f
C527 VTAIL.n435 VSUBS 1.1151f
C528 VTAIL.n436 VSUBS 0.025569f
C529 VTAIL.n437 VSUBS 0.01374f
C530 VTAIL.n438 VSUBS 0.014548f
C531 VTAIL.n439 VSUBS 0.032476f
C532 VTAIL.n440 VSUBS 0.032476f
C533 VTAIL.n441 VSUBS 0.014548f
C534 VTAIL.n442 VSUBS 0.01374f
C535 VTAIL.n443 VSUBS 0.025569f
C536 VTAIL.n444 VSUBS 0.025569f
C537 VTAIL.n445 VSUBS 0.01374f
C538 VTAIL.n446 VSUBS 0.014548f
C539 VTAIL.n447 VSUBS 0.032476f
C540 VTAIL.n448 VSUBS 0.032476f
C541 VTAIL.n449 VSUBS 0.032476f
C542 VTAIL.n450 VSUBS 0.014548f
C543 VTAIL.n451 VSUBS 0.01374f
C544 VTAIL.n452 VSUBS 0.025569f
C545 VTAIL.n453 VSUBS 0.025569f
C546 VTAIL.n454 VSUBS 0.01374f
C547 VTAIL.n455 VSUBS 0.014144f
C548 VTAIL.n456 VSUBS 0.014144f
C549 VTAIL.n457 VSUBS 0.032476f
C550 VTAIL.n458 VSUBS 0.032476f
C551 VTAIL.n459 VSUBS 0.014548f
C552 VTAIL.n460 VSUBS 0.01374f
C553 VTAIL.n461 VSUBS 0.025569f
C554 VTAIL.n462 VSUBS 0.025569f
C555 VTAIL.n463 VSUBS 0.01374f
C556 VTAIL.n464 VSUBS 0.014548f
C557 VTAIL.n465 VSUBS 0.032476f
C558 VTAIL.n466 VSUBS 0.077517f
C559 VTAIL.n467 VSUBS 0.014548f
C560 VTAIL.n468 VSUBS 0.01374f
C561 VTAIL.n469 VSUBS 0.061197f
C562 VTAIL.n470 VSUBS 0.038997f
C563 VTAIL.n471 VSUBS 1.26757f
C564 VP.n0 VSUBS 0.095277f
C565 VP.t5 VSUBS 1.14168f
C566 VP.n1 VSUBS 0.466249f
C567 VP.n2 VSUBS 0.285907f
C568 VP.t2 VSUBS 1.14168f
C569 VP.t6 VSUBS 1.14168f
C570 VP.t7 VSUBS 1.14168f
C571 VP.t1 VSUBS 1.16741f
C572 VP.n3 VSUBS 0.442304f
C573 VP.n4 VSUBS 0.47923f
C574 VP.n5 VSUBS 0.47923f
C575 VP.n6 VSUBS 0.466249f
C576 VP.n7 VSUBS 2.27957f
C577 VP.n8 VSUBS 2.32967f
C578 VP.n9 VSUBS 0.095277f
C579 VP.t4 VSUBS 1.14168f
C580 VP.n10 VSUBS 0.47923f
C581 VP.t3 VSUBS 1.14168f
C582 VP.n11 VSUBS 0.47923f
C583 VP.t0 VSUBS 1.14168f
C584 VP.n12 VSUBS 0.466249f
C585 VP.n13 VSUBS 0.063456f
C586 B.n0 VSUBS 0.007412f
C587 B.n1 VSUBS 0.007412f
C588 B.n2 VSUBS 0.010962f
C589 B.n3 VSUBS 0.0084f
C590 B.n4 VSUBS 0.0084f
C591 B.n5 VSUBS 0.0084f
C592 B.n6 VSUBS 0.0084f
C593 B.n7 VSUBS 0.0084f
C594 B.n8 VSUBS 0.0084f
C595 B.n9 VSUBS 0.0084f
C596 B.n10 VSUBS 0.0084f
C597 B.n11 VSUBS 0.0084f
C598 B.n12 VSUBS 0.0084f
C599 B.n13 VSUBS 0.020813f
C600 B.n14 VSUBS 0.0084f
C601 B.n15 VSUBS 0.0084f
C602 B.n16 VSUBS 0.0084f
C603 B.n17 VSUBS 0.0084f
C604 B.n18 VSUBS 0.0084f
C605 B.n19 VSUBS 0.0084f
C606 B.n20 VSUBS 0.0084f
C607 B.n21 VSUBS 0.0084f
C608 B.n22 VSUBS 0.0084f
C609 B.n23 VSUBS 0.0084f
C610 B.n24 VSUBS 0.0084f
C611 B.n25 VSUBS 0.0084f
C612 B.n26 VSUBS 0.0084f
C613 B.n27 VSUBS 0.0084f
C614 B.n28 VSUBS 0.0084f
C615 B.n29 VSUBS 0.0084f
C616 B.n30 VSUBS 0.0084f
C617 B.n31 VSUBS 0.0084f
C618 B.t1 VSUBS 0.220102f
C619 B.t2 VSUBS 0.233334f
C620 B.t0 VSUBS 0.346175f
C621 B.n32 VSUBS 0.336555f
C622 B.n33 VSUBS 0.270972f
C623 B.n34 VSUBS 0.019462f
C624 B.n35 VSUBS 0.0084f
C625 B.n36 VSUBS 0.0084f
C626 B.n37 VSUBS 0.0084f
C627 B.n38 VSUBS 0.0084f
C628 B.n39 VSUBS 0.0084f
C629 B.t7 VSUBS 0.220105f
C630 B.t8 VSUBS 0.233338f
C631 B.t6 VSUBS 0.346175f
C632 B.n40 VSUBS 0.336552f
C633 B.n41 VSUBS 0.270969f
C634 B.n42 VSUBS 0.0084f
C635 B.n43 VSUBS 0.0084f
C636 B.n44 VSUBS 0.0084f
C637 B.n45 VSUBS 0.0084f
C638 B.n46 VSUBS 0.0084f
C639 B.n47 VSUBS 0.0084f
C640 B.n48 VSUBS 0.0084f
C641 B.n49 VSUBS 0.0084f
C642 B.n50 VSUBS 0.0084f
C643 B.n51 VSUBS 0.0084f
C644 B.n52 VSUBS 0.0084f
C645 B.n53 VSUBS 0.0084f
C646 B.n54 VSUBS 0.0084f
C647 B.n55 VSUBS 0.0084f
C648 B.n56 VSUBS 0.0084f
C649 B.n57 VSUBS 0.0084f
C650 B.n58 VSUBS 0.0084f
C651 B.n59 VSUBS 0.0084f
C652 B.n60 VSUBS 0.020199f
C653 B.n61 VSUBS 0.0084f
C654 B.n62 VSUBS 0.0084f
C655 B.n63 VSUBS 0.0084f
C656 B.n64 VSUBS 0.0084f
C657 B.n65 VSUBS 0.0084f
C658 B.n66 VSUBS 0.0084f
C659 B.n67 VSUBS 0.0084f
C660 B.n68 VSUBS 0.0084f
C661 B.n69 VSUBS 0.0084f
C662 B.n70 VSUBS 0.0084f
C663 B.n71 VSUBS 0.0084f
C664 B.n72 VSUBS 0.0084f
C665 B.n73 VSUBS 0.0084f
C666 B.n74 VSUBS 0.0084f
C667 B.n75 VSUBS 0.0084f
C668 B.n76 VSUBS 0.0084f
C669 B.n77 VSUBS 0.0084f
C670 B.n78 VSUBS 0.0084f
C671 B.n79 VSUBS 0.0084f
C672 B.n80 VSUBS 0.0084f
C673 B.n81 VSUBS 0.0084f
C674 B.n82 VSUBS 0.0084f
C675 B.n83 VSUBS 0.020813f
C676 B.n84 VSUBS 0.0084f
C677 B.n85 VSUBS 0.0084f
C678 B.n86 VSUBS 0.0084f
C679 B.n87 VSUBS 0.0084f
C680 B.n88 VSUBS 0.0084f
C681 B.n89 VSUBS 0.0084f
C682 B.n90 VSUBS 0.0084f
C683 B.n91 VSUBS 0.0084f
C684 B.n92 VSUBS 0.0084f
C685 B.n93 VSUBS 0.0084f
C686 B.n94 VSUBS 0.0084f
C687 B.n95 VSUBS 0.0084f
C688 B.n96 VSUBS 0.0084f
C689 B.n97 VSUBS 0.0084f
C690 B.n98 VSUBS 0.0084f
C691 B.n99 VSUBS 0.0084f
C692 B.n100 VSUBS 0.0084f
C693 B.n101 VSUBS 0.0084f
C694 B.t11 VSUBS 0.220105f
C695 B.t10 VSUBS 0.233338f
C696 B.t9 VSUBS 0.346175f
C697 B.n102 VSUBS 0.336552f
C698 B.n103 VSUBS 0.270969f
C699 B.n104 VSUBS 0.019462f
C700 B.n105 VSUBS 0.0084f
C701 B.n106 VSUBS 0.0084f
C702 B.n107 VSUBS 0.0084f
C703 B.n108 VSUBS 0.0084f
C704 B.n109 VSUBS 0.0084f
C705 B.t5 VSUBS 0.220102f
C706 B.t4 VSUBS 0.233334f
C707 B.t3 VSUBS 0.346175f
C708 B.n110 VSUBS 0.336555f
C709 B.n111 VSUBS 0.270972f
C710 B.n112 VSUBS 0.0084f
C711 B.n113 VSUBS 0.0084f
C712 B.n114 VSUBS 0.0084f
C713 B.n115 VSUBS 0.0084f
C714 B.n116 VSUBS 0.0084f
C715 B.n117 VSUBS 0.0084f
C716 B.n118 VSUBS 0.0084f
C717 B.n119 VSUBS 0.0084f
C718 B.n120 VSUBS 0.0084f
C719 B.n121 VSUBS 0.0084f
C720 B.n122 VSUBS 0.0084f
C721 B.n123 VSUBS 0.0084f
C722 B.n124 VSUBS 0.0084f
C723 B.n125 VSUBS 0.0084f
C724 B.n126 VSUBS 0.0084f
C725 B.n127 VSUBS 0.0084f
C726 B.n128 VSUBS 0.0084f
C727 B.n129 VSUBS 0.0084f
C728 B.n130 VSUBS 0.020199f
C729 B.n131 VSUBS 0.0084f
C730 B.n132 VSUBS 0.0084f
C731 B.n133 VSUBS 0.0084f
C732 B.n134 VSUBS 0.0084f
C733 B.n135 VSUBS 0.0084f
C734 B.n136 VSUBS 0.0084f
C735 B.n137 VSUBS 0.0084f
C736 B.n138 VSUBS 0.0084f
C737 B.n139 VSUBS 0.0084f
C738 B.n140 VSUBS 0.0084f
C739 B.n141 VSUBS 0.0084f
C740 B.n142 VSUBS 0.0084f
C741 B.n143 VSUBS 0.0084f
C742 B.n144 VSUBS 0.0084f
C743 B.n145 VSUBS 0.0084f
C744 B.n146 VSUBS 0.0084f
C745 B.n147 VSUBS 0.0084f
C746 B.n148 VSUBS 0.0084f
C747 B.n149 VSUBS 0.0084f
C748 B.n150 VSUBS 0.0084f
C749 B.n151 VSUBS 0.0084f
C750 B.n152 VSUBS 0.0084f
C751 B.n153 VSUBS 0.0084f
C752 B.n154 VSUBS 0.0084f
C753 B.n155 VSUBS 0.0084f
C754 B.n156 VSUBS 0.0084f
C755 B.n157 VSUBS 0.0084f
C756 B.n158 VSUBS 0.0084f
C757 B.n159 VSUBS 0.0084f
C758 B.n160 VSUBS 0.0084f
C759 B.n161 VSUBS 0.0084f
C760 B.n162 VSUBS 0.0084f
C761 B.n163 VSUBS 0.0084f
C762 B.n164 VSUBS 0.0084f
C763 B.n165 VSUBS 0.0084f
C764 B.n166 VSUBS 0.0084f
C765 B.n167 VSUBS 0.0084f
C766 B.n168 VSUBS 0.0084f
C767 B.n169 VSUBS 0.0084f
C768 B.n170 VSUBS 0.0084f
C769 B.n171 VSUBS 0.020199f
C770 B.n172 VSUBS 0.020813f
C771 B.n173 VSUBS 0.020813f
C772 B.n174 VSUBS 0.0084f
C773 B.n175 VSUBS 0.0084f
C774 B.n176 VSUBS 0.0084f
C775 B.n177 VSUBS 0.0084f
C776 B.n178 VSUBS 0.0084f
C777 B.n179 VSUBS 0.0084f
C778 B.n180 VSUBS 0.0084f
C779 B.n181 VSUBS 0.0084f
C780 B.n182 VSUBS 0.0084f
C781 B.n183 VSUBS 0.0084f
C782 B.n184 VSUBS 0.0084f
C783 B.n185 VSUBS 0.0084f
C784 B.n186 VSUBS 0.0084f
C785 B.n187 VSUBS 0.0084f
C786 B.n188 VSUBS 0.0084f
C787 B.n189 VSUBS 0.0084f
C788 B.n190 VSUBS 0.0084f
C789 B.n191 VSUBS 0.0084f
C790 B.n192 VSUBS 0.0084f
C791 B.n193 VSUBS 0.0084f
C792 B.n194 VSUBS 0.0084f
C793 B.n195 VSUBS 0.0084f
C794 B.n196 VSUBS 0.0084f
C795 B.n197 VSUBS 0.0084f
C796 B.n198 VSUBS 0.0084f
C797 B.n199 VSUBS 0.0084f
C798 B.n200 VSUBS 0.0084f
C799 B.n201 VSUBS 0.0084f
C800 B.n202 VSUBS 0.0084f
C801 B.n203 VSUBS 0.0084f
C802 B.n204 VSUBS 0.0084f
C803 B.n205 VSUBS 0.0084f
C804 B.n206 VSUBS 0.0084f
C805 B.n207 VSUBS 0.0084f
C806 B.n208 VSUBS 0.0084f
C807 B.n209 VSUBS 0.0084f
C808 B.n210 VSUBS 0.0084f
C809 B.n211 VSUBS 0.0084f
C810 B.n212 VSUBS 0.0084f
C811 B.n213 VSUBS 0.0084f
C812 B.n214 VSUBS 0.0084f
C813 B.n215 VSUBS 0.0084f
C814 B.n216 VSUBS 0.0084f
C815 B.n217 VSUBS 0.0084f
C816 B.n218 VSUBS 0.0084f
C817 B.n219 VSUBS 0.0084f
C818 B.n220 VSUBS 0.0084f
C819 B.n221 VSUBS 0.0084f
C820 B.n222 VSUBS 0.0084f
C821 B.n223 VSUBS 0.0084f
C822 B.n224 VSUBS 0.0084f
C823 B.n225 VSUBS 0.0084f
C824 B.n226 VSUBS 0.0084f
C825 B.n227 VSUBS 0.0084f
C826 B.n228 VSUBS 0.005806f
C827 B.n229 VSUBS 0.019462f
C828 B.n230 VSUBS 0.006794f
C829 B.n231 VSUBS 0.0084f
C830 B.n232 VSUBS 0.0084f
C831 B.n233 VSUBS 0.0084f
C832 B.n234 VSUBS 0.0084f
C833 B.n235 VSUBS 0.0084f
C834 B.n236 VSUBS 0.0084f
C835 B.n237 VSUBS 0.0084f
C836 B.n238 VSUBS 0.0084f
C837 B.n239 VSUBS 0.0084f
C838 B.n240 VSUBS 0.0084f
C839 B.n241 VSUBS 0.0084f
C840 B.n242 VSUBS 0.006794f
C841 B.n243 VSUBS 0.0084f
C842 B.n244 VSUBS 0.0084f
C843 B.n245 VSUBS 0.005806f
C844 B.n246 VSUBS 0.0084f
C845 B.n247 VSUBS 0.0084f
C846 B.n248 VSUBS 0.0084f
C847 B.n249 VSUBS 0.0084f
C848 B.n250 VSUBS 0.0084f
C849 B.n251 VSUBS 0.0084f
C850 B.n252 VSUBS 0.0084f
C851 B.n253 VSUBS 0.0084f
C852 B.n254 VSUBS 0.0084f
C853 B.n255 VSUBS 0.0084f
C854 B.n256 VSUBS 0.0084f
C855 B.n257 VSUBS 0.0084f
C856 B.n258 VSUBS 0.0084f
C857 B.n259 VSUBS 0.0084f
C858 B.n260 VSUBS 0.0084f
C859 B.n261 VSUBS 0.0084f
C860 B.n262 VSUBS 0.0084f
C861 B.n263 VSUBS 0.0084f
C862 B.n264 VSUBS 0.0084f
C863 B.n265 VSUBS 0.0084f
C864 B.n266 VSUBS 0.0084f
C865 B.n267 VSUBS 0.0084f
C866 B.n268 VSUBS 0.0084f
C867 B.n269 VSUBS 0.0084f
C868 B.n270 VSUBS 0.0084f
C869 B.n271 VSUBS 0.0084f
C870 B.n272 VSUBS 0.0084f
C871 B.n273 VSUBS 0.0084f
C872 B.n274 VSUBS 0.0084f
C873 B.n275 VSUBS 0.0084f
C874 B.n276 VSUBS 0.0084f
C875 B.n277 VSUBS 0.0084f
C876 B.n278 VSUBS 0.0084f
C877 B.n279 VSUBS 0.0084f
C878 B.n280 VSUBS 0.0084f
C879 B.n281 VSUBS 0.0084f
C880 B.n282 VSUBS 0.0084f
C881 B.n283 VSUBS 0.0084f
C882 B.n284 VSUBS 0.0084f
C883 B.n285 VSUBS 0.0084f
C884 B.n286 VSUBS 0.0084f
C885 B.n287 VSUBS 0.0084f
C886 B.n288 VSUBS 0.0084f
C887 B.n289 VSUBS 0.0084f
C888 B.n290 VSUBS 0.0084f
C889 B.n291 VSUBS 0.0084f
C890 B.n292 VSUBS 0.0084f
C891 B.n293 VSUBS 0.0084f
C892 B.n294 VSUBS 0.0084f
C893 B.n295 VSUBS 0.0084f
C894 B.n296 VSUBS 0.0084f
C895 B.n297 VSUBS 0.0084f
C896 B.n298 VSUBS 0.0084f
C897 B.n299 VSUBS 0.0084f
C898 B.n300 VSUBS 0.019881f
C899 B.n301 VSUBS 0.021131f
C900 B.n302 VSUBS 0.020199f
C901 B.n303 VSUBS 0.0084f
C902 B.n304 VSUBS 0.0084f
C903 B.n305 VSUBS 0.0084f
C904 B.n306 VSUBS 0.0084f
C905 B.n307 VSUBS 0.0084f
C906 B.n308 VSUBS 0.0084f
C907 B.n309 VSUBS 0.0084f
C908 B.n310 VSUBS 0.0084f
C909 B.n311 VSUBS 0.0084f
C910 B.n312 VSUBS 0.0084f
C911 B.n313 VSUBS 0.0084f
C912 B.n314 VSUBS 0.0084f
C913 B.n315 VSUBS 0.0084f
C914 B.n316 VSUBS 0.0084f
C915 B.n317 VSUBS 0.0084f
C916 B.n318 VSUBS 0.0084f
C917 B.n319 VSUBS 0.0084f
C918 B.n320 VSUBS 0.0084f
C919 B.n321 VSUBS 0.0084f
C920 B.n322 VSUBS 0.0084f
C921 B.n323 VSUBS 0.0084f
C922 B.n324 VSUBS 0.0084f
C923 B.n325 VSUBS 0.0084f
C924 B.n326 VSUBS 0.0084f
C925 B.n327 VSUBS 0.0084f
C926 B.n328 VSUBS 0.0084f
C927 B.n329 VSUBS 0.0084f
C928 B.n330 VSUBS 0.0084f
C929 B.n331 VSUBS 0.0084f
C930 B.n332 VSUBS 0.0084f
C931 B.n333 VSUBS 0.0084f
C932 B.n334 VSUBS 0.0084f
C933 B.n335 VSUBS 0.0084f
C934 B.n336 VSUBS 0.0084f
C935 B.n337 VSUBS 0.0084f
C936 B.n338 VSUBS 0.0084f
C937 B.n339 VSUBS 0.0084f
C938 B.n340 VSUBS 0.0084f
C939 B.n341 VSUBS 0.0084f
C940 B.n342 VSUBS 0.0084f
C941 B.n343 VSUBS 0.0084f
C942 B.n344 VSUBS 0.0084f
C943 B.n345 VSUBS 0.0084f
C944 B.n346 VSUBS 0.0084f
C945 B.n347 VSUBS 0.0084f
C946 B.n348 VSUBS 0.0084f
C947 B.n349 VSUBS 0.0084f
C948 B.n350 VSUBS 0.0084f
C949 B.n351 VSUBS 0.0084f
C950 B.n352 VSUBS 0.0084f
C951 B.n353 VSUBS 0.0084f
C952 B.n354 VSUBS 0.0084f
C953 B.n355 VSUBS 0.0084f
C954 B.n356 VSUBS 0.0084f
C955 B.n357 VSUBS 0.0084f
C956 B.n358 VSUBS 0.0084f
C957 B.n359 VSUBS 0.0084f
C958 B.n360 VSUBS 0.0084f
C959 B.n361 VSUBS 0.0084f
C960 B.n362 VSUBS 0.0084f
C961 B.n363 VSUBS 0.0084f
C962 B.n364 VSUBS 0.0084f
C963 B.n365 VSUBS 0.0084f
C964 B.n366 VSUBS 0.0084f
C965 B.n367 VSUBS 0.0084f
C966 B.n368 VSUBS 0.0084f
C967 B.n369 VSUBS 0.020199f
C968 B.n370 VSUBS 0.020813f
C969 B.n371 VSUBS 0.020813f
C970 B.n372 VSUBS 0.0084f
C971 B.n373 VSUBS 0.0084f
C972 B.n374 VSUBS 0.0084f
C973 B.n375 VSUBS 0.0084f
C974 B.n376 VSUBS 0.0084f
C975 B.n377 VSUBS 0.0084f
C976 B.n378 VSUBS 0.0084f
C977 B.n379 VSUBS 0.0084f
C978 B.n380 VSUBS 0.0084f
C979 B.n381 VSUBS 0.0084f
C980 B.n382 VSUBS 0.0084f
C981 B.n383 VSUBS 0.0084f
C982 B.n384 VSUBS 0.0084f
C983 B.n385 VSUBS 0.0084f
C984 B.n386 VSUBS 0.0084f
C985 B.n387 VSUBS 0.0084f
C986 B.n388 VSUBS 0.0084f
C987 B.n389 VSUBS 0.0084f
C988 B.n390 VSUBS 0.0084f
C989 B.n391 VSUBS 0.0084f
C990 B.n392 VSUBS 0.0084f
C991 B.n393 VSUBS 0.0084f
C992 B.n394 VSUBS 0.0084f
C993 B.n395 VSUBS 0.0084f
C994 B.n396 VSUBS 0.0084f
C995 B.n397 VSUBS 0.0084f
C996 B.n398 VSUBS 0.0084f
C997 B.n399 VSUBS 0.0084f
C998 B.n400 VSUBS 0.0084f
C999 B.n401 VSUBS 0.0084f
C1000 B.n402 VSUBS 0.0084f
C1001 B.n403 VSUBS 0.0084f
C1002 B.n404 VSUBS 0.0084f
C1003 B.n405 VSUBS 0.0084f
C1004 B.n406 VSUBS 0.0084f
C1005 B.n407 VSUBS 0.0084f
C1006 B.n408 VSUBS 0.0084f
C1007 B.n409 VSUBS 0.0084f
C1008 B.n410 VSUBS 0.0084f
C1009 B.n411 VSUBS 0.0084f
C1010 B.n412 VSUBS 0.0084f
C1011 B.n413 VSUBS 0.0084f
C1012 B.n414 VSUBS 0.0084f
C1013 B.n415 VSUBS 0.0084f
C1014 B.n416 VSUBS 0.0084f
C1015 B.n417 VSUBS 0.0084f
C1016 B.n418 VSUBS 0.0084f
C1017 B.n419 VSUBS 0.0084f
C1018 B.n420 VSUBS 0.0084f
C1019 B.n421 VSUBS 0.0084f
C1020 B.n422 VSUBS 0.0084f
C1021 B.n423 VSUBS 0.0084f
C1022 B.n424 VSUBS 0.0084f
C1023 B.n425 VSUBS 0.0084f
C1024 B.n426 VSUBS 0.005806f
C1025 B.n427 VSUBS 0.019462f
C1026 B.n428 VSUBS 0.006794f
C1027 B.n429 VSUBS 0.0084f
C1028 B.n430 VSUBS 0.0084f
C1029 B.n431 VSUBS 0.0084f
C1030 B.n432 VSUBS 0.0084f
C1031 B.n433 VSUBS 0.0084f
C1032 B.n434 VSUBS 0.0084f
C1033 B.n435 VSUBS 0.0084f
C1034 B.n436 VSUBS 0.0084f
C1035 B.n437 VSUBS 0.0084f
C1036 B.n438 VSUBS 0.0084f
C1037 B.n439 VSUBS 0.0084f
C1038 B.n440 VSUBS 0.006794f
C1039 B.n441 VSUBS 0.0084f
C1040 B.n442 VSUBS 0.0084f
C1041 B.n443 VSUBS 0.005806f
C1042 B.n444 VSUBS 0.0084f
C1043 B.n445 VSUBS 0.0084f
C1044 B.n446 VSUBS 0.0084f
C1045 B.n447 VSUBS 0.0084f
C1046 B.n448 VSUBS 0.0084f
C1047 B.n449 VSUBS 0.0084f
C1048 B.n450 VSUBS 0.0084f
C1049 B.n451 VSUBS 0.0084f
C1050 B.n452 VSUBS 0.0084f
C1051 B.n453 VSUBS 0.0084f
C1052 B.n454 VSUBS 0.0084f
C1053 B.n455 VSUBS 0.0084f
C1054 B.n456 VSUBS 0.0084f
C1055 B.n457 VSUBS 0.0084f
C1056 B.n458 VSUBS 0.0084f
C1057 B.n459 VSUBS 0.0084f
C1058 B.n460 VSUBS 0.0084f
C1059 B.n461 VSUBS 0.0084f
C1060 B.n462 VSUBS 0.0084f
C1061 B.n463 VSUBS 0.0084f
C1062 B.n464 VSUBS 0.0084f
C1063 B.n465 VSUBS 0.0084f
C1064 B.n466 VSUBS 0.0084f
C1065 B.n467 VSUBS 0.0084f
C1066 B.n468 VSUBS 0.0084f
C1067 B.n469 VSUBS 0.0084f
C1068 B.n470 VSUBS 0.0084f
C1069 B.n471 VSUBS 0.0084f
C1070 B.n472 VSUBS 0.0084f
C1071 B.n473 VSUBS 0.0084f
C1072 B.n474 VSUBS 0.0084f
C1073 B.n475 VSUBS 0.0084f
C1074 B.n476 VSUBS 0.0084f
C1075 B.n477 VSUBS 0.0084f
C1076 B.n478 VSUBS 0.0084f
C1077 B.n479 VSUBS 0.0084f
C1078 B.n480 VSUBS 0.0084f
C1079 B.n481 VSUBS 0.0084f
C1080 B.n482 VSUBS 0.0084f
C1081 B.n483 VSUBS 0.0084f
C1082 B.n484 VSUBS 0.0084f
C1083 B.n485 VSUBS 0.0084f
C1084 B.n486 VSUBS 0.0084f
C1085 B.n487 VSUBS 0.0084f
C1086 B.n488 VSUBS 0.0084f
C1087 B.n489 VSUBS 0.0084f
C1088 B.n490 VSUBS 0.0084f
C1089 B.n491 VSUBS 0.0084f
C1090 B.n492 VSUBS 0.0084f
C1091 B.n493 VSUBS 0.0084f
C1092 B.n494 VSUBS 0.0084f
C1093 B.n495 VSUBS 0.0084f
C1094 B.n496 VSUBS 0.0084f
C1095 B.n497 VSUBS 0.0084f
C1096 B.n498 VSUBS 0.020813f
C1097 B.n499 VSUBS 0.020199f
C1098 B.n500 VSUBS 0.020199f
C1099 B.n501 VSUBS 0.0084f
C1100 B.n502 VSUBS 0.0084f
C1101 B.n503 VSUBS 0.0084f
C1102 B.n504 VSUBS 0.0084f
C1103 B.n505 VSUBS 0.0084f
C1104 B.n506 VSUBS 0.0084f
C1105 B.n507 VSUBS 0.0084f
C1106 B.n508 VSUBS 0.0084f
C1107 B.n509 VSUBS 0.0084f
C1108 B.n510 VSUBS 0.0084f
C1109 B.n511 VSUBS 0.0084f
C1110 B.n512 VSUBS 0.0084f
C1111 B.n513 VSUBS 0.0084f
C1112 B.n514 VSUBS 0.0084f
C1113 B.n515 VSUBS 0.0084f
C1114 B.n516 VSUBS 0.0084f
C1115 B.n517 VSUBS 0.0084f
C1116 B.n518 VSUBS 0.0084f
C1117 B.n519 VSUBS 0.0084f
C1118 B.n520 VSUBS 0.0084f
C1119 B.n521 VSUBS 0.0084f
C1120 B.n522 VSUBS 0.0084f
C1121 B.n523 VSUBS 0.0084f
C1122 B.n524 VSUBS 0.0084f
C1123 B.n525 VSUBS 0.0084f
C1124 B.n526 VSUBS 0.0084f
C1125 B.n527 VSUBS 0.0084f
C1126 B.n528 VSUBS 0.0084f
C1127 B.n529 VSUBS 0.0084f
C1128 B.n530 VSUBS 0.0084f
C1129 B.n531 VSUBS 0.010962f
C1130 B.n532 VSUBS 0.011677f
C1131 B.n533 VSUBS 0.023221f
.ends

