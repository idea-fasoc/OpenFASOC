* NGSPICE file created from diff_pair_sample_0398.ext - technology: sky130A

.subckt diff_pair_sample_0398 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=1.71
X1 VDD1.t9 VP.t0 VTAIL.t13 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X2 VTAIL.t9 VN.t0 VDD2.t9 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X3 VDD2.t8 VN.t1 VTAIL.t3 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X4 B.t8 B.t6 B.t7 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=1.71
X5 B.t5 B.t3 B.t4 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=1.71
X6 VDD2.t7 VN.t2 VTAIL.t8 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=1.71
X7 VDD2.t6 VN.t3 VTAIL.t1 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=1.71
X8 VDD2.t5 VN.t4 VTAIL.t7 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=1.71
X9 VDD1.t8 VP.t1 VTAIL.t14 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=1.71
X10 VTAIL.t6 VN.t5 VDD2.t4 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X11 VDD1.t7 VP.t2 VTAIL.t12 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=4.7229 ps=25 w=12.11 l=1.71
X12 VTAIL.t11 VP.t3 VDD1.t6 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X13 VDD1.t5 VP.t4 VTAIL.t16 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=1.71
X14 VTAIL.t19 VP.t5 VDD1.t4 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X15 VTAIL.t17 VP.t6 VDD1.t3 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X16 VTAIL.t0 VN.t6 VDD2.t3 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X17 B.t2 B.t0 B.t1 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=0 ps=0 w=12.11 l=1.71
X18 VDD1.t2 VP.t7 VTAIL.t18 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X19 VDD1.t1 VP.t8 VTAIL.t15 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=1.71
X20 VDD2.t2 VN.t7 VTAIL.t5 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X21 VTAIL.t2 VN.t8 VDD2.t1 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X22 VTAIL.t10 VP.t9 VDD1.t0 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=1.99815 pd=12.44 as=1.99815 ps=12.44 w=12.11 l=1.71
X23 VDD2.t0 VN.t9 VTAIL.t4 w_n3418_n3390# sky130_fd_pr__pfet_01v8 ad=4.7229 pd=25 as=1.99815 ps=12.44 w=12.11 l=1.71
R0 B.n531 B.n74 585
R1 B.n533 B.n532 585
R2 B.n534 B.n73 585
R3 B.n536 B.n535 585
R4 B.n537 B.n72 585
R5 B.n539 B.n538 585
R6 B.n540 B.n71 585
R7 B.n542 B.n541 585
R8 B.n543 B.n70 585
R9 B.n545 B.n544 585
R10 B.n546 B.n69 585
R11 B.n548 B.n547 585
R12 B.n549 B.n68 585
R13 B.n551 B.n550 585
R14 B.n552 B.n67 585
R15 B.n554 B.n553 585
R16 B.n555 B.n66 585
R17 B.n557 B.n556 585
R18 B.n558 B.n65 585
R19 B.n560 B.n559 585
R20 B.n561 B.n64 585
R21 B.n563 B.n562 585
R22 B.n564 B.n63 585
R23 B.n566 B.n565 585
R24 B.n567 B.n62 585
R25 B.n569 B.n568 585
R26 B.n570 B.n61 585
R27 B.n572 B.n571 585
R28 B.n573 B.n60 585
R29 B.n575 B.n574 585
R30 B.n576 B.n59 585
R31 B.n578 B.n577 585
R32 B.n579 B.n58 585
R33 B.n581 B.n580 585
R34 B.n582 B.n57 585
R35 B.n584 B.n583 585
R36 B.n585 B.n56 585
R37 B.n587 B.n586 585
R38 B.n588 B.n55 585
R39 B.n590 B.n589 585
R40 B.n591 B.n54 585
R41 B.n593 B.n592 585
R42 B.n595 B.n51 585
R43 B.n597 B.n596 585
R44 B.n598 B.n50 585
R45 B.n600 B.n599 585
R46 B.n601 B.n49 585
R47 B.n603 B.n602 585
R48 B.n604 B.n48 585
R49 B.n606 B.n605 585
R50 B.n607 B.n45 585
R51 B.n610 B.n609 585
R52 B.n611 B.n44 585
R53 B.n613 B.n612 585
R54 B.n614 B.n43 585
R55 B.n616 B.n615 585
R56 B.n617 B.n42 585
R57 B.n619 B.n618 585
R58 B.n620 B.n41 585
R59 B.n622 B.n621 585
R60 B.n623 B.n40 585
R61 B.n625 B.n624 585
R62 B.n626 B.n39 585
R63 B.n628 B.n627 585
R64 B.n629 B.n38 585
R65 B.n631 B.n630 585
R66 B.n632 B.n37 585
R67 B.n634 B.n633 585
R68 B.n635 B.n36 585
R69 B.n637 B.n636 585
R70 B.n638 B.n35 585
R71 B.n640 B.n639 585
R72 B.n641 B.n34 585
R73 B.n643 B.n642 585
R74 B.n644 B.n33 585
R75 B.n646 B.n645 585
R76 B.n647 B.n32 585
R77 B.n649 B.n648 585
R78 B.n650 B.n31 585
R79 B.n652 B.n651 585
R80 B.n653 B.n30 585
R81 B.n655 B.n654 585
R82 B.n656 B.n29 585
R83 B.n658 B.n657 585
R84 B.n659 B.n28 585
R85 B.n661 B.n660 585
R86 B.n662 B.n27 585
R87 B.n664 B.n663 585
R88 B.n665 B.n26 585
R89 B.n667 B.n666 585
R90 B.n668 B.n25 585
R91 B.n670 B.n669 585
R92 B.n671 B.n24 585
R93 B.n530 B.n529 585
R94 B.n528 B.n75 585
R95 B.n527 B.n526 585
R96 B.n525 B.n76 585
R97 B.n524 B.n523 585
R98 B.n522 B.n77 585
R99 B.n521 B.n520 585
R100 B.n519 B.n78 585
R101 B.n518 B.n517 585
R102 B.n516 B.n79 585
R103 B.n515 B.n514 585
R104 B.n513 B.n80 585
R105 B.n512 B.n511 585
R106 B.n510 B.n81 585
R107 B.n509 B.n508 585
R108 B.n507 B.n82 585
R109 B.n506 B.n505 585
R110 B.n504 B.n83 585
R111 B.n503 B.n502 585
R112 B.n501 B.n84 585
R113 B.n500 B.n499 585
R114 B.n498 B.n85 585
R115 B.n497 B.n496 585
R116 B.n495 B.n86 585
R117 B.n494 B.n493 585
R118 B.n492 B.n87 585
R119 B.n491 B.n490 585
R120 B.n489 B.n88 585
R121 B.n488 B.n487 585
R122 B.n486 B.n89 585
R123 B.n485 B.n484 585
R124 B.n483 B.n90 585
R125 B.n482 B.n481 585
R126 B.n480 B.n91 585
R127 B.n479 B.n478 585
R128 B.n477 B.n92 585
R129 B.n476 B.n475 585
R130 B.n474 B.n93 585
R131 B.n473 B.n472 585
R132 B.n471 B.n94 585
R133 B.n470 B.n469 585
R134 B.n468 B.n95 585
R135 B.n467 B.n466 585
R136 B.n465 B.n96 585
R137 B.n464 B.n463 585
R138 B.n462 B.n97 585
R139 B.n461 B.n460 585
R140 B.n459 B.n98 585
R141 B.n458 B.n457 585
R142 B.n456 B.n99 585
R143 B.n455 B.n454 585
R144 B.n453 B.n100 585
R145 B.n452 B.n451 585
R146 B.n450 B.n101 585
R147 B.n449 B.n448 585
R148 B.n447 B.n102 585
R149 B.n446 B.n445 585
R150 B.n444 B.n103 585
R151 B.n443 B.n442 585
R152 B.n441 B.n104 585
R153 B.n440 B.n439 585
R154 B.n438 B.n105 585
R155 B.n437 B.n436 585
R156 B.n435 B.n106 585
R157 B.n434 B.n433 585
R158 B.n432 B.n107 585
R159 B.n431 B.n430 585
R160 B.n429 B.n108 585
R161 B.n428 B.n427 585
R162 B.n426 B.n109 585
R163 B.n425 B.n424 585
R164 B.n423 B.n110 585
R165 B.n422 B.n421 585
R166 B.n420 B.n111 585
R167 B.n419 B.n418 585
R168 B.n417 B.n112 585
R169 B.n416 B.n415 585
R170 B.n414 B.n113 585
R171 B.n413 B.n412 585
R172 B.n411 B.n114 585
R173 B.n410 B.n409 585
R174 B.n408 B.n115 585
R175 B.n407 B.n406 585
R176 B.n405 B.n116 585
R177 B.n404 B.n403 585
R178 B.n402 B.n117 585
R179 B.n401 B.n400 585
R180 B.n399 B.n118 585
R181 B.n398 B.n397 585
R182 B.n257 B.n256 585
R183 B.n258 B.n169 585
R184 B.n260 B.n259 585
R185 B.n261 B.n168 585
R186 B.n263 B.n262 585
R187 B.n264 B.n167 585
R188 B.n266 B.n265 585
R189 B.n267 B.n166 585
R190 B.n269 B.n268 585
R191 B.n270 B.n165 585
R192 B.n272 B.n271 585
R193 B.n273 B.n164 585
R194 B.n275 B.n274 585
R195 B.n276 B.n163 585
R196 B.n278 B.n277 585
R197 B.n279 B.n162 585
R198 B.n281 B.n280 585
R199 B.n282 B.n161 585
R200 B.n284 B.n283 585
R201 B.n285 B.n160 585
R202 B.n287 B.n286 585
R203 B.n288 B.n159 585
R204 B.n290 B.n289 585
R205 B.n291 B.n158 585
R206 B.n293 B.n292 585
R207 B.n294 B.n157 585
R208 B.n296 B.n295 585
R209 B.n297 B.n156 585
R210 B.n299 B.n298 585
R211 B.n300 B.n155 585
R212 B.n302 B.n301 585
R213 B.n303 B.n154 585
R214 B.n305 B.n304 585
R215 B.n306 B.n153 585
R216 B.n308 B.n307 585
R217 B.n309 B.n152 585
R218 B.n311 B.n310 585
R219 B.n312 B.n151 585
R220 B.n314 B.n313 585
R221 B.n315 B.n150 585
R222 B.n317 B.n316 585
R223 B.n318 B.n147 585
R224 B.n321 B.n320 585
R225 B.n322 B.n146 585
R226 B.n324 B.n323 585
R227 B.n325 B.n145 585
R228 B.n327 B.n326 585
R229 B.n328 B.n144 585
R230 B.n330 B.n329 585
R231 B.n331 B.n143 585
R232 B.n333 B.n332 585
R233 B.n335 B.n334 585
R234 B.n336 B.n139 585
R235 B.n338 B.n337 585
R236 B.n339 B.n138 585
R237 B.n341 B.n340 585
R238 B.n342 B.n137 585
R239 B.n344 B.n343 585
R240 B.n345 B.n136 585
R241 B.n347 B.n346 585
R242 B.n348 B.n135 585
R243 B.n350 B.n349 585
R244 B.n351 B.n134 585
R245 B.n353 B.n352 585
R246 B.n354 B.n133 585
R247 B.n356 B.n355 585
R248 B.n357 B.n132 585
R249 B.n359 B.n358 585
R250 B.n360 B.n131 585
R251 B.n362 B.n361 585
R252 B.n363 B.n130 585
R253 B.n365 B.n364 585
R254 B.n366 B.n129 585
R255 B.n368 B.n367 585
R256 B.n369 B.n128 585
R257 B.n371 B.n370 585
R258 B.n372 B.n127 585
R259 B.n374 B.n373 585
R260 B.n375 B.n126 585
R261 B.n377 B.n376 585
R262 B.n378 B.n125 585
R263 B.n380 B.n379 585
R264 B.n381 B.n124 585
R265 B.n383 B.n382 585
R266 B.n384 B.n123 585
R267 B.n386 B.n385 585
R268 B.n387 B.n122 585
R269 B.n389 B.n388 585
R270 B.n390 B.n121 585
R271 B.n392 B.n391 585
R272 B.n393 B.n120 585
R273 B.n395 B.n394 585
R274 B.n396 B.n119 585
R275 B.n255 B.n170 585
R276 B.n254 B.n253 585
R277 B.n252 B.n171 585
R278 B.n251 B.n250 585
R279 B.n249 B.n172 585
R280 B.n248 B.n247 585
R281 B.n246 B.n173 585
R282 B.n245 B.n244 585
R283 B.n243 B.n174 585
R284 B.n242 B.n241 585
R285 B.n240 B.n175 585
R286 B.n239 B.n238 585
R287 B.n237 B.n176 585
R288 B.n236 B.n235 585
R289 B.n234 B.n177 585
R290 B.n233 B.n232 585
R291 B.n231 B.n178 585
R292 B.n230 B.n229 585
R293 B.n228 B.n179 585
R294 B.n227 B.n226 585
R295 B.n225 B.n180 585
R296 B.n224 B.n223 585
R297 B.n222 B.n181 585
R298 B.n221 B.n220 585
R299 B.n219 B.n182 585
R300 B.n218 B.n217 585
R301 B.n216 B.n183 585
R302 B.n215 B.n214 585
R303 B.n213 B.n184 585
R304 B.n212 B.n211 585
R305 B.n210 B.n185 585
R306 B.n209 B.n208 585
R307 B.n207 B.n186 585
R308 B.n206 B.n205 585
R309 B.n204 B.n187 585
R310 B.n203 B.n202 585
R311 B.n201 B.n188 585
R312 B.n200 B.n199 585
R313 B.n198 B.n189 585
R314 B.n197 B.n196 585
R315 B.n195 B.n190 585
R316 B.n194 B.n193 585
R317 B.n192 B.n191 585
R318 B.n2 B.n0 585
R319 B.n737 B.n1 585
R320 B.n736 B.n735 585
R321 B.n734 B.n3 585
R322 B.n733 B.n732 585
R323 B.n731 B.n4 585
R324 B.n730 B.n729 585
R325 B.n728 B.n5 585
R326 B.n727 B.n726 585
R327 B.n725 B.n6 585
R328 B.n724 B.n723 585
R329 B.n722 B.n7 585
R330 B.n721 B.n720 585
R331 B.n719 B.n8 585
R332 B.n718 B.n717 585
R333 B.n716 B.n9 585
R334 B.n715 B.n714 585
R335 B.n713 B.n10 585
R336 B.n712 B.n711 585
R337 B.n710 B.n11 585
R338 B.n709 B.n708 585
R339 B.n707 B.n12 585
R340 B.n706 B.n705 585
R341 B.n704 B.n13 585
R342 B.n703 B.n702 585
R343 B.n701 B.n14 585
R344 B.n700 B.n699 585
R345 B.n698 B.n15 585
R346 B.n697 B.n696 585
R347 B.n695 B.n16 585
R348 B.n694 B.n693 585
R349 B.n692 B.n17 585
R350 B.n691 B.n690 585
R351 B.n689 B.n18 585
R352 B.n688 B.n687 585
R353 B.n686 B.n19 585
R354 B.n685 B.n684 585
R355 B.n683 B.n20 585
R356 B.n682 B.n681 585
R357 B.n680 B.n21 585
R358 B.n679 B.n678 585
R359 B.n677 B.n22 585
R360 B.n676 B.n675 585
R361 B.n674 B.n23 585
R362 B.n673 B.n672 585
R363 B.n739 B.n738 585
R364 B.n256 B.n255 554.963
R365 B.n672 B.n671 554.963
R366 B.n398 B.n119 554.963
R367 B.n531 B.n530 554.963
R368 B.n140 B.t2 417.228
R369 B.n52 B.t4 417.228
R370 B.n148 B.t11 417.226
R371 B.n46 B.t7 417.226
R372 B.n141 B.t1 377.663
R373 B.n53 B.t5 377.663
R374 B.n149 B.t10 377.663
R375 B.n47 B.t8 377.663
R376 B.n140 B.t0 376.818
R377 B.n148 B.t9 376.818
R378 B.n46 B.t6 376.818
R379 B.n52 B.t3 376.818
R380 B.n255 B.n254 163.367
R381 B.n254 B.n171 163.367
R382 B.n250 B.n171 163.367
R383 B.n250 B.n249 163.367
R384 B.n249 B.n248 163.367
R385 B.n248 B.n173 163.367
R386 B.n244 B.n173 163.367
R387 B.n244 B.n243 163.367
R388 B.n243 B.n242 163.367
R389 B.n242 B.n175 163.367
R390 B.n238 B.n175 163.367
R391 B.n238 B.n237 163.367
R392 B.n237 B.n236 163.367
R393 B.n236 B.n177 163.367
R394 B.n232 B.n177 163.367
R395 B.n232 B.n231 163.367
R396 B.n231 B.n230 163.367
R397 B.n230 B.n179 163.367
R398 B.n226 B.n179 163.367
R399 B.n226 B.n225 163.367
R400 B.n225 B.n224 163.367
R401 B.n224 B.n181 163.367
R402 B.n220 B.n181 163.367
R403 B.n220 B.n219 163.367
R404 B.n219 B.n218 163.367
R405 B.n218 B.n183 163.367
R406 B.n214 B.n183 163.367
R407 B.n214 B.n213 163.367
R408 B.n213 B.n212 163.367
R409 B.n212 B.n185 163.367
R410 B.n208 B.n185 163.367
R411 B.n208 B.n207 163.367
R412 B.n207 B.n206 163.367
R413 B.n206 B.n187 163.367
R414 B.n202 B.n187 163.367
R415 B.n202 B.n201 163.367
R416 B.n201 B.n200 163.367
R417 B.n200 B.n189 163.367
R418 B.n196 B.n189 163.367
R419 B.n196 B.n195 163.367
R420 B.n195 B.n194 163.367
R421 B.n194 B.n191 163.367
R422 B.n191 B.n2 163.367
R423 B.n738 B.n2 163.367
R424 B.n738 B.n737 163.367
R425 B.n737 B.n736 163.367
R426 B.n736 B.n3 163.367
R427 B.n732 B.n3 163.367
R428 B.n732 B.n731 163.367
R429 B.n731 B.n730 163.367
R430 B.n730 B.n5 163.367
R431 B.n726 B.n5 163.367
R432 B.n726 B.n725 163.367
R433 B.n725 B.n724 163.367
R434 B.n724 B.n7 163.367
R435 B.n720 B.n7 163.367
R436 B.n720 B.n719 163.367
R437 B.n719 B.n718 163.367
R438 B.n718 B.n9 163.367
R439 B.n714 B.n9 163.367
R440 B.n714 B.n713 163.367
R441 B.n713 B.n712 163.367
R442 B.n712 B.n11 163.367
R443 B.n708 B.n11 163.367
R444 B.n708 B.n707 163.367
R445 B.n707 B.n706 163.367
R446 B.n706 B.n13 163.367
R447 B.n702 B.n13 163.367
R448 B.n702 B.n701 163.367
R449 B.n701 B.n700 163.367
R450 B.n700 B.n15 163.367
R451 B.n696 B.n15 163.367
R452 B.n696 B.n695 163.367
R453 B.n695 B.n694 163.367
R454 B.n694 B.n17 163.367
R455 B.n690 B.n17 163.367
R456 B.n690 B.n689 163.367
R457 B.n689 B.n688 163.367
R458 B.n688 B.n19 163.367
R459 B.n684 B.n19 163.367
R460 B.n684 B.n683 163.367
R461 B.n683 B.n682 163.367
R462 B.n682 B.n21 163.367
R463 B.n678 B.n21 163.367
R464 B.n678 B.n677 163.367
R465 B.n677 B.n676 163.367
R466 B.n676 B.n23 163.367
R467 B.n672 B.n23 163.367
R468 B.n256 B.n169 163.367
R469 B.n260 B.n169 163.367
R470 B.n261 B.n260 163.367
R471 B.n262 B.n261 163.367
R472 B.n262 B.n167 163.367
R473 B.n266 B.n167 163.367
R474 B.n267 B.n266 163.367
R475 B.n268 B.n267 163.367
R476 B.n268 B.n165 163.367
R477 B.n272 B.n165 163.367
R478 B.n273 B.n272 163.367
R479 B.n274 B.n273 163.367
R480 B.n274 B.n163 163.367
R481 B.n278 B.n163 163.367
R482 B.n279 B.n278 163.367
R483 B.n280 B.n279 163.367
R484 B.n280 B.n161 163.367
R485 B.n284 B.n161 163.367
R486 B.n285 B.n284 163.367
R487 B.n286 B.n285 163.367
R488 B.n286 B.n159 163.367
R489 B.n290 B.n159 163.367
R490 B.n291 B.n290 163.367
R491 B.n292 B.n291 163.367
R492 B.n292 B.n157 163.367
R493 B.n296 B.n157 163.367
R494 B.n297 B.n296 163.367
R495 B.n298 B.n297 163.367
R496 B.n298 B.n155 163.367
R497 B.n302 B.n155 163.367
R498 B.n303 B.n302 163.367
R499 B.n304 B.n303 163.367
R500 B.n304 B.n153 163.367
R501 B.n308 B.n153 163.367
R502 B.n309 B.n308 163.367
R503 B.n310 B.n309 163.367
R504 B.n310 B.n151 163.367
R505 B.n314 B.n151 163.367
R506 B.n315 B.n314 163.367
R507 B.n316 B.n315 163.367
R508 B.n316 B.n147 163.367
R509 B.n321 B.n147 163.367
R510 B.n322 B.n321 163.367
R511 B.n323 B.n322 163.367
R512 B.n323 B.n145 163.367
R513 B.n327 B.n145 163.367
R514 B.n328 B.n327 163.367
R515 B.n329 B.n328 163.367
R516 B.n329 B.n143 163.367
R517 B.n333 B.n143 163.367
R518 B.n334 B.n333 163.367
R519 B.n334 B.n139 163.367
R520 B.n338 B.n139 163.367
R521 B.n339 B.n338 163.367
R522 B.n340 B.n339 163.367
R523 B.n340 B.n137 163.367
R524 B.n344 B.n137 163.367
R525 B.n345 B.n344 163.367
R526 B.n346 B.n345 163.367
R527 B.n346 B.n135 163.367
R528 B.n350 B.n135 163.367
R529 B.n351 B.n350 163.367
R530 B.n352 B.n351 163.367
R531 B.n352 B.n133 163.367
R532 B.n356 B.n133 163.367
R533 B.n357 B.n356 163.367
R534 B.n358 B.n357 163.367
R535 B.n358 B.n131 163.367
R536 B.n362 B.n131 163.367
R537 B.n363 B.n362 163.367
R538 B.n364 B.n363 163.367
R539 B.n364 B.n129 163.367
R540 B.n368 B.n129 163.367
R541 B.n369 B.n368 163.367
R542 B.n370 B.n369 163.367
R543 B.n370 B.n127 163.367
R544 B.n374 B.n127 163.367
R545 B.n375 B.n374 163.367
R546 B.n376 B.n375 163.367
R547 B.n376 B.n125 163.367
R548 B.n380 B.n125 163.367
R549 B.n381 B.n380 163.367
R550 B.n382 B.n381 163.367
R551 B.n382 B.n123 163.367
R552 B.n386 B.n123 163.367
R553 B.n387 B.n386 163.367
R554 B.n388 B.n387 163.367
R555 B.n388 B.n121 163.367
R556 B.n392 B.n121 163.367
R557 B.n393 B.n392 163.367
R558 B.n394 B.n393 163.367
R559 B.n394 B.n119 163.367
R560 B.n399 B.n398 163.367
R561 B.n400 B.n399 163.367
R562 B.n400 B.n117 163.367
R563 B.n404 B.n117 163.367
R564 B.n405 B.n404 163.367
R565 B.n406 B.n405 163.367
R566 B.n406 B.n115 163.367
R567 B.n410 B.n115 163.367
R568 B.n411 B.n410 163.367
R569 B.n412 B.n411 163.367
R570 B.n412 B.n113 163.367
R571 B.n416 B.n113 163.367
R572 B.n417 B.n416 163.367
R573 B.n418 B.n417 163.367
R574 B.n418 B.n111 163.367
R575 B.n422 B.n111 163.367
R576 B.n423 B.n422 163.367
R577 B.n424 B.n423 163.367
R578 B.n424 B.n109 163.367
R579 B.n428 B.n109 163.367
R580 B.n429 B.n428 163.367
R581 B.n430 B.n429 163.367
R582 B.n430 B.n107 163.367
R583 B.n434 B.n107 163.367
R584 B.n435 B.n434 163.367
R585 B.n436 B.n435 163.367
R586 B.n436 B.n105 163.367
R587 B.n440 B.n105 163.367
R588 B.n441 B.n440 163.367
R589 B.n442 B.n441 163.367
R590 B.n442 B.n103 163.367
R591 B.n446 B.n103 163.367
R592 B.n447 B.n446 163.367
R593 B.n448 B.n447 163.367
R594 B.n448 B.n101 163.367
R595 B.n452 B.n101 163.367
R596 B.n453 B.n452 163.367
R597 B.n454 B.n453 163.367
R598 B.n454 B.n99 163.367
R599 B.n458 B.n99 163.367
R600 B.n459 B.n458 163.367
R601 B.n460 B.n459 163.367
R602 B.n460 B.n97 163.367
R603 B.n464 B.n97 163.367
R604 B.n465 B.n464 163.367
R605 B.n466 B.n465 163.367
R606 B.n466 B.n95 163.367
R607 B.n470 B.n95 163.367
R608 B.n471 B.n470 163.367
R609 B.n472 B.n471 163.367
R610 B.n472 B.n93 163.367
R611 B.n476 B.n93 163.367
R612 B.n477 B.n476 163.367
R613 B.n478 B.n477 163.367
R614 B.n478 B.n91 163.367
R615 B.n482 B.n91 163.367
R616 B.n483 B.n482 163.367
R617 B.n484 B.n483 163.367
R618 B.n484 B.n89 163.367
R619 B.n488 B.n89 163.367
R620 B.n489 B.n488 163.367
R621 B.n490 B.n489 163.367
R622 B.n490 B.n87 163.367
R623 B.n494 B.n87 163.367
R624 B.n495 B.n494 163.367
R625 B.n496 B.n495 163.367
R626 B.n496 B.n85 163.367
R627 B.n500 B.n85 163.367
R628 B.n501 B.n500 163.367
R629 B.n502 B.n501 163.367
R630 B.n502 B.n83 163.367
R631 B.n506 B.n83 163.367
R632 B.n507 B.n506 163.367
R633 B.n508 B.n507 163.367
R634 B.n508 B.n81 163.367
R635 B.n512 B.n81 163.367
R636 B.n513 B.n512 163.367
R637 B.n514 B.n513 163.367
R638 B.n514 B.n79 163.367
R639 B.n518 B.n79 163.367
R640 B.n519 B.n518 163.367
R641 B.n520 B.n519 163.367
R642 B.n520 B.n77 163.367
R643 B.n524 B.n77 163.367
R644 B.n525 B.n524 163.367
R645 B.n526 B.n525 163.367
R646 B.n526 B.n75 163.367
R647 B.n530 B.n75 163.367
R648 B.n671 B.n670 163.367
R649 B.n670 B.n25 163.367
R650 B.n666 B.n25 163.367
R651 B.n666 B.n665 163.367
R652 B.n665 B.n664 163.367
R653 B.n664 B.n27 163.367
R654 B.n660 B.n27 163.367
R655 B.n660 B.n659 163.367
R656 B.n659 B.n658 163.367
R657 B.n658 B.n29 163.367
R658 B.n654 B.n29 163.367
R659 B.n654 B.n653 163.367
R660 B.n653 B.n652 163.367
R661 B.n652 B.n31 163.367
R662 B.n648 B.n31 163.367
R663 B.n648 B.n647 163.367
R664 B.n647 B.n646 163.367
R665 B.n646 B.n33 163.367
R666 B.n642 B.n33 163.367
R667 B.n642 B.n641 163.367
R668 B.n641 B.n640 163.367
R669 B.n640 B.n35 163.367
R670 B.n636 B.n35 163.367
R671 B.n636 B.n635 163.367
R672 B.n635 B.n634 163.367
R673 B.n634 B.n37 163.367
R674 B.n630 B.n37 163.367
R675 B.n630 B.n629 163.367
R676 B.n629 B.n628 163.367
R677 B.n628 B.n39 163.367
R678 B.n624 B.n39 163.367
R679 B.n624 B.n623 163.367
R680 B.n623 B.n622 163.367
R681 B.n622 B.n41 163.367
R682 B.n618 B.n41 163.367
R683 B.n618 B.n617 163.367
R684 B.n617 B.n616 163.367
R685 B.n616 B.n43 163.367
R686 B.n612 B.n43 163.367
R687 B.n612 B.n611 163.367
R688 B.n611 B.n610 163.367
R689 B.n610 B.n45 163.367
R690 B.n605 B.n45 163.367
R691 B.n605 B.n604 163.367
R692 B.n604 B.n603 163.367
R693 B.n603 B.n49 163.367
R694 B.n599 B.n49 163.367
R695 B.n599 B.n598 163.367
R696 B.n598 B.n597 163.367
R697 B.n597 B.n51 163.367
R698 B.n592 B.n51 163.367
R699 B.n592 B.n591 163.367
R700 B.n591 B.n590 163.367
R701 B.n590 B.n55 163.367
R702 B.n586 B.n55 163.367
R703 B.n586 B.n585 163.367
R704 B.n585 B.n584 163.367
R705 B.n584 B.n57 163.367
R706 B.n580 B.n57 163.367
R707 B.n580 B.n579 163.367
R708 B.n579 B.n578 163.367
R709 B.n578 B.n59 163.367
R710 B.n574 B.n59 163.367
R711 B.n574 B.n573 163.367
R712 B.n573 B.n572 163.367
R713 B.n572 B.n61 163.367
R714 B.n568 B.n61 163.367
R715 B.n568 B.n567 163.367
R716 B.n567 B.n566 163.367
R717 B.n566 B.n63 163.367
R718 B.n562 B.n63 163.367
R719 B.n562 B.n561 163.367
R720 B.n561 B.n560 163.367
R721 B.n560 B.n65 163.367
R722 B.n556 B.n65 163.367
R723 B.n556 B.n555 163.367
R724 B.n555 B.n554 163.367
R725 B.n554 B.n67 163.367
R726 B.n550 B.n67 163.367
R727 B.n550 B.n549 163.367
R728 B.n549 B.n548 163.367
R729 B.n548 B.n69 163.367
R730 B.n544 B.n69 163.367
R731 B.n544 B.n543 163.367
R732 B.n543 B.n542 163.367
R733 B.n542 B.n71 163.367
R734 B.n538 B.n71 163.367
R735 B.n538 B.n537 163.367
R736 B.n537 B.n536 163.367
R737 B.n536 B.n73 163.367
R738 B.n532 B.n73 163.367
R739 B.n532 B.n531 163.367
R740 B.n142 B.n141 59.5399
R741 B.n319 B.n149 59.5399
R742 B.n608 B.n47 59.5399
R743 B.n594 B.n53 59.5399
R744 B.n141 B.n140 39.5641
R745 B.n149 B.n148 39.5641
R746 B.n47 B.n46 39.5641
R747 B.n53 B.n52 39.5641
R748 B.n673 B.n24 36.059
R749 B.n397 B.n396 36.059
R750 B.n257 B.n170 36.059
R751 B.n529 B.n74 36.059
R752 B B.n739 18.0485
R753 B.n669 B.n24 10.6151
R754 B.n669 B.n668 10.6151
R755 B.n668 B.n667 10.6151
R756 B.n667 B.n26 10.6151
R757 B.n663 B.n26 10.6151
R758 B.n663 B.n662 10.6151
R759 B.n662 B.n661 10.6151
R760 B.n661 B.n28 10.6151
R761 B.n657 B.n28 10.6151
R762 B.n657 B.n656 10.6151
R763 B.n656 B.n655 10.6151
R764 B.n655 B.n30 10.6151
R765 B.n651 B.n30 10.6151
R766 B.n651 B.n650 10.6151
R767 B.n650 B.n649 10.6151
R768 B.n649 B.n32 10.6151
R769 B.n645 B.n32 10.6151
R770 B.n645 B.n644 10.6151
R771 B.n644 B.n643 10.6151
R772 B.n643 B.n34 10.6151
R773 B.n639 B.n34 10.6151
R774 B.n639 B.n638 10.6151
R775 B.n638 B.n637 10.6151
R776 B.n637 B.n36 10.6151
R777 B.n633 B.n36 10.6151
R778 B.n633 B.n632 10.6151
R779 B.n632 B.n631 10.6151
R780 B.n631 B.n38 10.6151
R781 B.n627 B.n38 10.6151
R782 B.n627 B.n626 10.6151
R783 B.n626 B.n625 10.6151
R784 B.n625 B.n40 10.6151
R785 B.n621 B.n40 10.6151
R786 B.n621 B.n620 10.6151
R787 B.n620 B.n619 10.6151
R788 B.n619 B.n42 10.6151
R789 B.n615 B.n42 10.6151
R790 B.n615 B.n614 10.6151
R791 B.n614 B.n613 10.6151
R792 B.n613 B.n44 10.6151
R793 B.n609 B.n44 10.6151
R794 B.n607 B.n606 10.6151
R795 B.n606 B.n48 10.6151
R796 B.n602 B.n48 10.6151
R797 B.n602 B.n601 10.6151
R798 B.n601 B.n600 10.6151
R799 B.n600 B.n50 10.6151
R800 B.n596 B.n50 10.6151
R801 B.n596 B.n595 10.6151
R802 B.n593 B.n54 10.6151
R803 B.n589 B.n54 10.6151
R804 B.n589 B.n588 10.6151
R805 B.n588 B.n587 10.6151
R806 B.n587 B.n56 10.6151
R807 B.n583 B.n56 10.6151
R808 B.n583 B.n582 10.6151
R809 B.n582 B.n581 10.6151
R810 B.n581 B.n58 10.6151
R811 B.n577 B.n58 10.6151
R812 B.n577 B.n576 10.6151
R813 B.n576 B.n575 10.6151
R814 B.n575 B.n60 10.6151
R815 B.n571 B.n60 10.6151
R816 B.n571 B.n570 10.6151
R817 B.n570 B.n569 10.6151
R818 B.n569 B.n62 10.6151
R819 B.n565 B.n62 10.6151
R820 B.n565 B.n564 10.6151
R821 B.n564 B.n563 10.6151
R822 B.n563 B.n64 10.6151
R823 B.n559 B.n64 10.6151
R824 B.n559 B.n558 10.6151
R825 B.n558 B.n557 10.6151
R826 B.n557 B.n66 10.6151
R827 B.n553 B.n66 10.6151
R828 B.n553 B.n552 10.6151
R829 B.n552 B.n551 10.6151
R830 B.n551 B.n68 10.6151
R831 B.n547 B.n68 10.6151
R832 B.n547 B.n546 10.6151
R833 B.n546 B.n545 10.6151
R834 B.n545 B.n70 10.6151
R835 B.n541 B.n70 10.6151
R836 B.n541 B.n540 10.6151
R837 B.n540 B.n539 10.6151
R838 B.n539 B.n72 10.6151
R839 B.n535 B.n72 10.6151
R840 B.n535 B.n534 10.6151
R841 B.n534 B.n533 10.6151
R842 B.n533 B.n74 10.6151
R843 B.n397 B.n118 10.6151
R844 B.n401 B.n118 10.6151
R845 B.n402 B.n401 10.6151
R846 B.n403 B.n402 10.6151
R847 B.n403 B.n116 10.6151
R848 B.n407 B.n116 10.6151
R849 B.n408 B.n407 10.6151
R850 B.n409 B.n408 10.6151
R851 B.n409 B.n114 10.6151
R852 B.n413 B.n114 10.6151
R853 B.n414 B.n413 10.6151
R854 B.n415 B.n414 10.6151
R855 B.n415 B.n112 10.6151
R856 B.n419 B.n112 10.6151
R857 B.n420 B.n419 10.6151
R858 B.n421 B.n420 10.6151
R859 B.n421 B.n110 10.6151
R860 B.n425 B.n110 10.6151
R861 B.n426 B.n425 10.6151
R862 B.n427 B.n426 10.6151
R863 B.n427 B.n108 10.6151
R864 B.n431 B.n108 10.6151
R865 B.n432 B.n431 10.6151
R866 B.n433 B.n432 10.6151
R867 B.n433 B.n106 10.6151
R868 B.n437 B.n106 10.6151
R869 B.n438 B.n437 10.6151
R870 B.n439 B.n438 10.6151
R871 B.n439 B.n104 10.6151
R872 B.n443 B.n104 10.6151
R873 B.n444 B.n443 10.6151
R874 B.n445 B.n444 10.6151
R875 B.n445 B.n102 10.6151
R876 B.n449 B.n102 10.6151
R877 B.n450 B.n449 10.6151
R878 B.n451 B.n450 10.6151
R879 B.n451 B.n100 10.6151
R880 B.n455 B.n100 10.6151
R881 B.n456 B.n455 10.6151
R882 B.n457 B.n456 10.6151
R883 B.n457 B.n98 10.6151
R884 B.n461 B.n98 10.6151
R885 B.n462 B.n461 10.6151
R886 B.n463 B.n462 10.6151
R887 B.n463 B.n96 10.6151
R888 B.n467 B.n96 10.6151
R889 B.n468 B.n467 10.6151
R890 B.n469 B.n468 10.6151
R891 B.n469 B.n94 10.6151
R892 B.n473 B.n94 10.6151
R893 B.n474 B.n473 10.6151
R894 B.n475 B.n474 10.6151
R895 B.n475 B.n92 10.6151
R896 B.n479 B.n92 10.6151
R897 B.n480 B.n479 10.6151
R898 B.n481 B.n480 10.6151
R899 B.n481 B.n90 10.6151
R900 B.n485 B.n90 10.6151
R901 B.n486 B.n485 10.6151
R902 B.n487 B.n486 10.6151
R903 B.n487 B.n88 10.6151
R904 B.n491 B.n88 10.6151
R905 B.n492 B.n491 10.6151
R906 B.n493 B.n492 10.6151
R907 B.n493 B.n86 10.6151
R908 B.n497 B.n86 10.6151
R909 B.n498 B.n497 10.6151
R910 B.n499 B.n498 10.6151
R911 B.n499 B.n84 10.6151
R912 B.n503 B.n84 10.6151
R913 B.n504 B.n503 10.6151
R914 B.n505 B.n504 10.6151
R915 B.n505 B.n82 10.6151
R916 B.n509 B.n82 10.6151
R917 B.n510 B.n509 10.6151
R918 B.n511 B.n510 10.6151
R919 B.n511 B.n80 10.6151
R920 B.n515 B.n80 10.6151
R921 B.n516 B.n515 10.6151
R922 B.n517 B.n516 10.6151
R923 B.n517 B.n78 10.6151
R924 B.n521 B.n78 10.6151
R925 B.n522 B.n521 10.6151
R926 B.n523 B.n522 10.6151
R927 B.n523 B.n76 10.6151
R928 B.n527 B.n76 10.6151
R929 B.n528 B.n527 10.6151
R930 B.n529 B.n528 10.6151
R931 B.n258 B.n257 10.6151
R932 B.n259 B.n258 10.6151
R933 B.n259 B.n168 10.6151
R934 B.n263 B.n168 10.6151
R935 B.n264 B.n263 10.6151
R936 B.n265 B.n264 10.6151
R937 B.n265 B.n166 10.6151
R938 B.n269 B.n166 10.6151
R939 B.n270 B.n269 10.6151
R940 B.n271 B.n270 10.6151
R941 B.n271 B.n164 10.6151
R942 B.n275 B.n164 10.6151
R943 B.n276 B.n275 10.6151
R944 B.n277 B.n276 10.6151
R945 B.n277 B.n162 10.6151
R946 B.n281 B.n162 10.6151
R947 B.n282 B.n281 10.6151
R948 B.n283 B.n282 10.6151
R949 B.n283 B.n160 10.6151
R950 B.n287 B.n160 10.6151
R951 B.n288 B.n287 10.6151
R952 B.n289 B.n288 10.6151
R953 B.n289 B.n158 10.6151
R954 B.n293 B.n158 10.6151
R955 B.n294 B.n293 10.6151
R956 B.n295 B.n294 10.6151
R957 B.n295 B.n156 10.6151
R958 B.n299 B.n156 10.6151
R959 B.n300 B.n299 10.6151
R960 B.n301 B.n300 10.6151
R961 B.n301 B.n154 10.6151
R962 B.n305 B.n154 10.6151
R963 B.n306 B.n305 10.6151
R964 B.n307 B.n306 10.6151
R965 B.n307 B.n152 10.6151
R966 B.n311 B.n152 10.6151
R967 B.n312 B.n311 10.6151
R968 B.n313 B.n312 10.6151
R969 B.n313 B.n150 10.6151
R970 B.n317 B.n150 10.6151
R971 B.n318 B.n317 10.6151
R972 B.n320 B.n146 10.6151
R973 B.n324 B.n146 10.6151
R974 B.n325 B.n324 10.6151
R975 B.n326 B.n325 10.6151
R976 B.n326 B.n144 10.6151
R977 B.n330 B.n144 10.6151
R978 B.n331 B.n330 10.6151
R979 B.n332 B.n331 10.6151
R980 B.n336 B.n335 10.6151
R981 B.n337 B.n336 10.6151
R982 B.n337 B.n138 10.6151
R983 B.n341 B.n138 10.6151
R984 B.n342 B.n341 10.6151
R985 B.n343 B.n342 10.6151
R986 B.n343 B.n136 10.6151
R987 B.n347 B.n136 10.6151
R988 B.n348 B.n347 10.6151
R989 B.n349 B.n348 10.6151
R990 B.n349 B.n134 10.6151
R991 B.n353 B.n134 10.6151
R992 B.n354 B.n353 10.6151
R993 B.n355 B.n354 10.6151
R994 B.n355 B.n132 10.6151
R995 B.n359 B.n132 10.6151
R996 B.n360 B.n359 10.6151
R997 B.n361 B.n360 10.6151
R998 B.n361 B.n130 10.6151
R999 B.n365 B.n130 10.6151
R1000 B.n366 B.n365 10.6151
R1001 B.n367 B.n366 10.6151
R1002 B.n367 B.n128 10.6151
R1003 B.n371 B.n128 10.6151
R1004 B.n372 B.n371 10.6151
R1005 B.n373 B.n372 10.6151
R1006 B.n373 B.n126 10.6151
R1007 B.n377 B.n126 10.6151
R1008 B.n378 B.n377 10.6151
R1009 B.n379 B.n378 10.6151
R1010 B.n379 B.n124 10.6151
R1011 B.n383 B.n124 10.6151
R1012 B.n384 B.n383 10.6151
R1013 B.n385 B.n384 10.6151
R1014 B.n385 B.n122 10.6151
R1015 B.n389 B.n122 10.6151
R1016 B.n390 B.n389 10.6151
R1017 B.n391 B.n390 10.6151
R1018 B.n391 B.n120 10.6151
R1019 B.n395 B.n120 10.6151
R1020 B.n396 B.n395 10.6151
R1021 B.n253 B.n170 10.6151
R1022 B.n253 B.n252 10.6151
R1023 B.n252 B.n251 10.6151
R1024 B.n251 B.n172 10.6151
R1025 B.n247 B.n172 10.6151
R1026 B.n247 B.n246 10.6151
R1027 B.n246 B.n245 10.6151
R1028 B.n245 B.n174 10.6151
R1029 B.n241 B.n174 10.6151
R1030 B.n241 B.n240 10.6151
R1031 B.n240 B.n239 10.6151
R1032 B.n239 B.n176 10.6151
R1033 B.n235 B.n176 10.6151
R1034 B.n235 B.n234 10.6151
R1035 B.n234 B.n233 10.6151
R1036 B.n233 B.n178 10.6151
R1037 B.n229 B.n178 10.6151
R1038 B.n229 B.n228 10.6151
R1039 B.n228 B.n227 10.6151
R1040 B.n227 B.n180 10.6151
R1041 B.n223 B.n180 10.6151
R1042 B.n223 B.n222 10.6151
R1043 B.n222 B.n221 10.6151
R1044 B.n221 B.n182 10.6151
R1045 B.n217 B.n182 10.6151
R1046 B.n217 B.n216 10.6151
R1047 B.n216 B.n215 10.6151
R1048 B.n215 B.n184 10.6151
R1049 B.n211 B.n184 10.6151
R1050 B.n211 B.n210 10.6151
R1051 B.n210 B.n209 10.6151
R1052 B.n209 B.n186 10.6151
R1053 B.n205 B.n186 10.6151
R1054 B.n205 B.n204 10.6151
R1055 B.n204 B.n203 10.6151
R1056 B.n203 B.n188 10.6151
R1057 B.n199 B.n188 10.6151
R1058 B.n199 B.n198 10.6151
R1059 B.n198 B.n197 10.6151
R1060 B.n197 B.n190 10.6151
R1061 B.n193 B.n190 10.6151
R1062 B.n193 B.n192 10.6151
R1063 B.n192 B.n0 10.6151
R1064 B.n735 B.n1 10.6151
R1065 B.n735 B.n734 10.6151
R1066 B.n734 B.n733 10.6151
R1067 B.n733 B.n4 10.6151
R1068 B.n729 B.n4 10.6151
R1069 B.n729 B.n728 10.6151
R1070 B.n728 B.n727 10.6151
R1071 B.n727 B.n6 10.6151
R1072 B.n723 B.n6 10.6151
R1073 B.n723 B.n722 10.6151
R1074 B.n722 B.n721 10.6151
R1075 B.n721 B.n8 10.6151
R1076 B.n717 B.n8 10.6151
R1077 B.n717 B.n716 10.6151
R1078 B.n716 B.n715 10.6151
R1079 B.n715 B.n10 10.6151
R1080 B.n711 B.n10 10.6151
R1081 B.n711 B.n710 10.6151
R1082 B.n710 B.n709 10.6151
R1083 B.n709 B.n12 10.6151
R1084 B.n705 B.n12 10.6151
R1085 B.n705 B.n704 10.6151
R1086 B.n704 B.n703 10.6151
R1087 B.n703 B.n14 10.6151
R1088 B.n699 B.n14 10.6151
R1089 B.n699 B.n698 10.6151
R1090 B.n698 B.n697 10.6151
R1091 B.n697 B.n16 10.6151
R1092 B.n693 B.n16 10.6151
R1093 B.n693 B.n692 10.6151
R1094 B.n692 B.n691 10.6151
R1095 B.n691 B.n18 10.6151
R1096 B.n687 B.n18 10.6151
R1097 B.n687 B.n686 10.6151
R1098 B.n686 B.n685 10.6151
R1099 B.n685 B.n20 10.6151
R1100 B.n681 B.n20 10.6151
R1101 B.n681 B.n680 10.6151
R1102 B.n680 B.n679 10.6151
R1103 B.n679 B.n22 10.6151
R1104 B.n675 B.n22 10.6151
R1105 B.n675 B.n674 10.6151
R1106 B.n674 B.n673 10.6151
R1107 B.n608 B.n607 6.5566
R1108 B.n595 B.n594 6.5566
R1109 B.n320 B.n319 6.5566
R1110 B.n332 B.n142 6.5566
R1111 B.n609 B.n608 4.05904
R1112 B.n594 B.n593 4.05904
R1113 B.n319 B.n318 4.05904
R1114 B.n335 B.n142 4.05904
R1115 B.n739 B.n0 2.81026
R1116 B.n739 B.n1 2.81026
R1117 VP.n16 VP.t8 200.415
R1118 VP.n41 VP.n40 181.852
R1119 VP.n70 VP.n69 181.852
R1120 VP.n39 VP.n38 181.852
R1121 VP.n55 VP.t7 170.673
R1122 VP.n41 VP.t4 170.673
R1123 VP.n48 VP.t6 170.673
R1124 VP.n62 VP.t3 170.673
R1125 VP.n69 VP.t2 170.673
R1126 VP.n24 VP.t0 170.673
R1127 VP.n38 VP.t1 170.673
R1128 VP.n31 VP.t5 170.673
R1129 VP.n17 VP.t9 170.673
R1130 VP.n18 VP.n15 161.3
R1131 VP.n20 VP.n19 161.3
R1132 VP.n21 VP.n14 161.3
R1133 VP.n23 VP.n22 161.3
R1134 VP.n24 VP.n13 161.3
R1135 VP.n26 VP.n25 161.3
R1136 VP.n27 VP.n12 161.3
R1137 VP.n29 VP.n28 161.3
R1138 VP.n30 VP.n11 161.3
R1139 VP.n33 VP.n32 161.3
R1140 VP.n34 VP.n10 161.3
R1141 VP.n36 VP.n35 161.3
R1142 VP.n37 VP.n9 161.3
R1143 VP.n68 VP.n0 161.3
R1144 VP.n67 VP.n66 161.3
R1145 VP.n65 VP.n1 161.3
R1146 VP.n64 VP.n63 161.3
R1147 VP.n61 VP.n2 161.3
R1148 VP.n60 VP.n59 161.3
R1149 VP.n58 VP.n3 161.3
R1150 VP.n57 VP.n56 161.3
R1151 VP.n55 VP.n4 161.3
R1152 VP.n54 VP.n53 161.3
R1153 VP.n52 VP.n5 161.3
R1154 VP.n51 VP.n50 161.3
R1155 VP.n49 VP.n6 161.3
R1156 VP.n47 VP.n46 161.3
R1157 VP.n45 VP.n7 161.3
R1158 VP.n44 VP.n43 161.3
R1159 VP.n42 VP.n8 161.3
R1160 VP.n17 VP.n16 66.2588
R1161 VP.n40 VP.n39 48.2429
R1162 VP.n43 VP.n7 46.321
R1163 VP.n67 VP.n1 46.321
R1164 VP.n36 VP.n10 46.321
R1165 VP.n50 VP.n5 42.4359
R1166 VP.n60 VP.n3 42.4359
R1167 VP.n29 VP.n12 42.4359
R1168 VP.n19 VP.n14 42.4359
R1169 VP.n54 VP.n5 38.5509
R1170 VP.n56 VP.n3 38.5509
R1171 VP.n25 VP.n12 38.5509
R1172 VP.n23 VP.n14 38.5509
R1173 VP.n47 VP.n7 34.6658
R1174 VP.n63 VP.n1 34.6658
R1175 VP.n32 VP.n10 34.6658
R1176 VP.n43 VP.n42 24.4675
R1177 VP.n50 VP.n49 24.4675
R1178 VP.n55 VP.n54 24.4675
R1179 VP.n56 VP.n55 24.4675
R1180 VP.n61 VP.n60 24.4675
R1181 VP.n68 VP.n67 24.4675
R1182 VP.n37 VP.n36 24.4675
R1183 VP.n30 VP.n29 24.4675
R1184 VP.n24 VP.n23 24.4675
R1185 VP.n25 VP.n24 24.4675
R1186 VP.n19 VP.n18 24.4675
R1187 VP.n48 VP.n47 22.5101
R1188 VP.n63 VP.n62 22.5101
R1189 VP.n32 VP.n31 22.5101
R1190 VP.n16 VP.n15 18.5717
R1191 VP.n42 VP.n41 3.91522
R1192 VP.n69 VP.n68 3.91522
R1193 VP.n38 VP.n37 3.91522
R1194 VP.n49 VP.n48 1.95786
R1195 VP.n62 VP.n61 1.95786
R1196 VP.n31 VP.n30 1.95786
R1197 VP.n18 VP.n17 1.95786
R1198 VP.n20 VP.n15 0.189894
R1199 VP.n21 VP.n20 0.189894
R1200 VP.n22 VP.n21 0.189894
R1201 VP.n22 VP.n13 0.189894
R1202 VP.n26 VP.n13 0.189894
R1203 VP.n27 VP.n26 0.189894
R1204 VP.n28 VP.n27 0.189894
R1205 VP.n28 VP.n11 0.189894
R1206 VP.n33 VP.n11 0.189894
R1207 VP.n34 VP.n33 0.189894
R1208 VP.n35 VP.n34 0.189894
R1209 VP.n35 VP.n9 0.189894
R1210 VP.n39 VP.n9 0.189894
R1211 VP.n40 VP.n8 0.189894
R1212 VP.n44 VP.n8 0.189894
R1213 VP.n45 VP.n44 0.189894
R1214 VP.n46 VP.n45 0.189894
R1215 VP.n46 VP.n6 0.189894
R1216 VP.n51 VP.n6 0.189894
R1217 VP.n52 VP.n51 0.189894
R1218 VP.n53 VP.n52 0.189894
R1219 VP.n53 VP.n4 0.189894
R1220 VP.n57 VP.n4 0.189894
R1221 VP.n58 VP.n57 0.189894
R1222 VP.n59 VP.n58 0.189894
R1223 VP.n59 VP.n2 0.189894
R1224 VP.n64 VP.n2 0.189894
R1225 VP.n65 VP.n64 0.189894
R1226 VP.n66 VP.n65 0.189894
R1227 VP.n66 VP.n0 0.189894
R1228 VP.n70 VP.n0 0.189894
R1229 VP VP.n70 0.0516364
R1230 VTAIL.n272 VTAIL.n212 756.745
R1231 VTAIL.n62 VTAIL.n2 756.745
R1232 VTAIL.n206 VTAIL.n146 756.745
R1233 VTAIL.n136 VTAIL.n76 756.745
R1234 VTAIL.n232 VTAIL.n231 585
R1235 VTAIL.n237 VTAIL.n236 585
R1236 VTAIL.n239 VTAIL.n238 585
R1237 VTAIL.n228 VTAIL.n227 585
R1238 VTAIL.n245 VTAIL.n244 585
R1239 VTAIL.n247 VTAIL.n246 585
R1240 VTAIL.n224 VTAIL.n223 585
R1241 VTAIL.n254 VTAIL.n253 585
R1242 VTAIL.n255 VTAIL.n222 585
R1243 VTAIL.n257 VTAIL.n256 585
R1244 VTAIL.n220 VTAIL.n219 585
R1245 VTAIL.n263 VTAIL.n262 585
R1246 VTAIL.n265 VTAIL.n264 585
R1247 VTAIL.n216 VTAIL.n215 585
R1248 VTAIL.n271 VTAIL.n270 585
R1249 VTAIL.n273 VTAIL.n272 585
R1250 VTAIL.n22 VTAIL.n21 585
R1251 VTAIL.n27 VTAIL.n26 585
R1252 VTAIL.n29 VTAIL.n28 585
R1253 VTAIL.n18 VTAIL.n17 585
R1254 VTAIL.n35 VTAIL.n34 585
R1255 VTAIL.n37 VTAIL.n36 585
R1256 VTAIL.n14 VTAIL.n13 585
R1257 VTAIL.n44 VTAIL.n43 585
R1258 VTAIL.n45 VTAIL.n12 585
R1259 VTAIL.n47 VTAIL.n46 585
R1260 VTAIL.n10 VTAIL.n9 585
R1261 VTAIL.n53 VTAIL.n52 585
R1262 VTAIL.n55 VTAIL.n54 585
R1263 VTAIL.n6 VTAIL.n5 585
R1264 VTAIL.n61 VTAIL.n60 585
R1265 VTAIL.n63 VTAIL.n62 585
R1266 VTAIL.n207 VTAIL.n206 585
R1267 VTAIL.n205 VTAIL.n204 585
R1268 VTAIL.n150 VTAIL.n149 585
R1269 VTAIL.n199 VTAIL.n198 585
R1270 VTAIL.n197 VTAIL.n196 585
R1271 VTAIL.n154 VTAIL.n153 585
R1272 VTAIL.n191 VTAIL.n190 585
R1273 VTAIL.n189 VTAIL.n156 585
R1274 VTAIL.n188 VTAIL.n187 585
R1275 VTAIL.n159 VTAIL.n157 585
R1276 VTAIL.n182 VTAIL.n181 585
R1277 VTAIL.n180 VTAIL.n179 585
R1278 VTAIL.n163 VTAIL.n162 585
R1279 VTAIL.n174 VTAIL.n173 585
R1280 VTAIL.n172 VTAIL.n171 585
R1281 VTAIL.n167 VTAIL.n166 585
R1282 VTAIL.n137 VTAIL.n136 585
R1283 VTAIL.n135 VTAIL.n134 585
R1284 VTAIL.n80 VTAIL.n79 585
R1285 VTAIL.n129 VTAIL.n128 585
R1286 VTAIL.n127 VTAIL.n126 585
R1287 VTAIL.n84 VTAIL.n83 585
R1288 VTAIL.n121 VTAIL.n120 585
R1289 VTAIL.n119 VTAIL.n86 585
R1290 VTAIL.n118 VTAIL.n117 585
R1291 VTAIL.n89 VTAIL.n87 585
R1292 VTAIL.n112 VTAIL.n111 585
R1293 VTAIL.n110 VTAIL.n109 585
R1294 VTAIL.n93 VTAIL.n92 585
R1295 VTAIL.n104 VTAIL.n103 585
R1296 VTAIL.n102 VTAIL.n101 585
R1297 VTAIL.n97 VTAIL.n96 585
R1298 VTAIL.n233 VTAIL.t1 329.036
R1299 VTAIL.n23 VTAIL.t12 329.036
R1300 VTAIL.n168 VTAIL.t14 329.036
R1301 VTAIL.n98 VTAIL.t7 329.036
R1302 VTAIL.n237 VTAIL.n231 171.744
R1303 VTAIL.n238 VTAIL.n237 171.744
R1304 VTAIL.n238 VTAIL.n227 171.744
R1305 VTAIL.n245 VTAIL.n227 171.744
R1306 VTAIL.n246 VTAIL.n245 171.744
R1307 VTAIL.n246 VTAIL.n223 171.744
R1308 VTAIL.n254 VTAIL.n223 171.744
R1309 VTAIL.n255 VTAIL.n254 171.744
R1310 VTAIL.n256 VTAIL.n255 171.744
R1311 VTAIL.n256 VTAIL.n219 171.744
R1312 VTAIL.n263 VTAIL.n219 171.744
R1313 VTAIL.n264 VTAIL.n263 171.744
R1314 VTAIL.n264 VTAIL.n215 171.744
R1315 VTAIL.n271 VTAIL.n215 171.744
R1316 VTAIL.n272 VTAIL.n271 171.744
R1317 VTAIL.n27 VTAIL.n21 171.744
R1318 VTAIL.n28 VTAIL.n27 171.744
R1319 VTAIL.n28 VTAIL.n17 171.744
R1320 VTAIL.n35 VTAIL.n17 171.744
R1321 VTAIL.n36 VTAIL.n35 171.744
R1322 VTAIL.n36 VTAIL.n13 171.744
R1323 VTAIL.n44 VTAIL.n13 171.744
R1324 VTAIL.n45 VTAIL.n44 171.744
R1325 VTAIL.n46 VTAIL.n45 171.744
R1326 VTAIL.n46 VTAIL.n9 171.744
R1327 VTAIL.n53 VTAIL.n9 171.744
R1328 VTAIL.n54 VTAIL.n53 171.744
R1329 VTAIL.n54 VTAIL.n5 171.744
R1330 VTAIL.n61 VTAIL.n5 171.744
R1331 VTAIL.n62 VTAIL.n61 171.744
R1332 VTAIL.n206 VTAIL.n205 171.744
R1333 VTAIL.n205 VTAIL.n149 171.744
R1334 VTAIL.n198 VTAIL.n149 171.744
R1335 VTAIL.n198 VTAIL.n197 171.744
R1336 VTAIL.n197 VTAIL.n153 171.744
R1337 VTAIL.n190 VTAIL.n153 171.744
R1338 VTAIL.n190 VTAIL.n189 171.744
R1339 VTAIL.n189 VTAIL.n188 171.744
R1340 VTAIL.n188 VTAIL.n157 171.744
R1341 VTAIL.n181 VTAIL.n157 171.744
R1342 VTAIL.n181 VTAIL.n180 171.744
R1343 VTAIL.n180 VTAIL.n162 171.744
R1344 VTAIL.n173 VTAIL.n162 171.744
R1345 VTAIL.n173 VTAIL.n172 171.744
R1346 VTAIL.n172 VTAIL.n166 171.744
R1347 VTAIL.n136 VTAIL.n135 171.744
R1348 VTAIL.n135 VTAIL.n79 171.744
R1349 VTAIL.n128 VTAIL.n79 171.744
R1350 VTAIL.n128 VTAIL.n127 171.744
R1351 VTAIL.n127 VTAIL.n83 171.744
R1352 VTAIL.n120 VTAIL.n83 171.744
R1353 VTAIL.n120 VTAIL.n119 171.744
R1354 VTAIL.n119 VTAIL.n118 171.744
R1355 VTAIL.n118 VTAIL.n87 171.744
R1356 VTAIL.n111 VTAIL.n87 171.744
R1357 VTAIL.n111 VTAIL.n110 171.744
R1358 VTAIL.n110 VTAIL.n92 171.744
R1359 VTAIL.n103 VTAIL.n92 171.744
R1360 VTAIL.n103 VTAIL.n102 171.744
R1361 VTAIL.n102 VTAIL.n96 171.744
R1362 VTAIL.t1 VTAIL.n231 85.8723
R1363 VTAIL.t12 VTAIL.n21 85.8723
R1364 VTAIL.t14 VTAIL.n166 85.8723
R1365 VTAIL.t7 VTAIL.n96 85.8723
R1366 VTAIL.n145 VTAIL.n144 56.9665
R1367 VTAIL.n143 VTAIL.n142 56.9665
R1368 VTAIL.n75 VTAIL.n74 56.9665
R1369 VTAIL.n73 VTAIL.n72 56.9665
R1370 VTAIL.n279 VTAIL.n278 56.9663
R1371 VTAIL.n1 VTAIL.n0 56.9663
R1372 VTAIL.n69 VTAIL.n68 56.9663
R1373 VTAIL.n71 VTAIL.n70 56.9663
R1374 VTAIL.n277 VTAIL.n276 31.9914
R1375 VTAIL.n67 VTAIL.n66 31.9914
R1376 VTAIL.n211 VTAIL.n210 31.9914
R1377 VTAIL.n141 VTAIL.n140 31.9914
R1378 VTAIL.n73 VTAIL.n71 26.3238
R1379 VTAIL.n277 VTAIL.n211 24.5652
R1380 VTAIL.n257 VTAIL.n222 13.1884
R1381 VTAIL.n47 VTAIL.n12 13.1884
R1382 VTAIL.n191 VTAIL.n156 13.1884
R1383 VTAIL.n121 VTAIL.n86 13.1884
R1384 VTAIL.n253 VTAIL.n252 12.8005
R1385 VTAIL.n258 VTAIL.n220 12.8005
R1386 VTAIL.n43 VTAIL.n42 12.8005
R1387 VTAIL.n48 VTAIL.n10 12.8005
R1388 VTAIL.n192 VTAIL.n154 12.8005
R1389 VTAIL.n187 VTAIL.n158 12.8005
R1390 VTAIL.n122 VTAIL.n84 12.8005
R1391 VTAIL.n117 VTAIL.n88 12.8005
R1392 VTAIL.n251 VTAIL.n224 12.0247
R1393 VTAIL.n262 VTAIL.n261 12.0247
R1394 VTAIL.n41 VTAIL.n14 12.0247
R1395 VTAIL.n52 VTAIL.n51 12.0247
R1396 VTAIL.n196 VTAIL.n195 12.0247
R1397 VTAIL.n186 VTAIL.n159 12.0247
R1398 VTAIL.n126 VTAIL.n125 12.0247
R1399 VTAIL.n116 VTAIL.n89 12.0247
R1400 VTAIL.n248 VTAIL.n247 11.249
R1401 VTAIL.n265 VTAIL.n218 11.249
R1402 VTAIL.n38 VTAIL.n37 11.249
R1403 VTAIL.n55 VTAIL.n8 11.249
R1404 VTAIL.n199 VTAIL.n152 11.249
R1405 VTAIL.n183 VTAIL.n182 11.249
R1406 VTAIL.n129 VTAIL.n82 11.249
R1407 VTAIL.n113 VTAIL.n112 11.249
R1408 VTAIL.n233 VTAIL.n232 10.7239
R1409 VTAIL.n23 VTAIL.n22 10.7239
R1410 VTAIL.n168 VTAIL.n167 10.7239
R1411 VTAIL.n98 VTAIL.n97 10.7239
R1412 VTAIL.n244 VTAIL.n226 10.4732
R1413 VTAIL.n266 VTAIL.n216 10.4732
R1414 VTAIL.n34 VTAIL.n16 10.4732
R1415 VTAIL.n56 VTAIL.n6 10.4732
R1416 VTAIL.n200 VTAIL.n150 10.4732
R1417 VTAIL.n179 VTAIL.n161 10.4732
R1418 VTAIL.n130 VTAIL.n80 10.4732
R1419 VTAIL.n109 VTAIL.n91 10.4732
R1420 VTAIL.n243 VTAIL.n228 9.69747
R1421 VTAIL.n270 VTAIL.n269 9.69747
R1422 VTAIL.n33 VTAIL.n18 9.69747
R1423 VTAIL.n60 VTAIL.n59 9.69747
R1424 VTAIL.n204 VTAIL.n203 9.69747
R1425 VTAIL.n178 VTAIL.n163 9.69747
R1426 VTAIL.n134 VTAIL.n133 9.69747
R1427 VTAIL.n108 VTAIL.n93 9.69747
R1428 VTAIL.n276 VTAIL.n275 9.45567
R1429 VTAIL.n66 VTAIL.n65 9.45567
R1430 VTAIL.n210 VTAIL.n209 9.45567
R1431 VTAIL.n140 VTAIL.n139 9.45567
R1432 VTAIL.n275 VTAIL.n274 9.3005
R1433 VTAIL.n214 VTAIL.n213 9.3005
R1434 VTAIL.n269 VTAIL.n268 9.3005
R1435 VTAIL.n267 VTAIL.n266 9.3005
R1436 VTAIL.n218 VTAIL.n217 9.3005
R1437 VTAIL.n261 VTAIL.n260 9.3005
R1438 VTAIL.n259 VTAIL.n258 9.3005
R1439 VTAIL.n235 VTAIL.n234 9.3005
R1440 VTAIL.n230 VTAIL.n229 9.3005
R1441 VTAIL.n241 VTAIL.n240 9.3005
R1442 VTAIL.n243 VTAIL.n242 9.3005
R1443 VTAIL.n226 VTAIL.n225 9.3005
R1444 VTAIL.n249 VTAIL.n248 9.3005
R1445 VTAIL.n251 VTAIL.n250 9.3005
R1446 VTAIL.n252 VTAIL.n221 9.3005
R1447 VTAIL.n65 VTAIL.n64 9.3005
R1448 VTAIL.n4 VTAIL.n3 9.3005
R1449 VTAIL.n59 VTAIL.n58 9.3005
R1450 VTAIL.n57 VTAIL.n56 9.3005
R1451 VTAIL.n8 VTAIL.n7 9.3005
R1452 VTAIL.n51 VTAIL.n50 9.3005
R1453 VTAIL.n49 VTAIL.n48 9.3005
R1454 VTAIL.n25 VTAIL.n24 9.3005
R1455 VTAIL.n20 VTAIL.n19 9.3005
R1456 VTAIL.n31 VTAIL.n30 9.3005
R1457 VTAIL.n33 VTAIL.n32 9.3005
R1458 VTAIL.n16 VTAIL.n15 9.3005
R1459 VTAIL.n39 VTAIL.n38 9.3005
R1460 VTAIL.n41 VTAIL.n40 9.3005
R1461 VTAIL.n42 VTAIL.n11 9.3005
R1462 VTAIL.n170 VTAIL.n169 9.3005
R1463 VTAIL.n165 VTAIL.n164 9.3005
R1464 VTAIL.n176 VTAIL.n175 9.3005
R1465 VTAIL.n178 VTAIL.n177 9.3005
R1466 VTAIL.n161 VTAIL.n160 9.3005
R1467 VTAIL.n184 VTAIL.n183 9.3005
R1468 VTAIL.n186 VTAIL.n185 9.3005
R1469 VTAIL.n158 VTAIL.n155 9.3005
R1470 VTAIL.n209 VTAIL.n208 9.3005
R1471 VTAIL.n148 VTAIL.n147 9.3005
R1472 VTAIL.n203 VTAIL.n202 9.3005
R1473 VTAIL.n201 VTAIL.n200 9.3005
R1474 VTAIL.n152 VTAIL.n151 9.3005
R1475 VTAIL.n195 VTAIL.n194 9.3005
R1476 VTAIL.n193 VTAIL.n192 9.3005
R1477 VTAIL.n100 VTAIL.n99 9.3005
R1478 VTAIL.n95 VTAIL.n94 9.3005
R1479 VTAIL.n106 VTAIL.n105 9.3005
R1480 VTAIL.n108 VTAIL.n107 9.3005
R1481 VTAIL.n91 VTAIL.n90 9.3005
R1482 VTAIL.n114 VTAIL.n113 9.3005
R1483 VTAIL.n116 VTAIL.n115 9.3005
R1484 VTAIL.n88 VTAIL.n85 9.3005
R1485 VTAIL.n139 VTAIL.n138 9.3005
R1486 VTAIL.n78 VTAIL.n77 9.3005
R1487 VTAIL.n133 VTAIL.n132 9.3005
R1488 VTAIL.n131 VTAIL.n130 9.3005
R1489 VTAIL.n82 VTAIL.n81 9.3005
R1490 VTAIL.n125 VTAIL.n124 9.3005
R1491 VTAIL.n123 VTAIL.n122 9.3005
R1492 VTAIL.n240 VTAIL.n239 8.92171
R1493 VTAIL.n273 VTAIL.n214 8.92171
R1494 VTAIL.n30 VTAIL.n29 8.92171
R1495 VTAIL.n63 VTAIL.n4 8.92171
R1496 VTAIL.n207 VTAIL.n148 8.92171
R1497 VTAIL.n175 VTAIL.n174 8.92171
R1498 VTAIL.n137 VTAIL.n78 8.92171
R1499 VTAIL.n105 VTAIL.n104 8.92171
R1500 VTAIL.n236 VTAIL.n230 8.14595
R1501 VTAIL.n274 VTAIL.n212 8.14595
R1502 VTAIL.n26 VTAIL.n20 8.14595
R1503 VTAIL.n64 VTAIL.n2 8.14595
R1504 VTAIL.n208 VTAIL.n146 8.14595
R1505 VTAIL.n171 VTAIL.n165 8.14595
R1506 VTAIL.n138 VTAIL.n76 8.14595
R1507 VTAIL.n101 VTAIL.n95 8.14595
R1508 VTAIL.n235 VTAIL.n232 7.3702
R1509 VTAIL.n25 VTAIL.n22 7.3702
R1510 VTAIL.n170 VTAIL.n167 7.3702
R1511 VTAIL.n100 VTAIL.n97 7.3702
R1512 VTAIL.n236 VTAIL.n235 5.81868
R1513 VTAIL.n276 VTAIL.n212 5.81868
R1514 VTAIL.n26 VTAIL.n25 5.81868
R1515 VTAIL.n66 VTAIL.n2 5.81868
R1516 VTAIL.n210 VTAIL.n146 5.81868
R1517 VTAIL.n171 VTAIL.n170 5.81868
R1518 VTAIL.n140 VTAIL.n76 5.81868
R1519 VTAIL.n101 VTAIL.n100 5.81868
R1520 VTAIL.n239 VTAIL.n230 5.04292
R1521 VTAIL.n274 VTAIL.n273 5.04292
R1522 VTAIL.n29 VTAIL.n20 5.04292
R1523 VTAIL.n64 VTAIL.n63 5.04292
R1524 VTAIL.n208 VTAIL.n207 5.04292
R1525 VTAIL.n174 VTAIL.n165 5.04292
R1526 VTAIL.n138 VTAIL.n137 5.04292
R1527 VTAIL.n104 VTAIL.n95 5.04292
R1528 VTAIL.n240 VTAIL.n228 4.26717
R1529 VTAIL.n270 VTAIL.n214 4.26717
R1530 VTAIL.n30 VTAIL.n18 4.26717
R1531 VTAIL.n60 VTAIL.n4 4.26717
R1532 VTAIL.n204 VTAIL.n148 4.26717
R1533 VTAIL.n175 VTAIL.n163 4.26717
R1534 VTAIL.n134 VTAIL.n78 4.26717
R1535 VTAIL.n105 VTAIL.n93 4.26717
R1536 VTAIL.n244 VTAIL.n243 3.49141
R1537 VTAIL.n269 VTAIL.n216 3.49141
R1538 VTAIL.n34 VTAIL.n33 3.49141
R1539 VTAIL.n59 VTAIL.n6 3.49141
R1540 VTAIL.n203 VTAIL.n150 3.49141
R1541 VTAIL.n179 VTAIL.n178 3.49141
R1542 VTAIL.n133 VTAIL.n80 3.49141
R1543 VTAIL.n109 VTAIL.n108 3.49141
R1544 VTAIL.n247 VTAIL.n226 2.71565
R1545 VTAIL.n266 VTAIL.n265 2.71565
R1546 VTAIL.n37 VTAIL.n16 2.71565
R1547 VTAIL.n56 VTAIL.n55 2.71565
R1548 VTAIL.n200 VTAIL.n199 2.71565
R1549 VTAIL.n182 VTAIL.n161 2.71565
R1550 VTAIL.n130 VTAIL.n129 2.71565
R1551 VTAIL.n112 VTAIL.n91 2.71565
R1552 VTAIL.n278 VTAIL.t3 2.68465
R1553 VTAIL.n278 VTAIL.t6 2.68465
R1554 VTAIL.n0 VTAIL.t4 2.68465
R1555 VTAIL.n0 VTAIL.t2 2.68465
R1556 VTAIL.n68 VTAIL.t18 2.68465
R1557 VTAIL.n68 VTAIL.t11 2.68465
R1558 VTAIL.n70 VTAIL.t16 2.68465
R1559 VTAIL.n70 VTAIL.t17 2.68465
R1560 VTAIL.n144 VTAIL.t13 2.68465
R1561 VTAIL.n144 VTAIL.t19 2.68465
R1562 VTAIL.n142 VTAIL.t15 2.68465
R1563 VTAIL.n142 VTAIL.t10 2.68465
R1564 VTAIL.n74 VTAIL.t5 2.68465
R1565 VTAIL.n74 VTAIL.t0 2.68465
R1566 VTAIL.n72 VTAIL.t8 2.68465
R1567 VTAIL.n72 VTAIL.t9 2.68465
R1568 VTAIL.n169 VTAIL.n168 2.41282
R1569 VTAIL.n99 VTAIL.n98 2.41282
R1570 VTAIL.n234 VTAIL.n233 2.41282
R1571 VTAIL.n24 VTAIL.n23 2.41282
R1572 VTAIL.n248 VTAIL.n224 1.93989
R1573 VTAIL.n262 VTAIL.n218 1.93989
R1574 VTAIL.n38 VTAIL.n14 1.93989
R1575 VTAIL.n52 VTAIL.n8 1.93989
R1576 VTAIL.n196 VTAIL.n152 1.93989
R1577 VTAIL.n183 VTAIL.n159 1.93989
R1578 VTAIL.n126 VTAIL.n82 1.93989
R1579 VTAIL.n113 VTAIL.n89 1.93989
R1580 VTAIL.n75 VTAIL.n73 1.75912
R1581 VTAIL.n141 VTAIL.n75 1.75912
R1582 VTAIL.n145 VTAIL.n143 1.75912
R1583 VTAIL.n211 VTAIL.n145 1.75912
R1584 VTAIL.n71 VTAIL.n69 1.75912
R1585 VTAIL.n69 VTAIL.n67 1.75912
R1586 VTAIL.n279 VTAIL.n277 1.75912
R1587 VTAIL VTAIL.n1 1.37766
R1588 VTAIL.n143 VTAIL.n141 1.34964
R1589 VTAIL.n67 VTAIL.n1 1.34964
R1590 VTAIL.n253 VTAIL.n251 1.16414
R1591 VTAIL.n261 VTAIL.n220 1.16414
R1592 VTAIL.n43 VTAIL.n41 1.16414
R1593 VTAIL.n51 VTAIL.n10 1.16414
R1594 VTAIL.n195 VTAIL.n154 1.16414
R1595 VTAIL.n187 VTAIL.n186 1.16414
R1596 VTAIL.n125 VTAIL.n84 1.16414
R1597 VTAIL.n117 VTAIL.n116 1.16414
R1598 VTAIL.n252 VTAIL.n222 0.388379
R1599 VTAIL.n258 VTAIL.n257 0.388379
R1600 VTAIL.n42 VTAIL.n12 0.388379
R1601 VTAIL.n48 VTAIL.n47 0.388379
R1602 VTAIL.n192 VTAIL.n191 0.388379
R1603 VTAIL.n158 VTAIL.n156 0.388379
R1604 VTAIL.n122 VTAIL.n121 0.388379
R1605 VTAIL.n88 VTAIL.n86 0.388379
R1606 VTAIL VTAIL.n279 0.381966
R1607 VTAIL.n234 VTAIL.n229 0.155672
R1608 VTAIL.n241 VTAIL.n229 0.155672
R1609 VTAIL.n242 VTAIL.n241 0.155672
R1610 VTAIL.n242 VTAIL.n225 0.155672
R1611 VTAIL.n249 VTAIL.n225 0.155672
R1612 VTAIL.n250 VTAIL.n249 0.155672
R1613 VTAIL.n250 VTAIL.n221 0.155672
R1614 VTAIL.n259 VTAIL.n221 0.155672
R1615 VTAIL.n260 VTAIL.n259 0.155672
R1616 VTAIL.n260 VTAIL.n217 0.155672
R1617 VTAIL.n267 VTAIL.n217 0.155672
R1618 VTAIL.n268 VTAIL.n267 0.155672
R1619 VTAIL.n268 VTAIL.n213 0.155672
R1620 VTAIL.n275 VTAIL.n213 0.155672
R1621 VTAIL.n24 VTAIL.n19 0.155672
R1622 VTAIL.n31 VTAIL.n19 0.155672
R1623 VTAIL.n32 VTAIL.n31 0.155672
R1624 VTAIL.n32 VTAIL.n15 0.155672
R1625 VTAIL.n39 VTAIL.n15 0.155672
R1626 VTAIL.n40 VTAIL.n39 0.155672
R1627 VTAIL.n40 VTAIL.n11 0.155672
R1628 VTAIL.n49 VTAIL.n11 0.155672
R1629 VTAIL.n50 VTAIL.n49 0.155672
R1630 VTAIL.n50 VTAIL.n7 0.155672
R1631 VTAIL.n57 VTAIL.n7 0.155672
R1632 VTAIL.n58 VTAIL.n57 0.155672
R1633 VTAIL.n58 VTAIL.n3 0.155672
R1634 VTAIL.n65 VTAIL.n3 0.155672
R1635 VTAIL.n209 VTAIL.n147 0.155672
R1636 VTAIL.n202 VTAIL.n147 0.155672
R1637 VTAIL.n202 VTAIL.n201 0.155672
R1638 VTAIL.n201 VTAIL.n151 0.155672
R1639 VTAIL.n194 VTAIL.n151 0.155672
R1640 VTAIL.n194 VTAIL.n193 0.155672
R1641 VTAIL.n193 VTAIL.n155 0.155672
R1642 VTAIL.n185 VTAIL.n155 0.155672
R1643 VTAIL.n185 VTAIL.n184 0.155672
R1644 VTAIL.n184 VTAIL.n160 0.155672
R1645 VTAIL.n177 VTAIL.n160 0.155672
R1646 VTAIL.n177 VTAIL.n176 0.155672
R1647 VTAIL.n176 VTAIL.n164 0.155672
R1648 VTAIL.n169 VTAIL.n164 0.155672
R1649 VTAIL.n139 VTAIL.n77 0.155672
R1650 VTAIL.n132 VTAIL.n77 0.155672
R1651 VTAIL.n132 VTAIL.n131 0.155672
R1652 VTAIL.n131 VTAIL.n81 0.155672
R1653 VTAIL.n124 VTAIL.n81 0.155672
R1654 VTAIL.n124 VTAIL.n123 0.155672
R1655 VTAIL.n123 VTAIL.n85 0.155672
R1656 VTAIL.n115 VTAIL.n85 0.155672
R1657 VTAIL.n115 VTAIL.n114 0.155672
R1658 VTAIL.n114 VTAIL.n90 0.155672
R1659 VTAIL.n107 VTAIL.n90 0.155672
R1660 VTAIL.n107 VTAIL.n106 0.155672
R1661 VTAIL.n106 VTAIL.n94 0.155672
R1662 VTAIL.n99 VTAIL.n94 0.155672
R1663 VDD1.n60 VDD1.n0 756.745
R1664 VDD1.n127 VDD1.n67 756.745
R1665 VDD1.n61 VDD1.n60 585
R1666 VDD1.n59 VDD1.n58 585
R1667 VDD1.n4 VDD1.n3 585
R1668 VDD1.n53 VDD1.n52 585
R1669 VDD1.n51 VDD1.n50 585
R1670 VDD1.n8 VDD1.n7 585
R1671 VDD1.n45 VDD1.n44 585
R1672 VDD1.n43 VDD1.n10 585
R1673 VDD1.n42 VDD1.n41 585
R1674 VDD1.n13 VDD1.n11 585
R1675 VDD1.n36 VDD1.n35 585
R1676 VDD1.n34 VDD1.n33 585
R1677 VDD1.n17 VDD1.n16 585
R1678 VDD1.n28 VDD1.n27 585
R1679 VDD1.n26 VDD1.n25 585
R1680 VDD1.n21 VDD1.n20 585
R1681 VDD1.n87 VDD1.n86 585
R1682 VDD1.n92 VDD1.n91 585
R1683 VDD1.n94 VDD1.n93 585
R1684 VDD1.n83 VDD1.n82 585
R1685 VDD1.n100 VDD1.n99 585
R1686 VDD1.n102 VDD1.n101 585
R1687 VDD1.n79 VDD1.n78 585
R1688 VDD1.n109 VDD1.n108 585
R1689 VDD1.n110 VDD1.n77 585
R1690 VDD1.n112 VDD1.n111 585
R1691 VDD1.n75 VDD1.n74 585
R1692 VDD1.n118 VDD1.n117 585
R1693 VDD1.n120 VDD1.n119 585
R1694 VDD1.n71 VDD1.n70 585
R1695 VDD1.n126 VDD1.n125 585
R1696 VDD1.n128 VDD1.n127 585
R1697 VDD1.n22 VDD1.t1 329.036
R1698 VDD1.n88 VDD1.t5 329.036
R1699 VDD1.n60 VDD1.n59 171.744
R1700 VDD1.n59 VDD1.n3 171.744
R1701 VDD1.n52 VDD1.n3 171.744
R1702 VDD1.n52 VDD1.n51 171.744
R1703 VDD1.n51 VDD1.n7 171.744
R1704 VDD1.n44 VDD1.n7 171.744
R1705 VDD1.n44 VDD1.n43 171.744
R1706 VDD1.n43 VDD1.n42 171.744
R1707 VDD1.n42 VDD1.n11 171.744
R1708 VDD1.n35 VDD1.n11 171.744
R1709 VDD1.n35 VDD1.n34 171.744
R1710 VDD1.n34 VDD1.n16 171.744
R1711 VDD1.n27 VDD1.n16 171.744
R1712 VDD1.n27 VDD1.n26 171.744
R1713 VDD1.n26 VDD1.n20 171.744
R1714 VDD1.n92 VDD1.n86 171.744
R1715 VDD1.n93 VDD1.n92 171.744
R1716 VDD1.n93 VDD1.n82 171.744
R1717 VDD1.n100 VDD1.n82 171.744
R1718 VDD1.n101 VDD1.n100 171.744
R1719 VDD1.n101 VDD1.n78 171.744
R1720 VDD1.n109 VDD1.n78 171.744
R1721 VDD1.n110 VDD1.n109 171.744
R1722 VDD1.n111 VDD1.n110 171.744
R1723 VDD1.n111 VDD1.n74 171.744
R1724 VDD1.n118 VDD1.n74 171.744
R1725 VDD1.n119 VDD1.n118 171.744
R1726 VDD1.n119 VDD1.n70 171.744
R1727 VDD1.n126 VDD1.n70 171.744
R1728 VDD1.n127 VDD1.n126 171.744
R1729 VDD1.t1 VDD1.n20 85.8723
R1730 VDD1.t5 VDD1.n86 85.8723
R1731 VDD1.n135 VDD1.n134 74.9087
R1732 VDD1.n66 VDD1.n65 73.6453
R1733 VDD1.n137 VDD1.n136 73.6451
R1734 VDD1.n133 VDD1.n132 73.6451
R1735 VDD1.n66 VDD1.n64 50.4288
R1736 VDD1.n133 VDD1.n131 50.4288
R1737 VDD1.n137 VDD1.n135 43.9707
R1738 VDD1.n45 VDD1.n10 13.1884
R1739 VDD1.n112 VDD1.n77 13.1884
R1740 VDD1.n46 VDD1.n8 12.8005
R1741 VDD1.n41 VDD1.n12 12.8005
R1742 VDD1.n108 VDD1.n107 12.8005
R1743 VDD1.n113 VDD1.n75 12.8005
R1744 VDD1.n50 VDD1.n49 12.0247
R1745 VDD1.n40 VDD1.n13 12.0247
R1746 VDD1.n106 VDD1.n79 12.0247
R1747 VDD1.n117 VDD1.n116 12.0247
R1748 VDD1.n53 VDD1.n6 11.249
R1749 VDD1.n37 VDD1.n36 11.249
R1750 VDD1.n103 VDD1.n102 11.249
R1751 VDD1.n120 VDD1.n73 11.249
R1752 VDD1.n22 VDD1.n21 10.7239
R1753 VDD1.n88 VDD1.n87 10.7239
R1754 VDD1.n54 VDD1.n4 10.4732
R1755 VDD1.n33 VDD1.n15 10.4732
R1756 VDD1.n99 VDD1.n81 10.4732
R1757 VDD1.n121 VDD1.n71 10.4732
R1758 VDD1.n58 VDD1.n57 9.69747
R1759 VDD1.n32 VDD1.n17 9.69747
R1760 VDD1.n98 VDD1.n83 9.69747
R1761 VDD1.n125 VDD1.n124 9.69747
R1762 VDD1.n64 VDD1.n63 9.45567
R1763 VDD1.n131 VDD1.n130 9.45567
R1764 VDD1.n24 VDD1.n23 9.3005
R1765 VDD1.n19 VDD1.n18 9.3005
R1766 VDD1.n30 VDD1.n29 9.3005
R1767 VDD1.n32 VDD1.n31 9.3005
R1768 VDD1.n15 VDD1.n14 9.3005
R1769 VDD1.n38 VDD1.n37 9.3005
R1770 VDD1.n40 VDD1.n39 9.3005
R1771 VDD1.n12 VDD1.n9 9.3005
R1772 VDD1.n63 VDD1.n62 9.3005
R1773 VDD1.n2 VDD1.n1 9.3005
R1774 VDD1.n57 VDD1.n56 9.3005
R1775 VDD1.n55 VDD1.n54 9.3005
R1776 VDD1.n6 VDD1.n5 9.3005
R1777 VDD1.n49 VDD1.n48 9.3005
R1778 VDD1.n47 VDD1.n46 9.3005
R1779 VDD1.n130 VDD1.n129 9.3005
R1780 VDD1.n69 VDD1.n68 9.3005
R1781 VDD1.n124 VDD1.n123 9.3005
R1782 VDD1.n122 VDD1.n121 9.3005
R1783 VDD1.n73 VDD1.n72 9.3005
R1784 VDD1.n116 VDD1.n115 9.3005
R1785 VDD1.n114 VDD1.n113 9.3005
R1786 VDD1.n90 VDD1.n89 9.3005
R1787 VDD1.n85 VDD1.n84 9.3005
R1788 VDD1.n96 VDD1.n95 9.3005
R1789 VDD1.n98 VDD1.n97 9.3005
R1790 VDD1.n81 VDD1.n80 9.3005
R1791 VDD1.n104 VDD1.n103 9.3005
R1792 VDD1.n106 VDD1.n105 9.3005
R1793 VDD1.n107 VDD1.n76 9.3005
R1794 VDD1.n61 VDD1.n2 8.92171
R1795 VDD1.n29 VDD1.n28 8.92171
R1796 VDD1.n95 VDD1.n94 8.92171
R1797 VDD1.n128 VDD1.n69 8.92171
R1798 VDD1.n62 VDD1.n0 8.14595
R1799 VDD1.n25 VDD1.n19 8.14595
R1800 VDD1.n91 VDD1.n85 8.14595
R1801 VDD1.n129 VDD1.n67 8.14595
R1802 VDD1.n24 VDD1.n21 7.3702
R1803 VDD1.n90 VDD1.n87 7.3702
R1804 VDD1.n64 VDD1.n0 5.81868
R1805 VDD1.n25 VDD1.n24 5.81868
R1806 VDD1.n91 VDD1.n90 5.81868
R1807 VDD1.n131 VDD1.n67 5.81868
R1808 VDD1.n62 VDD1.n61 5.04292
R1809 VDD1.n28 VDD1.n19 5.04292
R1810 VDD1.n94 VDD1.n85 5.04292
R1811 VDD1.n129 VDD1.n128 5.04292
R1812 VDD1.n58 VDD1.n2 4.26717
R1813 VDD1.n29 VDD1.n17 4.26717
R1814 VDD1.n95 VDD1.n83 4.26717
R1815 VDD1.n125 VDD1.n69 4.26717
R1816 VDD1.n57 VDD1.n4 3.49141
R1817 VDD1.n33 VDD1.n32 3.49141
R1818 VDD1.n99 VDD1.n98 3.49141
R1819 VDD1.n124 VDD1.n71 3.49141
R1820 VDD1.n54 VDD1.n53 2.71565
R1821 VDD1.n36 VDD1.n15 2.71565
R1822 VDD1.n102 VDD1.n81 2.71565
R1823 VDD1.n121 VDD1.n120 2.71565
R1824 VDD1.n136 VDD1.t4 2.68465
R1825 VDD1.n136 VDD1.t8 2.68465
R1826 VDD1.n65 VDD1.t0 2.68465
R1827 VDD1.n65 VDD1.t9 2.68465
R1828 VDD1.n134 VDD1.t6 2.68465
R1829 VDD1.n134 VDD1.t7 2.68465
R1830 VDD1.n132 VDD1.t3 2.68465
R1831 VDD1.n132 VDD1.t2 2.68465
R1832 VDD1.n23 VDD1.n22 2.41282
R1833 VDD1.n89 VDD1.n88 2.41282
R1834 VDD1.n50 VDD1.n6 1.93989
R1835 VDD1.n37 VDD1.n13 1.93989
R1836 VDD1.n103 VDD1.n79 1.93989
R1837 VDD1.n117 VDD1.n73 1.93989
R1838 VDD1 VDD1.n137 1.26128
R1839 VDD1.n49 VDD1.n8 1.16414
R1840 VDD1.n41 VDD1.n40 1.16414
R1841 VDD1.n108 VDD1.n106 1.16414
R1842 VDD1.n116 VDD1.n75 1.16414
R1843 VDD1 VDD1.n66 0.498345
R1844 VDD1.n46 VDD1.n45 0.388379
R1845 VDD1.n12 VDD1.n10 0.388379
R1846 VDD1.n107 VDD1.n77 0.388379
R1847 VDD1.n113 VDD1.n112 0.388379
R1848 VDD1.n135 VDD1.n133 0.384809
R1849 VDD1.n63 VDD1.n1 0.155672
R1850 VDD1.n56 VDD1.n1 0.155672
R1851 VDD1.n56 VDD1.n55 0.155672
R1852 VDD1.n55 VDD1.n5 0.155672
R1853 VDD1.n48 VDD1.n5 0.155672
R1854 VDD1.n48 VDD1.n47 0.155672
R1855 VDD1.n47 VDD1.n9 0.155672
R1856 VDD1.n39 VDD1.n9 0.155672
R1857 VDD1.n39 VDD1.n38 0.155672
R1858 VDD1.n38 VDD1.n14 0.155672
R1859 VDD1.n31 VDD1.n14 0.155672
R1860 VDD1.n31 VDD1.n30 0.155672
R1861 VDD1.n30 VDD1.n18 0.155672
R1862 VDD1.n23 VDD1.n18 0.155672
R1863 VDD1.n89 VDD1.n84 0.155672
R1864 VDD1.n96 VDD1.n84 0.155672
R1865 VDD1.n97 VDD1.n96 0.155672
R1866 VDD1.n97 VDD1.n80 0.155672
R1867 VDD1.n104 VDD1.n80 0.155672
R1868 VDD1.n105 VDD1.n104 0.155672
R1869 VDD1.n105 VDD1.n76 0.155672
R1870 VDD1.n114 VDD1.n76 0.155672
R1871 VDD1.n115 VDD1.n114 0.155672
R1872 VDD1.n115 VDD1.n72 0.155672
R1873 VDD1.n122 VDD1.n72 0.155672
R1874 VDD1.n123 VDD1.n122 0.155672
R1875 VDD1.n123 VDD1.n68 0.155672
R1876 VDD1.n130 VDD1.n68 0.155672
R1877 VN.n7 VN.t9 200.415
R1878 VN.n38 VN.t4 200.415
R1879 VN.n30 VN.n29 181.852
R1880 VN.n61 VN.n60 181.852
R1881 VN.n15 VN.t1 170.673
R1882 VN.n8 VN.t8 170.673
R1883 VN.n22 VN.t5 170.673
R1884 VN.n29 VN.t3 170.673
R1885 VN.n46 VN.t7 170.673
R1886 VN.n39 VN.t6 170.673
R1887 VN.n53 VN.t0 170.673
R1888 VN.n60 VN.t2 170.673
R1889 VN.n59 VN.n31 161.3
R1890 VN.n58 VN.n57 161.3
R1891 VN.n56 VN.n32 161.3
R1892 VN.n55 VN.n54 161.3
R1893 VN.n52 VN.n33 161.3
R1894 VN.n51 VN.n50 161.3
R1895 VN.n49 VN.n34 161.3
R1896 VN.n48 VN.n47 161.3
R1897 VN.n46 VN.n35 161.3
R1898 VN.n45 VN.n44 161.3
R1899 VN.n43 VN.n36 161.3
R1900 VN.n42 VN.n41 161.3
R1901 VN.n40 VN.n37 161.3
R1902 VN.n28 VN.n0 161.3
R1903 VN.n27 VN.n26 161.3
R1904 VN.n25 VN.n1 161.3
R1905 VN.n24 VN.n23 161.3
R1906 VN.n21 VN.n2 161.3
R1907 VN.n20 VN.n19 161.3
R1908 VN.n18 VN.n3 161.3
R1909 VN.n17 VN.n16 161.3
R1910 VN.n15 VN.n4 161.3
R1911 VN.n14 VN.n13 161.3
R1912 VN.n12 VN.n5 161.3
R1913 VN.n11 VN.n10 161.3
R1914 VN.n9 VN.n6 161.3
R1915 VN.n8 VN.n7 66.2588
R1916 VN.n39 VN.n38 66.2588
R1917 VN VN.n61 48.6236
R1918 VN.n27 VN.n1 46.321
R1919 VN.n58 VN.n32 46.321
R1920 VN.n10 VN.n5 42.4359
R1921 VN.n20 VN.n3 42.4359
R1922 VN.n41 VN.n36 42.4359
R1923 VN.n51 VN.n34 42.4359
R1924 VN.n14 VN.n5 38.5509
R1925 VN.n16 VN.n3 38.5509
R1926 VN.n45 VN.n36 38.5509
R1927 VN.n47 VN.n34 38.5509
R1928 VN.n23 VN.n1 34.6658
R1929 VN.n54 VN.n32 34.6658
R1930 VN.n10 VN.n9 24.4675
R1931 VN.n15 VN.n14 24.4675
R1932 VN.n16 VN.n15 24.4675
R1933 VN.n21 VN.n20 24.4675
R1934 VN.n28 VN.n27 24.4675
R1935 VN.n41 VN.n40 24.4675
R1936 VN.n47 VN.n46 24.4675
R1937 VN.n46 VN.n45 24.4675
R1938 VN.n52 VN.n51 24.4675
R1939 VN.n59 VN.n58 24.4675
R1940 VN.n23 VN.n22 22.5101
R1941 VN.n54 VN.n53 22.5101
R1942 VN.n38 VN.n37 18.5717
R1943 VN.n7 VN.n6 18.5717
R1944 VN.n29 VN.n28 3.91522
R1945 VN.n60 VN.n59 3.91522
R1946 VN.n9 VN.n8 1.95786
R1947 VN.n22 VN.n21 1.95786
R1948 VN.n40 VN.n39 1.95786
R1949 VN.n53 VN.n52 1.95786
R1950 VN.n61 VN.n31 0.189894
R1951 VN.n57 VN.n31 0.189894
R1952 VN.n57 VN.n56 0.189894
R1953 VN.n56 VN.n55 0.189894
R1954 VN.n55 VN.n33 0.189894
R1955 VN.n50 VN.n33 0.189894
R1956 VN.n50 VN.n49 0.189894
R1957 VN.n49 VN.n48 0.189894
R1958 VN.n48 VN.n35 0.189894
R1959 VN.n44 VN.n35 0.189894
R1960 VN.n44 VN.n43 0.189894
R1961 VN.n43 VN.n42 0.189894
R1962 VN.n42 VN.n37 0.189894
R1963 VN.n11 VN.n6 0.189894
R1964 VN.n12 VN.n11 0.189894
R1965 VN.n13 VN.n12 0.189894
R1966 VN.n13 VN.n4 0.189894
R1967 VN.n17 VN.n4 0.189894
R1968 VN.n18 VN.n17 0.189894
R1969 VN.n19 VN.n18 0.189894
R1970 VN.n19 VN.n2 0.189894
R1971 VN.n24 VN.n2 0.189894
R1972 VN.n25 VN.n24 0.189894
R1973 VN.n26 VN.n25 0.189894
R1974 VN.n26 VN.n0 0.189894
R1975 VN.n30 VN.n0 0.189894
R1976 VN VN.n30 0.0516364
R1977 VDD2.n129 VDD2.n69 756.745
R1978 VDD2.n60 VDD2.n0 756.745
R1979 VDD2.n130 VDD2.n129 585
R1980 VDD2.n128 VDD2.n127 585
R1981 VDD2.n73 VDD2.n72 585
R1982 VDD2.n122 VDD2.n121 585
R1983 VDD2.n120 VDD2.n119 585
R1984 VDD2.n77 VDD2.n76 585
R1985 VDD2.n114 VDD2.n113 585
R1986 VDD2.n112 VDD2.n79 585
R1987 VDD2.n111 VDD2.n110 585
R1988 VDD2.n82 VDD2.n80 585
R1989 VDD2.n105 VDD2.n104 585
R1990 VDD2.n103 VDD2.n102 585
R1991 VDD2.n86 VDD2.n85 585
R1992 VDD2.n97 VDD2.n96 585
R1993 VDD2.n95 VDD2.n94 585
R1994 VDD2.n90 VDD2.n89 585
R1995 VDD2.n20 VDD2.n19 585
R1996 VDD2.n25 VDD2.n24 585
R1997 VDD2.n27 VDD2.n26 585
R1998 VDD2.n16 VDD2.n15 585
R1999 VDD2.n33 VDD2.n32 585
R2000 VDD2.n35 VDD2.n34 585
R2001 VDD2.n12 VDD2.n11 585
R2002 VDD2.n42 VDD2.n41 585
R2003 VDD2.n43 VDD2.n10 585
R2004 VDD2.n45 VDD2.n44 585
R2005 VDD2.n8 VDD2.n7 585
R2006 VDD2.n51 VDD2.n50 585
R2007 VDD2.n53 VDD2.n52 585
R2008 VDD2.n4 VDD2.n3 585
R2009 VDD2.n59 VDD2.n58 585
R2010 VDD2.n61 VDD2.n60 585
R2011 VDD2.n91 VDD2.t7 329.036
R2012 VDD2.n21 VDD2.t0 329.036
R2013 VDD2.n129 VDD2.n128 171.744
R2014 VDD2.n128 VDD2.n72 171.744
R2015 VDD2.n121 VDD2.n72 171.744
R2016 VDD2.n121 VDD2.n120 171.744
R2017 VDD2.n120 VDD2.n76 171.744
R2018 VDD2.n113 VDD2.n76 171.744
R2019 VDD2.n113 VDD2.n112 171.744
R2020 VDD2.n112 VDD2.n111 171.744
R2021 VDD2.n111 VDD2.n80 171.744
R2022 VDD2.n104 VDD2.n80 171.744
R2023 VDD2.n104 VDD2.n103 171.744
R2024 VDD2.n103 VDD2.n85 171.744
R2025 VDD2.n96 VDD2.n85 171.744
R2026 VDD2.n96 VDD2.n95 171.744
R2027 VDD2.n95 VDD2.n89 171.744
R2028 VDD2.n25 VDD2.n19 171.744
R2029 VDD2.n26 VDD2.n25 171.744
R2030 VDD2.n26 VDD2.n15 171.744
R2031 VDD2.n33 VDD2.n15 171.744
R2032 VDD2.n34 VDD2.n33 171.744
R2033 VDD2.n34 VDD2.n11 171.744
R2034 VDD2.n42 VDD2.n11 171.744
R2035 VDD2.n43 VDD2.n42 171.744
R2036 VDD2.n44 VDD2.n43 171.744
R2037 VDD2.n44 VDD2.n7 171.744
R2038 VDD2.n51 VDD2.n7 171.744
R2039 VDD2.n52 VDD2.n51 171.744
R2040 VDD2.n52 VDD2.n3 171.744
R2041 VDD2.n59 VDD2.n3 171.744
R2042 VDD2.n60 VDD2.n59 171.744
R2043 VDD2.t7 VDD2.n89 85.8723
R2044 VDD2.t0 VDD2.n19 85.8723
R2045 VDD2.n68 VDD2.n67 74.9087
R2046 VDD2 VDD2.n137 74.9059
R2047 VDD2.n136 VDD2.n135 73.6453
R2048 VDD2.n66 VDD2.n65 73.6451
R2049 VDD2.n66 VDD2.n64 50.4288
R2050 VDD2.n134 VDD2.n133 48.6702
R2051 VDD2.n134 VDD2.n68 42.5084
R2052 VDD2.n114 VDD2.n79 13.1884
R2053 VDD2.n45 VDD2.n10 13.1884
R2054 VDD2.n115 VDD2.n77 12.8005
R2055 VDD2.n110 VDD2.n81 12.8005
R2056 VDD2.n41 VDD2.n40 12.8005
R2057 VDD2.n46 VDD2.n8 12.8005
R2058 VDD2.n119 VDD2.n118 12.0247
R2059 VDD2.n109 VDD2.n82 12.0247
R2060 VDD2.n39 VDD2.n12 12.0247
R2061 VDD2.n50 VDD2.n49 12.0247
R2062 VDD2.n122 VDD2.n75 11.249
R2063 VDD2.n106 VDD2.n105 11.249
R2064 VDD2.n36 VDD2.n35 11.249
R2065 VDD2.n53 VDD2.n6 11.249
R2066 VDD2.n91 VDD2.n90 10.7239
R2067 VDD2.n21 VDD2.n20 10.7239
R2068 VDD2.n123 VDD2.n73 10.4732
R2069 VDD2.n102 VDD2.n84 10.4732
R2070 VDD2.n32 VDD2.n14 10.4732
R2071 VDD2.n54 VDD2.n4 10.4732
R2072 VDD2.n127 VDD2.n126 9.69747
R2073 VDD2.n101 VDD2.n86 9.69747
R2074 VDD2.n31 VDD2.n16 9.69747
R2075 VDD2.n58 VDD2.n57 9.69747
R2076 VDD2.n133 VDD2.n132 9.45567
R2077 VDD2.n64 VDD2.n63 9.45567
R2078 VDD2.n93 VDD2.n92 9.3005
R2079 VDD2.n88 VDD2.n87 9.3005
R2080 VDD2.n99 VDD2.n98 9.3005
R2081 VDD2.n101 VDD2.n100 9.3005
R2082 VDD2.n84 VDD2.n83 9.3005
R2083 VDD2.n107 VDD2.n106 9.3005
R2084 VDD2.n109 VDD2.n108 9.3005
R2085 VDD2.n81 VDD2.n78 9.3005
R2086 VDD2.n132 VDD2.n131 9.3005
R2087 VDD2.n71 VDD2.n70 9.3005
R2088 VDD2.n126 VDD2.n125 9.3005
R2089 VDD2.n124 VDD2.n123 9.3005
R2090 VDD2.n75 VDD2.n74 9.3005
R2091 VDD2.n118 VDD2.n117 9.3005
R2092 VDD2.n116 VDD2.n115 9.3005
R2093 VDD2.n63 VDD2.n62 9.3005
R2094 VDD2.n2 VDD2.n1 9.3005
R2095 VDD2.n57 VDD2.n56 9.3005
R2096 VDD2.n55 VDD2.n54 9.3005
R2097 VDD2.n6 VDD2.n5 9.3005
R2098 VDD2.n49 VDD2.n48 9.3005
R2099 VDD2.n47 VDD2.n46 9.3005
R2100 VDD2.n23 VDD2.n22 9.3005
R2101 VDD2.n18 VDD2.n17 9.3005
R2102 VDD2.n29 VDD2.n28 9.3005
R2103 VDD2.n31 VDD2.n30 9.3005
R2104 VDD2.n14 VDD2.n13 9.3005
R2105 VDD2.n37 VDD2.n36 9.3005
R2106 VDD2.n39 VDD2.n38 9.3005
R2107 VDD2.n40 VDD2.n9 9.3005
R2108 VDD2.n130 VDD2.n71 8.92171
R2109 VDD2.n98 VDD2.n97 8.92171
R2110 VDD2.n28 VDD2.n27 8.92171
R2111 VDD2.n61 VDD2.n2 8.92171
R2112 VDD2.n131 VDD2.n69 8.14595
R2113 VDD2.n94 VDD2.n88 8.14595
R2114 VDD2.n24 VDD2.n18 8.14595
R2115 VDD2.n62 VDD2.n0 8.14595
R2116 VDD2.n93 VDD2.n90 7.3702
R2117 VDD2.n23 VDD2.n20 7.3702
R2118 VDD2.n133 VDD2.n69 5.81868
R2119 VDD2.n94 VDD2.n93 5.81868
R2120 VDD2.n24 VDD2.n23 5.81868
R2121 VDD2.n64 VDD2.n0 5.81868
R2122 VDD2.n131 VDD2.n130 5.04292
R2123 VDD2.n97 VDD2.n88 5.04292
R2124 VDD2.n27 VDD2.n18 5.04292
R2125 VDD2.n62 VDD2.n61 5.04292
R2126 VDD2.n127 VDD2.n71 4.26717
R2127 VDD2.n98 VDD2.n86 4.26717
R2128 VDD2.n28 VDD2.n16 4.26717
R2129 VDD2.n58 VDD2.n2 4.26717
R2130 VDD2.n126 VDD2.n73 3.49141
R2131 VDD2.n102 VDD2.n101 3.49141
R2132 VDD2.n32 VDD2.n31 3.49141
R2133 VDD2.n57 VDD2.n4 3.49141
R2134 VDD2.n123 VDD2.n122 2.71565
R2135 VDD2.n105 VDD2.n84 2.71565
R2136 VDD2.n35 VDD2.n14 2.71565
R2137 VDD2.n54 VDD2.n53 2.71565
R2138 VDD2.n137 VDD2.t3 2.68465
R2139 VDD2.n137 VDD2.t5 2.68465
R2140 VDD2.n135 VDD2.t9 2.68465
R2141 VDD2.n135 VDD2.t2 2.68465
R2142 VDD2.n67 VDD2.t4 2.68465
R2143 VDD2.n67 VDD2.t6 2.68465
R2144 VDD2.n65 VDD2.t1 2.68465
R2145 VDD2.n65 VDD2.t8 2.68465
R2146 VDD2.n92 VDD2.n91 2.41282
R2147 VDD2.n22 VDD2.n21 2.41282
R2148 VDD2.n119 VDD2.n75 1.93989
R2149 VDD2.n106 VDD2.n82 1.93989
R2150 VDD2.n36 VDD2.n12 1.93989
R2151 VDD2.n50 VDD2.n6 1.93989
R2152 VDD2.n136 VDD2.n134 1.75912
R2153 VDD2.n118 VDD2.n77 1.16414
R2154 VDD2.n110 VDD2.n109 1.16414
R2155 VDD2.n41 VDD2.n39 1.16414
R2156 VDD2.n49 VDD2.n8 1.16414
R2157 VDD2 VDD2.n136 0.498345
R2158 VDD2.n115 VDD2.n114 0.388379
R2159 VDD2.n81 VDD2.n79 0.388379
R2160 VDD2.n40 VDD2.n10 0.388379
R2161 VDD2.n46 VDD2.n45 0.388379
R2162 VDD2.n68 VDD2.n66 0.384809
R2163 VDD2.n132 VDD2.n70 0.155672
R2164 VDD2.n125 VDD2.n70 0.155672
R2165 VDD2.n125 VDD2.n124 0.155672
R2166 VDD2.n124 VDD2.n74 0.155672
R2167 VDD2.n117 VDD2.n74 0.155672
R2168 VDD2.n117 VDD2.n116 0.155672
R2169 VDD2.n116 VDD2.n78 0.155672
R2170 VDD2.n108 VDD2.n78 0.155672
R2171 VDD2.n108 VDD2.n107 0.155672
R2172 VDD2.n107 VDD2.n83 0.155672
R2173 VDD2.n100 VDD2.n83 0.155672
R2174 VDD2.n100 VDD2.n99 0.155672
R2175 VDD2.n99 VDD2.n87 0.155672
R2176 VDD2.n92 VDD2.n87 0.155672
R2177 VDD2.n22 VDD2.n17 0.155672
R2178 VDD2.n29 VDD2.n17 0.155672
R2179 VDD2.n30 VDD2.n29 0.155672
R2180 VDD2.n30 VDD2.n13 0.155672
R2181 VDD2.n37 VDD2.n13 0.155672
R2182 VDD2.n38 VDD2.n37 0.155672
R2183 VDD2.n38 VDD2.n9 0.155672
R2184 VDD2.n47 VDD2.n9 0.155672
R2185 VDD2.n48 VDD2.n47 0.155672
R2186 VDD2.n48 VDD2.n5 0.155672
R2187 VDD2.n55 VDD2.n5 0.155672
R2188 VDD2.n56 VDD2.n55 0.155672
R2189 VDD2.n56 VDD2.n1 0.155672
R2190 VDD2.n63 VDD2.n1 0.155672
C0 w_n3418_n3390# VDD1 2.45201f
C1 B VP 1.79695f
C2 VP w_n3418_n3390# 7.492471f
C3 VP VDD1 10.040999f
C4 B VDD2 2.21856f
C5 B VTAIL 3.3466f
C6 w_n3418_n3390# VDD2 2.54941f
C7 w_n3418_n3390# VTAIL 3.10697f
C8 VDD1 VDD2 1.5934f
C9 VTAIL VDD1 10.717f
C10 VP VDD2 0.469815f
C11 VP VTAIL 10.0041f
C12 B VN 1.05818f
C13 VTAIL VDD2 10.7606f
C14 w_n3418_n3390# VN 7.05021f
C15 VN VDD1 0.15101f
C16 VP VN 7.10728f
C17 VN VDD2 9.72626f
C18 VN VTAIL 9.98974f
C19 B w_n3418_n3390# 9.08087f
C20 B VDD1 2.13531f
C21 VDD2 VSUBS 1.814292f
C22 VDD1 VSUBS 1.591292f
C23 VTAIL VSUBS 1.080834f
C24 VN VSUBS 6.24882f
C25 VP VSUBS 3.090647f
C26 B VSUBS 4.271712f
C27 w_n3418_n3390# VSUBS 0.142613p
C28 VDD2.n0 VSUBS 0.029963f
C29 VDD2.n1 VSUBS 0.02748f
C30 VDD2.n2 VSUBS 0.014767f
C31 VDD2.n3 VSUBS 0.034903f
C32 VDD2.n4 VSUBS 0.015635f
C33 VDD2.n5 VSUBS 0.02748f
C34 VDD2.n6 VSUBS 0.014767f
C35 VDD2.n7 VSUBS 0.034903f
C36 VDD2.n8 VSUBS 0.015635f
C37 VDD2.n9 VSUBS 0.02748f
C38 VDD2.n10 VSUBS 0.015201f
C39 VDD2.n11 VSUBS 0.034903f
C40 VDD2.n12 VSUBS 0.015635f
C41 VDD2.n13 VSUBS 0.02748f
C42 VDD2.n14 VSUBS 0.014767f
C43 VDD2.n15 VSUBS 0.034903f
C44 VDD2.n16 VSUBS 0.015635f
C45 VDD2.n17 VSUBS 0.02748f
C46 VDD2.n18 VSUBS 0.014767f
C47 VDD2.n19 VSUBS 0.026177f
C48 VDD2.n20 VSUBS 0.026256f
C49 VDD2.t0 VSUBS 0.075223f
C50 VDD2.n21 VSUBS 0.21779f
C51 VDD2.n22 VSUBS 1.36344f
C52 VDD2.n23 VSUBS 0.014767f
C53 VDD2.n24 VSUBS 0.015635f
C54 VDD2.n25 VSUBS 0.034903f
C55 VDD2.n26 VSUBS 0.034903f
C56 VDD2.n27 VSUBS 0.015635f
C57 VDD2.n28 VSUBS 0.014767f
C58 VDD2.n29 VSUBS 0.02748f
C59 VDD2.n30 VSUBS 0.02748f
C60 VDD2.n31 VSUBS 0.014767f
C61 VDD2.n32 VSUBS 0.015635f
C62 VDD2.n33 VSUBS 0.034903f
C63 VDD2.n34 VSUBS 0.034903f
C64 VDD2.n35 VSUBS 0.015635f
C65 VDD2.n36 VSUBS 0.014767f
C66 VDD2.n37 VSUBS 0.02748f
C67 VDD2.n38 VSUBS 0.02748f
C68 VDD2.n39 VSUBS 0.014767f
C69 VDD2.n40 VSUBS 0.014767f
C70 VDD2.n41 VSUBS 0.015635f
C71 VDD2.n42 VSUBS 0.034903f
C72 VDD2.n43 VSUBS 0.034903f
C73 VDD2.n44 VSUBS 0.034903f
C74 VDD2.n45 VSUBS 0.015201f
C75 VDD2.n46 VSUBS 0.014767f
C76 VDD2.n47 VSUBS 0.02748f
C77 VDD2.n48 VSUBS 0.02748f
C78 VDD2.n49 VSUBS 0.014767f
C79 VDD2.n50 VSUBS 0.015635f
C80 VDD2.n51 VSUBS 0.034903f
C81 VDD2.n52 VSUBS 0.034903f
C82 VDD2.n53 VSUBS 0.015635f
C83 VDD2.n54 VSUBS 0.014767f
C84 VDD2.n55 VSUBS 0.02748f
C85 VDD2.n56 VSUBS 0.02748f
C86 VDD2.n57 VSUBS 0.014767f
C87 VDD2.n58 VSUBS 0.015635f
C88 VDD2.n59 VSUBS 0.034903f
C89 VDD2.n60 VSUBS 0.083708f
C90 VDD2.n61 VSUBS 0.015635f
C91 VDD2.n62 VSUBS 0.014767f
C92 VDD2.n63 VSUBS 0.063144f
C93 VDD2.n64 VSUBS 0.068296f
C94 VDD2.t1 VSUBS 0.262977f
C95 VDD2.t8 VSUBS 0.262977f
C96 VDD2.n65 VSUBS 2.05399f
C97 VDD2.n66 VSUBS 0.910767f
C98 VDD2.t4 VSUBS 0.262977f
C99 VDD2.t6 VSUBS 0.262977f
C100 VDD2.n67 VSUBS 2.06744f
C101 VDD2.n68 VSUBS 2.97664f
C102 VDD2.n69 VSUBS 0.029963f
C103 VDD2.n70 VSUBS 0.02748f
C104 VDD2.n71 VSUBS 0.014767f
C105 VDD2.n72 VSUBS 0.034903f
C106 VDD2.n73 VSUBS 0.015635f
C107 VDD2.n74 VSUBS 0.02748f
C108 VDD2.n75 VSUBS 0.014767f
C109 VDD2.n76 VSUBS 0.034903f
C110 VDD2.n77 VSUBS 0.015635f
C111 VDD2.n78 VSUBS 0.02748f
C112 VDD2.n79 VSUBS 0.015201f
C113 VDD2.n80 VSUBS 0.034903f
C114 VDD2.n81 VSUBS 0.014767f
C115 VDD2.n82 VSUBS 0.015635f
C116 VDD2.n83 VSUBS 0.02748f
C117 VDD2.n84 VSUBS 0.014767f
C118 VDD2.n85 VSUBS 0.034903f
C119 VDD2.n86 VSUBS 0.015635f
C120 VDD2.n87 VSUBS 0.02748f
C121 VDD2.n88 VSUBS 0.014767f
C122 VDD2.n89 VSUBS 0.026177f
C123 VDD2.n90 VSUBS 0.026256f
C124 VDD2.t7 VSUBS 0.075223f
C125 VDD2.n91 VSUBS 0.21779f
C126 VDD2.n92 VSUBS 1.36344f
C127 VDD2.n93 VSUBS 0.014767f
C128 VDD2.n94 VSUBS 0.015635f
C129 VDD2.n95 VSUBS 0.034903f
C130 VDD2.n96 VSUBS 0.034903f
C131 VDD2.n97 VSUBS 0.015635f
C132 VDD2.n98 VSUBS 0.014767f
C133 VDD2.n99 VSUBS 0.02748f
C134 VDD2.n100 VSUBS 0.02748f
C135 VDD2.n101 VSUBS 0.014767f
C136 VDD2.n102 VSUBS 0.015635f
C137 VDD2.n103 VSUBS 0.034903f
C138 VDD2.n104 VSUBS 0.034903f
C139 VDD2.n105 VSUBS 0.015635f
C140 VDD2.n106 VSUBS 0.014767f
C141 VDD2.n107 VSUBS 0.02748f
C142 VDD2.n108 VSUBS 0.02748f
C143 VDD2.n109 VSUBS 0.014767f
C144 VDD2.n110 VSUBS 0.015635f
C145 VDD2.n111 VSUBS 0.034903f
C146 VDD2.n112 VSUBS 0.034903f
C147 VDD2.n113 VSUBS 0.034903f
C148 VDD2.n114 VSUBS 0.015201f
C149 VDD2.n115 VSUBS 0.014767f
C150 VDD2.n116 VSUBS 0.02748f
C151 VDD2.n117 VSUBS 0.02748f
C152 VDD2.n118 VSUBS 0.014767f
C153 VDD2.n119 VSUBS 0.015635f
C154 VDD2.n120 VSUBS 0.034903f
C155 VDD2.n121 VSUBS 0.034903f
C156 VDD2.n122 VSUBS 0.015635f
C157 VDD2.n123 VSUBS 0.014767f
C158 VDD2.n124 VSUBS 0.02748f
C159 VDD2.n125 VSUBS 0.02748f
C160 VDD2.n126 VSUBS 0.014767f
C161 VDD2.n127 VSUBS 0.015635f
C162 VDD2.n128 VSUBS 0.034903f
C163 VDD2.n129 VSUBS 0.083708f
C164 VDD2.n130 VSUBS 0.015635f
C165 VDD2.n131 VSUBS 0.014767f
C166 VDD2.n132 VSUBS 0.063144f
C167 VDD2.n133 VSUBS 0.061027f
C168 VDD2.n134 VSUBS 2.80619f
C169 VDD2.t9 VSUBS 0.262977f
C170 VDD2.t2 VSUBS 0.262977f
C171 VDD2.n135 VSUBS 2.054f
C172 VDD2.n136 VSUBS 0.717999f
C173 VDD2.t3 VSUBS 0.262977f
C174 VDD2.t5 VSUBS 0.262977f
C175 VDD2.n137 VSUBS 2.0674f
C176 VN.n0 VSUBS 0.035076f
C177 VN.t3 VSUBS 1.97953f
C178 VN.n1 VSUBS 0.030011f
C179 VN.n2 VSUBS 0.035076f
C180 VN.t5 VSUBS 1.97953f
C181 VN.n3 VSUBS 0.028536f
C182 VN.n4 VSUBS 0.035076f
C183 VN.t1 VSUBS 1.97953f
C184 VN.n5 VSUBS 0.028536f
C185 VN.n6 VSUBS 0.224302f
C186 VN.t8 VSUBS 1.97953f
C187 VN.t9 VSUBS 2.10712f
C188 VN.n7 VSUBS 0.803725f
C189 VN.n8 VSUBS 0.771974f
C190 VN.n9 VSUBS 0.035679f
C191 VN.n10 VSUBS 0.068922f
C192 VN.n11 VSUBS 0.035076f
C193 VN.n12 VSUBS 0.035076f
C194 VN.n13 VSUBS 0.035076f
C195 VN.n14 VSUBS 0.070321f
C196 VN.n15 VSUBS 0.743892f
C197 VN.n16 VSUBS 0.070321f
C198 VN.n17 VSUBS 0.035076f
C199 VN.n18 VSUBS 0.035076f
C200 VN.n19 VSUBS 0.035076f
C201 VN.n20 VSUBS 0.068922f
C202 VN.n21 VSUBS 0.035679f
C203 VN.n22 VSUBS 0.710795f
C204 VN.n23 VSUBS 0.068295f
C205 VN.n24 VSUBS 0.035076f
C206 VN.n25 VSUBS 0.035076f
C207 VN.n26 VSUBS 0.035076f
C208 VN.n27 VSUBS 0.066892f
C209 VN.n28 VSUBS 0.038261f
C210 VN.n29 VSUBS 0.785382f
C211 VN.n30 VSUBS 0.036686f
C212 VN.n31 VSUBS 0.035076f
C213 VN.t2 VSUBS 1.97953f
C214 VN.n32 VSUBS 0.030011f
C215 VN.n33 VSUBS 0.035076f
C216 VN.t0 VSUBS 1.97953f
C217 VN.n34 VSUBS 0.028536f
C218 VN.n35 VSUBS 0.035076f
C219 VN.t7 VSUBS 1.97953f
C220 VN.n36 VSUBS 0.028536f
C221 VN.n37 VSUBS 0.224302f
C222 VN.t6 VSUBS 1.97953f
C223 VN.t4 VSUBS 2.10712f
C224 VN.n38 VSUBS 0.803725f
C225 VN.n39 VSUBS 0.771974f
C226 VN.n40 VSUBS 0.035679f
C227 VN.n41 VSUBS 0.068922f
C228 VN.n42 VSUBS 0.035076f
C229 VN.n43 VSUBS 0.035076f
C230 VN.n44 VSUBS 0.035076f
C231 VN.n45 VSUBS 0.070321f
C232 VN.n46 VSUBS 0.743892f
C233 VN.n47 VSUBS 0.070321f
C234 VN.n48 VSUBS 0.035076f
C235 VN.n49 VSUBS 0.035076f
C236 VN.n50 VSUBS 0.035076f
C237 VN.n51 VSUBS 0.068922f
C238 VN.n52 VSUBS 0.035679f
C239 VN.n53 VSUBS 0.710795f
C240 VN.n54 VSUBS 0.068295f
C241 VN.n55 VSUBS 0.035076f
C242 VN.n56 VSUBS 0.035076f
C243 VN.n57 VSUBS 0.035076f
C244 VN.n58 VSUBS 0.066892f
C245 VN.n59 VSUBS 0.038261f
C246 VN.n60 VSUBS 0.785382f
C247 VN.n61 VSUBS 1.83851f
C248 VDD1.n0 VSUBS 0.029962f
C249 VDD1.n1 VSUBS 0.027479f
C250 VDD1.n2 VSUBS 0.014766f
C251 VDD1.n3 VSUBS 0.034901f
C252 VDD1.n4 VSUBS 0.015634f
C253 VDD1.n5 VSUBS 0.027479f
C254 VDD1.n6 VSUBS 0.014766f
C255 VDD1.n7 VSUBS 0.034901f
C256 VDD1.n8 VSUBS 0.015634f
C257 VDD1.n9 VSUBS 0.027479f
C258 VDD1.n10 VSUBS 0.0152f
C259 VDD1.n11 VSUBS 0.034901f
C260 VDD1.n12 VSUBS 0.014766f
C261 VDD1.n13 VSUBS 0.015634f
C262 VDD1.n14 VSUBS 0.027479f
C263 VDD1.n15 VSUBS 0.014766f
C264 VDD1.n16 VSUBS 0.034901f
C265 VDD1.n17 VSUBS 0.015634f
C266 VDD1.n18 VSUBS 0.027479f
C267 VDD1.n19 VSUBS 0.014766f
C268 VDD1.n20 VSUBS 0.026176f
C269 VDD1.n21 VSUBS 0.026254f
C270 VDD1.t1 VSUBS 0.075218f
C271 VDD1.n22 VSUBS 0.217777f
C272 VDD1.n23 VSUBS 1.36336f
C273 VDD1.n24 VSUBS 0.014766f
C274 VDD1.n25 VSUBS 0.015634f
C275 VDD1.n26 VSUBS 0.034901f
C276 VDD1.n27 VSUBS 0.034901f
C277 VDD1.n28 VSUBS 0.015634f
C278 VDD1.n29 VSUBS 0.014766f
C279 VDD1.n30 VSUBS 0.027479f
C280 VDD1.n31 VSUBS 0.027479f
C281 VDD1.n32 VSUBS 0.014766f
C282 VDD1.n33 VSUBS 0.015634f
C283 VDD1.n34 VSUBS 0.034901f
C284 VDD1.n35 VSUBS 0.034901f
C285 VDD1.n36 VSUBS 0.015634f
C286 VDD1.n37 VSUBS 0.014766f
C287 VDD1.n38 VSUBS 0.027479f
C288 VDD1.n39 VSUBS 0.027479f
C289 VDD1.n40 VSUBS 0.014766f
C290 VDD1.n41 VSUBS 0.015634f
C291 VDD1.n42 VSUBS 0.034901f
C292 VDD1.n43 VSUBS 0.034901f
C293 VDD1.n44 VSUBS 0.034901f
C294 VDD1.n45 VSUBS 0.0152f
C295 VDD1.n46 VSUBS 0.014766f
C296 VDD1.n47 VSUBS 0.027479f
C297 VDD1.n48 VSUBS 0.027479f
C298 VDD1.n49 VSUBS 0.014766f
C299 VDD1.n50 VSUBS 0.015634f
C300 VDD1.n51 VSUBS 0.034901f
C301 VDD1.n52 VSUBS 0.034901f
C302 VDD1.n53 VSUBS 0.015634f
C303 VDD1.n54 VSUBS 0.014766f
C304 VDD1.n55 VSUBS 0.027479f
C305 VDD1.n56 VSUBS 0.027479f
C306 VDD1.n57 VSUBS 0.014766f
C307 VDD1.n58 VSUBS 0.015634f
C308 VDD1.n59 VSUBS 0.034901f
C309 VDD1.n60 VSUBS 0.083703f
C310 VDD1.n61 VSUBS 0.015634f
C311 VDD1.n62 VSUBS 0.014766f
C312 VDD1.n63 VSUBS 0.06314f
C313 VDD1.n64 VSUBS 0.068291f
C314 VDD1.t0 VSUBS 0.262962f
C315 VDD1.t9 VSUBS 0.262962f
C316 VDD1.n65 VSUBS 2.05388f
C317 VDD1.n66 VSUBS 0.919098f
C318 VDD1.n67 VSUBS 0.029962f
C319 VDD1.n68 VSUBS 0.027479f
C320 VDD1.n69 VSUBS 0.014766f
C321 VDD1.n70 VSUBS 0.034901f
C322 VDD1.n71 VSUBS 0.015634f
C323 VDD1.n72 VSUBS 0.027479f
C324 VDD1.n73 VSUBS 0.014766f
C325 VDD1.n74 VSUBS 0.034901f
C326 VDD1.n75 VSUBS 0.015634f
C327 VDD1.n76 VSUBS 0.027479f
C328 VDD1.n77 VSUBS 0.0152f
C329 VDD1.n78 VSUBS 0.034901f
C330 VDD1.n79 VSUBS 0.015634f
C331 VDD1.n80 VSUBS 0.027479f
C332 VDD1.n81 VSUBS 0.014766f
C333 VDD1.n82 VSUBS 0.034901f
C334 VDD1.n83 VSUBS 0.015634f
C335 VDD1.n84 VSUBS 0.027479f
C336 VDD1.n85 VSUBS 0.014766f
C337 VDD1.n86 VSUBS 0.026176f
C338 VDD1.n87 VSUBS 0.026254f
C339 VDD1.t5 VSUBS 0.075218f
C340 VDD1.n88 VSUBS 0.217777f
C341 VDD1.n89 VSUBS 1.36336f
C342 VDD1.n90 VSUBS 0.014766f
C343 VDD1.n91 VSUBS 0.015634f
C344 VDD1.n92 VSUBS 0.034901f
C345 VDD1.n93 VSUBS 0.034901f
C346 VDD1.n94 VSUBS 0.015634f
C347 VDD1.n95 VSUBS 0.014766f
C348 VDD1.n96 VSUBS 0.027479f
C349 VDD1.n97 VSUBS 0.027479f
C350 VDD1.n98 VSUBS 0.014766f
C351 VDD1.n99 VSUBS 0.015634f
C352 VDD1.n100 VSUBS 0.034901f
C353 VDD1.n101 VSUBS 0.034901f
C354 VDD1.n102 VSUBS 0.015634f
C355 VDD1.n103 VSUBS 0.014766f
C356 VDD1.n104 VSUBS 0.027479f
C357 VDD1.n105 VSUBS 0.027479f
C358 VDD1.n106 VSUBS 0.014766f
C359 VDD1.n107 VSUBS 0.014766f
C360 VDD1.n108 VSUBS 0.015634f
C361 VDD1.n109 VSUBS 0.034901f
C362 VDD1.n110 VSUBS 0.034901f
C363 VDD1.n111 VSUBS 0.034901f
C364 VDD1.n112 VSUBS 0.0152f
C365 VDD1.n113 VSUBS 0.014766f
C366 VDD1.n114 VSUBS 0.027479f
C367 VDD1.n115 VSUBS 0.027479f
C368 VDD1.n116 VSUBS 0.014766f
C369 VDD1.n117 VSUBS 0.015634f
C370 VDD1.n118 VSUBS 0.034901f
C371 VDD1.n119 VSUBS 0.034901f
C372 VDD1.n120 VSUBS 0.015634f
C373 VDD1.n121 VSUBS 0.014766f
C374 VDD1.n122 VSUBS 0.027479f
C375 VDD1.n123 VSUBS 0.027479f
C376 VDD1.n124 VSUBS 0.014766f
C377 VDD1.n125 VSUBS 0.015634f
C378 VDD1.n126 VSUBS 0.034901f
C379 VDD1.n127 VSUBS 0.083703f
C380 VDD1.n128 VSUBS 0.015634f
C381 VDD1.n129 VSUBS 0.014766f
C382 VDD1.n130 VSUBS 0.06314f
C383 VDD1.n131 VSUBS 0.068291f
C384 VDD1.t3 VSUBS 0.262962f
C385 VDD1.t2 VSUBS 0.262962f
C386 VDD1.n132 VSUBS 2.05387f
C387 VDD1.n133 VSUBS 0.910713f
C388 VDD1.t6 VSUBS 0.262962f
C389 VDD1.t7 VSUBS 0.262962f
C390 VDD1.n134 VSUBS 2.06732f
C391 VDD1.n135 VSUBS 3.08836f
C392 VDD1.t4 VSUBS 0.262962f
C393 VDD1.t8 VSUBS 0.262962f
C394 VDD1.n136 VSUBS 2.05387f
C395 VDD1.n137 VSUBS 3.38379f
C396 VTAIL.t4 VSUBS 0.270377f
C397 VTAIL.t2 VSUBS 0.270377f
C398 VTAIL.n0 VSUBS 1.95737f
C399 VTAIL.n1 VSUBS 0.897f
C400 VTAIL.n2 VSUBS 0.030807f
C401 VTAIL.n3 VSUBS 0.028253f
C402 VTAIL.n4 VSUBS 0.015182f
C403 VTAIL.n5 VSUBS 0.035885f
C404 VTAIL.n6 VSUBS 0.016075f
C405 VTAIL.n7 VSUBS 0.028253f
C406 VTAIL.n8 VSUBS 0.015182f
C407 VTAIL.n9 VSUBS 0.035885f
C408 VTAIL.n10 VSUBS 0.016075f
C409 VTAIL.n11 VSUBS 0.028253f
C410 VTAIL.n12 VSUBS 0.015629f
C411 VTAIL.n13 VSUBS 0.035885f
C412 VTAIL.n14 VSUBS 0.016075f
C413 VTAIL.n15 VSUBS 0.028253f
C414 VTAIL.n16 VSUBS 0.015182f
C415 VTAIL.n17 VSUBS 0.035885f
C416 VTAIL.n18 VSUBS 0.016075f
C417 VTAIL.n19 VSUBS 0.028253f
C418 VTAIL.n20 VSUBS 0.015182f
C419 VTAIL.n21 VSUBS 0.026914f
C420 VTAIL.n22 VSUBS 0.026995f
C421 VTAIL.t12 VSUBS 0.077339f
C422 VTAIL.n23 VSUBS 0.223918f
C423 VTAIL.n24 VSUBS 1.4018f
C424 VTAIL.n25 VSUBS 0.015182f
C425 VTAIL.n26 VSUBS 0.016075f
C426 VTAIL.n27 VSUBS 0.035885f
C427 VTAIL.n28 VSUBS 0.035885f
C428 VTAIL.n29 VSUBS 0.016075f
C429 VTAIL.n30 VSUBS 0.015182f
C430 VTAIL.n31 VSUBS 0.028253f
C431 VTAIL.n32 VSUBS 0.028253f
C432 VTAIL.n33 VSUBS 0.015182f
C433 VTAIL.n34 VSUBS 0.016075f
C434 VTAIL.n35 VSUBS 0.035885f
C435 VTAIL.n36 VSUBS 0.035885f
C436 VTAIL.n37 VSUBS 0.016075f
C437 VTAIL.n38 VSUBS 0.015182f
C438 VTAIL.n39 VSUBS 0.028253f
C439 VTAIL.n40 VSUBS 0.028253f
C440 VTAIL.n41 VSUBS 0.015182f
C441 VTAIL.n42 VSUBS 0.015182f
C442 VTAIL.n43 VSUBS 0.016075f
C443 VTAIL.n44 VSUBS 0.035885f
C444 VTAIL.n45 VSUBS 0.035885f
C445 VTAIL.n46 VSUBS 0.035885f
C446 VTAIL.n47 VSUBS 0.015629f
C447 VTAIL.n48 VSUBS 0.015182f
C448 VTAIL.n49 VSUBS 0.028253f
C449 VTAIL.n50 VSUBS 0.028253f
C450 VTAIL.n51 VSUBS 0.015182f
C451 VTAIL.n52 VSUBS 0.016075f
C452 VTAIL.n53 VSUBS 0.035885f
C453 VTAIL.n54 VSUBS 0.035885f
C454 VTAIL.n55 VSUBS 0.016075f
C455 VTAIL.n56 VSUBS 0.015182f
C456 VTAIL.n57 VSUBS 0.028253f
C457 VTAIL.n58 VSUBS 0.028253f
C458 VTAIL.n59 VSUBS 0.015182f
C459 VTAIL.n60 VSUBS 0.016075f
C460 VTAIL.n61 VSUBS 0.035885f
C461 VTAIL.n62 VSUBS 0.086064f
C462 VTAIL.n63 VSUBS 0.016075f
C463 VTAIL.n64 VSUBS 0.015182f
C464 VTAIL.n65 VSUBS 0.064921f
C465 VTAIL.n66 VSUBS 0.043233f
C466 VTAIL.n67 VSUBS 0.30684f
C467 VTAIL.t18 VSUBS 0.270377f
C468 VTAIL.t11 VSUBS 0.270377f
C469 VTAIL.n68 VSUBS 1.95737f
C470 VTAIL.n69 VSUBS 0.969007f
C471 VTAIL.t16 VSUBS 0.270377f
C472 VTAIL.t17 VSUBS 0.270377f
C473 VTAIL.n70 VSUBS 1.95737f
C474 VTAIL.n71 VSUBS 2.46332f
C475 VTAIL.t8 VSUBS 0.270377f
C476 VTAIL.t9 VSUBS 0.270377f
C477 VTAIL.n72 VSUBS 1.95738f
C478 VTAIL.n73 VSUBS 2.4633f
C479 VTAIL.t5 VSUBS 0.270377f
C480 VTAIL.t0 VSUBS 0.270377f
C481 VTAIL.n74 VSUBS 1.95738f
C482 VTAIL.n75 VSUBS 0.968993f
C483 VTAIL.n76 VSUBS 0.030807f
C484 VTAIL.n77 VSUBS 0.028253f
C485 VTAIL.n78 VSUBS 0.015182f
C486 VTAIL.n79 VSUBS 0.035885f
C487 VTAIL.n80 VSUBS 0.016075f
C488 VTAIL.n81 VSUBS 0.028253f
C489 VTAIL.n82 VSUBS 0.015182f
C490 VTAIL.n83 VSUBS 0.035885f
C491 VTAIL.n84 VSUBS 0.016075f
C492 VTAIL.n85 VSUBS 0.028253f
C493 VTAIL.n86 VSUBS 0.015629f
C494 VTAIL.n87 VSUBS 0.035885f
C495 VTAIL.n88 VSUBS 0.015182f
C496 VTAIL.n89 VSUBS 0.016075f
C497 VTAIL.n90 VSUBS 0.028253f
C498 VTAIL.n91 VSUBS 0.015182f
C499 VTAIL.n92 VSUBS 0.035885f
C500 VTAIL.n93 VSUBS 0.016075f
C501 VTAIL.n94 VSUBS 0.028253f
C502 VTAIL.n95 VSUBS 0.015182f
C503 VTAIL.n96 VSUBS 0.026914f
C504 VTAIL.n97 VSUBS 0.026995f
C505 VTAIL.t7 VSUBS 0.077339f
C506 VTAIL.n98 VSUBS 0.223918f
C507 VTAIL.n99 VSUBS 1.4018f
C508 VTAIL.n100 VSUBS 0.015182f
C509 VTAIL.n101 VSUBS 0.016075f
C510 VTAIL.n102 VSUBS 0.035885f
C511 VTAIL.n103 VSUBS 0.035885f
C512 VTAIL.n104 VSUBS 0.016075f
C513 VTAIL.n105 VSUBS 0.015182f
C514 VTAIL.n106 VSUBS 0.028253f
C515 VTAIL.n107 VSUBS 0.028253f
C516 VTAIL.n108 VSUBS 0.015182f
C517 VTAIL.n109 VSUBS 0.016075f
C518 VTAIL.n110 VSUBS 0.035885f
C519 VTAIL.n111 VSUBS 0.035885f
C520 VTAIL.n112 VSUBS 0.016075f
C521 VTAIL.n113 VSUBS 0.015182f
C522 VTAIL.n114 VSUBS 0.028253f
C523 VTAIL.n115 VSUBS 0.028253f
C524 VTAIL.n116 VSUBS 0.015182f
C525 VTAIL.n117 VSUBS 0.016075f
C526 VTAIL.n118 VSUBS 0.035885f
C527 VTAIL.n119 VSUBS 0.035885f
C528 VTAIL.n120 VSUBS 0.035885f
C529 VTAIL.n121 VSUBS 0.015629f
C530 VTAIL.n122 VSUBS 0.015182f
C531 VTAIL.n123 VSUBS 0.028253f
C532 VTAIL.n124 VSUBS 0.028253f
C533 VTAIL.n125 VSUBS 0.015182f
C534 VTAIL.n126 VSUBS 0.016075f
C535 VTAIL.n127 VSUBS 0.035885f
C536 VTAIL.n128 VSUBS 0.035885f
C537 VTAIL.n129 VSUBS 0.016075f
C538 VTAIL.n130 VSUBS 0.015182f
C539 VTAIL.n131 VSUBS 0.028253f
C540 VTAIL.n132 VSUBS 0.028253f
C541 VTAIL.n133 VSUBS 0.015182f
C542 VTAIL.n134 VSUBS 0.016075f
C543 VTAIL.n135 VSUBS 0.035885f
C544 VTAIL.n136 VSUBS 0.086064f
C545 VTAIL.n137 VSUBS 0.016075f
C546 VTAIL.n138 VSUBS 0.015182f
C547 VTAIL.n139 VSUBS 0.064921f
C548 VTAIL.n140 VSUBS 0.043233f
C549 VTAIL.n141 VSUBS 0.30684f
C550 VTAIL.t15 VSUBS 0.270377f
C551 VTAIL.t10 VSUBS 0.270377f
C552 VTAIL.n142 VSUBS 1.95738f
C553 VTAIL.n143 VSUBS 0.931714f
C554 VTAIL.t13 VSUBS 0.270377f
C555 VTAIL.t19 VSUBS 0.270377f
C556 VTAIL.n144 VSUBS 1.95738f
C557 VTAIL.n145 VSUBS 0.968993f
C558 VTAIL.n146 VSUBS 0.030807f
C559 VTAIL.n147 VSUBS 0.028253f
C560 VTAIL.n148 VSUBS 0.015182f
C561 VTAIL.n149 VSUBS 0.035885f
C562 VTAIL.n150 VSUBS 0.016075f
C563 VTAIL.n151 VSUBS 0.028253f
C564 VTAIL.n152 VSUBS 0.015182f
C565 VTAIL.n153 VSUBS 0.035885f
C566 VTAIL.n154 VSUBS 0.016075f
C567 VTAIL.n155 VSUBS 0.028253f
C568 VTAIL.n156 VSUBS 0.015629f
C569 VTAIL.n157 VSUBS 0.035885f
C570 VTAIL.n158 VSUBS 0.015182f
C571 VTAIL.n159 VSUBS 0.016075f
C572 VTAIL.n160 VSUBS 0.028253f
C573 VTAIL.n161 VSUBS 0.015182f
C574 VTAIL.n162 VSUBS 0.035885f
C575 VTAIL.n163 VSUBS 0.016075f
C576 VTAIL.n164 VSUBS 0.028253f
C577 VTAIL.n165 VSUBS 0.015182f
C578 VTAIL.n166 VSUBS 0.026914f
C579 VTAIL.n167 VSUBS 0.026995f
C580 VTAIL.t14 VSUBS 0.077339f
C581 VTAIL.n168 VSUBS 0.223918f
C582 VTAIL.n169 VSUBS 1.4018f
C583 VTAIL.n170 VSUBS 0.015182f
C584 VTAIL.n171 VSUBS 0.016075f
C585 VTAIL.n172 VSUBS 0.035885f
C586 VTAIL.n173 VSUBS 0.035885f
C587 VTAIL.n174 VSUBS 0.016075f
C588 VTAIL.n175 VSUBS 0.015182f
C589 VTAIL.n176 VSUBS 0.028253f
C590 VTAIL.n177 VSUBS 0.028253f
C591 VTAIL.n178 VSUBS 0.015182f
C592 VTAIL.n179 VSUBS 0.016075f
C593 VTAIL.n180 VSUBS 0.035885f
C594 VTAIL.n181 VSUBS 0.035885f
C595 VTAIL.n182 VSUBS 0.016075f
C596 VTAIL.n183 VSUBS 0.015182f
C597 VTAIL.n184 VSUBS 0.028253f
C598 VTAIL.n185 VSUBS 0.028253f
C599 VTAIL.n186 VSUBS 0.015182f
C600 VTAIL.n187 VSUBS 0.016075f
C601 VTAIL.n188 VSUBS 0.035885f
C602 VTAIL.n189 VSUBS 0.035885f
C603 VTAIL.n190 VSUBS 0.035885f
C604 VTAIL.n191 VSUBS 0.015629f
C605 VTAIL.n192 VSUBS 0.015182f
C606 VTAIL.n193 VSUBS 0.028253f
C607 VTAIL.n194 VSUBS 0.028253f
C608 VTAIL.n195 VSUBS 0.015182f
C609 VTAIL.n196 VSUBS 0.016075f
C610 VTAIL.n197 VSUBS 0.035885f
C611 VTAIL.n198 VSUBS 0.035885f
C612 VTAIL.n199 VSUBS 0.016075f
C613 VTAIL.n200 VSUBS 0.015182f
C614 VTAIL.n201 VSUBS 0.028253f
C615 VTAIL.n202 VSUBS 0.028253f
C616 VTAIL.n203 VSUBS 0.015182f
C617 VTAIL.n204 VSUBS 0.016075f
C618 VTAIL.n205 VSUBS 0.035885f
C619 VTAIL.n206 VSUBS 0.086064f
C620 VTAIL.n207 VSUBS 0.016075f
C621 VTAIL.n208 VSUBS 0.015182f
C622 VTAIL.n209 VSUBS 0.064921f
C623 VTAIL.n210 VSUBS 0.043233f
C624 VTAIL.n211 VSUBS 1.67832f
C625 VTAIL.n212 VSUBS 0.030807f
C626 VTAIL.n213 VSUBS 0.028253f
C627 VTAIL.n214 VSUBS 0.015182f
C628 VTAIL.n215 VSUBS 0.035885f
C629 VTAIL.n216 VSUBS 0.016075f
C630 VTAIL.n217 VSUBS 0.028253f
C631 VTAIL.n218 VSUBS 0.015182f
C632 VTAIL.n219 VSUBS 0.035885f
C633 VTAIL.n220 VSUBS 0.016075f
C634 VTAIL.n221 VSUBS 0.028253f
C635 VTAIL.n222 VSUBS 0.015629f
C636 VTAIL.n223 VSUBS 0.035885f
C637 VTAIL.n224 VSUBS 0.016075f
C638 VTAIL.n225 VSUBS 0.028253f
C639 VTAIL.n226 VSUBS 0.015182f
C640 VTAIL.n227 VSUBS 0.035885f
C641 VTAIL.n228 VSUBS 0.016075f
C642 VTAIL.n229 VSUBS 0.028253f
C643 VTAIL.n230 VSUBS 0.015182f
C644 VTAIL.n231 VSUBS 0.026914f
C645 VTAIL.n232 VSUBS 0.026995f
C646 VTAIL.t1 VSUBS 0.077339f
C647 VTAIL.n233 VSUBS 0.223918f
C648 VTAIL.n234 VSUBS 1.4018f
C649 VTAIL.n235 VSUBS 0.015182f
C650 VTAIL.n236 VSUBS 0.016075f
C651 VTAIL.n237 VSUBS 0.035885f
C652 VTAIL.n238 VSUBS 0.035885f
C653 VTAIL.n239 VSUBS 0.016075f
C654 VTAIL.n240 VSUBS 0.015182f
C655 VTAIL.n241 VSUBS 0.028253f
C656 VTAIL.n242 VSUBS 0.028253f
C657 VTAIL.n243 VSUBS 0.015182f
C658 VTAIL.n244 VSUBS 0.016075f
C659 VTAIL.n245 VSUBS 0.035885f
C660 VTAIL.n246 VSUBS 0.035885f
C661 VTAIL.n247 VSUBS 0.016075f
C662 VTAIL.n248 VSUBS 0.015182f
C663 VTAIL.n249 VSUBS 0.028253f
C664 VTAIL.n250 VSUBS 0.028253f
C665 VTAIL.n251 VSUBS 0.015182f
C666 VTAIL.n252 VSUBS 0.015182f
C667 VTAIL.n253 VSUBS 0.016075f
C668 VTAIL.n254 VSUBS 0.035885f
C669 VTAIL.n255 VSUBS 0.035885f
C670 VTAIL.n256 VSUBS 0.035885f
C671 VTAIL.n257 VSUBS 0.015629f
C672 VTAIL.n258 VSUBS 0.015182f
C673 VTAIL.n259 VSUBS 0.028253f
C674 VTAIL.n260 VSUBS 0.028253f
C675 VTAIL.n261 VSUBS 0.015182f
C676 VTAIL.n262 VSUBS 0.016075f
C677 VTAIL.n263 VSUBS 0.035885f
C678 VTAIL.n264 VSUBS 0.035885f
C679 VTAIL.n265 VSUBS 0.016075f
C680 VTAIL.n266 VSUBS 0.015182f
C681 VTAIL.n267 VSUBS 0.028253f
C682 VTAIL.n268 VSUBS 0.028253f
C683 VTAIL.n269 VSUBS 0.015182f
C684 VTAIL.n270 VSUBS 0.016075f
C685 VTAIL.n271 VSUBS 0.035885f
C686 VTAIL.n272 VSUBS 0.086064f
C687 VTAIL.n273 VSUBS 0.016075f
C688 VTAIL.n274 VSUBS 0.015182f
C689 VTAIL.n275 VSUBS 0.064921f
C690 VTAIL.n276 VSUBS 0.043233f
C691 VTAIL.n277 VSUBS 1.67832f
C692 VTAIL.t3 VSUBS 0.270377f
C693 VTAIL.t6 VSUBS 0.270377f
C694 VTAIL.n278 VSUBS 1.95737f
C695 VTAIL.n279 VSUBS 0.843632f
C696 VP.n0 VSUBS 0.035852f
C697 VP.t2 VSUBS 2.02335f
C698 VP.n1 VSUBS 0.030676f
C699 VP.n2 VSUBS 0.035852f
C700 VP.t3 VSUBS 2.02335f
C701 VP.n3 VSUBS 0.029167f
C702 VP.n4 VSUBS 0.035852f
C703 VP.t7 VSUBS 2.02335f
C704 VP.n5 VSUBS 0.029167f
C705 VP.n6 VSUBS 0.035852f
C706 VP.t6 VSUBS 2.02335f
C707 VP.n7 VSUBS 0.030676f
C708 VP.n8 VSUBS 0.035852f
C709 VP.t4 VSUBS 2.02335f
C710 VP.n9 VSUBS 0.035852f
C711 VP.t1 VSUBS 2.02335f
C712 VP.n10 VSUBS 0.030676f
C713 VP.n11 VSUBS 0.035852f
C714 VP.t5 VSUBS 2.02335f
C715 VP.n12 VSUBS 0.029167f
C716 VP.n13 VSUBS 0.035852f
C717 VP.t0 VSUBS 2.02335f
C718 VP.n14 VSUBS 0.029167f
C719 VP.n15 VSUBS 0.229267f
C720 VP.t9 VSUBS 2.02335f
C721 VP.t8 VSUBS 2.15377f
C722 VP.n16 VSUBS 0.821516f
C723 VP.n17 VSUBS 0.789062f
C724 VP.n18 VSUBS 0.036469f
C725 VP.n19 VSUBS 0.070448f
C726 VP.n20 VSUBS 0.035852f
C727 VP.n21 VSUBS 0.035852f
C728 VP.n22 VSUBS 0.035852f
C729 VP.n23 VSUBS 0.071878f
C730 VP.n24 VSUBS 0.760359f
C731 VP.n25 VSUBS 0.071878f
C732 VP.n26 VSUBS 0.035852f
C733 VP.n27 VSUBS 0.035852f
C734 VP.n28 VSUBS 0.035852f
C735 VP.n29 VSUBS 0.070448f
C736 VP.n30 VSUBS 0.036469f
C737 VP.n31 VSUBS 0.726529f
C738 VP.n32 VSUBS 0.069806f
C739 VP.n33 VSUBS 0.035852f
C740 VP.n34 VSUBS 0.035852f
C741 VP.n35 VSUBS 0.035852f
C742 VP.n36 VSUBS 0.068372f
C743 VP.n37 VSUBS 0.039108f
C744 VP.n38 VSUBS 0.802767f
C745 VP.n39 VSUBS 1.85586f
C746 VP.n40 VSUBS 1.88258f
C747 VP.n41 VSUBS 0.802767f
C748 VP.n42 VSUBS 0.039108f
C749 VP.n43 VSUBS 0.068372f
C750 VP.n44 VSUBS 0.035852f
C751 VP.n45 VSUBS 0.035852f
C752 VP.n46 VSUBS 0.035852f
C753 VP.n47 VSUBS 0.069806f
C754 VP.n48 VSUBS 0.726529f
C755 VP.n49 VSUBS 0.036469f
C756 VP.n50 VSUBS 0.070448f
C757 VP.n51 VSUBS 0.035852f
C758 VP.n52 VSUBS 0.035852f
C759 VP.n53 VSUBS 0.035852f
C760 VP.n54 VSUBS 0.071878f
C761 VP.n55 VSUBS 0.760359f
C762 VP.n56 VSUBS 0.071878f
C763 VP.n57 VSUBS 0.035852f
C764 VP.n58 VSUBS 0.035852f
C765 VP.n59 VSUBS 0.035852f
C766 VP.n60 VSUBS 0.070448f
C767 VP.n61 VSUBS 0.036469f
C768 VP.n62 VSUBS 0.726529f
C769 VP.n63 VSUBS 0.069806f
C770 VP.n64 VSUBS 0.035852f
C771 VP.n65 VSUBS 0.035852f
C772 VP.n66 VSUBS 0.035852f
C773 VP.n67 VSUBS 0.068372f
C774 VP.n68 VSUBS 0.039108f
C775 VP.n69 VSUBS 0.802767f
C776 VP.n70 VSUBS 0.037498f
C777 B.n0 VSUBS 0.005583f
C778 B.n1 VSUBS 0.005583f
C779 B.n2 VSUBS 0.008828f
C780 B.n3 VSUBS 0.008828f
C781 B.n4 VSUBS 0.008828f
C782 B.n5 VSUBS 0.008828f
C783 B.n6 VSUBS 0.008828f
C784 B.n7 VSUBS 0.008828f
C785 B.n8 VSUBS 0.008828f
C786 B.n9 VSUBS 0.008828f
C787 B.n10 VSUBS 0.008828f
C788 B.n11 VSUBS 0.008828f
C789 B.n12 VSUBS 0.008828f
C790 B.n13 VSUBS 0.008828f
C791 B.n14 VSUBS 0.008828f
C792 B.n15 VSUBS 0.008828f
C793 B.n16 VSUBS 0.008828f
C794 B.n17 VSUBS 0.008828f
C795 B.n18 VSUBS 0.008828f
C796 B.n19 VSUBS 0.008828f
C797 B.n20 VSUBS 0.008828f
C798 B.n21 VSUBS 0.008828f
C799 B.n22 VSUBS 0.008828f
C800 B.n23 VSUBS 0.008828f
C801 B.n24 VSUBS 0.022428f
C802 B.n25 VSUBS 0.008828f
C803 B.n26 VSUBS 0.008828f
C804 B.n27 VSUBS 0.008828f
C805 B.n28 VSUBS 0.008828f
C806 B.n29 VSUBS 0.008828f
C807 B.n30 VSUBS 0.008828f
C808 B.n31 VSUBS 0.008828f
C809 B.n32 VSUBS 0.008828f
C810 B.n33 VSUBS 0.008828f
C811 B.n34 VSUBS 0.008828f
C812 B.n35 VSUBS 0.008828f
C813 B.n36 VSUBS 0.008828f
C814 B.n37 VSUBS 0.008828f
C815 B.n38 VSUBS 0.008828f
C816 B.n39 VSUBS 0.008828f
C817 B.n40 VSUBS 0.008828f
C818 B.n41 VSUBS 0.008828f
C819 B.n42 VSUBS 0.008828f
C820 B.n43 VSUBS 0.008828f
C821 B.n44 VSUBS 0.008828f
C822 B.n45 VSUBS 0.008828f
C823 B.t8 VSUBS 0.2693f
C824 B.t7 VSUBS 0.297958f
C825 B.t6 VSUBS 1.15322f
C826 B.n46 VSUBS 0.460003f
C827 B.n47 VSUBS 0.314812f
C828 B.n48 VSUBS 0.008828f
C829 B.n49 VSUBS 0.008828f
C830 B.n50 VSUBS 0.008828f
C831 B.n51 VSUBS 0.008828f
C832 B.t5 VSUBS 0.269304f
C833 B.t4 VSUBS 0.297961f
C834 B.t3 VSUBS 1.15322f
C835 B.n52 VSUBS 0.459999f
C836 B.n53 VSUBS 0.314808f
C837 B.n54 VSUBS 0.008828f
C838 B.n55 VSUBS 0.008828f
C839 B.n56 VSUBS 0.008828f
C840 B.n57 VSUBS 0.008828f
C841 B.n58 VSUBS 0.008828f
C842 B.n59 VSUBS 0.008828f
C843 B.n60 VSUBS 0.008828f
C844 B.n61 VSUBS 0.008828f
C845 B.n62 VSUBS 0.008828f
C846 B.n63 VSUBS 0.008828f
C847 B.n64 VSUBS 0.008828f
C848 B.n65 VSUBS 0.008828f
C849 B.n66 VSUBS 0.008828f
C850 B.n67 VSUBS 0.008828f
C851 B.n68 VSUBS 0.008828f
C852 B.n69 VSUBS 0.008828f
C853 B.n70 VSUBS 0.008828f
C854 B.n71 VSUBS 0.008828f
C855 B.n72 VSUBS 0.008828f
C856 B.n73 VSUBS 0.008828f
C857 B.n74 VSUBS 0.021483f
C858 B.n75 VSUBS 0.008828f
C859 B.n76 VSUBS 0.008828f
C860 B.n77 VSUBS 0.008828f
C861 B.n78 VSUBS 0.008828f
C862 B.n79 VSUBS 0.008828f
C863 B.n80 VSUBS 0.008828f
C864 B.n81 VSUBS 0.008828f
C865 B.n82 VSUBS 0.008828f
C866 B.n83 VSUBS 0.008828f
C867 B.n84 VSUBS 0.008828f
C868 B.n85 VSUBS 0.008828f
C869 B.n86 VSUBS 0.008828f
C870 B.n87 VSUBS 0.008828f
C871 B.n88 VSUBS 0.008828f
C872 B.n89 VSUBS 0.008828f
C873 B.n90 VSUBS 0.008828f
C874 B.n91 VSUBS 0.008828f
C875 B.n92 VSUBS 0.008828f
C876 B.n93 VSUBS 0.008828f
C877 B.n94 VSUBS 0.008828f
C878 B.n95 VSUBS 0.008828f
C879 B.n96 VSUBS 0.008828f
C880 B.n97 VSUBS 0.008828f
C881 B.n98 VSUBS 0.008828f
C882 B.n99 VSUBS 0.008828f
C883 B.n100 VSUBS 0.008828f
C884 B.n101 VSUBS 0.008828f
C885 B.n102 VSUBS 0.008828f
C886 B.n103 VSUBS 0.008828f
C887 B.n104 VSUBS 0.008828f
C888 B.n105 VSUBS 0.008828f
C889 B.n106 VSUBS 0.008828f
C890 B.n107 VSUBS 0.008828f
C891 B.n108 VSUBS 0.008828f
C892 B.n109 VSUBS 0.008828f
C893 B.n110 VSUBS 0.008828f
C894 B.n111 VSUBS 0.008828f
C895 B.n112 VSUBS 0.008828f
C896 B.n113 VSUBS 0.008828f
C897 B.n114 VSUBS 0.008828f
C898 B.n115 VSUBS 0.008828f
C899 B.n116 VSUBS 0.008828f
C900 B.n117 VSUBS 0.008828f
C901 B.n118 VSUBS 0.008828f
C902 B.n119 VSUBS 0.022428f
C903 B.n120 VSUBS 0.008828f
C904 B.n121 VSUBS 0.008828f
C905 B.n122 VSUBS 0.008828f
C906 B.n123 VSUBS 0.008828f
C907 B.n124 VSUBS 0.008828f
C908 B.n125 VSUBS 0.008828f
C909 B.n126 VSUBS 0.008828f
C910 B.n127 VSUBS 0.008828f
C911 B.n128 VSUBS 0.008828f
C912 B.n129 VSUBS 0.008828f
C913 B.n130 VSUBS 0.008828f
C914 B.n131 VSUBS 0.008828f
C915 B.n132 VSUBS 0.008828f
C916 B.n133 VSUBS 0.008828f
C917 B.n134 VSUBS 0.008828f
C918 B.n135 VSUBS 0.008828f
C919 B.n136 VSUBS 0.008828f
C920 B.n137 VSUBS 0.008828f
C921 B.n138 VSUBS 0.008828f
C922 B.n139 VSUBS 0.008828f
C923 B.t1 VSUBS 0.269304f
C924 B.t2 VSUBS 0.297961f
C925 B.t0 VSUBS 1.15322f
C926 B.n140 VSUBS 0.459999f
C927 B.n141 VSUBS 0.314808f
C928 B.n142 VSUBS 0.020454f
C929 B.n143 VSUBS 0.008828f
C930 B.n144 VSUBS 0.008828f
C931 B.n145 VSUBS 0.008828f
C932 B.n146 VSUBS 0.008828f
C933 B.n147 VSUBS 0.008828f
C934 B.t10 VSUBS 0.2693f
C935 B.t11 VSUBS 0.297958f
C936 B.t9 VSUBS 1.15322f
C937 B.n148 VSUBS 0.460003f
C938 B.n149 VSUBS 0.314812f
C939 B.n150 VSUBS 0.008828f
C940 B.n151 VSUBS 0.008828f
C941 B.n152 VSUBS 0.008828f
C942 B.n153 VSUBS 0.008828f
C943 B.n154 VSUBS 0.008828f
C944 B.n155 VSUBS 0.008828f
C945 B.n156 VSUBS 0.008828f
C946 B.n157 VSUBS 0.008828f
C947 B.n158 VSUBS 0.008828f
C948 B.n159 VSUBS 0.008828f
C949 B.n160 VSUBS 0.008828f
C950 B.n161 VSUBS 0.008828f
C951 B.n162 VSUBS 0.008828f
C952 B.n163 VSUBS 0.008828f
C953 B.n164 VSUBS 0.008828f
C954 B.n165 VSUBS 0.008828f
C955 B.n166 VSUBS 0.008828f
C956 B.n167 VSUBS 0.008828f
C957 B.n168 VSUBS 0.008828f
C958 B.n169 VSUBS 0.008828f
C959 B.n170 VSUBS 0.021713f
C960 B.n171 VSUBS 0.008828f
C961 B.n172 VSUBS 0.008828f
C962 B.n173 VSUBS 0.008828f
C963 B.n174 VSUBS 0.008828f
C964 B.n175 VSUBS 0.008828f
C965 B.n176 VSUBS 0.008828f
C966 B.n177 VSUBS 0.008828f
C967 B.n178 VSUBS 0.008828f
C968 B.n179 VSUBS 0.008828f
C969 B.n180 VSUBS 0.008828f
C970 B.n181 VSUBS 0.008828f
C971 B.n182 VSUBS 0.008828f
C972 B.n183 VSUBS 0.008828f
C973 B.n184 VSUBS 0.008828f
C974 B.n185 VSUBS 0.008828f
C975 B.n186 VSUBS 0.008828f
C976 B.n187 VSUBS 0.008828f
C977 B.n188 VSUBS 0.008828f
C978 B.n189 VSUBS 0.008828f
C979 B.n190 VSUBS 0.008828f
C980 B.n191 VSUBS 0.008828f
C981 B.n192 VSUBS 0.008828f
C982 B.n193 VSUBS 0.008828f
C983 B.n194 VSUBS 0.008828f
C984 B.n195 VSUBS 0.008828f
C985 B.n196 VSUBS 0.008828f
C986 B.n197 VSUBS 0.008828f
C987 B.n198 VSUBS 0.008828f
C988 B.n199 VSUBS 0.008828f
C989 B.n200 VSUBS 0.008828f
C990 B.n201 VSUBS 0.008828f
C991 B.n202 VSUBS 0.008828f
C992 B.n203 VSUBS 0.008828f
C993 B.n204 VSUBS 0.008828f
C994 B.n205 VSUBS 0.008828f
C995 B.n206 VSUBS 0.008828f
C996 B.n207 VSUBS 0.008828f
C997 B.n208 VSUBS 0.008828f
C998 B.n209 VSUBS 0.008828f
C999 B.n210 VSUBS 0.008828f
C1000 B.n211 VSUBS 0.008828f
C1001 B.n212 VSUBS 0.008828f
C1002 B.n213 VSUBS 0.008828f
C1003 B.n214 VSUBS 0.008828f
C1004 B.n215 VSUBS 0.008828f
C1005 B.n216 VSUBS 0.008828f
C1006 B.n217 VSUBS 0.008828f
C1007 B.n218 VSUBS 0.008828f
C1008 B.n219 VSUBS 0.008828f
C1009 B.n220 VSUBS 0.008828f
C1010 B.n221 VSUBS 0.008828f
C1011 B.n222 VSUBS 0.008828f
C1012 B.n223 VSUBS 0.008828f
C1013 B.n224 VSUBS 0.008828f
C1014 B.n225 VSUBS 0.008828f
C1015 B.n226 VSUBS 0.008828f
C1016 B.n227 VSUBS 0.008828f
C1017 B.n228 VSUBS 0.008828f
C1018 B.n229 VSUBS 0.008828f
C1019 B.n230 VSUBS 0.008828f
C1020 B.n231 VSUBS 0.008828f
C1021 B.n232 VSUBS 0.008828f
C1022 B.n233 VSUBS 0.008828f
C1023 B.n234 VSUBS 0.008828f
C1024 B.n235 VSUBS 0.008828f
C1025 B.n236 VSUBS 0.008828f
C1026 B.n237 VSUBS 0.008828f
C1027 B.n238 VSUBS 0.008828f
C1028 B.n239 VSUBS 0.008828f
C1029 B.n240 VSUBS 0.008828f
C1030 B.n241 VSUBS 0.008828f
C1031 B.n242 VSUBS 0.008828f
C1032 B.n243 VSUBS 0.008828f
C1033 B.n244 VSUBS 0.008828f
C1034 B.n245 VSUBS 0.008828f
C1035 B.n246 VSUBS 0.008828f
C1036 B.n247 VSUBS 0.008828f
C1037 B.n248 VSUBS 0.008828f
C1038 B.n249 VSUBS 0.008828f
C1039 B.n250 VSUBS 0.008828f
C1040 B.n251 VSUBS 0.008828f
C1041 B.n252 VSUBS 0.008828f
C1042 B.n253 VSUBS 0.008828f
C1043 B.n254 VSUBS 0.008828f
C1044 B.n255 VSUBS 0.021713f
C1045 B.n256 VSUBS 0.022428f
C1046 B.n257 VSUBS 0.022428f
C1047 B.n258 VSUBS 0.008828f
C1048 B.n259 VSUBS 0.008828f
C1049 B.n260 VSUBS 0.008828f
C1050 B.n261 VSUBS 0.008828f
C1051 B.n262 VSUBS 0.008828f
C1052 B.n263 VSUBS 0.008828f
C1053 B.n264 VSUBS 0.008828f
C1054 B.n265 VSUBS 0.008828f
C1055 B.n266 VSUBS 0.008828f
C1056 B.n267 VSUBS 0.008828f
C1057 B.n268 VSUBS 0.008828f
C1058 B.n269 VSUBS 0.008828f
C1059 B.n270 VSUBS 0.008828f
C1060 B.n271 VSUBS 0.008828f
C1061 B.n272 VSUBS 0.008828f
C1062 B.n273 VSUBS 0.008828f
C1063 B.n274 VSUBS 0.008828f
C1064 B.n275 VSUBS 0.008828f
C1065 B.n276 VSUBS 0.008828f
C1066 B.n277 VSUBS 0.008828f
C1067 B.n278 VSUBS 0.008828f
C1068 B.n279 VSUBS 0.008828f
C1069 B.n280 VSUBS 0.008828f
C1070 B.n281 VSUBS 0.008828f
C1071 B.n282 VSUBS 0.008828f
C1072 B.n283 VSUBS 0.008828f
C1073 B.n284 VSUBS 0.008828f
C1074 B.n285 VSUBS 0.008828f
C1075 B.n286 VSUBS 0.008828f
C1076 B.n287 VSUBS 0.008828f
C1077 B.n288 VSUBS 0.008828f
C1078 B.n289 VSUBS 0.008828f
C1079 B.n290 VSUBS 0.008828f
C1080 B.n291 VSUBS 0.008828f
C1081 B.n292 VSUBS 0.008828f
C1082 B.n293 VSUBS 0.008828f
C1083 B.n294 VSUBS 0.008828f
C1084 B.n295 VSUBS 0.008828f
C1085 B.n296 VSUBS 0.008828f
C1086 B.n297 VSUBS 0.008828f
C1087 B.n298 VSUBS 0.008828f
C1088 B.n299 VSUBS 0.008828f
C1089 B.n300 VSUBS 0.008828f
C1090 B.n301 VSUBS 0.008828f
C1091 B.n302 VSUBS 0.008828f
C1092 B.n303 VSUBS 0.008828f
C1093 B.n304 VSUBS 0.008828f
C1094 B.n305 VSUBS 0.008828f
C1095 B.n306 VSUBS 0.008828f
C1096 B.n307 VSUBS 0.008828f
C1097 B.n308 VSUBS 0.008828f
C1098 B.n309 VSUBS 0.008828f
C1099 B.n310 VSUBS 0.008828f
C1100 B.n311 VSUBS 0.008828f
C1101 B.n312 VSUBS 0.008828f
C1102 B.n313 VSUBS 0.008828f
C1103 B.n314 VSUBS 0.008828f
C1104 B.n315 VSUBS 0.008828f
C1105 B.n316 VSUBS 0.008828f
C1106 B.n317 VSUBS 0.008828f
C1107 B.n318 VSUBS 0.006102f
C1108 B.n319 VSUBS 0.020454f
C1109 B.n320 VSUBS 0.00714f
C1110 B.n321 VSUBS 0.008828f
C1111 B.n322 VSUBS 0.008828f
C1112 B.n323 VSUBS 0.008828f
C1113 B.n324 VSUBS 0.008828f
C1114 B.n325 VSUBS 0.008828f
C1115 B.n326 VSUBS 0.008828f
C1116 B.n327 VSUBS 0.008828f
C1117 B.n328 VSUBS 0.008828f
C1118 B.n329 VSUBS 0.008828f
C1119 B.n330 VSUBS 0.008828f
C1120 B.n331 VSUBS 0.008828f
C1121 B.n332 VSUBS 0.00714f
C1122 B.n333 VSUBS 0.008828f
C1123 B.n334 VSUBS 0.008828f
C1124 B.n335 VSUBS 0.006102f
C1125 B.n336 VSUBS 0.008828f
C1126 B.n337 VSUBS 0.008828f
C1127 B.n338 VSUBS 0.008828f
C1128 B.n339 VSUBS 0.008828f
C1129 B.n340 VSUBS 0.008828f
C1130 B.n341 VSUBS 0.008828f
C1131 B.n342 VSUBS 0.008828f
C1132 B.n343 VSUBS 0.008828f
C1133 B.n344 VSUBS 0.008828f
C1134 B.n345 VSUBS 0.008828f
C1135 B.n346 VSUBS 0.008828f
C1136 B.n347 VSUBS 0.008828f
C1137 B.n348 VSUBS 0.008828f
C1138 B.n349 VSUBS 0.008828f
C1139 B.n350 VSUBS 0.008828f
C1140 B.n351 VSUBS 0.008828f
C1141 B.n352 VSUBS 0.008828f
C1142 B.n353 VSUBS 0.008828f
C1143 B.n354 VSUBS 0.008828f
C1144 B.n355 VSUBS 0.008828f
C1145 B.n356 VSUBS 0.008828f
C1146 B.n357 VSUBS 0.008828f
C1147 B.n358 VSUBS 0.008828f
C1148 B.n359 VSUBS 0.008828f
C1149 B.n360 VSUBS 0.008828f
C1150 B.n361 VSUBS 0.008828f
C1151 B.n362 VSUBS 0.008828f
C1152 B.n363 VSUBS 0.008828f
C1153 B.n364 VSUBS 0.008828f
C1154 B.n365 VSUBS 0.008828f
C1155 B.n366 VSUBS 0.008828f
C1156 B.n367 VSUBS 0.008828f
C1157 B.n368 VSUBS 0.008828f
C1158 B.n369 VSUBS 0.008828f
C1159 B.n370 VSUBS 0.008828f
C1160 B.n371 VSUBS 0.008828f
C1161 B.n372 VSUBS 0.008828f
C1162 B.n373 VSUBS 0.008828f
C1163 B.n374 VSUBS 0.008828f
C1164 B.n375 VSUBS 0.008828f
C1165 B.n376 VSUBS 0.008828f
C1166 B.n377 VSUBS 0.008828f
C1167 B.n378 VSUBS 0.008828f
C1168 B.n379 VSUBS 0.008828f
C1169 B.n380 VSUBS 0.008828f
C1170 B.n381 VSUBS 0.008828f
C1171 B.n382 VSUBS 0.008828f
C1172 B.n383 VSUBS 0.008828f
C1173 B.n384 VSUBS 0.008828f
C1174 B.n385 VSUBS 0.008828f
C1175 B.n386 VSUBS 0.008828f
C1176 B.n387 VSUBS 0.008828f
C1177 B.n388 VSUBS 0.008828f
C1178 B.n389 VSUBS 0.008828f
C1179 B.n390 VSUBS 0.008828f
C1180 B.n391 VSUBS 0.008828f
C1181 B.n392 VSUBS 0.008828f
C1182 B.n393 VSUBS 0.008828f
C1183 B.n394 VSUBS 0.008828f
C1184 B.n395 VSUBS 0.008828f
C1185 B.n396 VSUBS 0.022428f
C1186 B.n397 VSUBS 0.021713f
C1187 B.n398 VSUBS 0.021713f
C1188 B.n399 VSUBS 0.008828f
C1189 B.n400 VSUBS 0.008828f
C1190 B.n401 VSUBS 0.008828f
C1191 B.n402 VSUBS 0.008828f
C1192 B.n403 VSUBS 0.008828f
C1193 B.n404 VSUBS 0.008828f
C1194 B.n405 VSUBS 0.008828f
C1195 B.n406 VSUBS 0.008828f
C1196 B.n407 VSUBS 0.008828f
C1197 B.n408 VSUBS 0.008828f
C1198 B.n409 VSUBS 0.008828f
C1199 B.n410 VSUBS 0.008828f
C1200 B.n411 VSUBS 0.008828f
C1201 B.n412 VSUBS 0.008828f
C1202 B.n413 VSUBS 0.008828f
C1203 B.n414 VSUBS 0.008828f
C1204 B.n415 VSUBS 0.008828f
C1205 B.n416 VSUBS 0.008828f
C1206 B.n417 VSUBS 0.008828f
C1207 B.n418 VSUBS 0.008828f
C1208 B.n419 VSUBS 0.008828f
C1209 B.n420 VSUBS 0.008828f
C1210 B.n421 VSUBS 0.008828f
C1211 B.n422 VSUBS 0.008828f
C1212 B.n423 VSUBS 0.008828f
C1213 B.n424 VSUBS 0.008828f
C1214 B.n425 VSUBS 0.008828f
C1215 B.n426 VSUBS 0.008828f
C1216 B.n427 VSUBS 0.008828f
C1217 B.n428 VSUBS 0.008828f
C1218 B.n429 VSUBS 0.008828f
C1219 B.n430 VSUBS 0.008828f
C1220 B.n431 VSUBS 0.008828f
C1221 B.n432 VSUBS 0.008828f
C1222 B.n433 VSUBS 0.008828f
C1223 B.n434 VSUBS 0.008828f
C1224 B.n435 VSUBS 0.008828f
C1225 B.n436 VSUBS 0.008828f
C1226 B.n437 VSUBS 0.008828f
C1227 B.n438 VSUBS 0.008828f
C1228 B.n439 VSUBS 0.008828f
C1229 B.n440 VSUBS 0.008828f
C1230 B.n441 VSUBS 0.008828f
C1231 B.n442 VSUBS 0.008828f
C1232 B.n443 VSUBS 0.008828f
C1233 B.n444 VSUBS 0.008828f
C1234 B.n445 VSUBS 0.008828f
C1235 B.n446 VSUBS 0.008828f
C1236 B.n447 VSUBS 0.008828f
C1237 B.n448 VSUBS 0.008828f
C1238 B.n449 VSUBS 0.008828f
C1239 B.n450 VSUBS 0.008828f
C1240 B.n451 VSUBS 0.008828f
C1241 B.n452 VSUBS 0.008828f
C1242 B.n453 VSUBS 0.008828f
C1243 B.n454 VSUBS 0.008828f
C1244 B.n455 VSUBS 0.008828f
C1245 B.n456 VSUBS 0.008828f
C1246 B.n457 VSUBS 0.008828f
C1247 B.n458 VSUBS 0.008828f
C1248 B.n459 VSUBS 0.008828f
C1249 B.n460 VSUBS 0.008828f
C1250 B.n461 VSUBS 0.008828f
C1251 B.n462 VSUBS 0.008828f
C1252 B.n463 VSUBS 0.008828f
C1253 B.n464 VSUBS 0.008828f
C1254 B.n465 VSUBS 0.008828f
C1255 B.n466 VSUBS 0.008828f
C1256 B.n467 VSUBS 0.008828f
C1257 B.n468 VSUBS 0.008828f
C1258 B.n469 VSUBS 0.008828f
C1259 B.n470 VSUBS 0.008828f
C1260 B.n471 VSUBS 0.008828f
C1261 B.n472 VSUBS 0.008828f
C1262 B.n473 VSUBS 0.008828f
C1263 B.n474 VSUBS 0.008828f
C1264 B.n475 VSUBS 0.008828f
C1265 B.n476 VSUBS 0.008828f
C1266 B.n477 VSUBS 0.008828f
C1267 B.n478 VSUBS 0.008828f
C1268 B.n479 VSUBS 0.008828f
C1269 B.n480 VSUBS 0.008828f
C1270 B.n481 VSUBS 0.008828f
C1271 B.n482 VSUBS 0.008828f
C1272 B.n483 VSUBS 0.008828f
C1273 B.n484 VSUBS 0.008828f
C1274 B.n485 VSUBS 0.008828f
C1275 B.n486 VSUBS 0.008828f
C1276 B.n487 VSUBS 0.008828f
C1277 B.n488 VSUBS 0.008828f
C1278 B.n489 VSUBS 0.008828f
C1279 B.n490 VSUBS 0.008828f
C1280 B.n491 VSUBS 0.008828f
C1281 B.n492 VSUBS 0.008828f
C1282 B.n493 VSUBS 0.008828f
C1283 B.n494 VSUBS 0.008828f
C1284 B.n495 VSUBS 0.008828f
C1285 B.n496 VSUBS 0.008828f
C1286 B.n497 VSUBS 0.008828f
C1287 B.n498 VSUBS 0.008828f
C1288 B.n499 VSUBS 0.008828f
C1289 B.n500 VSUBS 0.008828f
C1290 B.n501 VSUBS 0.008828f
C1291 B.n502 VSUBS 0.008828f
C1292 B.n503 VSUBS 0.008828f
C1293 B.n504 VSUBS 0.008828f
C1294 B.n505 VSUBS 0.008828f
C1295 B.n506 VSUBS 0.008828f
C1296 B.n507 VSUBS 0.008828f
C1297 B.n508 VSUBS 0.008828f
C1298 B.n509 VSUBS 0.008828f
C1299 B.n510 VSUBS 0.008828f
C1300 B.n511 VSUBS 0.008828f
C1301 B.n512 VSUBS 0.008828f
C1302 B.n513 VSUBS 0.008828f
C1303 B.n514 VSUBS 0.008828f
C1304 B.n515 VSUBS 0.008828f
C1305 B.n516 VSUBS 0.008828f
C1306 B.n517 VSUBS 0.008828f
C1307 B.n518 VSUBS 0.008828f
C1308 B.n519 VSUBS 0.008828f
C1309 B.n520 VSUBS 0.008828f
C1310 B.n521 VSUBS 0.008828f
C1311 B.n522 VSUBS 0.008828f
C1312 B.n523 VSUBS 0.008828f
C1313 B.n524 VSUBS 0.008828f
C1314 B.n525 VSUBS 0.008828f
C1315 B.n526 VSUBS 0.008828f
C1316 B.n527 VSUBS 0.008828f
C1317 B.n528 VSUBS 0.008828f
C1318 B.n529 VSUBS 0.022658f
C1319 B.n530 VSUBS 0.021713f
C1320 B.n531 VSUBS 0.022428f
C1321 B.n532 VSUBS 0.008828f
C1322 B.n533 VSUBS 0.008828f
C1323 B.n534 VSUBS 0.008828f
C1324 B.n535 VSUBS 0.008828f
C1325 B.n536 VSUBS 0.008828f
C1326 B.n537 VSUBS 0.008828f
C1327 B.n538 VSUBS 0.008828f
C1328 B.n539 VSUBS 0.008828f
C1329 B.n540 VSUBS 0.008828f
C1330 B.n541 VSUBS 0.008828f
C1331 B.n542 VSUBS 0.008828f
C1332 B.n543 VSUBS 0.008828f
C1333 B.n544 VSUBS 0.008828f
C1334 B.n545 VSUBS 0.008828f
C1335 B.n546 VSUBS 0.008828f
C1336 B.n547 VSUBS 0.008828f
C1337 B.n548 VSUBS 0.008828f
C1338 B.n549 VSUBS 0.008828f
C1339 B.n550 VSUBS 0.008828f
C1340 B.n551 VSUBS 0.008828f
C1341 B.n552 VSUBS 0.008828f
C1342 B.n553 VSUBS 0.008828f
C1343 B.n554 VSUBS 0.008828f
C1344 B.n555 VSUBS 0.008828f
C1345 B.n556 VSUBS 0.008828f
C1346 B.n557 VSUBS 0.008828f
C1347 B.n558 VSUBS 0.008828f
C1348 B.n559 VSUBS 0.008828f
C1349 B.n560 VSUBS 0.008828f
C1350 B.n561 VSUBS 0.008828f
C1351 B.n562 VSUBS 0.008828f
C1352 B.n563 VSUBS 0.008828f
C1353 B.n564 VSUBS 0.008828f
C1354 B.n565 VSUBS 0.008828f
C1355 B.n566 VSUBS 0.008828f
C1356 B.n567 VSUBS 0.008828f
C1357 B.n568 VSUBS 0.008828f
C1358 B.n569 VSUBS 0.008828f
C1359 B.n570 VSUBS 0.008828f
C1360 B.n571 VSUBS 0.008828f
C1361 B.n572 VSUBS 0.008828f
C1362 B.n573 VSUBS 0.008828f
C1363 B.n574 VSUBS 0.008828f
C1364 B.n575 VSUBS 0.008828f
C1365 B.n576 VSUBS 0.008828f
C1366 B.n577 VSUBS 0.008828f
C1367 B.n578 VSUBS 0.008828f
C1368 B.n579 VSUBS 0.008828f
C1369 B.n580 VSUBS 0.008828f
C1370 B.n581 VSUBS 0.008828f
C1371 B.n582 VSUBS 0.008828f
C1372 B.n583 VSUBS 0.008828f
C1373 B.n584 VSUBS 0.008828f
C1374 B.n585 VSUBS 0.008828f
C1375 B.n586 VSUBS 0.008828f
C1376 B.n587 VSUBS 0.008828f
C1377 B.n588 VSUBS 0.008828f
C1378 B.n589 VSUBS 0.008828f
C1379 B.n590 VSUBS 0.008828f
C1380 B.n591 VSUBS 0.008828f
C1381 B.n592 VSUBS 0.008828f
C1382 B.n593 VSUBS 0.006102f
C1383 B.n594 VSUBS 0.020454f
C1384 B.n595 VSUBS 0.00714f
C1385 B.n596 VSUBS 0.008828f
C1386 B.n597 VSUBS 0.008828f
C1387 B.n598 VSUBS 0.008828f
C1388 B.n599 VSUBS 0.008828f
C1389 B.n600 VSUBS 0.008828f
C1390 B.n601 VSUBS 0.008828f
C1391 B.n602 VSUBS 0.008828f
C1392 B.n603 VSUBS 0.008828f
C1393 B.n604 VSUBS 0.008828f
C1394 B.n605 VSUBS 0.008828f
C1395 B.n606 VSUBS 0.008828f
C1396 B.n607 VSUBS 0.00714f
C1397 B.n608 VSUBS 0.020454f
C1398 B.n609 VSUBS 0.006102f
C1399 B.n610 VSUBS 0.008828f
C1400 B.n611 VSUBS 0.008828f
C1401 B.n612 VSUBS 0.008828f
C1402 B.n613 VSUBS 0.008828f
C1403 B.n614 VSUBS 0.008828f
C1404 B.n615 VSUBS 0.008828f
C1405 B.n616 VSUBS 0.008828f
C1406 B.n617 VSUBS 0.008828f
C1407 B.n618 VSUBS 0.008828f
C1408 B.n619 VSUBS 0.008828f
C1409 B.n620 VSUBS 0.008828f
C1410 B.n621 VSUBS 0.008828f
C1411 B.n622 VSUBS 0.008828f
C1412 B.n623 VSUBS 0.008828f
C1413 B.n624 VSUBS 0.008828f
C1414 B.n625 VSUBS 0.008828f
C1415 B.n626 VSUBS 0.008828f
C1416 B.n627 VSUBS 0.008828f
C1417 B.n628 VSUBS 0.008828f
C1418 B.n629 VSUBS 0.008828f
C1419 B.n630 VSUBS 0.008828f
C1420 B.n631 VSUBS 0.008828f
C1421 B.n632 VSUBS 0.008828f
C1422 B.n633 VSUBS 0.008828f
C1423 B.n634 VSUBS 0.008828f
C1424 B.n635 VSUBS 0.008828f
C1425 B.n636 VSUBS 0.008828f
C1426 B.n637 VSUBS 0.008828f
C1427 B.n638 VSUBS 0.008828f
C1428 B.n639 VSUBS 0.008828f
C1429 B.n640 VSUBS 0.008828f
C1430 B.n641 VSUBS 0.008828f
C1431 B.n642 VSUBS 0.008828f
C1432 B.n643 VSUBS 0.008828f
C1433 B.n644 VSUBS 0.008828f
C1434 B.n645 VSUBS 0.008828f
C1435 B.n646 VSUBS 0.008828f
C1436 B.n647 VSUBS 0.008828f
C1437 B.n648 VSUBS 0.008828f
C1438 B.n649 VSUBS 0.008828f
C1439 B.n650 VSUBS 0.008828f
C1440 B.n651 VSUBS 0.008828f
C1441 B.n652 VSUBS 0.008828f
C1442 B.n653 VSUBS 0.008828f
C1443 B.n654 VSUBS 0.008828f
C1444 B.n655 VSUBS 0.008828f
C1445 B.n656 VSUBS 0.008828f
C1446 B.n657 VSUBS 0.008828f
C1447 B.n658 VSUBS 0.008828f
C1448 B.n659 VSUBS 0.008828f
C1449 B.n660 VSUBS 0.008828f
C1450 B.n661 VSUBS 0.008828f
C1451 B.n662 VSUBS 0.008828f
C1452 B.n663 VSUBS 0.008828f
C1453 B.n664 VSUBS 0.008828f
C1454 B.n665 VSUBS 0.008828f
C1455 B.n666 VSUBS 0.008828f
C1456 B.n667 VSUBS 0.008828f
C1457 B.n668 VSUBS 0.008828f
C1458 B.n669 VSUBS 0.008828f
C1459 B.n670 VSUBS 0.008828f
C1460 B.n671 VSUBS 0.022428f
C1461 B.n672 VSUBS 0.021713f
C1462 B.n673 VSUBS 0.021713f
C1463 B.n674 VSUBS 0.008828f
C1464 B.n675 VSUBS 0.008828f
C1465 B.n676 VSUBS 0.008828f
C1466 B.n677 VSUBS 0.008828f
C1467 B.n678 VSUBS 0.008828f
C1468 B.n679 VSUBS 0.008828f
C1469 B.n680 VSUBS 0.008828f
C1470 B.n681 VSUBS 0.008828f
C1471 B.n682 VSUBS 0.008828f
C1472 B.n683 VSUBS 0.008828f
C1473 B.n684 VSUBS 0.008828f
C1474 B.n685 VSUBS 0.008828f
C1475 B.n686 VSUBS 0.008828f
C1476 B.n687 VSUBS 0.008828f
C1477 B.n688 VSUBS 0.008828f
C1478 B.n689 VSUBS 0.008828f
C1479 B.n690 VSUBS 0.008828f
C1480 B.n691 VSUBS 0.008828f
C1481 B.n692 VSUBS 0.008828f
C1482 B.n693 VSUBS 0.008828f
C1483 B.n694 VSUBS 0.008828f
C1484 B.n695 VSUBS 0.008828f
C1485 B.n696 VSUBS 0.008828f
C1486 B.n697 VSUBS 0.008828f
C1487 B.n698 VSUBS 0.008828f
C1488 B.n699 VSUBS 0.008828f
C1489 B.n700 VSUBS 0.008828f
C1490 B.n701 VSUBS 0.008828f
C1491 B.n702 VSUBS 0.008828f
C1492 B.n703 VSUBS 0.008828f
C1493 B.n704 VSUBS 0.008828f
C1494 B.n705 VSUBS 0.008828f
C1495 B.n706 VSUBS 0.008828f
C1496 B.n707 VSUBS 0.008828f
C1497 B.n708 VSUBS 0.008828f
C1498 B.n709 VSUBS 0.008828f
C1499 B.n710 VSUBS 0.008828f
C1500 B.n711 VSUBS 0.008828f
C1501 B.n712 VSUBS 0.008828f
C1502 B.n713 VSUBS 0.008828f
C1503 B.n714 VSUBS 0.008828f
C1504 B.n715 VSUBS 0.008828f
C1505 B.n716 VSUBS 0.008828f
C1506 B.n717 VSUBS 0.008828f
C1507 B.n718 VSUBS 0.008828f
C1508 B.n719 VSUBS 0.008828f
C1509 B.n720 VSUBS 0.008828f
C1510 B.n721 VSUBS 0.008828f
C1511 B.n722 VSUBS 0.008828f
C1512 B.n723 VSUBS 0.008828f
C1513 B.n724 VSUBS 0.008828f
C1514 B.n725 VSUBS 0.008828f
C1515 B.n726 VSUBS 0.008828f
C1516 B.n727 VSUBS 0.008828f
C1517 B.n728 VSUBS 0.008828f
C1518 B.n729 VSUBS 0.008828f
C1519 B.n730 VSUBS 0.008828f
C1520 B.n731 VSUBS 0.008828f
C1521 B.n732 VSUBS 0.008828f
C1522 B.n733 VSUBS 0.008828f
C1523 B.n734 VSUBS 0.008828f
C1524 B.n735 VSUBS 0.008828f
C1525 B.n736 VSUBS 0.008828f
C1526 B.n737 VSUBS 0.008828f
C1527 B.n738 VSUBS 0.008828f
C1528 B.n739 VSUBS 0.01999f
.ends

