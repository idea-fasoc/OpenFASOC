* NGSPICE file created from diff_pair_sample_1427.ext - technology: sky130A

.subckt diff_pair_sample_1427 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=3.3696 ps=18.06 w=8.64 l=3.78
X1 VTAIL.t0 VN.t0 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=1.4256 ps=8.97 w=8.64 l=3.78
X2 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.78
X3 VDD2.t4 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=3.3696 ps=18.06 w=8.64 l=3.78
X4 VDD1.t4 VP.t1 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=3.3696 ps=18.06 w=8.64 l=3.78
X5 VDD1.t3 VP.t2 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=1.4256 ps=8.97 w=8.64 l=3.78
X6 VTAIL.t5 VN.t2 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=1.4256 ps=8.97 w=8.64 l=3.78
X7 VTAIL.t9 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=1.4256 ps=8.97 w=8.64 l=3.78
X8 VDD1.t1 VP.t4 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=1.4256 ps=8.97 w=8.64 l=3.78
X9 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=1.4256 ps=8.97 w=8.64 l=3.78
X10 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.78
X11 VDD2.t1 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=3.3696 ps=18.06 w=8.64 l=3.78
X12 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.78
X13 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=0 ps=0 w=8.64 l=3.78
X14 VDD2.t0 VN.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.3696 pd=18.06 as=1.4256 ps=8.97 w=8.64 l=3.78
X15 VTAIL.t6 VP.t5 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.4256 pd=8.97 as=1.4256 ps=8.97 w=8.64 l=3.78
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n56 VP.n55 161.3
R9 VP.n54 VP.n1 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n2 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n3 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n45 VP.n4 161.3
R16 VP.n44 VP.n43 161.3
R17 VP.n42 VP.n5 161.3
R18 VP.n41 VP.n40 161.3
R19 VP.n39 VP.n6 161.3
R20 VP.n38 VP.n37 161.3
R21 VP.n36 VP.n7 161.3
R22 VP.n35 VP.n34 161.3
R23 VP.n33 VP.n8 161.3
R24 VP.n32 VP.n31 161.3
R25 VP.n15 VP.t2 88.5049
R26 VP.n30 VP.n29 84.5354
R27 VP.n57 VP.n0 84.5354
R28 VP.n28 VP.n9 84.5354
R29 VP.n43 VP.t3 55.0862
R30 VP.n30 VP.t4 55.0862
R31 VP.n0 VP.t1 55.0862
R32 VP.n14 VP.t5 55.0862
R33 VP.n9 VP.t0 55.0862
R34 VP.n29 VP.n28 50.8438
R35 VP.n15 VP.n14 50.3788
R36 VP.n37 VP.n36 45.7662
R37 VP.n49 VP.n2 45.7662
R38 VP.n20 VP.n11 45.7662
R39 VP.n37 VP.n6 35.055
R40 VP.n49 VP.n48 35.055
R41 VP.n20 VP.n19 35.055
R42 VP.n31 VP.n8 24.3439
R43 VP.n35 VP.n8 24.3439
R44 VP.n36 VP.n35 24.3439
R45 VP.n41 VP.n6 24.3439
R46 VP.n42 VP.n41 24.3439
R47 VP.n43 VP.n42 24.3439
R48 VP.n43 VP.n4 24.3439
R49 VP.n47 VP.n4 24.3439
R50 VP.n48 VP.n47 24.3439
R51 VP.n53 VP.n2 24.3439
R52 VP.n54 VP.n53 24.3439
R53 VP.n55 VP.n54 24.3439
R54 VP.n24 VP.n11 24.3439
R55 VP.n25 VP.n24 24.3439
R56 VP.n26 VP.n25 24.3439
R57 VP.n14 VP.n13 24.3439
R58 VP.n18 VP.n13 24.3439
R59 VP.n19 VP.n18 24.3439
R60 VP.n31 VP.n30 5.35606
R61 VP.n55 VP.n0 5.35606
R62 VP.n26 VP.n9 5.35606
R63 VP.n16 VP.n15 2.42076
R64 VP.n28 VP.n27 0.355081
R65 VP.n32 VP.n29 0.355081
R66 VP.n57 VP.n56 0.355081
R67 VP VP.n57 0.26685
R68 VP.n17 VP.n16 0.189894
R69 VP.n17 VP.n12 0.189894
R70 VP.n21 VP.n12 0.189894
R71 VP.n22 VP.n21 0.189894
R72 VP.n23 VP.n22 0.189894
R73 VP.n23 VP.n10 0.189894
R74 VP.n27 VP.n10 0.189894
R75 VP.n33 VP.n32 0.189894
R76 VP.n34 VP.n33 0.189894
R77 VP.n34 VP.n7 0.189894
R78 VP.n38 VP.n7 0.189894
R79 VP.n39 VP.n38 0.189894
R80 VP.n40 VP.n39 0.189894
R81 VP.n40 VP.n5 0.189894
R82 VP.n44 VP.n5 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n46 VP.n45 0.189894
R85 VP.n46 VP.n3 0.189894
R86 VP.n50 VP.n3 0.189894
R87 VP.n51 VP.n50 0.189894
R88 VP.n52 VP.n51 0.189894
R89 VP.n52 VP.n1 0.189894
R90 VP.n56 VP.n1 0.189894
R91 VTAIL.n186 VTAIL.n146 289.615
R92 VTAIL.n42 VTAIL.n2 289.615
R93 VTAIL.n140 VTAIL.n100 289.615
R94 VTAIL.n92 VTAIL.n52 289.615
R95 VTAIL.n161 VTAIL.n160 185
R96 VTAIL.n158 VTAIL.n157 185
R97 VTAIL.n167 VTAIL.n166 185
R98 VTAIL.n169 VTAIL.n168 185
R99 VTAIL.n154 VTAIL.n153 185
R100 VTAIL.n175 VTAIL.n174 185
R101 VTAIL.n178 VTAIL.n177 185
R102 VTAIL.n176 VTAIL.n150 185
R103 VTAIL.n183 VTAIL.n149 185
R104 VTAIL.n185 VTAIL.n184 185
R105 VTAIL.n187 VTAIL.n186 185
R106 VTAIL.n17 VTAIL.n16 185
R107 VTAIL.n14 VTAIL.n13 185
R108 VTAIL.n23 VTAIL.n22 185
R109 VTAIL.n25 VTAIL.n24 185
R110 VTAIL.n10 VTAIL.n9 185
R111 VTAIL.n31 VTAIL.n30 185
R112 VTAIL.n34 VTAIL.n33 185
R113 VTAIL.n32 VTAIL.n6 185
R114 VTAIL.n39 VTAIL.n5 185
R115 VTAIL.n41 VTAIL.n40 185
R116 VTAIL.n43 VTAIL.n42 185
R117 VTAIL.n141 VTAIL.n140 185
R118 VTAIL.n139 VTAIL.n138 185
R119 VTAIL.n137 VTAIL.n103 185
R120 VTAIL.n107 VTAIL.n104 185
R121 VTAIL.n132 VTAIL.n131 185
R122 VTAIL.n130 VTAIL.n129 185
R123 VTAIL.n109 VTAIL.n108 185
R124 VTAIL.n124 VTAIL.n123 185
R125 VTAIL.n122 VTAIL.n121 185
R126 VTAIL.n113 VTAIL.n112 185
R127 VTAIL.n116 VTAIL.n115 185
R128 VTAIL.n93 VTAIL.n92 185
R129 VTAIL.n91 VTAIL.n90 185
R130 VTAIL.n89 VTAIL.n55 185
R131 VTAIL.n59 VTAIL.n56 185
R132 VTAIL.n84 VTAIL.n83 185
R133 VTAIL.n82 VTAIL.n81 185
R134 VTAIL.n61 VTAIL.n60 185
R135 VTAIL.n76 VTAIL.n75 185
R136 VTAIL.n74 VTAIL.n73 185
R137 VTAIL.n65 VTAIL.n64 185
R138 VTAIL.n68 VTAIL.n67 185
R139 VTAIL.t2 VTAIL.n159 149.524
R140 VTAIL.t10 VTAIL.n15 149.524
R141 VTAIL.t8 VTAIL.n114 149.524
R142 VTAIL.t3 VTAIL.n66 149.524
R143 VTAIL.n160 VTAIL.n157 104.615
R144 VTAIL.n167 VTAIL.n157 104.615
R145 VTAIL.n168 VTAIL.n167 104.615
R146 VTAIL.n168 VTAIL.n153 104.615
R147 VTAIL.n175 VTAIL.n153 104.615
R148 VTAIL.n177 VTAIL.n175 104.615
R149 VTAIL.n177 VTAIL.n176 104.615
R150 VTAIL.n176 VTAIL.n149 104.615
R151 VTAIL.n185 VTAIL.n149 104.615
R152 VTAIL.n186 VTAIL.n185 104.615
R153 VTAIL.n16 VTAIL.n13 104.615
R154 VTAIL.n23 VTAIL.n13 104.615
R155 VTAIL.n24 VTAIL.n23 104.615
R156 VTAIL.n24 VTAIL.n9 104.615
R157 VTAIL.n31 VTAIL.n9 104.615
R158 VTAIL.n33 VTAIL.n31 104.615
R159 VTAIL.n33 VTAIL.n32 104.615
R160 VTAIL.n32 VTAIL.n5 104.615
R161 VTAIL.n41 VTAIL.n5 104.615
R162 VTAIL.n42 VTAIL.n41 104.615
R163 VTAIL.n140 VTAIL.n139 104.615
R164 VTAIL.n139 VTAIL.n103 104.615
R165 VTAIL.n107 VTAIL.n103 104.615
R166 VTAIL.n131 VTAIL.n107 104.615
R167 VTAIL.n131 VTAIL.n130 104.615
R168 VTAIL.n130 VTAIL.n108 104.615
R169 VTAIL.n123 VTAIL.n108 104.615
R170 VTAIL.n123 VTAIL.n122 104.615
R171 VTAIL.n122 VTAIL.n112 104.615
R172 VTAIL.n115 VTAIL.n112 104.615
R173 VTAIL.n92 VTAIL.n91 104.615
R174 VTAIL.n91 VTAIL.n55 104.615
R175 VTAIL.n59 VTAIL.n55 104.615
R176 VTAIL.n83 VTAIL.n59 104.615
R177 VTAIL.n83 VTAIL.n82 104.615
R178 VTAIL.n82 VTAIL.n60 104.615
R179 VTAIL.n75 VTAIL.n60 104.615
R180 VTAIL.n75 VTAIL.n74 104.615
R181 VTAIL.n74 VTAIL.n64 104.615
R182 VTAIL.n67 VTAIL.n64 104.615
R183 VTAIL.n160 VTAIL.t2 52.3082
R184 VTAIL.n16 VTAIL.t10 52.3082
R185 VTAIL.n115 VTAIL.t8 52.3082
R186 VTAIL.n67 VTAIL.t3 52.3082
R187 VTAIL.n99 VTAIL.n98 49.0897
R188 VTAIL.n51 VTAIL.n50 49.0897
R189 VTAIL.n1 VTAIL.n0 49.0895
R190 VTAIL.n49 VTAIL.n48 49.0895
R191 VTAIL.n191 VTAIL.n190 34.5126
R192 VTAIL.n47 VTAIL.n46 34.5126
R193 VTAIL.n145 VTAIL.n144 34.5126
R194 VTAIL.n97 VTAIL.n96 34.5126
R195 VTAIL.n51 VTAIL.n49 26.9014
R196 VTAIL.n191 VTAIL.n145 23.3583
R197 VTAIL.n184 VTAIL.n183 13.1884
R198 VTAIL.n40 VTAIL.n39 13.1884
R199 VTAIL.n138 VTAIL.n137 13.1884
R200 VTAIL.n90 VTAIL.n89 13.1884
R201 VTAIL.n182 VTAIL.n150 12.8005
R202 VTAIL.n187 VTAIL.n148 12.8005
R203 VTAIL.n38 VTAIL.n6 12.8005
R204 VTAIL.n43 VTAIL.n4 12.8005
R205 VTAIL.n141 VTAIL.n102 12.8005
R206 VTAIL.n136 VTAIL.n104 12.8005
R207 VTAIL.n93 VTAIL.n54 12.8005
R208 VTAIL.n88 VTAIL.n56 12.8005
R209 VTAIL.n179 VTAIL.n178 12.0247
R210 VTAIL.n188 VTAIL.n146 12.0247
R211 VTAIL.n35 VTAIL.n34 12.0247
R212 VTAIL.n44 VTAIL.n2 12.0247
R213 VTAIL.n142 VTAIL.n100 12.0247
R214 VTAIL.n133 VTAIL.n132 12.0247
R215 VTAIL.n94 VTAIL.n52 12.0247
R216 VTAIL.n85 VTAIL.n84 12.0247
R217 VTAIL.n174 VTAIL.n152 11.249
R218 VTAIL.n30 VTAIL.n8 11.249
R219 VTAIL.n129 VTAIL.n106 11.249
R220 VTAIL.n81 VTAIL.n58 11.249
R221 VTAIL.n173 VTAIL.n154 10.4732
R222 VTAIL.n29 VTAIL.n10 10.4732
R223 VTAIL.n128 VTAIL.n109 10.4732
R224 VTAIL.n80 VTAIL.n61 10.4732
R225 VTAIL.n161 VTAIL.n159 10.2747
R226 VTAIL.n17 VTAIL.n15 10.2747
R227 VTAIL.n116 VTAIL.n114 10.2747
R228 VTAIL.n68 VTAIL.n66 10.2747
R229 VTAIL.n170 VTAIL.n169 9.69747
R230 VTAIL.n26 VTAIL.n25 9.69747
R231 VTAIL.n125 VTAIL.n124 9.69747
R232 VTAIL.n77 VTAIL.n76 9.69747
R233 VTAIL.n190 VTAIL.n189 9.45567
R234 VTAIL.n46 VTAIL.n45 9.45567
R235 VTAIL.n144 VTAIL.n143 9.45567
R236 VTAIL.n96 VTAIL.n95 9.45567
R237 VTAIL.n189 VTAIL.n188 9.3005
R238 VTAIL.n148 VTAIL.n147 9.3005
R239 VTAIL.n163 VTAIL.n162 9.3005
R240 VTAIL.n165 VTAIL.n164 9.3005
R241 VTAIL.n156 VTAIL.n155 9.3005
R242 VTAIL.n171 VTAIL.n170 9.3005
R243 VTAIL.n173 VTAIL.n172 9.3005
R244 VTAIL.n152 VTAIL.n151 9.3005
R245 VTAIL.n180 VTAIL.n179 9.3005
R246 VTAIL.n182 VTAIL.n181 9.3005
R247 VTAIL.n45 VTAIL.n44 9.3005
R248 VTAIL.n4 VTAIL.n3 9.3005
R249 VTAIL.n19 VTAIL.n18 9.3005
R250 VTAIL.n21 VTAIL.n20 9.3005
R251 VTAIL.n12 VTAIL.n11 9.3005
R252 VTAIL.n27 VTAIL.n26 9.3005
R253 VTAIL.n29 VTAIL.n28 9.3005
R254 VTAIL.n8 VTAIL.n7 9.3005
R255 VTAIL.n36 VTAIL.n35 9.3005
R256 VTAIL.n38 VTAIL.n37 9.3005
R257 VTAIL.n118 VTAIL.n117 9.3005
R258 VTAIL.n120 VTAIL.n119 9.3005
R259 VTAIL.n111 VTAIL.n110 9.3005
R260 VTAIL.n126 VTAIL.n125 9.3005
R261 VTAIL.n128 VTAIL.n127 9.3005
R262 VTAIL.n106 VTAIL.n105 9.3005
R263 VTAIL.n134 VTAIL.n133 9.3005
R264 VTAIL.n136 VTAIL.n135 9.3005
R265 VTAIL.n143 VTAIL.n142 9.3005
R266 VTAIL.n102 VTAIL.n101 9.3005
R267 VTAIL.n70 VTAIL.n69 9.3005
R268 VTAIL.n72 VTAIL.n71 9.3005
R269 VTAIL.n63 VTAIL.n62 9.3005
R270 VTAIL.n78 VTAIL.n77 9.3005
R271 VTAIL.n80 VTAIL.n79 9.3005
R272 VTAIL.n58 VTAIL.n57 9.3005
R273 VTAIL.n86 VTAIL.n85 9.3005
R274 VTAIL.n88 VTAIL.n87 9.3005
R275 VTAIL.n95 VTAIL.n94 9.3005
R276 VTAIL.n54 VTAIL.n53 9.3005
R277 VTAIL.n166 VTAIL.n156 8.92171
R278 VTAIL.n22 VTAIL.n12 8.92171
R279 VTAIL.n121 VTAIL.n111 8.92171
R280 VTAIL.n73 VTAIL.n63 8.92171
R281 VTAIL.n165 VTAIL.n158 8.14595
R282 VTAIL.n21 VTAIL.n14 8.14595
R283 VTAIL.n120 VTAIL.n113 8.14595
R284 VTAIL.n72 VTAIL.n65 8.14595
R285 VTAIL.n162 VTAIL.n161 7.3702
R286 VTAIL.n18 VTAIL.n17 7.3702
R287 VTAIL.n117 VTAIL.n116 7.3702
R288 VTAIL.n69 VTAIL.n68 7.3702
R289 VTAIL.n162 VTAIL.n158 5.81868
R290 VTAIL.n18 VTAIL.n14 5.81868
R291 VTAIL.n117 VTAIL.n113 5.81868
R292 VTAIL.n69 VTAIL.n65 5.81868
R293 VTAIL.n166 VTAIL.n165 5.04292
R294 VTAIL.n22 VTAIL.n21 5.04292
R295 VTAIL.n121 VTAIL.n120 5.04292
R296 VTAIL.n73 VTAIL.n72 5.04292
R297 VTAIL.n169 VTAIL.n156 4.26717
R298 VTAIL.n25 VTAIL.n12 4.26717
R299 VTAIL.n124 VTAIL.n111 4.26717
R300 VTAIL.n76 VTAIL.n63 4.26717
R301 VTAIL.n97 VTAIL.n51 3.5436
R302 VTAIL.n145 VTAIL.n99 3.5436
R303 VTAIL.n49 VTAIL.n47 3.5436
R304 VTAIL.n170 VTAIL.n154 3.49141
R305 VTAIL.n26 VTAIL.n10 3.49141
R306 VTAIL.n125 VTAIL.n109 3.49141
R307 VTAIL.n77 VTAIL.n61 3.49141
R308 VTAIL.n163 VTAIL.n159 2.84303
R309 VTAIL.n19 VTAIL.n15 2.84303
R310 VTAIL.n118 VTAIL.n114 2.84303
R311 VTAIL.n70 VTAIL.n66 2.84303
R312 VTAIL.n174 VTAIL.n173 2.71565
R313 VTAIL.n30 VTAIL.n29 2.71565
R314 VTAIL.n129 VTAIL.n128 2.71565
R315 VTAIL.n81 VTAIL.n80 2.71565
R316 VTAIL VTAIL.n191 2.59964
R317 VTAIL.n0 VTAIL.t1 2.29217
R318 VTAIL.n0 VTAIL.t5 2.29217
R319 VTAIL.n48 VTAIL.t7 2.29217
R320 VTAIL.n48 VTAIL.t9 2.29217
R321 VTAIL.n98 VTAIL.t11 2.29217
R322 VTAIL.n98 VTAIL.t6 2.29217
R323 VTAIL.n50 VTAIL.t4 2.29217
R324 VTAIL.n50 VTAIL.t0 2.29217
R325 VTAIL.n99 VTAIL.n97 2.24188
R326 VTAIL.n47 VTAIL.n1 2.24188
R327 VTAIL.n178 VTAIL.n152 1.93989
R328 VTAIL.n190 VTAIL.n146 1.93989
R329 VTAIL.n34 VTAIL.n8 1.93989
R330 VTAIL.n46 VTAIL.n2 1.93989
R331 VTAIL.n144 VTAIL.n100 1.93989
R332 VTAIL.n132 VTAIL.n106 1.93989
R333 VTAIL.n96 VTAIL.n52 1.93989
R334 VTAIL.n84 VTAIL.n58 1.93989
R335 VTAIL.n179 VTAIL.n150 1.16414
R336 VTAIL.n188 VTAIL.n187 1.16414
R337 VTAIL.n35 VTAIL.n6 1.16414
R338 VTAIL.n44 VTAIL.n43 1.16414
R339 VTAIL.n142 VTAIL.n141 1.16414
R340 VTAIL.n133 VTAIL.n104 1.16414
R341 VTAIL.n94 VTAIL.n93 1.16414
R342 VTAIL.n85 VTAIL.n56 1.16414
R343 VTAIL VTAIL.n1 0.944465
R344 VTAIL.n183 VTAIL.n182 0.388379
R345 VTAIL.n184 VTAIL.n148 0.388379
R346 VTAIL.n39 VTAIL.n38 0.388379
R347 VTAIL.n40 VTAIL.n4 0.388379
R348 VTAIL.n138 VTAIL.n102 0.388379
R349 VTAIL.n137 VTAIL.n136 0.388379
R350 VTAIL.n90 VTAIL.n54 0.388379
R351 VTAIL.n89 VTAIL.n88 0.388379
R352 VTAIL.n164 VTAIL.n163 0.155672
R353 VTAIL.n164 VTAIL.n155 0.155672
R354 VTAIL.n171 VTAIL.n155 0.155672
R355 VTAIL.n172 VTAIL.n171 0.155672
R356 VTAIL.n172 VTAIL.n151 0.155672
R357 VTAIL.n180 VTAIL.n151 0.155672
R358 VTAIL.n181 VTAIL.n180 0.155672
R359 VTAIL.n181 VTAIL.n147 0.155672
R360 VTAIL.n189 VTAIL.n147 0.155672
R361 VTAIL.n20 VTAIL.n19 0.155672
R362 VTAIL.n20 VTAIL.n11 0.155672
R363 VTAIL.n27 VTAIL.n11 0.155672
R364 VTAIL.n28 VTAIL.n27 0.155672
R365 VTAIL.n28 VTAIL.n7 0.155672
R366 VTAIL.n36 VTAIL.n7 0.155672
R367 VTAIL.n37 VTAIL.n36 0.155672
R368 VTAIL.n37 VTAIL.n3 0.155672
R369 VTAIL.n45 VTAIL.n3 0.155672
R370 VTAIL.n143 VTAIL.n101 0.155672
R371 VTAIL.n135 VTAIL.n101 0.155672
R372 VTAIL.n135 VTAIL.n134 0.155672
R373 VTAIL.n134 VTAIL.n105 0.155672
R374 VTAIL.n127 VTAIL.n105 0.155672
R375 VTAIL.n127 VTAIL.n126 0.155672
R376 VTAIL.n126 VTAIL.n110 0.155672
R377 VTAIL.n119 VTAIL.n110 0.155672
R378 VTAIL.n119 VTAIL.n118 0.155672
R379 VTAIL.n95 VTAIL.n53 0.155672
R380 VTAIL.n87 VTAIL.n53 0.155672
R381 VTAIL.n87 VTAIL.n86 0.155672
R382 VTAIL.n86 VTAIL.n57 0.155672
R383 VTAIL.n79 VTAIL.n57 0.155672
R384 VTAIL.n79 VTAIL.n78 0.155672
R385 VTAIL.n78 VTAIL.n62 0.155672
R386 VTAIL.n71 VTAIL.n62 0.155672
R387 VTAIL.n71 VTAIL.n70 0.155672
R388 VDD1.n40 VDD1.n0 289.615
R389 VDD1.n85 VDD1.n45 289.615
R390 VDD1.n41 VDD1.n40 185
R391 VDD1.n39 VDD1.n38 185
R392 VDD1.n37 VDD1.n3 185
R393 VDD1.n7 VDD1.n4 185
R394 VDD1.n32 VDD1.n31 185
R395 VDD1.n30 VDD1.n29 185
R396 VDD1.n9 VDD1.n8 185
R397 VDD1.n24 VDD1.n23 185
R398 VDD1.n22 VDD1.n21 185
R399 VDD1.n13 VDD1.n12 185
R400 VDD1.n16 VDD1.n15 185
R401 VDD1.n60 VDD1.n59 185
R402 VDD1.n57 VDD1.n56 185
R403 VDD1.n66 VDD1.n65 185
R404 VDD1.n68 VDD1.n67 185
R405 VDD1.n53 VDD1.n52 185
R406 VDD1.n74 VDD1.n73 185
R407 VDD1.n77 VDD1.n76 185
R408 VDD1.n75 VDD1.n49 185
R409 VDD1.n82 VDD1.n48 185
R410 VDD1.n84 VDD1.n83 185
R411 VDD1.n86 VDD1.n85 185
R412 VDD1.t3 VDD1.n14 149.524
R413 VDD1.t1 VDD1.n58 149.524
R414 VDD1.n40 VDD1.n39 104.615
R415 VDD1.n39 VDD1.n3 104.615
R416 VDD1.n7 VDD1.n3 104.615
R417 VDD1.n31 VDD1.n7 104.615
R418 VDD1.n31 VDD1.n30 104.615
R419 VDD1.n30 VDD1.n8 104.615
R420 VDD1.n23 VDD1.n8 104.615
R421 VDD1.n23 VDD1.n22 104.615
R422 VDD1.n22 VDD1.n12 104.615
R423 VDD1.n15 VDD1.n12 104.615
R424 VDD1.n59 VDD1.n56 104.615
R425 VDD1.n66 VDD1.n56 104.615
R426 VDD1.n67 VDD1.n66 104.615
R427 VDD1.n67 VDD1.n52 104.615
R428 VDD1.n74 VDD1.n52 104.615
R429 VDD1.n76 VDD1.n74 104.615
R430 VDD1.n76 VDD1.n75 104.615
R431 VDD1.n75 VDD1.n48 104.615
R432 VDD1.n84 VDD1.n48 104.615
R433 VDD1.n85 VDD1.n84 104.615
R434 VDD1.n91 VDD1.n90 66.5987
R435 VDD1.n93 VDD1.n92 65.7683
R436 VDD1 VDD1.n44 53.9069
R437 VDD1.n91 VDD1.n89 53.7934
R438 VDD1.n15 VDD1.t3 52.3082
R439 VDD1.n59 VDD1.t1 52.3082
R440 VDD1.n93 VDD1.n91 45.0332
R441 VDD1.n38 VDD1.n37 13.1884
R442 VDD1.n83 VDD1.n82 13.1884
R443 VDD1.n41 VDD1.n2 12.8005
R444 VDD1.n36 VDD1.n4 12.8005
R445 VDD1.n81 VDD1.n49 12.8005
R446 VDD1.n86 VDD1.n47 12.8005
R447 VDD1.n42 VDD1.n0 12.0247
R448 VDD1.n33 VDD1.n32 12.0247
R449 VDD1.n78 VDD1.n77 12.0247
R450 VDD1.n87 VDD1.n45 12.0247
R451 VDD1.n29 VDD1.n6 11.249
R452 VDD1.n73 VDD1.n51 11.249
R453 VDD1.n28 VDD1.n9 10.4732
R454 VDD1.n72 VDD1.n53 10.4732
R455 VDD1.n16 VDD1.n14 10.2747
R456 VDD1.n60 VDD1.n58 10.2747
R457 VDD1.n25 VDD1.n24 9.69747
R458 VDD1.n69 VDD1.n68 9.69747
R459 VDD1.n44 VDD1.n43 9.45567
R460 VDD1.n89 VDD1.n88 9.45567
R461 VDD1.n18 VDD1.n17 9.3005
R462 VDD1.n20 VDD1.n19 9.3005
R463 VDD1.n11 VDD1.n10 9.3005
R464 VDD1.n26 VDD1.n25 9.3005
R465 VDD1.n28 VDD1.n27 9.3005
R466 VDD1.n6 VDD1.n5 9.3005
R467 VDD1.n34 VDD1.n33 9.3005
R468 VDD1.n36 VDD1.n35 9.3005
R469 VDD1.n43 VDD1.n42 9.3005
R470 VDD1.n2 VDD1.n1 9.3005
R471 VDD1.n88 VDD1.n87 9.3005
R472 VDD1.n47 VDD1.n46 9.3005
R473 VDD1.n62 VDD1.n61 9.3005
R474 VDD1.n64 VDD1.n63 9.3005
R475 VDD1.n55 VDD1.n54 9.3005
R476 VDD1.n70 VDD1.n69 9.3005
R477 VDD1.n72 VDD1.n71 9.3005
R478 VDD1.n51 VDD1.n50 9.3005
R479 VDD1.n79 VDD1.n78 9.3005
R480 VDD1.n81 VDD1.n80 9.3005
R481 VDD1.n21 VDD1.n11 8.92171
R482 VDD1.n65 VDD1.n55 8.92171
R483 VDD1.n20 VDD1.n13 8.14595
R484 VDD1.n64 VDD1.n57 8.14595
R485 VDD1.n17 VDD1.n16 7.3702
R486 VDD1.n61 VDD1.n60 7.3702
R487 VDD1.n17 VDD1.n13 5.81868
R488 VDD1.n61 VDD1.n57 5.81868
R489 VDD1.n21 VDD1.n20 5.04292
R490 VDD1.n65 VDD1.n64 5.04292
R491 VDD1.n24 VDD1.n11 4.26717
R492 VDD1.n68 VDD1.n55 4.26717
R493 VDD1.n25 VDD1.n9 3.49141
R494 VDD1.n69 VDD1.n53 3.49141
R495 VDD1.n62 VDD1.n58 2.84303
R496 VDD1.n18 VDD1.n14 2.84303
R497 VDD1.n29 VDD1.n28 2.71565
R498 VDD1.n73 VDD1.n72 2.71565
R499 VDD1.n92 VDD1.t0 2.29217
R500 VDD1.n92 VDD1.t5 2.29217
R501 VDD1.n90 VDD1.t2 2.29217
R502 VDD1.n90 VDD1.t4 2.29217
R503 VDD1.n44 VDD1.n0 1.93989
R504 VDD1.n32 VDD1.n6 1.93989
R505 VDD1.n77 VDD1.n51 1.93989
R506 VDD1.n89 VDD1.n45 1.93989
R507 VDD1.n42 VDD1.n41 1.16414
R508 VDD1.n33 VDD1.n4 1.16414
R509 VDD1.n78 VDD1.n49 1.16414
R510 VDD1.n87 VDD1.n86 1.16414
R511 VDD1 VDD1.n93 0.828086
R512 VDD1.n38 VDD1.n2 0.388379
R513 VDD1.n37 VDD1.n36 0.388379
R514 VDD1.n82 VDD1.n81 0.388379
R515 VDD1.n83 VDD1.n47 0.388379
R516 VDD1.n43 VDD1.n1 0.155672
R517 VDD1.n35 VDD1.n1 0.155672
R518 VDD1.n35 VDD1.n34 0.155672
R519 VDD1.n34 VDD1.n5 0.155672
R520 VDD1.n27 VDD1.n5 0.155672
R521 VDD1.n27 VDD1.n26 0.155672
R522 VDD1.n26 VDD1.n10 0.155672
R523 VDD1.n19 VDD1.n10 0.155672
R524 VDD1.n19 VDD1.n18 0.155672
R525 VDD1.n63 VDD1.n62 0.155672
R526 VDD1.n63 VDD1.n54 0.155672
R527 VDD1.n70 VDD1.n54 0.155672
R528 VDD1.n71 VDD1.n70 0.155672
R529 VDD1.n71 VDD1.n50 0.155672
R530 VDD1.n79 VDD1.n50 0.155672
R531 VDD1.n80 VDD1.n79 0.155672
R532 VDD1.n80 VDD1.n46 0.155672
R533 VDD1.n88 VDD1.n46 0.155672
R534 B.n829 B.n828 585
R535 B.n830 B.n829 585
R536 B.n288 B.n141 585
R537 B.n287 B.n286 585
R538 B.n285 B.n284 585
R539 B.n283 B.n282 585
R540 B.n281 B.n280 585
R541 B.n279 B.n278 585
R542 B.n277 B.n276 585
R543 B.n275 B.n274 585
R544 B.n273 B.n272 585
R545 B.n271 B.n270 585
R546 B.n269 B.n268 585
R547 B.n267 B.n266 585
R548 B.n265 B.n264 585
R549 B.n263 B.n262 585
R550 B.n261 B.n260 585
R551 B.n259 B.n258 585
R552 B.n257 B.n256 585
R553 B.n255 B.n254 585
R554 B.n253 B.n252 585
R555 B.n251 B.n250 585
R556 B.n249 B.n248 585
R557 B.n247 B.n246 585
R558 B.n245 B.n244 585
R559 B.n243 B.n242 585
R560 B.n241 B.n240 585
R561 B.n239 B.n238 585
R562 B.n237 B.n236 585
R563 B.n235 B.n234 585
R564 B.n233 B.n232 585
R565 B.n231 B.n230 585
R566 B.n229 B.n228 585
R567 B.n226 B.n225 585
R568 B.n224 B.n223 585
R569 B.n222 B.n221 585
R570 B.n220 B.n219 585
R571 B.n218 B.n217 585
R572 B.n216 B.n215 585
R573 B.n214 B.n213 585
R574 B.n212 B.n211 585
R575 B.n210 B.n209 585
R576 B.n208 B.n207 585
R577 B.n206 B.n205 585
R578 B.n204 B.n203 585
R579 B.n202 B.n201 585
R580 B.n200 B.n199 585
R581 B.n198 B.n197 585
R582 B.n196 B.n195 585
R583 B.n194 B.n193 585
R584 B.n192 B.n191 585
R585 B.n190 B.n189 585
R586 B.n188 B.n187 585
R587 B.n186 B.n185 585
R588 B.n184 B.n183 585
R589 B.n182 B.n181 585
R590 B.n180 B.n179 585
R591 B.n178 B.n177 585
R592 B.n176 B.n175 585
R593 B.n174 B.n173 585
R594 B.n172 B.n171 585
R595 B.n170 B.n169 585
R596 B.n168 B.n167 585
R597 B.n166 B.n165 585
R598 B.n164 B.n163 585
R599 B.n162 B.n161 585
R600 B.n160 B.n159 585
R601 B.n158 B.n157 585
R602 B.n156 B.n155 585
R603 B.n154 B.n153 585
R604 B.n152 B.n151 585
R605 B.n150 B.n149 585
R606 B.n148 B.n147 585
R607 B.n103 B.n102 585
R608 B.n827 B.n104 585
R609 B.n831 B.n104 585
R610 B.n826 B.n825 585
R611 B.n825 B.n100 585
R612 B.n824 B.n99 585
R613 B.n837 B.n99 585
R614 B.n823 B.n98 585
R615 B.n838 B.n98 585
R616 B.n822 B.n97 585
R617 B.n839 B.n97 585
R618 B.n821 B.n820 585
R619 B.n820 B.n93 585
R620 B.n819 B.n92 585
R621 B.n845 B.n92 585
R622 B.n818 B.n91 585
R623 B.n846 B.n91 585
R624 B.n817 B.n90 585
R625 B.n847 B.n90 585
R626 B.n816 B.n815 585
R627 B.n815 B.n89 585
R628 B.n814 B.n85 585
R629 B.n853 B.n85 585
R630 B.n813 B.n84 585
R631 B.n854 B.n84 585
R632 B.n812 B.n83 585
R633 B.n855 B.n83 585
R634 B.n811 B.n810 585
R635 B.n810 B.n79 585
R636 B.n809 B.n78 585
R637 B.n861 B.n78 585
R638 B.n808 B.n77 585
R639 B.n862 B.n77 585
R640 B.n807 B.n76 585
R641 B.n863 B.n76 585
R642 B.n806 B.n805 585
R643 B.n805 B.n72 585
R644 B.n804 B.n71 585
R645 B.n869 B.n71 585
R646 B.n803 B.n70 585
R647 B.n870 B.n70 585
R648 B.n802 B.n69 585
R649 B.n871 B.n69 585
R650 B.n801 B.n800 585
R651 B.n800 B.n65 585
R652 B.n799 B.n64 585
R653 B.n877 B.n64 585
R654 B.n798 B.n63 585
R655 B.n878 B.n63 585
R656 B.n797 B.n62 585
R657 B.n879 B.n62 585
R658 B.n796 B.n795 585
R659 B.n795 B.n58 585
R660 B.n794 B.n57 585
R661 B.n885 B.n57 585
R662 B.n793 B.n56 585
R663 B.n886 B.n56 585
R664 B.n792 B.n55 585
R665 B.n887 B.n55 585
R666 B.n791 B.n790 585
R667 B.n790 B.n51 585
R668 B.n789 B.n50 585
R669 B.n893 B.n50 585
R670 B.n788 B.n49 585
R671 B.n894 B.n49 585
R672 B.n787 B.n48 585
R673 B.n895 B.n48 585
R674 B.n786 B.n785 585
R675 B.n785 B.n44 585
R676 B.n784 B.n43 585
R677 B.n901 B.n43 585
R678 B.n783 B.n42 585
R679 B.n902 B.n42 585
R680 B.n782 B.n41 585
R681 B.n903 B.n41 585
R682 B.n781 B.n780 585
R683 B.n780 B.n37 585
R684 B.n779 B.n36 585
R685 B.n909 B.n36 585
R686 B.n778 B.n35 585
R687 B.n910 B.n35 585
R688 B.n777 B.n34 585
R689 B.n911 B.n34 585
R690 B.n776 B.n775 585
R691 B.n775 B.n30 585
R692 B.n774 B.n29 585
R693 B.n917 B.n29 585
R694 B.n773 B.n28 585
R695 B.n918 B.n28 585
R696 B.n772 B.n27 585
R697 B.n919 B.n27 585
R698 B.n771 B.n770 585
R699 B.n770 B.n23 585
R700 B.n769 B.n22 585
R701 B.n925 B.n22 585
R702 B.n768 B.n21 585
R703 B.n926 B.n21 585
R704 B.n767 B.n20 585
R705 B.n927 B.n20 585
R706 B.n766 B.n765 585
R707 B.n765 B.n16 585
R708 B.n764 B.n15 585
R709 B.n933 B.n15 585
R710 B.n763 B.n14 585
R711 B.n934 B.n14 585
R712 B.n762 B.n13 585
R713 B.n935 B.n13 585
R714 B.n761 B.n760 585
R715 B.n760 B.n12 585
R716 B.n759 B.n758 585
R717 B.n759 B.n8 585
R718 B.n757 B.n7 585
R719 B.n942 B.n7 585
R720 B.n756 B.n6 585
R721 B.n943 B.n6 585
R722 B.n755 B.n5 585
R723 B.n944 B.n5 585
R724 B.n754 B.n753 585
R725 B.n753 B.n4 585
R726 B.n752 B.n289 585
R727 B.n752 B.n751 585
R728 B.n742 B.n290 585
R729 B.n291 B.n290 585
R730 B.n744 B.n743 585
R731 B.n745 B.n744 585
R732 B.n741 B.n296 585
R733 B.n296 B.n295 585
R734 B.n740 B.n739 585
R735 B.n739 B.n738 585
R736 B.n298 B.n297 585
R737 B.n299 B.n298 585
R738 B.n731 B.n730 585
R739 B.n732 B.n731 585
R740 B.n729 B.n304 585
R741 B.n304 B.n303 585
R742 B.n728 B.n727 585
R743 B.n727 B.n726 585
R744 B.n306 B.n305 585
R745 B.n307 B.n306 585
R746 B.n719 B.n718 585
R747 B.n720 B.n719 585
R748 B.n717 B.n312 585
R749 B.n312 B.n311 585
R750 B.n716 B.n715 585
R751 B.n715 B.n714 585
R752 B.n314 B.n313 585
R753 B.n315 B.n314 585
R754 B.n707 B.n706 585
R755 B.n708 B.n707 585
R756 B.n705 B.n320 585
R757 B.n320 B.n319 585
R758 B.n704 B.n703 585
R759 B.n703 B.n702 585
R760 B.n322 B.n321 585
R761 B.n323 B.n322 585
R762 B.n695 B.n694 585
R763 B.n696 B.n695 585
R764 B.n693 B.n328 585
R765 B.n328 B.n327 585
R766 B.n692 B.n691 585
R767 B.n691 B.n690 585
R768 B.n330 B.n329 585
R769 B.n331 B.n330 585
R770 B.n683 B.n682 585
R771 B.n684 B.n683 585
R772 B.n681 B.n336 585
R773 B.n336 B.n335 585
R774 B.n680 B.n679 585
R775 B.n679 B.n678 585
R776 B.n338 B.n337 585
R777 B.n339 B.n338 585
R778 B.n671 B.n670 585
R779 B.n672 B.n671 585
R780 B.n669 B.n344 585
R781 B.n344 B.n343 585
R782 B.n668 B.n667 585
R783 B.n667 B.n666 585
R784 B.n346 B.n345 585
R785 B.n347 B.n346 585
R786 B.n659 B.n658 585
R787 B.n660 B.n659 585
R788 B.n657 B.n352 585
R789 B.n352 B.n351 585
R790 B.n656 B.n655 585
R791 B.n655 B.n654 585
R792 B.n354 B.n353 585
R793 B.n355 B.n354 585
R794 B.n647 B.n646 585
R795 B.n648 B.n647 585
R796 B.n645 B.n360 585
R797 B.n360 B.n359 585
R798 B.n644 B.n643 585
R799 B.n643 B.n642 585
R800 B.n362 B.n361 585
R801 B.n363 B.n362 585
R802 B.n635 B.n634 585
R803 B.n636 B.n635 585
R804 B.n633 B.n368 585
R805 B.n368 B.n367 585
R806 B.n632 B.n631 585
R807 B.n631 B.n630 585
R808 B.n370 B.n369 585
R809 B.n371 B.n370 585
R810 B.n623 B.n622 585
R811 B.n624 B.n623 585
R812 B.n621 B.n376 585
R813 B.n376 B.n375 585
R814 B.n620 B.n619 585
R815 B.n619 B.n618 585
R816 B.n378 B.n377 585
R817 B.n611 B.n378 585
R818 B.n610 B.n609 585
R819 B.n612 B.n610 585
R820 B.n608 B.n383 585
R821 B.n383 B.n382 585
R822 B.n607 B.n606 585
R823 B.n606 B.n605 585
R824 B.n385 B.n384 585
R825 B.n386 B.n385 585
R826 B.n598 B.n597 585
R827 B.n599 B.n598 585
R828 B.n596 B.n391 585
R829 B.n391 B.n390 585
R830 B.n595 B.n594 585
R831 B.n594 B.n593 585
R832 B.n393 B.n392 585
R833 B.n394 B.n393 585
R834 B.n586 B.n585 585
R835 B.n587 B.n586 585
R836 B.n397 B.n396 585
R837 B.n441 B.n439 585
R838 B.n442 B.n438 585
R839 B.n442 B.n398 585
R840 B.n445 B.n444 585
R841 B.n446 B.n437 585
R842 B.n448 B.n447 585
R843 B.n450 B.n436 585
R844 B.n453 B.n452 585
R845 B.n454 B.n435 585
R846 B.n456 B.n455 585
R847 B.n458 B.n434 585
R848 B.n461 B.n460 585
R849 B.n462 B.n433 585
R850 B.n464 B.n463 585
R851 B.n466 B.n432 585
R852 B.n469 B.n468 585
R853 B.n470 B.n431 585
R854 B.n472 B.n471 585
R855 B.n474 B.n430 585
R856 B.n477 B.n476 585
R857 B.n478 B.n429 585
R858 B.n480 B.n479 585
R859 B.n482 B.n428 585
R860 B.n485 B.n484 585
R861 B.n486 B.n427 585
R862 B.n488 B.n487 585
R863 B.n490 B.n426 585
R864 B.n493 B.n492 585
R865 B.n494 B.n425 585
R866 B.n496 B.n495 585
R867 B.n498 B.n424 585
R868 B.n501 B.n500 585
R869 B.n503 B.n421 585
R870 B.n505 B.n504 585
R871 B.n507 B.n420 585
R872 B.n510 B.n509 585
R873 B.n511 B.n419 585
R874 B.n513 B.n512 585
R875 B.n515 B.n418 585
R876 B.n518 B.n517 585
R877 B.n519 B.n415 585
R878 B.n522 B.n521 585
R879 B.n524 B.n414 585
R880 B.n527 B.n526 585
R881 B.n528 B.n413 585
R882 B.n530 B.n529 585
R883 B.n532 B.n412 585
R884 B.n535 B.n534 585
R885 B.n536 B.n411 585
R886 B.n538 B.n537 585
R887 B.n540 B.n410 585
R888 B.n543 B.n542 585
R889 B.n544 B.n409 585
R890 B.n546 B.n545 585
R891 B.n548 B.n408 585
R892 B.n551 B.n550 585
R893 B.n552 B.n407 585
R894 B.n554 B.n553 585
R895 B.n556 B.n406 585
R896 B.n559 B.n558 585
R897 B.n560 B.n405 585
R898 B.n562 B.n561 585
R899 B.n564 B.n404 585
R900 B.n567 B.n566 585
R901 B.n568 B.n403 585
R902 B.n570 B.n569 585
R903 B.n572 B.n402 585
R904 B.n575 B.n574 585
R905 B.n576 B.n401 585
R906 B.n578 B.n577 585
R907 B.n580 B.n400 585
R908 B.n583 B.n582 585
R909 B.n584 B.n399 585
R910 B.n589 B.n588 585
R911 B.n588 B.n587 585
R912 B.n590 B.n395 585
R913 B.n395 B.n394 585
R914 B.n592 B.n591 585
R915 B.n593 B.n592 585
R916 B.n389 B.n388 585
R917 B.n390 B.n389 585
R918 B.n601 B.n600 585
R919 B.n600 B.n599 585
R920 B.n602 B.n387 585
R921 B.n387 B.n386 585
R922 B.n604 B.n603 585
R923 B.n605 B.n604 585
R924 B.n381 B.n380 585
R925 B.n382 B.n381 585
R926 B.n614 B.n613 585
R927 B.n613 B.n612 585
R928 B.n615 B.n379 585
R929 B.n611 B.n379 585
R930 B.n617 B.n616 585
R931 B.n618 B.n617 585
R932 B.n374 B.n373 585
R933 B.n375 B.n374 585
R934 B.n626 B.n625 585
R935 B.n625 B.n624 585
R936 B.n627 B.n372 585
R937 B.n372 B.n371 585
R938 B.n629 B.n628 585
R939 B.n630 B.n629 585
R940 B.n366 B.n365 585
R941 B.n367 B.n366 585
R942 B.n638 B.n637 585
R943 B.n637 B.n636 585
R944 B.n639 B.n364 585
R945 B.n364 B.n363 585
R946 B.n641 B.n640 585
R947 B.n642 B.n641 585
R948 B.n358 B.n357 585
R949 B.n359 B.n358 585
R950 B.n650 B.n649 585
R951 B.n649 B.n648 585
R952 B.n651 B.n356 585
R953 B.n356 B.n355 585
R954 B.n653 B.n652 585
R955 B.n654 B.n653 585
R956 B.n350 B.n349 585
R957 B.n351 B.n350 585
R958 B.n662 B.n661 585
R959 B.n661 B.n660 585
R960 B.n663 B.n348 585
R961 B.n348 B.n347 585
R962 B.n665 B.n664 585
R963 B.n666 B.n665 585
R964 B.n342 B.n341 585
R965 B.n343 B.n342 585
R966 B.n674 B.n673 585
R967 B.n673 B.n672 585
R968 B.n675 B.n340 585
R969 B.n340 B.n339 585
R970 B.n677 B.n676 585
R971 B.n678 B.n677 585
R972 B.n334 B.n333 585
R973 B.n335 B.n334 585
R974 B.n686 B.n685 585
R975 B.n685 B.n684 585
R976 B.n687 B.n332 585
R977 B.n332 B.n331 585
R978 B.n689 B.n688 585
R979 B.n690 B.n689 585
R980 B.n326 B.n325 585
R981 B.n327 B.n326 585
R982 B.n698 B.n697 585
R983 B.n697 B.n696 585
R984 B.n699 B.n324 585
R985 B.n324 B.n323 585
R986 B.n701 B.n700 585
R987 B.n702 B.n701 585
R988 B.n318 B.n317 585
R989 B.n319 B.n318 585
R990 B.n710 B.n709 585
R991 B.n709 B.n708 585
R992 B.n711 B.n316 585
R993 B.n316 B.n315 585
R994 B.n713 B.n712 585
R995 B.n714 B.n713 585
R996 B.n310 B.n309 585
R997 B.n311 B.n310 585
R998 B.n722 B.n721 585
R999 B.n721 B.n720 585
R1000 B.n723 B.n308 585
R1001 B.n308 B.n307 585
R1002 B.n725 B.n724 585
R1003 B.n726 B.n725 585
R1004 B.n302 B.n301 585
R1005 B.n303 B.n302 585
R1006 B.n734 B.n733 585
R1007 B.n733 B.n732 585
R1008 B.n735 B.n300 585
R1009 B.n300 B.n299 585
R1010 B.n737 B.n736 585
R1011 B.n738 B.n737 585
R1012 B.n294 B.n293 585
R1013 B.n295 B.n294 585
R1014 B.n747 B.n746 585
R1015 B.n746 B.n745 585
R1016 B.n748 B.n292 585
R1017 B.n292 B.n291 585
R1018 B.n750 B.n749 585
R1019 B.n751 B.n750 585
R1020 B.n3 B.n0 585
R1021 B.n4 B.n3 585
R1022 B.n941 B.n1 585
R1023 B.n942 B.n941 585
R1024 B.n940 B.n939 585
R1025 B.n940 B.n8 585
R1026 B.n938 B.n9 585
R1027 B.n12 B.n9 585
R1028 B.n937 B.n936 585
R1029 B.n936 B.n935 585
R1030 B.n11 B.n10 585
R1031 B.n934 B.n11 585
R1032 B.n932 B.n931 585
R1033 B.n933 B.n932 585
R1034 B.n930 B.n17 585
R1035 B.n17 B.n16 585
R1036 B.n929 B.n928 585
R1037 B.n928 B.n927 585
R1038 B.n19 B.n18 585
R1039 B.n926 B.n19 585
R1040 B.n924 B.n923 585
R1041 B.n925 B.n924 585
R1042 B.n922 B.n24 585
R1043 B.n24 B.n23 585
R1044 B.n921 B.n920 585
R1045 B.n920 B.n919 585
R1046 B.n26 B.n25 585
R1047 B.n918 B.n26 585
R1048 B.n916 B.n915 585
R1049 B.n917 B.n916 585
R1050 B.n914 B.n31 585
R1051 B.n31 B.n30 585
R1052 B.n913 B.n912 585
R1053 B.n912 B.n911 585
R1054 B.n33 B.n32 585
R1055 B.n910 B.n33 585
R1056 B.n908 B.n907 585
R1057 B.n909 B.n908 585
R1058 B.n906 B.n38 585
R1059 B.n38 B.n37 585
R1060 B.n905 B.n904 585
R1061 B.n904 B.n903 585
R1062 B.n40 B.n39 585
R1063 B.n902 B.n40 585
R1064 B.n900 B.n899 585
R1065 B.n901 B.n900 585
R1066 B.n898 B.n45 585
R1067 B.n45 B.n44 585
R1068 B.n897 B.n896 585
R1069 B.n896 B.n895 585
R1070 B.n47 B.n46 585
R1071 B.n894 B.n47 585
R1072 B.n892 B.n891 585
R1073 B.n893 B.n892 585
R1074 B.n890 B.n52 585
R1075 B.n52 B.n51 585
R1076 B.n889 B.n888 585
R1077 B.n888 B.n887 585
R1078 B.n54 B.n53 585
R1079 B.n886 B.n54 585
R1080 B.n884 B.n883 585
R1081 B.n885 B.n884 585
R1082 B.n882 B.n59 585
R1083 B.n59 B.n58 585
R1084 B.n881 B.n880 585
R1085 B.n880 B.n879 585
R1086 B.n61 B.n60 585
R1087 B.n878 B.n61 585
R1088 B.n876 B.n875 585
R1089 B.n877 B.n876 585
R1090 B.n874 B.n66 585
R1091 B.n66 B.n65 585
R1092 B.n873 B.n872 585
R1093 B.n872 B.n871 585
R1094 B.n68 B.n67 585
R1095 B.n870 B.n68 585
R1096 B.n868 B.n867 585
R1097 B.n869 B.n868 585
R1098 B.n866 B.n73 585
R1099 B.n73 B.n72 585
R1100 B.n865 B.n864 585
R1101 B.n864 B.n863 585
R1102 B.n75 B.n74 585
R1103 B.n862 B.n75 585
R1104 B.n860 B.n859 585
R1105 B.n861 B.n860 585
R1106 B.n858 B.n80 585
R1107 B.n80 B.n79 585
R1108 B.n857 B.n856 585
R1109 B.n856 B.n855 585
R1110 B.n82 B.n81 585
R1111 B.n854 B.n82 585
R1112 B.n852 B.n851 585
R1113 B.n853 B.n852 585
R1114 B.n850 B.n86 585
R1115 B.n89 B.n86 585
R1116 B.n849 B.n848 585
R1117 B.n848 B.n847 585
R1118 B.n88 B.n87 585
R1119 B.n846 B.n88 585
R1120 B.n844 B.n843 585
R1121 B.n845 B.n844 585
R1122 B.n842 B.n94 585
R1123 B.n94 B.n93 585
R1124 B.n841 B.n840 585
R1125 B.n840 B.n839 585
R1126 B.n96 B.n95 585
R1127 B.n838 B.n96 585
R1128 B.n836 B.n835 585
R1129 B.n837 B.n836 585
R1130 B.n834 B.n101 585
R1131 B.n101 B.n100 585
R1132 B.n833 B.n832 585
R1133 B.n832 B.n831 585
R1134 B.n945 B.n944 585
R1135 B.n943 B.n2 585
R1136 B.n832 B.n103 497.305
R1137 B.n829 B.n104 497.305
R1138 B.n586 B.n399 497.305
R1139 B.n588 B.n397 497.305
R1140 B.n142 B.t18 303.933
R1141 B.n416 B.t13 303.933
R1142 B.n144 B.t8 303.933
R1143 B.n422 B.t16 303.933
R1144 B.n144 B.t6 264.414
R1145 B.n142 B.t17 264.414
R1146 B.n416 B.t10 264.414
R1147 B.n422 B.t14 264.414
R1148 B.n830 B.n140 256.663
R1149 B.n830 B.n139 256.663
R1150 B.n830 B.n138 256.663
R1151 B.n830 B.n137 256.663
R1152 B.n830 B.n136 256.663
R1153 B.n830 B.n135 256.663
R1154 B.n830 B.n134 256.663
R1155 B.n830 B.n133 256.663
R1156 B.n830 B.n132 256.663
R1157 B.n830 B.n131 256.663
R1158 B.n830 B.n130 256.663
R1159 B.n830 B.n129 256.663
R1160 B.n830 B.n128 256.663
R1161 B.n830 B.n127 256.663
R1162 B.n830 B.n126 256.663
R1163 B.n830 B.n125 256.663
R1164 B.n830 B.n124 256.663
R1165 B.n830 B.n123 256.663
R1166 B.n830 B.n122 256.663
R1167 B.n830 B.n121 256.663
R1168 B.n830 B.n120 256.663
R1169 B.n830 B.n119 256.663
R1170 B.n830 B.n118 256.663
R1171 B.n830 B.n117 256.663
R1172 B.n830 B.n116 256.663
R1173 B.n830 B.n115 256.663
R1174 B.n830 B.n114 256.663
R1175 B.n830 B.n113 256.663
R1176 B.n830 B.n112 256.663
R1177 B.n830 B.n111 256.663
R1178 B.n830 B.n110 256.663
R1179 B.n830 B.n109 256.663
R1180 B.n830 B.n108 256.663
R1181 B.n830 B.n107 256.663
R1182 B.n830 B.n106 256.663
R1183 B.n830 B.n105 256.663
R1184 B.n440 B.n398 256.663
R1185 B.n443 B.n398 256.663
R1186 B.n449 B.n398 256.663
R1187 B.n451 B.n398 256.663
R1188 B.n457 B.n398 256.663
R1189 B.n459 B.n398 256.663
R1190 B.n465 B.n398 256.663
R1191 B.n467 B.n398 256.663
R1192 B.n473 B.n398 256.663
R1193 B.n475 B.n398 256.663
R1194 B.n481 B.n398 256.663
R1195 B.n483 B.n398 256.663
R1196 B.n489 B.n398 256.663
R1197 B.n491 B.n398 256.663
R1198 B.n497 B.n398 256.663
R1199 B.n499 B.n398 256.663
R1200 B.n506 B.n398 256.663
R1201 B.n508 B.n398 256.663
R1202 B.n514 B.n398 256.663
R1203 B.n516 B.n398 256.663
R1204 B.n523 B.n398 256.663
R1205 B.n525 B.n398 256.663
R1206 B.n531 B.n398 256.663
R1207 B.n533 B.n398 256.663
R1208 B.n539 B.n398 256.663
R1209 B.n541 B.n398 256.663
R1210 B.n547 B.n398 256.663
R1211 B.n549 B.n398 256.663
R1212 B.n555 B.n398 256.663
R1213 B.n557 B.n398 256.663
R1214 B.n563 B.n398 256.663
R1215 B.n565 B.n398 256.663
R1216 B.n571 B.n398 256.663
R1217 B.n573 B.n398 256.663
R1218 B.n579 B.n398 256.663
R1219 B.n581 B.n398 256.663
R1220 B.n947 B.n946 256.663
R1221 B.n143 B.t19 224.225
R1222 B.n417 B.t12 224.225
R1223 B.n145 B.t9 224.225
R1224 B.n423 B.t15 224.225
R1225 B.n149 B.n148 163.367
R1226 B.n153 B.n152 163.367
R1227 B.n157 B.n156 163.367
R1228 B.n161 B.n160 163.367
R1229 B.n165 B.n164 163.367
R1230 B.n169 B.n168 163.367
R1231 B.n173 B.n172 163.367
R1232 B.n177 B.n176 163.367
R1233 B.n181 B.n180 163.367
R1234 B.n185 B.n184 163.367
R1235 B.n189 B.n188 163.367
R1236 B.n193 B.n192 163.367
R1237 B.n197 B.n196 163.367
R1238 B.n201 B.n200 163.367
R1239 B.n205 B.n204 163.367
R1240 B.n209 B.n208 163.367
R1241 B.n213 B.n212 163.367
R1242 B.n217 B.n216 163.367
R1243 B.n221 B.n220 163.367
R1244 B.n225 B.n224 163.367
R1245 B.n230 B.n229 163.367
R1246 B.n234 B.n233 163.367
R1247 B.n238 B.n237 163.367
R1248 B.n242 B.n241 163.367
R1249 B.n246 B.n245 163.367
R1250 B.n250 B.n249 163.367
R1251 B.n254 B.n253 163.367
R1252 B.n258 B.n257 163.367
R1253 B.n262 B.n261 163.367
R1254 B.n266 B.n265 163.367
R1255 B.n270 B.n269 163.367
R1256 B.n274 B.n273 163.367
R1257 B.n278 B.n277 163.367
R1258 B.n282 B.n281 163.367
R1259 B.n286 B.n285 163.367
R1260 B.n829 B.n141 163.367
R1261 B.n586 B.n393 163.367
R1262 B.n594 B.n393 163.367
R1263 B.n594 B.n391 163.367
R1264 B.n598 B.n391 163.367
R1265 B.n598 B.n385 163.367
R1266 B.n606 B.n385 163.367
R1267 B.n606 B.n383 163.367
R1268 B.n610 B.n383 163.367
R1269 B.n610 B.n378 163.367
R1270 B.n619 B.n378 163.367
R1271 B.n619 B.n376 163.367
R1272 B.n623 B.n376 163.367
R1273 B.n623 B.n370 163.367
R1274 B.n631 B.n370 163.367
R1275 B.n631 B.n368 163.367
R1276 B.n635 B.n368 163.367
R1277 B.n635 B.n362 163.367
R1278 B.n643 B.n362 163.367
R1279 B.n643 B.n360 163.367
R1280 B.n647 B.n360 163.367
R1281 B.n647 B.n354 163.367
R1282 B.n655 B.n354 163.367
R1283 B.n655 B.n352 163.367
R1284 B.n659 B.n352 163.367
R1285 B.n659 B.n346 163.367
R1286 B.n667 B.n346 163.367
R1287 B.n667 B.n344 163.367
R1288 B.n671 B.n344 163.367
R1289 B.n671 B.n338 163.367
R1290 B.n679 B.n338 163.367
R1291 B.n679 B.n336 163.367
R1292 B.n683 B.n336 163.367
R1293 B.n683 B.n330 163.367
R1294 B.n691 B.n330 163.367
R1295 B.n691 B.n328 163.367
R1296 B.n695 B.n328 163.367
R1297 B.n695 B.n322 163.367
R1298 B.n703 B.n322 163.367
R1299 B.n703 B.n320 163.367
R1300 B.n707 B.n320 163.367
R1301 B.n707 B.n314 163.367
R1302 B.n715 B.n314 163.367
R1303 B.n715 B.n312 163.367
R1304 B.n719 B.n312 163.367
R1305 B.n719 B.n306 163.367
R1306 B.n727 B.n306 163.367
R1307 B.n727 B.n304 163.367
R1308 B.n731 B.n304 163.367
R1309 B.n731 B.n298 163.367
R1310 B.n739 B.n298 163.367
R1311 B.n739 B.n296 163.367
R1312 B.n744 B.n296 163.367
R1313 B.n744 B.n290 163.367
R1314 B.n752 B.n290 163.367
R1315 B.n753 B.n752 163.367
R1316 B.n753 B.n5 163.367
R1317 B.n6 B.n5 163.367
R1318 B.n7 B.n6 163.367
R1319 B.n759 B.n7 163.367
R1320 B.n760 B.n759 163.367
R1321 B.n760 B.n13 163.367
R1322 B.n14 B.n13 163.367
R1323 B.n15 B.n14 163.367
R1324 B.n765 B.n15 163.367
R1325 B.n765 B.n20 163.367
R1326 B.n21 B.n20 163.367
R1327 B.n22 B.n21 163.367
R1328 B.n770 B.n22 163.367
R1329 B.n770 B.n27 163.367
R1330 B.n28 B.n27 163.367
R1331 B.n29 B.n28 163.367
R1332 B.n775 B.n29 163.367
R1333 B.n775 B.n34 163.367
R1334 B.n35 B.n34 163.367
R1335 B.n36 B.n35 163.367
R1336 B.n780 B.n36 163.367
R1337 B.n780 B.n41 163.367
R1338 B.n42 B.n41 163.367
R1339 B.n43 B.n42 163.367
R1340 B.n785 B.n43 163.367
R1341 B.n785 B.n48 163.367
R1342 B.n49 B.n48 163.367
R1343 B.n50 B.n49 163.367
R1344 B.n790 B.n50 163.367
R1345 B.n790 B.n55 163.367
R1346 B.n56 B.n55 163.367
R1347 B.n57 B.n56 163.367
R1348 B.n795 B.n57 163.367
R1349 B.n795 B.n62 163.367
R1350 B.n63 B.n62 163.367
R1351 B.n64 B.n63 163.367
R1352 B.n800 B.n64 163.367
R1353 B.n800 B.n69 163.367
R1354 B.n70 B.n69 163.367
R1355 B.n71 B.n70 163.367
R1356 B.n805 B.n71 163.367
R1357 B.n805 B.n76 163.367
R1358 B.n77 B.n76 163.367
R1359 B.n78 B.n77 163.367
R1360 B.n810 B.n78 163.367
R1361 B.n810 B.n83 163.367
R1362 B.n84 B.n83 163.367
R1363 B.n85 B.n84 163.367
R1364 B.n815 B.n85 163.367
R1365 B.n815 B.n90 163.367
R1366 B.n91 B.n90 163.367
R1367 B.n92 B.n91 163.367
R1368 B.n820 B.n92 163.367
R1369 B.n820 B.n97 163.367
R1370 B.n98 B.n97 163.367
R1371 B.n99 B.n98 163.367
R1372 B.n825 B.n99 163.367
R1373 B.n825 B.n104 163.367
R1374 B.n442 B.n441 163.367
R1375 B.n444 B.n442 163.367
R1376 B.n448 B.n437 163.367
R1377 B.n452 B.n450 163.367
R1378 B.n456 B.n435 163.367
R1379 B.n460 B.n458 163.367
R1380 B.n464 B.n433 163.367
R1381 B.n468 B.n466 163.367
R1382 B.n472 B.n431 163.367
R1383 B.n476 B.n474 163.367
R1384 B.n480 B.n429 163.367
R1385 B.n484 B.n482 163.367
R1386 B.n488 B.n427 163.367
R1387 B.n492 B.n490 163.367
R1388 B.n496 B.n425 163.367
R1389 B.n500 B.n498 163.367
R1390 B.n505 B.n421 163.367
R1391 B.n509 B.n507 163.367
R1392 B.n513 B.n419 163.367
R1393 B.n517 B.n515 163.367
R1394 B.n522 B.n415 163.367
R1395 B.n526 B.n524 163.367
R1396 B.n530 B.n413 163.367
R1397 B.n534 B.n532 163.367
R1398 B.n538 B.n411 163.367
R1399 B.n542 B.n540 163.367
R1400 B.n546 B.n409 163.367
R1401 B.n550 B.n548 163.367
R1402 B.n554 B.n407 163.367
R1403 B.n558 B.n556 163.367
R1404 B.n562 B.n405 163.367
R1405 B.n566 B.n564 163.367
R1406 B.n570 B.n403 163.367
R1407 B.n574 B.n572 163.367
R1408 B.n578 B.n401 163.367
R1409 B.n582 B.n580 163.367
R1410 B.n588 B.n395 163.367
R1411 B.n592 B.n395 163.367
R1412 B.n592 B.n389 163.367
R1413 B.n600 B.n389 163.367
R1414 B.n600 B.n387 163.367
R1415 B.n604 B.n387 163.367
R1416 B.n604 B.n381 163.367
R1417 B.n613 B.n381 163.367
R1418 B.n613 B.n379 163.367
R1419 B.n617 B.n379 163.367
R1420 B.n617 B.n374 163.367
R1421 B.n625 B.n374 163.367
R1422 B.n625 B.n372 163.367
R1423 B.n629 B.n372 163.367
R1424 B.n629 B.n366 163.367
R1425 B.n637 B.n366 163.367
R1426 B.n637 B.n364 163.367
R1427 B.n641 B.n364 163.367
R1428 B.n641 B.n358 163.367
R1429 B.n649 B.n358 163.367
R1430 B.n649 B.n356 163.367
R1431 B.n653 B.n356 163.367
R1432 B.n653 B.n350 163.367
R1433 B.n661 B.n350 163.367
R1434 B.n661 B.n348 163.367
R1435 B.n665 B.n348 163.367
R1436 B.n665 B.n342 163.367
R1437 B.n673 B.n342 163.367
R1438 B.n673 B.n340 163.367
R1439 B.n677 B.n340 163.367
R1440 B.n677 B.n334 163.367
R1441 B.n685 B.n334 163.367
R1442 B.n685 B.n332 163.367
R1443 B.n689 B.n332 163.367
R1444 B.n689 B.n326 163.367
R1445 B.n697 B.n326 163.367
R1446 B.n697 B.n324 163.367
R1447 B.n701 B.n324 163.367
R1448 B.n701 B.n318 163.367
R1449 B.n709 B.n318 163.367
R1450 B.n709 B.n316 163.367
R1451 B.n713 B.n316 163.367
R1452 B.n713 B.n310 163.367
R1453 B.n721 B.n310 163.367
R1454 B.n721 B.n308 163.367
R1455 B.n725 B.n308 163.367
R1456 B.n725 B.n302 163.367
R1457 B.n733 B.n302 163.367
R1458 B.n733 B.n300 163.367
R1459 B.n737 B.n300 163.367
R1460 B.n737 B.n294 163.367
R1461 B.n746 B.n294 163.367
R1462 B.n746 B.n292 163.367
R1463 B.n750 B.n292 163.367
R1464 B.n750 B.n3 163.367
R1465 B.n945 B.n3 163.367
R1466 B.n941 B.n2 163.367
R1467 B.n941 B.n940 163.367
R1468 B.n940 B.n9 163.367
R1469 B.n936 B.n9 163.367
R1470 B.n936 B.n11 163.367
R1471 B.n932 B.n11 163.367
R1472 B.n932 B.n17 163.367
R1473 B.n928 B.n17 163.367
R1474 B.n928 B.n19 163.367
R1475 B.n924 B.n19 163.367
R1476 B.n924 B.n24 163.367
R1477 B.n920 B.n24 163.367
R1478 B.n920 B.n26 163.367
R1479 B.n916 B.n26 163.367
R1480 B.n916 B.n31 163.367
R1481 B.n912 B.n31 163.367
R1482 B.n912 B.n33 163.367
R1483 B.n908 B.n33 163.367
R1484 B.n908 B.n38 163.367
R1485 B.n904 B.n38 163.367
R1486 B.n904 B.n40 163.367
R1487 B.n900 B.n40 163.367
R1488 B.n900 B.n45 163.367
R1489 B.n896 B.n45 163.367
R1490 B.n896 B.n47 163.367
R1491 B.n892 B.n47 163.367
R1492 B.n892 B.n52 163.367
R1493 B.n888 B.n52 163.367
R1494 B.n888 B.n54 163.367
R1495 B.n884 B.n54 163.367
R1496 B.n884 B.n59 163.367
R1497 B.n880 B.n59 163.367
R1498 B.n880 B.n61 163.367
R1499 B.n876 B.n61 163.367
R1500 B.n876 B.n66 163.367
R1501 B.n872 B.n66 163.367
R1502 B.n872 B.n68 163.367
R1503 B.n868 B.n68 163.367
R1504 B.n868 B.n73 163.367
R1505 B.n864 B.n73 163.367
R1506 B.n864 B.n75 163.367
R1507 B.n860 B.n75 163.367
R1508 B.n860 B.n80 163.367
R1509 B.n856 B.n80 163.367
R1510 B.n856 B.n82 163.367
R1511 B.n852 B.n82 163.367
R1512 B.n852 B.n86 163.367
R1513 B.n848 B.n86 163.367
R1514 B.n848 B.n88 163.367
R1515 B.n844 B.n88 163.367
R1516 B.n844 B.n94 163.367
R1517 B.n840 B.n94 163.367
R1518 B.n840 B.n96 163.367
R1519 B.n836 B.n96 163.367
R1520 B.n836 B.n101 163.367
R1521 B.n832 B.n101 163.367
R1522 B.n587 B.n398 95.6527
R1523 B.n831 B.n830 95.6527
R1524 B.n145 B.n144 79.7096
R1525 B.n143 B.n142 79.7096
R1526 B.n417 B.n416 79.7096
R1527 B.n423 B.n422 79.7096
R1528 B.n105 B.n103 71.676
R1529 B.n149 B.n106 71.676
R1530 B.n153 B.n107 71.676
R1531 B.n157 B.n108 71.676
R1532 B.n161 B.n109 71.676
R1533 B.n165 B.n110 71.676
R1534 B.n169 B.n111 71.676
R1535 B.n173 B.n112 71.676
R1536 B.n177 B.n113 71.676
R1537 B.n181 B.n114 71.676
R1538 B.n185 B.n115 71.676
R1539 B.n189 B.n116 71.676
R1540 B.n193 B.n117 71.676
R1541 B.n197 B.n118 71.676
R1542 B.n201 B.n119 71.676
R1543 B.n205 B.n120 71.676
R1544 B.n209 B.n121 71.676
R1545 B.n213 B.n122 71.676
R1546 B.n217 B.n123 71.676
R1547 B.n221 B.n124 71.676
R1548 B.n225 B.n125 71.676
R1549 B.n230 B.n126 71.676
R1550 B.n234 B.n127 71.676
R1551 B.n238 B.n128 71.676
R1552 B.n242 B.n129 71.676
R1553 B.n246 B.n130 71.676
R1554 B.n250 B.n131 71.676
R1555 B.n254 B.n132 71.676
R1556 B.n258 B.n133 71.676
R1557 B.n262 B.n134 71.676
R1558 B.n266 B.n135 71.676
R1559 B.n270 B.n136 71.676
R1560 B.n274 B.n137 71.676
R1561 B.n278 B.n138 71.676
R1562 B.n282 B.n139 71.676
R1563 B.n286 B.n140 71.676
R1564 B.n141 B.n140 71.676
R1565 B.n285 B.n139 71.676
R1566 B.n281 B.n138 71.676
R1567 B.n277 B.n137 71.676
R1568 B.n273 B.n136 71.676
R1569 B.n269 B.n135 71.676
R1570 B.n265 B.n134 71.676
R1571 B.n261 B.n133 71.676
R1572 B.n257 B.n132 71.676
R1573 B.n253 B.n131 71.676
R1574 B.n249 B.n130 71.676
R1575 B.n245 B.n129 71.676
R1576 B.n241 B.n128 71.676
R1577 B.n237 B.n127 71.676
R1578 B.n233 B.n126 71.676
R1579 B.n229 B.n125 71.676
R1580 B.n224 B.n124 71.676
R1581 B.n220 B.n123 71.676
R1582 B.n216 B.n122 71.676
R1583 B.n212 B.n121 71.676
R1584 B.n208 B.n120 71.676
R1585 B.n204 B.n119 71.676
R1586 B.n200 B.n118 71.676
R1587 B.n196 B.n117 71.676
R1588 B.n192 B.n116 71.676
R1589 B.n188 B.n115 71.676
R1590 B.n184 B.n114 71.676
R1591 B.n180 B.n113 71.676
R1592 B.n176 B.n112 71.676
R1593 B.n172 B.n111 71.676
R1594 B.n168 B.n110 71.676
R1595 B.n164 B.n109 71.676
R1596 B.n160 B.n108 71.676
R1597 B.n156 B.n107 71.676
R1598 B.n152 B.n106 71.676
R1599 B.n148 B.n105 71.676
R1600 B.n440 B.n397 71.676
R1601 B.n444 B.n443 71.676
R1602 B.n449 B.n448 71.676
R1603 B.n452 B.n451 71.676
R1604 B.n457 B.n456 71.676
R1605 B.n460 B.n459 71.676
R1606 B.n465 B.n464 71.676
R1607 B.n468 B.n467 71.676
R1608 B.n473 B.n472 71.676
R1609 B.n476 B.n475 71.676
R1610 B.n481 B.n480 71.676
R1611 B.n484 B.n483 71.676
R1612 B.n489 B.n488 71.676
R1613 B.n492 B.n491 71.676
R1614 B.n497 B.n496 71.676
R1615 B.n500 B.n499 71.676
R1616 B.n506 B.n505 71.676
R1617 B.n509 B.n508 71.676
R1618 B.n514 B.n513 71.676
R1619 B.n517 B.n516 71.676
R1620 B.n523 B.n522 71.676
R1621 B.n526 B.n525 71.676
R1622 B.n531 B.n530 71.676
R1623 B.n534 B.n533 71.676
R1624 B.n539 B.n538 71.676
R1625 B.n542 B.n541 71.676
R1626 B.n547 B.n546 71.676
R1627 B.n550 B.n549 71.676
R1628 B.n555 B.n554 71.676
R1629 B.n558 B.n557 71.676
R1630 B.n563 B.n562 71.676
R1631 B.n566 B.n565 71.676
R1632 B.n571 B.n570 71.676
R1633 B.n574 B.n573 71.676
R1634 B.n579 B.n578 71.676
R1635 B.n582 B.n581 71.676
R1636 B.n441 B.n440 71.676
R1637 B.n443 B.n437 71.676
R1638 B.n450 B.n449 71.676
R1639 B.n451 B.n435 71.676
R1640 B.n458 B.n457 71.676
R1641 B.n459 B.n433 71.676
R1642 B.n466 B.n465 71.676
R1643 B.n467 B.n431 71.676
R1644 B.n474 B.n473 71.676
R1645 B.n475 B.n429 71.676
R1646 B.n482 B.n481 71.676
R1647 B.n483 B.n427 71.676
R1648 B.n490 B.n489 71.676
R1649 B.n491 B.n425 71.676
R1650 B.n498 B.n497 71.676
R1651 B.n499 B.n421 71.676
R1652 B.n507 B.n506 71.676
R1653 B.n508 B.n419 71.676
R1654 B.n515 B.n514 71.676
R1655 B.n516 B.n415 71.676
R1656 B.n524 B.n523 71.676
R1657 B.n525 B.n413 71.676
R1658 B.n532 B.n531 71.676
R1659 B.n533 B.n411 71.676
R1660 B.n540 B.n539 71.676
R1661 B.n541 B.n409 71.676
R1662 B.n548 B.n547 71.676
R1663 B.n549 B.n407 71.676
R1664 B.n556 B.n555 71.676
R1665 B.n557 B.n405 71.676
R1666 B.n564 B.n563 71.676
R1667 B.n565 B.n403 71.676
R1668 B.n572 B.n571 71.676
R1669 B.n573 B.n401 71.676
R1670 B.n580 B.n579 71.676
R1671 B.n581 B.n399 71.676
R1672 B.n946 B.n945 71.676
R1673 B.n946 B.n2 71.676
R1674 B.n146 B.n145 59.5399
R1675 B.n227 B.n143 59.5399
R1676 B.n520 B.n417 59.5399
R1677 B.n502 B.n423 59.5399
R1678 B.n587 B.n394 53.7554
R1679 B.n593 B.n394 53.7554
R1680 B.n593 B.n390 53.7554
R1681 B.n599 B.n390 53.7554
R1682 B.n599 B.n386 53.7554
R1683 B.n605 B.n386 53.7554
R1684 B.n605 B.n382 53.7554
R1685 B.n612 B.n382 53.7554
R1686 B.n612 B.n611 53.7554
R1687 B.n618 B.n375 53.7554
R1688 B.n624 B.n375 53.7554
R1689 B.n624 B.n371 53.7554
R1690 B.n630 B.n371 53.7554
R1691 B.n630 B.n367 53.7554
R1692 B.n636 B.n367 53.7554
R1693 B.n636 B.n363 53.7554
R1694 B.n642 B.n363 53.7554
R1695 B.n642 B.n359 53.7554
R1696 B.n648 B.n359 53.7554
R1697 B.n648 B.n355 53.7554
R1698 B.n654 B.n355 53.7554
R1699 B.n654 B.n351 53.7554
R1700 B.n660 B.n351 53.7554
R1701 B.n666 B.n347 53.7554
R1702 B.n666 B.n343 53.7554
R1703 B.n672 B.n343 53.7554
R1704 B.n672 B.n339 53.7554
R1705 B.n678 B.n339 53.7554
R1706 B.n678 B.n335 53.7554
R1707 B.n684 B.n335 53.7554
R1708 B.n684 B.n331 53.7554
R1709 B.n690 B.n331 53.7554
R1710 B.n690 B.n327 53.7554
R1711 B.n696 B.n327 53.7554
R1712 B.n702 B.n323 53.7554
R1713 B.n702 B.n319 53.7554
R1714 B.n708 B.n319 53.7554
R1715 B.n708 B.n315 53.7554
R1716 B.n714 B.n315 53.7554
R1717 B.n714 B.n311 53.7554
R1718 B.n720 B.n311 53.7554
R1719 B.n720 B.n307 53.7554
R1720 B.n726 B.n307 53.7554
R1721 B.n726 B.n303 53.7554
R1722 B.n732 B.n303 53.7554
R1723 B.n738 B.n299 53.7554
R1724 B.n738 B.n295 53.7554
R1725 B.n745 B.n295 53.7554
R1726 B.n745 B.n291 53.7554
R1727 B.n751 B.n291 53.7554
R1728 B.n751 B.n4 53.7554
R1729 B.n944 B.n4 53.7554
R1730 B.n944 B.n943 53.7554
R1731 B.n943 B.n942 53.7554
R1732 B.n942 B.n8 53.7554
R1733 B.n12 B.n8 53.7554
R1734 B.n935 B.n12 53.7554
R1735 B.n935 B.n934 53.7554
R1736 B.n934 B.n933 53.7554
R1737 B.n933 B.n16 53.7554
R1738 B.n927 B.n926 53.7554
R1739 B.n926 B.n925 53.7554
R1740 B.n925 B.n23 53.7554
R1741 B.n919 B.n23 53.7554
R1742 B.n919 B.n918 53.7554
R1743 B.n918 B.n917 53.7554
R1744 B.n917 B.n30 53.7554
R1745 B.n911 B.n30 53.7554
R1746 B.n911 B.n910 53.7554
R1747 B.n910 B.n909 53.7554
R1748 B.n909 B.n37 53.7554
R1749 B.n903 B.n902 53.7554
R1750 B.n902 B.n901 53.7554
R1751 B.n901 B.n44 53.7554
R1752 B.n895 B.n44 53.7554
R1753 B.n895 B.n894 53.7554
R1754 B.n894 B.n893 53.7554
R1755 B.n893 B.n51 53.7554
R1756 B.n887 B.n51 53.7554
R1757 B.n887 B.n886 53.7554
R1758 B.n886 B.n885 53.7554
R1759 B.n885 B.n58 53.7554
R1760 B.n879 B.n878 53.7554
R1761 B.n878 B.n877 53.7554
R1762 B.n877 B.n65 53.7554
R1763 B.n871 B.n65 53.7554
R1764 B.n871 B.n870 53.7554
R1765 B.n870 B.n869 53.7554
R1766 B.n869 B.n72 53.7554
R1767 B.n863 B.n72 53.7554
R1768 B.n863 B.n862 53.7554
R1769 B.n862 B.n861 53.7554
R1770 B.n861 B.n79 53.7554
R1771 B.n855 B.n79 53.7554
R1772 B.n855 B.n854 53.7554
R1773 B.n854 B.n853 53.7554
R1774 B.n847 B.n89 53.7554
R1775 B.n847 B.n846 53.7554
R1776 B.n846 B.n845 53.7554
R1777 B.n845 B.n93 53.7554
R1778 B.n839 B.n93 53.7554
R1779 B.n839 B.n838 53.7554
R1780 B.n838 B.n837 53.7554
R1781 B.n837 B.n100 53.7554
R1782 B.n831 B.n100 53.7554
R1783 B.n732 B.t3 45.8503
R1784 B.n927 B.t1 45.8503
R1785 B.n696 B.t0 41.1072
R1786 B.n903 B.t5 41.1072
R1787 B.n660 B.t4 36.3641
R1788 B.n879 B.t2 36.3641
R1789 B.n618 B.t11 33.2021
R1790 B.n853 B.t7 33.2021
R1791 B.n589 B.n396 32.3127
R1792 B.n585 B.n584 32.3127
R1793 B.n828 B.n827 32.3127
R1794 B.n833 B.n102 32.3127
R1795 B.n611 B.t11 20.5539
R1796 B.n89 B.t7 20.5539
R1797 B B.n947 18.0485
R1798 B.t4 B.n347 17.3918
R1799 B.t2 B.n58 17.3918
R1800 B.t0 B.n323 12.6487
R1801 B.t5 B.n37 12.6487
R1802 B.n590 B.n589 10.6151
R1803 B.n591 B.n590 10.6151
R1804 B.n591 B.n388 10.6151
R1805 B.n601 B.n388 10.6151
R1806 B.n602 B.n601 10.6151
R1807 B.n603 B.n602 10.6151
R1808 B.n603 B.n380 10.6151
R1809 B.n614 B.n380 10.6151
R1810 B.n615 B.n614 10.6151
R1811 B.n616 B.n615 10.6151
R1812 B.n616 B.n373 10.6151
R1813 B.n626 B.n373 10.6151
R1814 B.n627 B.n626 10.6151
R1815 B.n628 B.n627 10.6151
R1816 B.n628 B.n365 10.6151
R1817 B.n638 B.n365 10.6151
R1818 B.n639 B.n638 10.6151
R1819 B.n640 B.n639 10.6151
R1820 B.n640 B.n357 10.6151
R1821 B.n650 B.n357 10.6151
R1822 B.n651 B.n650 10.6151
R1823 B.n652 B.n651 10.6151
R1824 B.n652 B.n349 10.6151
R1825 B.n662 B.n349 10.6151
R1826 B.n663 B.n662 10.6151
R1827 B.n664 B.n663 10.6151
R1828 B.n664 B.n341 10.6151
R1829 B.n674 B.n341 10.6151
R1830 B.n675 B.n674 10.6151
R1831 B.n676 B.n675 10.6151
R1832 B.n676 B.n333 10.6151
R1833 B.n686 B.n333 10.6151
R1834 B.n687 B.n686 10.6151
R1835 B.n688 B.n687 10.6151
R1836 B.n688 B.n325 10.6151
R1837 B.n698 B.n325 10.6151
R1838 B.n699 B.n698 10.6151
R1839 B.n700 B.n699 10.6151
R1840 B.n700 B.n317 10.6151
R1841 B.n710 B.n317 10.6151
R1842 B.n711 B.n710 10.6151
R1843 B.n712 B.n711 10.6151
R1844 B.n712 B.n309 10.6151
R1845 B.n722 B.n309 10.6151
R1846 B.n723 B.n722 10.6151
R1847 B.n724 B.n723 10.6151
R1848 B.n724 B.n301 10.6151
R1849 B.n734 B.n301 10.6151
R1850 B.n735 B.n734 10.6151
R1851 B.n736 B.n735 10.6151
R1852 B.n736 B.n293 10.6151
R1853 B.n747 B.n293 10.6151
R1854 B.n748 B.n747 10.6151
R1855 B.n749 B.n748 10.6151
R1856 B.n749 B.n0 10.6151
R1857 B.n439 B.n396 10.6151
R1858 B.n439 B.n438 10.6151
R1859 B.n445 B.n438 10.6151
R1860 B.n446 B.n445 10.6151
R1861 B.n447 B.n446 10.6151
R1862 B.n447 B.n436 10.6151
R1863 B.n453 B.n436 10.6151
R1864 B.n454 B.n453 10.6151
R1865 B.n455 B.n454 10.6151
R1866 B.n455 B.n434 10.6151
R1867 B.n461 B.n434 10.6151
R1868 B.n462 B.n461 10.6151
R1869 B.n463 B.n462 10.6151
R1870 B.n463 B.n432 10.6151
R1871 B.n469 B.n432 10.6151
R1872 B.n470 B.n469 10.6151
R1873 B.n471 B.n470 10.6151
R1874 B.n471 B.n430 10.6151
R1875 B.n477 B.n430 10.6151
R1876 B.n478 B.n477 10.6151
R1877 B.n479 B.n478 10.6151
R1878 B.n479 B.n428 10.6151
R1879 B.n485 B.n428 10.6151
R1880 B.n486 B.n485 10.6151
R1881 B.n487 B.n486 10.6151
R1882 B.n487 B.n426 10.6151
R1883 B.n493 B.n426 10.6151
R1884 B.n494 B.n493 10.6151
R1885 B.n495 B.n494 10.6151
R1886 B.n495 B.n424 10.6151
R1887 B.n501 B.n424 10.6151
R1888 B.n504 B.n503 10.6151
R1889 B.n504 B.n420 10.6151
R1890 B.n510 B.n420 10.6151
R1891 B.n511 B.n510 10.6151
R1892 B.n512 B.n511 10.6151
R1893 B.n512 B.n418 10.6151
R1894 B.n518 B.n418 10.6151
R1895 B.n519 B.n518 10.6151
R1896 B.n521 B.n414 10.6151
R1897 B.n527 B.n414 10.6151
R1898 B.n528 B.n527 10.6151
R1899 B.n529 B.n528 10.6151
R1900 B.n529 B.n412 10.6151
R1901 B.n535 B.n412 10.6151
R1902 B.n536 B.n535 10.6151
R1903 B.n537 B.n536 10.6151
R1904 B.n537 B.n410 10.6151
R1905 B.n543 B.n410 10.6151
R1906 B.n544 B.n543 10.6151
R1907 B.n545 B.n544 10.6151
R1908 B.n545 B.n408 10.6151
R1909 B.n551 B.n408 10.6151
R1910 B.n552 B.n551 10.6151
R1911 B.n553 B.n552 10.6151
R1912 B.n553 B.n406 10.6151
R1913 B.n559 B.n406 10.6151
R1914 B.n560 B.n559 10.6151
R1915 B.n561 B.n560 10.6151
R1916 B.n561 B.n404 10.6151
R1917 B.n567 B.n404 10.6151
R1918 B.n568 B.n567 10.6151
R1919 B.n569 B.n568 10.6151
R1920 B.n569 B.n402 10.6151
R1921 B.n575 B.n402 10.6151
R1922 B.n576 B.n575 10.6151
R1923 B.n577 B.n576 10.6151
R1924 B.n577 B.n400 10.6151
R1925 B.n583 B.n400 10.6151
R1926 B.n584 B.n583 10.6151
R1927 B.n585 B.n392 10.6151
R1928 B.n595 B.n392 10.6151
R1929 B.n596 B.n595 10.6151
R1930 B.n597 B.n596 10.6151
R1931 B.n597 B.n384 10.6151
R1932 B.n607 B.n384 10.6151
R1933 B.n608 B.n607 10.6151
R1934 B.n609 B.n608 10.6151
R1935 B.n609 B.n377 10.6151
R1936 B.n620 B.n377 10.6151
R1937 B.n621 B.n620 10.6151
R1938 B.n622 B.n621 10.6151
R1939 B.n622 B.n369 10.6151
R1940 B.n632 B.n369 10.6151
R1941 B.n633 B.n632 10.6151
R1942 B.n634 B.n633 10.6151
R1943 B.n634 B.n361 10.6151
R1944 B.n644 B.n361 10.6151
R1945 B.n645 B.n644 10.6151
R1946 B.n646 B.n645 10.6151
R1947 B.n646 B.n353 10.6151
R1948 B.n656 B.n353 10.6151
R1949 B.n657 B.n656 10.6151
R1950 B.n658 B.n657 10.6151
R1951 B.n658 B.n345 10.6151
R1952 B.n668 B.n345 10.6151
R1953 B.n669 B.n668 10.6151
R1954 B.n670 B.n669 10.6151
R1955 B.n670 B.n337 10.6151
R1956 B.n680 B.n337 10.6151
R1957 B.n681 B.n680 10.6151
R1958 B.n682 B.n681 10.6151
R1959 B.n682 B.n329 10.6151
R1960 B.n692 B.n329 10.6151
R1961 B.n693 B.n692 10.6151
R1962 B.n694 B.n693 10.6151
R1963 B.n694 B.n321 10.6151
R1964 B.n704 B.n321 10.6151
R1965 B.n705 B.n704 10.6151
R1966 B.n706 B.n705 10.6151
R1967 B.n706 B.n313 10.6151
R1968 B.n716 B.n313 10.6151
R1969 B.n717 B.n716 10.6151
R1970 B.n718 B.n717 10.6151
R1971 B.n718 B.n305 10.6151
R1972 B.n728 B.n305 10.6151
R1973 B.n729 B.n728 10.6151
R1974 B.n730 B.n729 10.6151
R1975 B.n730 B.n297 10.6151
R1976 B.n740 B.n297 10.6151
R1977 B.n741 B.n740 10.6151
R1978 B.n743 B.n741 10.6151
R1979 B.n743 B.n742 10.6151
R1980 B.n742 B.n289 10.6151
R1981 B.n754 B.n289 10.6151
R1982 B.n755 B.n754 10.6151
R1983 B.n756 B.n755 10.6151
R1984 B.n757 B.n756 10.6151
R1985 B.n758 B.n757 10.6151
R1986 B.n761 B.n758 10.6151
R1987 B.n762 B.n761 10.6151
R1988 B.n763 B.n762 10.6151
R1989 B.n764 B.n763 10.6151
R1990 B.n766 B.n764 10.6151
R1991 B.n767 B.n766 10.6151
R1992 B.n768 B.n767 10.6151
R1993 B.n769 B.n768 10.6151
R1994 B.n771 B.n769 10.6151
R1995 B.n772 B.n771 10.6151
R1996 B.n773 B.n772 10.6151
R1997 B.n774 B.n773 10.6151
R1998 B.n776 B.n774 10.6151
R1999 B.n777 B.n776 10.6151
R2000 B.n778 B.n777 10.6151
R2001 B.n779 B.n778 10.6151
R2002 B.n781 B.n779 10.6151
R2003 B.n782 B.n781 10.6151
R2004 B.n783 B.n782 10.6151
R2005 B.n784 B.n783 10.6151
R2006 B.n786 B.n784 10.6151
R2007 B.n787 B.n786 10.6151
R2008 B.n788 B.n787 10.6151
R2009 B.n789 B.n788 10.6151
R2010 B.n791 B.n789 10.6151
R2011 B.n792 B.n791 10.6151
R2012 B.n793 B.n792 10.6151
R2013 B.n794 B.n793 10.6151
R2014 B.n796 B.n794 10.6151
R2015 B.n797 B.n796 10.6151
R2016 B.n798 B.n797 10.6151
R2017 B.n799 B.n798 10.6151
R2018 B.n801 B.n799 10.6151
R2019 B.n802 B.n801 10.6151
R2020 B.n803 B.n802 10.6151
R2021 B.n804 B.n803 10.6151
R2022 B.n806 B.n804 10.6151
R2023 B.n807 B.n806 10.6151
R2024 B.n808 B.n807 10.6151
R2025 B.n809 B.n808 10.6151
R2026 B.n811 B.n809 10.6151
R2027 B.n812 B.n811 10.6151
R2028 B.n813 B.n812 10.6151
R2029 B.n814 B.n813 10.6151
R2030 B.n816 B.n814 10.6151
R2031 B.n817 B.n816 10.6151
R2032 B.n818 B.n817 10.6151
R2033 B.n819 B.n818 10.6151
R2034 B.n821 B.n819 10.6151
R2035 B.n822 B.n821 10.6151
R2036 B.n823 B.n822 10.6151
R2037 B.n824 B.n823 10.6151
R2038 B.n826 B.n824 10.6151
R2039 B.n827 B.n826 10.6151
R2040 B.n939 B.n1 10.6151
R2041 B.n939 B.n938 10.6151
R2042 B.n938 B.n937 10.6151
R2043 B.n937 B.n10 10.6151
R2044 B.n931 B.n10 10.6151
R2045 B.n931 B.n930 10.6151
R2046 B.n930 B.n929 10.6151
R2047 B.n929 B.n18 10.6151
R2048 B.n923 B.n18 10.6151
R2049 B.n923 B.n922 10.6151
R2050 B.n922 B.n921 10.6151
R2051 B.n921 B.n25 10.6151
R2052 B.n915 B.n25 10.6151
R2053 B.n915 B.n914 10.6151
R2054 B.n914 B.n913 10.6151
R2055 B.n913 B.n32 10.6151
R2056 B.n907 B.n32 10.6151
R2057 B.n907 B.n906 10.6151
R2058 B.n906 B.n905 10.6151
R2059 B.n905 B.n39 10.6151
R2060 B.n899 B.n39 10.6151
R2061 B.n899 B.n898 10.6151
R2062 B.n898 B.n897 10.6151
R2063 B.n897 B.n46 10.6151
R2064 B.n891 B.n46 10.6151
R2065 B.n891 B.n890 10.6151
R2066 B.n890 B.n889 10.6151
R2067 B.n889 B.n53 10.6151
R2068 B.n883 B.n53 10.6151
R2069 B.n883 B.n882 10.6151
R2070 B.n882 B.n881 10.6151
R2071 B.n881 B.n60 10.6151
R2072 B.n875 B.n60 10.6151
R2073 B.n875 B.n874 10.6151
R2074 B.n874 B.n873 10.6151
R2075 B.n873 B.n67 10.6151
R2076 B.n867 B.n67 10.6151
R2077 B.n867 B.n866 10.6151
R2078 B.n866 B.n865 10.6151
R2079 B.n865 B.n74 10.6151
R2080 B.n859 B.n74 10.6151
R2081 B.n859 B.n858 10.6151
R2082 B.n858 B.n857 10.6151
R2083 B.n857 B.n81 10.6151
R2084 B.n851 B.n81 10.6151
R2085 B.n851 B.n850 10.6151
R2086 B.n850 B.n849 10.6151
R2087 B.n849 B.n87 10.6151
R2088 B.n843 B.n87 10.6151
R2089 B.n843 B.n842 10.6151
R2090 B.n842 B.n841 10.6151
R2091 B.n841 B.n95 10.6151
R2092 B.n835 B.n95 10.6151
R2093 B.n835 B.n834 10.6151
R2094 B.n834 B.n833 10.6151
R2095 B.n147 B.n102 10.6151
R2096 B.n150 B.n147 10.6151
R2097 B.n151 B.n150 10.6151
R2098 B.n154 B.n151 10.6151
R2099 B.n155 B.n154 10.6151
R2100 B.n158 B.n155 10.6151
R2101 B.n159 B.n158 10.6151
R2102 B.n162 B.n159 10.6151
R2103 B.n163 B.n162 10.6151
R2104 B.n166 B.n163 10.6151
R2105 B.n167 B.n166 10.6151
R2106 B.n170 B.n167 10.6151
R2107 B.n171 B.n170 10.6151
R2108 B.n174 B.n171 10.6151
R2109 B.n175 B.n174 10.6151
R2110 B.n178 B.n175 10.6151
R2111 B.n179 B.n178 10.6151
R2112 B.n182 B.n179 10.6151
R2113 B.n183 B.n182 10.6151
R2114 B.n186 B.n183 10.6151
R2115 B.n187 B.n186 10.6151
R2116 B.n190 B.n187 10.6151
R2117 B.n191 B.n190 10.6151
R2118 B.n194 B.n191 10.6151
R2119 B.n195 B.n194 10.6151
R2120 B.n198 B.n195 10.6151
R2121 B.n199 B.n198 10.6151
R2122 B.n202 B.n199 10.6151
R2123 B.n203 B.n202 10.6151
R2124 B.n206 B.n203 10.6151
R2125 B.n207 B.n206 10.6151
R2126 B.n211 B.n210 10.6151
R2127 B.n214 B.n211 10.6151
R2128 B.n215 B.n214 10.6151
R2129 B.n218 B.n215 10.6151
R2130 B.n219 B.n218 10.6151
R2131 B.n222 B.n219 10.6151
R2132 B.n223 B.n222 10.6151
R2133 B.n226 B.n223 10.6151
R2134 B.n231 B.n228 10.6151
R2135 B.n232 B.n231 10.6151
R2136 B.n235 B.n232 10.6151
R2137 B.n236 B.n235 10.6151
R2138 B.n239 B.n236 10.6151
R2139 B.n240 B.n239 10.6151
R2140 B.n243 B.n240 10.6151
R2141 B.n244 B.n243 10.6151
R2142 B.n247 B.n244 10.6151
R2143 B.n248 B.n247 10.6151
R2144 B.n251 B.n248 10.6151
R2145 B.n252 B.n251 10.6151
R2146 B.n255 B.n252 10.6151
R2147 B.n256 B.n255 10.6151
R2148 B.n259 B.n256 10.6151
R2149 B.n260 B.n259 10.6151
R2150 B.n263 B.n260 10.6151
R2151 B.n264 B.n263 10.6151
R2152 B.n267 B.n264 10.6151
R2153 B.n268 B.n267 10.6151
R2154 B.n271 B.n268 10.6151
R2155 B.n272 B.n271 10.6151
R2156 B.n275 B.n272 10.6151
R2157 B.n276 B.n275 10.6151
R2158 B.n279 B.n276 10.6151
R2159 B.n280 B.n279 10.6151
R2160 B.n283 B.n280 10.6151
R2161 B.n284 B.n283 10.6151
R2162 B.n287 B.n284 10.6151
R2163 B.n288 B.n287 10.6151
R2164 B.n828 B.n288 10.6151
R2165 B.n947 B.n0 8.11757
R2166 B.n947 B.n1 8.11757
R2167 B.t3 B.n299 7.90564
R2168 B.t1 B.n16 7.90564
R2169 B.n503 B.n502 6.5566
R2170 B.n520 B.n519 6.5566
R2171 B.n210 B.n146 6.5566
R2172 B.n227 B.n226 6.5566
R2173 B.n502 B.n501 4.05904
R2174 B.n521 B.n520 4.05904
R2175 B.n207 B.n146 4.05904
R2176 B.n228 B.n227 4.05904
R2177 VN.n38 VN.n37 161.3
R2178 VN.n36 VN.n21 161.3
R2179 VN.n35 VN.n34 161.3
R2180 VN.n33 VN.n22 161.3
R2181 VN.n32 VN.n31 161.3
R2182 VN.n30 VN.n23 161.3
R2183 VN.n29 VN.n28 161.3
R2184 VN.n27 VN.n24 161.3
R2185 VN.n18 VN.n17 161.3
R2186 VN.n16 VN.n1 161.3
R2187 VN.n15 VN.n14 161.3
R2188 VN.n13 VN.n2 161.3
R2189 VN.n12 VN.n11 161.3
R2190 VN.n10 VN.n3 161.3
R2191 VN.n9 VN.n8 161.3
R2192 VN.n7 VN.n4 161.3
R2193 VN.n26 VN.t4 88.505
R2194 VN.n6 VN.t5 88.505
R2195 VN.n19 VN.n0 84.5354
R2196 VN.n39 VN.n20 84.5354
R2197 VN.n5 VN.t2 55.0862
R2198 VN.n0 VN.t1 55.0862
R2199 VN.n25 VN.t0 55.0862
R2200 VN.n20 VN.t3 55.0862
R2201 VN VN.n39 51.0093
R2202 VN.n6 VN.n5 50.3788
R2203 VN.n26 VN.n25 50.3788
R2204 VN.n11 VN.n2 45.7662
R2205 VN.n31 VN.n22 45.7662
R2206 VN.n11 VN.n10 35.055
R2207 VN.n31 VN.n30 35.055
R2208 VN.n5 VN.n4 24.3439
R2209 VN.n9 VN.n4 24.3439
R2210 VN.n10 VN.n9 24.3439
R2211 VN.n15 VN.n2 24.3439
R2212 VN.n16 VN.n15 24.3439
R2213 VN.n17 VN.n16 24.3439
R2214 VN.n30 VN.n29 24.3439
R2215 VN.n29 VN.n24 24.3439
R2216 VN.n25 VN.n24 24.3439
R2217 VN.n37 VN.n36 24.3439
R2218 VN.n36 VN.n35 24.3439
R2219 VN.n35 VN.n22 24.3439
R2220 VN.n17 VN.n0 5.35606
R2221 VN.n37 VN.n20 5.35606
R2222 VN.n27 VN.n26 2.42077
R2223 VN.n7 VN.n6 2.42077
R2224 VN.n39 VN.n38 0.355081
R2225 VN.n19 VN.n18 0.355081
R2226 VN VN.n19 0.26685
R2227 VN.n38 VN.n21 0.189894
R2228 VN.n34 VN.n21 0.189894
R2229 VN.n34 VN.n33 0.189894
R2230 VN.n33 VN.n32 0.189894
R2231 VN.n32 VN.n23 0.189894
R2232 VN.n28 VN.n23 0.189894
R2233 VN.n28 VN.n27 0.189894
R2234 VN.n8 VN.n7 0.189894
R2235 VN.n8 VN.n3 0.189894
R2236 VN.n12 VN.n3 0.189894
R2237 VN.n13 VN.n12 0.189894
R2238 VN.n14 VN.n13 0.189894
R2239 VN.n14 VN.n1 0.189894
R2240 VN.n18 VN.n1 0.189894
R2241 VDD2.n87 VDD2.n47 289.615
R2242 VDD2.n40 VDD2.n0 289.615
R2243 VDD2.n88 VDD2.n87 185
R2244 VDD2.n86 VDD2.n85 185
R2245 VDD2.n84 VDD2.n50 185
R2246 VDD2.n54 VDD2.n51 185
R2247 VDD2.n79 VDD2.n78 185
R2248 VDD2.n77 VDD2.n76 185
R2249 VDD2.n56 VDD2.n55 185
R2250 VDD2.n71 VDD2.n70 185
R2251 VDD2.n69 VDD2.n68 185
R2252 VDD2.n60 VDD2.n59 185
R2253 VDD2.n63 VDD2.n62 185
R2254 VDD2.n15 VDD2.n14 185
R2255 VDD2.n12 VDD2.n11 185
R2256 VDD2.n21 VDD2.n20 185
R2257 VDD2.n23 VDD2.n22 185
R2258 VDD2.n8 VDD2.n7 185
R2259 VDD2.n29 VDD2.n28 185
R2260 VDD2.n32 VDD2.n31 185
R2261 VDD2.n30 VDD2.n4 185
R2262 VDD2.n37 VDD2.n3 185
R2263 VDD2.n39 VDD2.n38 185
R2264 VDD2.n41 VDD2.n40 185
R2265 VDD2.t2 VDD2.n61 149.524
R2266 VDD2.t0 VDD2.n13 149.524
R2267 VDD2.n87 VDD2.n86 104.615
R2268 VDD2.n86 VDD2.n50 104.615
R2269 VDD2.n54 VDD2.n50 104.615
R2270 VDD2.n78 VDD2.n54 104.615
R2271 VDD2.n78 VDD2.n77 104.615
R2272 VDD2.n77 VDD2.n55 104.615
R2273 VDD2.n70 VDD2.n55 104.615
R2274 VDD2.n70 VDD2.n69 104.615
R2275 VDD2.n69 VDD2.n59 104.615
R2276 VDD2.n62 VDD2.n59 104.615
R2277 VDD2.n14 VDD2.n11 104.615
R2278 VDD2.n21 VDD2.n11 104.615
R2279 VDD2.n22 VDD2.n21 104.615
R2280 VDD2.n22 VDD2.n7 104.615
R2281 VDD2.n29 VDD2.n7 104.615
R2282 VDD2.n31 VDD2.n29 104.615
R2283 VDD2.n31 VDD2.n30 104.615
R2284 VDD2.n30 VDD2.n3 104.615
R2285 VDD2.n39 VDD2.n3 104.615
R2286 VDD2.n40 VDD2.n39 104.615
R2287 VDD2.n46 VDD2.n45 66.5987
R2288 VDD2 VDD2.n93 66.5959
R2289 VDD2.n46 VDD2.n44 53.7934
R2290 VDD2.n62 VDD2.t2 52.3082
R2291 VDD2.n14 VDD2.t0 52.3082
R2292 VDD2.n92 VDD2.n91 51.1914
R2293 VDD2.n92 VDD2.n46 42.6787
R2294 VDD2.n85 VDD2.n84 13.1884
R2295 VDD2.n38 VDD2.n37 13.1884
R2296 VDD2.n88 VDD2.n49 12.8005
R2297 VDD2.n83 VDD2.n51 12.8005
R2298 VDD2.n36 VDD2.n4 12.8005
R2299 VDD2.n41 VDD2.n2 12.8005
R2300 VDD2.n89 VDD2.n47 12.0247
R2301 VDD2.n80 VDD2.n79 12.0247
R2302 VDD2.n33 VDD2.n32 12.0247
R2303 VDD2.n42 VDD2.n0 12.0247
R2304 VDD2.n76 VDD2.n53 11.249
R2305 VDD2.n28 VDD2.n6 11.249
R2306 VDD2.n75 VDD2.n56 10.4732
R2307 VDD2.n27 VDD2.n8 10.4732
R2308 VDD2.n63 VDD2.n61 10.2747
R2309 VDD2.n15 VDD2.n13 10.2747
R2310 VDD2.n72 VDD2.n71 9.69747
R2311 VDD2.n24 VDD2.n23 9.69747
R2312 VDD2.n91 VDD2.n90 9.45567
R2313 VDD2.n44 VDD2.n43 9.45567
R2314 VDD2.n65 VDD2.n64 9.3005
R2315 VDD2.n67 VDD2.n66 9.3005
R2316 VDD2.n58 VDD2.n57 9.3005
R2317 VDD2.n73 VDD2.n72 9.3005
R2318 VDD2.n75 VDD2.n74 9.3005
R2319 VDD2.n53 VDD2.n52 9.3005
R2320 VDD2.n81 VDD2.n80 9.3005
R2321 VDD2.n83 VDD2.n82 9.3005
R2322 VDD2.n90 VDD2.n89 9.3005
R2323 VDD2.n49 VDD2.n48 9.3005
R2324 VDD2.n43 VDD2.n42 9.3005
R2325 VDD2.n2 VDD2.n1 9.3005
R2326 VDD2.n17 VDD2.n16 9.3005
R2327 VDD2.n19 VDD2.n18 9.3005
R2328 VDD2.n10 VDD2.n9 9.3005
R2329 VDD2.n25 VDD2.n24 9.3005
R2330 VDD2.n27 VDD2.n26 9.3005
R2331 VDD2.n6 VDD2.n5 9.3005
R2332 VDD2.n34 VDD2.n33 9.3005
R2333 VDD2.n36 VDD2.n35 9.3005
R2334 VDD2.n68 VDD2.n58 8.92171
R2335 VDD2.n20 VDD2.n10 8.92171
R2336 VDD2.n67 VDD2.n60 8.14595
R2337 VDD2.n19 VDD2.n12 8.14595
R2338 VDD2.n64 VDD2.n63 7.3702
R2339 VDD2.n16 VDD2.n15 7.3702
R2340 VDD2.n64 VDD2.n60 5.81868
R2341 VDD2.n16 VDD2.n12 5.81868
R2342 VDD2.n68 VDD2.n67 5.04292
R2343 VDD2.n20 VDD2.n19 5.04292
R2344 VDD2.n71 VDD2.n58 4.26717
R2345 VDD2.n23 VDD2.n10 4.26717
R2346 VDD2.n72 VDD2.n56 3.49141
R2347 VDD2.n24 VDD2.n8 3.49141
R2348 VDD2.n17 VDD2.n13 2.84303
R2349 VDD2.n65 VDD2.n61 2.84303
R2350 VDD2 VDD2.n92 2.71602
R2351 VDD2.n76 VDD2.n75 2.71565
R2352 VDD2.n28 VDD2.n27 2.71565
R2353 VDD2.n93 VDD2.t5 2.29217
R2354 VDD2.n93 VDD2.t1 2.29217
R2355 VDD2.n45 VDD2.t3 2.29217
R2356 VDD2.n45 VDD2.t4 2.29217
R2357 VDD2.n91 VDD2.n47 1.93989
R2358 VDD2.n79 VDD2.n53 1.93989
R2359 VDD2.n32 VDD2.n6 1.93989
R2360 VDD2.n44 VDD2.n0 1.93989
R2361 VDD2.n89 VDD2.n88 1.16414
R2362 VDD2.n80 VDD2.n51 1.16414
R2363 VDD2.n33 VDD2.n4 1.16414
R2364 VDD2.n42 VDD2.n41 1.16414
R2365 VDD2.n85 VDD2.n49 0.388379
R2366 VDD2.n84 VDD2.n83 0.388379
R2367 VDD2.n37 VDD2.n36 0.388379
R2368 VDD2.n38 VDD2.n2 0.388379
R2369 VDD2.n90 VDD2.n48 0.155672
R2370 VDD2.n82 VDD2.n48 0.155672
R2371 VDD2.n82 VDD2.n81 0.155672
R2372 VDD2.n81 VDD2.n52 0.155672
R2373 VDD2.n74 VDD2.n52 0.155672
R2374 VDD2.n74 VDD2.n73 0.155672
R2375 VDD2.n73 VDD2.n57 0.155672
R2376 VDD2.n66 VDD2.n57 0.155672
R2377 VDD2.n66 VDD2.n65 0.155672
R2378 VDD2.n18 VDD2.n17 0.155672
R2379 VDD2.n18 VDD2.n9 0.155672
R2380 VDD2.n25 VDD2.n9 0.155672
R2381 VDD2.n26 VDD2.n25 0.155672
R2382 VDD2.n26 VDD2.n5 0.155672
R2383 VDD2.n34 VDD2.n5 0.155672
R2384 VDD2.n35 VDD2.n34 0.155672
R2385 VDD2.n35 VDD2.n1 0.155672
R2386 VDD2.n43 VDD2.n1 0.155672
C0 VTAIL VDD1 7.08182f
C1 VP VN 7.457211f
C2 VDD2 VN 5.25678f
C3 VDD2 VP 0.557435f
C4 VN VTAIL 5.86094f
C5 VN VDD1 0.151914f
C6 VP VTAIL 5.875451f
C7 VDD2 VTAIL 7.14204f
C8 VP VDD1 5.66f
C9 VDD2 VDD1 1.86647f
C10 VDD2 B 6.285424f
C11 VDD1 B 6.47915f
C12 VTAIL B 7.190857f
C13 VN B 16.13677f
C14 VP B 14.86338f
C15 VDD2.n0 B 0.029189f
C16 VDD2.n1 B 0.021596f
C17 VDD2.n2 B 0.011605f
C18 VDD2.n3 B 0.027429f
C19 VDD2.n4 B 0.012287f
C20 VDD2.n5 B 0.021596f
C21 VDD2.n6 B 0.011605f
C22 VDD2.n7 B 0.027429f
C23 VDD2.n8 B 0.012287f
C24 VDD2.n9 B 0.021596f
C25 VDD2.n10 B 0.011605f
C26 VDD2.n11 B 0.027429f
C27 VDD2.n12 B 0.012287f
C28 VDD2.n13 B 0.12786f
C29 VDD2.t0 B 0.045943f
C30 VDD2.n14 B 0.020572f
C31 VDD2.n15 B 0.01939f
C32 VDD2.n16 B 0.011605f
C33 VDD2.n17 B 0.766713f
C34 VDD2.n18 B 0.021596f
C35 VDD2.n19 B 0.011605f
C36 VDD2.n20 B 0.012287f
C37 VDD2.n21 B 0.027429f
C38 VDD2.n22 B 0.027429f
C39 VDD2.n23 B 0.012287f
C40 VDD2.n24 B 0.011605f
C41 VDD2.n25 B 0.021596f
C42 VDD2.n26 B 0.021596f
C43 VDD2.n27 B 0.011605f
C44 VDD2.n28 B 0.012287f
C45 VDD2.n29 B 0.027429f
C46 VDD2.n30 B 0.027429f
C47 VDD2.n31 B 0.027429f
C48 VDD2.n32 B 0.012287f
C49 VDD2.n33 B 0.011605f
C50 VDD2.n34 B 0.021596f
C51 VDD2.n35 B 0.021596f
C52 VDD2.n36 B 0.011605f
C53 VDD2.n37 B 0.011946f
C54 VDD2.n38 B 0.011946f
C55 VDD2.n39 B 0.027429f
C56 VDD2.n40 B 0.057319f
C57 VDD2.n41 B 0.012287f
C58 VDD2.n42 B 0.011605f
C59 VDD2.n43 B 0.053458f
C60 VDD2.n44 B 0.057728f
C61 VDD2.t3 B 0.147449f
C62 VDD2.t4 B 0.147449f
C63 VDD2.n45 B 1.2916f
C64 VDD2.n46 B 2.57104f
C65 VDD2.n47 B 0.029189f
C66 VDD2.n48 B 0.021596f
C67 VDD2.n49 B 0.011605f
C68 VDD2.n50 B 0.027429f
C69 VDD2.n51 B 0.012287f
C70 VDD2.n52 B 0.021596f
C71 VDD2.n53 B 0.011605f
C72 VDD2.n54 B 0.027429f
C73 VDD2.n55 B 0.027429f
C74 VDD2.n56 B 0.012287f
C75 VDD2.n57 B 0.021596f
C76 VDD2.n58 B 0.011605f
C77 VDD2.n59 B 0.027429f
C78 VDD2.n60 B 0.012287f
C79 VDD2.n61 B 0.12786f
C80 VDD2.t2 B 0.045943f
C81 VDD2.n62 B 0.020572f
C82 VDD2.n63 B 0.01939f
C83 VDD2.n64 B 0.011605f
C84 VDD2.n65 B 0.766713f
C85 VDD2.n66 B 0.021596f
C86 VDD2.n67 B 0.011605f
C87 VDD2.n68 B 0.012287f
C88 VDD2.n69 B 0.027429f
C89 VDD2.n70 B 0.027429f
C90 VDD2.n71 B 0.012287f
C91 VDD2.n72 B 0.011605f
C92 VDD2.n73 B 0.021596f
C93 VDD2.n74 B 0.021596f
C94 VDD2.n75 B 0.011605f
C95 VDD2.n76 B 0.012287f
C96 VDD2.n77 B 0.027429f
C97 VDD2.n78 B 0.027429f
C98 VDD2.n79 B 0.012287f
C99 VDD2.n80 B 0.011605f
C100 VDD2.n81 B 0.021596f
C101 VDD2.n82 B 0.021596f
C102 VDD2.n83 B 0.011605f
C103 VDD2.n84 B 0.011946f
C104 VDD2.n85 B 0.011946f
C105 VDD2.n86 B 0.027429f
C106 VDD2.n87 B 0.057319f
C107 VDD2.n88 B 0.012287f
C108 VDD2.n89 B 0.011605f
C109 VDD2.n90 B 0.053458f
C110 VDD2.n91 B 0.046851f
C111 VDD2.n92 B 2.269f
C112 VDD2.t5 B 0.147449f
C113 VDD2.t1 B 0.147449f
C114 VDD2.n93 B 1.29157f
C115 VN.t1 B 1.72404f
C116 VN.n0 B 0.69222f
C117 VN.n1 B 0.019592f
C118 VN.n2 B 0.037716f
C119 VN.n3 B 0.019592f
C120 VN.n4 B 0.036698f
C121 VN.t2 B 1.72404f
C122 VN.n5 B 0.696995f
C123 VN.t5 B 2.0161f
C124 VN.n6 B 0.659171f
C125 VN.n7 B 0.250557f
C126 VN.n8 B 0.019592f
C127 VN.n9 B 0.036698f
C128 VN.n10 B 0.039799f
C129 VN.n11 B 0.016635f
C130 VN.n12 B 0.019592f
C131 VN.n13 B 0.019592f
C132 VN.n14 B 0.019592f
C133 VN.n15 B 0.036698f
C134 VN.n16 B 0.036698f
C135 VN.n17 B 0.022565f
C136 VN.n18 B 0.031627f
C137 VN.n19 B 0.058535f
C138 VN.t3 B 1.72404f
C139 VN.n20 B 0.69222f
C140 VN.n21 B 0.019592f
C141 VN.n22 B 0.037716f
C142 VN.n23 B 0.019592f
C143 VN.n24 B 0.036698f
C144 VN.t4 B 2.0161f
C145 VN.t0 B 1.72404f
C146 VN.n25 B 0.696995f
C147 VN.n26 B 0.659171f
C148 VN.n27 B 0.250557f
C149 VN.n28 B 0.019592f
C150 VN.n29 B 0.036698f
C151 VN.n30 B 0.039799f
C152 VN.n31 B 0.016635f
C153 VN.n32 B 0.019592f
C154 VN.n33 B 0.019592f
C155 VN.n34 B 0.019592f
C156 VN.n35 B 0.036698f
C157 VN.n36 B 0.036698f
C158 VN.n37 B 0.022565f
C159 VN.n38 B 0.031627f
C160 VN.n39 B 1.16148f
C161 VDD1.n0 B 0.029938f
C162 VDD1.n1 B 0.02215f
C163 VDD1.n2 B 0.011902f
C164 VDD1.n3 B 0.028133f
C165 VDD1.n4 B 0.012603f
C166 VDD1.n5 B 0.02215f
C167 VDD1.n6 B 0.011902f
C168 VDD1.n7 B 0.028133f
C169 VDD1.n8 B 0.028133f
C170 VDD1.n9 B 0.012603f
C171 VDD1.n10 B 0.02215f
C172 VDD1.n11 B 0.011902f
C173 VDD1.n12 B 0.028133f
C174 VDD1.n13 B 0.012603f
C175 VDD1.n14 B 0.131141f
C176 VDD1.t3 B 0.047122f
C177 VDD1.n15 B 0.0211f
C178 VDD1.n16 B 0.019888f
C179 VDD1.n17 B 0.011902f
C180 VDD1.n18 B 0.786387f
C181 VDD1.n19 B 0.02215f
C182 VDD1.n20 B 0.011902f
C183 VDD1.n21 B 0.012603f
C184 VDD1.n22 B 0.028133f
C185 VDD1.n23 B 0.028133f
C186 VDD1.n24 B 0.012603f
C187 VDD1.n25 B 0.011902f
C188 VDD1.n26 B 0.02215f
C189 VDD1.n27 B 0.02215f
C190 VDD1.n28 B 0.011902f
C191 VDD1.n29 B 0.012603f
C192 VDD1.n30 B 0.028133f
C193 VDD1.n31 B 0.028133f
C194 VDD1.n32 B 0.012603f
C195 VDD1.n33 B 0.011902f
C196 VDD1.n34 B 0.02215f
C197 VDD1.n35 B 0.02215f
C198 VDD1.n36 B 0.011902f
C199 VDD1.n37 B 0.012253f
C200 VDD1.n38 B 0.012253f
C201 VDD1.n39 B 0.028133f
C202 VDD1.n40 B 0.05879f
C203 VDD1.n41 B 0.012603f
C204 VDD1.n42 B 0.011902f
C205 VDD1.n43 B 0.05483f
C206 VDD1.n44 B 0.06007f
C207 VDD1.n45 B 0.029938f
C208 VDD1.n46 B 0.02215f
C209 VDD1.n47 B 0.011902f
C210 VDD1.n48 B 0.028133f
C211 VDD1.n49 B 0.012603f
C212 VDD1.n50 B 0.02215f
C213 VDD1.n51 B 0.011902f
C214 VDD1.n52 B 0.028133f
C215 VDD1.n53 B 0.012603f
C216 VDD1.n54 B 0.02215f
C217 VDD1.n55 B 0.011902f
C218 VDD1.n56 B 0.028133f
C219 VDD1.n57 B 0.012603f
C220 VDD1.n58 B 0.131141f
C221 VDD1.t1 B 0.047122f
C222 VDD1.n59 B 0.0211f
C223 VDD1.n60 B 0.019888f
C224 VDD1.n61 B 0.011902f
C225 VDD1.n62 B 0.786387f
C226 VDD1.n63 B 0.02215f
C227 VDD1.n64 B 0.011902f
C228 VDD1.n65 B 0.012603f
C229 VDD1.n66 B 0.028133f
C230 VDD1.n67 B 0.028133f
C231 VDD1.n68 B 0.012603f
C232 VDD1.n69 B 0.011902f
C233 VDD1.n70 B 0.02215f
C234 VDD1.n71 B 0.02215f
C235 VDD1.n72 B 0.011902f
C236 VDD1.n73 B 0.012603f
C237 VDD1.n74 B 0.028133f
C238 VDD1.n75 B 0.028133f
C239 VDD1.n76 B 0.028133f
C240 VDD1.n77 B 0.012603f
C241 VDD1.n78 B 0.011902f
C242 VDD1.n79 B 0.02215f
C243 VDD1.n80 B 0.02215f
C244 VDD1.n81 B 0.011902f
C245 VDD1.n82 B 0.012253f
C246 VDD1.n83 B 0.012253f
C247 VDD1.n84 B 0.028133f
C248 VDD1.n85 B 0.05879f
C249 VDD1.n86 B 0.012603f
C250 VDD1.n87 B 0.011902f
C251 VDD1.n88 B 0.05483f
C252 VDD1.n89 B 0.05921f
C253 VDD1.t2 B 0.151232f
C254 VDD1.t4 B 0.151232f
C255 VDD1.n90 B 1.32475f
C256 VDD1.n91 B 2.77184f
C257 VDD1.t0 B 0.151232f
C258 VDD1.t5 B 0.151232f
C259 VDD1.n92 B 1.31853f
C260 VDD1.n93 B 2.53336f
C261 VTAIL.t1 B 0.177986f
C262 VTAIL.t5 B 0.177986f
C263 VTAIL.n0 B 1.48276f
C264 VTAIL.n1 B 0.50927f
C265 VTAIL.n2 B 0.035235f
C266 VTAIL.n3 B 0.026069f
C267 VTAIL.n4 B 0.014008f
C268 VTAIL.n5 B 0.03311f
C269 VTAIL.n6 B 0.014832f
C270 VTAIL.n7 B 0.026069f
C271 VTAIL.n8 B 0.014008f
C272 VTAIL.n9 B 0.03311f
C273 VTAIL.n10 B 0.014832f
C274 VTAIL.n11 B 0.026069f
C275 VTAIL.n12 B 0.014008f
C276 VTAIL.n13 B 0.03311f
C277 VTAIL.n14 B 0.014832f
C278 VTAIL.n15 B 0.15434f
C279 VTAIL.t10 B 0.055458f
C280 VTAIL.n16 B 0.024833f
C281 VTAIL.n17 B 0.023406f
C282 VTAIL.n18 B 0.014008f
C283 VTAIL.n19 B 0.9255f
C284 VTAIL.n20 B 0.026069f
C285 VTAIL.n21 B 0.014008f
C286 VTAIL.n22 B 0.014832f
C287 VTAIL.n23 B 0.03311f
C288 VTAIL.n24 B 0.03311f
C289 VTAIL.n25 B 0.014832f
C290 VTAIL.n26 B 0.014008f
C291 VTAIL.n27 B 0.026069f
C292 VTAIL.n28 B 0.026069f
C293 VTAIL.n29 B 0.014008f
C294 VTAIL.n30 B 0.014832f
C295 VTAIL.n31 B 0.03311f
C296 VTAIL.n32 B 0.03311f
C297 VTAIL.n33 B 0.03311f
C298 VTAIL.n34 B 0.014832f
C299 VTAIL.n35 B 0.014008f
C300 VTAIL.n36 B 0.026069f
C301 VTAIL.n37 B 0.026069f
C302 VTAIL.n38 B 0.014008f
C303 VTAIL.n39 B 0.01442f
C304 VTAIL.n40 B 0.01442f
C305 VTAIL.n41 B 0.03311f
C306 VTAIL.n42 B 0.06919f
C307 VTAIL.n43 B 0.014832f
C308 VTAIL.n44 B 0.014008f
C309 VTAIL.n45 B 0.06453f
C310 VTAIL.n46 B 0.038586f
C311 VTAIL.n47 B 0.51057f
C312 VTAIL.t7 B 0.177986f
C313 VTAIL.t9 B 0.177986f
C314 VTAIL.n48 B 1.48276f
C315 VTAIL.n49 B 2.11431f
C316 VTAIL.t4 B 0.177986f
C317 VTAIL.t0 B 0.177986f
C318 VTAIL.n50 B 1.48277f
C319 VTAIL.n51 B 2.1143f
C320 VTAIL.n52 B 0.035235f
C321 VTAIL.n53 B 0.026069f
C322 VTAIL.n54 B 0.014008f
C323 VTAIL.n55 B 0.03311f
C324 VTAIL.n56 B 0.014832f
C325 VTAIL.n57 B 0.026069f
C326 VTAIL.n58 B 0.014008f
C327 VTAIL.n59 B 0.03311f
C328 VTAIL.n60 B 0.03311f
C329 VTAIL.n61 B 0.014832f
C330 VTAIL.n62 B 0.026069f
C331 VTAIL.n63 B 0.014008f
C332 VTAIL.n64 B 0.03311f
C333 VTAIL.n65 B 0.014832f
C334 VTAIL.n66 B 0.15434f
C335 VTAIL.t3 B 0.055458f
C336 VTAIL.n67 B 0.024833f
C337 VTAIL.n68 B 0.023406f
C338 VTAIL.n69 B 0.014008f
C339 VTAIL.n70 B 0.9255f
C340 VTAIL.n71 B 0.026069f
C341 VTAIL.n72 B 0.014008f
C342 VTAIL.n73 B 0.014832f
C343 VTAIL.n74 B 0.03311f
C344 VTAIL.n75 B 0.03311f
C345 VTAIL.n76 B 0.014832f
C346 VTAIL.n77 B 0.014008f
C347 VTAIL.n78 B 0.026069f
C348 VTAIL.n79 B 0.026069f
C349 VTAIL.n80 B 0.014008f
C350 VTAIL.n81 B 0.014832f
C351 VTAIL.n82 B 0.03311f
C352 VTAIL.n83 B 0.03311f
C353 VTAIL.n84 B 0.014832f
C354 VTAIL.n85 B 0.014008f
C355 VTAIL.n86 B 0.026069f
C356 VTAIL.n87 B 0.026069f
C357 VTAIL.n88 B 0.014008f
C358 VTAIL.n89 B 0.01442f
C359 VTAIL.n90 B 0.01442f
C360 VTAIL.n91 B 0.03311f
C361 VTAIL.n92 B 0.06919f
C362 VTAIL.n93 B 0.014832f
C363 VTAIL.n94 B 0.014008f
C364 VTAIL.n95 B 0.06453f
C365 VTAIL.n96 B 0.038586f
C366 VTAIL.n97 B 0.51057f
C367 VTAIL.t11 B 0.177986f
C368 VTAIL.t6 B 0.177986f
C369 VTAIL.n98 B 1.48277f
C370 VTAIL.n99 B 0.727585f
C371 VTAIL.n100 B 0.035235f
C372 VTAIL.n101 B 0.026069f
C373 VTAIL.n102 B 0.014008f
C374 VTAIL.n103 B 0.03311f
C375 VTAIL.n104 B 0.014832f
C376 VTAIL.n105 B 0.026069f
C377 VTAIL.n106 B 0.014008f
C378 VTAIL.n107 B 0.03311f
C379 VTAIL.n108 B 0.03311f
C380 VTAIL.n109 B 0.014832f
C381 VTAIL.n110 B 0.026069f
C382 VTAIL.n111 B 0.014008f
C383 VTAIL.n112 B 0.03311f
C384 VTAIL.n113 B 0.014832f
C385 VTAIL.n114 B 0.15434f
C386 VTAIL.t8 B 0.055458f
C387 VTAIL.n115 B 0.024833f
C388 VTAIL.n116 B 0.023406f
C389 VTAIL.n117 B 0.014008f
C390 VTAIL.n118 B 0.9255f
C391 VTAIL.n119 B 0.026069f
C392 VTAIL.n120 B 0.014008f
C393 VTAIL.n121 B 0.014832f
C394 VTAIL.n122 B 0.03311f
C395 VTAIL.n123 B 0.03311f
C396 VTAIL.n124 B 0.014832f
C397 VTAIL.n125 B 0.014008f
C398 VTAIL.n126 B 0.026069f
C399 VTAIL.n127 B 0.026069f
C400 VTAIL.n128 B 0.014008f
C401 VTAIL.n129 B 0.014832f
C402 VTAIL.n130 B 0.03311f
C403 VTAIL.n131 B 0.03311f
C404 VTAIL.n132 B 0.014832f
C405 VTAIL.n133 B 0.014008f
C406 VTAIL.n134 B 0.026069f
C407 VTAIL.n135 B 0.026069f
C408 VTAIL.n136 B 0.014008f
C409 VTAIL.n137 B 0.01442f
C410 VTAIL.n138 B 0.01442f
C411 VTAIL.n139 B 0.03311f
C412 VTAIL.n140 B 0.06919f
C413 VTAIL.n141 B 0.014832f
C414 VTAIL.n142 B 0.014008f
C415 VTAIL.n143 B 0.06453f
C416 VTAIL.n144 B 0.038586f
C417 VTAIL.n145 B 1.59967f
C418 VTAIL.n146 B 0.035235f
C419 VTAIL.n147 B 0.026069f
C420 VTAIL.n148 B 0.014008f
C421 VTAIL.n149 B 0.03311f
C422 VTAIL.n150 B 0.014832f
C423 VTAIL.n151 B 0.026069f
C424 VTAIL.n152 B 0.014008f
C425 VTAIL.n153 B 0.03311f
C426 VTAIL.n154 B 0.014832f
C427 VTAIL.n155 B 0.026069f
C428 VTAIL.n156 B 0.014008f
C429 VTAIL.n157 B 0.03311f
C430 VTAIL.n158 B 0.014832f
C431 VTAIL.n159 B 0.15434f
C432 VTAIL.t2 B 0.055458f
C433 VTAIL.n160 B 0.024833f
C434 VTAIL.n161 B 0.023406f
C435 VTAIL.n162 B 0.014008f
C436 VTAIL.n163 B 0.9255f
C437 VTAIL.n164 B 0.026069f
C438 VTAIL.n165 B 0.014008f
C439 VTAIL.n166 B 0.014832f
C440 VTAIL.n167 B 0.03311f
C441 VTAIL.n168 B 0.03311f
C442 VTAIL.n169 B 0.014832f
C443 VTAIL.n170 B 0.014008f
C444 VTAIL.n171 B 0.026069f
C445 VTAIL.n172 B 0.026069f
C446 VTAIL.n173 B 0.014008f
C447 VTAIL.n174 B 0.014832f
C448 VTAIL.n175 B 0.03311f
C449 VTAIL.n176 B 0.03311f
C450 VTAIL.n177 B 0.03311f
C451 VTAIL.n178 B 0.014832f
C452 VTAIL.n179 B 0.014008f
C453 VTAIL.n180 B 0.026069f
C454 VTAIL.n181 B 0.026069f
C455 VTAIL.n182 B 0.014008f
C456 VTAIL.n183 B 0.01442f
C457 VTAIL.n184 B 0.01442f
C458 VTAIL.n185 B 0.03311f
C459 VTAIL.n186 B 0.06919f
C460 VTAIL.n187 B 0.014832f
C461 VTAIL.n188 B 0.014008f
C462 VTAIL.n189 B 0.06453f
C463 VTAIL.n190 B 0.038586f
C464 VTAIL.n191 B 1.52038f
C465 VP.t1 B 1.76352f
C466 VP.n0 B 0.70807f
C467 VP.n1 B 0.020041f
C468 VP.n2 B 0.03858f
C469 VP.n3 B 0.020041f
C470 VP.n4 B 0.037539f
C471 VP.n5 B 0.020041f
C472 VP.t3 B 1.76352f
C473 VP.n6 B 0.04071f
C474 VP.n7 B 0.020041f
C475 VP.n8 B 0.037539f
C476 VP.t0 B 1.76352f
C477 VP.n9 B 0.70807f
C478 VP.n10 B 0.020041f
C479 VP.n11 B 0.03858f
C480 VP.n12 B 0.020041f
C481 VP.n13 B 0.037539f
C482 VP.t2 B 2.06226f
C483 VP.t5 B 1.76352f
C484 VP.n14 B 0.712954f
C485 VP.n15 B 0.674264f
C486 VP.n16 B 0.256295f
C487 VP.n17 B 0.020041f
C488 VP.n18 B 0.037539f
C489 VP.n19 B 0.04071f
C490 VP.n20 B 0.017016f
C491 VP.n21 B 0.020041f
C492 VP.n22 B 0.020041f
C493 VP.n23 B 0.020041f
C494 VP.n24 B 0.037539f
C495 VP.n25 B 0.037539f
C496 VP.n26 B 0.023082f
C497 VP.n27 B 0.032351f
C498 VP.n28 B 1.17993f
C499 VP.n29 B 1.19406f
C500 VP.t4 B 1.76352f
C501 VP.n30 B 0.70807f
C502 VP.n31 B 0.023082f
C503 VP.n32 B 0.032351f
C504 VP.n33 B 0.020041f
C505 VP.n34 B 0.020041f
C506 VP.n35 B 0.037539f
C507 VP.n36 B 0.03858f
C508 VP.n37 B 0.017016f
C509 VP.n38 B 0.020041f
C510 VP.n39 B 0.020041f
C511 VP.n40 B 0.020041f
C512 VP.n41 B 0.037539f
C513 VP.n42 B 0.037539f
C514 VP.n43 B 0.648966f
C515 VP.n44 B 0.020041f
C516 VP.n45 B 0.020041f
C517 VP.n46 B 0.020041f
C518 VP.n47 B 0.037539f
C519 VP.n48 B 0.04071f
C520 VP.n49 B 0.017016f
C521 VP.n50 B 0.020041f
C522 VP.n51 B 0.020041f
C523 VP.n52 B 0.020041f
C524 VP.n53 B 0.037539f
C525 VP.n54 B 0.037539f
C526 VP.n55 B 0.023082f
C527 VP.n56 B 0.032351f
C528 VP.n57 B 0.059876f
.ends

