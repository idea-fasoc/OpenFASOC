* NGSPICE file created from diff_pair_sample_1377.ext - technology: sky130A

.subckt diff_pair_sample_1377 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t10 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0.4026 ps=2.77 w=2.44 l=1.68
X1 VDD1.t5 VP.t0 VTAIL.t5 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.9516 ps=5.66 w=2.44 l=1.68
X2 B.t11 B.t9 B.t10 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0 ps=0 w=2.44 l=1.68
X3 VDD1.t4 VP.t1 VTAIL.t2 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0.4026 ps=2.77 w=2.44 l=1.68
X4 VDD2.t4 VN.t1 VTAIL.t7 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.9516 ps=5.66 w=2.44 l=1.68
X5 VDD2.t3 VN.t2 VTAIL.t11 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.9516 ps=5.66 w=2.44 l=1.68
X6 B.t8 B.t6 B.t7 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0 ps=0 w=2.44 l=1.68
X7 VTAIL.t3 VP.t2 VDD1.t3 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.4026 ps=2.77 w=2.44 l=1.68
X8 VTAIL.t9 VN.t3 VDD2.t2 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.4026 ps=2.77 w=2.44 l=1.68
X9 VTAIL.t8 VN.t4 VDD2.t1 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.4026 ps=2.77 w=2.44 l=1.68
X10 VDD1.t2 VP.t3 VTAIL.t4 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0.4026 ps=2.77 w=2.44 l=1.68
X11 VDD2.t0 VN.t5 VTAIL.t6 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0.4026 ps=2.77 w=2.44 l=1.68
X12 B.t5 B.t3 B.t4 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0 ps=0 w=2.44 l=1.68
X13 VTAIL.t0 VP.t4 VDD1.t1 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.4026 ps=2.77 w=2.44 l=1.68
X14 VDD1.t0 VP.t5 VTAIL.t1 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.4026 pd=2.77 as=0.9516 ps=5.66 w=2.44 l=1.68
X15 B.t2 B.t0 B.t1 w_n2578_n1456# sky130_fd_pr__pfet_01v8 ad=0.9516 pd=5.66 as=0 ps=0 w=2.44 l=1.68
R0 VN.n11 VN.n10 185.4
R1 VN.n23 VN.n22 185.4
R2 VN.n21 VN.n12 161.3
R3 VN.n20 VN.n19 161.3
R4 VN.n18 VN.n13 161.3
R5 VN.n17 VN.n16 161.3
R6 VN.n9 VN.n0 161.3
R7 VN.n8 VN.n7 161.3
R8 VN.n6 VN.n1 161.3
R9 VN.n5 VN.n4 161.3
R10 VN.n2 VN.t0 67.6592
R11 VN.n14 VN.t2 67.6592
R12 VN.n15 VN.n14 44.7528
R13 VN.n3 VN.n2 44.7528
R14 VN.n8 VN.n1 41.0614
R15 VN.n20 VN.n13 41.0614
R16 VN.n4 VN.n1 40.0926
R17 VN.n16 VN.n13 40.0926
R18 VN VN.n23 38.0289
R19 VN.n3 VN.t3 35.0029
R20 VN.n10 VN.t1 35.0029
R21 VN.n15 VN.t4 35.0029
R22 VN.n22 VN.t5 35.0029
R23 VN.n4 VN.n3 24.5923
R24 VN.n9 VN.n8 24.5923
R25 VN.n16 VN.n15 24.5923
R26 VN.n21 VN.n20 24.5923
R27 VN.n17 VN.n14 12.4791
R28 VN.n5 VN.n2 12.4791
R29 VN.n10 VN.n9 0.492337
R30 VN.n22 VN.n21 0.492337
R31 VN.n23 VN.n12 0.189894
R32 VN.n19 VN.n12 0.189894
R33 VN.n19 VN.n18 0.189894
R34 VN.n18 VN.n17 0.189894
R35 VN.n6 VN.n5 0.189894
R36 VN.n7 VN.n6 0.189894
R37 VN.n7 VN.n0 0.189894
R38 VN.n11 VN.n0 0.189894
R39 VN VN.n11 0.0516364
R40 VTAIL.n50 VTAIL.n44 756.745
R41 VTAIL.n8 VTAIL.n2 756.745
R42 VTAIL.n38 VTAIL.n32 756.745
R43 VTAIL.n24 VTAIL.n18 756.745
R44 VTAIL.n49 VTAIL.n48 585
R45 VTAIL.n51 VTAIL.n50 585
R46 VTAIL.n7 VTAIL.n6 585
R47 VTAIL.n9 VTAIL.n8 585
R48 VTAIL.n39 VTAIL.n38 585
R49 VTAIL.n37 VTAIL.n36 585
R50 VTAIL.n25 VTAIL.n24 585
R51 VTAIL.n23 VTAIL.n22 585
R52 VTAIL.n47 VTAIL.t7 355.474
R53 VTAIL.n5 VTAIL.t5 355.474
R54 VTAIL.n35 VTAIL.t1 355.474
R55 VTAIL.n21 VTAIL.t11 355.474
R56 VTAIL.n50 VTAIL.n49 171.744
R57 VTAIL.n8 VTAIL.n7 171.744
R58 VTAIL.n38 VTAIL.n37 171.744
R59 VTAIL.n24 VTAIL.n23 171.744
R60 VTAIL.n31 VTAIL.n30 135.817
R61 VTAIL.n17 VTAIL.n16 135.817
R62 VTAIL.n1 VTAIL.n0 135.817
R63 VTAIL.n15 VTAIL.n14 135.817
R64 VTAIL.n49 VTAIL.t7 85.8723
R65 VTAIL.n7 VTAIL.t5 85.8723
R66 VTAIL.n37 VTAIL.t1 85.8723
R67 VTAIL.n23 VTAIL.t11 85.8723
R68 VTAIL.n55 VTAIL.n54 32.9611
R69 VTAIL.n13 VTAIL.n12 32.9611
R70 VTAIL.n43 VTAIL.n42 32.9611
R71 VTAIL.n29 VTAIL.n28 32.9611
R72 VTAIL.n17 VTAIL.n15 17.9358
R73 VTAIL.n55 VTAIL.n43 16.2031
R74 VTAIL.n48 VTAIL.n47 15.8418
R75 VTAIL.n6 VTAIL.n5 15.8418
R76 VTAIL.n36 VTAIL.n35 15.8418
R77 VTAIL.n22 VTAIL.n21 15.8418
R78 VTAIL.n0 VTAIL.t10 13.3222
R79 VTAIL.n0 VTAIL.t9 13.3222
R80 VTAIL.n14 VTAIL.t2 13.3222
R81 VTAIL.n14 VTAIL.t3 13.3222
R82 VTAIL.n30 VTAIL.t4 13.3222
R83 VTAIL.n30 VTAIL.t0 13.3222
R84 VTAIL.n16 VTAIL.t6 13.3222
R85 VTAIL.n16 VTAIL.t8 13.3222
R86 VTAIL.n51 VTAIL.n46 12.8005
R87 VTAIL.n9 VTAIL.n4 12.8005
R88 VTAIL.n39 VTAIL.n34 12.8005
R89 VTAIL.n25 VTAIL.n20 12.8005
R90 VTAIL.n52 VTAIL.n44 12.0247
R91 VTAIL.n10 VTAIL.n2 12.0247
R92 VTAIL.n40 VTAIL.n32 12.0247
R93 VTAIL.n26 VTAIL.n18 12.0247
R94 VTAIL.n54 VTAIL.n53 9.45567
R95 VTAIL.n12 VTAIL.n11 9.45567
R96 VTAIL.n42 VTAIL.n41 9.45567
R97 VTAIL.n28 VTAIL.n27 9.45567
R98 VTAIL.n53 VTAIL.n52 9.3005
R99 VTAIL.n46 VTAIL.n45 9.3005
R100 VTAIL.n11 VTAIL.n10 9.3005
R101 VTAIL.n4 VTAIL.n3 9.3005
R102 VTAIL.n41 VTAIL.n40 9.3005
R103 VTAIL.n34 VTAIL.n33 9.3005
R104 VTAIL.n27 VTAIL.n26 9.3005
R105 VTAIL.n20 VTAIL.n19 9.3005
R106 VTAIL.n35 VTAIL.n33 4.29255
R107 VTAIL.n21 VTAIL.n19 4.29255
R108 VTAIL.n47 VTAIL.n45 4.29255
R109 VTAIL.n5 VTAIL.n3 4.29255
R110 VTAIL.n54 VTAIL.n44 1.93989
R111 VTAIL.n12 VTAIL.n2 1.93989
R112 VTAIL.n42 VTAIL.n32 1.93989
R113 VTAIL.n28 VTAIL.n18 1.93989
R114 VTAIL.n29 VTAIL.n17 1.73326
R115 VTAIL.n43 VTAIL.n31 1.73326
R116 VTAIL.n15 VTAIL.n13 1.73326
R117 VTAIL.n31 VTAIL.n29 1.33671
R118 VTAIL.n13 VTAIL.n1 1.33671
R119 VTAIL VTAIL.n55 1.24188
R120 VTAIL.n52 VTAIL.n51 1.16414
R121 VTAIL.n10 VTAIL.n9 1.16414
R122 VTAIL.n40 VTAIL.n39 1.16414
R123 VTAIL.n26 VTAIL.n25 1.16414
R124 VTAIL VTAIL.n1 0.491879
R125 VTAIL.n48 VTAIL.n46 0.388379
R126 VTAIL.n6 VTAIL.n4 0.388379
R127 VTAIL.n36 VTAIL.n34 0.388379
R128 VTAIL.n22 VTAIL.n20 0.388379
R129 VTAIL.n53 VTAIL.n45 0.155672
R130 VTAIL.n11 VTAIL.n3 0.155672
R131 VTAIL.n41 VTAIL.n33 0.155672
R132 VTAIL.n27 VTAIL.n19 0.155672
R133 VDD2.n19 VDD2.n13 756.745
R134 VDD2.n6 VDD2.n0 756.745
R135 VDD2.n20 VDD2.n19 585
R136 VDD2.n18 VDD2.n17 585
R137 VDD2.n5 VDD2.n4 585
R138 VDD2.n7 VDD2.n6 585
R139 VDD2.n16 VDD2.t0 355.474
R140 VDD2.n3 VDD2.t5 355.474
R141 VDD2.n19 VDD2.n18 171.744
R142 VDD2.n6 VDD2.n5 171.744
R143 VDD2.n12 VDD2.n11 152.874
R144 VDD2 VDD2.n25 152.87
R145 VDD2.n18 VDD2.t0 85.8723
R146 VDD2.n5 VDD2.t5 85.8723
R147 VDD2.n12 VDD2.n10 50.8841
R148 VDD2.n24 VDD2.n23 49.6399
R149 VDD2.n24 VDD2.n12 31.4502
R150 VDD2.n17 VDD2.n16 15.8418
R151 VDD2.n4 VDD2.n3 15.8418
R152 VDD2.n25 VDD2.t1 13.3222
R153 VDD2.n25 VDD2.t3 13.3222
R154 VDD2.n11 VDD2.t2 13.3222
R155 VDD2.n11 VDD2.t4 13.3222
R156 VDD2.n20 VDD2.n15 12.8005
R157 VDD2.n7 VDD2.n2 12.8005
R158 VDD2.n21 VDD2.n13 12.0247
R159 VDD2.n8 VDD2.n0 12.0247
R160 VDD2.n23 VDD2.n22 9.45567
R161 VDD2.n10 VDD2.n9 9.45567
R162 VDD2.n22 VDD2.n21 9.3005
R163 VDD2.n15 VDD2.n14 9.3005
R164 VDD2.n9 VDD2.n8 9.3005
R165 VDD2.n2 VDD2.n1 9.3005
R166 VDD2.n16 VDD2.n14 4.29255
R167 VDD2.n3 VDD2.n1 4.29255
R168 VDD2.n23 VDD2.n13 1.93989
R169 VDD2.n10 VDD2.n0 1.93989
R170 VDD2 VDD2.n24 1.35826
R171 VDD2.n21 VDD2.n20 1.16414
R172 VDD2.n8 VDD2.n7 1.16414
R173 VDD2.n17 VDD2.n15 0.388379
R174 VDD2.n4 VDD2.n2 0.388379
R175 VDD2.n22 VDD2.n14 0.155672
R176 VDD2.n9 VDD2.n1 0.155672
R177 VP.n18 VP.n17 185.4
R178 VP.n33 VP.n32 185.4
R179 VP.n16 VP.n15 185.4
R180 VP.n10 VP.n9 161.3
R181 VP.n11 VP.n6 161.3
R182 VP.n13 VP.n12 161.3
R183 VP.n14 VP.n5 161.3
R184 VP.n31 VP.n0 161.3
R185 VP.n30 VP.n29 161.3
R186 VP.n28 VP.n1 161.3
R187 VP.n27 VP.n26 161.3
R188 VP.n25 VP.n2 161.3
R189 VP.n24 VP.n23 161.3
R190 VP.n22 VP.n3 161.3
R191 VP.n21 VP.n20 161.3
R192 VP.n19 VP.n4 161.3
R193 VP.n7 VP.t3 67.6592
R194 VP.n8 VP.n7 44.7528
R195 VP.n20 VP.n3 41.0614
R196 VP.n30 VP.n1 41.0614
R197 VP.n13 VP.n6 41.0614
R198 VP.n24 VP.n3 40.0926
R199 VP.n26 VP.n1 40.0926
R200 VP.n9 VP.n6 40.0926
R201 VP.n17 VP.n16 37.6482
R202 VP.n25 VP.t2 35.0029
R203 VP.n18 VP.t1 35.0029
R204 VP.n32 VP.t0 35.0029
R205 VP.n8 VP.t4 35.0029
R206 VP.n15 VP.t5 35.0029
R207 VP.n20 VP.n19 24.5923
R208 VP.n25 VP.n24 24.5923
R209 VP.n26 VP.n25 24.5923
R210 VP.n31 VP.n30 24.5923
R211 VP.n14 VP.n13 24.5923
R212 VP.n9 VP.n8 24.5923
R213 VP.n10 VP.n7 12.4791
R214 VP.n19 VP.n18 0.492337
R215 VP.n32 VP.n31 0.492337
R216 VP.n15 VP.n14 0.492337
R217 VP.n11 VP.n10 0.189894
R218 VP.n12 VP.n11 0.189894
R219 VP.n12 VP.n5 0.189894
R220 VP.n16 VP.n5 0.189894
R221 VP.n17 VP.n4 0.189894
R222 VP.n21 VP.n4 0.189894
R223 VP.n22 VP.n21 0.189894
R224 VP.n23 VP.n22 0.189894
R225 VP.n23 VP.n2 0.189894
R226 VP.n27 VP.n2 0.189894
R227 VP.n28 VP.n27 0.189894
R228 VP.n29 VP.n28 0.189894
R229 VP.n29 VP.n0 0.189894
R230 VP.n33 VP.n0 0.189894
R231 VP VP.n33 0.0516364
R232 VDD1.n6 VDD1.n0 756.745
R233 VDD1.n17 VDD1.n11 756.745
R234 VDD1.n7 VDD1.n6 585
R235 VDD1.n5 VDD1.n4 585
R236 VDD1.n16 VDD1.n15 585
R237 VDD1.n18 VDD1.n17 585
R238 VDD1.n3 VDD1.t2 355.474
R239 VDD1.n14 VDD1.t4 355.474
R240 VDD1.n6 VDD1.n5 171.744
R241 VDD1.n17 VDD1.n16 171.744
R242 VDD1.n23 VDD1.n22 152.874
R243 VDD1.n25 VDD1.n24 152.495
R244 VDD1.n5 VDD1.t2 85.8723
R245 VDD1.n16 VDD1.t4 85.8723
R246 VDD1 VDD1.n10 50.9977
R247 VDD1.n23 VDD1.n21 50.8841
R248 VDD1.n25 VDD1.n23 32.8996
R249 VDD1.n4 VDD1.n3 15.8418
R250 VDD1.n15 VDD1.n14 15.8418
R251 VDD1.n24 VDD1.t1 13.3222
R252 VDD1.n24 VDD1.t0 13.3222
R253 VDD1.n22 VDD1.t3 13.3222
R254 VDD1.n22 VDD1.t5 13.3222
R255 VDD1.n7 VDD1.n2 12.8005
R256 VDD1.n18 VDD1.n13 12.8005
R257 VDD1.n8 VDD1.n0 12.0247
R258 VDD1.n19 VDD1.n11 12.0247
R259 VDD1.n10 VDD1.n9 9.45567
R260 VDD1.n21 VDD1.n20 9.45567
R261 VDD1.n9 VDD1.n8 9.3005
R262 VDD1.n2 VDD1.n1 9.3005
R263 VDD1.n20 VDD1.n19 9.3005
R264 VDD1.n13 VDD1.n12 9.3005
R265 VDD1.n3 VDD1.n1 4.29255
R266 VDD1.n14 VDD1.n12 4.29255
R267 VDD1.n10 VDD1.n0 1.93989
R268 VDD1.n21 VDD1.n11 1.93989
R269 VDD1.n8 VDD1.n7 1.16414
R270 VDD1.n19 VDD1.n18 1.16414
R271 VDD1.n4 VDD1.n2 0.388379
R272 VDD1.n15 VDD1.n13 0.388379
R273 VDD1 VDD1.n25 0.3755
R274 VDD1.n9 VDD1.n1 0.155672
R275 VDD1.n20 VDD1.n12 0.155672
R276 B.n212 B.n73 585
R277 B.n211 B.n210 585
R278 B.n209 B.n74 585
R279 B.n208 B.n207 585
R280 B.n206 B.n75 585
R281 B.n205 B.n204 585
R282 B.n203 B.n76 585
R283 B.n202 B.n201 585
R284 B.n200 B.n77 585
R285 B.n199 B.n198 585
R286 B.n197 B.n78 585
R287 B.n196 B.n195 585
R288 B.n194 B.n79 585
R289 B.n193 B.n192 585
R290 B.n190 B.n80 585
R291 B.n189 B.n188 585
R292 B.n187 B.n83 585
R293 B.n186 B.n185 585
R294 B.n184 B.n84 585
R295 B.n183 B.n182 585
R296 B.n181 B.n85 585
R297 B.n180 B.n179 585
R298 B.n178 B.n86 585
R299 B.n176 B.n175 585
R300 B.n174 B.n89 585
R301 B.n173 B.n172 585
R302 B.n171 B.n90 585
R303 B.n170 B.n169 585
R304 B.n168 B.n91 585
R305 B.n167 B.n166 585
R306 B.n165 B.n92 585
R307 B.n164 B.n163 585
R308 B.n162 B.n93 585
R309 B.n161 B.n160 585
R310 B.n159 B.n94 585
R311 B.n158 B.n157 585
R312 B.n156 B.n95 585
R313 B.n214 B.n213 585
R314 B.n215 B.n72 585
R315 B.n217 B.n216 585
R316 B.n218 B.n71 585
R317 B.n220 B.n219 585
R318 B.n221 B.n70 585
R319 B.n223 B.n222 585
R320 B.n224 B.n69 585
R321 B.n226 B.n225 585
R322 B.n227 B.n68 585
R323 B.n229 B.n228 585
R324 B.n230 B.n67 585
R325 B.n232 B.n231 585
R326 B.n233 B.n66 585
R327 B.n235 B.n234 585
R328 B.n236 B.n65 585
R329 B.n238 B.n237 585
R330 B.n239 B.n64 585
R331 B.n241 B.n240 585
R332 B.n242 B.n63 585
R333 B.n244 B.n243 585
R334 B.n245 B.n62 585
R335 B.n247 B.n246 585
R336 B.n248 B.n61 585
R337 B.n250 B.n249 585
R338 B.n251 B.n60 585
R339 B.n253 B.n252 585
R340 B.n254 B.n59 585
R341 B.n256 B.n255 585
R342 B.n257 B.n58 585
R343 B.n259 B.n258 585
R344 B.n260 B.n57 585
R345 B.n262 B.n261 585
R346 B.n263 B.n56 585
R347 B.n265 B.n264 585
R348 B.n266 B.n55 585
R349 B.n268 B.n267 585
R350 B.n269 B.n54 585
R351 B.n271 B.n270 585
R352 B.n272 B.n53 585
R353 B.n274 B.n273 585
R354 B.n275 B.n52 585
R355 B.n277 B.n276 585
R356 B.n278 B.n51 585
R357 B.n280 B.n279 585
R358 B.n281 B.n50 585
R359 B.n283 B.n282 585
R360 B.n284 B.n49 585
R361 B.n286 B.n285 585
R362 B.n287 B.n48 585
R363 B.n289 B.n288 585
R364 B.n290 B.n47 585
R365 B.n292 B.n291 585
R366 B.n293 B.n46 585
R367 B.n295 B.n294 585
R368 B.n296 B.n45 585
R369 B.n298 B.n297 585
R370 B.n299 B.n44 585
R371 B.n301 B.n300 585
R372 B.n302 B.n43 585
R373 B.n304 B.n303 585
R374 B.n305 B.n42 585
R375 B.n307 B.n306 585
R376 B.n308 B.n41 585
R377 B.n365 B.n364 585
R378 B.n363 B.n18 585
R379 B.n362 B.n361 585
R380 B.n360 B.n19 585
R381 B.n359 B.n358 585
R382 B.n357 B.n20 585
R383 B.n356 B.n355 585
R384 B.n354 B.n21 585
R385 B.n353 B.n352 585
R386 B.n351 B.n22 585
R387 B.n350 B.n349 585
R388 B.n348 B.n23 585
R389 B.n347 B.n346 585
R390 B.n345 B.n24 585
R391 B.n344 B.n343 585
R392 B.n342 B.n25 585
R393 B.n341 B.n340 585
R394 B.n339 B.n29 585
R395 B.n338 B.n337 585
R396 B.n336 B.n30 585
R397 B.n335 B.n334 585
R398 B.n333 B.n31 585
R399 B.n332 B.n331 585
R400 B.n329 B.n32 585
R401 B.n328 B.n327 585
R402 B.n326 B.n35 585
R403 B.n325 B.n324 585
R404 B.n323 B.n36 585
R405 B.n322 B.n321 585
R406 B.n320 B.n37 585
R407 B.n319 B.n318 585
R408 B.n317 B.n38 585
R409 B.n316 B.n315 585
R410 B.n314 B.n39 585
R411 B.n313 B.n312 585
R412 B.n311 B.n40 585
R413 B.n310 B.n309 585
R414 B.n366 B.n17 585
R415 B.n368 B.n367 585
R416 B.n369 B.n16 585
R417 B.n371 B.n370 585
R418 B.n372 B.n15 585
R419 B.n374 B.n373 585
R420 B.n375 B.n14 585
R421 B.n377 B.n376 585
R422 B.n378 B.n13 585
R423 B.n380 B.n379 585
R424 B.n381 B.n12 585
R425 B.n383 B.n382 585
R426 B.n384 B.n11 585
R427 B.n386 B.n385 585
R428 B.n387 B.n10 585
R429 B.n389 B.n388 585
R430 B.n390 B.n9 585
R431 B.n392 B.n391 585
R432 B.n393 B.n8 585
R433 B.n395 B.n394 585
R434 B.n396 B.n7 585
R435 B.n398 B.n397 585
R436 B.n399 B.n6 585
R437 B.n401 B.n400 585
R438 B.n402 B.n5 585
R439 B.n404 B.n403 585
R440 B.n405 B.n4 585
R441 B.n407 B.n406 585
R442 B.n408 B.n3 585
R443 B.n410 B.n409 585
R444 B.n411 B.n0 585
R445 B.n2 B.n1 585
R446 B.n111 B.n110 585
R447 B.n113 B.n112 585
R448 B.n114 B.n109 585
R449 B.n116 B.n115 585
R450 B.n117 B.n108 585
R451 B.n119 B.n118 585
R452 B.n120 B.n107 585
R453 B.n122 B.n121 585
R454 B.n123 B.n106 585
R455 B.n125 B.n124 585
R456 B.n126 B.n105 585
R457 B.n128 B.n127 585
R458 B.n129 B.n104 585
R459 B.n131 B.n130 585
R460 B.n132 B.n103 585
R461 B.n134 B.n133 585
R462 B.n135 B.n102 585
R463 B.n137 B.n136 585
R464 B.n138 B.n101 585
R465 B.n140 B.n139 585
R466 B.n141 B.n100 585
R467 B.n143 B.n142 585
R468 B.n144 B.n99 585
R469 B.n146 B.n145 585
R470 B.n147 B.n98 585
R471 B.n149 B.n148 585
R472 B.n150 B.n97 585
R473 B.n152 B.n151 585
R474 B.n153 B.n96 585
R475 B.n155 B.n154 585
R476 B.n156 B.n155 506.916
R477 B.n213 B.n212 506.916
R478 B.n309 B.n308 506.916
R479 B.n364 B.n17 506.916
R480 B.n81 B.t10 262.07
R481 B.n33 B.t2 262.07
R482 B.n87 B.t4 262.07
R483 B.n26 B.t8 262.07
R484 B.n413 B.n412 256.663
R485 B.n87 B.t3 241.055
R486 B.n81 B.t9 241.055
R487 B.n33 B.t0 241.055
R488 B.n26 B.t6 241.055
R489 B.n412 B.n411 235.042
R490 B.n412 B.n2 235.042
R491 B.n82 B.t11 223.088
R492 B.n34 B.t1 223.088
R493 B.n88 B.t5 223.088
R494 B.n27 B.t7 223.088
R495 B.n157 B.n156 163.367
R496 B.n157 B.n94 163.367
R497 B.n161 B.n94 163.367
R498 B.n162 B.n161 163.367
R499 B.n163 B.n162 163.367
R500 B.n163 B.n92 163.367
R501 B.n167 B.n92 163.367
R502 B.n168 B.n167 163.367
R503 B.n169 B.n168 163.367
R504 B.n169 B.n90 163.367
R505 B.n173 B.n90 163.367
R506 B.n174 B.n173 163.367
R507 B.n175 B.n174 163.367
R508 B.n175 B.n86 163.367
R509 B.n180 B.n86 163.367
R510 B.n181 B.n180 163.367
R511 B.n182 B.n181 163.367
R512 B.n182 B.n84 163.367
R513 B.n186 B.n84 163.367
R514 B.n187 B.n186 163.367
R515 B.n188 B.n187 163.367
R516 B.n188 B.n80 163.367
R517 B.n193 B.n80 163.367
R518 B.n194 B.n193 163.367
R519 B.n195 B.n194 163.367
R520 B.n195 B.n78 163.367
R521 B.n199 B.n78 163.367
R522 B.n200 B.n199 163.367
R523 B.n201 B.n200 163.367
R524 B.n201 B.n76 163.367
R525 B.n205 B.n76 163.367
R526 B.n206 B.n205 163.367
R527 B.n207 B.n206 163.367
R528 B.n207 B.n74 163.367
R529 B.n211 B.n74 163.367
R530 B.n212 B.n211 163.367
R531 B.n308 B.n307 163.367
R532 B.n307 B.n42 163.367
R533 B.n303 B.n42 163.367
R534 B.n303 B.n302 163.367
R535 B.n302 B.n301 163.367
R536 B.n301 B.n44 163.367
R537 B.n297 B.n44 163.367
R538 B.n297 B.n296 163.367
R539 B.n296 B.n295 163.367
R540 B.n295 B.n46 163.367
R541 B.n291 B.n46 163.367
R542 B.n291 B.n290 163.367
R543 B.n290 B.n289 163.367
R544 B.n289 B.n48 163.367
R545 B.n285 B.n48 163.367
R546 B.n285 B.n284 163.367
R547 B.n284 B.n283 163.367
R548 B.n283 B.n50 163.367
R549 B.n279 B.n50 163.367
R550 B.n279 B.n278 163.367
R551 B.n278 B.n277 163.367
R552 B.n277 B.n52 163.367
R553 B.n273 B.n52 163.367
R554 B.n273 B.n272 163.367
R555 B.n272 B.n271 163.367
R556 B.n271 B.n54 163.367
R557 B.n267 B.n54 163.367
R558 B.n267 B.n266 163.367
R559 B.n266 B.n265 163.367
R560 B.n265 B.n56 163.367
R561 B.n261 B.n56 163.367
R562 B.n261 B.n260 163.367
R563 B.n260 B.n259 163.367
R564 B.n259 B.n58 163.367
R565 B.n255 B.n58 163.367
R566 B.n255 B.n254 163.367
R567 B.n254 B.n253 163.367
R568 B.n253 B.n60 163.367
R569 B.n249 B.n60 163.367
R570 B.n249 B.n248 163.367
R571 B.n248 B.n247 163.367
R572 B.n247 B.n62 163.367
R573 B.n243 B.n62 163.367
R574 B.n243 B.n242 163.367
R575 B.n242 B.n241 163.367
R576 B.n241 B.n64 163.367
R577 B.n237 B.n64 163.367
R578 B.n237 B.n236 163.367
R579 B.n236 B.n235 163.367
R580 B.n235 B.n66 163.367
R581 B.n231 B.n66 163.367
R582 B.n231 B.n230 163.367
R583 B.n230 B.n229 163.367
R584 B.n229 B.n68 163.367
R585 B.n225 B.n68 163.367
R586 B.n225 B.n224 163.367
R587 B.n224 B.n223 163.367
R588 B.n223 B.n70 163.367
R589 B.n219 B.n70 163.367
R590 B.n219 B.n218 163.367
R591 B.n218 B.n217 163.367
R592 B.n217 B.n72 163.367
R593 B.n213 B.n72 163.367
R594 B.n364 B.n363 163.367
R595 B.n363 B.n362 163.367
R596 B.n362 B.n19 163.367
R597 B.n358 B.n19 163.367
R598 B.n358 B.n357 163.367
R599 B.n357 B.n356 163.367
R600 B.n356 B.n21 163.367
R601 B.n352 B.n21 163.367
R602 B.n352 B.n351 163.367
R603 B.n351 B.n350 163.367
R604 B.n350 B.n23 163.367
R605 B.n346 B.n23 163.367
R606 B.n346 B.n345 163.367
R607 B.n345 B.n344 163.367
R608 B.n344 B.n25 163.367
R609 B.n340 B.n25 163.367
R610 B.n340 B.n339 163.367
R611 B.n339 B.n338 163.367
R612 B.n338 B.n30 163.367
R613 B.n334 B.n30 163.367
R614 B.n334 B.n333 163.367
R615 B.n333 B.n332 163.367
R616 B.n332 B.n32 163.367
R617 B.n327 B.n32 163.367
R618 B.n327 B.n326 163.367
R619 B.n326 B.n325 163.367
R620 B.n325 B.n36 163.367
R621 B.n321 B.n36 163.367
R622 B.n321 B.n320 163.367
R623 B.n320 B.n319 163.367
R624 B.n319 B.n38 163.367
R625 B.n315 B.n38 163.367
R626 B.n315 B.n314 163.367
R627 B.n314 B.n313 163.367
R628 B.n313 B.n40 163.367
R629 B.n309 B.n40 163.367
R630 B.n368 B.n17 163.367
R631 B.n369 B.n368 163.367
R632 B.n370 B.n369 163.367
R633 B.n370 B.n15 163.367
R634 B.n374 B.n15 163.367
R635 B.n375 B.n374 163.367
R636 B.n376 B.n375 163.367
R637 B.n376 B.n13 163.367
R638 B.n380 B.n13 163.367
R639 B.n381 B.n380 163.367
R640 B.n382 B.n381 163.367
R641 B.n382 B.n11 163.367
R642 B.n386 B.n11 163.367
R643 B.n387 B.n386 163.367
R644 B.n388 B.n387 163.367
R645 B.n388 B.n9 163.367
R646 B.n392 B.n9 163.367
R647 B.n393 B.n392 163.367
R648 B.n394 B.n393 163.367
R649 B.n394 B.n7 163.367
R650 B.n398 B.n7 163.367
R651 B.n399 B.n398 163.367
R652 B.n400 B.n399 163.367
R653 B.n400 B.n5 163.367
R654 B.n404 B.n5 163.367
R655 B.n405 B.n404 163.367
R656 B.n406 B.n405 163.367
R657 B.n406 B.n3 163.367
R658 B.n410 B.n3 163.367
R659 B.n411 B.n410 163.367
R660 B.n110 B.n2 163.367
R661 B.n113 B.n110 163.367
R662 B.n114 B.n113 163.367
R663 B.n115 B.n114 163.367
R664 B.n115 B.n108 163.367
R665 B.n119 B.n108 163.367
R666 B.n120 B.n119 163.367
R667 B.n121 B.n120 163.367
R668 B.n121 B.n106 163.367
R669 B.n125 B.n106 163.367
R670 B.n126 B.n125 163.367
R671 B.n127 B.n126 163.367
R672 B.n127 B.n104 163.367
R673 B.n131 B.n104 163.367
R674 B.n132 B.n131 163.367
R675 B.n133 B.n132 163.367
R676 B.n133 B.n102 163.367
R677 B.n137 B.n102 163.367
R678 B.n138 B.n137 163.367
R679 B.n139 B.n138 163.367
R680 B.n139 B.n100 163.367
R681 B.n143 B.n100 163.367
R682 B.n144 B.n143 163.367
R683 B.n145 B.n144 163.367
R684 B.n145 B.n98 163.367
R685 B.n149 B.n98 163.367
R686 B.n150 B.n149 163.367
R687 B.n151 B.n150 163.367
R688 B.n151 B.n96 163.367
R689 B.n155 B.n96 163.367
R690 B.n177 B.n88 59.5399
R691 B.n191 B.n82 59.5399
R692 B.n330 B.n34 59.5399
R693 B.n28 B.n27 59.5399
R694 B.n88 B.n87 38.9823
R695 B.n82 B.n81 38.9823
R696 B.n34 B.n33 38.9823
R697 B.n27 B.n26 38.9823
R698 B.n366 B.n365 32.9371
R699 B.n310 B.n41 32.9371
R700 B.n214 B.n73 32.9371
R701 B.n154 B.n95 32.9371
R702 B B.n413 18.0485
R703 B.n367 B.n366 10.6151
R704 B.n367 B.n16 10.6151
R705 B.n371 B.n16 10.6151
R706 B.n372 B.n371 10.6151
R707 B.n373 B.n372 10.6151
R708 B.n373 B.n14 10.6151
R709 B.n377 B.n14 10.6151
R710 B.n378 B.n377 10.6151
R711 B.n379 B.n378 10.6151
R712 B.n379 B.n12 10.6151
R713 B.n383 B.n12 10.6151
R714 B.n384 B.n383 10.6151
R715 B.n385 B.n384 10.6151
R716 B.n385 B.n10 10.6151
R717 B.n389 B.n10 10.6151
R718 B.n390 B.n389 10.6151
R719 B.n391 B.n390 10.6151
R720 B.n391 B.n8 10.6151
R721 B.n395 B.n8 10.6151
R722 B.n396 B.n395 10.6151
R723 B.n397 B.n396 10.6151
R724 B.n397 B.n6 10.6151
R725 B.n401 B.n6 10.6151
R726 B.n402 B.n401 10.6151
R727 B.n403 B.n402 10.6151
R728 B.n403 B.n4 10.6151
R729 B.n407 B.n4 10.6151
R730 B.n408 B.n407 10.6151
R731 B.n409 B.n408 10.6151
R732 B.n409 B.n0 10.6151
R733 B.n365 B.n18 10.6151
R734 B.n361 B.n18 10.6151
R735 B.n361 B.n360 10.6151
R736 B.n360 B.n359 10.6151
R737 B.n359 B.n20 10.6151
R738 B.n355 B.n20 10.6151
R739 B.n355 B.n354 10.6151
R740 B.n354 B.n353 10.6151
R741 B.n353 B.n22 10.6151
R742 B.n349 B.n22 10.6151
R743 B.n349 B.n348 10.6151
R744 B.n348 B.n347 10.6151
R745 B.n347 B.n24 10.6151
R746 B.n343 B.n342 10.6151
R747 B.n342 B.n341 10.6151
R748 B.n341 B.n29 10.6151
R749 B.n337 B.n29 10.6151
R750 B.n337 B.n336 10.6151
R751 B.n336 B.n335 10.6151
R752 B.n335 B.n31 10.6151
R753 B.n331 B.n31 10.6151
R754 B.n329 B.n328 10.6151
R755 B.n328 B.n35 10.6151
R756 B.n324 B.n35 10.6151
R757 B.n324 B.n323 10.6151
R758 B.n323 B.n322 10.6151
R759 B.n322 B.n37 10.6151
R760 B.n318 B.n37 10.6151
R761 B.n318 B.n317 10.6151
R762 B.n317 B.n316 10.6151
R763 B.n316 B.n39 10.6151
R764 B.n312 B.n39 10.6151
R765 B.n312 B.n311 10.6151
R766 B.n311 B.n310 10.6151
R767 B.n306 B.n41 10.6151
R768 B.n306 B.n305 10.6151
R769 B.n305 B.n304 10.6151
R770 B.n304 B.n43 10.6151
R771 B.n300 B.n43 10.6151
R772 B.n300 B.n299 10.6151
R773 B.n299 B.n298 10.6151
R774 B.n298 B.n45 10.6151
R775 B.n294 B.n45 10.6151
R776 B.n294 B.n293 10.6151
R777 B.n293 B.n292 10.6151
R778 B.n292 B.n47 10.6151
R779 B.n288 B.n47 10.6151
R780 B.n288 B.n287 10.6151
R781 B.n287 B.n286 10.6151
R782 B.n286 B.n49 10.6151
R783 B.n282 B.n49 10.6151
R784 B.n282 B.n281 10.6151
R785 B.n281 B.n280 10.6151
R786 B.n280 B.n51 10.6151
R787 B.n276 B.n51 10.6151
R788 B.n276 B.n275 10.6151
R789 B.n275 B.n274 10.6151
R790 B.n274 B.n53 10.6151
R791 B.n270 B.n53 10.6151
R792 B.n270 B.n269 10.6151
R793 B.n269 B.n268 10.6151
R794 B.n268 B.n55 10.6151
R795 B.n264 B.n55 10.6151
R796 B.n264 B.n263 10.6151
R797 B.n263 B.n262 10.6151
R798 B.n262 B.n57 10.6151
R799 B.n258 B.n57 10.6151
R800 B.n258 B.n257 10.6151
R801 B.n257 B.n256 10.6151
R802 B.n256 B.n59 10.6151
R803 B.n252 B.n59 10.6151
R804 B.n252 B.n251 10.6151
R805 B.n251 B.n250 10.6151
R806 B.n250 B.n61 10.6151
R807 B.n246 B.n61 10.6151
R808 B.n246 B.n245 10.6151
R809 B.n245 B.n244 10.6151
R810 B.n244 B.n63 10.6151
R811 B.n240 B.n63 10.6151
R812 B.n240 B.n239 10.6151
R813 B.n239 B.n238 10.6151
R814 B.n238 B.n65 10.6151
R815 B.n234 B.n65 10.6151
R816 B.n234 B.n233 10.6151
R817 B.n233 B.n232 10.6151
R818 B.n232 B.n67 10.6151
R819 B.n228 B.n67 10.6151
R820 B.n228 B.n227 10.6151
R821 B.n227 B.n226 10.6151
R822 B.n226 B.n69 10.6151
R823 B.n222 B.n69 10.6151
R824 B.n222 B.n221 10.6151
R825 B.n221 B.n220 10.6151
R826 B.n220 B.n71 10.6151
R827 B.n216 B.n71 10.6151
R828 B.n216 B.n215 10.6151
R829 B.n215 B.n214 10.6151
R830 B.n111 B.n1 10.6151
R831 B.n112 B.n111 10.6151
R832 B.n112 B.n109 10.6151
R833 B.n116 B.n109 10.6151
R834 B.n117 B.n116 10.6151
R835 B.n118 B.n117 10.6151
R836 B.n118 B.n107 10.6151
R837 B.n122 B.n107 10.6151
R838 B.n123 B.n122 10.6151
R839 B.n124 B.n123 10.6151
R840 B.n124 B.n105 10.6151
R841 B.n128 B.n105 10.6151
R842 B.n129 B.n128 10.6151
R843 B.n130 B.n129 10.6151
R844 B.n130 B.n103 10.6151
R845 B.n134 B.n103 10.6151
R846 B.n135 B.n134 10.6151
R847 B.n136 B.n135 10.6151
R848 B.n136 B.n101 10.6151
R849 B.n140 B.n101 10.6151
R850 B.n141 B.n140 10.6151
R851 B.n142 B.n141 10.6151
R852 B.n142 B.n99 10.6151
R853 B.n146 B.n99 10.6151
R854 B.n147 B.n146 10.6151
R855 B.n148 B.n147 10.6151
R856 B.n148 B.n97 10.6151
R857 B.n152 B.n97 10.6151
R858 B.n153 B.n152 10.6151
R859 B.n154 B.n153 10.6151
R860 B.n158 B.n95 10.6151
R861 B.n159 B.n158 10.6151
R862 B.n160 B.n159 10.6151
R863 B.n160 B.n93 10.6151
R864 B.n164 B.n93 10.6151
R865 B.n165 B.n164 10.6151
R866 B.n166 B.n165 10.6151
R867 B.n166 B.n91 10.6151
R868 B.n170 B.n91 10.6151
R869 B.n171 B.n170 10.6151
R870 B.n172 B.n171 10.6151
R871 B.n172 B.n89 10.6151
R872 B.n176 B.n89 10.6151
R873 B.n179 B.n178 10.6151
R874 B.n179 B.n85 10.6151
R875 B.n183 B.n85 10.6151
R876 B.n184 B.n183 10.6151
R877 B.n185 B.n184 10.6151
R878 B.n185 B.n83 10.6151
R879 B.n189 B.n83 10.6151
R880 B.n190 B.n189 10.6151
R881 B.n192 B.n79 10.6151
R882 B.n196 B.n79 10.6151
R883 B.n197 B.n196 10.6151
R884 B.n198 B.n197 10.6151
R885 B.n198 B.n77 10.6151
R886 B.n202 B.n77 10.6151
R887 B.n203 B.n202 10.6151
R888 B.n204 B.n203 10.6151
R889 B.n204 B.n75 10.6151
R890 B.n208 B.n75 10.6151
R891 B.n209 B.n208 10.6151
R892 B.n210 B.n209 10.6151
R893 B.n210 B.n73 10.6151
R894 B.n413 B.n0 8.11757
R895 B.n413 B.n1 8.11757
R896 B.n343 B.n28 6.5566
R897 B.n331 B.n330 6.5566
R898 B.n178 B.n177 6.5566
R899 B.n191 B.n190 6.5566
R900 B.n28 B.n24 4.05904
R901 B.n330 B.n329 4.05904
R902 B.n177 B.n176 4.05904
R903 B.n192 B.n191 4.05904
C0 VDD2 w_n2578_n1456# 1.43319f
C1 VDD2 VP 0.386026f
C2 w_n2578_n1456# VP 4.80517f
C3 VDD1 VN 0.155375f
C4 VTAIL VDD2 3.74685f
C5 B VN 0.85625f
C6 VTAIL w_n2578_n1456# 1.4798f
C7 B VDD1 1.10967f
C8 VTAIL VP 2.04961f
C9 VN VDD2 1.53403f
C10 VDD1 VDD2 1.07198f
C11 VN w_n2578_n1456# 4.47778f
C12 VN VP 4.26867f
C13 VDD1 w_n2578_n1456# 1.37826f
C14 VDD1 VP 1.76253f
C15 B VDD2 1.16198f
C16 B w_n2578_n1456# 5.73915f
C17 B VP 1.40322f
C18 VTAIL VN 2.03545f
C19 VTAIL VDD1 3.70026f
C20 B VTAIL 1.24627f
C21 VDD2 VSUBS 0.859204f
C22 VDD1 VSUBS 1.042151f
C23 VTAIL VSUBS 0.442702f
C24 VN VSUBS 4.48067f
C25 VP VSUBS 1.690943f
C26 B VSUBS 2.762212f
C27 w_n2578_n1456# VSUBS 47.7342f
C28 B.n0 VSUBS 0.007301f
C29 B.n1 VSUBS 0.007301f
C30 B.n2 VSUBS 0.010798f
C31 B.n3 VSUBS 0.008274f
C32 B.n4 VSUBS 0.008274f
C33 B.n5 VSUBS 0.008274f
C34 B.n6 VSUBS 0.008274f
C35 B.n7 VSUBS 0.008274f
C36 B.n8 VSUBS 0.008274f
C37 B.n9 VSUBS 0.008274f
C38 B.n10 VSUBS 0.008274f
C39 B.n11 VSUBS 0.008274f
C40 B.n12 VSUBS 0.008274f
C41 B.n13 VSUBS 0.008274f
C42 B.n14 VSUBS 0.008274f
C43 B.n15 VSUBS 0.008274f
C44 B.n16 VSUBS 0.008274f
C45 B.n17 VSUBS 0.01863f
C46 B.n18 VSUBS 0.008274f
C47 B.n19 VSUBS 0.008274f
C48 B.n20 VSUBS 0.008274f
C49 B.n21 VSUBS 0.008274f
C50 B.n22 VSUBS 0.008274f
C51 B.n23 VSUBS 0.008274f
C52 B.n24 VSUBS 0.005719f
C53 B.n25 VSUBS 0.008274f
C54 B.t7 VSUBS 0.044609f
C55 B.t8 VSUBS 0.056158f
C56 B.t6 VSUBS 0.234587f
C57 B.n26 VSUBS 0.100971f
C58 B.n27 VSUBS 0.089443f
C59 B.n28 VSUBS 0.019171f
C60 B.n29 VSUBS 0.008274f
C61 B.n30 VSUBS 0.008274f
C62 B.n31 VSUBS 0.008274f
C63 B.n32 VSUBS 0.008274f
C64 B.t1 VSUBS 0.044609f
C65 B.t2 VSUBS 0.056158f
C66 B.t0 VSUBS 0.234587f
C67 B.n33 VSUBS 0.100971f
C68 B.n34 VSUBS 0.089443f
C69 B.n35 VSUBS 0.008274f
C70 B.n36 VSUBS 0.008274f
C71 B.n37 VSUBS 0.008274f
C72 B.n38 VSUBS 0.008274f
C73 B.n39 VSUBS 0.008274f
C74 B.n40 VSUBS 0.008274f
C75 B.n41 VSUBS 0.01863f
C76 B.n42 VSUBS 0.008274f
C77 B.n43 VSUBS 0.008274f
C78 B.n44 VSUBS 0.008274f
C79 B.n45 VSUBS 0.008274f
C80 B.n46 VSUBS 0.008274f
C81 B.n47 VSUBS 0.008274f
C82 B.n48 VSUBS 0.008274f
C83 B.n49 VSUBS 0.008274f
C84 B.n50 VSUBS 0.008274f
C85 B.n51 VSUBS 0.008274f
C86 B.n52 VSUBS 0.008274f
C87 B.n53 VSUBS 0.008274f
C88 B.n54 VSUBS 0.008274f
C89 B.n55 VSUBS 0.008274f
C90 B.n56 VSUBS 0.008274f
C91 B.n57 VSUBS 0.008274f
C92 B.n58 VSUBS 0.008274f
C93 B.n59 VSUBS 0.008274f
C94 B.n60 VSUBS 0.008274f
C95 B.n61 VSUBS 0.008274f
C96 B.n62 VSUBS 0.008274f
C97 B.n63 VSUBS 0.008274f
C98 B.n64 VSUBS 0.008274f
C99 B.n65 VSUBS 0.008274f
C100 B.n66 VSUBS 0.008274f
C101 B.n67 VSUBS 0.008274f
C102 B.n68 VSUBS 0.008274f
C103 B.n69 VSUBS 0.008274f
C104 B.n70 VSUBS 0.008274f
C105 B.n71 VSUBS 0.008274f
C106 B.n72 VSUBS 0.008274f
C107 B.n73 VSUBS 0.019339f
C108 B.n74 VSUBS 0.008274f
C109 B.n75 VSUBS 0.008274f
C110 B.n76 VSUBS 0.008274f
C111 B.n77 VSUBS 0.008274f
C112 B.n78 VSUBS 0.008274f
C113 B.n79 VSUBS 0.008274f
C114 B.n80 VSUBS 0.008274f
C115 B.t11 VSUBS 0.044609f
C116 B.t10 VSUBS 0.056158f
C117 B.t9 VSUBS 0.234587f
C118 B.n81 VSUBS 0.100971f
C119 B.n82 VSUBS 0.089443f
C120 B.n83 VSUBS 0.008274f
C121 B.n84 VSUBS 0.008274f
C122 B.n85 VSUBS 0.008274f
C123 B.n86 VSUBS 0.008274f
C124 B.t5 VSUBS 0.044609f
C125 B.t4 VSUBS 0.056158f
C126 B.t3 VSUBS 0.234587f
C127 B.n87 VSUBS 0.100971f
C128 B.n88 VSUBS 0.089443f
C129 B.n89 VSUBS 0.008274f
C130 B.n90 VSUBS 0.008274f
C131 B.n91 VSUBS 0.008274f
C132 B.n92 VSUBS 0.008274f
C133 B.n93 VSUBS 0.008274f
C134 B.n94 VSUBS 0.008274f
C135 B.n95 VSUBS 0.020309f
C136 B.n96 VSUBS 0.008274f
C137 B.n97 VSUBS 0.008274f
C138 B.n98 VSUBS 0.008274f
C139 B.n99 VSUBS 0.008274f
C140 B.n100 VSUBS 0.008274f
C141 B.n101 VSUBS 0.008274f
C142 B.n102 VSUBS 0.008274f
C143 B.n103 VSUBS 0.008274f
C144 B.n104 VSUBS 0.008274f
C145 B.n105 VSUBS 0.008274f
C146 B.n106 VSUBS 0.008274f
C147 B.n107 VSUBS 0.008274f
C148 B.n108 VSUBS 0.008274f
C149 B.n109 VSUBS 0.008274f
C150 B.n110 VSUBS 0.008274f
C151 B.n111 VSUBS 0.008274f
C152 B.n112 VSUBS 0.008274f
C153 B.n113 VSUBS 0.008274f
C154 B.n114 VSUBS 0.008274f
C155 B.n115 VSUBS 0.008274f
C156 B.n116 VSUBS 0.008274f
C157 B.n117 VSUBS 0.008274f
C158 B.n118 VSUBS 0.008274f
C159 B.n119 VSUBS 0.008274f
C160 B.n120 VSUBS 0.008274f
C161 B.n121 VSUBS 0.008274f
C162 B.n122 VSUBS 0.008274f
C163 B.n123 VSUBS 0.008274f
C164 B.n124 VSUBS 0.008274f
C165 B.n125 VSUBS 0.008274f
C166 B.n126 VSUBS 0.008274f
C167 B.n127 VSUBS 0.008274f
C168 B.n128 VSUBS 0.008274f
C169 B.n129 VSUBS 0.008274f
C170 B.n130 VSUBS 0.008274f
C171 B.n131 VSUBS 0.008274f
C172 B.n132 VSUBS 0.008274f
C173 B.n133 VSUBS 0.008274f
C174 B.n134 VSUBS 0.008274f
C175 B.n135 VSUBS 0.008274f
C176 B.n136 VSUBS 0.008274f
C177 B.n137 VSUBS 0.008274f
C178 B.n138 VSUBS 0.008274f
C179 B.n139 VSUBS 0.008274f
C180 B.n140 VSUBS 0.008274f
C181 B.n141 VSUBS 0.008274f
C182 B.n142 VSUBS 0.008274f
C183 B.n143 VSUBS 0.008274f
C184 B.n144 VSUBS 0.008274f
C185 B.n145 VSUBS 0.008274f
C186 B.n146 VSUBS 0.008274f
C187 B.n147 VSUBS 0.008274f
C188 B.n148 VSUBS 0.008274f
C189 B.n149 VSUBS 0.008274f
C190 B.n150 VSUBS 0.008274f
C191 B.n151 VSUBS 0.008274f
C192 B.n152 VSUBS 0.008274f
C193 B.n153 VSUBS 0.008274f
C194 B.n154 VSUBS 0.01863f
C195 B.n155 VSUBS 0.01863f
C196 B.n156 VSUBS 0.020309f
C197 B.n157 VSUBS 0.008274f
C198 B.n158 VSUBS 0.008274f
C199 B.n159 VSUBS 0.008274f
C200 B.n160 VSUBS 0.008274f
C201 B.n161 VSUBS 0.008274f
C202 B.n162 VSUBS 0.008274f
C203 B.n163 VSUBS 0.008274f
C204 B.n164 VSUBS 0.008274f
C205 B.n165 VSUBS 0.008274f
C206 B.n166 VSUBS 0.008274f
C207 B.n167 VSUBS 0.008274f
C208 B.n168 VSUBS 0.008274f
C209 B.n169 VSUBS 0.008274f
C210 B.n170 VSUBS 0.008274f
C211 B.n171 VSUBS 0.008274f
C212 B.n172 VSUBS 0.008274f
C213 B.n173 VSUBS 0.008274f
C214 B.n174 VSUBS 0.008274f
C215 B.n175 VSUBS 0.008274f
C216 B.n176 VSUBS 0.005719f
C217 B.n177 VSUBS 0.019171f
C218 B.n178 VSUBS 0.006692f
C219 B.n179 VSUBS 0.008274f
C220 B.n180 VSUBS 0.008274f
C221 B.n181 VSUBS 0.008274f
C222 B.n182 VSUBS 0.008274f
C223 B.n183 VSUBS 0.008274f
C224 B.n184 VSUBS 0.008274f
C225 B.n185 VSUBS 0.008274f
C226 B.n186 VSUBS 0.008274f
C227 B.n187 VSUBS 0.008274f
C228 B.n188 VSUBS 0.008274f
C229 B.n189 VSUBS 0.008274f
C230 B.n190 VSUBS 0.006692f
C231 B.n191 VSUBS 0.019171f
C232 B.n192 VSUBS 0.005719f
C233 B.n193 VSUBS 0.008274f
C234 B.n194 VSUBS 0.008274f
C235 B.n195 VSUBS 0.008274f
C236 B.n196 VSUBS 0.008274f
C237 B.n197 VSUBS 0.008274f
C238 B.n198 VSUBS 0.008274f
C239 B.n199 VSUBS 0.008274f
C240 B.n200 VSUBS 0.008274f
C241 B.n201 VSUBS 0.008274f
C242 B.n202 VSUBS 0.008274f
C243 B.n203 VSUBS 0.008274f
C244 B.n204 VSUBS 0.008274f
C245 B.n205 VSUBS 0.008274f
C246 B.n206 VSUBS 0.008274f
C247 B.n207 VSUBS 0.008274f
C248 B.n208 VSUBS 0.008274f
C249 B.n209 VSUBS 0.008274f
C250 B.n210 VSUBS 0.008274f
C251 B.n211 VSUBS 0.008274f
C252 B.n212 VSUBS 0.020309f
C253 B.n213 VSUBS 0.01863f
C254 B.n214 VSUBS 0.019599f
C255 B.n215 VSUBS 0.008274f
C256 B.n216 VSUBS 0.008274f
C257 B.n217 VSUBS 0.008274f
C258 B.n218 VSUBS 0.008274f
C259 B.n219 VSUBS 0.008274f
C260 B.n220 VSUBS 0.008274f
C261 B.n221 VSUBS 0.008274f
C262 B.n222 VSUBS 0.008274f
C263 B.n223 VSUBS 0.008274f
C264 B.n224 VSUBS 0.008274f
C265 B.n225 VSUBS 0.008274f
C266 B.n226 VSUBS 0.008274f
C267 B.n227 VSUBS 0.008274f
C268 B.n228 VSUBS 0.008274f
C269 B.n229 VSUBS 0.008274f
C270 B.n230 VSUBS 0.008274f
C271 B.n231 VSUBS 0.008274f
C272 B.n232 VSUBS 0.008274f
C273 B.n233 VSUBS 0.008274f
C274 B.n234 VSUBS 0.008274f
C275 B.n235 VSUBS 0.008274f
C276 B.n236 VSUBS 0.008274f
C277 B.n237 VSUBS 0.008274f
C278 B.n238 VSUBS 0.008274f
C279 B.n239 VSUBS 0.008274f
C280 B.n240 VSUBS 0.008274f
C281 B.n241 VSUBS 0.008274f
C282 B.n242 VSUBS 0.008274f
C283 B.n243 VSUBS 0.008274f
C284 B.n244 VSUBS 0.008274f
C285 B.n245 VSUBS 0.008274f
C286 B.n246 VSUBS 0.008274f
C287 B.n247 VSUBS 0.008274f
C288 B.n248 VSUBS 0.008274f
C289 B.n249 VSUBS 0.008274f
C290 B.n250 VSUBS 0.008274f
C291 B.n251 VSUBS 0.008274f
C292 B.n252 VSUBS 0.008274f
C293 B.n253 VSUBS 0.008274f
C294 B.n254 VSUBS 0.008274f
C295 B.n255 VSUBS 0.008274f
C296 B.n256 VSUBS 0.008274f
C297 B.n257 VSUBS 0.008274f
C298 B.n258 VSUBS 0.008274f
C299 B.n259 VSUBS 0.008274f
C300 B.n260 VSUBS 0.008274f
C301 B.n261 VSUBS 0.008274f
C302 B.n262 VSUBS 0.008274f
C303 B.n263 VSUBS 0.008274f
C304 B.n264 VSUBS 0.008274f
C305 B.n265 VSUBS 0.008274f
C306 B.n266 VSUBS 0.008274f
C307 B.n267 VSUBS 0.008274f
C308 B.n268 VSUBS 0.008274f
C309 B.n269 VSUBS 0.008274f
C310 B.n270 VSUBS 0.008274f
C311 B.n271 VSUBS 0.008274f
C312 B.n272 VSUBS 0.008274f
C313 B.n273 VSUBS 0.008274f
C314 B.n274 VSUBS 0.008274f
C315 B.n275 VSUBS 0.008274f
C316 B.n276 VSUBS 0.008274f
C317 B.n277 VSUBS 0.008274f
C318 B.n278 VSUBS 0.008274f
C319 B.n279 VSUBS 0.008274f
C320 B.n280 VSUBS 0.008274f
C321 B.n281 VSUBS 0.008274f
C322 B.n282 VSUBS 0.008274f
C323 B.n283 VSUBS 0.008274f
C324 B.n284 VSUBS 0.008274f
C325 B.n285 VSUBS 0.008274f
C326 B.n286 VSUBS 0.008274f
C327 B.n287 VSUBS 0.008274f
C328 B.n288 VSUBS 0.008274f
C329 B.n289 VSUBS 0.008274f
C330 B.n290 VSUBS 0.008274f
C331 B.n291 VSUBS 0.008274f
C332 B.n292 VSUBS 0.008274f
C333 B.n293 VSUBS 0.008274f
C334 B.n294 VSUBS 0.008274f
C335 B.n295 VSUBS 0.008274f
C336 B.n296 VSUBS 0.008274f
C337 B.n297 VSUBS 0.008274f
C338 B.n298 VSUBS 0.008274f
C339 B.n299 VSUBS 0.008274f
C340 B.n300 VSUBS 0.008274f
C341 B.n301 VSUBS 0.008274f
C342 B.n302 VSUBS 0.008274f
C343 B.n303 VSUBS 0.008274f
C344 B.n304 VSUBS 0.008274f
C345 B.n305 VSUBS 0.008274f
C346 B.n306 VSUBS 0.008274f
C347 B.n307 VSUBS 0.008274f
C348 B.n308 VSUBS 0.01863f
C349 B.n309 VSUBS 0.020309f
C350 B.n310 VSUBS 0.020309f
C351 B.n311 VSUBS 0.008274f
C352 B.n312 VSUBS 0.008274f
C353 B.n313 VSUBS 0.008274f
C354 B.n314 VSUBS 0.008274f
C355 B.n315 VSUBS 0.008274f
C356 B.n316 VSUBS 0.008274f
C357 B.n317 VSUBS 0.008274f
C358 B.n318 VSUBS 0.008274f
C359 B.n319 VSUBS 0.008274f
C360 B.n320 VSUBS 0.008274f
C361 B.n321 VSUBS 0.008274f
C362 B.n322 VSUBS 0.008274f
C363 B.n323 VSUBS 0.008274f
C364 B.n324 VSUBS 0.008274f
C365 B.n325 VSUBS 0.008274f
C366 B.n326 VSUBS 0.008274f
C367 B.n327 VSUBS 0.008274f
C368 B.n328 VSUBS 0.008274f
C369 B.n329 VSUBS 0.005719f
C370 B.n330 VSUBS 0.019171f
C371 B.n331 VSUBS 0.006692f
C372 B.n332 VSUBS 0.008274f
C373 B.n333 VSUBS 0.008274f
C374 B.n334 VSUBS 0.008274f
C375 B.n335 VSUBS 0.008274f
C376 B.n336 VSUBS 0.008274f
C377 B.n337 VSUBS 0.008274f
C378 B.n338 VSUBS 0.008274f
C379 B.n339 VSUBS 0.008274f
C380 B.n340 VSUBS 0.008274f
C381 B.n341 VSUBS 0.008274f
C382 B.n342 VSUBS 0.008274f
C383 B.n343 VSUBS 0.006692f
C384 B.n344 VSUBS 0.008274f
C385 B.n345 VSUBS 0.008274f
C386 B.n346 VSUBS 0.008274f
C387 B.n347 VSUBS 0.008274f
C388 B.n348 VSUBS 0.008274f
C389 B.n349 VSUBS 0.008274f
C390 B.n350 VSUBS 0.008274f
C391 B.n351 VSUBS 0.008274f
C392 B.n352 VSUBS 0.008274f
C393 B.n353 VSUBS 0.008274f
C394 B.n354 VSUBS 0.008274f
C395 B.n355 VSUBS 0.008274f
C396 B.n356 VSUBS 0.008274f
C397 B.n357 VSUBS 0.008274f
C398 B.n358 VSUBS 0.008274f
C399 B.n359 VSUBS 0.008274f
C400 B.n360 VSUBS 0.008274f
C401 B.n361 VSUBS 0.008274f
C402 B.n362 VSUBS 0.008274f
C403 B.n363 VSUBS 0.008274f
C404 B.n364 VSUBS 0.020309f
C405 B.n365 VSUBS 0.020309f
C406 B.n366 VSUBS 0.01863f
C407 B.n367 VSUBS 0.008274f
C408 B.n368 VSUBS 0.008274f
C409 B.n369 VSUBS 0.008274f
C410 B.n370 VSUBS 0.008274f
C411 B.n371 VSUBS 0.008274f
C412 B.n372 VSUBS 0.008274f
C413 B.n373 VSUBS 0.008274f
C414 B.n374 VSUBS 0.008274f
C415 B.n375 VSUBS 0.008274f
C416 B.n376 VSUBS 0.008274f
C417 B.n377 VSUBS 0.008274f
C418 B.n378 VSUBS 0.008274f
C419 B.n379 VSUBS 0.008274f
C420 B.n380 VSUBS 0.008274f
C421 B.n381 VSUBS 0.008274f
C422 B.n382 VSUBS 0.008274f
C423 B.n383 VSUBS 0.008274f
C424 B.n384 VSUBS 0.008274f
C425 B.n385 VSUBS 0.008274f
C426 B.n386 VSUBS 0.008274f
C427 B.n387 VSUBS 0.008274f
C428 B.n388 VSUBS 0.008274f
C429 B.n389 VSUBS 0.008274f
C430 B.n390 VSUBS 0.008274f
C431 B.n391 VSUBS 0.008274f
C432 B.n392 VSUBS 0.008274f
C433 B.n393 VSUBS 0.008274f
C434 B.n394 VSUBS 0.008274f
C435 B.n395 VSUBS 0.008274f
C436 B.n396 VSUBS 0.008274f
C437 B.n397 VSUBS 0.008274f
C438 B.n398 VSUBS 0.008274f
C439 B.n399 VSUBS 0.008274f
C440 B.n400 VSUBS 0.008274f
C441 B.n401 VSUBS 0.008274f
C442 B.n402 VSUBS 0.008274f
C443 B.n403 VSUBS 0.008274f
C444 B.n404 VSUBS 0.008274f
C445 B.n405 VSUBS 0.008274f
C446 B.n406 VSUBS 0.008274f
C447 B.n407 VSUBS 0.008274f
C448 B.n408 VSUBS 0.008274f
C449 B.n409 VSUBS 0.008274f
C450 B.n410 VSUBS 0.008274f
C451 B.n411 VSUBS 0.010798f
C452 B.n412 VSUBS 0.011502f
C453 B.n413 VSUBS 0.022873f
C454 VDD1.n0 VSUBS 0.015982f
C455 VDD1.n1 VSUBS 0.107022f
C456 VDD1.n2 VSUBS 0.008364f
C457 VDD1.t2 VSUBS 0.043384f
C458 VDD1.n3 VSUBS 0.050762f
C459 VDD1.n4 VSUBS 0.011657f
C460 VDD1.n5 VSUBS 0.014827f
C461 VDD1.n6 VSUBS 0.044041f
C462 VDD1.n7 VSUBS 0.008856f
C463 VDD1.n8 VSUBS 0.008364f
C464 VDD1.n9 VSUBS 0.036828f
C465 VDD1.n10 VSUBS 0.035369f
C466 VDD1.n11 VSUBS 0.015982f
C467 VDD1.n12 VSUBS 0.107022f
C468 VDD1.n13 VSUBS 0.008364f
C469 VDD1.t4 VSUBS 0.043384f
C470 VDD1.n14 VSUBS 0.050762f
C471 VDD1.n15 VSUBS 0.011657f
C472 VDD1.n16 VSUBS 0.014827f
C473 VDD1.n17 VSUBS 0.044041f
C474 VDD1.n18 VSUBS 0.008856f
C475 VDD1.n19 VSUBS 0.008364f
C476 VDD1.n20 VSUBS 0.036828f
C477 VDD1.n21 VSUBS 0.035023f
C478 VDD1.t3 VSUBS 0.030011f
C479 VDD1.t5 VSUBS 0.030011f
C480 VDD1.n22 VSUBS 0.146551f
C481 VDD1.n23 VSUBS 1.17758f
C482 VDD1.t1 VSUBS 0.030011f
C483 VDD1.t0 VSUBS 0.030011f
C484 VDD1.n24 VSUBS 0.145828f
C485 VDD1.n25 VSUBS 1.15659f
C486 VP.n0 VSUBS 0.052599f
C487 VP.t0 VSUBS 0.521699f
C488 VP.n1 VSUBS 0.042499f
C489 VP.n2 VSUBS 0.052599f
C490 VP.t2 VSUBS 0.521699f
C491 VP.n3 VSUBS 0.042499f
C492 VP.n4 VSUBS 0.052599f
C493 VP.t1 VSUBS 0.521699f
C494 VP.n5 VSUBS 0.052599f
C495 VP.t5 VSUBS 0.521699f
C496 VP.n6 VSUBS 0.042499f
C497 VP.t3 VSUBS 0.75499f
C498 VP.n7 VSUBS 0.340385f
C499 VP.t4 VSUBS 0.521699f
C500 VP.n8 VSUBS 0.386708f
C501 VP.n9 VSUBS 0.104241f
C502 VP.n10 VSUBS 0.379462f
C503 VP.n11 VSUBS 0.052599f
C504 VP.n12 VSUBS 0.052599f
C505 VP.n13 VSUBS 0.10372f
C506 VP.n14 VSUBS 0.05035f
C507 VP.n15 VSUBS 0.350348f
C508 VP.n16 VSUBS 1.81092f
C509 VP.n17 VSUBS 1.86129f
C510 VP.n18 VSUBS 0.350348f
C511 VP.n19 VSUBS 0.05035f
C512 VP.n20 VSUBS 0.10372f
C513 VP.n21 VSUBS 0.052599f
C514 VP.n22 VSUBS 0.052599f
C515 VP.n23 VSUBS 0.052599f
C516 VP.n24 VSUBS 0.104241f
C517 VP.n25 VSUBS 0.298955f
C518 VP.n26 VSUBS 0.104241f
C519 VP.n27 VSUBS 0.052599f
C520 VP.n28 VSUBS 0.052599f
C521 VP.n29 VSUBS 0.052599f
C522 VP.n30 VSUBS 0.10372f
C523 VP.n31 VSUBS 0.05035f
C524 VP.n32 VSUBS 0.350348f
C525 VP.n33 VSUBS 0.055819f
C526 VDD2.n0 VSUBS 0.016234f
C527 VDD2.n1 VSUBS 0.108711f
C528 VDD2.n2 VSUBS 0.008496f
C529 VDD2.t5 VSUBS 0.044068f
C530 VDD2.n3 VSUBS 0.051563f
C531 VDD2.n4 VSUBS 0.01184f
C532 VDD2.n5 VSUBS 0.015061f
C533 VDD2.n6 VSUBS 0.044736f
C534 VDD2.n7 VSUBS 0.008996f
C535 VDD2.n8 VSUBS 0.008496f
C536 VDD2.n9 VSUBS 0.037409f
C537 VDD2.n10 VSUBS 0.035575f
C538 VDD2.t2 VSUBS 0.030485f
C539 VDD2.t4 VSUBS 0.030485f
C540 VDD2.n11 VSUBS 0.148864f
C541 VDD2.n12 VSUBS 1.13754f
C542 VDD2.n13 VSUBS 0.016234f
C543 VDD2.n14 VSUBS 0.108711f
C544 VDD2.n15 VSUBS 0.008496f
C545 VDD2.t0 VSUBS 0.044068f
C546 VDD2.n16 VSUBS 0.051563f
C547 VDD2.n17 VSUBS 0.01184f
C548 VDD2.n18 VSUBS 0.015061f
C549 VDD2.n19 VSUBS 0.044736f
C550 VDD2.n20 VSUBS 0.008996f
C551 VDD2.n21 VSUBS 0.008496f
C552 VDD2.n22 VSUBS 0.037409f
C553 VDD2.n23 VSUBS 0.033262f
C554 VDD2.n24 VSUBS 0.979274f
C555 VDD2.t1 VSUBS 0.030485f
C556 VDD2.t3 VSUBS 0.030485f
C557 VDD2.n25 VSUBS 0.148856f
C558 VTAIL.t10 VSUBS 0.05948f
C559 VTAIL.t9 VSUBS 0.05948f
C560 VTAIL.n0 VSUBS 0.246091f
C561 VTAIL.n1 VSUBS 0.5381f
C562 VTAIL.n2 VSUBS 0.031674f
C563 VTAIL.n3 VSUBS 0.212109f
C564 VTAIL.n4 VSUBS 0.016576f
C565 VTAIL.t5 VSUBS 0.085982f
C566 VTAIL.n5 VSUBS 0.100605f
C567 VTAIL.n6 VSUBS 0.023102f
C568 VTAIL.n7 VSUBS 0.029386f
C569 VTAIL.n8 VSUBS 0.087286f
C570 VTAIL.n9 VSUBS 0.017552f
C571 VTAIL.n10 VSUBS 0.016576f
C572 VTAIL.n11 VSUBS 0.07299f
C573 VTAIL.n12 VSUBS 0.043611f
C574 VTAIL.n13 VSUBS 0.332353f
C575 VTAIL.t2 VSUBS 0.05948f
C576 VTAIL.t3 VSUBS 0.05948f
C577 VTAIL.n14 VSUBS 0.246091f
C578 VTAIL.n15 VSUBS 1.50126f
C579 VTAIL.t6 VSUBS 0.05948f
C580 VTAIL.t8 VSUBS 0.05948f
C581 VTAIL.n16 VSUBS 0.246092f
C582 VTAIL.n17 VSUBS 1.50126f
C583 VTAIL.n18 VSUBS 0.031674f
C584 VTAIL.n19 VSUBS 0.212109f
C585 VTAIL.n20 VSUBS 0.016576f
C586 VTAIL.t11 VSUBS 0.085982f
C587 VTAIL.n21 VSUBS 0.100605f
C588 VTAIL.n22 VSUBS 0.023102f
C589 VTAIL.n23 VSUBS 0.029386f
C590 VTAIL.n24 VSUBS 0.087286f
C591 VTAIL.n25 VSUBS 0.017552f
C592 VTAIL.n26 VSUBS 0.016576f
C593 VTAIL.n27 VSUBS 0.07299f
C594 VTAIL.n28 VSUBS 0.043611f
C595 VTAIL.n29 VSUBS 0.332353f
C596 VTAIL.t4 VSUBS 0.05948f
C597 VTAIL.t0 VSUBS 0.05948f
C598 VTAIL.n30 VSUBS 0.246092f
C599 VTAIL.n31 VSUBS 0.661491f
C600 VTAIL.n32 VSUBS 0.031674f
C601 VTAIL.n33 VSUBS 0.212109f
C602 VTAIL.n34 VSUBS 0.016576f
C603 VTAIL.t1 VSUBS 0.085982f
C604 VTAIL.n35 VSUBS 0.100605f
C605 VTAIL.n36 VSUBS 0.023102f
C606 VTAIL.n37 VSUBS 0.029386f
C607 VTAIL.n38 VSUBS 0.087286f
C608 VTAIL.n39 VSUBS 0.017552f
C609 VTAIL.n40 VSUBS 0.016576f
C610 VTAIL.n41 VSUBS 0.07299f
C611 VTAIL.n42 VSUBS 0.043611f
C612 VTAIL.n43 VSUBS 0.999888f
C613 VTAIL.n44 VSUBS 0.031674f
C614 VTAIL.n45 VSUBS 0.212109f
C615 VTAIL.n46 VSUBS 0.016576f
C616 VTAIL.t7 VSUBS 0.085982f
C617 VTAIL.n47 VSUBS 0.100605f
C618 VTAIL.n48 VSUBS 0.023102f
C619 VTAIL.n49 VSUBS 0.029386f
C620 VTAIL.n50 VSUBS 0.087286f
C621 VTAIL.n51 VSUBS 0.017552f
C622 VTAIL.n52 VSUBS 0.016576f
C623 VTAIL.n53 VSUBS 0.07299f
C624 VTAIL.n54 VSUBS 0.043611f
C625 VTAIL.n55 VSUBS 0.951045f
C626 VN.n0 VSUBS 0.050838f
C627 VN.t1 VSUBS 0.50424f
C628 VN.n1 VSUBS 0.041077f
C629 VN.t0 VSUBS 0.729724f
C630 VN.n2 VSUBS 0.328994f
C631 VN.t3 VSUBS 0.50424f
C632 VN.n3 VSUBS 0.373766f
C633 VN.n4 VSUBS 0.100753f
C634 VN.n5 VSUBS 0.366764f
C635 VN.n6 VSUBS 0.050838f
C636 VN.n7 VSUBS 0.050838f
C637 VN.n8 VSUBS 0.100249f
C638 VN.n9 VSUBS 0.048665f
C639 VN.n10 VSUBS 0.338623f
C640 VN.n11 VSUBS 0.053951f
C641 VN.n12 VSUBS 0.050838f
C642 VN.t5 VSUBS 0.50424f
C643 VN.n13 VSUBS 0.041077f
C644 VN.t2 VSUBS 0.729724f
C645 VN.n14 VSUBS 0.328994f
C646 VN.t4 VSUBS 0.50424f
C647 VN.n15 VSUBS 0.373766f
C648 VN.n16 VSUBS 0.100753f
C649 VN.n17 VSUBS 0.366764f
C650 VN.n18 VSUBS 0.050838f
C651 VN.n19 VSUBS 0.050838f
C652 VN.n20 VSUBS 0.100249f
C653 VN.n21 VSUBS 0.048665f
C654 VN.n22 VSUBS 0.338623f
C655 VN.n23 VSUBS 1.78393f
.ends

