* NGSPICE file created from diff_pair_sample_0688.ext - technology: sky130A

.subckt diff_pair_sample_0688 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0 ps=0 w=1.42 l=1.22
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0.5538 ps=3.62 w=1.42 l=1.22
X2 VDD1.t0 VP.t1 VTAIL.t2 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0.5538 ps=3.62 w=1.42 l=1.22
X3 VDD2.t1 VN.t0 VTAIL.t1 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0.5538 ps=3.62 w=1.42 l=1.22
X4 B.t8 B.t6 B.t7 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0 ps=0 w=1.42 l=1.22
X5 VDD2.t0 VN.t1 VTAIL.t0 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0.5538 ps=3.62 w=1.42 l=1.22
X6 B.t5 B.t3 B.t4 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0 ps=0 w=1.42 l=1.22
X7 B.t2 B.t0 B.t1 w_n1590_n1252# sky130_fd_pr__pfet_01v8 ad=0.5538 pd=3.62 as=0 ps=0 w=1.42 l=1.22
R0 B.n201 B.n30 585
R1 B.n203 B.n202 585
R2 B.n204 B.n29 585
R3 B.n206 B.n205 585
R4 B.n207 B.n28 585
R5 B.n209 B.n208 585
R6 B.n210 B.n27 585
R7 B.n212 B.n211 585
R8 B.n213 B.n26 585
R9 B.n215 B.n214 585
R10 B.n216 B.n23 585
R11 B.n219 B.n218 585
R12 B.n220 B.n22 585
R13 B.n222 B.n221 585
R14 B.n223 B.n21 585
R15 B.n225 B.n224 585
R16 B.n226 B.n20 585
R17 B.n228 B.n227 585
R18 B.n229 B.n19 585
R19 B.n231 B.n230 585
R20 B.n233 B.n232 585
R21 B.n234 B.n15 585
R22 B.n236 B.n235 585
R23 B.n237 B.n14 585
R24 B.n239 B.n238 585
R25 B.n240 B.n13 585
R26 B.n242 B.n241 585
R27 B.n243 B.n12 585
R28 B.n245 B.n244 585
R29 B.n246 B.n11 585
R30 B.n248 B.n247 585
R31 B.n200 B.n199 585
R32 B.n198 B.n31 585
R33 B.n197 B.n196 585
R34 B.n195 B.n32 585
R35 B.n194 B.n193 585
R36 B.n192 B.n33 585
R37 B.n191 B.n190 585
R38 B.n189 B.n34 585
R39 B.n188 B.n187 585
R40 B.n186 B.n35 585
R41 B.n185 B.n184 585
R42 B.n183 B.n36 585
R43 B.n182 B.n181 585
R44 B.n180 B.n37 585
R45 B.n179 B.n178 585
R46 B.n177 B.n38 585
R47 B.n176 B.n175 585
R48 B.n174 B.n39 585
R49 B.n173 B.n172 585
R50 B.n171 B.n40 585
R51 B.n170 B.n169 585
R52 B.n168 B.n41 585
R53 B.n167 B.n166 585
R54 B.n165 B.n42 585
R55 B.n164 B.n163 585
R56 B.n162 B.n43 585
R57 B.n161 B.n160 585
R58 B.n159 B.n44 585
R59 B.n158 B.n157 585
R60 B.n156 B.n45 585
R61 B.n155 B.n154 585
R62 B.n153 B.n46 585
R63 B.n152 B.n151 585
R64 B.n150 B.n47 585
R65 B.n149 B.n148 585
R66 B.n101 B.n100 585
R67 B.n102 B.n67 585
R68 B.n104 B.n103 585
R69 B.n105 B.n66 585
R70 B.n107 B.n106 585
R71 B.n108 B.n65 585
R72 B.n110 B.n109 585
R73 B.n111 B.n64 585
R74 B.n113 B.n112 585
R75 B.n114 B.n63 585
R76 B.n116 B.n115 585
R77 B.n118 B.n117 585
R78 B.n119 B.n59 585
R79 B.n121 B.n120 585
R80 B.n122 B.n58 585
R81 B.n124 B.n123 585
R82 B.n125 B.n57 585
R83 B.n127 B.n126 585
R84 B.n128 B.n56 585
R85 B.n130 B.n129 585
R86 B.n132 B.n53 585
R87 B.n134 B.n133 585
R88 B.n135 B.n52 585
R89 B.n137 B.n136 585
R90 B.n138 B.n51 585
R91 B.n140 B.n139 585
R92 B.n141 B.n50 585
R93 B.n143 B.n142 585
R94 B.n144 B.n49 585
R95 B.n146 B.n145 585
R96 B.n147 B.n48 585
R97 B.n99 B.n68 585
R98 B.n98 B.n97 585
R99 B.n96 B.n69 585
R100 B.n95 B.n94 585
R101 B.n93 B.n70 585
R102 B.n92 B.n91 585
R103 B.n90 B.n71 585
R104 B.n89 B.n88 585
R105 B.n87 B.n72 585
R106 B.n86 B.n85 585
R107 B.n84 B.n73 585
R108 B.n83 B.n82 585
R109 B.n81 B.n74 585
R110 B.n80 B.n79 585
R111 B.n78 B.n75 585
R112 B.n77 B.n76 585
R113 B.n2 B.n0 585
R114 B.n273 B.n1 585
R115 B.n272 B.n271 585
R116 B.n270 B.n3 585
R117 B.n269 B.n268 585
R118 B.n267 B.n4 585
R119 B.n266 B.n265 585
R120 B.n264 B.n5 585
R121 B.n263 B.n262 585
R122 B.n261 B.n6 585
R123 B.n260 B.n259 585
R124 B.n258 B.n7 585
R125 B.n257 B.n256 585
R126 B.n255 B.n8 585
R127 B.n254 B.n253 585
R128 B.n252 B.n9 585
R129 B.n251 B.n250 585
R130 B.n249 B.n10 585
R131 B.n275 B.n274 585
R132 B.n100 B.n99 502.111
R133 B.n249 B.n248 502.111
R134 B.n148 B.n147 502.111
R135 B.n201 B.n200 502.111
R136 B.n54 B.t8 279.178
R137 B.n24 B.t1 279.178
R138 B.n60 B.t5 279.178
R139 B.n16 B.t10 279.178
R140 B.n55 B.t7 249.118
R141 B.n25 B.t2 249.118
R142 B.n61 B.t4 249.117
R143 B.n17 B.t11 249.117
R144 B.n54 B.t6 232.27
R145 B.n60 B.t3 232.27
R146 B.n16 B.t9 232.27
R147 B.n24 B.t0 232.27
R148 B.n99 B.n98 163.367
R149 B.n98 B.n69 163.367
R150 B.n94 B.n69 163.367
R151 B.n94 B.n93 163.367
R152 B.n93 B.n92 163.367
R153 B.n92 B.n71 163.367
R154 B.n88 B.n71 163.367
R155 B.n88 B.n87 163.367
R156 B.n87 B.n86 163.367
R157 B.n86 B.n73 163.367
R158 B.n82 B.n73 163.367
R159 B.n82 B.n81 163.367
R160 B.n81 B.n80 163.367
R161 B.n80 B.n75 163.367
R162 B.n76 B.n75 163.367
R163 B.n76 B.n2 163.367
R164 B.n274 B.n2 163.367
R165 B.n274 B.n273 163.367
R166 B.n273 B.n272 163.367
R167 B.n272 B.n3 163.367
R168 B.n268 B.n3 163.367
R169 B.n268 B.n267 163.367
R170 B.n267 B.n266 163.367
R171 B.n266 B.n5 163.367
R172 B.n262 B.n5 163.367
R173 B.n262 B.n261 163.367
R174 B.n261 B.n260 163.367
R175 B.n260 B.n7 163.367
R176 B.n256 B.n7 163.367
R177 B.n256 B.n255 163.367
R178 B.n255 B.n254 163.367
R179 B.n254 B.n9 163.367
R180 B.n250 B.n9 163.367
R181 B.n250 B.n249 163.367
R182 B.n100 B.n67 163.367
R183 B.n104 B.n67 163.367
R184 B.n105 B.n104 163.367
R185 B.n106 B.n105 163.367
R186 B.n106 B.n65 163.367
R187 B.n110 B.n65 163.367
R188 B.n111 B.n110 163.367
R189 B.n112 B.n111 163.367
R190 B.n112 B.n63 163.367
R191 B.n116 B.n63 163.367
R192 B.n117 B.n116 163.367
R193 B.n117 B.n59 163.367
R194 B.n121 B.n59 163.367
R195 B.n122 B.n121 163.367
R196 B.n123 B.n122 163.367
R197 B.n123 B.n57 163.367
R198 B.n127 B.n57 163.367
R199 B.n128 B.n127 163.367
R200 B.n129 B.n128 163.367
R201 B.n129 B.n53 163.367
R202 B.n134 B.n53 163.367
R203 B.n135 B.n134 163.367
R204 B.n136 B.n135 163.367
R205 B.n136 B.n51 163.367
R206 B.n140 B.n51 163.367
R207 B.n141 B.n140 163.367
R208 B.n142 B.n141 163.367
R209 B.n142 B.n49 163.367
R210 B.n146 B.n49 163.367
R211 B.n147 B.n146 163.367
R212 B.n148 B.n47 163.367
R213 B.n152 B.n47 163.367
R214 B.n153 B.n152 163.367
R215 B.n154 B.n153 163.367
R216 B.n154 B.n45 163.367
R217 B.n158 B.n45 163.367
R218 B.n159 B.n158 163.367
R219 B.n160 B.n159 163.367
R220 B.n160 B.n43 163.367
R221 B.n164 B.n43 163.367
R222 B.n165 B.n164 163.367
R223 B.n166 B.n165 163.367
R224 B.n166 B.n41 163.367
R225 B.n170 B.n41 163.367
R226 B.n171 B.n170 163.367
R227 B.n172 B.n171 163.367
R228 B.n172 B.n39 163.367
R229 B.n176 B.n39 163.367
R230 B.n177 B.n176 163.367
R231 B.n178 B.n177 163.367
R232 B.n178 B.n37 163.367
R233 B.n182 B.n37 163.367
R234 B.n183 B.n182 163.367
R235 B.n184 B.n183 163.367
R236 B.n184 B.n35 163.367
R237 B.n188 B.n35 163.367
R238 B.n189 B.n188 163.367
R239 B.n190 B.n189 163.367
R240 B.n190 B.n33 163.367
R241 B.n194 B.n33 163.367
R242 B.n195 B.n194 163.367
R243 B.n196 B.n195 163.367
R244 B.n196 B.n31 163.367
R245 B.n200 B.n31 163.367
R246 B.n248 B.n11 163.367
R247 B.n244 B.n11 163.367
R248 B.n244 B.n243 163.367
R249 B.n243 B.n242 163.367
R250 B.n242 B.n13 163.367
R251 B.n238 B.n13 163.367
R252 B.n238 B.n237 163.367
R253 B.n237 B.n236 163.367
R254 B.n236 B.n15 163.367
R255 B.n232 B.n15 163.367
R256 B.n232 B.n231 163.367
R257 B.n231 B.n19 163.367
R258 B.n227 B.n19 163.367
R259 B.n227 B.n226 163.367
R260 B.n226 B.n225 163.367
R261 B.n225 B.n21 163.367
R262 B.n221 B.n21 163.367
R263 B.n221 B.n220 163.367
R264 B.n220 B.n219 163.367
R265 B.n219 B.n23 163.367
R266 B.n214 B.n23 163.367
R267 B.n214 B.n213 163.367
R268 B.n213 B.n212 163.367
R269 B.n212 B.n27 163.367
R270 B.n208 B.n27 163.367
R271 B.n208 B.n207 163.367
R272 B.n207 B.n206 163.367
R273 B.n206 B.n29 163.367
R274 B.n202 B.n29 163.367
R275 B.n202 B.n201 163.367
R276 B.n131 B.n55 59.5399
R277 B.n62 B.n61 59.5399
R278 B.n18 B.n17 59.5399
R279 B.n217 B.n25 59.5399
R280 B.n247 B.n10 32.6249
R281 B.n199 B.n30 32.6249
R282 B.n149 B.n48 32.6249
R283 B.n101 B.n68 32.6249
R284 B.n55 B.n54 30.0611
R285 B.n61 B.n60 30.0611
R286 B.n17 B.n16 30.0611
R287 B.n25 B.n24 30.0611
R288 B B.n275 18.0485
R289 B.n247 B.n246 10.6151
R290 B.n246 B.n245 10.6151
R291 B.n245 B.n12 10.6151
R292 B.n241 B.n12 10.6151
R293 B.n241 B.n240 10.6151
R294 B.n240 B.n239 10.6151
R295 B.n239 B.n14 10.6151
R296 B.n235 B.n14 10.6151
R297 B.n235 B.n234 10.6151
R298 B.n234 B.n233 10.6151
R299 B.n230 B.n229 10.6151
R300 B.n229 B.n228 10.6151
R301 B.n228 B.n20 10.6151
R302 B.n224 B.n20 10.6151
R303 B.n224 B.n223 10.6151
R304 B.n223 B.n222 10.6151
R305 B.n222 B.n22 10.6151
R306 B.n218 B.n22 10.6151
R307 B.n216 B.n215 10.6151
R308 B.n215 B.n26 10.6151
R309 B.n211 B.n26 10.6151
R310 B.n211 B.n210 10.6151
R311 B.n210 B.n209 10.6151
R312 B.n209 B.n28 10.6151
R313 B.n205 B.n28 10.6151
R314 B.n205 B.n204 10.6151
R315 B.n204 B.n203 10.6151
R316 B.n203 B.n30 10.6151
R317 B.n150 B.n149 10.6151
R318 B.n151 B.n150 10.6151
R319 B.n151 B.n46 10.6151
R320 B.n155 B.n46 10.6151
R321 B.n156 B.n155 10.6151
R322 B.n157 B.n156 10.6151
R323 B.n157 B.n44 10.6151
R324 B.n161 B.n44 10.6151
R325 B.n162 B.n161 10.6151
R326 B.n163 B.n162 10.6151
R327 B.n163 B.n42 10.6151
R328 B.n167 B.n42 10.6151
R329 B.n168 B.n167 10.6151
R330 B.n169 B.n168 10.6151
R331 B.n169 B.n40 10.6151
R332 B.n173 B.n40 10.6151
R333 B.n174 B.n173 10.6151
R334 B.n175 B.n174 10.6151
R335 B.n175 B.n38 10.6151
R336 B.n179 B.n38 10.6151
R337 B.n180 B.n179 10.6151
R338 B.n181 B.n180 10.6151
R339 B.n181 B.n36 10.6151
R340 B.n185 B.n36 10.6151
R341 B.n186 B.n185 10.6151
R342 B.n187 B.n186 10.6151
R343 B.n187 B.n34 10.6151
R344 B.n191 B.n34 10.6151
R345 B.n192 B.n191 10.6151
R346 B.n193 B.n192 10.6151
R347 B.n193 B.n32 10.6151
R348 B.n197 B.n32 10.6151
R349 B.n198 B.n197 10.6151
R350 B.n199 B.n198 10.6151
R351 B.n102 B.n101 10.6151
R352 B.n103 B.n102 10.6151
R353 B.n103 B.n66 10.6151
R354 B.n107 B.n66 10.6151
R355 B.n108 B.n107 10.6151
R356 B.n109 B.n108 10.6151
R357 B.n109 B.n64 10.6151
R358 B.n113 B.n64 10.6151
R359 B.n114 B.n113 10.6151
R360 B.n115 B.n114 10.6151
R361 B.n119 B.n118 10.6151
R362 B.n120 B.n119 10.6151
R363 B.n120 B.n58 10.6151
R364 B.n124 B.n58 10.6151
R365 B.n125 B.n124 10.6151
R366 B.n126 B.n125 10.6151
R367 B.n126 B.n56 10.6151
R368 B.n130 B.n56 10.6151
R369 B.n133 B.n132 10.6151
R370 B.n133 B.n52 10.6151
R371 B.n137 B.n52 10.6151
R372 B.n138 B.n137 10.6151
R373 B.n139 B.n138 10.6151
R374 B.n139 B.n50 10.6151
R375 B.n143 B.n50 10.6151
R376 B.n144 B.n143 10.6151
R377 B.n145 B.n144 10.6151
R378 B.n145 B.n48 10.6151
R379 B.n97 B.n68 10.6151
R380 B.n97 B.n96 10.6151
R381 B.n96 B.n95 10.6151
R382 B.n95 B.n70 10.6151
R383 B.n91 B.n70 10.6151
R384 B.n91 B.n90 10.6151
R385 B.n90 B.n89 10.6151
R386 B.n89 B.n72 10.6151
R387 B.n85 B.n72 10.6151
R388 B.n85 B.n84 10.6151
R389 B.n84 B.n83 10.6151
R390 B.n83 B.n74 10.6151
R391 B.n79 B.n74 10.6151
R392 B.n79 B.n78 10.6151
R393 B.n78 B.n77 10.6151
R394 B.n77 B.n0 10.6151
R395 B.n271 B.n1 10.6151
R396 B.n271 B.n270 10.6151
R397 B.n270 B.n269 10.6151
R398 B.n269 B.n4 10.6151
R399 B.n265 B.n4 10.6151
R400 B.n265 B.n264 10.6151
R401 B.n264 B.n263 10.6151
R402 B.n263 B.n6 10.6151
R403 B.n259 B.n6 10.6151
R404 B.n259 B.n258 10.6151
R405 B.n258 B.n257 10.6151
R406 B.n257 B.n8 10.6151
R407 B.n253 B.n8 10.6151
R408 B.n253 B.n252 10.6151
R409 B.n252 B.n251 10.6151
R410 B.n251 B.n10 10.6151
R411 B.n230 B.n18 6.5566
R412 B.n218 B.n217 6.5566
R413 B.n118 B.n62 6.5566
R414 B.n131 B.n130 6.5566
R415 B.n233 B.n18 4.05904
R416 B.n217 B.n216 4.05904
R417 B.n115 B.n62 4.05904
R418 B.n132 B.n131 4.05904
R419 B.n275 B.n0 2.81026
R420 B.n275 B.n1 2.81026
R421 VP.n0 VP.t1 173.835
R422 VP.n0 VP.t0 140.853
R423 VP VP.n0 0.146778
R424 VTAIL.n1 VTAIL.t1 255.613
R425 VTAIL.n3 VTAIL.t0 255.613
R426 VTAIL.n0 VTAIL.t3 255.613
R427 VTAIL.n2 VTAIL.t2 255.613
R428 VTAIL.n1 VTAIL.n0 16.2634
R429 VTAIL.n3 VTAIL.n2 14.9272
R430 VTAIL.n2 VTAIL.n1 1.13843
R431 VTAIL VTAIL.n0 0.862569
R432 VTAIL VTAIL.n3 0.276362
R433 VDD1 VDD1.t1 300.707
R434 VDD1 VDD1.t0 272.683
R435 VN VN.t0 174.121
R436 VN VN.t1 141
R437 VDD2.n0 VDD2.t0 299.848
R438 VDD2.n0 VDD2.t1 272.291
R439 VDD2 VDD2.n0 0.392741
C0 VDD2 VN 0.496742f
C1 VP VDD2 0.282375f
C2 B VDD2 0.724981f
C3 w_n1590_n1252# VDD2 0.865125f
C4 VP VN 2.85652f
C5 B VN 0.663322f
C6 B VP 0.984861f
C7 w_n1590_n1252# VN 1.83437f
C8 w_n1590_n1252# VP 2.02752f
C9 w_n1590_n1252# B 4.34531f
C10 VTAIL VDD1 1.84948f
C11 VTAIL VDD2 1.89295f
C12 VDD1 VDD2 0.513188f
C13 VTAIL VN 0.651792f
C14 VDD1 VN 0.155006f
C15 VTAIL VP 0.665942f
C16 VTAIL B 0.867351f
C17 VDD1 VP 0.622523f
C18 B VDD1 0.706405f
C19 VTAIL w_n1590_n1252# 1.11732f
C20 w_n1590_n1252# VDD1 0.856207f
C21 VDD2 VSUBS 0.35768f
C22 VDD1 VSUBS 0.53347f
C23 VTAIL VSUBS 0.208963f
C24 VN VSUBS 3.45685f
C25 VP VSUBS 0.795691f
C26 B VSUBS 1.882441f
C27 w_n1590_n1252# VSUBS 25.5481f
C28 VN.t1 VSUBS 0.302911f
C29 VN.t0 VSUBS 0.517201f
C30 VP.t1 VSUBS 0.880365f
C31 VP.t0 VSUBS 0.521138f
C32 VP.n0 VSUBS 3.4423f
C33 B.n0 VSUBS 0.006262f
C34 B.n1 VSUBS 0.006262f
C35 B.n2 VSUBS 0.009903f
C36 B.n3 VSUBS 0.009903f
C37 B.n4 VSUBS 0.009903f
C38 B.n5 VSUBS 0.009903f
C39 B.n6 VSUBS 0.009903f
C40 B.n7 VSUBS 0.009903f
C41 B.n8 VSUBS 0.009903f
C42 B.n9 VSUBS 0.009903f
C43 B.n10 VSUBS 0.022169f
C44 B.n11 VSUBS 0.009903f
C45 B.n12 VSUBS 0.009903f
C46 B.n13 VSUBS 0.009903f
C47 B.n14 VSUBS 0.009903f
C48 B.n15 VSUBS 0.009903f
C49 B.t11 VSUBS 0.0405f
C50 B.t10 VSUBS 0.045985f
C51 B.t9 VSUBS 0.121528f
C52 B.n16 VSUBS 0.0729f
C53 B.n17 VSUBS 0.065066f
C54 B.n18 VSUBS 0.022944f
C55 B.n19 VSUBS 0.009903f
C56 B.n20 VSUBS 0.009903f
C57 B.n21 VSUBS 0.009903f
C58 B.n22 VSUBS 0.009903f
C59 B.n23 VSUBS 0.009903f
C60 B.t2 VSUBS 0.0405f
C61 B.t1 VSUBS 0.045985f
C62 B.t0 VSUBS 0.121528f
C63 B.n24 VSUBS 0.0729f
C64 B.n25 VSUBS 0.065066f
C65 B.n26 VSUBS 0.009903f
C66 B.n27 VSUBS 0.009903f
C67 B.n28 VSUBS 0.009903f
C68 B.n29 VSUBS 0.009903f
C69 B.n30 VSUBS 0.022969f
C70 B.n31 VSUBS 0.009903f
C71 B.n32 VSUBS 0.009903f
C72 B.n33 VSUBS 0.009903f
C73 B.n34 VSUBS 0.009903f
C74 B.n35 VSUBS 0.009903f
C75 B.n36 VSUBS 0.009903f
C76 B.n37 VSUBS 0.009903f
C77 B.n38 VSUBS 0.009903f
C78 B.n39 VSUBS 0.009903f
C79 B.n40 VSUBS 0.009903f
C80 B.n41 VSUBS 0.009903f
C81 B.n42 VSUBS 0.009903f
C82 B.n43 VSUBS 0.009903f
C83 B.n44 VSUBS 0.009903f
C84 B.n45 VSUBS 0.009903f
C85 B.n46 VSUBS 0.009903f
C86 B.n47 VSUBS 0.009903f
C87 B.n48 VSUBS 0.02414f
C88 B.n49 VSUBS 0.009903f
C89 B.n50 VSUBS 0.009903f
C90 B.n51 VSUBS 0.009903f
C91 B.n52 VSUBS 0.009903f
C92 B.n53 VSUBS 0.009903f
C93 B.t7 VSUBS 0.0405f
C94 B.t8 VSUBS 0.045985f
C95 B.t6 VSUBS 0.121528f
C96 B.n54 VSUBS 0.0729f
C97 B.n55 VSUBS 0.065066f
C98 B.n56 VSUBS 0.009903f
C99 B.n57 VSUBS 0.009903f
C100 B.n58 VSUBS 0.009903f
C101 B.n59 VSUBS 0.009903f
C102 B.t4 VSUBS 0.0405f
C103 B.t5 VSUBS 0.045985f
C104 B.t3 VSUBS 0.121528f
C105 B.n60 VSUBS 0.0729f
C106 B.n61 VSUBS 0.065066f
C107 B.n62 VSUBS 0.022944f
C108 B.n63 VSUBS 0.009903f
C109 B.n64 VSUBS 0.009903f
C110 B.n65 VSUBS 0.009903f
C111 B.n66 VSUBS 0.009903f
C112 B.n67 VSUBS 0.009903f
C113 B.n68 VSUBS 0.022169f
C114 B.n69 VSUBS 0.009903f
C115 B.n70 VSUBS 0.009903f
C116 B.n71 VSUBS 0.009903f
C117 B.n72 VSUBS 0.009903f
C118 B.n73 VSUBS 0.009903f
C119 B.n74 VSUBS 0.009903f
C120 B.n75 VSUBS 0.009903f
C121 B.n76 VSUBS 0.009903f
C122 B.n77 VSUBS 0.009903f
C123 B.n78 VSUBS 0.009903f
C124 B.n79 VSUBS 0.009903f
C125 B.n80 VSUBS 0.009903f
C126 B.n81 VSUBS 0.009903f
C127 B.n82 VSUBS 0.009903f
C128 B.n83 VSUBS 0.009903f
C129 B.n84 VSUBS 0.009903f
C130 B.n85 VSUBS 0.009903f
C131 B.n86 VSUBS 0.009903f
C132 B.n87 VSUBS 0.009903f
C133 B.n88 VSUBS 0.009903f
C134 B.n89 VSUBS 0.009903f
C135 B.n90 VSUBS 0.009903f
C136 B.n91 VSUBS 0.009903f
C137 B.n92 VSUBS 0.009903f
C138 B.n93 VSUBS 0.009903f
C139 B.n94 VSUBS 0.009903f
C140 B.n95 VSUBS 0.009903f
C141 B.n96 VSUBS 0.009903f
C142 B.n97 VSUBS 0.009903f
C143 B.n98 VSUBS 0.009903f
C144 B.n99 VSUBS 0.022169f
C145 B.n100 VSUBS 0.02414f
C146 B.n101 VSUBS 0.02414f
C147 B.n102 VSUBS 0.009903f
C148 B.n103 VSUBS 0.009903f
C149 B.n104 VSUBS 0.009903f
C150 B.n105 VSUBS 0.009903f
C151 B.n106 VSUBS 0.009903f
C152 B.n107 VSUBS 0.009903f
C153 B.n108 VSUBS 0.009903f
C154 B.n109 VSUBS 0.009903f
C155 B.n110 VSUBS 0.009903f
C156 B.n111 VSUBS 0.009903f
C157 B.n112 VSUBS 0.009903f
C158 B.n113 VSUBS 0.009903f
C159 B.n114 VSUBS 0.009903f
C160 B.n115 VSUBS 0.006845f
C161 B.n116 VSUBS 0.009903f
C162 B.n117 VSUBS 0.009903f
C163 B.n118 VSUBS 0.00801f
C164 B.n119 VSUBS 0.009903f
C165 B.n120 VSUBS 0.009903f
C166 B.n121 VSUBS 0.009903f
C167 B.n122 VSUBS 0.009903f
C168 B.n123 VSUBS 0.009903f
C169 B.n124 VSUBS 0.009903f
C170 B.n125 VSUBS 0.009903f
C171 B.n126 VSUBS 0.009903f
C172 B.n127 VSUBS 0.009903f
C173 B.n128 VSUBS 0.009903f
C174 B.n129 VSUBS 0.009903f
C175 B.n130 VSUBS 0.00801f
C176 B.n131 VSUBS 0.022944f
C177 B.n132 VSUBS 0.006845f
C178 B.n133 VSUBS 0.009903f
C179 B.n134 VSUBS 0.009903f
C180 B.n135 VSUBS 0.009903f
C181 B.n136 VSUBS 0.009903f
C182 B.n137 VSUBS 0.009903f
C183 B.n138 VSUBS 0.009903f
C184 B.n139 VSUBS 0.009903f
C185 B.n140 VSUBS 0.009903f
C186 B.n141 VSUBS 0.009903f
C187 B.n142 VSUBS 0.009903f
C188 B.n143 VSUBS 0.009903f
C189 B.n144 VSUBS 0.009903f
C190 B.n145 VSUBS 0.009903f
C191 B.n146 VSUBS 0.009903f
C192 B.n147 VSUBS 0.02414f
C193 B.n148 VSUBS 0.022169f
C194 B.n149 VSUBS 0.022169f
C195 B.n150 VSUBS 0.009903f
C196 B.n151 VSUBS 0.009903f
C197 B.n152 VSUBS 0.009903f
C198 B.n153 VSUBS 0.009903f
C199 B.n154 VSUBS 0.009903f
C200 B.n155 VSUBS 0.009903f
C201 B.n156 VSUBS 0.009903f
C202 B.n157 VSUBS 0.009903f
C203 B.n158 VSUBS 0.009903f
C204 B.n159 VSUBS 0.009903f
C205 B.n160 VSUBS 0.009903f
C206 B.n161 VSUBS 0.009903f
C207 B.n162 VSUBS 0.009903f
C208 B.n163 VSUBS 0.009903f
C209 B.n164 VSUBS 0.009903f
C210 B.n165 VSUBS 0.009903f
C211 B.n166 VSUBS 0.009903f
C212 B.n167 VSUBS 0.009903f
C213 B.n168 VSUBS 0.009903f
C214 B.n169 VSUBS 0.009903f
C215 B.n170 VSUBS 0.009903f
C216 B.n171 VSUBS 0.009903f
C217 B.n172 VSUBS 0.009903f
C218 B.n173 VSUBS 0.009903f
C219 B.n174 VSUBS 0.009903f
C220 B.n175 VSUBS 0.009903f
C221 B.n176 VSUBS 0.009903f
C222 B.n177 VSUBS 0.009903f
C223 B.n178 VSUBS 0.009903f
C224 B.n179 VSUBS 0.009903f
C225 B.n180 VSUBS 0.009903f
C226 B.n181 VSUBS 0.009903f
C227 B.n182 VSUBS 0.009903f
C228 B.n183 VSUBS 0.009903f
C229 B.n184 VSUBS 0.009903f
C230 B.n185 VSUBS 0.009903f
C231 B.n186 VSUBS 0.009903f
C232 B.n187 VSUBS 0.009903f
C233 B.n188 VSUBS 0.009903f
C234 B.n189 VSUBS 0.009903f
C235 B.n190 VSUBS 0.009903f
C236 B.n191 VSUBS 0.009903f
C237 B.n192 VSUBS 0.009903f
C238 B.n193 VSUBS 0.009903f
C239 B.n194 VSUBS 0.009903f
C240 B.n195 VSUBS 0.009903f
C241 B.n196 VSUBS 0.009903f
C242 B.n197 VSUBS 0.009903f
C243 B.n198 VSUBS 0.009903f
C244 B.n199 VSUBS 0.023341f
C245 B.n200 VSUBS 0.022169f
C246 B.n201 VSUBS 0.02414f
C247 B.n202 VSUBS 0.009903f
C248 B.n203 VSUBS 0.009903f
C249 B.n204 VSUBS 0.009903f
C250 B.n205 VSUBS 0.009903f
C251 B.n206 VSUBS 0.009903f
C252 B.n207 VSUBS 0.009903f
C253 B.n208 VSUBS 0.009903f
C254 B.n209 VSUBS 0.009903f
C255 B.n210 VSUBS 0.009903f
C256 B.n211 VSUBS 0.009903f
C257 B.n212 VSUBS 0.009903f
C258 B.n213 VSUBS 0.009903f
C259 B.n214 VSUBS 0.009903f
C260 B.n215 VSUBS 0.009903f
C261 B.n216 VSUBS 0.006845f
C262 B.n217 VSUBS 0.022944f
C263 B.n218 VSUBS 0.00801f
C264 B.n219 VSUBS 0.009903f
C265 B.n220 VSUBS 0.009903f
C266 B.n221 VSUBS 0.009903f
C267 B.n222 VSUBS 0.009903f
C268 B.n223 VSUBS 0.009903f
C269 B.n224 VSUBS 0.009903f
C270 B.n225 VSUBS 0.009903f
C271 B.n226 VSUBS 0.009903f
C272 B.n227 VSUBS 0.009903f
C273 B.n228 VSUBS 0.009903f
C274 B.n229 VSUBS 0.009903f
C275 B.n230 VSUBS 0.00801f
C276 B.n231 VSUBS 0.009903f
C277 B.n232 VSUBS 0.009903f
C278 B.n233 VSUBS 0.006845f
C279 B.n234 VSUBS 0.009903f
C280 B.n235 VSUBS 0.009903f
C281 B.n236 VSUBS 0.009903f
C282 B.n237 VSUBS 0.009903f
C283 B.n238 VSUBS 0.009903f
C284 B.n239 VSUBS 0.009903f
C285 B.n240 VSUBS 0.009903f
C286 B.n241 VSUBS 0.009903f
C287 B.n242 VSUBS 0.009903f
C288 B.n243 VSUBS 0.009903f
C289 B.n244 VSUBS 0.009903f
C290 B.n245 VSUBS 0.009903f
C291 B.n246 VSUBS 0.009903f
C292 B.n247 VSUBS 0.02414f
C293 B.n248 VSUBS 0.02414f
C294 B.n249 VSUBS 0.022169f
C295 B.n250 VSUBS 0.009903f
C296 B.n251 VSUBS 0.009903f
C297 B.n252 VSUBS 0.009903f
C298 B.n253 VSUBS 0.009903f
C299 B.n254 VSUBS 0.009903f
C300 B.n255 VSUBS 0.009903f
C301 B.n256 VSUBS 0.009903f
C302 B.n257 VSUBS 0.009903f
C303 B.n258 VSUBS 0.009903f
C304 B.n259 VSUBS 0.009903f
C305 B.n260 VSUBS 0.009903f
C306 B.n261 VSUBS 0.009903f
C307 B.n262 VSUBS 0.009903f
C308 B.n263 VSUBS 0.009903f
C309 B.n264 VSUBS 0.009903f
C310 B.n265 VSUBS 0.009903f
C311 B.n266 VSUBS 0.009903f
C312 B.n267 VSUBS 0.009903f
C313 B.n268 VSUBS 0.009903f
C314 B.n269 VSUBS 0.009903f
C315 B.n270 VSUBS 0.009903f
C316 B.n271 VSUBS 0.009903f
C317 B.n272 VSUBS 0.009903f
C318 B.n273 VSUBS 0.009903f
C319 B.n274 VSUBS 0.009903f
C320 B.n275 VSUBS 0.022423f
.ends

