* NGSPICE file created from diff_pair_sample_1262.ext - technology: sky130A

.subckt diff_pair_sample_1262 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=0.43
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=4.4343 ps=23.52 w=11.37 l=0.43
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=4.4343 ps=23.52 w=11.37 l=0.43
X3 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=4.4343 ps=23.52 w=11.37 l=0.43
X4 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=0.43
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=0.43
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=0 ps=0 w=11.37 l=0.43
X7 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=4.4343 pd=23.52 as=4.4343 ps=23.52 w=11.37 l=0.43
R0 B.n75 B.t6 845.619
R1 B.n73 B.t13 845.619
R2 B.n295 B.t10 845.619
R3 B.n301 B.t2 845.619
R4 B.n557 B.n556 585
R5 B.n558 B.n557 585
R6 B.n251 B.n72 585
R7 B.n250 B.n249 585
R8 B.n248 B.n247 585
R9 B.n246 B.n245 585
R10 B.n244 B.n243 585
R11 B.n242 B.n241 585
R12 B.n240 B.n239 585
R13 B.n238 B.n237 585
R14 B.n236 B.n235 585
R15 B.n234 B.n233 585
R16 B.n232 B.n231 585
R17 B.n230 B.n229 585
R18 B.n228 B.n227 585
R19 B.n226 B.n225 585
R20 B.n224 B.n223 585
R21 B.n222 B.n221 585
R22 B.n220 B.n219 585
R23 B.n218 B.n217 585
R24 B.n216 B.n215 585
R25 B.n214 B.n213 585
R26 B.n212 B.n211 585
R27 B.n210 B.n209 585
R28 B.n208 B.n207 585
R29 B.n206 B.n205 585
R30 B.n204 B.n203 585
R31 B.n202 B.n201 585
R32 B.n200 B.n199 585
R33 B.n198 B.n197 585
R34 B.n196 B.n195 585
R35 B.n194 B.n193 585
R36 B.n192 B.n191 585
R37 B.n190 B.n189 585
R38 B.n188 B.n187 585
R39 B.n186 B.n185 585
R40 B.n184 B.n183 585
R41 B.n182 B.n181 585
R42 B.n180 B.n179 585
R43 B.n178 B.n177 585
R44 B.n176 B.n175 585
R45 B.n173 B.n172 585
R46 B.n171 B.n170 585
R47 B.n169 B.n168 585
R48 B.n167 B.n166 585
R49 B.n165 B.n164 585
R50 B.n163 B.n162 585
R51 B.n161 B.n160 585
R52 B.n159 B.n158 585
R53 B.n157 B.n156 585
R54 B.n155 B.n154 585
R55 B.n153 B.n152 585
R56 B.n151 B.n150 585
R57 B.n149 B.n148 585
R58 B.n147 B.n146 585
R59 B.n145 B.n144 585
R60 B.n143 B.n142 585
R61 B.n141 B.n140 585
R62 B.n139 B.n138 585
R63 B.n137 B.n136 585
R64 B.n135 B.n134 585
R65 B.n133 B.n132 585
R66 B.n131 B.n130 585
R67 B.n129 B.n128 585
R68 B.n127 B.n126 585
R69 B.n125 B.n124 585
R70 B.n123 B.n122 585
R71 B.n121 B.n120 585
R72 B.n119 B.n118 585
R73 B.n117 B.n116 585
R74 B.n115 B.n114 585
R75 B.n113 B.n112 585
R76 B.n111 B.n110 585
R77 B.n109 B.n108 585
R78 B.n107 B.n106 585
R79 B.n105 B.n104 585
R80 B.n103 B.n102 585
R81 B.n101 B.n100 585
R82 B.n99 B.n98 585
R83 B.n97 B.n96 585
R84 B.n95 B.n94 585
R85 B.n93 B.n92 585
R86 B.n91 B.n90 585
R87 B.n89 B.n88 585
R88 B.n87 B.n86 585
R89 B.n85 B.n84 585
R90 B.n83 B.n82 585
R91 B.n81 B.n80 585
R92 B.n79 B.n78 585
R93 B.n26 B.n25 585
R94 B.n555 B.n27 585
R95 B.n559 B.n27 585
R96 B.n554 B.n553 585
R97 B.n553 B.n23 585
R98 B.n552 B.n22 585
R99 B.n565 B.n22 585
R100 B.n551 B.n21 585
R101 B.n566 B.n21 585
R102 B.n550 B.n20 585
R103 B.n567 B.n20 585
R104 B.n549 B.n548 585
R105 B.n548 B.n16 585
R106 B.n547 B.n15 585
R107 B.n573 B.n15 585
R108 B.n546 B.n14 585
R109 B.n574 B.n14 585
R110 B.n545 B.n13 585
R111 B.n575 B.n13 585
R112 B.n544 B.n543 585
R113 B.n543 B.n12 585
R114 B.n542 B.n541 585
R115 B.n542 B.n8 585
R116 B.n540 B.n7 585
R117 B.n582 B.n7 585
R118 B.n539 B.n6 585
R119 B.n583 B.n6 585
R120 B.n538 B.n5 585
R121 B.n584 B.n5 585
R122 B.n537 B.n536 585
R123 B.n536 B.n4 585
R124 B.n535 B.n252 585
R125 B.n535 B.n534 585
R126 B.n524 B.n253 585
R127 B.n527 B.n253 585
R128 B.n526 B.n525 585
R129 B.n528 B.n526 585
R130 B.n523 B.n258 585
R131 B.n258 B.n257 585
R132 B.n522 B.n521 585
R133 B.n521 B.n520 585
R134 B.n260 B.n259 585
R135 B.n261 B.n260 585
R136 B.n513 B.n512 585
R137 B.n514 B.n513 585
R138 B.n511 B.n266 585
R139 B.n266 B.n265 585
R140 B.n510 B.n509 585
R141 B.n509 B.n508 585
R142 B.n268 B.n267 585
R143 B.n269 B.n268 585
R144 B.n501 B.n500 585
R145 B.n502 B.n501 585
R146 B.n272 B.n271 585
R147 B.n324 B.n322 585
R148 B.n325 B.n321 585
R149 B.n325 B.n273 585
R150 B.n328 B.n327 585
R151 B.n329 B.n320 585
R152 B.n331 B.n330 585
R153 B.n333 B.n319 585
R154 B.n336 B.n335 585
R155 B.n337 B.n318 585
R156 B.n339 B.n338 585
R157 B.n341 B.n317 585
R158 B.n344 B.n343 585
R159 B.n345 B.n316 585
R160 B.n347 B.n346 585
R161 B.n349 B.n315 585
R162 B.n352 B.n351 585
R163 B.n353 B.n314 585
R164 B.n355 B.n354 585
R165 B.n357 B.n313 585
R166 B.n360 B.n359 585
R167 B.n361 B.n312 585
R168 B.n363 B.n362 585
R169 B.n365 B.n311 585
R170 B.n368 B.n367 585
R171 B.n369 B.n310 585
R172 B.n371 B.n370 585
R173 B.n373 B.n309 585
R174 B.n376 B.n375 585
R175 B.n377 B.n308 585
R176 B.n379 B.n378 585
R177 B.n381 B.n307 585
R178 B.n384 B.n383 585
R179 B.n385 B.n306 585
R180 B.n387 B.n386 585
R181 B.n389 B.n305 585
R182 B.n392 B.n391 585
R183 B.n393 B.n304 585
R184 B.n395 B.n394 585
R185 B.n397 B.n303 585
R186 B.n400 B.n399 585
R187 B.n402 B.n300 585
R188 B.n404 B.n403 585
R189 B.n406 B.n299 585
R190 B.n409 B.n408 585
R191 B.n410 B.n298 585
R192 B.n412 B.n411 585
R193 B.n414 B.n297 585
R194 B.n417 B.n416 585
R195 B.n418 B.n294 585
R196 B.n421 B.n420 585
R197 B.n423 B.n293 585
R198 B.n426 B.n425 585
R199 B.n427 B.n292 585
R200 B.n429 B.n428 585
R201 B.n431 B.n291 585
R202 B.n434 B.n433 585
R203 B.n435 B.n290 585
R204 B.n437 B.n436 585
R205 B.n439 B.n289 585
R206 B.n442 B.n441 585
R207 B.n443 B.n288 585
R208 B.n445 B.n444 585
R209 B.n447 B.n287 585
R210 B.n450 B.n449 585
R211 B.n451 B.n286 585
R212 B.n453 B.n452 585
R213 B.n455 B.n285 585
R214 B.n458 B.n457 585
R215 B.n459 B.n284 585
R216 B.n461 B.n460 585
R217 B.n463 B.n283 585
R218 B.n466 B.n465 585
R219 B.n467 B.n282 585
R220 B.n469 B.n468 585
R221 B.n471 B.n281 585
R222 B.n474 B.n473 585
R223 B.n475 B.n280 585
R224 B.n477 B.n476 585
R225 B.n479 B.n279 585
R226 B.n482 B.n481 585
R227 B.n483 B.n278 585
R228 B.n485 B.n484 585
R229 B.n487 B.n277 585
R230 B.n490 B.n489 585
R231 B.n491 B.n276 585
R232 B.n493 B.n492 585
R233 B.n495 B.n275 585
R234 B.n498 B.n497 585
R235 B.n499 B.n274 585
R236 B.n504 B.n503 585
R237 B.n503 B.n502 585
R238 B.n505 B.n270 585
R239 B.n270 B.n269 585
R240 B.n507 B.n506 585
R241 B.n508 B.n507 585
R242 B.n264 B.n263 585
R243 B.n265 B.n264 585
R244 B.n516 B.n515 585
R245 B.n515 B.n514 585
R246 B.n517 B.n262 585
R247 B.n262 B.n261 585
R248 B.n519 B.n518 585
R249 B.n520 B.n519 585
R250 B.n256 B.n255 585
R251 B.n257 B.n256 585
R252 B.n530 B.n529 585
R253 B.n529 B.n528 585
R254 B.n531 B.n254 585
R255 B.n527 B.n254 585
R256 B.n533 B.n532 585
R257 B.n534 B.n533 585
R258 B.n3 B.n0 585
R259 B.n4 B.n3 585
R260 B.n581 B.n1 585
R261 B.n582 B.n581 585
R262 B.n580 B.n579 585
R263 B.n580 B.n8 585
R264 B.n578 B.n9 585
R265 B.n12 B.n9 585
R266 B.n577 B.n576 585
R267 B.n576 B.n575 585
R268 B.n11 B.n10 585
R269 B.n574 B.n11 585
R270 B.n572 B.n571 585
R271 B.n573 B.n572 585
R272 B.n570 B.n17 585
R273 B.n17 B.n16 585
R274 B.n569 B.n568 585
R275 B.n568 B.n567 585
R276 B.n19 B.n18 585
R277 B.n566 B.n19 585
R278 B.n564 B.n563 585
R279 B.n565 B.n564 585
R280 B.n562 B.n24 585
R281 B.n24 B.n23 585
R282 B.n561 B.n560 585
R283 B.n560 B.n559 585
R284 B.n585 B.n584 585
R285 B.n583 B.n2 585
R286 B.n560 B.n26 530.939
R287 B.n557 B.n27 530.939
R288 B.n501 B.n274 530.939
R289 B.n503 B.n272 530.939
R290 B.n73 B.t14 286.005
R291 B.n295 B.t12 286.005
R292 B.n75 B.t8 286.005
R293 B.n301 B.t5 286.005
R294 B.n74 B.t15 271.265
R295 B.n296 B.t11 271.265
R296 B.n76 B.t9 271.265
R297 B.n302 B.t4 271.265
R298 B.n558 B.n71 256.663
R299 B.n558 B.n70 256.663
R300 B.n558 B.n69 256.663
R301 B.n558 B.n68 256.663
R302 B.n558 B.n67 256.663
R303 B.n558 B.n66 256.663
R304 B.n558 B.n65 256.663
R305 B.n558 B.n64 256.663
R306 B.n558 B.n63 256.663
R307 B.n558 B.n62 256.663
R308 B.n558 B.n61 256.663
R309 B.n558 B.n60 256.663
R310 B.n558 B.n59 256.663
R311 B.n558 B.n58 256.663
R312 B.n558 B.n57 256.663
R313 B.n558 B.n56 256.663
R314 B.n558 B.n55 256.663
R315 B.n558 B.n54 256.663
R316 B.n558 B.n53 256.663
R317 B.n558 B.n52 256.663
R318 B.n558 B.n51 256.663
R319 B.n558 B.n50 256.663
R320 B.n558 B.n49 256.663
R321 B.n558 B.n48 256.663
R322 B.n558 B.n47 256.663
R323 B.n558 B.n46 256.663
R324 B.n558 B.n45 256.663
R325 B.n558 B.n44 256.663
R326 B.n558 B.n43 256.663
R327 B.n558 B.n42 256.663
R328 B.n558 B.n41 256.663
R329 B.n558 B.n40 256.663
R330 B.n558 B.n39 256.663
R331 B.n558 B.n38 256.663
R332 B.n558 B.n37 256.663
R333 B.n558 B.n36 256.663
R334 B.n558 B.n35 256.663
R335 B.n558 B.n34 256.663
R336 B.n558 B.n33 256.663
R337 B.n558 B.n32 256.663
R338 B.n558 B.n31 256.663
R339 B.n558 B.n30 256.663
R340 B.n558 B.n29 256.663
R341 B.n558 B.n28 256.663
R342 B.n323 B.n273 256.663
R343 B.n326 B.n273 256.663
R344 B.n332 B.n273 256.663
R345 B.n334 B.n273 256.663
R346 B.n340 B.n273 256.663
R347 B.n342 B.n273 256.663
R348 B.n348 B.n273 256.663
R349 B.n350 B.n273 256.663
R350 B.n356 B.n273 256.663
R351 B.n358 B.n273 256.663
R352 B.n364 B.n273 256.663
R353 B.n366 B.n273 256.663
R354 B.n372 B.n273 256.663
R355 B.n374 B.n273 256.663
R356 B.n380 B.n273 256.663
R357 B.n382 B.n273 256.663
R358 B.n388 B.n273 256.663
R359 B.n390 B.n273 256.663
R360 B.n396 B.n273 256.663
R361 B.n398 B.n273 256.663
R362 B.n405 B.n273 256.663
R363 B.n407 B.n273 256.663
R364 B.n413 B.n273 256.663
R365 B.n415 B.n273 256.663
R366 B.n422 B.n273 256.663
R367 B.n424 B.n273 256.663
R368 B.n430 B.n273 256.663
R369 B.n432 B.n273 256.663
R370 B.n438 B.n273 256.663
R371 B.n440 B.n273 256.663
R372 B.n446 B.n273 256.663
R373 B.n448 B.n273 256.663
R374 B.n454 B.n273 256.663
R375 B.n456 B.n273 256.663
R376 B.n462 B.n273 256.663
R377 B.n464 B.n273 256.663
R378 B.n470 B.n273 256.663
R379 B.n472 B.n273 256.663
R380 B.n478 B.n273 256.663
R381 B.n480 B.n273 256.663
R382 B.n486 B.n273 256.663
R383 B.n488 B.n273 256.663
R384 B.n494 B.n273 256.663
R385 B.n496 B.n273 256.663
R386 B.n587 B.n586 256.663
R387 B.n80 B.n79 163.367
R388 B.n84 B.n83 163.367
R389 B.n88 B.n87 163.367
R390 B.n92 B.n91 163.367
R391 B.n96 B.n95 163.367
R392 B.n100 B.n99 163.367
R393 B.n104 B.n103 163.367
R394 B.n108 B.n107 163.367
R395 B.n112 B.n111 163.367
R396 B.n116 B.n115 163.367
R397 B.n120 B.n119 163.367
R398 B.n124 B.n123 163.367
R399 B.n128 B.n127 163.367
R400 B.n132 B.n131 163.367
R401 B.n136 B.n135 163.367
R402 B.n140 B.n139 163.367
R403 B.n144 B.n143 163.367
R404 B.n148 B.n147 163.367
R405 B.n152 B.n151 163.367
R406 B.n156 B.n155 163.367
R407 B.n160 B.n159 163.367
R408 B.n164 B.n163 163.367
R409 B.n168 B.n167 163.367
R410 B.n172 B.n171 163.367
R411 B.n177 B.n176 163.367
R412 B.n181 B.n180 163.367
R413 B.n185 B.n184 163.367
R414 B.n189 B.n188 163.367
R415 B.n193 B.n192 163.367
R416 B.n197 B.n196 163.367
R417 B.n201 B.n200 163.367
R418 B.n205 B.n204 163.367
R419 B.n209 B.n208 163.367
R420 B.n213 B.n212 163.367
R421 B.n217 B.n216 163.367
R422 B.n221 B.n220 163.367
R423 B.n225 B.n224 163.367
R424 B.n229 B.n228 163.367
R425 B.n233 B.n232 163.367
R426 B.n237 B.n236 163.367
R427 B.n241 B.n240 163.367
R428 B.n245 B.n244 163.367
R429 B.n249 B.n248 163.367
R430 B.n557 B.n72 163.367
R431 B.n501 B.n268 163.367
R432 B.n509 B.n268 163.367
R433 B.n509 B.n266 163.367
R434 B.n513 B.n266 163.367
R435 B.n513 B.n260 163.367
R436 B.n521 B.n260 163.367
R437 B.n521 B.n258 163.367
R438 B.n526 B.n258 163.367
R439 B.n526 B.n253 163.367
R440 B.n535 B.n253 163.367
R441 B.n536 B.n535 163.367
R442 B.n536 B.n5 163.367
R443 B.n6 B.n5 163.367
R444 B.n7 B.n6 163.367
R445 B.n542 B.n7 163.367
R446 B.n543 B.n542 163.367
R447 B.n543 B.n13 163.367
R448 B.n14 B.n13 163.367
R449 B.n15 B.n14 163.367
R450 B.n548 B.n15 163.367
R451 B.n548 B.n20 163.367
R452 B.n21 B.n20 163.367
R453 B.n22 B.n21 163.367
R454 B.n553 B.n22 163.367
R455 B.n553 B.n27 163.367
R456 B.n325 B.n324 163.367
R457 B.n327 B.n325 163.367
R458 B.n331 B.n320 163.367
R459 B.n335 B.n333 163.367
R460 B.n339 B.n318 163.367
R461 B.n343 B.n341 163.367
R462 B.n347 B.n316 163.367
R463 B.n351 B.n349 163.367
R464 B.n355 B.n314 163.367
R465 B.n359 B.n357 163.367
R466 B.n363 B.n312 163.367
R467 B.n367 B.n365 163.367
R468 B.n371 B.n310 163.367
R469 B.n375 B.n373 163.367
R470 B.n379 B.n308 163.367
R471 B.n383 B.n381 163.367
R472 B.n387 B.n306 163.367
R473 B.n391 B.n389 163.367
R474 B.n395 B.n304 163.367
R475 B.n399 B.n397 163.367
R476 B.n404 B.n300 163.367
R477 B.n408 B.n406 163.367
R478 B.n412 B.n298 163.367
R479 B.n416 B.n414 163.367
R480 B.n421 B.n294 163.367
R481 B.n425 B.n423 163.367
R482 B.n429 B.n292 163.367
R483 B.n433 B.n431 163.367
R484 B.n437 B.n290 163.367
R485 B.n441 B.n439 163.367
R486 B.n445 B.n288 163.367
R487 B.n449 B.n447 163.367
R488 B.n453 B.n286 163.367
R489 B.n457 B.n455 163.367
R490 B.n461 B.n284 163.367
R491 B.n465 B.n463 163.367
R492 B.n469 B.n282 163.367
R493 B.n473 B.n471 163.367
R494 B.n477 B.n280 163.367
R495 B.n481 B.n479 163.367
R496 B.n485 B.n278 163.367
R497 B.n489 B.n487 163.367
R498 B.n493 B.n276 163.367
R499 B.n497 B.n495 163.367
R500 B.n503 B.n270 163.367
R501 B.n507 B.n270 163.367
R502 B.n507 B.n264 163.367
R503 B.n515 B.n264 163.367
R504 B.n515 B.n262 163.367
R505 B.n519 B.n262 163.367
R506 B.n519 B.n256 163.367
R507 B.n529 B.n256 163.367
R508 B.n529 B.n254 163.367
R509 B.n533 B.n254 163.367
R510 B.n533 B.n3 163.367
R511 B.n585 B.n3 163.367
R512 B.n581 B.n2 163.367
R513 B.n581 B.n580 163.367
R514 B.n580 B.n9 163.367
R515 B.n576 B.n9 163.367
R516 B.n576 B.n11 163.367
R517 B.n572 B.n11 163.367
R518 B.n572 B.n17 163.367
R519 B.n568 B.n17 163.367
R520 B.n568 B.n19 163.367
R521 B.n564 B.n19 163.367
R522 B.n564 B.n24 163.367
R523 B.n560 B.n24 163.367
R524 B.n502 B.n273 85.149
R525 B.n559 B.n558 85.149
R526 B.n28 B.n26 71.676
R527 B.n80 B.n29 71.676
R528 B.n84 B.n30 71.676
R529 B.n88 B.n31 71.676
R530 B.n92 B.n32 71.676
R531 B.n96 B.n33 71.676
R532 B.n100 B.n34 71.676
R533 B.n104 B.n35 71.676
R534 B.n108 B.n36 71.676
R535 B.n112 B.n37 71.676
R536 B.n116 B.n38 71.676
R537 B.n120 B.n39 71.676
R538 B.n124 B.n40 71.676
R539 B.n128 B.n41 71.676
R540 B.n132 B.n42 71.676
R541 B.n136 B.n43 71.676
R542 B.n140 B.n44 71.676
R543 B.n144 B.n45 71.676
R544 B.n148 B.n46 71.676
R545 B.n152 B.n47 71.676
R546 B.n156 B.n48 71.676
R547 B.n160 B.n49 71.676
R548 B.n164 B.n50 71.676
R549 B.n168 B.n51 71.676
R550 B.n172 B.n52 71.676
R551 B.n177 B.n53 71.676
R552 B.n181 B.n54 71.676
R553 B.n185 B.n55 71.676
R554 B.n189 B.n56 71.676
R555 B.n193 B.n57 71.676
R556 B.n197 B.n58 71.676
R557 B.n201 B.n59 71.676
R558 B.n205 B.n60 71.676
R559 B.n209 B.n61 71.676
R560 B.n213 B.n62 71.676
R561 B.n217 B.n63 71.676
R562 B.n221 B.n64 71.676
R563 B.n225 B.n65 71.676
R564 B.n229 B.n66 71.676
R565 B.n233 B.n67 71.676
R566 B.n237 B.n68 71.676
R567 B.n241 B.n69 71.676
R568 B.n245 B.n70 71.676
R569 B.n249 B.n71 71.676
R570 B.n72 B.n71 71.676
R571 B.n248 B.n70 71.676
R572 B.n244 B.n69 71.676
R573 B.n240 B.n68 71.676
R574 B.n236 B.n67 71.676
R575 B.n232 B.n66 71.676
R576 B.n228 B.n65 71.676
R577 B.n224 B.n64 71.676
R578 B.n220 B.n63 71.676
R579 B.n216 B.n62 71.676
R580 B.n212 B.n61 71.676
R581 B.n208 B.n60 71.676
R582 B.n204 B.n59 71.676
R583 B.n200 B.n58 71.676
R584 B.n196 B.n57 71.676
R585 B.n192 B.n56 71.676
R586 B.n188 B.n55 71.676
R587 B.n184 B.n54 71.676
R588 B.n180 B.n53 71.676
R589 B.n176 B.n52 71.676
R590 B.n171 B.n51 71.676
R591 B.n167 B.n50 71.676
R592 B.n163 B.n49 71.676
R593 B.n159 B.n48 71.676
R594 B.n155 B.n47 71.676
R595 B.n151 B.n46 71.676
R596 B.n147 B.n45 71.676
R597 B.n143 B.n44 71.676
R598 B.n139 B.n43 71.676
R599 B.n135 B.n42 71.676
R600 B.n131 B.n41 71.676
R601 B.n127 B.n40 71.676
R602 B.n123 B.n39 71.676
R603 B.n119 B.n38 71.676
R604 B.n115 B.n37 71.676
R605 B.n111 B.n36 71.676
R606 B.n107 B.n35 71.676
R607 B.n103 B.n34 71.676
R608 B.n99 B.n33 71.676
R609 B.n95 B.n32 71.676
R610 B.n91 B.n31 71.676
R611 B.n87 B.n30 71.676
R612 B.n83 B.n29 71.676
R613 B.n79 B.n28 71.676
R614 B.n323 B.n272 71.676
R615 B.n327 B.n326 71.676
R616 B.n332 B.n331 71.676
R617 B.n335 B.n334 71.676
R618 B.n340 B.n339 71.676
R619 B.n343 B.n342 71.676
R620 B.n348 B.n347 71.676
R621 B.n351 B.n350 71.676
R622 B.n356 B.n355 71.676
R623 B.n359 B.n358 71.676
R624 B.n364 B.n363 71.676
R625 B.n367 B.n366 71.676
R626 B.n372 B.n371 71.676
R627 B.n375 B.n374 71.676
R628 B.n380 B.n379 71.676
R629 B.n383 B.n382 71.676
R630 B.n388 B.n387 71.676
R631 B.n391 B.n390 71.676
R632 B.n396 B.n395 71.676
R633 B.n399 B.n398 71.676
R634 B.n405 B.n404 71.676
R635 B.n408 B.n407 71.676
R636 B.n413 B.n412 71.676
R637 B.n416 B.n415 71.676
R638 B.n422 B.n421 71.676
R639 B.n425 B.n424 71.676
R640 B.n430 B.n429 71.676
R641 B.n433 B.n432 71.676
R642 B.n438 B.n437 71.676
R643 B.n441 B.n440 71.676
R644 B.n446 B.n445 71.676
R645 B.n449 B.n448 71.676
R646 B.n454 B.n453 71.676
R647 B.n457 B.n456 71.676
R648 B.n462 B.n461 71.676
R649 B.n465 B.n464 71.676
R650 B.n470 B.n469 71.676
R651 B.n473 B.n472 71.676
R652 B.n478 B.n477 71.676
R653 B.n481 B.n480 71.676
R654 B.n486 B.n485 71.676
R655 B.n489 B.n488 71.676
R656 B.n494 B.n493 71.676
R657 B.n497 B.n496 71.676
R658 B.n324 B.n323 71.676
R659 B.n326 B.n320 71.676
R660 B.n333 B.n332 71.676
R661 B.n334 B.n318 71.676
R662 B.n341 B.n340 71.676
R663 B.n342 B.n316 71.676
R664 B.n349 B.n348 71.676
R665 B.n350 B.n314 71.676
R666 B.n357 B.n356 71.676
R667 B.n358 B.n312 71.676
R668 B.n365 B.n364 71.676
R669 B.n366 B.n310 71.676
R670 B.n373 B.n372 71.676
R671 B.n374 B.n308 71.676
R672 B.n381 B.n380 71.676
R673 B.n382 B.n306 71.676
R674 B.n389 B.n388 71.676
R675 B.n390 B.n304 71.676
R676 B.n397 B.n396 71.676
R677 B.n398 B.n300 71.676
R678 B.n406 B.n405 71.676
R679 B.n407 B.n298 71.676
R680 B.n414 B.n413 71.676
R681 B.n415 B.n294 71.676
R682 B.n423 B.n422 71.676
R683 B.n424 B.n292 71.676
R684 B.n431 B.n430 71.676
R685 B.n432 B.n290 71.676
R686 B.n439 B.n438 71.676
R687 B.n440 B.n288 71.676
R688 B.n447 B.n446 71.676
R689 B.n448 B.n286 71.676
R690 B.n455 B.n454 71.676
R691 B.n456 B.n284 71.676
R692 B.n463 B.n462 71.676
R693 B.n464 B.n282 71.676
R694 B.n471 B.n470 71.676
R695 B.n472 B.n280 71.676
R696 B.n479 B.n478 71.676
R697 B.n480 B.n278 71.676
R698 B.n487 B.n486 71.676
R699 B.n488 B.n276 71.676
R700 B.n495 B.n494 71.676
R701 B.n496 B.n274 71.676
R702 B.n586 B.n585 71.676
R703 B.n586 B.n2 71.676
R704 B.n77 B.n76 59.5399
R705 B.n174 B.n74 59.5399
R706 B.n419 B.n296 59.5399
R707 B.n401 B.n302 59.5399
R708 B.n502 B.n269 44.885
R709 B.n508 B.n269 44.885
R710 B.n508 B.n265 44.885
R711 B.n514 B.n265 44.885
R712 B.n520 B.n261 44.885
R713 B.n520 B.n257 44.885
R714 B.n528 B.n257 44.885
R715 B.n528 B.n527 44.885
R716 B.n534 B.n4 44.885
R717 B.n584 B.n4 44.885
R718 B.n584 B.n583 44.885
R719 B.n583 B.n582 44.885
R720 B.n582 B.n8 44.885
R721 B.n575 B.n12 44.885
R722 B.n575 B.n574 44.885
R723 B.n574 B.n573 44.885
R724 B.n573 B.n16 44.885
R725 B.n567 B.n566 44.885
R726 B.n566 B.n565 44.885
R727 B.n565 B.n23 44.885
R728 B.n559 B.n23 44.885
R729 B.n527 B.t1 34.984
R730 B.n12 B.t0 34.984
R731 B.n504 B.n271 34.4981
R732 B.n500 B.n499 34.4981
R733 B.n556 B.n555 34.4981
R734 B.n561 B.n25 34.4981
R735 B.t3 B.n261 29.7035
R736 B.t7 B.n16 29.7035
R737 B B.n587 18.0485
R738 B.n514 B.t3 15.182
R739 B.n567 B.t7 15.182
R740 B.n76 B.n75 14.7399
R741 B.n74 B.n73 14.7399
R742 B.n296 B.n295 14.7399
R743 B.n302 B.n301 14.7399
R744 B.n505 B.n504 10.6151
R745 B.n506 B.n505 10.6151
R746 B.n506 B.n263 10.6151
R747 B.n516 B.n263 10.6151
R748 B.n517 B.n516 10.6151
R749 B.n518 B.n517 10.6151
R750 B.n518 B.n255 10.6151
R751 B.n530 B.n255 10.6151
R752 B.n531 B.n530 10.6151
R753 B.n532 B.n531 10.6151
R754 B.n532 B.n0 10.6151
R755 B.n322 B.n271 10.6151
R756 B.n322 B.n321 10.6151
R757 B.n328 B.n321 10.6151
R758 B.n329 B.n328 10.6151
R759 B.n330 B.n329 10.6151
R760 B.n330 B.n319 10.6151
R761 B.n336 B.n319 10.6151
R762 B.n337 B.n336 10.6151
R763 B.n338 B.n337 10.6151
R764 B.n338 B.n317 10.6151
R765 B.n344 B.n317 10.6151
R766 B.n345 B.n344 10.6151
R767 B.n346 B.n345 10.6151
R768 B.n346 B.n315 10.6151
R769 B.n352 B.n315 10.6151
R770 B.n353 B.n352 10.6151
R771 B.n354 B.n353 10.6151
R772 B.n354 B.n313 10.6151
R773 B.n360 B.n313 10.6151
R774 B.n361 B.n360 10.6151
R775 B.n362 B.n361 10.6151
R776 B.n362 B.n311 10.6151
R777 B.n368 B.n311 10.6151
R778 B.n369 B.n368 10.6151
R779 B.n370 B.n369 10.6151
R780 B.n370 B.n309 10.6151
R781 B.n376 B.n309 10.6151
R782 B.n377 B.n376 10.6151
R783 B.n378 B.n377 10.6151
R784 B.n378 B.n307 10.6151
R785 B.n384 B.n307 10.6151
R786 B.n385 B.n384 10.6151
R787 B.n386 B.n385 10.6151
R788 B.n386 B.n305 10.6151
R789 B.n392 B.n305 10.6151
R790 B.n393 B.n392 10.6151
R791 B.n394 B.n393 10.6151
R792 B.n394 B.n303 10.6151
R793 B.n400 B.n303 10.6151
R794 B.n403 B.n402 10.6151
R795 B.n403 B.n299 10.6151
R796 B.n409 B.n299 10.6151
R797 B.n410 B.n409 10.6151
R798 B.n411 B.n410 10.6151
R799 B.n411 B.n297 10.6151
R800 B.n417 B.n297 10.6151
R801 B.n418 B.n417 10.6151
R802 B.n420 B.n293 10.6151
R803 B.n426 B.n293 10.6151
R804 B.n427 B.n426 10.6151
R805 B.n428 B.n427 10.6151
R806 B.n428 B.n291 10.6151
R807 B.n434 B.n291 10.6151
R808 B.n435 B.n434 10.6151
R809 B.n436 B.n435 10.6151
R810 B.n436 B.n289 10.6151
R811 B.n442 B.n289 10.6151
R812 B.n443 B.n442 10.6151
R813 B.n444 B.n443 10.6151
R814 B.n444 B.n287 10.6151
R815 B.n450 B.n287 10.6151
R816 B.n451 B.n450 10.6151
R817 B.n452 B.n451 10.6151
R818 B.n452 B.n285 10.6151
R819 B.n458 B.n285 10.6151
R820 B.n459 B.n458 10.6151
R821 B.n460 B.n459 10.6151
R822 B.n460 B.n283 10.6151
R823 B.n466 B.n283 10.6151
R824 B.n467 B.n466 10.6151
R825 B.n468 B.n467 10.6151
R826 B.n468 B.n281 10.6151
R827 B.n474 B.n281 10.6151
R828 B.n475 B.n474 10.6151
R829 B.n476 B.n475 10.6151
R830 B.n476 B.n279 10.6151
R831 B.n482 B.n279 10.6151
R832 B.n483 B.n482 10.6151
R833 B.n484 B.n483 10.6151
R834 B.n484 B.n277 10.6151
R835 B.n490 B.n277 10.6151
R836 B.n491 B.n490 10.6151
R837 B.n492 B.n491 10.6151
R838 B.n492 B.n275 10.6151
R839 B.n498 B.n275 10.6151
R840 B.n499 B.n498 10.6151
R841 B.n500 B.n267 10.6151
R842 B.n510 B.n267 10.6151
R843 B.n511 B.n510 10.6151
R844 B.n512 B.n511 10.6151
R845 B.n512 B.n259 10.6151
R846 B.n522 B.n259 10.6151
R847 B.n523 B.n522 10.6151
R848 B.n525 B.n523 10.6151
R849 B.n525 B.n524 10.6151
R850 B.n524 B.n252 10.6151
R851 B.n537 B.n252 10.6151
R852 B.n538 B.n537 10.6151
R853 B.n539 B.n538 10.6151
R854 B.n540 B.n539 10.6151
R855 B.n541 B.n540 10.6151
R856 B.n544 B.n541 10.6151
R857 B.n545 B.n544 10.6151
R858 B.n546 B.n545 10.6151
R859 B.n547 B.n546 10.6151
R860 B.n549 B.n547 10.6151
R861 B.n550 B.n549 10.6151
R862 B.n551 B.n550 10.6151
R863 B.n552 B.n551 10.6151
R864 B.n554 B.n552 10.6151
R865 B.n555 B.n554 10.6151
R866 B.n579 B.n1 10.6151
R867 B.n579 B.n578 10.6151
R868 B.n578 B.n577 10.6151
R869 B.n577 B.n10 10.6151
R870 B.n571 B.n10 10.6151
R871 B.n571 B.n570 10.6151
R872 B.n570 B.n569 10.6151
R873 B.n569 B.n18 10.6151
R874 B.n563 B.n18 10.6151
R875 B.n563 B.n562 10.6151
R876 B.n562 B.n561 10.6151
R877 B.n78 B.n25 10.6151
R878 B.n81 B.n78 10.6151
R879 B.n82 B.n81 10.6151
R880 B.n85 B.n82 10.6151
R881 B.n86 B.n85 10.6151
R882 B.n89 B.n86 10.6151
R883 B.n90 B.n89 10.6151
R884 B.n93 B.n90 10.6151
R885 B.n94 B.n93 10.6151
R886 B.n97 B.n94 10.6151
R887 B.n98 B.n97 10.6151
R888 B.n101 B.n98 10.6151
R889 B.n102 B.n101 10.6151
R890 B.n105 B.n102 10.6151
R891 B.n106 B.n105 10.6151
R892 B.n109 B.n106 10.6151
R893 B.n110 B.n109 10.6151
R894 B.n113 B.n110 10.6151
R895 B.n114 B.n113 10.6151
R896 B.n117 B.n114 10.6151
R897 B.n118 B.n117 10.6151
R898 B.n121 B.n118 10.6151
R899 B.n122 B.n121 10.6151
R900 B.n125 B.n122 10.6151
R901 B.n126 B.n125 10.6151
R902 B.n129 B.n126 10.6151
R903 B.n130 B.n129 10.6151
R904 B.n133 B.n130 10.6151
R905 B.n134 B.n133 10.6151
R906 B.n137 B.n134 10.6151
R907 B.n138 B.n137 10.6151
R908 B.n141 B.n138 10.6151
R909 B.n142 B.n141 10.6151
R910 B.n145 B.n142 10.6151
R911 B.n146 B.n145 10.6151
R912 B.n149 B.n146 10.6151
R913 B.n150 B.n149 10.6151
R914 B.n153 B.n150 10.6151
R915 B.n154 B.n153 10.6151
R916 B.n158 B.n157 10.6151
R917 B.n161 B.n158 10.6151
R918 B.n162 B.n161 10.6151
R919 B.n165 B.n162 10.6151
R920 B.n166 B.n165 10.6151
R921 B.n169 B.n166 10.6151
R922 B.n170 B.n169 10.6151
R923 B.n173 B.n170 10.6151
R924 B.n178 B.n175 10.6151
R925 B.n179 B.n178 10.6151
R926 B.n182 B.n179 10.6151
R927 B.n183 B.n182 10.6151
R928 B.n186 B.n183 10.6151
R929 B.n187 B.n186 10.6151
R930 B.n190 B.n187 10.6151
R931 B.n191 B.n190 10.6151
R932 B.n194 B.n191 10.6151
R933 B.n195 B.n194 10.6151
R934 B.n198 B.n195 10.6151
R935 B.n199 B.n198 10.6151
R936 B.n202 B.n199 10.6151
R937 B.n203 B.n202 10.6151
R938 B.n206 B.n203 10.6151
R939 B.n207 B.n206 10.6151
R940 B.n210 B.n207 10.6151
R941 B.n211 B.n210 10.6151
R942 B.n214 B.n211 10.6151
R943 B.n215 B.n214 10.6151
R944 B.n218 B.n215 10.6151
R945 B.n219 B.n218 10.6151
R946 B.n222 B.n219 10.6151
R947 B.n223 B.n222 10.6151
R948 B.n226 B.n223 10.6151
R949 B.n227 B.n226 10.6151
R950 B.n230 B.n227 10.6151
R951 B.n231 B.n230 10.6151
R952 B.n234 B.n231 10.6151
R953 B.n235 B.n234 10.6151
R954 B.n238 B.n235 10.6151
R955 B.n239 B.n238 10.6151
R956 B.n242 B.n239 10.6151
R957 B.n243 B.n242 10.6151
R958 B.n246 B.n243 10.6151
R959 B.n247 B.n246 10.6151
R960 B.n250 B.n247 10.6151
R961 B.n251 B.n250 10.6151
R962 B.n556 B.n251 10.6151
R963 B.n534 B.t1 9.90149
R964 B.t0 B.n8 9.90149
R965 B.n587 B.n0 8.11757
R966 B.n587 B.n1 8.11757
R967 B.n402 B.n401 7.18099
R968 B.n419 B.n418 7.18099
R969 B.n157 B.n77 7.18099
R970 B.n174 B.n173 7.18099
R971 B.n401 B.n400 3.43465
R972 B.n420 B.n419 3.43465
R973 B.n154 B.n77 3.43465
R974 B.n175 B.n174 3.43465
R975 VN VN.t0 929.285
R976 VN VN.t1 890.516
R977 VTAIL.n242 VTAIL.n186 289.615
R978 VTAIL.n56 VTAIL.n0 289.615
R979 VTAIL.n180 VTAIL.n124 289.615
R980 VTAIL.n118 VTAIL.n62 289.615
R981 VTAIL.n207 VTAIL.n206 185
R982 VTAIL.n209 VTAIL.n208 185
R983 VTAIL.n202 VTAIL.n201 185
R984 VTAIL.n215 VTAIL.n214 185
R985 VTAIL.n217 VTAIL.n216 185
R986 VTAIL.n198 VTAIL.n197 185
R987 VTAIL.n224 VTAIL.n223 185
R988 VTAIL.n225 VTAIL.n196 185
R989 VTAIL.n227 VTAIL.n226 185
R990 VTAIL.n194 VTAIL.n193 185
R991 VTAIL.n233 VTAIL.n232 185
R992 VTAIL.n235 VTAIL.n234 185
R993 VTAIL.n190 VTAIL.n189 185
R994 VTAIL.n241 VTAIL.n240 185
R995 VTAIL.n243 VTAIL.n242 185
R996 VTAIL.n21 VTAIL.n20 185
R997 VTAIL.n23 VTAIL.n22 185
R998 VTAIL.n16 VTAIL.n15 185
R999 VTAIL.n29 VTAIL.n28 185
R1000 VTAIL.n31 VTAIL.n30 185
R1001 VTAIL.n12 VTAIL.n11 185
R1002 VTAIL.n38 VTAIL.n37 185
R1003 VTAIL.n39 VTAIL.n10 185
R1004 VTAIL.n41 VTAIL.n40 185
R1005 VTAIL.n8 VTAIL.n7 185
R1006 VTAIL.n47 VTAIL.n46 185
R1007 VTAIL.n49 VTAIL.n48 185
R1008 VTAIL.n4 VTAIL.n3 185
R1009 VTAIL.n55 VTAIL.n54 185
R1010 VTAIL.n57 VTAIL.n56 185
R1011 VTAIL.n181 VTAIL.n180 185
R1012 VTAIL.n179 VTAIL.n178 185
R1013 VTAIL.n128 VTAIL.n127 185
R1014 VTAIL.n173 VTAIL.n172 185
R1015 VTAIL.n171 VTAIL.n170 185
R1016 VTAIL.n132 VTAIL.n131 185
R1017 VTAIL.n136 VTAIL.n134 185
R1018 VTAIL.n165 VTAIL.n164 185
R1019 VTAIL.n163 VTAIL.n162 185
R1020 VTAIL.n138 VTAIL.n137 185
R1021 VTAIL.n157 VTAIL.n156 185
R1022 VTAIL.n155 VTAIL.n154 185
R1023 VTAIL.n142 VTAIL.n141 185
R1024 VTAIL.n149 VTAIL.n148 185
R1025 VTAIL.n147 VTAIL.n146 185
R1026 VTAIL.n119 VTAIL.n118 185
R1027 VTAIL.n117 VTAIL.n116 185
R1028 VTAIL.n66 VTAIL.n65 185
R1029 VTAIL.n111 VTAIL.n110 185
R1030 VTAIL.n109 VTAIL.n108 185
R1031 VTAIL.n70 VTAIL.n69 185
R1032 VTAIL.n74 VTAIL.n72 185
R1033 VTAIL.n103 VTAIL.n102 185
R1034 VTAIL.n101 VTAIL.n100 185
R1035 VTAIL.n76 VTAIL.n75 185
R1036 VTAIL.n95 VTAIL.n94 185
R1037 VTAIL.n93 VTAIL.n92 185
R1038 VTAIL.n80 VTAIL.n79 185
R1039 VTAIL.n87 VTAIL.n86 185
R1040 VTAIL.n85 VTAIL.n84 185
R1041 VTAIL.n205 VTAIL.t2 149.524
R1042 VTAIL.n19 VTAIL.t1 149.524
R1043 VTAIL.n145 VTAIL.t0 149.524
R1044 VTAIL.n83 VTAIL.t3 149.524
R1045 VTAIL.n208 VTAIL.n207 104.615
R1046 VTAIL.n208 VTAIL.n201 104.615
R1047 VTAIL.n215 VTAIL.n201 104.615
R1048 VTAIL.n216 VTAIL.n215 104.615
R1049 VTAIL.n216 VTAIL.n197 104.615
R1050 VTAIL.n224 VTAIL.n197 104.615
R1051 VTAIL.n225 VTAIL.n224 104.615
R1052 VTAIL.n226 VTAIL.n225 104.615
R1053 VTAIL.n226 VTAIL.n193 104.615
R1054 VTAIL.n233 VTAIL.n193 104.615
R1055 VTAIL.n234 VTAIL.n233 104.615
R1056 VTAIL.n234 VTAIL.n189 104.615
R1057 VTAIL.n241 VTAIL.n189 104.615
R1058 VTAIL.n242 VTAIL.n241 104.615
R1059 VTAIL.n22 VTAIL.n21 104.615
R1060 VTAIL.n22 VTAIL.n15 104.615
R1061 VTAIL.n29 VTAIL.n15 104.615
R1062 VTAIL.n30 VTAIL.n29 104.615
R1063 VTAIL.n30 VTAIL.n11 104.615
R1064 VTAIL.n38 VTAIL.n11 104.615
R1065 VTAIL.n39 VTAIL.n38 104.615
R1066 VTAIL.n40 VTAIL.n39 104.615
R1067 VTAIL.n40 VTAIL.n7 104.615
R1068 VTAIL.n47 VTAIL.n7 104.615
R1069 VTAIL.n48 VTAIL.n47 104.615
R1070 VTAIL.n48 VTAIL.n3 104.615
R1071 VTAIL.n55 VTAIL.n3 104.615
R1072 VTAIL.n56 VTAIL.n55 104.615
R1073 VTAIL.n180 VTAIL.n179 104.615
R1074 VTAIL.n179 VTAIL.n127 104.615
R1075 VTAIL.n172 VTAIL.n127 104.615
R1076 VTAIL.n172 VTAIL.n171 104.615
R1077 VTAIL.n171 VTAIL.n131 104.615
R1078 VTAIL.n136 VTAIL.n131 104.615
R1079 VTAIL.n164 VTAIL.n136 104.615
R1080 VTAIL.n164 VTAIL.n163 104.615
R1081 VTAIL.n163 VTAIL.n137 104.615
R1082 VTAIL.n156 VTAIL.n137 104.615
R1083 VTAIL.n156 VTAIL.n155 104.615
R1084 VTAIL.n155 VTAIL.n141 104.615
R1085 VTAIL.n148 VTAIL.n141 104.615
R1086 VTAIL.n148 VTAIL.n147 104.615
R1087 VTAIL.n118 VTAIL.n117 104.615
R1088 VTAIL.n117 VTAIL.n65 104.615
R1089 VTAIL.n110 VTAIL.n65 104.615
R1090 VTAIL.n110 VTAIL.n109 104.615
R1091 VTAIL.n109 VTAIL.n69 104.615
R1092 VTAIL.n74 VTAIL.n69 104.615
R1093 VTAIL.n102 VTAIL.n74 104.615
R1094 VTAIL.n102 VTAIL.n101 104.615
R1095 VTAIL.n101 VTAIL.n75 104.615
R1096 VTAIL.n94 VTAIL.n75 104.615
R1097 VTAIL.n94 VTAIL.n93 104.615
R1098 VTAIL.n93 VTAIL.n79 104.615
R1099 VTAIL.n86 VTAIL.n79 104.615
R1100 VTAIL.n86 VTAIL.n85 104.615
R1101 VTAIL.n207 VTAIL.t2 52.3082
R1102 VTAIL.n21 VTAIL.t1 52.3082
R1103 VTAIL.n147 VTAIL.t0 52.3082
R1104 VTAIL.n85 VTAIL.t3 52.3082
R1105 VTAIL.n247 VTAIL.n246 31.6035
R1106 VTAIL.n61 VTAIL.n60 31.6035
R1107 VTAIL.n185 VTAIL.n184 31.6035
R1108 VTAIL.n123 VTAIL.n122 31.6035
R1109 VTAIL.n123 VTAIL.n61 23.4962
R1110 VTAIL.n247 VTAIL.n185 22.841
R1111 VTAIL.n227 VTAIL.n194 13.1884
R1112 VTAIL.n41 VTAIL.n8 13.1884
R1113 VTAIL.n134 VTAIL.n132 13.1884
R1114 VTAIL.n72 VTAIL.n70 13.1884
R1115 VTAIL.n228 VTAIL.n196 12.8005
R1116 VTAIL.n232 VTAIL.n231 12.8005
R1117 VTAIL.n42 VTAIL.n10 12.8005
R1118 VTAIL.n46 VTAIL.n45 12.8005
R1119 VTAIL.n170 VTAIL.n169 12.8005
R1120 VTAIL.n166 VTAIL.n165 12.8005
R1121 VTAIL.n108 VTAIL.n107 12.8005
R1122 VTAIL.n104 VTAIL.n103 12.8005
R1123 VTAIL.n223 VTAIL.n222 12.0247
R1124 VTAIL.n235 VTAIL.n192 12.0247
R1125 VTAIL.n37 VTAIL.n36 12.0247
R1126 VTAIL.n49 VTAIL.n6 12.0247
R1127 VTAIL.n173 VTAIL.n130 12.0247
R1128 VTAIL.n162 VTAIL.n135 12.0247
R1129 VTAIL.n111 VTAIL.n68 12.0247
R1130 VTAIL.n100 VTAIL.n73 12.0247
R1131 VTAIL.n221 VTAIL.n198 11.249
R1132 VTAIL.n236 VTAIL.n190 11.249
R1133 VTAIL.n35 VTAIL.n12 11.249
R1134 VTAIL.n50 VTAIL.n4 11.249
R1135 VTAIL.n174 VTAIL.n128 11.249
R1136 VTAIL.n161 VTAIL.n138 11.249
R1137 VTAIL.n112 VTAIL.n66 11.249
R1138 VTAIL.n99 VTAIL.n76 11.249
R1139 VTAIL.n218 VTAIL.n217 10.4732
R1140 VTAIL.n240 VTAIL.n239 10.4732
R1141 VTAIL.n32 VTAIL.n31 10.4732
R1142 VTAIL.n54 VTAIL.n53 10.4732
R1143 VTAIL.n178 VTAIL.n177 10.4732
R1144 VTAIL.n158 VTAIL.n157 10.4732
R1145 VTAIL.n116 VTAIL.n115 10.4732
R1146 VTAIL.n96 VTAIL.n95 10.4732
R1147 VTAIL.n206 VTAIL.n205 10.2747
R1148 VTAIL.n20 VTAIL.n19 10.2747
R1149 VTAIL.n146 VTAIL.n145 10.2747
R1150 VTAIL.n84 VTAIL.n83 10.2747
R1151 VTAIL.n214 VTAIL.n200 9.69747
R1152 VTAIL.n243 VTAIL.n188 9.69747
R1153 VTAIL.n28 VTAIL.n14 9.69747
R1154 VTAIL.n57 VTAIL.n2 9.69747
R1155 VTAIL.n181 VTAIL.n126 9.69747
R1156 VTAIL.n154 VTAIL.n140 9.69747
R1157 VTAIL.n119 VTAIL.n64 9.69747
R1158 VTAIL.n92 VTAIL.n78 9.69747
R1159 VTAIL.n246 VTAIL.n245 9.45567
R1160 VTAIL.n60 VTAIL.n59 9.45567
R1161 VTAIL.n184 VTAIL.n183 9.45567
R1162 VTAIL.n122 VTAIL.n121 9.45567
R1163 VTAIL.n245 VTAIL.n244 9.3005
R1164 VTAIL.n188 VTAIL.n187 9.3005
R1165 VTAIL.n239 VTAIL.n238 9.3005
R1166 VTAIL.n237 VTAIL.n236 9.3005
R1167 VTAIL.n192 VTAIL.n191 9.3005
R1168 VTAIL.n231 VTAIL.n230 9.3005
R1169 VTAIL.n204 VTAIL.n203 9.3005
R1170 VTAIL.n211 VTAIL.n210 9.3005
R1171 VTAIL.n213 VTAIL.n212 9.3005
R1172 VTAIL.n200 VTAIL.n199 9.3005
R1173 VTAIL.n219 VTAIL.n218 9.3005
R1174 VTAIL.n221 VTAIL.n220 9.3005
R1175 VTAIL.n222 VTAIL.n195 9.3005
R1176 VTAIL.n229 VTAIL.n228 9.3005
R1177 VTAIL.n59 VTAIL.n58 9.3005
R1178 VTAIL.n2 VTAIL.n1 9.3005
R1179 VTAIL.n53 VTAIL.n52 9.3005
R1180 VTAIL.n51 VTAIL.n50 9.3005
R1181 VTAIL.n6 VTAIL.n5 9.3005
R1182 VTAIL.n45 VTAIL.n44 9.3005
R1183 VTAIL.n18 VTAIL.n17 9.3005
R1184 VTAIL.n25 VTAIL.n24 9.3005
R1185 VTAIL.n27 VTAIL.n26 9.3005
R1186 VTAIL.n14 VTAIL.n13 9.3005
R1187 VTAIL.n33 VTAIL.n32 9.3005
R1188 VTAIL.n35 VTAIL.n34 9.3005
R1189 VTAIL.n36 VTAIL.n9 9.3005
R1190 VTAIL.n43 VTAIL.n42 9.3005
R1191 VTAIL.n144 VTAIL.n143 9.3005
R1192 VTAIL.n151 VTAIL.n150 9.3005
R1193 VTAIL.n153 VTAIL.n152 9.3005
R1194 VTAIL.n140 VTAIL.n139 9.3005
R1195 VTAIL.n159 VTAIL.n158 9.3005
R1196 VTAIL.n161 VTAIL.n160 9.3005
R1197 VTAIL.n135 VTAIL.n133 9.3005
R1198 VTAIL.n167 VTAIL.n166 9.3005
R1199 VTAIL.n183 VTAIL.n182 9.3005
R1200 VTAIL.n126 VTAIL.n125 9.3005
R1201 VTAIL.n177 VTAIL.n176 9.3005
R1202 VTAIL.n175 VTAIL.n174 9.3005
R1203 VTAIL.n130 VTAIL.n129 9.3005
R1204 VTAIL.n169 VTAIL.n168 9.3005
R1205 VTAIL.n82 VTAIL.n81 9.3005
R1206 VTAIL.n89 VTAIL.n88 9.3005
R1207 VTAIL.n91 VTAIL.n90 9.3005
R1208 VTAIL.n78 VTAIL.n77 9.3005
R1209 VTAIL.n97 VTAIL.n96 9.3005
R1210 VTAIL.n99 VTAIL.n98 9.3005
R1211 VTAIL.n73 VTAIL.n71 9.3005
R1212 VTAIL.n105 VTAIL.n104 9.3005
R1213 VTAIL.n121 VTAIL.n120 9.3005
R1214 VTAIL.n64 VTAIL.n63 9.3005
R1215 VTAIL.n115 VTAIL.n114 9.3005
R1216 VTAIL.n113 VTAIL.n112 9.3005
R1217 VTAIL.n68 VTAIL.n67 9.3005
R1218 VTAIL.n107 VTAIL.n106 9.3005
R1219 VTAIL.n213 VTAIL.n202 8.92171
R1220 VTAIL.n244 VTAIL.n186 8.92171
R1221 VTAIL.n27 VTAIL.n16 8.92171
R1222 VTAIL.n58 VTAIL.n0 8.92171
R1223 VTAIL.n182 VTAIL.n124 8.92171
R1224 VTAIL.n153 VTAIL.n142 8.92171
R1225 VTAIL.n120 VTAIL.n62 8.92171
R1226 VTAIL.n91 VTAIL.n80 8.92171
R1227 VTAIL.n210 VTAIL.n209 8.14595
R1228 VTAIL.n24 VTAIL.n23 8.14595
R1229 VTAIL.n150 VTAIL.n149 8.14595
R1230 VTAIL.n88 VTAIL.n87 8.14595
R1231 VTAIL.n206 VTAIL.n204 7.3702
R1232 VTAIL.n20 VTAIL.n18 7.3702
R1233 VTAIL.n146 VTAIL.n144 7.3702
R1234 VTAIL.n84 VTAIL.n82 7.3702
R1235 VTAIL.n209 VTAIL.n204 5.81868
R1236 VTAIL.n23 VTAIL.n18 5.81868
R1237 VTAIL.n149 VTAIL.n144 5.81868
R1238 VTAIL.n87 VTAIL.n82 5.81868
R1239 VTAIL.n210 VTAIL.n202 5.04292
R1240 VTAIL.n246 VTAIL.n186 5.04292
R1241 VTAIL.n24 VTAIL.n16 5.04292
R1242 VTAIL.n60 VTAIL.n0 5.04292
R1243 VTAIL.n184 VTAIL.n124 5.04292
R1244 VTAIL.n150 VTAIL.n142 5.04292
R1245 VTAIL.n122 VTAIL.n62 5.04292
R1246 VTAIL.n88 VTAIL.n80 5.04292
R1247 VTAIL.n214 VTAIL.n213 4.26717
R1248 VTAIL.n244 VTAIL.n243 4.26717
R1249 VTAIL.n28 VTAIL.n27 4.26717
R1250 VTAIL.n58 VTAIL.n57 4.26717
R1251 VTAIL.n182 VTAIL.n181 4.26717
R1252 VTAIL.n154 VTAIL.n153 4.26717
R1253 VTAIL.n120 VTAIL.n119 4.26717
R1254 VTAIL.n92 VTAIL.n91 4.26717
R1255 VTAIL.n217 VTAIL.n200 3.49141
R1256 VTAIL.n240 VTAIL.n188 3.49141
R1257 VTAIL.n31 VTAIL.n14 3.49141
R1258 VTAIL.n54 VTAIL.n2 3.49141
R1259 VTAIL.n178 VTAIL.n126 3.49141
R1260 VTAIL.n157 VTAIL.n140 3.49141
R1261 VTAIL.n116 VTAIL.n64 3.49141
R1262 VTAIL.n95 VTAIL.n78 3.49141
R1263 VTAIL.n205 VTAIL.n203 2.84303
R1264 VTAIL.n19 VTAIL.n17 2.84303
R1265 VTAIL.n145 VTAIL.n143 2.84303
R1266 VTAIL.n83 VTAIL.n81 2.84303
R1267 VTAIL.n218 VTAIL.n198 2.71565
R1268 VTAIL.n239 VTAIL.n190 2.71565
R1269 VTAIL.n32 VTAIL.n12 2.71565
R1270 VTAIL.n53 VTAIL.n4 2.71565
R1271 VTAIL.n177 VTAIL.n128 2.71565
R1272 VTAIL.n158 VTAIL.n138 2.71565
R1273 VTAIL.n115 VTAIL.n66 2.71565
R1274 VTAIL.n96 VTAIL.n76 2.71565
R1275 VTAIL.n223 VTAIL.n221 1.93989
R1276 VTAIL.n236 VTAIL.n235 1.93989
R1277 VTAIL.n37 VTAIL.n35 1.93989
R1278 VTAIL.n50 VTAIL.n49 1.93989
R1279 VTAIL.n174 VTAIL.n173 1.93989
R1280 VTAIL.n162 VTAIL.n161 1.93989
R1281 VTAIL.n112 VTAIL.n111 1.93989
R1282 VTAIL.n100 VTAIL.n99 1.93989
R1283 VTAIL.n222 VTAIL.n196 1.16414
R1284 VTAIL.n232 VTAIL.n192 1.16414
R1285 VTAIL.n36 VTAIL.n10 1.16414
R1286 VTAIL.n46 VTAIL.n6 1.16414
R1287 VTAIL.n170 VTAIL.n130 1.16414
R1288 VTAIL.n165 VTAIL.n135 1.16414
R1289 VTAIL.n108 VTAIL.n68 1.16414
R1290 VTAIL.n103 VTAIL.n73 1.16414
R1291 VTAIL.n185 VTAIL.n123 0.797914
R1292 VTAIL VTAIL.n61 0.69231
R1293 VTAIL.n228 VTAIL.n227 0.388379
R1294 VTAIL.n231 VTAIL.n194 0.388379
R1295 VTAIL.n42 VTAIL.n41 0.388379
R1296 VTAIL.n45 VTAIL.n8 0.388379
R1297 VTAIL.n169 VTAIL.n132 0.388379
R1298 VTAIL.n166 VTAIL.n134 0.388379
R1299 VTAIL.n107 VTAIL.n70 0.388379
R1300 VTAIL.n104 VTAIL.n72 0.388379
R1301 VTAIL.n211 VTAIL.n203 0.155672
R1302 VTAIL.n212 VTAIL.n211 0.155672
R1303 VTAIL.n212 VTAIL.n199 0.155672
R1304 VTAIL.n219 VTAIL.n199 0.155672
R1305 VTAIL.n220 VTAIL.n219 0.155672
R1306 VTAIL.n220 VTAIL.n195 0.155672
R1307 VTAIL.n229 VTAIL.n195 0.155672
R1308 VTAIL.n230 VTAIL.n229 0.155672
R1309 VTAIL.n230 VTAIL.n191 0.155672
R1310 VTAIL.n237 VTAIL.n191 0.155672
R1311 VTAIL.n238 VTAIL.n237 0.155672
R1312 VTAIL.n238 VTAIL.n187 0.155672
R1313 VTAIL.n245 VTAIL.n187 0.155672
R1314 VTAIL.n25 VTAIL.n17 0.155672
R1315 VTAIL.n26 VTAIL.n25 0.155672
R1316 VTAIL.n26 VTAIL.n13 0.155672
R1317 VTAIL.n33 VTAIL.n13 0.155672
R1318 VTAIL.n34 VTAIL.n33 0.155672
R1319 VTAIL.n34 VTAIL.n9 0.155672
R1320 VTAIL.n43 VTAIL.n9 0.155672
R1321 VTAIL.n44 VTAIL.n43 0.155672
R1322 VTAIL.n44 VTAIL.n5 0.155672
R1323 VTAIL.n51 VTAIL.n5 0.155672
R1324 VTAIL.n52 VTAIL.n51 0.155672
R1325 VTAIL.n52 VTAIL.n1 0.155672
R1326 VTAIL.n59 VTAIL.n1 0.155672
R1327 VTAIL.n183 VTAIL.n125 0.155672
R1328 VTAIL.n176 VTAIL.n125 0.155672
R1329 VTAIL.n176 VTAIL.n175 0.155672
R1330 VTAIL.n175 VTAIL.n129 0.155672
R1331 VTAIL.n168 VTAIL.n129 0.155672
R1332 VTAIL.n168 VTAIL.n167 0.155672
R1333 VTAIL.n167 VTAIL.n133 0.155672
R1334 VTAIL.n160 VTAIL.n133 0.155672
R1335 VTAIL.n160 VTAIL.n159 0.155672
R1336 VTAIL.n159 VTAIL.n139 0.155672
R1337 VTAIL.n152 VTAIL.n139 0.155672
R1338 VTAIL.n152 VTAIL.n151 0.155672
R1339 VTAIL.n151 VTAIL.n143 0.155672
R1340 VTAIL.n121 VTAIL.n63 0.155672
R1341 VTAIL.n114 VTAIL.n63 0.155672
R1342 VTAIL.n114 VTAIL.n113 0.155672
R1343 VTAIL.n113 VTAIL.n67 0.155672
R1344 VTAIL.n106 VTAIL.n67 0.155672
R1345 VTAIL.n106 VTAIL.n105 0.155672
R1346 VTAIL.n105 VTAIL.n71 0.155672
R1347 VTAIL.n98 VTAIL.n71 0.155672
R1348 VTAIL.n98 VTAIL.n97 0.155672
R1349 VTAIL.n97 VTAIL.n77 0.155672
R1350 VTAIL.n90 VTAIL.n77 0.155672
R1351 VTAIL.n90 VTAIL.n89 0.155672
R1352 VTAIL.n89 VTAIL.n81 0.155672
R1353 VTAIL VTAIL.n247 0.106103
R1354 VDD2.n117 VDD2.n61 289.615
R1355 VDD2.n56 VDD2.n0 289.615
R1356 VDD2.n118 VDD2.n117 185
R1357 VDD2.n116 VDD2.n115 185
R1358 VDD2.n65 VDD2.n64 185
R1359 VDD2.n110 VDD2.n109 185
R1360 VDD2.n108 VDD2.n107 185
R1361 VDD2.n69 VDD2.n68 185
R1362 VDD2.n73 VDD2.n71 185
R1363 VDD2.n102 VDD2.n101 185
R1364 VDD2.n100 VDD2.n99 185
R1365 VDD2.n75 VDD2.n74 185
R1366 VDD2.n94 VDD2.n93 185
R1367 VDD2.n92 VDD2.n91 185
R1368 VDD2.n79 VDD2.n78 185
R1369 VDD2.n86 VDD2.n85 185
R1370 VDD2.n84 VDD2.n83 185
R1371 VDD2.n21 VDD2.n20 185
R1372 VDD2.n23 VDD2.n22 185
R1373 VDD2.n16 VDD2.n15 185
R1374 VDD2.n29 VDD2.n28 185
R1375 VDD2.n31 VDD2.n30 185
R1376 VDD2.n12 VDD2.n11 185
R1377 VDD2.n38 VDD2.n37 185
R1378 VDD2.n39 VDD2.n10 185
R1379 VDD2.n41 VDD2.n40 185
R1380 VDD2.n8 VDD2.n7 185
R1381 VDD2.n47 VDD2.n46 185
R1382 VDD2.n49 VDD2.n48 185
R1383 VDD2.n4 VDD2.n3 185
R1384 VDD2.n55 VDD2.n54 185
R1385 VDD2.n57 VDD2.n56 185
R1386 VDD2.n82 VDD2.t1 149.524
R1387 VDD2.n19 VDD2.t0 149.524
R1388 VDD2.n117 VDD2.n116 104.615
R1389 VDD2.n116 VDD2.n64 104.615
R1390 VDD2.n109 VDD2.n64 104.615
R1391 VDD2.n109 VDD2.n108 104.615
R1392 VDD2.n108 VDD2.n68 104.615
R1393 VDD2.n73 VDD2.n68 104.615
R1394 VDD2.n101 VDD2.n73 104.615
R1395 VDD2.n101 VDD2.n100 104.615
R1396 VDD2.n100 VDD2.n74 104.615
R1397 VDD2.n93 VDD2.n74 104.615
R1398 VDD2.n93 VDD2.n92 104.615
R1399 VDD2.n92 VDD2.n78 104.615
R1400 VDD2.n85 VDD2.n78 104.615
R1401 VDD2.n85 VDD2.n84 104.615
R1402 VDD2.n22 VDD2.n21 104.615
R1403 VDD2.n22 VDD2.n15 104.615
R1404 VDD2.n29 VDD2.n15 104.615
R1405 VDD2.n30 VDD2.n29 104.615
R1406 VDD2.n30 VDD2.n11 104.615
R1407 VDD2.n38 VDD2.n11 104.615
R1408 VDD2.n39 VDD2.n38 104.615
R1409 VDD2.n40 VDD2.n39 104.615
R1410 VDD2.n40 VDD2.n7 104.615
R1411 VDD2.n47 VDD2.n7 104.615
R1412 VDD2.n48 VDD2.n47 104.615
R1413 VDD2.n48 VDD2.n3 104.615
R1414 VDD2.n55 VDD2.n3 104.615
R1415 VDD2.n56 VDD2.n55 104.615
R1416 VDD2.n122 VDD2.n60 83.0711
R1417 VDD2.n84 VDD2.t1 52.3082
R1418 VDD2.n21 VDD2.t0 52.3082
R1419 VDD2.n122 VDD2.n121 48.2823
R1420 VDD2.n71 VDD2.n69 13.1884
R1421 VDD2.n41 VDD2.n8 13.1884
R1422 VDD2.n107 VDD2.n106 12.8005
R1423 VDD2.n103 VDD2.n102 12.8005
R1424 VDD2.n42 VDD2.n10 12.8005
R1425 VDD2.n46 VDD2.n45 12.8005
R1426 VDD2.n110 VDD2.n67 12.0247
R1427 VDD2.n99 VDD2.n72 12.0247
R1428 VDD2.n37 VDD2.n36 12.0247
R1429 VDD2.n49 VDD2.n6 12.0247
R1430 VDD2.n111 VDD2.n65 11.249
R1431 VDD2.n98 VDD2.n75 11.249
R1432 VDD2.n35 VDD2.n12 11.249
R1433 VDD2.n50 VDD2.n4 11.249
R1434 VDD2.n115 VDD2.n114 10.4732
R1435 VDD2.n95 VDD2.n94 10.4732
R1436 VDD2.n32 VDD2.n31 10.4732
R1437 VDD2.n54 VDD2.n53 10.4732
R1438 VDD2.n83 VDD2.n82 10.2747
R1439 VDD2.n20 VDD2.n19 10.2747
R1440 VDD2.n118 VDD2.n63 9.69747
R1441 VDD2.n91 VDD2.n77 9.69747
R1442 VDD2.n28 VDD2.n14 9.69747
R1443 VDD2.n57 VDD2.n2 9.69747
R1444 VDD2.n121 VDD2.n120 9.45567
R1445 VDD2.n60 VDD2.n59 9.45567
R1446 VDD2.n81 VDD2.n80 9.3005
R1447 VDD2.n88 VDD2.n87 9.3005
R1448 VDD2.n90 VDD2.n89 9.3005
R1449 VDD2.n77 VDD2.n76 9.3005
R1450 VDD2.n96 VDD2.n95 9.3005
R1451 VDD2.n98 VDD2.n97 9.3005
R1452 VDD2.n72 VDD2.n70 9.3005
R1453 VDD2.n104 VDD2.n103 9.3005
R1454 VDD2.n120 VDD2.n119 9.3005
R1455 VDD2.n63 VDD2.n62 9.3005
R1456 VDD2.n114 VDD2.n113 9.3005
R1457 VDD2.n112 VDD2.n111 9.3005
R1458 VDD2.n67 VDD2.n66 9.3005
R1459 VDD2.n106 VDD2.n105 9.3005
R1460 VDD2.n59 VDD2.n58 9.3005
R1461 VDD2.n2 VDD2.n1 9.3005
R1462 VDD2.n53 VDD2.n52 9.3005
R1463 VDD2.n51 VDD2.n50 9.3005
R1464 VDD2.n6 VDD2.n5 9.3005
R1465 VDD2.n45 VDD2.n44 9.3005
R1466 VDD2.n18 VDD2.n17 9.3005
R1467 VDD2.n25 VDD2.n24 9.3005
R1468 VDD2.n27 VDD2.n26 9.3005
R1469 VDD2.n14 VDD2.n13 9.3005
R1470 VDD2.n33 VDD2.n32 9.3005
R1471 VDD2.n35 VDD2.n34 9.3005
R1472 VDD2.n36 VDD2.n9 9.3005
R1473 VDD2.n43 VDD2.n42 9.3005
R1474 VDD2.n119 VDD2.n61 8.92171
R1475 VDD2.n90 VDD2.n79 8.92171
R1476 VDD2.n27 VDD2.n16 8.92171
R1477 VDD2.n58 VDD2.n0 8.92171
R1478 VDD2.n87 VDD2.n86 8.14595
R1479 VDD2.n24 VDD2.n23 8.14595
R1480 VDD2.n83 VDD2.n81 7.3702
R1481 VDD2.n20 VDD2.n18 7.3702
R1482 VDD2.n86 VDD2.n81 5.81868
R1483 VDD2.n23 VDD2.n18 5.81868
R1484 VDD2.n121 VDD2.n61 5.04292
R1485 VDD2.n87 VDD2.n79 5.04292
R1486 VDD2.n24 VDD2.n16 5.04292
R1487 VDD2.n60 VDD2.n0 5.04292
R1488 VDD2.n119 VDD2.n118 4.26717
R1489 VDD2.n91 VDD2.n90 4.26717
R1490 VDD2.n28 VDD2.n27 4.26717
R1491 VDD2.n58 VDD2.n57 4.26717
R1492 VDD2.n115 VDD2.n63 3.49141
R1493 VDD2.n94 VDD2.n77 3.49141
R1494 VDD2.n31 VDD2.n14 3.49141
R1495 VDD2.n54 VDD2.n2 3.49141
R1496 VDD2.n82 VDD2.n80 2.84303
R1497 VDD2.n19 VDD2.n17 2.84303
R1498 VDD2.n114 VDD2.n65 2.71565
R1499 VDD2.n95 VDD2.n75 2.71565
R1500 VDD2.n32 VDD2.n12 2.71565
R1501 VDD2.n53 VDD2.n4 2.71565
R1502 VDD2.n111 VDD2.n110 1.93989
R1503 VDD2.n99 VDD2.n98 1.93989
R1504 VDD2.n37 VDD2.n35 1.93989
R1505 VDD2.n50 VDD2.n49 1.93989
R1506 VDD2.n107 VDD2.n67 1.16414
R1507 VDD2.n102 VDD2.n72 1.16414
R1508 VDD2.n36 VDD2.n10 1.16414
R1509 VDD2.n46 VDD2.n6 1.16414
R1510 VDD2.n106 VDD2.n69 0.388379
R1511 VDD2.n103 VDD2.n71 0.388379
R1512 VDD2.n42 VDD2.n41 0.388379
R1513 VDD2.n45 VDD2.n8 0.388379
R1514 VDD2 VDD2.n122 0.222483
R1515 VDD2.n120 VDD2.n62 0.155672
R1516 VDD2.n113 VDD2.n62 0.155672
R1517 VDD2.n113 VDD2.n112 0.155672
R1518 VDD2.n112 VDD2.n66 0.155672
R1519 VDD2.n105 VDD2.n66 0.155672
R1520 VDD2.n105 VDD2.n104 0.155672
R1521 VDD2.n104 VDD2.n70 0.155672
R1522 VDD2.n97 VDD2.n70 0.155672
R1523 VDD2.n97 VDD2.n96 0.155672
R1524 VDD2.n96 VDD2.n76 0.155672
R1525 VDD2.n89 VDD2.n76 0.155672
R1526 VDD2.n89 VDD2.n88 0.155672
R1527 VDD2.n88 VDD2.n80 0.155672
R1528 VDD2.n25 VDD2.n17 0.155672
R1529 VDD2.n26 VDD2.n25 0.155672
R1530 VDD2.n26 VDD2.n13 0.155672
R1531 VDD2.n33 VDD2.n13 0.155672
R1532 VDD2.n34 VDD2.n33 0.155672
R1533 VDD2.n34 VDD2.n9 0.155672
R1534 VDD2.n43 VDD2.n9 0.155672
R1535 VDD2.n44 VDD2.n43 0.155672
R1536 VDD2.n44 VDD2.n5 0.155672
R1537 VDD2.n51 VDD2.n5 0.155672
R1538 VDD2.n52 VDD2.n51 0.155672
R1539 VDD2.n52 VDD2.n1 0.155672
R1540 VDD2.n59 VDD2.n1 0.155672
R1541 VP.n0 VP.t1 928.904
R1542 VP.n0 VP.t0 890.466
R1543 VP VP.n0 0.0516364
R1544 VDD1.n56 VDD1.n0 289.615
R1545 VDD1.n117 VDD1.n61 289.615
R1546 VDD1.n57 VDD1.n56 185
R1547 VDD1.n55 VDD1.n54 185
R1548 VDD1.n4 VDD1.n3 185
R1549 VDD1.n49 VDD1.n48 185
R1550 VDD1.n47 VDD1.n46 185
R1551 VDD1.n8 VDD1.n7 185
R1552 VDD1.n12 VDD1.n10 185
R1553 VDD1.n41 VDD1.n40 185
R1554 VDD1.n39 VDD1.n38 185
R1555 VDD1.n14 VDD1.n13 185
R1556 VDD1.n33 VDD1.n32 185
R1557 VDD1.n31 VDD1.n30 185
R1558 VDD1.n18 VDD1.n17 185
R1559 VDD1.n25 VDD1.n24 185
R1560 VDD1.n23 VDD1.n22 185
R1561 VDD1.n82 VDD1.n81 185
R1562 VDD1.n84 VDD1.n83 185
R1563 VDD1.n77 VDD1.n76 185
R1564 VDD1.n90 VDD1.n89 185
R1565 VDD1.n92 VDD1.n91 185
R1566 VDD1.n73 VDD1.n72 185
R1567 VDD1.n99 VDD1.n98 185
R1568 VDD1.n100 VDD1.n71 185
R1569 VDD1.n102 VDD1.n101 185
R1570 VDD1.n69 VDD1.n68 185
R1571 VDD1.n108 VDD1.n107 185
R1572 VDD1.n110 VDD1.n109 185
R1573 VDD1.n65 VDD1.n64 185
R1574 VDD1.n116 VDD1.n115 185
R1575 VDD1.n118 VDD1.n117 185
R1576 VDD1.n21 VDD1.t0 149.524
R1577 VDD1.n80 VDD1.t1 149.524
R1578 VDD1.n56 VDD1.n55 104.615
R1579 VDD1.n55 VDD1.n3 104.615
R1580 VDD1.n48 VDD1.n3 104.615
R1581 VDD1.n48 VDD1.n47 104.615
R1582 VDD1.n47 VDD1.n7 104.615
R1583 VDD1.n12 VDD1.n7 104.615
R1584 VDD1.n40 VDD1.n12 104.615
R1585 VDD1.n40 VDD1.n39 104.615
R1586 VDD1.n39 VDD1.n13 104.615
R1587 VDD1.n32 VDD1.n13 104.615
R1588 VDD1.n32 VDD1.n31 104.615
R1589 VDD1.n31 VDD1.n17 104.615
R1590 VDD1.n24 VDD1.n17 104.615
R1591 VDD1.n24 VDD1.n23 104.615
R1592 VDD1.n83 VDD1.n82 104.615
R1593 VDD1.n83 VDD1.n76 104.615
R1594 VDD1.n90 VDD1.n76 104.615
R1595 VDD1.n91 VDD1.n90 104.615
R1596 VDD1.n91 VDD1.n72 104.615
R1597 VDD1.n99 VDD1.n72 104.615
R1598 VDD1.n100 VDD1.n99 104.615
R1599 VDD1.n101 VDD1.n100 104.615
R1600 VDD1.n101 VDD1.n68 104.615
R1601 VDD1.n108 VDD1.n68 104.615
R1602 VDD1.n109 VDD1.n108 104.615
R1603 VDD1.n109 VDD1.n64 104.615
R1604 VDD1.n116 VDD1.n64 104.615
R1605 VDD1.n117 VDD1.n116 104.615
R1606 VDD1 VDD1.n121 83.7597
R1607 VDD1.n23 VDD1.t0 52.3082
R1608 VDD1.n82 VDD1.t1 52.3082
R1609 VDD1 VDD1.n60 48.5043
R1610 VDD1.n10 VDD1.n8 13.1884
R1611 VDD1.n102 VDD1.n69 13.1884
R1612 VDD1.n46 VDD1.n45 12.8005
R1613 VDD1.n42 VDD1.n41 12.8005
R1614 VDD1.n103 VDD1.n71 12.8005
R1615 VDD1.n107 VDD1.n106 12.8005
R1616 VDD1.n49 VDD1.n6 12.0247
R1617 VDD1.n38 VDD1.n11 12.0247
R1618 VDD1.n98 VDD1.n97 12.0247
R1619 VDD1.n110 VDD1.n67 12.0247
R1620 VDD1.n50 VDD1.n4 11.249
R1621 VDD1.n37 VDD1.n14 11.249
R1622 VDD1.n96 VDD1.n73 11.249
R1623 VDD1.n111 VDD1.n65 11.249
R1624 VDD1.n54 VDD1.n53 10.4732
R1625 VDD1.n34 VDD1.n33 10.4732
R1626 VDD1.n93 VDD1.n92 10.4732
R1627 VDD1.n115 VDD1.n114 10.4732
R1628 VDD1.n22 VDD1.n21 10.2747
R1629 VDD1.n81 VDD1.n80 10.2747
R1630 VDD1.n57 VDD1.n2 9.69747
R1631 VDD1.n30 VDD1.n16 9.69747
R1632 VDD1.n89 VDD1.n75 9.69747
R1633 VDD1.n118 VDD1.n63 9.69747
R1634 VDD1.n60 VDD1.n59 9.45567
R1635 VDD1.n121 VDD1.n120 9.45567
R1636 VDD1.n20 VDD1.n19 9.3005
R1637 VDD1.n27 VDD1.n26 9.3005
R1638 VDD1.n29 VDD1.n28 9.3005
R1639 VDD1.n16 VDD1.n15 9.3005
R1640 VDD1.n35 VDD1.n34 9.3005
R1641 VDD1.n37 VDD1.n36 9.3005
R1642 VDD1.n11 VDD1.n9 9.3005
R1643 VDD1.n43 VDD1.n42 9.3005
R1644 VDD1.n59 VDD1.n58 9.3005
R1645 VDD1.n2 VDD1.n1 9.3005
R1646 VDD1.n53 VDD1.n52 9.3005
R1647 VDD1.n51 VDD1.n50 9.3005
R1648 VDD1.n6 VDD1.n5 9.3005
R1649 VDD1.n45 VDD1.n44 9.3005
R1650 VDD1.n120 VDD1.n119 9.3005
R1651 VDD1.n63 VDD1.n62 9.3005
R1652 VDD1.n114 VDD1.n113 9.3005
R1653 VDD1.n112 VDD1.n111 9.3005
R1654 VDD1.n67 VDD1.n66 9.3005
R1655 VDD1.n106 VDD1.n105 9.3005
R1656 VDD1.n79 VDD1.n78 9.3005
R1657 VDD1.n86 VDD1.n85 9.3005
R1658 VDD1.n88 VDD1.n87 9.3005
R1659 VDD1.n75 VDD1.n74 9.3005
R1660 VDD1.n94 VDD1.n93 9.3005
R1661 VDD1.n96 VDD1.n95 9.3005
R1662 VDD1.n97 VDD1.n70 9.3005
R1663 VDD1.n104 VDD1.n103 9.3005
R1664 VDD1.n58 VDD1.n0 8.92171
R1665 VDD1.n29 VDD1.n18 8.92171
R1666 VDD1.n88 VDD1.n77 8.92171
R1667 VDD1.n119 VDD1.n61 8.92171
R1668 VDD1.n26 VDD1.n25 8.14595
R1669 VDD1.n85 VDD1.n84 8.14595
R1670 VDD1.n22 VDD1.n20 7.3702
R1671 VDD1.n81 VDD1.n79 7.3702
R1672 VDD1.n25 VDD1.n20 5.81868
R1673 VDD1.n84 VDD1.n79 5.81868
R1674 VDD1.n60 VDD1.n0 5.04292
R1675 VDD1.n26 VDD1.n18 5.04292
R1676 VDD1.n85 VDD1.n77 5.04292
R1677 VDD1.n121 VDD1.n61 5.04292
R1678 VDD1.n58 VDD1.n57 4.26717
R1679 VDD1.n30 VDD1.n29 4.26717
R1680 VDD1.n89 VDD1.n88 4.26717
R1681 VDD1.n119 VDD1.n118 4.26717
R1682 VDD1.n54 VDD1.n2 3.49141
R1683 VDD1.n33 VDD1.n16 3.49141
R1684 VDD1.n92 VDD1.n75 3.49141
R1685 VDD1.n115 VDD1.n63 3.49141
R1686 VDD1.n21 VDD1.n19 2.84303
R1687 VDD1.n80 VDD1.n78 2.84303
R1688 VDD1.n53 VDD1.n4 2.71565
R1689 VDD1.n34 VDD1.n14 2.71565
R1690 VDD1.n93 VDD1.n73 2.71565
R1691 VDD1.n114 VDD1.n65 2.71565
R1692 VDD1.n50 VDD1.n49 1.93989
R1693 VDD1.n38 VDD1.n37 1.93989
R1694 VDD1.n98 VDD1.n96 1.93989
R1695 VDD1.n111 VDD1.n110 1.93989
R1696 VDD1.n46 VDD1.n6 1.16414
R1697 VDD1.n41 VDD1.n11 1.16414
R1698 VDD1.n97 VDD1.n71 1.16414
R1699 VDD1.n107 VDD1.n67 1.16414
R1700 VDD1.n45 VDD1.n8 0.388379
R1701 VDD1.n42 VDD1.n10 0.388379
R1702 VDD1.n103 VDD1.n102 0.388379
R1703 VDD1.n106 VDD1.n69 0.388379
R1704 VDD1.n59 VDD1.n1 0.155672
R1705 VDD1.n52 VDD1.n1 0.155672
R1706 VDD1.n52 VDD1.n51 0.155672
R1707 VDD1.n51 VDD1.n5 0.155672
R1708 VDD1.n44 VDD1.n5 0.155672
R1709 VDD1.n44 VDD1.n43 0.155672
R1710 VDD1.n43 VDD1.n9 0.155672
R1711 VDD1.n36 VDD1.n9 0.155672
R1712 VDD1.n36 VDD1.n35 0.155672
R1713 VDD1.n35 VDD1.n15 0.155672
R1714 VDD1.n28 VDD1.n15 0.155672
R1715 VDD1.n28 VDD1.n27 0.155672
R1716 VDD1.n27 VDD1.n19 0.155672
R1717 VDD1.n86 VDD1.n78 0.155672
R1718 VDD1.n87 VDD1.n86 0.155672
R1719 VDD1.n87 VDD1.n74 0.155672
R1720 VDD1.n94 VDD1.n74 0.155672
R1721 VDD1.n95 VDD1.n94 0.155672
R1722 VDD1.n95 VDD1.n70 0.155672
R1723 VDD1.n104 VDD1.n70 0.155672
R1724 VDD1.n105 VDD1.n104 0.155672
R1725 VDD1.n105 VDD1.n66 0.155672
R1726 VDD1.n112 VDD1.n66 0.155672
R1727 VDD1.n113 VDD1.n112 0.155672
R1728 VDD1.n113 VDD1.n62 0.155672
R1729 VDD1.n120 VDD1.n62 0.155672
C0 VP VN 4.32292f
C1 VDD2 VTAIL 6.09746f
C2 VP VDD1 1.66926f
C3 VN VTAIL 1.0516f
C4 VN VDD2 1.57861f
C5 VDD1 VTAIL 6.06622f
C6 VP VTAIL 1.06628f
C7 VDD1 VDD2 0.437386f
C8 VP VDD2 0.243699f
C9 VN VDD1 0.148466f
C10 VDD2 B 3.534746f
C11 VDD1 B 5.47736f
C12 VTAIL B 5.544043f
C13 VN B 6.833549f
C14 VP B 3.659746f
C15 VDD1.n0 B 0.023619f
C16 VDD1.n1 B 0.017388f
C17 VDD1.n2 B 0.009343f
C18 VDD1.n3 B 0.022084f
C19 VDD1.n4 B 0.009893f
C20 VDD1.n5 B 0.017388f
C21 VDD1.n6 B 0.009343f
C22 VDD1.n7 B 0.022084f
C23 VDD1.n8 B 0.009618f
C24 VDD1.n9 B 0.017388f
C25 VDD1.n10 B 0.009618f
C26 VDD1.n11 B 0.009343f
C27 VDD1.n12 B 0.022084f
C28 VDD1.n13 B 0.022084f
C29 VDD1.n14 B 0.009893f
C30 VDD1.n15 B 0.017388f
C31 VDD1.n16 B 0.009343f
C32 VDD1.n17 B 0.022084f
C33 VDD1.n18 B 0.009893f
C34 VDD1.n19 B 0.828456f
C35 VDD1.n20 B 0.009343f
C36 VDD1.t0 B 0.03724f
C37 VDD1.n21 B 0.121158f
C38 VDD1.n22 B 0.015612f
C39 VDD1.n23 B 0.016563f
C40 VDD1.n24 B 0.022084f
C41 VDD1.n25 B 0.009893f
C42 VDD1.n26 B 0.009343f
C43 VDD1.n27 B 0.017388f
C44 VDD1.n28 B 0.017388f
C45 VDD1.n29 B 0.009343f
C46 VDD1.n30 B 0.009893f
C47 VDD1.n31 B 0.022084f
C48 VDD1.n32 B 0.022084f
C49 VDD1.n33 B 0.009893f
C50 VDD1.n34 B 0.009343f
C51 VDD1.n35 B 0.017388f
C52 VDD1.n36 B 0.017388f
C53 VDD1.n37 B 0.009343f
C54 VDD1.n38 B 0.009893f
C55 VDD1.n39 B 0.022084f
C56 VDD1.n40 B 0.022084f
C57 VDD1.n41 B 0.009893f
C58 VDD1.n42 B 0.009343f
C59 VDD1.n43 B 0.017388f
C60 VDD1.n44 B 0.017388f
C61 VDD1.n45 B 0.009343f
C62 VDD1.n46 B 0.009893f
C63 VDD1.n47 B 0.022084f
C64 VDD1.n48 B 0.022084f
C65 VDD1.n49 B 0.009893f
C66 VDD1.n50 B 0.009343f
C67 VDD1.n51 B 0.017388f
C68 VDD1.n52 B 0.017388f
C69 VDD1.n53 B 0.009343f
C70 VDD1.n54 B 0.009893f
C71 VDD1.n55 B 0.022084f
C72 VDD1.n56 B 0.046357f
C73 VDD1.n57 B 0.009893f
C74 VDD1.n58 B 0.009343f
C75 VDD1.n59 B 0.039478f
C76 VDD1.n60 B 0.037987f
C77 VDD1.n61 B 0.023619f
C78 VDD1.n62 B 0.017388f
C79 VDD1.n63 B 0.009343f
C80 VDD1.n64 B 0.022084f
C81 VDD1.n65 B 0.009893f
C82 VDD1.n66 B 0.017388f
C83 VDD1.n67 B 0.009343f
C84 VDD1.n68 B 0.022084f
C85 VDD1.n69 B 0.009618f
C86 VDD1.n70 B 0.017388f
C87 VDD1.n71 B 0.009893f
C88 VDD1.n72 B 0.022084f
C89 VDD1.n73 B 0.009893f
C90 VDD1.n74 B 0.017388f
C91 VDD1.n75 B 0.009343f
C92 VDD1.n76 B 0.022084f
C93 VDD1.n77 B 0.009893f
C94 VDD1.n78 B 0.828456f
C95 VDD1.n79 B 0.009343f
C96 VDD1.t1 B 0.03724f
C97 VDD1.n80 B 0.121158f
C98 VDD1.n81 B 0.015612f
C99 VDD1.n82 B 0.016563f
C100 VDD1.n83 B 0.022084f
C101 VDD1.n84 B 0.009893f
C102 VDD1.n85 B 0.009343f
C103 VDD1.n86 B 0.017388f
C104 VDD1.n87 B 0.017388f
C105 VDD1.n88 B 0.009343f
C106 VDD1.n89 B 0.009893f
C107 VDD1.n90 B 0.022084f
C108 VDD1.n91 B 0.022084f
C109 VDD1.n92 B 0.009893f
C110 VDD1.n93 B 0.009343f
C111 VDD1.n94 B 0.017388f
C112 VDD1.n95 B 0.017388f
C113 VDD1.n96 B 0.009343f
C114 VDD1.n97 B 0.009343f
C115 VDD1.n98 B 0.009893f
C116 VDD1.n99 B 0.022084f
C117 VDD1.n100 B 0.022084f
C118 VDD1.n101 B 0.022084f
C119 VDD1.n102 B 0.009618f
C120 VDD1.n103 B 0.009343f
C121 VDD1.n104 B 0.017388f
C122 VDD1.n105 B 0.017388f
C123 VDD1.n106 B 0.009343f
C124 VDD1.n107 B 0.009893f
C125 VDD1.n108 B 0.022084f
C126 VDD1.n109 B 0.022084f
C127 VDD1.n110 B 0.009893f
C128 VDD1.n111 B 0.009343f
C129 VDD1.n112 B 0.017388f
C130 VDD1.n113 B 0.017388f
C131 VDD1.n114 B 0.009343f
C132 VDD1.n115 B 0.009893f
C133 VDD1.n116 B 0.022084f
C134 VDD1.n117 B 0.046357f
C135 VDD1.n118 B 0.009893f
C136 VDD1.n119 B 0.009343f
C137 VDD1.n120 B 0.039478f
C138 VDD1.n121 B 0.424301f
C139 VP.t1 B 0.645272f
C140 VP.t0 B 0.58111f
C141 VP.n0 B 3.06655f
C142 VDD2.n0 B 0.02387f
C143 VDD2.n1 B 0.017573f
C144 VDD2.n2 B 0.009443f
C145 VDD2.n3 B 0.022319f
C146 VDD2.n4 B 0.009998f
C147 VDD2.n5 B 0.017573f
C148 VDD2.n6 B 0.009443f
C149 VDD2.n7 B 0.022319f
C150 VDD2.n8 B 0.009721f
C151 VDD2.n9 B 0.017573f
C152 VDD2.n10 B 0.009998f
C153 VDD2.n11 B 0.022319f
C154 VDD2.n12 B 0.009998f
C155 VDD2.n13 B 0.017573f
C156 VDD2.n14 B 0.009443f
C157 VDD2.n15 B 0.022319f
C158 VDD2.n16 B 0.009998f
C159 VDD2.n17 B 0.83727f
C160 VDD2.n18 B 0.009443f
C161 VDD2.t0 B 0.037637f
C162 VDD2.n19 B 0.122447f
C163 VDD2.n20 B 0.015778f
C164 VDD2.n21 B 0.01674f
C165 VDD2.n22 B 0.022319f
C166 VDD2.n23 B 0.009998f
C167 VDD2.n24 B 0.009443f
C168 VDD2.n25 B 0.017573f
C169 VDD2.n26 B 0.017573f
C170 VDD2.n27 B 0.009443f
C171 VDD2.n28 B 0.009998f
C172 VDD2.n29 B 0.022319f
C173 VDD2.n30 B 0.022319f
C174 VDD2.n31 B 0.009998f
C175 VDD2.n32 B 0.009443f
C176 VDD2.n33 B 0.017573f
C177 VDD2.n34 B 0.017573f
C178 VDD2.n35 B 0.009443f
C179 VDD2.n36 B 0.009443f
C180 VDD2.n37 B 0.009998f
C181 VDD2.n38 B 0.022319f
C182 VDD2.n39 B 0.022319f
C183 VDD2.n40 B 0.022319f
C184 VDD2.n41 B 0.009721f
C185 VDD2.n42 B 0.009443f
C186 VDD2.n43 B 0.017573f
C187 VDD2.n44 B 0.017573f
C188 VDD2.n45 B 0.009443f
C189 VDD2.n46 B 0.009998f
C190 VDD2.n47 B 0.022319f
C191 VDD2.n48 B 0.022319f
C192 VDD2.n49 B 0.009998f
C193 VDD2.n50 B 0.009443f
C194 VDD2.n51 B 0.017573f
C195 VDD2.n52 B 0.017573f
C196 VDD2.n53 B 0.009443f
C197 VDD2.n54 B 0.009998f
C198 VDD2.n55 B 0.022319f
C199 VDD2.n56 B 0.04685f
C200 VDD2.n57 B 0.009998f
C201 VDD2.n58 B 0.009443f
C202 VDD2.n59 B 0.039898f
C203 VDD2.n60 B 0.406929f
C204 VDD2.n61 B 0.02387f
C205 VDD2.n62 B 0.017573f
C206 VDD2.n63 B 0.009443f
C207 VDD2.n64 B 0.022319f
C208 VDD2.n65 B 0.009998f
C209 VDD2.n66 B 0.017573f
C210 VDD2.n67 B 0.009443f
C211 VDD2.n68 B 0.022319f
C212 VDD2.n69 B 0.009721f
C213 VDD2.n70 B 0.017573f
C214 VDD2.n71 B 0.009721f
C215 VDD2.n72 B 0.009443f
C216 VDD2.n73 B 0.022319f
C217 VDD2.n74 B 0.022319f
C218 VDD2.n75 B 0.009998f
C219 VDD2.n76 B 0.017573f
C220 VDD2.n77 B 0.009443f
C221 VDD2.n78 B 0.022319f
C222 VDD2.n79 B 0.009998f
C223 VDD2.n80 B 0.83727f
C224 VDD2.n81 B 0.009443f
C225 VDD2.t1 B 0.037637f
C226 VDD2.n82 B 0.122447f
C227 VDD2.n83 B 0.015778f
C228 VDD2.n84 B 0.01674f
C229 VDD2.n85 B 0.022319f
C230 VDD2.n86 B 0.009998f
C231 VDD2.n87 B 0.009443f
C232 VDD2.n88 B 0.017573f
C233 VDD2.n89 B 0.017573f
C234 VDD2.n90 B 0.009443f
C235 VDD2.n91 B 0.009998f
C236 VDD2.n92 B 0.022319f
C237 VDD2.n93 B 0.022319f
C238 VDD2.n94 B 0.009998f
C239 VDD2.n95 B 0.009443f
C240 VDD2.n96 B 0.017573f
C241 VDD2.n97 B 0.017573f
C242 VDD2.n98 B 0.009443f
C243 VDD2.n99 B 0.009998f
C244 VDD2.n100 B 0.022319f
C245 VDD2.n101 B 0.022319f
C246 VDD2.n102 B 0.009998f
C247 VDD2.n103 B 0.009443f
C248 VDD2.n104 B 0.017573f
C249 VDD2.n105 B 0.017573f
C250 VDD2.n106 B 0.009443f
C251 VDD2.n107 B 0.009998f
C252 VDD2.n108 B 0.022319f
C253 VDD2.n109 B 0.022319f
C254 VDD2.n110 B 0.009998f
C255 VDD2.n111 B 0.009443f
C256 VDD2.n112 B 0.017573f
C257 VDD2.n113 B 0.017573f
C258 VDD2.n114 B 0.009443f
C259 VDD2.n115 B 0.009998f
C260 VDD2.n116 B 0.022319f
C261 VDD2.n117 B 0.04685f
C262 VDD2.n118 B 0.009998f
C263 VDD2.n119 B 0.009443f
C264 VDD2.n120 B 0.039898f
C265 VDD2.n121 B 0.038181f
C266 VDD2.n122 B 1.79702f
C267 VTAIL.n0 B 0.025552f
C268 VTAIL.n1 B 0.018811f
C269 VTAIL.n2 B 0.010108f
C270 VTAIL.n3 B 0.023892f
C271 VTAIL.n4 B 0.010703f
C272 VTAIL.n5 B 0.018811f
C273 VTAIL.n6 B 0.010108f
C274 VTAIL.n7 B 0.023892f
C275 VTAIL.n8 B 0.010405f
C276 VTAIL.n9 B 0.018811f
C277 VTAIL.n10 B 0.010703f
C278 VTAIL.n11 B 0.023892f
C279 VTAIL.n12 B 0.010703f
C280 VTAIL.n13 B 0.018811f
C281 VTAIL.n14 B 0.010108f
C282 VTAIL.n15 B 0.023892f
C283 VTAIL.n16 B 0.010703f
C284 VTAIL.n17 B 0.896259f
C285 VTAIL.n18 B 0.010108f
C286 VTAIL.t1 B 0.040288f
C287 VTAIL.n19 B 0.131074f
C288 VTAIL.n20 B 0.01689f
C289 VTAIL.n21 B 0.017919f
C290 VTAIL.n22 B 0.023892f
C291 VTAIL.n23 B 0.010703f
C292 VTAIL.n24 B 0.010108f
C293 VTAIL.n25 B 0.018811f
C294 VTAIL.n26 B 0.018811f
C295 VTAIL.n27 B 0.010108f
C296 VTAIL.n28 B 0.010703f
C297 VTAIL.n29 B 0.023892f
C298 VTAIL.n30 B 0.023892f
C299 VTAIL.n31 B 0.010703f
C300 VTAIL.n32 B 0.010108f
C301 VTAIL.n33 B 0.018811f
C302 VTAIL.n34 B 0.018811f
C303 VTAIL.n35 B 0.010108f
C304 VTAIL.n36 B 0.010108f
C305 VTAIL.n37 B 0.010703f
C306 VTAIL.n38 B 0.023892f
C307 VTAIL.n39 B 0.023892f
C308 VTAIL.n40 B 0.023892f
C309 VTAIL.n41 B 0.010405f
C310 VTAIL.n42 B 0.010108f
C311 VTAIL.n43 B 0.018811f
C312 VTAIL.n44 B 0.018811f
C313 VTAIL.n45 B 0.010108f
C314 VTAIL.n46 B 0.010703f
C315 VTAIL.n47 B 0.023892f
C316 VTAIL.n48 B 0.023892f
C317 VTAIL.n49 B 0.010703f
C318 VTAIL.n50 B 0.010108f
C319 VTAIL.n51 B 0.018811f
C320 VTAIL.n52 B 0.018811f
C321 VTAIL.n53 B 0.010108f
C322 VTAIL.n54 B 0.010703f
C323 VTAIL.n55 B 0.023892f
C324 VTAIL.n56 B 0.050151f
C325 VTAIL.n57 B 0.010703f
C326 VTAIL.n58 B 0.010108f
C327 VTAIL.n59 B 0.042709f
C328 VTAIL.n60 B 0.027876f
C329 VTAIL.n61 B 0.987659f
C330 VTAIL.n62 B 0.025552f
C331 VTAIL.n63 B 0.018811f
C332 VTAIL.n64 B 0.010108f
C333 VTAIL.n65 B 0.023892f
C334 VTAIL.n66 B 0.010703f
C335 VTAIL.n67 B 0.018811f
C336 VTAIL.n68 B 0.010108f
C337 VTAIL.n69 B 0.023892f
C338 VTAIL.n70 B 0.010405f
C339 VTAIL.n71 B 0.018811f
C340 VTAIL.n72 B 0.010405f
C341 VTAIL.n73 B 0.010108f
C342 VTAIL.n74 B 0.023892f
C343 VTAIL.n75 B 0.023892f
C344 VTAIL.n76 B 0.010703f
C345 VTAIL.n77 B 0.018811f
C346 VTAIL.n78 B 0.010108f
C347 VTAIL.n79 B 0.023892f
C348 VTAIL.n80 B 0.010703f
C349 VTAIL.n81 B 0.896259f
C350 VTAIL.n82 B 0.010108f
C351 VTAIL.t3 B 0.040288f
C352 VTAIL.n83 B 0.131074f
C353 VTAIL.n84 B 0.01689f
C354 VTAIL.n85 B 0.017919f
C355 VTAIL.n86 B 0.023892f
C356 VTAIL.n87 B 0.010703f
C357 VTAIL.n88 B 0.010108f
C358 VTAIL.n89 B 0.018811f
C359 VTAIL.n90 B 0.018811f
C360 VTAIL.n91 B 0.010108f
C361 VTAIL.n92 B 0.010703f
C362 VTAIL.n93 B 0.023892f
C363 VTAIL.n94 B 0.023892f
C364 VTAIL.n95 B 0.010703f
C365 VTAIL.n96 B 0.010108f
C366 VTAIL.n97 B 0.018811f
C367 VTAIL.n98 B 0.018811f
C368 VTAIL.n99 B 0.010108f
C369 VTAIL.n100 B 0.010703f
C370 VTAIL.n101 B 0.023892f
C371 VTAIL.n102 B 0.023892f
C372 VTAIL.n103 B 0.010703f
C373 VTAIL.n104 B 0.010108f
C374 VTAIL.n105 B 0.018811f
C375 VTAIL.n106 B 0.018811f
C376 VTAIL.n107 B 0.010108f
C377 VTAIL.n108 B 0.010703f
C378 VTAIL.n109 B 0.023892f
C379 VTAIL.n110 B 0.023892f
C380 VTAIL.n111 B 0.010703f
C381 VTAIL.n112 B 0.010108f
C382 VTAIL.n113 B 0.018811f
C383 VTAIL.n114 B 0.018811f
C384 VTAIL.n115 B 0.010108f
C385 VTAIL.n116 B 0.010703f
C386 VTAIL.n117 B 0.023892f
C387 VTAIL.n118 B 0.050151f
C388 VTAIL.n119 B 0.010703f
C389 VTAIL.n120 B 0.010108f
C390 VTAIL.n121 B 0.042709f
C391 VTAIL.n122 B 0.027876f
C392 VTAIL.n123 B 0.99406f
C393 VTAIL.n124 B 0.025552f
C394 VTAIL.n125 B 0.018811f
C395 VTAIL.n126 B 0.010108f
C396 VTAIL.n127 B 0.023892f
C397 VTAIL.n128 B 0.010703f
C398 VTAIL.n129 B 0.018811f
C399 VTAIL.n130 B 0.010108f
C400 VTAIL.n131 B 0.023892f
C401 VTAIL.n132 B 0.010405f
C402 VTAIL.n133 B 0.018811f
C403 VTAIL.n134 B 0.010405f
C404 VTAIL.n135 B 0.010108f
C405 VTAIL.n136 B 0.023892f
C406 VTAIL.n137 B 0.023892f
C407 VTAIL.n138 B 0.010703f
C408 VTAIL.n139 B 0.018811f
C409 VTAIL.n140 B 0.010108f
C410 VTAIL.n141 B 0.023892f
C411 VTAIL.n142 B 0.010703f
C412 VTAIL.n143 B 0.896259f
C413 VTAIL.n144 B 0.010108f
C414 VTAIL.t0 B 0.040288f
C415 VTAIL.n145 B 0.131074f
C416 VTAIL.n146 B 0.01689f
C417 VTAIL.n147 B 0.017919f
C418 VTAIL.n148 B 0.023892f
C419 VTAIL.n149 B 0.010703f
C420 VTAIL.n150 B 0.010108f
C421 VTAIL.n151 B 0.018811f
C422 VTAIL.n152 B 0.018811f
C423 VTAIL.n153 B 0.010108f
C424 VTAIL.n154 B 0.010703f
C425 VTAIL.n155 B 0.023892f
C426 VTAIL.n156 B 0.023892f
C427 VTAIL.n157 B 0.010703f
C428 VTAIL.n158 B 0.010108f
C429 VTAIL.n159 B 0.018811f
C430 VTAIL.n160 B 0.018811f
C431 VTAIL.n161 B 0.010108f
C432 VTAIL.n162 B 0.010703f
C433 VTAIL.n163 B 0.023892f
C434 VTAIL.n164 B 0.023892f
C435 VTAIL.n165 B 0.010703f
C436 VTAIL.n166 B 0.010108f
C437 VTAIL.n167 B 0.018811f
C438 VTAIL.n168 B 0.018811f
C439 VTAIL.n169 B 0.010108f
C440 VTAIL.n170 B 0.010703f
C441 VTAIL.n171 B 0.023892f
C442 VTAIL.n172 B 0.023892f
C443 VTAIL.n173 B 0.010703f
C444 VTAIL.n174 B 0.010108f
C445 VTAIL.n175 B 0.018811f
C446 VTAIL.n176 B 0.018811f
C447 VTAIL.n177 B 0.010108f
C448 VTAIL.n178 B 0.010703f
C449 VTAIL.n179 B 0.023892f
C450 VTAIL.n180 B 0.050151f
C451 VTAIL.n181 B 0.010703f
C452 VTAIL.n182 B 0.010108f
C453 VTAIL.n183 B 0.042709f
C454 VTAIL.n184 B 0.027876f
C455 VTAIL.n185 B 0.954349f
C456 VTAIL.n186 B 0.025552f
C457 VTAIL.n187 B 0.018811f
C458 VTAIL.n188 B 0.010108f
C459 VTAIL.n189 B 0.023892f
C460 VTAIL.n190 B 0.010703f
C461 VTAIL.n191 B 0.018811f
C462 VTAIL.n192 B 0.010108f
C463 VTAIL.n193 B 0.023892f
C464 VTAIL.n194 B 0.010405f
C465 VTAIL.n195 B 0.018811f
C466 VTAIL.n196 B 0.010703f
C467 VTAIL.n197 B 0.023892f
C468 VTAIL.n198 B 0.010703f
C469 VTAIL.n199 B 0.018811f
C470 VTAIL.n200 B 0.010108f
C471 VTAIL.n201 B 0.023892f
C472 VTAIL.n202 B 0.010703f
C473 VTAIL.n203 B 0.896259f
C474 VTAIL.n204 B 0.010108f
C475 VTAIL.t2 B 0.040288f
C476 VTAIL.n205 B 0.131074f
C477 VTAIL.n206 B 0.01689f
C478 VTAIL.n207 B 0.017919f
C479 VTAIL.n208 B 0.023892f
C480 VTAIL.n209 B 0.010703f
C481 VTAIL.n210 B 0.010108f
C482 VTAIL.n211 B 0.018811f
C483 VTAIL.n212 B 0.018811f
C484 VTAIL.n213 B 0.010108f
C485 VTAIL.n214 B 0.010703f
C486 VTAIL.n215 B 0.023892f
C487 VTAIL.n216 B 0.023892f
C488 VTAIL.n217 B 0.010703f
C489 VTAIL.n218 B 0.010108f
C490 VTAIL.n219 B 0.018811f
C491 VTAIL.n220 B 0.018811f
C492 VTAIL.n221 B 0.010108f
C493 VTAIL.n222 B 0.010108f
C494 VTAIL.n223 B 0.010703f
C495 VTAIL.n224 B 0.023892f
C496 VTAIL.n225 B 0.023892f
C497 VTAIL.n226 B 0.023892f
C498 VTAIL.n227 B 0.010405f
C499 VTAIL.n228 B 0.010108f
C500 VTAIL.n229 B 0.018811f
C501 VTAIL.n230 B 0.018811f
C502 VTAIL.n231 B 0.010108f
C503 VTAIL.n232 B 0.010703f
C504 VTAIL.n233 B 0.023892f
C505 VTAIL.n234 B 0.023892f
C506 VTAIL.n235 B 0.010703f
C507 VTAIL.n236 B 0.010108f
C508 VTAIL.n237 B 0.018811f
C509 VTAIL.n238 B 0.018811f
C510 VTAIL.n239 B 0.010108f
C511 VTAIL.n240 B 0.010703f
C512 VTAIL.n241 B 0.023892f
C513 VTAIL.n242 B 0.050151f
C514 VTAIL.n243 B 0.010703f
C515 VTAIL.n244 B 0.010108f
C516 VTAIL.n245 B 0.042709f
C517 VTAIL.n246 B 0.027876f
C518 VTAIL.n247 B 0.912416f
C519 VN.t1 B 0.573833f
C520 VN.t0 B 0.638839f
.ends

