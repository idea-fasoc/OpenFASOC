* NGSPICE file created from diff_pair_sample_1124.ext - technology: sky130A

.subckt diff_pair_sample_1124 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0 ps=0 w=3.09 l=3.84
X1 B.t8 B.t6 B.t7 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0 ps=0 w=3.09 l=3.84
X2 B.t5 B.t3 B.t4 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0 ps=0 w=3.09 l=3.84
X3 VTAIL.t7 VP.t0 VDD1.t0 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0.50985 ps=3.42 w=3.09 l=3.84
X4 VDD2.t3 VN.t0 VTAIL.t2 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=0.50985 pd=3.42 as=1.2051 ps=6.96 w=3.09 l=3.84
X5 B.t2 B.t0 B.t1 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0 ps=0 w=3.09 l=3.84
X6 VDD1.t1 VP.t1 VTAIL.t6 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=0.50985 pd=3.42 as=1.2051 ps=6.96 w=3.09 l=3.84
X7 VTAIL.t3 VN.t1 VDD2.t2 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0.50985 ps=3.42 w=3.09 l=3.84
X8 VDD1.t2 VP.t2 VTAIL.t5 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=0.50985 pd=3.42 as=1.2051 ps=6.96 w=3.09 l=3.84
X9 VDD2.t1 VN.t2 VTAIL.t0 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=0.50985 pd=3.42 as=1.2051 ps=6.96 w=3.09 l=3.84
X10 VTAIL.t1 VN.t3 VDD2.t0 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0.50985 ps=3.42 w=3.09 l=3.84
X11 VTAIL.t4 VP.t3 VDD1.t3 w_n3472_n1586# sky130_fd_pr__pfet_01v8 ad=1.2051 pd=6.96 as=0.50985 ps=3.42 w=3.09 l=3.84
R0 B.n406 B.n405 585
R1 B.n407 B.n48 585
R2 B.n409 B.n408 585
R3 B.n410 B.n47 585
R4 B.n412 B.n411 585
R5 B.n413 B.n46 585
R6 B.n415 B.n414 585
R7 B.n416 B.n45 585
R8 B.n418 B.n417 585
R9 B.n419 B.n44 585
R10 B.n421 B.n420 585
R11 B.n422 B.n43 585
R12 B.n424 B.n423 585
R13 B.n425 B.n42 585
R14 B.n427 B.n426 585
R15 B.n429 B.n39 585
R16 B.n431 B.n430 585
R17 B.n432 B.n38 585
R18 B.n434 B.n433 585
R19 B.n435 B.n37 585
R20 B.n437 B.n436 585
R21 B.n438 B.n36 585
R22 B.n440 B.n439 585
R23 B.n441 B.n35 585
R24 B.n443 B.n442 585
R25 B.n445 B.n444 585
R26 B.n446 B.n31 585
R27 B.n448 B.n447 585
R28 B.n449 B.n30 585
R29 B.n451 B.n450 585
R30 B.n452 B.n29 585
R31 B.n454 B.n453 585
R32 B.n455 B.n28 585
R33 B.n457 B.n456 585
R34 B.n458 B.n27 585
R35 B.n460 B.n459 585
R36 B.n461 B.n26 585
R37 B.n463 B.n462 585
R38 B.n464 B.n25 585
R39 B.n466 B.n465 585
R40 B.n404 B.n49 585
R41 B.n403 B.n402 585
R42 B.n401 B.n50 585
R43 B.n400 B.n399 585
R44 B.n398 B.n51 585
R45 B.n397 B.n396 585
R46 B.n395 B.n52 585
R47 B.n394 B.n393 585
R48 B.n392 B.n53 585
R49 B.n391 B.n390 585
R50 B.n389 B.n54 585
R51 B.n388 B.n387 585
R52 B.n386 B.n55 585
R53 B.n385 B.n384 585
R54 B.n383 B.n56 585
R55 B.n382 B.n381 585
R56 B.n380 B.n57 585
R57 B.n379 B.n378 585
R58 B.n377 B.n58 585
R59 B.n376 B.n375 585
R60 B.n374 B.n59 585
R61 B.n373 B.n372 585
R62 B.n371 B.n60 585
R63 B.n370 B.n369 585
R64 B.n368 B.n61 585
R65 B.n367 B.n366 585
R66 B.n365 B.n62 585
R67 B.n364 B.n363 585
R68 B.n362 B.n63 585
R69 B.n361 B.n360 585
R70 B.n359 B.n64 585
R71 B.n358 B.n357 585
R72 B.n356 B.n65 585
R73 B.n355 B.n354 585
R74 B.n353 B.n66 585
R75 B.n352 B.n351 585
R76 B.n350 B.n67 585
R77 B.n349 B.n348 585
R78 B.n347 B.n68 585
R79 B.n346 B.n345 585
R80 B.n344 B.n69 585
R81 B.n343 B.n342 585
R82 B.n341 B.n70 585
R83 B.n340 B.n339 585
R84 B.n338 B.n71 585
R85 B.n337 B.n336 585
R86 B.n335 B.n72 585
R87 B.n334 B.n333 585
R88 B.n332 B.n73 585
R89 B.n331 B.n330 585
R90 B.n329 B.n74 585
R91 B.n328 B.n327 585
R92 B.n326 B.n75 585
R93 B.n325 B.n324 585
R94 B.n323 B.n76 585
R95 B.n322 B.n321 585
R96 B.n320 B.n77 585
R97 B.n319 B.n318 585
R98 B.n317 B.n78 585
R99 B.n316 B.n315 585
R100 B.n314 B.n79 585
R101 B.n313 B.n312 585
R102 B.n311 B.n80 585
R103 B.n310 B.n309 585
R104 B.n308 B.n81 585
R105 B.n307 B.n306 585
R106 B.n305 B.n82 585
R107 B.n304 B.n303 585
R108 B.n302 B.n83 585
R109 B.n301 B.n300 585
R110 B.n299 B.n84 585
R111 B.n298 B.n297 585
R112 B.n296 B.n85 585
R113 B.n295 B.n294 585
R114 B.n293 B.n86 585
R115 B.n292 B.n291 585
R116 B.n290 B.n87 585
R117 B.n289 B.n288 585
R118 B.n287 B.n88 585
R119 B.n286 B.n285 585
R120 B.n284 B.n89 585
R121 B.n283 B.n282 585
R122 B.n281 B.n90 585
R123 B.n280 B.n279 585
R124 B.n278 B.n91 585
R125 B.n277 B.n276 585
R126 B.n275 B.n92 585
R127 B.n274 B.n273 585
R128 B.n272 B.n93 585
R129 B.n271 B.n270 585
R130 B.n269 B.n94 585
R131 B.n208 B.n207 585
R132 B.n209 B.n118 585
R133 B.n211 B.n210 585
R134 B.n212 B.n117 585
R135 B.n214 B.n213 585
R136 B.n215 B.n116 585
R137 B.n217 B.n216 585
R138 B.n218 B.n115 585
R139 B.n220 B.n219 585
R140 B.n221 B.n114 585
R141 B.n223 B.n222 585
R142 B.n224 B.n113 585
R143 B.n226 B.n225 585
R144 B.n227 B.n112 585
R145 B.n229 B.n228 585
R146 B.n231 B.n109 585
R147 B.n233 B.n232 585
R148 B.n234 B.n108 585
R149 B.n236 B.n235 585
R150 B.n237 B.n107 585
R151 B.n239 B.n238 585
R152 B.n240 B.n106 585
R153 B.n242 B.n241 585
R154 B.n243 B.n105 585
R155 B.n245 B.n244 585
R156 B.n247 B.n246 585
R157 B.n248 B.n101 585
R158 B.n250 B.n249 585
R159 B.n251 B.n100 585
R160 B.n253 B.n252 585
R161 B.n254 B.n99 585
R162 B.n256 B.n255 585
R163 B.n257 B.n98 585
R164 B.n259 B.n258 585
R165 B.n260 B.n97 585
R166 B.n262 B.n261 585
R167 B.n263 B.n96 585
R168 B.n265 B.n264 585
R169 B.n266 B.n95 585
R170 B.n268 B.n267 585
R171 B.n206 B.n119 585
R172 B.n205 B.n204 585
R173 B.n203 B.n120 585
R174 B.n202 B.n201 585
R175 B.n200 B.n121 585
R176 B.n199 B.n198 585
R177 B.n197 B.n122 585
R178 B.n196 B.n195 585
R179 B.n194 B.n123 585
R180 B.n193 B.n192 585
R181 B.n191 B.n124 585
R182 B.n190 B.n189 585
R183 B.n188 B.n125 585
R184 B.n187 B.n186 585
R185 B.n185 B.n126 585
R186 B.n184 B.n183 585
R187 B.n182 B.n127 585
R188 B.n181 B.n180 585
R189 B.n179 B.n128 585
R190 B.n178 B.n177 585
R191 B.n176 B.n129 585
R192 B.n175 B.n174 585
R193 B.n173 B.n130 585
R194 B.n172 B.n171 585
R195 B.n170 B.n131 585
R196 B.n169 B.n168 585
R197 B.n167 B.n132 585
R198 B.n166 B.n165 585
R199 B.n164 B.n133 585
R200 B.n163 B.n162 585
R201 B.n161 B.n134 585
R202 B.n160 B.n159 585
R203 B.n158 B.n135 585
R204 B.n157 B.n156 585
R205 B.n155 B.n136 585
R206 B.n154 B.n153 585
R207 B.n152 B.n137 585
R208 B.n151 B.n150 585
R209 B.n149 B.n138 585
R210 B.n148 B.n147 585
R211 B.n146 B.n139 585
R212 B.n145 B.n144 585
R213 B.n143 B.n140 585
R214 B.n142 B.n141 585
R215 B.n2 B.n0 585
R216 B.n533 B.n1 585
R217 B.n532 B.n531 585
R218 B.n530 B.n3 585
R219 B.n529 B.n528 585
R220 B.n527 B.n4 585
R221 B.n526 B.n525 585
R222 B.n524 B.n5 585
R223 B.n523 B.n522 585
R224 B.n521 B.n6 585
R225 B.n520 B.n519 585
R226 B.n518 B.n7 585
R227 B.n517 B.n516 585
R228 B.n515 B.n8 585
R229 B.n514 B.n513 585
R230 B.n512 B.n9 585
R231 B.n511 B.n510 585
R232 B.n509 B.n10 585
R233 B.n508 B.n507 585
R234 B.n506 B.n11 585
R235 B.n505 B.n504 585
R236 B.n503 B.n12 585
R237 B.n502 B.n501 585
R238 B.n500 B.n13 585
R239 B.n499 B.n498 585
R240 B.n497 B.n14 585
R241 B.n496 B.n495 585
R242 B.n494 B.n15 585
R243 B.n493 B.n492 585
R244 B.n491 B.n16 585
R245 B.n490 B.n489 585
R246 B.n488 B.n17 585
R247 B.n487 B.n486 585
R248 B.n485 B.n18 585
R249 B.n484 B.n483 585
R250 B.n482 B.n19 585
R251 B.n481 B.n480 585
R252 B.n479 B.n20 585
R253 B.n478 B.n477 585
R254 B.n476 B.n21 585
R255 B.n475 B.n474 585
R256 B.n473 B.n22 585
R257 B.n472 B.n471 585
R258 B.n470 B.n23 585
R259 B.n469 B.n468 585
R260 B.n467 B.n24 585
R261 B.n535 B.n534 585
R262 B.n208 B.n119 516.524
R263 B.n467 B.n466 516.524
R264 B.n269 B.n268 516.524
R265 B.n406 B.n49 516.524
R266 B.n102 B.t5 304.3
R267 B.n40 B.t10 304.3
R268 B.n110 B.t8 304.3
R269 B.n32 B.t1 304.3
R270 B.n102 B.t3 228.768
R271 B.n110 B.t6 228.768
R272 B.n32 B.t0 228.768
R273 B.n40 B.t9 228.768
R274 B.n103 B.t4 223.428
R275 B.n41 B.t11 223.428
R276 B.n111 B.t7 223.428
R277 B.n33 B.t2 223.428
R278 B.n204 B.n119 163.367
R279 B.n204 B.n203 163.367
R280 B.n203 B.n202 163.367
R281 B.n202 B.n121 163.367
R282 B.n198 B.n121 163.367
R283 B.n198 B.n197 163.367
R284 B.n197 B.n196 163.367
R285 B.n196 B.n123 163.367
R286 B.n192 B.n123 163.367
R287 B.n192 B.n191 163.367
R288 B.n191 B.n190 163.367
R289 B.n190 B.n125 163.367
R290 B.n186 B.n125 163.367
R291 B.n186 B.n185 163.367
R292 B.n185 B.n184 163.367
R293 B.n184 B.n127 163.367
R294 B.n180 B.n127 163.367
R295 B.n180 B.n179 163.367
R296 B.n179 B.n178 163.367
R297 B.n178 B.n129 163.367
R298 B.n174 B.n129 163.367
R299 B.n174 B.n173 163.367
R300 B.n173 B.n172 163.367
R301 B.n172 B.n131 163.367
R302 B.n168 B.n131 163.367
R303 B.n168 B.n167 163.367
R304 B.n167 B.n166 163.367
R305 B.n166 B.n133 163.367
R306 B.n162 B.n133 163.367
R307 B.n162 B.n161 163.367
R308 B.n161 B.n160 163.367
R309 B.n160 B.n135 163.367
R310 B.n156 B.n135 163.367
R311 B.n156 B.n155 163.367
R312 B.n155 B.n154 163.367
R313 B.n154 B.n137 163.367
R314 B.n150 B.n137 163.367
R315 B.n150 B.n149 163.367
R316 B.n149 B.n148 163.367
R317 B.n148 B.n139 163.367
R318 B.n144 B.n139 163.367
R319 B.n144 B.n143 163.367
R320 B.n143 B.n142 163.367
R321 B.n142 B.n2 163.367
R322 B.n534 B.n2 163.367
R323 B.n534 B.n533 163.367
R324 B.n533 B.n532 163.367
R325 B.n532 B.n3 163.367
R326 B.n528 B.n3 163.367
R327 B.n528 B.n527 163.367
R328 B.n527 B.n526 163.367
R329 B.n526 B.n5 163.367
R330 B.n522 B.n5 163.367
R331 B.n522 B.n521 163.367
R332 B.n521 B.n520 163.367
R333 B.n520 B.n7 163.367
R334 B.n516 B.n7 163.367
R335 B.n516 B.n515 163.367
R336 B.n515 B.n514 163.367
R337 B.n514 B.n9 163.367
R338 B.n510 B.n9 163.367
R339 B.n510 B.n509 163.367
R340 B.n509 B.n508 163.367
R341 B.n508 B.n11 163.367
R342 B.n504 B.n11 163.367
R343 B.n504 B.n503 163.367
R344 B.n503 B.n502 163.367
R345 B.n502 B.n13 163.367
R346 B.n498 B.n13 163.367
R347 B.n498 B.n497 163.367
R348 B.n497 B.n496 163.367
R349 B.n496 B.n15 163.367
R350 B.n492 B.n15 163.367
R351 B.n492 B.n491 163.367
R352 B.n491 B.n490 163.367
R353 B.n490 B.n17 163.367
R354 B.n486 B.n17 163.367
R355 B.n486 B.n485 163.367
R356 B.n485 B.n484 163.367
R357 B.n484 B.n19 163.367
R358 B.n480 B.n19 163.367
R359 B.n480 B.n479 163.367
R360 B.n479 B.n478 163.367
R361 B.n478 B.n21 163.367
R362 B.n474 B.n21 163.367
R363 B.n474 B.n473 163.367
R364 B.n473 B.n472 163.367
R365 B.n472 B.n23 163.367
R366 B.n468 B.n23 163.367
R367 B.n468 B.n467 163.367
R368 B.n209 B.n208 163.367
R369 B.n210 B.n209 163.367
R370 B.n210 B.n117 163.367
R371 B.n214 B.n117 163.367
R372 B.n215 B.n214 163.367
R373 B.n216 B.n215 163.367
R374 B.n216 B.n115 163.367
R375 B.n220 B.n115 163.367
R376 B.n221 B.n220 163.367
R377 B.n222 B.n221 163.367
R378 B.n222 B.n113 163.367
R379 B.n226 B.n113 163.367
R380 B.n227 B.n226 163.367
R381 B.n228 B.n227 163.367
R382 B.n228 B.n109 163.367
R383 B.n233 B.n109 163.367
R384 B.n234 B.n233 163.367
R385 B.n235 B.n234 163.367
R386 B.n235 B.n107 163.367
R387 B.n239 B.n107 163.367
R388 B.n240 B.n239 163.367
R389 B.n241 B.n240 163.367
R390 B.n241 B.n105 163.367
R391 B.n245 B.n105 163.367
R392 B.n246 B.n245 163.367
R393 B.n246 B.n101 163.367
R394 B.n250 B.n101 163.367
R395 B.n251 B.n250 163.367
R396 B.n252 B.n251 163.367
R397 B.n252 B.n99 163.367
R398 B.n256 B.n99 163.367
R399 B.n257 B.n256 163.367
R400 B.n258 B.n257 163.367
R401 B.n258 B.n97 163.367
R402 B.n262 B.n97 163.367
R403 B.n263 B.n262 163.367
R404 B.n264 B.n263 163.367
R405 B.n264 B.n95 163.367
R406 B.n268 B.n95 163.367
R407 B.n270 B.n269 163.367
R408 B.n270 B.n93 163.367
R409 B.n274 B.n93 163.367
R410 B.n275 B.n274 163.367
R411 B.n276 B.n275 163.367
R412 B.n276 B.n91 163.367
R413 B.n280 B.n91 163.367
R414 B.n281 B.n280 163.367
R415 B.n282 B.n281 163.367
R416 B.n282 B.n89 163.367
R417 B.n286 B.n89 163.367
R418 B.n287 B.n286 163.367
R419 B.n288 B.n287 163.367
R420 B.n288 B.n87 163.367
R421 B.n292 B.n87 163.367
R422 B.n293 B.n292 163.367
R423 B.n294 B.n293 163.367
R424 B.n294 B.n85 163.367
R425 B.n298 B.n85 163.367
R426 B.n299 B.n298 163.367
R427 B.n300 B.n299 163.367
R428 B.n300 B.n83 163.367
R429 B.n304 B.n83 163.367
R430 B.n305 B.n304 163.367
R431 B.n306 B.n305 163.367
R432 B.n306 B.n81 163.367
R433 B.n310 B.n81 163.367
R434 B.n311 B.n310 163.367
R435 B.n312 B.n311 163.367
R436 B.n312 B.n79 163.367
R437 B.n316 B.n79 163.367
R438 B.n317 B.n316 163.367
R439 B.n318 B.n317 163.367
R440 B.n318 B.n77 163.367
R441 B.n322 B.n77 163.367
R442 B.n323 B.n322 163.367
R443 B.n324 B.n323 163.367
R444 B.n324 B.n75 163.367
R445 B.n328 B.n75 163.367
R446 B.n329 B.n328 163.367
R447 B.n330 B.n329 163.367
R448 B.n330 B.n73 163.367
R449 B.n334 B.n73 163.367
R450 B.n335 B.n334 163.367
R451 B.n336 B.n335 163.367
R452 B.n336 B.n71 163.367
R453 B.n340 B.n71 163.367
R454 B.n341 B.n340 163.367
R455 B.n342 B.n341 163.367
R456 B.n342 B.n69 163.367
R457 B.n346 B.n69 163.367
R458 B.n347 B.n346 163.367
R459 B.n348 B.n347 163.367
R460 B.n348 B.n67 163.367
R461 B.n352 B.n67 163.367
R462 B.n353 B.n352 163.367
R463 B.n354 B.n353 163.367
R464 B.n354 B.n65 163.367
R465 B.n358 B.n65 163.367
R466 B.n359 B.n358 163.367
R467 B.n360 B.n359 163.367
R468 B.n360 B.n63 163.367
R469 B.n364 B.n63 163.367
R470 B.n365 B.n364 163.367
R471 B.n366 B.n365 163.367
R472 B.n366 B.n61 163.367
R473 B.n370 B.n61 163.367
R474 B.n371 B.n370 163.367
R475 B.n372 B.n371 163.367
R476 B.n372 B.n59 163.367
R477 B.n376 B.n59 163.367
R478 B.n377 B.n376 163.367
R479 B.n378 B.n377 163.367
R480 B.n378 B.n57 163.367
R481 B.n382 B.n57 163.367
R482 B.n383 B.n382 163.367
R483 B.n384 B.n383 163.367
R484 B.n384 B.n55 163.367
R485 B.n388 B.n55 163.367
R486 B.n389 B.n388 163.367
R487 B.n390 B.n389 163.367
R488 B.n390 B.n53 163.367
R489 B.n394 B.n53 163.367
R490 B.n395 B.n394 163.367
R491 B.n396 B.n395 163.367
R492 B.n396 B.n51 163.367
R493 B.n400 B.n51 163.367
R494 B.n401 B.n400 163.367
R495 B.n402 B.n401 163.367
R496 B.n402 B.n49 163.367
R497 B.n466 B.n25 163.367
R498 B.n462 B.n25 163.367
R499 B.n462 B.n461 163.367
R500 B.n461 B.n460 163.367
R501 B.n460 B.n27 163.367
R502 B.n456 B.n27 163.367
R503 B.n456 B.n455 163.367
R504 B.n455 B.n454 163.367
R505 B.n454 B.n29 163.367
R506 B.n450 B.n29 163.367
R507 B.n450 B.n449 163.367
R508 B.n449 B.n448 163.367
R509 B.n448 B.n31 163.367
R510 B.n444 B.n31 163.367
R511 B.n444 B.n443 163.367
R512 B.n443 B.n35 163.367
R513 B.n439 B.n35 163.367
R514 B.n439 B.n438 163.367
R515 B.n438 B.n437 163.367
R516 B.n437 B.n37 163.367
R517 B.n433 B.n37 163.367
R518 B.n433 B.n432 163.367
R519 B.n432 B.n431 163.367
R520 B.n431 B.n39 163.367
R521 B.n426 B.n39 163.367
R522 B.n426 B.n425 163.367
R523 B.n425 B.n424 163.367
R524 B.n424 B.n43 163.367
R525 B.n420 B.n43 163.367
R526 B.n420 B.n419 163.367
R527 B.n419 B.n418 163.367
R528 B.n418 B.n45 163.367
R529 B.n414 B.n45 163.367
R530 B.n414 B.n413 163.367
R531 B.n413 B.n412 163.367
R532 B.n412 B.n47 163.367
R533 B.n408 B.n47 163.367
R534 B.n408 B.n407 163.367
R535 B.n407 B.n406 163.367
R536 B.n103 B.n102 80.8732
R537 B.n111 B.n110 80.8732
R538 B.n33 B.n32 80.8732
R539 B.n41 B.n40 80.8732
R540 B.n104 B.n103 59.5399
R541 B.n230 B.n111 59.5399
R542 B.n34 B.n33 59.5399
R543 B.n428 B.n41 59.5399
R544 B.n465 B.n24 33.5615
R545 B.n405 B.n404 33.5615
R546 B.n267 B.n94 33.5615
R547 B.n207 B.n206 33.5615
R548 B B.n535 18.0485
R549 B.n465 B.n464 10.6151
R550 B.n464 B.n463 10.6151
R551 B.n463 B.n26 10.6151
R552 B.n459 B.n26 10.6151
R553 B.n459 B.n458 10.6151
R554 B.n458 B.n457 10.6151
R555 B.n457 B.n28 10.6151
R556 B.n453 B.n28 10.6151
R557 B.n453 B.n452 10.6151
R558 B.n452 B.n451 10.6151
R559 B.n451 B.n30 10.6151
R560 B.n447 B.n30 10.6151
R561 B.n447 B.n446 10.6151
R562 B.n446 B.n445 10.6151
R563 B.n442 B.n441 10.6151
R564 B.n441 B.n440 10.6151
R565 B.n440 B.n36 10.6151
R566 B.n436 B.n36 10.6151
R567 B.n436 B.n435 10.6151
R568 B.n435 B.n434 10.6151
R569 B.n434 B.n38 10.6151
R570 B.n430 B.n38 10.6151
R571 B.n430 B.n429 10.6151
R572 B.n427 B.n42 10.6151
R573 B.n423 B.n42 10.6151
R574 B.n423 B.n422 10.6151
R575 B.n422 B.n421 10.6151
R576 B.n421 B.n44 10.6151
R577 B.n417 B.n44 10.6151
R578 B.n417 B.n416 10.6151
R579 B.n416 B.n415 10.6151
R580 B.n415 B.n46 10.6151
R581 B.n411 B.n46 10.6151
R582 B.n411 B.n410 10.6151
R583 B.n410 B.n409 10.6151
R584 B.n409 B.n48 10.6151
R585 B.n405 B.n48 10.6151
R586 B.n271 B.n94 10.6151
R587 B.n272 B.n271 10.6151
R588 B.n273 B.n272 10.6151
R589 B.n273 B.n92 10.6151
R590 B.n277 B.n92 10.6151
R591 B.n278 B.n277 10.6151
R592 B.n279 B.n278 10.6151
R593 B.n279 B.n90 10.6151
R594 B.n283 B.n90 10.6151
R595 B.n284 B.n283 10.6151
R596 B.n285 B.n284 10.6151
R597 B.n285 B.n88 10.6151
R598 B.n289 B.n88 10.6151
R599 B.n290 B.n289 10.6151
R600 B.n291 B.n290 10.6151
R601 B.n291 B.n86 10.6151
R602 B.n295 B.n86 10.6151
R603 B.n296 B.n295 10.6151
R604 B.n297 B.n296 10.6151
R605 B.n297 B.n84 10.6151
R606 B.n301 B.n84 10.6151
R607 B.n302 B.n301 10.6151
R608 B.n303 B.n302 10.6151
R609 B.n303 B.n82 10.6151
R610 B.n307 B.n82 10.6151
R611 B.n308 B.n307 10.6151
R612 B.n309 B.n308 10.6151
R613 B.n309 B.n80 10.6151
R614 B.n313 B.n80 10.6151
R615 B.n314 B.n313 10.6151
R616 B.n315 B.n314 10.6151
R617 B.n315 B.n78 10.6151
R618 B.n319 B.n78 10.6151
R619 B.n320 B.n319 10.6151
R620 B.n321 B.n320 10.6151
R621 B.n321 B.n76 10.6151
R622 B.n325 B.n76 10.6151
R623 B.n326 B.n325 10.6151
R624 B.n327 B.n326 10.6151
R625 B.n327 B.n74 10.6151
R626 B.n331 B.n74 10.6151
R627 B.n332 B.n331 10.6151
R628 B.n333 B.n332 10.6151
R629 B.n333 B.n72 10.6151
R630 B.n337 B.n72 10.6151
R631 B.n338 B.n337 10.6151
R632 B.n339 B.n338 10.6151
R633 B.n339 B.n70 10.6151
R634 B.n343 B.n70 10.6151
R635 B.n344 B.n343 10.6151
R636 B.n345 B.n344 10.6151
R637 B.n345 B.n68 10.6151
R638 B.n349 B.n68 10.6151
R639 B.n350 B.n349 10.6151
R640 B.n351 B.n350 10.6151
R641 B.n351 B.n66 10.6151
R642 B.n355 B.n66 10.6151
R643 B.n356 B.n355 10.6151
R644 B.n357 B.n356 10.6151
R645 B.n357 B.n64 10.6151
R646 B.n361 B.n64 10.6151
R647 B.n362 B.n361 10.6151
R648 B.n363 B.n362 10.6151
R649 B.n363 B.n62 10.6151
R650 B.n367 B.n62 10.6151
R651 B.n368 B.n367 10.6151
R652 B.n369 B.n368 10.6151
R653 B.n369 B.n60 10.6151
R654 B.n373 B.n60 10.6151
R655 B.n374 B.n373 10.6151
R656 B.n375 B.n374 10.6151
R657 B.n375 B.n58 10.6151
R658 B.n379 B.n58 10.6151
R659 B.n380 B.n379 10.6151
R660 B.n381 B.n380 10.6151
R661 B.n381 B.n56 10.6151
R662 B.n385 B.n56 10.6151
R663 B.n386 B.n385 10.6151
R664 B.n387 B.n386 10.6151
R665 B.n387 B.n54 10.6151
R666 B.n391 B.n54 10.6151
R667 B.n392 B.n391 10.6151
R668 B.n393 B.n392 10.6151
R669 B.n393 B.n52 10.6151
R670 B.n397 B.n52 10.6151
R671 B.n398 B.n397 10.6151
R672 B.n399 B.n398 10.6151
R673 B.n399 B.n50 10.6151
R674 B.n403 B.n50 10.6151
R675 B.n404 B.n403 10.6151
R676 B.n207 B.n118 10.6151
R677 B.n211 B.n118 10.6151
R678 B.n212 B.n211 10.6151
R679 B.n213 B.n212 10.6151
R680 B.n213 B.n116 10.6151
R681 B.n217 B.n116 10.6151
R682 B.n218 B.n217 10.6151
R683 B.n219 B.n218 10.6151
R684 B.n219 B.n114 10.6151
R685 B.n223 B.n114 10.6151
R686 B.n224 B.n223 10.6151
R687 B.n225 B.n224 10.6151
R688 B.n225 B.n112 10.6151
R689 B.n229 B.n112 10.6151
R690 B.n232 B.n231 10.6151
R691 B.n232 B.n108 10.6151
R692 B.n236 B.n108 10.6151
R693 B.n237 B.n236 10.6151
R694 B.n238 B.n237 10.6151
R695 B.n238 B.n106 10.6151
R696 B.n242 B.n106 10.6151
R697 B.n243 B.n242 10.6151
R698 B.n244 B.n243 10.6151
R699 B.n248 B.n247 10.6151
R700 B.n249 B.n248 10.6151
R701 B.n249 B.n100 10.6151
R702 B.n253 B.n100 10.6151
R703 B.n254 B.n253 10.6151
R704 B.n255 B.n254 10.6151
R705 B.n255 B.n98 10.6151
R706 B.n259 B.n98 10.6151
R707 B.n260 B.n259 10.6151
R708 B.n261 B.n260 10.6151
R709 B.n261 B.n96 10.6151
R710 B.n265 B.n96 10.6151
R711 B.n266 B.n265 10.6151
R712 B.n267 B.n266 10.6151
R713 B.n206 B.n205 10.6151
R714 B.n205 B.n120 10.6151
R715 B.n201 B.n120 10.6151
R716 B.n201 B.n200 10.6151
R717 B.n200 B.n199 10.6151
R718 B.n199 B.n122 10.6151
R719 B.n195 B.n122 10.6151
R720 B.n195 B.n194 10.6151
R721 B.n194 B.n193 10.6151
R722 B.n193 B.n124 10.6151
R723 B.n189 B.n124 10.6151
R724 B.n189 B.n188 10.6151
R725 B.n188 B.n187 10.6151
R726 B.n187 B.n126 10.6151
R727 B.n183 B.n126 10.6151
R728 B.n183 B.n182 10.6151
R729 B.n182 B.n181 10.6151
R730 B.n181 B.n128 10.6151
R731 B.n177 B.n128 10.6151
R732 B.n177 B.n176 10.6151
R733 B.n176 B.n175 10.6151
R734 B.n175 B.n130 10.6151
R735 B.n171 B.n130 10.6151
R736 B.n171 B.n170 10.6151
R737 B.n170 B.n169 10.6151
R738 B.n169 B.n132 10.6151
R739 B.n165 B.n132 10.6151
R740 B.n165 B.n164 10.6151
R741 B.n164 B.n163 10.6151
R742 B.n163 B.n134 10.6151
R743 B.n159 B.n134 10.6151
R744 B.n159 B.n158 10.6151
R745 B.n158 B.n157 10.6151
R746 B.n157 B.n136 10.6151
R747 B.n153 B.n136 10.6151
R748 B.n153 B.n152 10.6151
R749 B.n152 B.n151 10.6151
R750 B.n151 B.n138 10.6151
R751 B.n147 B.n138 10.6151
R752 B.n147 B.n146 10.6151
R753 B.n146 B.n145 10.6151
R754 B.n145 B.n140 10.6151
R755 B.n141 B.n140 10.6151
R756 B.n141 B.n0 10.6151
R757 B.n531 B.n1 10.6151
R758 B.n531 B.n530 10.6151
R759 B.n530 B.n529 10.6151
R760 B.n529 B.n4 10.6151
R761 B.n525 B.n4 10.6151
R762 B.n525 B.n524 10.6151
R763 B.n524 B.n523 10.6151
R764 B.n523 B.n6 10.6151
R765 B.n519 B.n6 10.6151
R766 B.n519 B.n518 10.6151
R767 B.n518 B.n517 10.6151
R768 B.n517 B.n8 10.6151
R769 B.n513 B.n8 10.6151
R770 B.n513 B.n512 10.6151
R771 B.n512 B.n511 10.6151
R772 B.n511 B.n10 10.6151
R773 B.n507 B.n10 10.6151
R774 B.n507 B.n506 10.6151
R775 B.n506 B.n505 10.6151
R776 B.n505 B.n12 10.6151
R777 B.n501 B.n12 10.6151
R778 B.n501 B.n500 10.6151
R779 B.n500 B.n499 10.6151
R780 B.n499 B.n14 10.6151
R781 B.n495 B.n14 10.6151
R782 B.n495 B.n494 10.6151
R783 B.n494 B.n493 10.6151
R784 B.n493 B.n16 10.6151
R785 B.n489 B.n16 10.6151
R786 B.n489 B.n488 10.6151
R787 B.n488 B.n487 10.6151
R788 B.n487 B.n18 10.6151
R789 B.n483 B.n18 10.6151
R790 B.n483 B.n482 10.6151
R791 B.n482 B.n481 10.6151
R792 B.n481 B.n20 10.6151
R793 B.n477 B.n20 10.6151
R794 B.n477 B.n476 10.6151
R795 B.n476 B.n475 10.6151
R796 B.n475 B.n22 10.6151
R797 B.n471 B.n22 10.6151
R798 B.n471 B.n470 10.6151
R799 B.n470 B.n469 10.6151
R800 B.n469 B.n24 10.6151
R801 B.n445 B.n34 9.36635
R802 B.n428 B.n427 9.36635
R803 B.n230 B.n229 9.36635
R804 B.n247 B.n104 9.36635
R805 B.n535 B.n0 2.81026
R806 B.n535 B.n1 2.81026
R807 B.n442 B.n34 1.24928
R808 B.n429 B.n428 1.24928
R809 B.n231 B.n230 1.24928
R810 B.n244 B.n104 1.24928
R811 VP.n21 VP.n20 161.3
R812 VP.n19 VP.n1 161.3
R813 VP.n18 VP.n17 161.3
R814 VP.n16 VP.n2 161.3
R815 VP.n15 VP.n14 161.3
R816 VP.n13 VP.n3 161.3
R817 VP.n12 VP.n11 161.3
R818 VP.n10 VP.n4 161.3
R819 VP.n9 VP.n8 161.3
R820 VP.n7 VP.n6 85.908
R821 VP.n22 VP.n0 85.908
R822 VP.n5 VP.t0 53.5776
R823 VP.n5 VP.t2 52.2179
R824 VP.n6 VP.n5 45.2713
R825 VP.n14 VP.n13 40.4934
R826 VP.n14 VP.n2 40.4934
R827 VP.n8 VP.n4 24.4675
R828 VP.n12 VP.n4 24.4675
R829 VP.n13 VP.n12 24.4675
R830 VP.n18 VP.n2 24.4675
R831 VP.n19 VP.n18 24.4675
R832 VP.n20 VP.n19 24.4675
R833 VP.n7 VP.t3 19.3935
R834 VP.n0 VP.t1 19.3935
R835 VP.n8 VP.n7 4.15989
R836 VP.n20 VP.n0 4.15989
R837 VP.n9 VP.n6 0.354971
R838 VP.n22 VP.n21 0.354971
R839 VP VP.n22 0.26696
R840 VP.n10 VP.n9 0.189894
R841 VP.n11 VP.n10 0.189894
R842 VP.n11 VP.n3 0.189894
R843 VP.n15 VP.n3 0.189894
R844 VP.n16 VP.n15 0.189894
R845 VP.n17 VP.n16 0.189894
R846 VP.n17 VP.n1 0.189894
R847 VP.n21 VP.n1 0.189894
R848 VDD1 VDD1.n1 164.957
R849 VDD1 VDD1.n0 127.328
R850 VDD1.n0 VDD1.t0 10.5199
R851 VDD1.n0 VDD1.t2 10.5199
R852 VDD1.n1 VDD1.t3 10.5199
R853 VDD1.n1 VDD1.t1 10.5199
R854 VTAIL.n122 VTAIL.n112 756.745
R855 VTAIL.n10 VTAIL.n0 756.745
R856 VTAIL.n26 VTAIL.n16 756.745
R857 VTAIL.n42 VTAIL.n32 756.745
R858 VTAIL.n106 VTAIL.n96 756.745
R859 VTAIL.n90 VTAIL.n80 756.745
R860 VTAIL.n74 VTAIL.n64 756.745
R861 VTAIL.n58 VTAIL.n48 756.745
R862 VTAIL.n116 VTAIL.n115 585
R863 VTAIL.n121 VTAIL.n120 585
R864 VTAIL.n123 VTAIL.n122 585
R865 VTAIL.n4 VTAIL.n3 585
R866 VTAIL.n9 VTAIL.n8 585
R867 VTAIL.n11 VTAIL.n10 585
R868 VTAIL.n20 VTAIL.n19 585
R869 VTAIL.n25 VTAIL.n24 585
R870 VTAIL.n27 VTAIL.n26 585
R871 VTAIL.n36 VTAIL.n35 585
R872 VTAIL.n41 VTAIL.n40 585
R873 VTAIL.n43 VTAIL.n42 585
R874 VTAIL.n107 VTAIL.n106 585
R875 VTAIL.n105 VTAIL.n104 585
R876 VTAIL.n100 VTAIL.n99 585
R877 VTAIL.n91 VTAIL.n90 585
R878 VTAIL.n89 VTAIL.n88 585
R879 VTAIL.n84 VTAIL.n83 585
R880 VTAIL.n75 VTAIL.n74 585
R881 VTAIL.n73 VTAIL.n72 585
R882 VTAIL.n68 VTAIL.n67 585
R883 VTAIL.n59 VTAIL.n58 585
R884 VTAIL.n57 VTAIL.n56 585
R885 VTAIL.n52 VTAIL.n51 585
R886 VTAIL.n117 VTAIL.t0 336.901
R887 VTAIL.n5 VTAIL.t3 336.901
R888 VTAIL.n21 VTAIL.t6 336.901
R889 VTAIL.n37 VTAIL.t4 336.901
R890 VTAIL.n101 VTAIL.t5 336.901
R891 VTAIL.n85 VTAIL.t7 336.901
R892 VTAIL.n69 VTAIL.t2 336.901
R893 VTAIL.n53 VTAIL.t1 336.901
R894 VTAIL.n121 VTAIL.n115 171.744
R895 VTAIL.n122 VTAIL.n121 171.744
R896 VTAIL.n9 VTAIL.n3 171.744
R897 VTAIL.n10 VTAIL.n9 171.744
R898 VTAIL.n25 VTAIL.n19 171.744
R899 VTAIL.n26 VTAIL.n25 171.744
R900 VTAIL.n41 VTAIL.n35 171.744
R901 VTAIL.n42 VTAIL.n41 171.744
R902 VTAIL.n106 VTAIL.n105 171.744
R903 VTAIL.n105 VTAIL.n99 171.744
R904 VTAIL.n90 VTAIL.n89 171.744
R905 VTAIL.n89 VTAIL.n83 171.744
R906 VTAIL.n74 VTAIL.n73 171.744
R907 VTAIL.n73 VTAIL.n67 171.744
R908 VTAIL.n58 VTAIL.n57 171.744
R909 VTAIL.n57 VTAIL.n51 171.744
R910 VTAIL.t0 VTAIL.n115 85.8723
R911 VTAIL.t3 VTAIL.n3 85.8723
R912 VTAIL.t6 VTAIL.n19 85.8723
R913 VTAIL.t4 VTAIL.n35 85.8723
R914 VTAIL.t5 VTAIL.n99 85.8723
R915 VTAIL.t7 VTAIL.n83 85.8723
R916 VTAIL.t2 VTAIL.n67 85.8723
R917 VTAIL.t1 VTAIL.n51 85.8723
R918 VTAIL.n127 VTAIL.n126 31.6035
R919 VTAIL.n15 VTAIL.n14 31.6035
R920 VTAIL.n31 VTAIL.n30 31.6035
R921 VTAIL.n47 VTAIL.n46 31.6035
R922 VTAIL.n111 VTAIL.n110 31.6035
R923 VTAIL.n95 VTAIL.n94 31.6035
R924 VTAIL.n79 VTAIL.n78 31.6035
R925 VTAIL.n63 VTAIL.n62 31.6035
R926 VTAIL.n127 VTAIL.n111 18.6255
R927 VTAIL.n63 VTAIL.n47 18.6255
R928 VTAIL.n117 VTAIL.n116 16.193
R929 VTAIL.n5 VTAIL.n4 16.193
R930 VTAIL.n21 VTAIL.n20 16.193
R931 VTAIL.n37 VTAIL.n36 16.193
R932 VTAIL.n101 VTAIL.n100 16.193
R933 VTAIL.n85 VTAIL.n84 16.193
R934 VTAIL.n69 VTAIL.n68 16.193
R935 VTAIL.n53 VTAIL.n52 16.193
R936 VTAIL.n120 VTAIL.n119 12.8005
R937 VTAIL.n8 VTAIL.n7 12.8005
R938 VTAIL.n24 VTAIL.n23 12.8005
R939 VTAIL.n40 VTAIL.n39 12.8005
R940 VTAIL.n104 VTAIL.n103 12.8005
R941 VTAIL.n88 VTAIL.n87 12.8005
R942 VTAIL.n72 VTAIL.n71 12.8005
R943 VTAIL.n56 VTAIL.n55 12.8005
R944 VTAIL.n123 VTAIL.n114 12.0247
R945 VTAIL.n11 VTAIL.n2 12.0247
R946 VTAIL.n27 VTAIL.n18 12.0247
R947 VTAIL.n43 VTAIL.n34 12.0247
R948 VTAIL.n107 VTAIL.n98 12.0247
R949 VTAIL.n91 VTAIL.n82 12.0247
R950 VTAIL.n75 VTAIL.n66 12.0247
R951 VTAIL.n59 VTAIL.n50 12.0247
R952 VTAIL.n124 VTAIL.n112 11.249
R953 VTAIL.n12 VTAIL.n0 11.249
R954 VTAIL.n28 VTAIL.n16 11.249
R955 VTAIL.n44 VTAIL.n32 11.249
R956 VTAIL.n108 VTAIL.n96 11.249
R957 VTAIL.n92 VTAIL.n80 11.249
R958 VTAIL.n76 VTAIL.n64 11.249
R959 VTAIL.n60 VTAIL.n48 11.249
R960 VTAIL.n126 VTAIL.n125 9.45567
R961 VTAIL.n14 VTAIL.n13 9.45567
R962 VTAIL.n30 VTAIL.n29 9.45567
R963 VTAIL.n46 VTAIL.n45 9.45567
R964 VTAIL.n110 VTAIL.n109 9.45567
R965 VTAIL.n94 VTAIL.n93 9.45567
R966 VTAIL.n78 VTAIL.n77 9.45567
R967 VTAIL.n62 VTAIL.n61 9.45567
R968 VTAIL.n125 VTAIL.n124 9.3005
R969 VTAIL.n114 VTAIL.n113 9.3005
R970 VTAIL.n119 VTAIL.n118 9.3005
R971 VTAIL.n13 VTAIL.n12 9.3005
R972 VTAIL.n2 VTAIL.n1 9.3005
R973 VTAIL.n7 VTAIL.n6 9.3005
R974 VTAIL.n29 VTAIL.n28 9.3005
R975 VTAIL.n18 VTAIL.n17 9.3005
R976 VTAIL.n23 VTAIL.n22 9.3005
R977 VTAIL.n45 VTAIL.n44 9.3005
R978 VTAIL.n34 VTAIL.n33 9.3005
R979 VTAIL.n39 VTAIL.n38 9.3005
R980 VTAIL.n109 VTAIL.n108 9.3005
R981 VTAIL.n98 VTAIL.n97 9.3005
R982 VTAIL.n103 VTAIL.n102 9.3005
R983 VTAIL.n93 VTAIL.n92 9.3005
R984 VTAIL.n82 VTAIL.n81 9.3005
R985 VTAIL.n87 VTAIL.n86 9.3005
R986 VTAIL.n77 VTAIL.n76 9.3005
R987 VTAIL.n66 VTAIL.n65 9.3005
R988 VTAIL.n71 VTAIL.n70 9.3005
R989 VTAIL.n61 VTAIL.n60 9.3005
R990 VTAIL.n50 VTAIL.n49 9.3005
R991 VTAIL.n55 VTAIL.n54 9.3005
R992 VTAIL.n102 VTAIL.n101 3.91276
R993 VTAIL.n86 VTAIL.n85 3.91276
R994 VTAIL.n70 VTAIL.n69 3.91276
R995 VTAIL.n54 VTAIL.n53 3.91276
R996 VTAIL.n118 VTAIL.n117 3.91276
R997 VTAIL.n6 VTAIL.n5 3.91276
R998 VTAIL.n22 VTAIL.n21 3.91276
R999 VTAIL.n38 VTAIL.n37 3.91276
R1000 VTAIL.n79 VTAIL.n63 3.59533
R1001 VTAIL.n111 VTAIL.n95 3.59533
R1002 VTAIL.n47 VTAIL.n31 3.59533
R1003 VTAIL.n126 VTAIL.n112 2.71565
R1004 VTAIL.n14 VTAIL.n0 2.71565
R1005 VTAIL.n30 VTAIL.n16 2.71565
R1006 VTAIL.n46 VTAIL.n32 2.71565
R1007 VTAIL.n110 VTAIL.n96 2.71565
R1008 VTAIL.n94 VTAIL.n80 2.71565
R1009 VTAIL.n78 VTAIL.n64 2.71565
R1010 VTAIL.n62 VTAIL.n48 2.71565
R1011 VTAIL.n124 VTAIL.n123 1.93989
R1012 VTAIL.n12 VTAIL.n11 1.93989
R1013 VTAIL.n28 VTAIL.n27 1.93989
R1014 VTAIL.n44 VTAIL.n43 1.93989
R1015 VTAIL.n108 VTAIL.n107 1.93989
R1016 VTAIL.n92 VTAIL.n91 1.93989
R1017 VTAIL.n76 VTAIL.n75 1.93989
R1018 VTAIL.n60 VTAIL.n59 1.93989
R1019 VTAIL VTAIL.n15 1.8561
R1020 VTAIL VTAIL.n127 1.73972
R1021 VTAIL.n120 VTAIL.n114 1.16414
R1022 VTAIL.n8 VTAIL.n2 1.16414
R1023 VTAIL.n24 VTAIL.n18 1.16414
R1024 VTAIL.n40 VTAIL.n34 1.16414
R1025 VTAIL.n104 VTAIL.n98 1.16414
R1026 VTAIL.n88 VTAIL.n82 1.16414
R1027 VTAIL.n72 VTAIL.n66 1.16414
R1028 VTAIL.n56 VTAIL.n50 1.16414
R1029 VTAIL.n95 VTAIL.n79 0.470328
R1030 VTAIL.n31 VTAIL.n15 0.470328
R1031 VTAIL.n119 VTAIL.n116 0.388379
R1032 VTAIL.n7 VTAIL.n4 0.388379
R1033 VTAIL.n23 VTAIL.n20 0.388379
R1034 VTAIL.n39 VTAIL.n36 0.388379
R1035 VTAIL.n103 VTAIL.n100 0.388379
R1036 VTAIL.n87 VTAIL.n84 0.388379
R1037 VTAIL.n71 VTAIL.n68 0.388379
R1038 VTAIL.n55 VTAIL.n52 0.388379
R1039 VTAIL.n118 VTAIL.n113 0.155672
R1040 VTAIL.n125 VTAIL.n113 0.155672
R1041 VTAIL.n6 VTAIL.n1 0.155672
R1042 VTAIL.n13 VTAIL.n1 0.155672
R1043 VTAIL.n22 VTAIL.n17 0.155672
R1044 VTAIL.n29 VTAIL.n17 0.155672
R1045 VTAIL.n38 VTAIL.n33 0.155672
R1046 VTAIL.n45 VTAIL.n33 0.155672
R1047 VTAIL.n109 VTAIL.n97 0.155672
R1048 VTAIL.n102 VTAIL.n97 0.155672
R1049 VTAIL.n93 VTAIL.n81 0.155672
R1050 VTAIL.n86 VTAIL.n81 0.155672
R1051 VTAIL.n77 VTAIL.n65 0.155672
R1052 VTAIL.n70 VTAIL.n65 0.155672
R1053 VTAIL.n61 VTAIL.n49 0.155672
R1054 VTAIL.n54 VTAIL.n49 0.155672
R1055 VN.n0 VN.t1 53.5778
R1056 VN.n1 VN.t0 53.5778
R1057 VN.n0 VN.t2 52.2179
R1058 VN.n1 VN.t3 52.2179
R1059 VN VN.n1 45.4367
R1060 VN VN.n0 1.82681
R1061 VDD2.n2 VDD2.n0 164.433
R1062 VDD2.n2 VDD2.n1 127.269
R1063 VDD2.n1 VDD2.t0 10.5199
R1064 VDD2.n1 VDD2.t3 10.5199
R1065 VDD2.n0 VDD2.t2 10.5199
R1066 VDD2.n0 VDD2.t1 10.5199
R1067 VDD2 VDD2.n2 0.0586897
C0 VTAIL B 2.26843f
C1 VDD2 VN 1.5528f
C2 VTAIL VDD2 3.97712f
C3 VDD1 VN 0.154812f
C4 w_n3472_n1586# VN 5.94156f
C5 B VP 1.98215f
C6 VTAIL VDD1 3.9146f
C7 VTAIL w_n3472_n1586# 2.05554f
C8 VDD2 VP 0.478581f
C9 B VDD2 1.31415f
C10 VDD1 VP 1.87472f
C11 VTAIL VN 2.29268f
C12 B VDD1 1.24119f
C13 w_n3472_n1586# VP 6.38885f
C14 B w_n3472_n1586# 8.31519f
C15 VDD2 VDD1 1.3281f
C16 VN VP 5.44011f
C17 VDD2 w_n3472_n1586# 1.52306f
C18 B VN 1.2309f
C19 VTAIL VP 2.30678f
C20 w_n3472_n1586# VDD1 1.44011f
C21 VDD2 VSUBS 0.855439f
C22 VDD1 VSUBS 4.02731f
C23 VTAIL VSUBS 0.734534f
C24 VN VSUBS 6.11601f
C25 VP VSUBS 2.395899f
C26 B VSUBS 4.331995f
C27 w_n3472_n1586# VSUBS 69.7039f
C28 VDD2.t2 VSUBS 0.052494f
C29 VDD2.t1 VSUBS 0.052494f
C30 VDD2.n0 VSUBS 0.513133f
C31 VDD2.t0 VSUBS 0.052494f
C32 VDD2.t3 VSUBS 0.052494f
C33 VDD2.n1 VSUBS 0.280242f
C34 VDD2.n2 VSUBS 2.743f
C35 VN.t2 VSUBS 1.69107f
C36 VN.t1 VSUBS 1.71238f
C37 VN.n0 VSUBS 1.07149f
C38 VN.t3 VSUBS 1.69107f
C39 VN.t0 VSUBS 1.71238f
C40 VN.n1 VSUBS 3.28722f
C41 VTAIL.n0 VSUBS 0.035529f
C42 VTAIL.n1 VSUBS 0.035036f
C43 VTAIL.n2 VSUBS 0.018827f
C44 VTAIL.n3 VSUBS 0.033375f
C45 VTAIL.n4 VSUBS 0.027473f
C46 VTAIL.t3 VSUBS 0.097494f
C47 VTAIL.n5 VSUBS 0.12447f
C48 VTAIL.n6 VSUBS 0.339788f
C49 VTAIL.n7 VSUBS 0.018827f
C50 VTAIL.n8 VSUBS 0.019934f
C51 VTAIL.n9 VSUBS 0.0445f
C52 VTAIL.n10 VSUBS 0.097619f
C53 VTAIL.n11 VSUBS 0.019934f
C54 VTAIL.n12 VSUBS 0.018827f
C55 VTAIL.n13 VSUBS 0.079549f
C56 VTAIL.n14 VSUBS 0.048598f
C57 VTAIL.n15 VSUBS 0.291643f
C58 VTAIL.n16 VSUBS 0.035529f
C59 VTAIL.n17 VSUBS 0.035036f
C60 VTAIL.n18 VSUBS 0.018827f
C61 VTAIL.n19 VSUBS 0.033375f
C62 VTAIL.n20 VSUBS 0.027473f
C63 VTAIL.t6 VSUBS 0.097494f
C64 VTAIL.n21 VSUBS 0.12447f
C65 VTAIL.n22 VSUBS 0.339788f
C66 VTAIL.n23 VSUBS 0.018827f
C67 VTAIL.n24 VSUBS 0.019934f
C68 VTAIL.n25 VSUBS 0.0445f
C69 VTAIL.n26 VSUBS 0.097619f
C70 VTAIL.n27 VSUBS 0.019934f
C71 VTAIL.n28 VSUBS 0.018827f
C72 VTAIL.n29 VSUBS 0.079549f
C73 VTAIL.n30 VSUBS 0.048598f
C74 VTAIL.n31 VSUBS 0.487992f
C75 VTAIL.n32 VSUBS 0.035529f
C76 VTAIL.n33 VSUBS 0.035036f
C77 VTAIL.n34 VSUBS 0.018827f
C78 VTAIL.n35 VSUBS 0.033375f
C79 VTAIL.n36 VSUBS 0.027473f
C80 VTAIL.t4 VSUBS 0.097494f
C81 VTAIL.n37 VSUBS 0.12447f
C82 VTAIL.n38 VSUBS 0.339788f
C83 VTAIL.n39 VSUBS 0.018827f
C84 VTAIL.n40 VSUBS 0.019934f
C85 VTAIL.n41 VSUBS 0.0445f
C86 VTAIL.n42 VSUBS 0.097619f
C87 VTAIL.n43 VSUBS 0.019934f
C88 VTAIL.n44 VSUBS 0.018827f
C89 VTAIL.n45 VSUBS 0.079549f
C90 VTAIL.n46 VSUBS 0.048598f
C91 VTAIL.n47 VSUBS 1.61744f
C92 VTAIL.n48 VSUBS 0.035529f
C93 VTAIL.n49 VSUBS 0.035036f
C94 VTAIL.n50 VSUBS 0.018827f
C95 VTAIL.n51 VSUBS 0.033375f
C96 VTAIL.n52 VSUBS 0.027473f
C97 VTAIL.t1 VSUBS 0.097494f
C98 VTAIL.n53 VSUBS 0.12447f
C99 VTAIL.n54 VSUBS 0.339788f
C100 VTAIL.n55 VSUBS 0.018827f
C101 VTAIL.n56 VSUBS 0.019934f
C102 VTAIL.n57 VSUBS 0.0445f
C103 VTAIL.n58 VSUBS 0.097619f
C104 VTAIL.n59 VSUBS 0.019934f
C105 VTAIL.n60 VSUBS 0.018827f
C106 VTAIL.n61 VSUBS 0.079549f
C107 VTAIL.n62 VSUBS 0.048598f
C108 VTAIL.n63 VSUBS 1.61744f
C109 VTAIL.n64 VSUBS 0.035529f
C110 VTAIL.n65 VSUBS 0.035036f
C111 VTAIL.n66 VSUBS 0.018827f
C112 VTAIL.n67 VSUBS 0.033375f
C113 VTAIL.n68 VSUBS 0.027473f
C114 VTAIL.t2 VSUBS 0.097494f
C115 VTAIL.n69 VSUBS 0.12447f
C116 VTAIL.n70 VSUBS 0.339788f
C117 VTAIL.n71 VSUBS 0.018827f
C118 VTAIL.n72 VSUBS 0.019934f
C119 VTAIL.n73 VSUBS 0.0445f
C120 VTAIL.n74 VSUBS 0.097619f
C121 VTAIL.n75 VSUBS 0.019934f
C122 VTAIL.n76 VSUBS 0.018827f
C123 VTAIL.n77 VSUBS 0.079549f
C124 VTAIL.n78 VSUBS 0.048598f
C125 VTAIL.n79 VSUBS 0.487992f
C126 VTAIL.n80 VSUBS 0.035529f
C127 VTAIL.n81 VSUBS 0.035036f
C128 VTAIL.n82 VSUBS 0.018827f
C129 VTAIL.n83 VSUBS 0.033375f
C130 VTAIL.n84 VSUBS 0.027473f
C131 VTAIL.t7 VSUBS 0.097494f
C132 VTAIL.n85 VSUBS 0.12447f
C133 VTAIL.n86 VSUBS 0.339788f
C134 VTAIL.n87 VSUBS 0.018827f
C135 VTAIL.n88 VSUBS 0.019934f
C136 VTAIL.n89 VSUBS 0.0445f
C137 VTAIL.n90 VSUBS 0.097619f
C138 VTAIL.n91 VSUBS 0.019934f
C139 VTAIL.n92 VSUBS 0.018827f
C140 VTAIL.n93 VSUBS 0.079549f
C141 VTAIL.n94 VSUBS 0.048598f
C142 VTAIL.n95 VSUBS 0.487992f
C143 VTAIL.n96 VSUBS 0.035529f
C144 VTAIL.n97 VSUBS 0.035036f
C145 VTAIL.n98 VSUBS 0.018827f
C146 VTAIL.n99 VSUBS 0.033375f
C147 VTAIL.n100 VSUBS 0.027473f
C148 VTAIL.t5 VSUBS 0.097494f
C149 VTAIL.n101 VSUBS 0.12447f
C150 VTAIL.n102 VSUBS 0.339788f
C151 VTAIL.n103 VSUBS 0.018827f
C152 VTAIL.n104 VSUBS 0.019934f
C153 VTAIL.n105 VSUBS 0.0445f
C154 VTAIL.n106 VSUBS 0.097619f
C155 VTAIL.n107 VSUBS 0.019934f
C156 VTAIL.n108 VSUBS 0.018827f
C157 VTAIL.n109 VSUBS 0.079549f
C158 VTAIL.n110 VSUBS 0.048598f
C159 VTAIL.n111 VSUBS 1.61744f
C160 VTAIL.n112 VSUBS 0.035529f
C161 VTAIL.n113 VSUBS 0.035036f
C162 VTAIL.n114 VSUBS 0.018827f
C163 VTAIL.n115 VSUBS 0.033375f
C164 VTAIL.n116 VSUBS 0.027473f
C165 VTAIL.t0 VSUBS 0.097494f
C166 VTAIL.n117 VSUBS 0.12447f
C167 VTAIL.n118 VSUBS 0.339788f
C168 VTAIL.n119 VSUBS 0.018827f
C169 VTAIL.n120 VSUBS 0.019934f
C170 VTAIL.n121 VSUBS 0.0445f
C171 VTAIL.n122 VSUBS 0.097619f
C172 VTAIL.n123 VSUBS 0.019934f
C173 VTAIL.n124 VSUBS 0.018827f
C174 VTAIL.n125 VSUBS 0.079549f
C175 VTAIL.n126 VSUBS 0.048598f
C176 VTAIL.n127 VSUBS 1.40796f
C177 VDD1.t0 VSUBS 0.050185f
C178 VDD1.t2 VSUBS 0.050185f
C179 VDD1.n0 VSUBS 0.268152f
C180 VDD1.t3 VSUBS 0.050185f
C181 VDD1.t1 VSUBS 0.050185f
C182 VDD1.n1 VSUBS 0.50238f
C183 VP.t1 VSUBS 1.24026f
C184 VP.n0 VSUBS 0.663255f
C185 VP.n1 VSUBS 0.041808f
C186 VP.n2 VSUBS 0.083092f
C187 VP.n3 VSUBS 0.041808f
C188 VP.n4 VSUBS 0.077919f
C189 VP.t0 VSUBS 1.78273f
C190 VP.t2 VSUBS 1.76054f
C191 VP.n5 VSUBS 3.40465f
C192 VP.n6 VSUBS 2.09584f
C193 VP.t3 VSUBS 1.24026f
C194 VP.n7 VSUBS 0.663255f
C195 VP.n8 VSUBS 0.045988f
C196 VP.n9 VSUBS 0.067477f
C197 VP.n10 VSUBS 0.041808f
C198 VP.n11 VSUBS 0.041808f
C199 VP.n12 VSUBS 0.077919f
C200 VP.n13 VSUBS 0.083092f
C201 VP.n14 VSUBS 0.033798f
C202 VP.n15 VSUBS 0.041808f
C203 VP.n16 VSUBS 0.041808f
C204 VP.n17 VSUBS 0.041808f
C205 VP.n18 VSUBS 0.077919f
C206 VP.n19 VSUBS 0.077919f
C207 VP.n20 VSUBS 0.045988f
C208 VP.n21 VSUBS 0.067477f
C209 VP.n22 VSUBS 0.127725f
C210 B.n0 VSUBS 0.006209f
C211 B.n1 VSUBS 0.006209f
C212 B.n2 VSUBS 0.009819f
C213 B.n3 VSUBS 0.009819f
C214 B.n4 VSUBS 0.009819f
C215 B.n5 VSUBS 0.009819f
C216 B.n6 VSUBS 0.009819f
C217 B.n7 VSUBS 0.009819f
C218 B.n8 VSUBS 0.009819f
C219 B.n9 VSUBS 0.009819f
C220 B.n10 VSUBS 0.009819f
C221 B.n11 VSUBS 0.009819f
C222 B.n12 VSUBS 0.009819f
C223 B.n13 VSUBS 0.009819f
C224 B.n14 VSUBS 0.009819f
C225 B.n15 VSUBS 0.009819f
C226 B.n16 VSUBS 0.009819f
C227 B.n17 VSUBS 0.009819f
C228 B.n18 VSUBS 0.009819f
C229 B.n19 VSUBS 0.009819f
C230 B.n20 VSUBS 0.009819f
C231 B.n21 VSUBS 0.009819f
C232 B.n22 VSUBS 0.009819f
C233 B.n23 VSUBS 0.009819f
C234 B.n24 VSUBS 0.023131f
C235 B.n25 VSUBS 0.009819f
C236 B.n26 VSUBS 0.009819f
C237 B.n27 VSUBS 0.009819f
C238 B.n28 VSUBS 0.009819f
C239 B.n29 VSUBS 0.009819f
C240 B.n30 VSUBS 0.009819f
C241 B.n31 VSUBS 0.009819f
C242 B.t2 VSUBS 0.063543f
C243 B.t1 VSUBS 0.097309f
C244 B.t0 VSUBS 0.816244f
C245 B.n32 VSUBS 0.168985f
C246 B.n33 VSUBS 0.141056f
C247 B.n34 VSUBS 0.02275f
C248 B.n35 VSUBS 0.009819f
C249 B.n36 VSUBS 0.009819f
C250 B.n37 VSUBS 0.009819f
C251 B.n38 VSUBS 0.009819f
C252 B.n39 VSUBS 0.009819f
C253 B.t11 VSUBS 0.063544f
C254 B.t10 VSUBS 0.097309f
C255 B.t9 VSUBS 0.816244f
C256 B.n40 VSUBS 0.168984f
C257 B.n41 VSUBS 0.141055f
C258 B.n42 VSUBS 0.009819f
C259 B.n43 VSUBS 0.009819f
C260 B.n44 VSUBS 0.009819f
C261 B.n45 VSUBS 0.009819f
C262 B.n46 VSUBS 0.009819f
C263 B.n47 VSUBS 0.009819f
C264 B.n48 VSUBS 0.009819f
C265 B.n49 VSUBS 0.023131f
C266 B.n50 VSUBS 0.009819f
C267 B.n51 VSUBS 0.009819f
C268 B.n52 VSUBS 0.009819f
C269 B.n53 VSUBS 0.009819f
C270 B.n54 VSUBS 0.009819f
C271 B.n55 VSUBS 0.009819f
C272 B.n56 VSUBS 0.009819f
C273 B.n57 VSUBS 0.009819f
C274 B.n58 VSUBS 0.009819f
C275 B.n59 VSUBS 0.009819f
C276 B.n60 VSUBS 0.009819f
C277 B.n61 VSUBS 0.009819f
C278 B.n62 VSUBS 0.009819f
C279 B.n63 VSUBS 0.009819f
C280 B.n64 VSUBS 0.009819f
C281 B.n65 VSUBS 0.009819f
C282 B.n66 VSUBS 0.009819f
C283 B.n67 VSUBS 0.009819f
C284 B.n68 VSUBS 0.009819f
C285 B.n69 VSUBS 0.009819f
C286 B.n70 VSUBS 0.009819f
C287 B.n71 VSUBS 0.009819f
C288 B.n72 VSUBS 0.009819f
C289 B.n73 VSUBS 0.009819f
C290 B.n74 VSUBS 0.009819f
C291 B.n75 VSUBS 0.009819f
C292 B.n76 VSUBS 0.009819f
C293 B.n77 VSUBS 0.009819f
C294 B.n78 VSUBS 0.009819f
C295 B.n79 VSUBS 0.009819f
C296 B.n80 VSUBS 0.009819f
C297 B.n81 VSUBS 0.009819f
C298 B.n82 VSUBS 0.009819f
C299 B.n83 VSUBS 0.009819f
C300 B.n84 VSUBS 0.009819f
C301 B.n85 VSUBS 0.009819f
C302 B.n86 VSUBS 0.009819f
C303 B.n87 VSUBS 0.009819f
C304 B.n88 VSUBS 0.009819f
C305 B.n89 VSUBS 0.009819f
C306 B.n90 VSUBS 0.009819f
C307 B.n91 VSUBS 0.009819f
C308 B.n92 VSUBS 0.009819f
C309 B.n93 VSUBS 0.009819f
C310 B.n94 VSUBS 0.023131f
C311 B.n95 VSUBS 0.009819f
C312 B.n96 VSUBS 0.009819f
C313 B.n97 VSUBS 0.009819f
C314 B.n98 VSUBS 0.009819f
C315 B.n99 VSUBS 0.009819f
C316 B.n100 VSUBS 0.009819f
C317 B.n101 VSUBS 0.009819f
C318 B.t4 VSUBS 0.063544f
C319 B.t5 VSUBS 0.097309f
C320 B.t3 VSUBS 0.816244f
C321 B.n102 VSUBS 0.168984f
C322 B.n103 VSUBS 0.141055f
C323 B.n104 VSUBS 0.02275f
C324 B.n105 VSUBS 0.009819f
C325 B.n106 VSUBS 0.009819f
C326 B.n107 VSUBS 0.009819f
C327 B.n108 VSUBS 0.009819f
C328 B.n109 VSUBS 0.009819f
C329 B.t7 VSUBS 0.063543f
C330 B.t8 VSUBS 0.097309f
C331 B.t6 VSUBS 0.816244f
C332 B.n110 VSUBS 0.168985f
C333 B.n111 VSUBS 0.141056f
C334 B.n112 VSUBS 0.009819f
C335 B.n113 VSUBS 0.009819f
C336 B.n114 VSUBS 0.009819f
C337 B.n115 VSUBS 0.009819f
C338 B.n116 VSUBS 0.009819f
C339 B.n117 VSUBS 0.009819f
C340 B.n118 VSUBS 0.009819f
C341 B.n119 VSUBS 0.023131f
C342 B.n120 VSUBS 0.009819f
C343 B.n121 VSUBS 0.009819f
C344 B.n122 VSUBS 0.009819f
C345 B.n123 VSUBS 0.009819f
C346 B.n124 VSUBS 0.009819f
C347 B.n125 VSUBS 0.009819f
C348 B.n126 VSUBS 0.009819f
C349 B.n127 VSUBS 0.009819f
C350 B.n128 VSUBS 0.009819f
C351 B.n129 VSUBS 0.009819f
C352 B.n130 VSUBS 0.009819f
C353 B.n131 VSUBS 0.009819f
C354 B.n132 VSUBS 0.009819f
C355 B.n133 VSUBS 0.009819f
C356 B.n134 VSUBS 0.009819f
C357 B.n135 VSUBS 0.009819f
C358 B.n136 VSUBS 0.009819f
C359 B.n137 VSUBS 0.009819f
C360 B.n138 VSUBS 0.009819f
C361 B.n139 VSUBS 0.009819f
C362 B.n140 VSUBS 0.009819f
C363 B.n141 VSUBS 0.009819f
C364 B.n142 VSUBS 0.009819f
C365 B.n143 VSUBS 0.009819f
C366 B.n144 VSUBS 0.009819f
C367 B.n145 VSUBS 0.009819f
C368 B.n146 VSUBS 0.009819f
C369 B.n147 VSUBS 0.009819f
C370 B.n148 VSUBS 0.009819f
C371 B.n149 VSUBS 0.009819f
C372 B.n150 VSUBS 0.009819f
C373 B.n151 VSUBS 0.009819f
C374 B.n152 VSUBS 0.009819f
C375 B.n153 VSUBS 0.009819f
C376 B.n154 VSUBS 0.009819f
C377 B.n155 VSUBS 0.009819f
C378 B.n156 VSUBS 0.009819f
C379 B.n157 VSUBS 0.009819f
C380 B.n158 VSUBS 0.009819f
C381 B.n159 VSUBS 0.009819f
C382 B.n160 VSUBS 0.009819f
C383 B.n161 VSUBS 0.009819f
C384 B.n162 VSUBS 0.009819f
C385 B.n163 VSUBS 0.009819f
C386 B.n164 VSUBS 0.009819f
C387 B.n165 VSUBS 0.009819f
C388 B.n166 VSUBS 0.009819f
C389 B.n167 VSUBS 0.009819f
C390 B.n168 VSUBS 0.009819f
C391 B.n169 VSUBS 0.009819f
C392 B.n170 VSUBS 0.009819f
C393 B.n171 VSUBS 0.009819f
C394 B.n172 VSUBS 0.009819f
C395 B.n173 VSUBS 0.009819f
C396 B.n174 VSUBS 0.009819f
C397 B.n175 VSUBS 0.009819f
C398 B.n176 VSUBS 0.009819f
C399 B.n177 VSUBS 0.009819f
C400 B.n178 VSUBS 0.009819f
C401 B.n179 VSUBS 0.009819f
C402 B.n180 VSUBS 0.009819f
C403 B.n181 VSUBS 0.009819f
C404 B.n182 VSUBS 0.009819f
C405 B.n183 VSUBS 0.009819f
C406 B.n184 VSUBS 0.009819f
C407 B.n185 VSUBS 0.009819f
C408 B.n186 VSUBS 0.009819f
C409 B.n187 VSUBS 0.009819f
C410 B.n188 VSUBS 0.009819f
C411 B.n189 VSUBS 0.009819f
C412 B.n190 VSUBS 0.009819f
C413 B.n191 VSUBS 0.009819f
C414 B.n192 VSUBS 0.009819f
C415 B.n193 VSUBS 0.009819f
C416 B.n194 VSUBS 0.009819f
C417 B.n195 VSUBS 0.009819f
C418 B.n196 VSUBS 0.009819f
C419 B.n197 VSUBS 0.009819f
C420 B.n198 VSUBS 0.009819f
C421 B.n199 VSUBS 0.009819f
C422 B.n200 VSUBS 0.009819f
C423 B.n201 VSUBS 0.009819f
C424 B.n202 VSUBS 0.009819f
C425 B.n203 VSUBS 0.009819f
C426 B.n204 VSUBS 0.009819f
C427 B.n205 VSUBS 0.009819f
C428 B.n206 VSUBS 0.023131f
C429 B.n207 VSUBS 0.023655f
C430 B.n208 VSUBS 0.023655f
C431 B.n209 VSUBS 0.009819f
C432 B.n210 VSUBS 0.009819f
C433 B.n211 VSUBS 0.009819f
C434 B.n212 VSUBS 0.009819f
C435 B.n213 VSUBS 0.009819f
C436 B.n214 VSUBS 0.009819f
C437 B.n215 VSUBS 0.009819f
C438 B.n216 VSUBS 0.009819f
C439 B.n217 VSUBS 0.009819f
C440 B.n218 VSUBS 0.009819f
C441 B.n219 VSUBS 0.009819f
C442 B.n220 VSUBS 0.009819f
C443 B.n221 VSUBS 0.009819f
C444 B.n222 VSUBS 0.009819f
C445 B.n223 VSUBS 0.009819f
C446 B.n224 VSUBS 0.009819f
C447 B.n225 VSUBS 0.009819f
C448 B.n226 VSUBS 0.009819f
C449 B.n227 VSUBS 0.009819f
C450 B.n228 VSUBS 0.009819f
C451 B.n229 VSUBS 0.009242f
C452 B.n230 VSUBS 0.02275f
C453 B.n231 VSUBS 0.005487f
C454 B.n232 VSUBS 0.009819f
C455 B.n233 VSUBS 0.009819f
C456 B.n234 VSUBS 0.009819f
C457 B.n235 VSUBS 0.009819f
C458 B.n236 VSUBS 0.009819f
C459 B.n237 VSUBS 0.009819f
C460 B.n238 VSUBS 0.009819f
C461 B.n239 VSUBS 0.009819f
C462 B.n240 VSUBS 0.009819f
C463 B.n241 VSUBS 0.009819f
C464 B.n242 VSUBS 0.009819f
C465 B.n243 VSUBS 0.009819f
C466 B.n244 VSUBS 0.005487f
C467 B.n245 VSUBS 0.009819f
C468 B.n246 VSUBS 0.009819f
C469 B.n247 VSUBS 0.009242f
C470 B.n248 VSUBS 0.009819f
C471 B.n249 VSUBS 0.009819f
C472 B.n250 VSUBS 0.009819f
C473 B.n251 VSUBS 0.009819f
C474 B.n252 VSUBS 0.009819f
C475 B.n253 VSUBS 0.009819f
C476 B.n254 VSUBS 0.009819f
C477 B.n255 VSUBS 0.009819f
C478 B.n256 VSUBS 0.009819f
C479 B.n257 VSUBS 0.009819f
C480 B.n258 VSUBS 0.009819f
C481 B.n259 VSUBS 0.009819f
C482 B.n260 VSUBS 0.009819f
C483 B.n261 VSUBS 0.009819f
C484 B.n262 VSUBS 0.009819f
C485 B.n263 VSUBS 0.009819f
C486 B.n264 VSUBS 0.009819f
C487 B.n265 VSUBS 0.009819f
C488 B.n266 VSUBS 0.009819f
C489 B.n267 VSUBS 0.023655f
C490 B.n268 VSUBS 0.023655f
C491 B.n269 VSUBS 0.023131f
C492 B.n270 VSUBS 0.009819f
C493 B.n271 VSUBS 0.009819f
C494 B.n272 VSUBS 0.009819f
C495 B.n273 VSUBS 0.009819f
C496 B.n274 VSUBS 0.009819f
C497 B.n275 VSUBS 0.009819f
C498 B.n276 VSUBS 0.009819f
C499 B.n277 VSUBS 0.009819f
C500 B.n278 VSUBS 0.009819f
C501 B.n279 VSUBS 0.009819f
C502 B.n280 VSUBS 0.009819f
C503 B.n281 VSUBS 0.009819f
C504 B.n282 VSUBS 0.009819f
C505 B.n283 VSUBS 0.009819f
C506 B.n284 VSUBS 0.009819f
C507 B.n285 VSUBS 0.009819f
C508 B.n286 VSUBS 0.009819f
C509 B.n287 VSUBS 0.009819f
C510 B.n288 VSUBS 0.009819f
C511 B.n289 VSUBS 0.009819f
C512 B.n290 VSUBS 0.009819f
C513 B.n291 VSUBS 0.009819f
C514 B.n292 VSUBS 0.009819f
C515 B.n293 VSUBS 0.009819f
C516 B.n294 VSUBS 0.009819f
C517 B.n295 VSUBS 0.009819f
C518 B.n296 VSUBS 0.009819f
C519 B.n297 VSUBS 0.009819f
C520 B.n298 VSUBS 0.009819f
C521 B.n299 VSUBS 0.009819f
C522 B.n300 VSUBS 0.009819f
C523 B.n301 VSUBS 0.009819f
C524 B.n302 VSUBS 0.009819f
C525 B.n303 VSUBS 0.009819f
C526 B.n304 VSUBS 0.009819f
C527 B.n305 VSUBS 0.009819f
C528 B.n306 VSUBS 0.009819f
C529 B.n307 VSUBS 0.009819f
C530 B.n308 VSUBS 0.009819f
C531 B.n309 VSUBS 0.009819f
C532 B.n310 VSUBS 0.009819f
C533 B.n311 VSUBS 0.009819f
C534 B.n312 VSUBS 0.009819f
C535 B.n313 VSUBS 0.009819f
C536 B.n314 VSUBS 0.009819f
C537 B.n315 VSUBS 0.009819f
C538 B.n316 VSUBS 0.009819f
C539 B.n317 VSUBS 0.009819f
C540 B.n318 VSUBS 0.009819f
C541 B.n319 VSUBS 0.009819f
C542 B.n320 VSUBS 0.009819f
C543 B.n321 VSUBS 0.009819f
C544 B.n322 VSUBS 0.009819f
C545 B.n323 VSUBS 0.009819f
C546 B.n324 VSUBS 0.009819f
C547 B.n325 VSUBS 0.009819f
C548 B.n326 VSUBS 0.009819f
C549 B.n327 VSUBS 0.009819f
C550 B.n328 VSUBS 0.009819f
C551 B.n329 VSUBS 0.009819f
C552 B.n330 VSUBS 0.009819f
C553 B.n331 VSUBS 0.009819f
C554 B.n332 VSUBS 0.009819f
C555 B.n333 VSUBS 0.009819f
C556 B.n334 VSUBS 0.009819f
C557 B.n335 VSUBS 0.009819f
C558 B.n336 VSUBS 0.009819f
C559 B.n337 VSUBS 0.009819f
C560 B.n338 VSUBS 0.009819f
C561 B.n339 VSUBS 0.009819f
C562 B.n340 VSUBS 0.009819f
C563 B.n341 VSUBS 0.009819f
C564 B.n342 VSUBS 0.009819f
C565 B.n343 VSUBS 0.009819f
C566 B.n344 VSUBS 0.009819f
C567 B.n345 VSUBS 0.009819f
C568 B.n346 VSUBS 0.009819f
C569 B.n347 VSUBS 0.009819f
C570 B.n348 VSUBS 0.009819f
C571 B.n349 VSUBS 0.009819f
C572 B.n350 VSUBS 0.009819f
C573 B.n351 VSUBS 0.009819f
C574 B.n352 VSUBS 0.009819f
C575 B.n353 VSUBS 0.009819f
C576 B.n354 VSUBS 0.009819f
C577 B.n355 VSUBS 0.009819f
C578 B.n356 VSUBS 0.009819f
C579 B.n357 VSUBS 0.009819f
C580 B.n358 VSUBS 0.009819f
C581 B.n359 VSUBS 0.009819f
C582 B.n360 VSUBS 0.009819f
C583 B.n361 VSUBS 0.009819f
C584 B.n362 VSUBS 0.009819f
C585 B.n363 VSUBS 0.009819f
C586 B.n364 VSUBS 0.009819f
C587 B.n365 VSUBS 0.009819f
C588 B.n366 VSUBS 0.009819f
C589 B.n367 VSUBS 0.009819f
C590 B.n368 VSUBS 0.009819f
C591 B.n369 VSUBS 0.009819f
C592 B.n370 VSUBS 0.009819f
C593 B.n371 VSUBS 0.009819f
C594 B.n372 VSUBS 0.009819f
C595 B.n373 VSUBS 0.009819f
C596 B.n374 VSUBS 0.009819f
C597 B.n375 VSUBS 0.009819f
C598 B.n376 VSUBS 0.009819f
C599 B.n377 VSUBS 0.009819f
C600 B.n378 VSUBS 0.009819f
C601 B.n379 VSUBS 0.009819f
C602 B.n380 VSUBS 0.009819f
C603 B.n381 VSUBS 0.009819f
C604 B.n382 VSUBS 0.009819f
C605 B.n383 VSUBS 0.009819f
C606 B.n384 VSUBS 0.009819f
C607 B.n385 VSUBS 0.009819f
C608 B.n386 VSUBS 0.009819f
C609 B.n387 VSUBS 0.009819f
C610 B.n388 VSUBS 0.009819f
C611 B.n389 VSUBS 0.009819f
C612 B.n390 VSUBS 0.009819f
C613 B.n391 VSUBS 0.009819f
C614 B.n392 VSUBS 0.009819f
C615 B.n393 VSUBS 0.009819f
C616 B.n394 VSUBS 0.009819f
C617 B.n395 VSUBS 0.009819f
C618 B.n396 VSUBS 0.009819f
C619 B.n397 VSUBS 0.009819f
C620 B.n398 VSUBS 0.009819f
C621 B.n399 VSUBS 0.009819f
C622 B.n400 VSUBS 0.009819f
C623 B.n401 VSUBS 0.009819f
C624 B.n402 VSUBS 0.009819f
C625 B.n403 VSUBS 0.009819f
C626 B.n404 VSUBS 0.02426f
C627 B.n405 VSUBS 0.022526f
C628 B.n406 VSUBS 0.023655f
C629 B.n407 VSUBS 0.009819f
C630 B.n408 VSUBS 0.009819f
C631 B.n409 VSUBS 0.009819f
C632 B.n410 VSUBS 0.009819f
C633 B.n411 VSUBS 0.009819f
C634 B.n412 VSUBS 0.009819f
C635 B.n413 VSUBS 0.009819f
C636 B.n414 VSUBS 0.009819f
C637 B.n415 VSUBS 0.009819f
C638 B.n416 VSUBS 0.009819f
C639 B.n417 VSUBS 0.009819f
C640 B.n418 VSUBS 0.009819f
C641 B.n419 VSUBS 0.009819f
C642 B.n420 VSUBS 0.009819f
C643 B.n421 VSUBS 0.009819f
C644 B.n422 VSUBS 0.009819f
C645 B.n423 VSUBS 0.009819f
C646 B.n424 VSUBS 0.009819f
C647 B.n425 VSUBS 0.009819f
C648 B.n426 VSUBS 0.009819f
C649 B.n427 VSUBS 0.009242f
C650 B.n428 VSUBS 0.02275f
C651 B.n429 VSUBS 0.005487f
C652 B.n430 VSUBS 0.009819f
C653 B.n431 VSUBS 0.009819f
C654 B.n432 VSUBS 0.009819f
C655 B.n433 VSUBS 0.009819f
C656 B.n434 VSUBS 0.009819f
C657 B.n435 VSUBS 0.009819f
C658 B.n436 VSUBS 0.009819f
C659 B.n437 VSUBS 0.009819f
C660 B.n438 VSUBS 0.009819f
C661 B.n439 VSUBS 0.009819f
C662 B.n440 VSUBS 0.009819f
C663 B.n441 VSUBS 0.009819f
C664 B.n442 VSUBS 0.005487f
C665 B.n443 VSUBS 0.009819f
C666 B.n444 VSUBS 0.009819f
C667 B.n445 VSUBS 0.009242f
C668 B.n446 VSUBS 0.009819f
C669 B.n447 VSUBS 0.009819f
C670 B.n448 VSUBS 0.009819f
C671 B.n449 VSUBS 0.009819f
C672 B.n450 VSUBS 0.009819f
C673 B.n451 VSUBS 0.009819f
C674 B.n452 VSUBS 0.009819f
C675 B.n453 VSUBS 0.009819f
C676 B.n454 VSUBS 0.009819f
C677 B.n455 VSUBS 0.009819f
C678 B.n456 VSUBS 0.009819f
C679 B.n457 VSUBS 0.009819f
C680 B.n458 VSUBS 0.009819f
C681 B.n459 VSUBS 0.009819f
C682 B.n460 VSUBS 0.009819f
C683 B.n461 VSUBS 0.009819f
C684 B.n462 VSUBS 0.009819f
C685 B.n463 VSUBS 0.009819f
C686 B.n464 VSUBS 0.009819f
C687 B.n465 VSUBS 0.023655f
C688 B.n466 VSUBS 0.023655f
C689 B.n467 VSUBS 0.023131f
C690 B.n468 VSUBS 0.009819f
C691 B.n469 VSUBS 0.009819f
C692 B.n470 VSUBS 0.009819f
C693 B.n471 VSUBS 0.009819f
C694 B.n472 VSUBS 0.009819f
C695 B.n473 VSUBS 0.009819f
C696 B.n474 VSUBS 0.009819f
C697 B.n475 VSUBS 0.009819f
C698 B.n476 VSUBS 0.009819f
C699 B.n477 VSUBS 0.009819f
C700 B.n478 VSUBS 0.009819f
C701 B.n479 VSUBS 0.009819f
C702 B.n480 VSUBS 0.009819f
C703 B.n481 VSUBS 0.009819f
C704 B.n482 VSUBS 0.009819f
C705 B.n483 VSUBS 0.009819f
C706 B.n484 VSUBS 0.009819f
C707 B.n485 VSUBS 0.009819f
C708 B.n486 VSUBS 0.009819f
C709 B.n487 VSUBS 0.009819f
C710 B.n488 VSUBS 0.009819f
C711 B.n489 VSUBS 0.009819f
C712 B.n490 VSUBS 0.009819f
C713 B.n491 VSUBS 0.009819f
C714 B.n492 VSUBS 0.009819f
C715 B.n493 VSUBS 0.009819f
C716 B.n494 VSUBS 0.009819f
C717 B.n495 VSUBS 0.009819f
C718 B.n496 VSUBS 0.009819f
C719 B.n497 VSUBS 0.009819f
C720 B.n498 VSUBS 0.009819f
C721 B.n499 VSUBS 0.009819f
C722 B.n500 VSUBS 0.009819f
C723 B.n501 VSUBS 0.009819f
C724 B.n502 VSUBS 0.009819f
C725 B.n503 VSUBS 0.009819f
C726 B.n504 VSUBS 0.009819f
C727 B.n505 VSUBS 0.009819f
C728 B.n506 VSUBS 0.009819f
C729 B.n507 VSUBS 0.009819f
C730 B.n508 VSUBS 0.009819f
C731 B.n509 VSUBS 0.009819f
C732 B.n510 VSUBS 0.009819f
C733 B.n511 VSUBS 0.009819f
C734 B.n512 VSUBS 0.009819f
C735 B.n513 VSUBS 0.009819f
C736 B.n514 VSUBS 0.009819f
C737 B.n515 VSUBS 0.009819f
C738 B.n516 VSUBS 0.009819f
C739 B.n517 VSUBS 0.009819f
C740 B.n518 VSUBS 0.009819f
C741 B.n519 VSUBS 0.009819f
C742 B.n520 VSUBS 0.009819f
C743 B.n521 VSUBS 0.009819f
C744 B.n522 VSUBS 0.009819f
C745 B.n523 VSUBS 0.009819f
C746 B.n524 VSUBS 0.009819f
C747 B.n525 VSUBS 0.009819f
C748 B.n526 VSUBS 0.009819f
C749 B.n527 VSUBS 0.009819f
C750 B.n528 VSUBS 0.009819f
C751 B.n529 VSUBS 0.009819f
C752 B.n530 VSUBS 0.009819f
C753 B.n531 VSUBS 0.009819f
C754 B.n532 VSUBS 0.009819f
C755 B.n533 VSUBS 0.009819f
C756 B.n534 VSUBS 0.009819f
C757 B.n535 VSUBS 0.022234f
.ends

