* NGSPICE file created from diff_pair_sample_0268.ext - technology: sky130A

.subckt diff_pair_sample_0268 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0 ps=0 w=2.64 l=2
X1 VDD1.t9 VP.t0 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=1.0296 ps=6.06 w=2.64 l=2
X2 VDD1.t8 VP.t1 VTAIL.t10 B.t6 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X3 VDD1.t7 VP.t2 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X4 VTAIL.t9 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X5 VTAIL.t1 VN.t1 VDD2.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X6 VTAIL.t18 VP.t3 VDD1.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X7 VDD1.t5 VP.t4 VTAIL.t19 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0.4356 ps=2.97 w=2.64 l=2
X8 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0 ps=0 w=2.64 l=2
X9 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0 ps=0 w=2.64 l=2
X10 VDD2.t7 VN.t2 VTAIL.t4 B.t6 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X11 VTAIL.t8 VN.t3 VDD2.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X12 VDD2.t5 VN.t4 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0.4356 ps=2.97 w=2.64 l=2
X13 VDD2.t4 VN.t5 VTAIL.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X14 VDD2.t3 VN.t6 VTAIL.t3 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=1.0296 ps=6.06 w=2.64 l=2
X15 VDD1.t4 VP.t5 VTAIL.t12 B.t0 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0.4356 ps=2.97 w=2.64 l=2
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0 ps=0 w=2.64 l=2
X17 VTAIL.t17 VP.t6 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X18 VDD1.t2 VP.t7 VTAIL.t15 B.t9 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=1.0296 ps=6.06 w=2.64 l=2
X19 VTAIL.t16 VP.t8 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X20 VTAIL.t7 VN.t7 VDD2.t2 B.t8 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X21 VTAIL.t11 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=0.4356 ps=2.97 w=2.64 l=2
X22 VDD2.t1 VN.t8 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=0.4356 pd=2.97 as=1.0296 ps=6.06 w=2.64 l=2
X23 VDD2.t0 VN.t9 VTAIL.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=1.0296 pd=6.06 as=0.4356 ps=2.97 w=2.64 l=2
R0 B.n595 B.n594 585
R1 B.n188 B.n109 585
R2 B.n187 B.n186 585
R3 B.n185 B.n184 585
R4 B.n183 B.n182 585
R5 B.n181 B.n180 585
R6 B.n179 B.n178 585
R7 B.n177 B.n176 585
R8 B.n175 B.n174 585
R9 B.n173 B.n172 585
R10 B.n171 B.n170 585
R11 B.n169 B.n168 585
R12 B.n167 B.n166 585
R13 B.n165 B.n164 585
R14 B.n163 B.n162 585
R15 B.n161 B.n160 585
R16 B.n159 B.n158 585
R17 B.n157 B.n156 585
R18 B.n155 B.n154 585
R19 B.n153 B.n152 585
R20 B.n151 B.n150 585
R21 B.n149 B.n148 585
R22 B.n147 B.n146 585
R23 B.n145 B.n144 585
R24 B.n143 B.n142 585
R25 B.n141 B.n140 585
R26 B.n139 B.n138 585
R27 B.n137 B.n136 585
R28 B.n135 B.n134 585
R29 B.n133 B.n132 585
R30 B.n131 B.n130 585
R31 B.n129 B.n128 585
R32 B.n127 B.n126 585
R33 B.n125 B.n124 585
R34 B.n123 B.n122 585
R35 B.n121 B.n120 585
R36 B.n119 B.n118 585
R37 B.n117 B.n116 585
R38 B.n593 B.n90 585
R39 B.n598 B.n90 585
R40 B.n592 B.n89 585
R41 B.n599 B.n89 585
R42 B.n591 B.n590 585
R43 B.n590 B.n85 585
R44 B.n589 B.n84 585
R45 B.n605 B.n84 585
R46 B.n588 B.n83 585
R47 B.n606 B.n83 585
R48 B.n587 B.n82 585
R49 B.n607 B.n82 585
R50 B.n586 B.n585 585
R51 B.n585 B.n81 585
R52 B.n584 B.n77 585
R53 B.n613 B.n77 585
R54 B.n583 B.n76 585
R55 B.n614 B.n76 585
R56 B.n582 B.n75 585
R57 B.n615 B.n75 585
R58 B.n581 B.n580 585
R59 B.n580 B.n71 585
R60 B.n579 B.n70 585
R61 B.n621 B.n70 585
R62 B.n578 B.n69 585
R63 B.n622 B.n69 585
R64 B.n577 B.n68 585
R65 B.n623 B.n68 585
R66 B.n576 B.n575 585
R67 B.n575 B.n64 585
R68 B.n574 B.n63 585
R69 B.n629 B.n63 585
R70 B.n573 B.n62 585
R71 B.n630 B.n62 585
R72 B.n572 B.n61 585
R73 B.n631 B.n61 585
R74 B.n571 B.n570 585
R75 B.n570 B.n57 585
R76 B.n569 B.n56 585
R77 B.n637 B.n56 585
R78 B.n568 B.n55 585
R79 B.n638 B.n55 585
R80 B.n567 B.n54 585
R81 B.n639 B.n54 585
R82 B.n566 B.n565 585
R83 B.n565 B.n50 585
R84 B.n564 B.n49 585
R85 B.n645 B.n49 585
R86 B.n563 B.n48 585
R87 B.n646 B.n48 585
R88 B.n562 B.n47 585
R89 B.n647 B.n47 585
R90 B.n561 B.n560 585
R91 B.n560 B.n43 585
R92 B.n559 B.n42 585
R93 B.n653 B.n42 585
R94 B.n558 B.n41 585
R95 B.n654 B.n41 585
R96 B.n557 B.n40 585
R97 B.n655 B.n40 585
R98 B.n556 B.n555 585
R99 B.n555 B.n39 585
R100 B.n554 B.n35 585
R101 B.n661 B.n35 585
R102 B.n553 B.n34 585
R103 B.n662 B.n34 585
R104 B.n552 B.n33 585
R105 B.n663 B.n33 585
R106 B.n551 B.n550 585
R107 B.n550 B.n29 585
R108 B.n549 B.n28 585
R109 B.n669 B.n28 585
R110 B.n548 B.n27 585
R111 B.n670 B.n27 585
R112 B.n547 B.n26 585
R113 B.n671 B.n26 585
R114 B.n546 B.n545 585
R115 B.n545 B.n22 585
R116 B.n544 B.n21 585
R117 B.n677 B.n21 585
R118 B.n543 B.n20 585
R119 B.n678 B.n20 585
R120 B.n542 B.n19 585
R121 B.n679 B.n19 585
R122 B.n541 B.n540 585
R123 B.n540 B.n15 585
R124 B.n539 B.n14 585
R125 B.n685 B.n14 585
R126 B.n538 B.n13 585
R127 B.n686 B.n13 585
R128 B.n537 B.n12 585
R129 B.n687 B.n12 585
R130 B.n536 B.n535 585
R131 B.n535 B.n8 585
R132 B.n534 B.n7 585
R133 B.n693 B.n7 585
R134 B.n533 B.n6 585
R135 B.n694 B.n6 585
R136 B.n532 B.n5 585
R137 B.n695 B.n5 585
R138 B.n531 B.n530 585
R139 B.n530 B.n4 585
R140 B.n529 B.n189 585
R141 B.n529 B.n528 585
R142 B.n519 B.n190 585
R143 B.n191 B.n190 585
R144 B.n521 B.n520 585
R145 B.n522 B.n521 585
R146 B.n518 B.n196 585
R147 B.n196 B.n195 585
R148 B.n517 B.n516 585
R149 B.n516 B.n515 585
R150 B.n198 B.n197 585
R151 B.n199 B.n198 585
R152 B.n508 B.n507 585
R153 B.n509 B.n508 585
R154 B.n506 B.n204 585
R155 B.n204 B.n203 585
R156 B.n505 B.n504 585
R157 B.n504 B.n503 585
R158 B.n206 B.n205 585
R159 B.n207 B.n206 585
R160 B.n496 B.n495 585
R161 B.n497 B.n496 585
R162 B.n494 B.n212 585
R163 B.n212 B.n211 585
R164 B.n493 B.n492 585
R165 B.n492 B.n491 585
R166 B.n214 B.n213 585
R167 B.n215 B.n214 585
R168 B.n484 B.n483 585
R169 B.n485 B.n484 585
R170 B.n482 B.n220 585
R171 B.n220 B.n219 585
R172 B.n481 B.n480 585
R173 B.n480 B.n479 585
R174 B.n222 B.n221 585
R175 B.n472 B.n222 585
R176 B.n471 B.n470 585
R177 B.n473 B.n471 585
R178 B.n469 B.n227 585
R179 B.n227 B.n226 585
R180 B.n468 B.n467 585
R181 B.n467 B.n466 585
R182 B.n229 B.n228 585
R183 B.n230 B.n229 585
R184 B.n459 B.n458 585
R185 B.n460 B.n459 585
R186 B.n457 B.n235 585
R187 B.n235 B.n234 585
R188 B.n456 B.n455 585
R189 B.n455 B.n454 585
R190 B.n237 B.n236 585
R191 B.n238 B.n237 585
R192 B.n447 B.n446 585
R193 B.n448 B.n447 585
R194 B.n445 B.n243 585
R195 B.n243 B.n242 585
R196 B.n444 B.n443 585
R197 B.n443 B.n442 585
R198 B.n245 B.n244 585
R199 B.n246 B.n245 585
R200 B.n435 B.n434 585
R201 B.n436 B.n435 585
R202 B.n433 B.n250 585
R203 B.n254 B.n250 585
R204 B.n432 B.n431 585
R205 B.n431 B.n430 585
R206 B.n252 B.n251 585
R207 B.n253 B.n252 585
R208 B.n423 B.n422 585
R209 B.n424 B.n423 585
R210 B.n421 B.n259 585
R211 B.n259 B.n258 585
R212 B.n420 B.n419 585
R213 B.n419 B.n418 585
R214 B.n261 B.n260 585
R215 B.n262 B.n261 585
R216 B.n411 B.n410 585
R217 B.n412 B.n411 585
R218 B.n409 B.n267 585
R219 B.n267 B.n266 585
R220 B.n408 B.n407 585
R221 B.n407 B.n406 585
R222 B.n269 B.n268 585
R223 B.n399 B.n269 585
R224 B.n398 B.n397 585
R225 B.n400 B.n398 585
R226 B.n396 B.n274 585
R227 B.n274 B.n273 585
R228 B.n395 B.n394 585
R229 B.n394 B.n393 585
R230 B.n276 B.n275 585
R231 B.n277 B.n276 585
R232 B.n386 B.n385 585
R233 B.n387 B.n386 585
R234 B.n384 B.n282 585
R235 B.n282 B.n281 585
R236 B.n379 B.n378 585
R237 B.n377 B.n303 585
R238 B.n376 B.n302 585
R239 B.n381 B.n302 585
R240 B.n375 B.n374 585
R241 B.n373 B.n372 585
R242 B.n371 B.n370 585
R243 B.n369 B.n368 585
R244 B.n367 B.n366 585
R245 B.n365 B.n364 585
R246 B.n363 B.n362 585
R247 B.n361 B.n360 585
R248 B.n359 B.n358 585
R249 B.n357 B.n356 585
R250 B.n355 B.n354 585
R251 B.n352 B.n351 585
R252 B.n350 B.n349 585
R253 B.n348 B.n347 585
R254 B.n346 B.n345 585
R255 B.n344 B.n343 585
R256 B.n342 B.n341 585
R257 B.n340 B.n339 585
R258 B.n338 B.n337 585
R259 B.n336 B.n335 585
R260 B.n334 B.n333 585
R261 B.n331 B.n330 585
R262 B.n329 B.n328 585
R263 B.n327 B.n326 585
R264 B.n325 B.n324 585
R265 B.n323 B.n322 585
R266 B.n321 B.n320 585
R267 B.n319 B.n318 585
R268 B.n317 B.n316 585
R269 B.n315 B.n314 585
R270 B.n313 B.n312 585
R271 B.n311 B.n310 585
R272 B.n309 B.n308 585
R273 B.n284 B.n283 585
R274 B.n383 B.n382 585
R275 B.n382 B.n381 585
R276 B.n280 B.n279 585
R277 B.n281 B.n280 585
R278 B.n389 B.n388 585
R279 B.n388 B.n387 585
R280 B.n390 B.n278 585
R281 B.n278 B.n277 585
R282 B.n392 B.n391 585
R283 B.n393 B.n392 585
R284 B.n272 B.n271 585
R285 B.n273 B.n272 585
R286 B.n402 B.n401 585
R287 B.n401 B.n400 585
R288 B.n403 B.n270 585
R289 B.n399 B.n270 585
R290 B.n405 B.n404 585
R291 B.n406 B.n405 585
R292 B.n265 B.n264 585
R293 B.n266 B.n265 585
R294 B.n414 B.n413 585
R295 B.n413 B.n412 585
R296 B.n415 B.n263 585
R297 B.n263 B.n262 585
R298 B.n417 B.n416 585
R299 B.n418 B.n417 585
R300 B.n257 B.n256 585
R301 B.n258 B.n257 585
R302 B.n426 B.n425 585
R303 B.n425 B.n424 585
R304 B.n427 B.n255 585
R305 B.n255 B.n253 585
R306 B.n429 B.n428 585
R307 B.n430 B.n429 585
R308 B.n249 B.n248 585
R309 B.n254 B.n249 585
R310 B.n438 B.n437 585
R311 B.n437 B.n436 585
R312 B.n439 B.n247 585
R313 B.n247 B.n246 585
R314 B.n441 B.n440 585
R315 B.n442 B.n441 585
R316 B.n241 B.n240 585
R317 B.n242 B.n241 585
R318 B.n450 B.n449 585
R319 B.n449 B.n448 585
R320 B.n451 B.n239 585
R321 B.n239 B.n238 585
R322 B.n453 B.n452 585
R323 B.n454 B.n453 585
R324 B.n233 B.n232 585
R325 B.n234 B.n233 585
R326 B.n462 B.n461 585
R327 B.n461 B.n460 585
R328 B.n463 B.n231 585
R329 B.n231 B.n230 585
R330 B.n465 B.n464 585
R331 B.n466 B.n465 585
R332 B.n225 B.n224 585
R333 B.n226 B.n225 585
R334 B.n475 B.n474 585
R335 B.n474 B.n473 585
R336 B.n476 B.n223 585
R337 B.n472 B.n223 585
R338 B.n478 B.n477 585
R339 B.n479 B.n478 585
R340 B.n218 B.n217 585
R341 B.n219 B.n218 585
R342 B.n487 B.n486 585
R343 B.n486 B.n485 585
R344 B.n488 B.n216 585
R345 B.n216 B.n215 585
R346 B.n490 B.n489 585
R347 B.n491 B.n490 585
R348 B.n210 B.n209 585
R349 B.n211 B.n210 585
R350 B.n499 B.n498 585
R351 B.n498 B.n497 585
R352 B.n500 B.n208 585
R353 B.n208 B.n207 585
R354 B.n502 B.n501 585
R355 B.n503 B.n502 585
R356 B.n202 B.n201 585
R357 B.n203 B.n202 585
R358 B.n511 B.n510 585
R359 B.n510 B.n509 585
R360 B.n512 B.n200 585
R361 B.n200 B.n199 585
R362 B.n514 B.n513 585
R363 B.n515 B.n514 585
R364 B.n194 B.n193 585
R365 B.n195 B.n194 585
R366 B.n524 B.n523 585
R367 B.n523 B.n522 585
R368 B.n525 B.n192 585
R369 B.n192 B.n191 585
R370 B.n527 B.n526 585
R371 B.n528 B.n527 585
R372 B.n2 B.n0 585
R373 B.n4 B.n2 585
R374 B.n3 B.n1 585
R375 B.n694 B.n3 585
R376 B.n692 B.n691 585
R377 B.n693 B.n692 585
R378 B.n690 B.n9 585
R379 B.n9 B.n8 585
R380 B.n689 B.n688 585
R381 B.n688 B.n687 585
R382 B.n11 B.n10 585
R383 B.n686 B.n11 585
R384 B.n684 B.n683 585
R385 B.n685 B.n684 585
R386 B.n682 B.n16 585
R387 B.n16 B.n15 585
R388 B.n681 B.n680 585
R389 B.n680 B.n679 585
R390 B.n18 B.n17 585
R391 B.n678 B.n18 585
R392 B.n676 B.n675 585
R393 B.n677 B.n676 585
R394 B.n674 B.n23 585
R395 B.n23 B.n22 585
R396 B.n673 B.n672 585
R397 B.n672 B.n671 585
R398 B.n25 B.n24 585
R399 B.n670 B.n25 585
R400 B.n668 B.n667 585
R401 B.n669 B.n668 585
R402 B.n666 B.n30 585
R403 B.n30 B.n29 585
R404 B.n665 B.n664 585
R405 B.n664 B.n663 585
R406 B.n32 B.n31 585
R407 B.n662 B.n32 585
R408 B.n660 B.n659 585
R409 B.n661 B.n660 585
R410 B.n658 B.n36 585
R411 B.n39 B.n36 585
R412 B.n657 B.n656 585
R413 B.n656 B.n655 585
R414 B.n38 B.n37 585
R415 B.n654 B.n38 585
R416 B.n652 B.n651 585
R417 B.n653 B.n652 585
R418 B.n650 B.n44 585
R419 B.n44 B.n43 585
R420 B.n649 B.n648 585
R421 B.n648 B.n647 585
R422 B.n46 B.n45 585
R423 B.n646 B.n46 585
R424 B.n644 B.n643 585
R425 B.n645 B.n644 585
R426 B.n642 B.n51 585
R427 B.n51 B.n50 585
R428 B.n641 B.n640 585
R429 B.n640 B.n639 585
R430 B.n53 B.n52 585
R431 B.n638 B.n53 585
R432 B.n636 B.n635 585
R433 B.n637 B.n636 585
R434 B.n634 B.n58 585
R435 B.n58 B.n57 585
R436 B.n633 B.n632 585
R437 B.n632 B.n631 585
R438 B.n60 B.n59 585
R439 B.n630 B.n60 585
R440 B.n628 B.n627 585
R441 B.n629 B.n628 585
R442 B.n626 B.n65 585
R443 B.n65 B.n64 585
R444 B.n625 B.n624 585
R445 B.n624 B.n623 585
R446 B.n67 B.n66 585
R447 B.n622 B.n67 585
R448 B.n620 B.n619 585
R449 B.n621 B.n620 585
R450 B.n618 B.n72 585
R451 B.n72 B.n71 585
R452 B.n617 B.n616 585
R453 B.n616 B.n615 585
R454 B.n74 B.n73 585
R455 B.n614 B.n74 585
R456 B.n612 B.n611 585
R457 B.n613 B.n612 585
R458 B.n610 B.n78 585
R459 B.n81 B.n78 585
R460 B.n609 B.n608 585
R461 B.n608 B.n607 585
R462 B.n80 B.n79 585
R463 B.n606 B.n80 585
R464 B.n604 B.n603 585
R465 B.n605 B.n604 585
R466 B.n602 B.n86 585
R467 B.n86 B.n85 585
R468 B.n601 B.n600 585
R469 B.n600 B.n599 585
R470 B.n88 B.n87 585
R471 B.n598 B.n88 585
R472 B.n697 B.n696 585
R473 B.n696 B.n695 585
R474 B.n379 B.n280 516.524
R475 B.n116 B.n88 516.524
R476 B.n382 B.n282 516.524
R477 B.n595 B.n90 516.524
R478 B.n597 B.n596 256.663
R479 B.n597 B.n108 256.663
R480 B.n597 B.n107 256.663
R481 B.n597 B.n106 256.663
R482 B.n597 B.n105 256.663
R483 B.n597 B.n104 256.663
R484 B.n597 B.n103 256.663
R485 B.n597 B.n102 256.663
R486 B.n597 B.n101 256.663
R487 B.n597 B.n100 256.663
R488 B.n597 B.n99 256.663
R489 B.n597 B.n98 256.663
R490 B.n597 B.n97 256.663
R491 B.n597 B.n96 256.663
R492 B.n597 B.n95 256.663
R493 B.n597 B.n94 256.663
R494 B.n597 B.n93 256.663
R495 B.n597 B.n92 256.663
R496 B.n597 B.n91 256.663
R497 B.n381 B.n380 256.663
R498 B.n381 B.n285 256.663
R499 B.n381 B.n286 256.663
R500 B.n381 B.n287 256.663
R501 B.n381 B.n288 256.663
R502 B.n381 B.n289 256.663
R503 B.n381 B.n290 256.663
R504 B.n381 B.n291 256.663
R505 B.n381 B.n292 256.663
R506 B.n381 B.n293 256.663
R507 B.n381 B.n294 256.663
R508 B.n381 B.n295 256.663
R509 B.n381 B.n296 256.663
R510 B.n381 B.n297 256.663
R511 B.n381 B.n298 256.663
R512 B.n381 B.n299 256.663
R513 B.n381 B.n300 256.663
R514 B.n381 B.n301 256.663
R515 B.n306 B.t21 238.73
R516 B.n304 B.t17 238.73
R517 B.n113 B.t10 238.73
R518 B.n110 B.t14 238.73
R519 B.n381 B.n281 193.179
R520 B.n598 B.n597 193.179
R521 B.n306 B.t23 170.602
R522 B.n110 B.t15 170.602
R523 B.n304 B.t20 170.602
R524 B.n113 B.t12 170.602
R525 B.n388 B.n280 163.367
R526 B.n388 B.n278 163.367
R527 B.n392 B.n278 163.367
R528 B.n392 B.n272 163.367
R529 B.n401 B.n272 163.367
R530 B.n401 B.n270 163.367
R531 B.n405 B.n270 163.367
R532 B.n405 B.n265 163.367
R533 B.n413 B.n265 163.367
R534 B.n413 B.n263 163.367
R535 B.n417 B.n263 163.367
R536 B.n417 B.n257 163.367
R537 B.n425 B.n257 163.367
R538 B.n425 B.n255 163.367
R539 B.n429 B.n255 163.367
R540 B.n429 B.n249 163.367
R541 B.n437 B.n249 163.367
R542 B.n437 B.n247 163.367
R543 B.n441 B.n247 163.367
R544 B.n441 B.n241 163.367
R545 B.n449 B.n241 163.367
R546 B.n449 B.n239 163.367
R547 B.n453 B.n239 163.367
R548 B.n453 B.n233 163.367
R549 B.n461 B.n233 163.367
R550 B.n461 B.n231 163.367
R551 B.n465 B.n231 163.367
R552 B.n465 B.n225 163.367
R553 B.n474 B.n225 163.367
R554 B.n474 B.n223 163.367
R555 B.n478 B.n223 163.367
R556 B.n478 B.n218 163.367
R557 B.n486 B.n218 163.367
R558 B.n486 B.n216 163.367
R559 B.n490 B.n216 163.367
R560 B.n490 B.n210 163.367
R561 B.n498 B.n210 163.367
R562 B.n498 B.n208 163.367
R563 B.n502 B.n208 163.367
R564 B.n502 B.n202 163.367
R565 B.n510 B.n202 163.367
R566 B.n510 B.n200 163.367
R567 B.n514 B.n200 163.367
R568 B.n514 B.n194 163.367
R569 B.n523 B.n194 163.367
R570 B.n523 B.n192 163.367
R571 B.n527 B.n192 163.367
R572 B.n527 B.n2 163.367
R573 B.n696 B.n2 163.367
R574 B.n696 B.n3 163.367
R575 B.n692 B.n3 163.367
R576 B.n692 B.n9 163.367
R577 B.n688 B.n9 163.367
R578 B.n688 B.n11 163.367
R579 B.n684 B.n11 163.367
R580 B.n684 B.n16 163.367
R581 B.n680 B.n16 163.367
R582 B.n680 B.n18 163.367
R583 B.n676 B.n18 163.367
R584 B.n676 B.n23 163.367
R585 B.n672 B.n23 163.367
R586 B.n672 B.n25 163.367
R587 B.n668 B.n25 163.367
R588 B.n668 B.n30 163.367
R589 B.n664 B.n30 163.367
R590 B.n664 B.n32 163.367
R591 B.n660 B.n32 163.367
R592 B.n660 B.n36 163.367
R593 B.n656 B.n36 163.367
R594 B.n656 B.n38 163.367
R595 B.n652 B.n38 163.367
R596 B.n652 B.n44 163.367
R597 B.n648 B.n44 163.367
R598 B.n648 B.n46 163.367
R599 B.n644 B.n46 163.367
R600 B.n644 B.n51 163.367
R601 B.n640 B.n51 163.367
R602 B.n640 B.n53 163.367
R603 B.n636 B.n53 163.367
R604 B.n636 B.n58 163.367
R605 B.n632 B.n58 163.367
R606 B.n632 B.n60 163.367
R607 B.n628 B.n60 163.367
R608 B.n628 B.n65 163.367
R609 B.n624 B.n65 163.367
R610 B.n624 B.n67 163.367
R611 B.n620 B.n67 163.367
R612 B.n620 B.n72 163.367
R613 B.n616 B.n72 163.367
R614 B.n616 B.n74 163.367
R615 B.n612 B.n74 163.367
R616 B.n612 B.n78 163.367
R617 B.n608 B.n78 163.367
R618 B.n608 B.n80 163.367
R619 B.n604 B.n80 163.367
R620 B.n604 B.n86 163.367
R621 B.n600 B.n86 163.367
R622 B.n600 B.n88 163.367
R623 B.n303 B.n302 163.367
R624 B.n374 B.n302 163.367
R625 B.n372 B.n371 163.367
R626 B.n368 B.n367 163.367
R627 B.n364 B.n363 163.367
R628 B.n360 B.n359 163.367
R629 B.n356 B.n355 163.367
R630 B.n351 B.n350 163.367
R631 B.n347 B.n346 163.367
R632 B.n343 B.n342 163.367
R633 B.n339 B.n338 163.367
R634 B.n335 B.n334 163.367
R635 B.n330 B.n329 163.367
R636 B.n326 B.n325 163.367
R637 B.n322 B.n321 163.367
R638 B.n318 B.n317 163.367
R639 B.n314 B.n313 163.367
R640 B.n310 B.n309 163.367
R641 B.n382 B.n284 163.367
R642 B.n386 B.n282 163.367
R643 B.n386 B.n276 163.367
R644 B.n394 B.n276 163.367
R645 B.n394 B.n274 163.367
R646 B.n398 B.n274 163.367
R647 B.n398 B.n269 163.367
R648 B.n407 B.n269 163.367
R649 B.n407 B.n267 163.367
R650 B.n411 B.n267 163.367
R651 B.n411 B.n261 163.367
R652 B.n419 B.n261 163.367
R653 B.n419 B.n259 163.367
R654 B.n423 B.n259 163.367
R655 B.n423 B.n252 163.367
R656 B.n431 B.n252 163.367
R657 B.n431 B.n250 163.367
R658 B.n435 B.n250 163.367
R659 B.n435 B.n245 163.367
R660 B.n443 B.n245 163.367
R661 B.n443 B.n243 163.367
R662 B.n447 B.n243 163.367
R663 B.n447 B.n237 163.367
R664 B.n455 B.n237 163.367
R665 B.n455 B.n235 163.367
R666 B.n459 B.n235 163.367
R667 B.n459 B.n229 163.367
R668 B.n467 B.n229 163.367
R669 B.n467 B.n227 163.367
R670 B.n471 B.n227 163.367
R671 B.n471 B.n222 163.367
R672 B.n480 B.n222 163.367
R673 B.n480 B.n220 163.367
R674 B.n484 B.n220 163.367
R675 B.n484 B.n214 163.367
R676 B.n492 B.n214 163.367
R677 B.n492 B.n212 163.367
R678 B.n496 B.n212 163.367
R679 B.n496 B.n206 163.367
R680 B.n504 B.n206 163.367
R681 B.n504 B.n204 163.367
R682 B.n508 B.n204 163.367
R683 B.n508 B.n198 163.367
R684 B.n516 B.n198 163.367
R685 B.n516 B.n196 163.367
R686 B.n521 B.n196 163.367
R687 B.n521 B.n190 163.367
R688 B.n529 B.n190 163.367
R689 B.n530 B.n529 163.367
R690 B.n530 B.n5 163.367
R691 B.n6 B.n5 163.367
R692 B.n7 B.n6 163.367
R693 B.n535 B.n7 163.367
R694 B.n535 B.n12 163.367
R695 B.n13 B.n12 163.367
R696 B.n14 B.n13 163.367
R697 B.n540 B.n14 163.367
R698 B.n540 B.n19 163.367
R699 B.n20 B.n19 163.367
R700 B.n21 B.n20 163.367
R701 B.n545 B.n21 163.367
R702 B.n545 B.n26 163.367
R703 B.n27 B.n26 163.367
R704 B.n28 B.n27 163.367
R705 B.n550 B.n28 163.367
R706 B.n550 B.n33 163.367
R707 B.n34 B.n33 163.367
R708 B.n35 B.n34 163.367
R709 B.n555 B.n35 163.367
R710 B.n555 B.n40 163.367
R711 B.n41 B.n40 163.367
R712 B.n42 B.n41 163.367
R713 B.n560 B.n42 163.367
R714 B.n560 B.n47 163.367
R715 B.n48 B.n47 163.367
R716 B.n49 B.n48 163.367
R717 B.n565 B.n49 163.367
R718 B.n565 B.n54 163.367
R719 B.n55 B.n54 163.367
R720 B.n56 B.n55 163.367
R721 B.n570 B.n56 163.367
R722 B.n570 B.n61 163.367
R723 B.n62 B.n61 163.367
R724 B.n63 B.n62 163.367
R725 B.n575 B.n63 163.367
R726 B.n575 B.n68 163.367
R727 B.n69 B.n68 163.367
R728 B.n70 B.n69 163.367
R729 B.n580 B.n70 163.367
R730 B.n580 B.n75 163.367
R731 B.n76 B.n75 163.367
R732 B.n77 B.n76 163.367
R733 B.n585 B.n77 163.367
R734 B.n585 B.n82 163.367
R735 B.n83 B.n82 163.367
R736 B.n84 B.n83 163.367
R737 B.n590 B.n84 163.367
R738 B.n590 B.n89 163.367
R739 B.n90 B.n89 163.367
R740 B.n120 B.n119 163.367
R741 B.n124 B.n123 163.367
R742 B.n128 B.n127 163.367
R743 B.n132 B.n131 163.367
R744 B.n136 B.n135 163.367
R745 B.n140 B.n139 163.367
R746 B.n144 B.n143 163.367
R747 B.n148 B.n147 163.367
R748 B.n152 B.n151 163.367
R749 B.n156 B.n155 163.367
R750 B.n160 B.n159 163.367
R751 B.n164 B.n163 163.367
R752 B.n168 B.n167 163.367
R753 B.n172 B.n171 163.367
R754 B.n176 B.n175 163.367
R755 B.n180 B.n179 163.367
R756 B.n184 B.n183 163.367
R757 B.n186 B.n109 163.367
R758 B.n307 B.t22 125.415
R759 B.n111 B.t16 125.415
R760 B.n305 B.t19 125.415
R761 B.n114 B.t13 125.415
R762 B.n387 B.n281 94.5046
R763 B.n387 B.n277 94.5046
R764 B.n393 B.n277 94.5046
R765 B.n393 B.n273 94.5046
R766 B.n400 B.n273 94.5046
R767 B.n400 B.n399 94.5046
R768 B.n406 B.n266 94.5046
R769 B.n412 B.n266 94.5046
R770 B.n412 B.n262 94.5046
R771 B.n418 B.n262 94.5046
R772 B.n418 B.n258 94.5046
R773 B.n424 B.n258 94.5046
R774 B.n424 B.n253 94.5046
R775 B.n430 B.n253 94.5046
R776 B.n430 B.n254 94.5046
R777 B.n436 B.n246 94.5046
R778 B.n442 B.n246 94.5046
R779 B.n442 B.n242 94.5046
R780 B.n448 B.n242 94.5046
R781 B.n448 B.n238 94.5046
R782 B.n454 B.n238 94.5046
R783 B.n460 B.n234 94.5046
R784 B.n460 B.n230 94.5046
R785 B.n466 B.n230 94.5046
R786 B.n466 B.n226 94.5046
R787 B.n473 B.n226 94.5046
R788 B.n473 B.n472 94.5046
R789 B.n479 B.n219 94.5046
R790 B.n485 B.n219 94.5046
R791 B.n485 B.n215 94.5046
R792 B.n491 B.n215 94.5046
R793 B.n491 B.n211 94.5046
R794 B.n497 B.n211 94.5046
R795 B.n503 B.n207 94.5046
R796 B.n503 B.n203 94.5046
R797 B.n509 B.n203 94.5046
R798 B.n509 B.n199 94.5046
R799 B.n515 B.n199 94.5046
R800 B.n522 B.n195 94.5046
R801 B.n522 B.n191 94.5046
R802 B.n528 B.n191 94.5046
R803 B.n528 B.n4 94.5046
R804 B.n695 B.n4 94.5046
R805 B.n695 B.n694 94.5046
R806 B.n694 B.n693 94.5046
R807 B.n693 B.n8 94.5046
R808 B.n687 B.n8 94.5046
R809 B.n687 B.n686 94.5046
R810 B.n685 B.n15 94.5046
R811 B.n679 B.n15 94.5046
R812 B.n679 B.n678 94.5046
R813 B.n678 B.n677 94.5046
R814 B.n677 B.n22 94.5046
R815 B.n671 B.n670 94.5046
R816 B.n670 B.n669 94.5046
R817 B.n669 B.n29 94.5046
R818 B.n663 B.n29 94.5046
R819 B.n663 B.n662 94.5046
R820 B.n662 B.n661 94.5046
R821 B.n655 B.n39 94.5046
R822 B.n655 B.n654 94.5046
R823 B.n654 B.n653 94.5046
R824 B.n653 B.n43 94.5046
R825 B.n647 B.n43 94.5046
R826 B.n647 B.n646 94.5046
R827 B.n645 B.n50 94.5046
R828 B.n639 B.n50 94.5046
R829 B.n639 B.n638 94.5046
R830 B.n638 B.n637 94.5046
R831 B.n637 B.n57 94.5046
R832 B.n631 B.n57 94.5046
R833 B.n630 B.n629 94.5046
R834 B.n629 B.n64 94.5046
R835 B.n623 B.n64 94.5046
R836 B.n623 B.n622 94.5046
R837 B.n622 B.n621 94.5046
R838 B.n621 B.n71 94.5046
R839 B.n615 B.n71 94.5046
R840 B.n615 B.n614 94.5046
R841 B.n614 B.n613 94.5046
R842 B.n607 B.n81 94.5046
R843 B.n607 B.n606 94.5046
R844 B.n606 B.n605 94.5046
R845 B.n605 B.n85 94.5046
R846 B.n599 B.n85 94.5046
R847 B.n599 B.n598 94.5046
R848 B.n515 B.t9 91.7251
R849 B.t7 B.n685 91.7251
R850 B.t3 B.n207 83.3865
R851 B.t1 B.n22 83.3865
R852 B.n380 B.n379 71.676
R853 B.n374 B.n285 71.676
R854 B.n371 B.n286 71.676
R855 B.n367 B.n287 71.676
R856 B.n363 B.n288 71.676
R857 B.n359 B.n289 71.676
R858 B.n355 B.n290 71.676
R859 B.n350 B.n291 71.676
R860 B.n346 B.n292 71.676
R861 B.n342 B.n293 71.676
R862 B.n338 B.n294 71.676
R863 B.n334 B.n295 71.676
R864 B.n329 B.n296 71.676
R865 B.n325 B.n297 71.676
R866 B.n321 B.n298 71.676
R867 B.n317 B.n299 71.676
R868 B.n313 B.n300 71.676
R869 B.n309 B.n301 71.676
R870 B.n116 B.n91 71.676
R871 B.n120 B.n92 71.676
R872 B.n124 B.n93 71.676
R873 B.n128 B.n94 71.676
R874 B.n132 B.n95 71.676
R875 B.n136 B.n96 71.676
R876 B.n140 B.n97 71.676
R877 B.n144 B.n98 71.676
R878 B.n148 B.n99 71.676
R879 B.n152 B.n100 71.676
R880 B.n156 B.n101 71.676
R881 B.n160 B.n102 71.676
R882 B.n164 B.n103 71.676
R883 B.n168 B.n104 71.676
R884 B.n172 B.n105 71.676
R885 B.n176 B.n106 71.676
R886 B.n180 B.n107 71.676
R887 B.n184 B.n108 71.676
R888 B.n596 B.n109 71.676
R889 B.n596 B.n595 71.676
R890 B.n186 B.n108 71.676
R891 B.n183 B.n107 71.676
R892 B.n179 B.n106 71.676
R893 B.n175 B.n105 71.676
R894 B.n171 B.n104 71.676
R895 B.n167 B.n103 71.676
R896 B.n163 B.n102 71.676
R897 B.n159 B.n101 71.676
R898 B.n155 B.n100 71.676
R899 B.n151 B.n99 71.676
R900 B.n147 B.n98 71.676
R901 B.n143 B.n97 71.676
R902 B.n139 B.n96 71.676
R903 B.n135 B.n95 71.676
R904 B.n131 B.n94 71.676
R905 B.n127 B.n93 71.676
R906 B.n123 B.n92 71.676
R907 B.n119 B.n91 71.676
R908 B.n380 B.n303 71.676
R909 B.n372 B.n285 71.676
R910 B.n368 B.n286 71.676
R911 B.n364 B.n287 71.676
R912 B.n360 B.n288 71.676
R913 B.n356 B.n289 71.676
R914 B.n351 B.n290 71.676
R915 B.n347 B.n291 71.676
R916 B.n343 B.n292 71.676
R917 B.n339 B.n293 71.676
R918 B.n335 B.n294 71.676
R919 B.n330 B.n295 71.676
R920 B.n326 B.n296 71.676
R921 B.n322 B.n297 71.676
R922 B.n318 B.n298 71.676
R923 B.n314 B.n299 71.676
R924 B.n310 B.n300 71.676
R925 B.n301 B.n284 71.676
R926 B.n479 B.t2 69.4888
R927 B.n661 B.t6 69.4888
R928 B.n332 B.n307 59.5399
R929 B.n353 B.n305 59.5399
R930 B.n115 B.n114 59.5399
R931 B.n112 B.n111 59.5399
R932 B.t5 B.n234 55.5912
R933 B.n646 B.t8 55.5912
R934 B.n254 B.t0 52.8116
R935 B.t4 B.n630 52.8116
R936 B.n399 B.t18 47.2526
R937 B.n406 B.t18 47.2526
R938 B.n613 B.t11 47.2526
R939 B.n81 B.t11 47.2526
R940 B.n307 B.n306 45.1884
R941 B.n305 B.n304 45.1884
R942 B.n114 B.n113 45.1884
R943 B.n111 B.n110 45.1884
R944 B.n436 B.t0 41.6935
R945 B.n631 B.t4 41.6935
R946 B.n454 B.t5 38.914
R947 B.t8 B.n645 38.914
R948 B.n117 B.n87 33.5615
R949 B.n594 B.n593 33.5615
R950 B.n384 B.n383 33.5615
R951 B.n378 B.n279 33.5615
R952 B.n472 B.t2 25.0163
R953 B.n39 B.t6 25.0163
R954 B B.n697 18.0485
R955 B.n497 B.t3 11.1186
R956 B.n671 B.t1 11.1186
R957 B.n118 B.n117 10.6151
R958 B.n121 B.n118 10.6151
R959 B.n122 B.n121 10.6151
R960 B.n125 B.n122 10.6151
R961 B.n126 B.n125 10.6151
R962 B.n129 B.n126 10.6151
R963 B.n130 B.n129 10.6151
R964 B.n133 B.n130 10.6151
R965 B.n134 B.n133 10.6151
R966 B.n137 B.n134 10.6151
R967 B.n138 B.n137 10.6151
R968 B.n141 B.n138 10.6151
R969 B.n142 B.n141 10.6151
R970 B.n146 B.n145 10.6151
R971 B.n149 B.n146 10.6151
R972 B.n150 B.n149 10.6151
R973 B.n153 B.n150 10.6151
R974 B.n154 B.n153 10.6151
R975 B.n157 B.n154 10.6151
R976 B.n158 B.n157 10.6151
R977 B.n161 B.n158 10.6151
R978 B.n162 B.n161 10.6151
R979 B.n166 B.n165 10.6151
R980 B.n169 B.n166 10.6151
R981 B.n170 B.n169 10.6151
R982 B.n173 B.n170 10.6151
R983 B.n174 B.n173 10.6151
R984 B.n177 B.n174 10.6151
R985 B.n178 B.n177 10.6151
R986 B.n181 B.n178 10.6151
R987 B.n182 B.n181 10.6151
R988 B.n185 B.n182 10.6151
R989 B.n187 B.n185 10.6151
R990 B.n188 B.n187 10.6151
R991 B.n594 B.n188 10.6151
R992 B.n385 B.n384 10.6151
R993 B.n385 B.n275 10.6151
R994 B.n395 B.n275 10.6151
R995 B.n396 B.n395 10.6151
R996 B.n397 B.n396 10.6151
R997 B.n397 B.n268 10.6151
R998 B.n408 B.n268 10.6151
R999 B.n409 B.n408 10.6151
R1000 B.n410 B.n409 10.6151
R1001 B.n410 B.n260 10.6151
R1002 B.n420 B.n260 10.6151
R1003 B.n421 B.n420 10.6151
R1004 B.n422 B.n421 10.6151
R1005 B.n422 B.n251 10.6151
R1006 B.n432 B.n251 10.6151
R1007 B.n433 B.n432 10.6151
R1008 B.n434 B.n433 10.6151
R1009 B.n434 B.n244 10.6151
R1010 B.n444 B.n244 10.6151
R1011 B.n445 B.n444 10.6151
R1012 B.n446 B.n445 10.6151
R1013 B.n446 B.n236 10.6151
R1014 B.n456 B.n236 10.6151
R1015 B.n457 B.n456 10.6151
R1016 B.n458 B.n457 10.6151
R1017 B.n458 B.n228 10.6151
R1018 B.n468 B.n228 10.6151
R1019 B.n469 B.n468 10.6151
R1020 B.n470 B.n469 10.6151
R1021 B.n470 B.n221 10.6151
R1022 B.n481 B.n221 10.6151
R1023 B.n482 B.n481 10.6151
R1024 B.n483 B.n482 10.6151
R1025 B.n483 B.n213 10.6151
R1026 B.n493 B.n213 10.6151
R1027 B.n494 B.n493 10.6151
R1028 B.n495 B.n494 10.6151
R1029 B.n495 B.n205 10.6151
R1030 B.n505 B.n205 10.6151
R1031 B.n506 B.n505 10.6151
R1032 B.n507 B.n506 10.6151
R1033 B.n507 B.n197 10.6151
R1034 B.n517 B.n197 10.6151
R1035 B.n518 B.n517 10.6151
R1036 B.n520 B.n518 10.6151
R1037 B.n520 B.n519 10.6151
R1038 B.n519 B.n189 10.6151
R1039 B.n531 B.n189 10.6151
R1040 B.n532 B.n531 10.6151
R1041 B.n533 B.n532 10.6151
R1042 B.n534 B.n533 10.6151
R1043 B.n536 B.n534 10.6151
R1044 B.n537 B.n536 10.6151
R1045 B.n538 B.n537 10.6151
R1046 B.n539 B.n538 10.6151
R1047 B.n541 B.n539 10.6151
R1048 B.n542 B.n541 10.6151
R1049 B.n543 B.n542 10.6151
R1050 B.n544 B.n543 10.6151
R1051 B.n546 B.n544 10.6151
R1052 B.n547 B.n546 10.6151
R1053 B.n548 B.n547 10.6151
R1054 B.n549 B.n548 10.6151
R1055 B.n551 B.n549 10.6151
R1056 B.n552 B.n551 10.6151
R1057 B.n553 B.n552 10.6151
R1058 B.n554 B.n553 10.6151
R1059 B.n556 B.n554 10.6151
R1060 B.n557 B.n556 10.6151
R1061 B.n558 B.n557 10.6151
R1062 B.n559 B.n558 10.6151
R1063 B.n561 B.n559 10.6151
R1064 B.n562 B.n561 10.6151
R1065 B.n563 B.n562 10.6151
R1066 B.n564 B.n563 10.6151
R1067 B.n566 B.n564 10.6151
R1068 B.n567 B.n566 10.6151
R1069 B.n568 B.n567 10.6151
R1070 B.n569 B.n568 10.6151
R1071 B.n571 B.n569 10.6151
R1072 B.n572 B.n571 10.6151
R1073 B.n573 B.n572 10.6151
R1074 B.n574 B.n573 10.6151
R1075 B.n576 B.n574 10.6151
R1076 B.n577 B.n576 10.6151
R1077 B.n578 B.n577 10.6151
R1078 B.n579 B.n578 10.6151
R1079 B.n581 B.n579 10.6151
R1080 B.n582 B.n581 10.6151
R1081 B.n583 B.n582 10.6151
R1082 B.n584 B.n583 10.6151
R1083 B.n586 B.n584 10.6151
R1084 B.n587 B.n586 10.6151
R1085 B.n588 B.n587 10.6151
R1086 B.n589 B.n588 10.6151
R1087 B.n591 B.n589 10.6151
R1088 B.n592 B.n591 10.6151
R1089 B.n593 B.n592 10.6151
R1090 B.n378 B.n377 10.6151
R1091 B.n377 B.n376 10.6151
R1092 B.n376 B.n375 10.6151
R1093 B.n375 B.n373 10.6151
R1094 B.n373 B.n370 10.6151
R1095 B.n370 B.n369 10.6151
R1096 B.n369 B.n366 10.6151
R1097 B.n366 B.n365 10.6151
R1098 B.n365 B.n362 10.6151
R1099 B.n362 B.n361 10.6151
R1100 B.n361 B.n358 10.6151
R1101 B.n358 B.n357 10.6151
R1102 B.n357 B.n354 10.6151
R1103 B.n352 B.n349 10.6151
R1104 B.n349 B.n348 10.6151
R1105 B.n348 B.n345 10.6151
R1106 B.n345 B.n344 10.6151
R1107 B.n344 B.n341 10.6151
R1108 B.n341 B.n340 10.6151
R1109 B.n340 B.n337 10.6151
R1110 B.n337 B.n336 10.6151
R1111 B.n336 B.n333 10.6151
R1112 B.n331 B.n328 10.6151
R1113 B.n328 B.n327 10.6151
R1114 B.n327 B.n324 10.6151
R1115 B.n324 B.n323 10.6151
R1116 B.n323 B.n320 10.6151
R1117 B.n320 B.n319 10.6151
R1118 B.n319 B.n316 10.6151
R1119 B.n316 B.n315 10.6151
R1120 B.n315 B.n312 10.6151
R1121 B.n312 B.n311 10.6151
R1122 B.n311 B.n308 10.6151
R1123 B.n308 B.n283 10.6151
R1124 B.n383 B.n283 10.6151
R1125 B.n389 B.n279 10.6151
R1126 B.n390 B.n389 10.6151
R1127 B.n391 B.n390 10.6151
R1128 B.n391 B.n271 10.6151
R1129 B.n402 B.n271 10.6151
R1130 B.n403 B.n402 10.6151
R1131 B.n404 B.n403 10.6151
R1132 B.n404 B.n264 10.6151
R1133 B.n414 B.n264 10.6151
R1134 B.n415 B.n414 10.6151
R1135 B.n416 B.n415 10.6151
R1136 B.n416 B.n256 10.6151
R1137 B.n426 B.n256 10.6151
R1138 B.n427 B.n426 10.6151
R1139 B.n428 B.n427 10.6151
R1140 B.n428 B.n248 10.6151
R1141 B.n438 B.n248 10.6151
R1142 B.n439 B.n438 10.6151
R1143 B.n440 B.n439 10.6151
R1144 B.n440 B.n240 10.6151
R1145 B.n450 B.n240 10.6151
R1146 B.n451 B.n450 10.6151
R1147 B.n452 B.n451 10.6151
R1148 B.n452 B.n232 10.6151
R1149 B.n462 B.n232 10.6151
R1150 B.n463 B.n462 10.6151
R1151 B.n464 B.n463 10.6151
R1152 B.n464 B.n224 10.6151
R1153 B.n475 B.n224 10.6151
R1154 B.n476 B.n475 10.6151
R1155 B.n477 B.n476 10.6151
R1156 B.n477 B.n217 10.6151
R1157 B.n487 B.n217 10.6151
R1158 B.n488 B.n487 10.6151
R1159 B.n489 B.n488 10.6151
R1160 B.n489 B.n209 10.6151
R1161 B.n499 B.n209 10.6151
R1162 B.n500 B.n499 10.6151
R1163 B.n501 B.n500 10.6151
R1164 B.n501 B.n201 10.6151
R1165 B.n511 B.n201 10.6151
R1166 B.n512 B.n511 10.6151
R1167 B.n513 B.n512 10.6151
R1168 B.n513 B.n193 10.6151
R1169 B.n524 B.n193 10.6151
R1170 B.n525 B.n524 10.6151
R1171 B.n526 B.n525 10.6151
R1172 B.n526 B.n0 10.6151
R1173 B.n691 B.n1 10.6151
R1174 B.n691 B.n690 10.6151
R1175 B.n690 B.n689 10.6151
R1176 B.n689 B.n10 10.6151
R1177 B.n683 B.n10 10.6151
R1178 B.n683 B.n682 10.6151
R1179 B.n682 B.n681 10.6151
R1180 B.n681 B.n17 10.6151
R1181 B.n675 B.n17 10.6151
R1182 B.n675 B.n674 10.6151
R1183 B.n674 B.n673 10.6151
R1184 B.n673 B.n24 10.6151
R1185 B.n667 B.n24 10.6151
R1186 B.n667 B.n666 10.6151
R1187 B.n666 B.n665 10.6151
R1188 B.n665 B.n31 10.6151
R1189 B.n659 B.n31 10.6151
R1190 B.n659 B.n658 10.6151
R1191 B.n658 B.n657 10.6151
R1192 B.n657 B.n37 10.6151
R1193 B.n651 B.n37 10.6151
R1194 B.n651 B.n650 10.6151
R1195 B.n650 B.n649 10.6151
R1196 B.n649 B.n45 10.6151
R1197 B.n643 B.n45 10.6151
R1198 B.n643 B.n642 10.6151
R1199 B.n642 B.n641 10.6151
R1200 B.n641 B.n52 10.6151
R1201 B.n635 B.n52 10.6151
R1202 B.n635 B.n634 10.6151
R1203 B.n634 B.n633 10.6151
R1204 B.n633 B.n59 10.6151
R1205 B.n627 B.n59 10.6151
R1206 B.n627 B.n626 10.6151
R1207 B.n626 B.n625 10.6151
R1208 B.n625 B.n66 10.6151
R1209 B.n619 B.n66 10.6151
R1210 B.n619 B.n618 10.6151
R1211 B.n618 B.n617 10.6151
R1212 B.n617 B.n73 10.6151
R1213 B.n611 B.n73 10.6151
R1214 B.n611 B.n610 10.6151
R1215 B.n610 B.n609 10.6151
R1216 B.n609 B.n79 10.6151
R1217 B.n603 B.n79 10.6151
R1218 B.n603 B.n602 10.6151
R1219 B.n602 B.n601 10.6151
R1220 B.n601 B.n87 10.6151
R1221 B.n142 B.n115 9.36635
R1222 B.n165 B.n112 9.36635
R1223 B.n354 B.n353 9.36635
R1224 B.n332 B.n331 9.36635
R1225 B.n697 B.n0 2.81026
R1226 B.n697 B.n1 2.81026
R1227 B.t9 B.n195 2.78003
R1228 B.n686 B.t7 2.78003
R1229 B.n145 B.n115 1.24928
R1230 B.n162 B.n112 1.24928
R1231 B.n353 B.n352 1.24928
R1232 B.n333 B.n332 1.24928
R1233 VP.n20 VP.n19 161.3
R1234 VP.n21 VP.n16 161.3
R1235 VP.n23 VP.n22 161.3
R1236 VP.n24 VP.n15 161.3
R1237 VP.n26 VP.n25 161.3
R1238 VP.n28 VP.n14 161.3
R1239 VP.n30 VP.n29 161.3
R1240 VP.n31 VP.n13 161.3
R1241 VP.n33 VP.n32 161.3
R1242 VP.n34 VP.n12 161.3
R1243 VP.n37 VP.n36 161.3
R1244 VP.n38 VP.n11 161.3
R1245 VP.n40 VP.n39 161.3
R1246 VP.n41 VP.n10 161.3
R1247 VP.n74 VP.n0 161.3
R1248 VP.n73 VP.n72 161.3
R1249 VP.n71 VP.n1 161.3
R1250 VP.n70 VP.n69 161.3
R1251 VP.n67 VP.n2 161.3
R1252 VP.n66 VP.n65 161.3
R1253 VP.n64 VP.n3 161.3
R1254 VP.n63 VP.n62 161.3
R1255 VP.n61 VP.n4 161.3
R1256 VP.n59 VP.n58 161.3
R1257 VP.n57 VP.n5 161.3
R1258 VP.n56 VP.n55 161.3
R1259 VP.n54 VP.n6 161.3
R1260 VP.n53 VP.n52 161.3
R1261 VP.n51 VP.n50 161.3
R1262 VP.n49 VP.n8 161.3
R1263 VP.n48 VP.n47 161.3
R1264 VP.n46 VP.n9 161.3
R1265 VP.n45 VP.n44 90.6446
R1266 VP.n76 VP.n75 90.6446
R1267 VP.n43 VP.n42 90.6446
R1268 VP.n18 VP.n17 65.7074
R1269 VP.n18 VP.t4 62.1016
R1270 VP.n73 VP.n1 56.4773
R1271 VP.n49 VP.n48 56.4773
R1272 VP.n40 VP.n11 56.4773
R1273 VP.n55 VP.n5 48.6874
R1274 VP.n62 VP.n3 48.6874
R1275 VP.n29 VP.n13 48.6874
R1276 VP.n22 VP.n15 48.6874
R1277 VP.n45 VP.n43 42.7912
R1278 VP.n55 VP.n54 32.1338
R1279 VP.n66 VP.n3 32.1338
R1280 VP.n33 VP.n13 32.1338
R1281 VP.n22 VP.n21 32.1338
R1282 VP.n44 VP.t5 31.8125
R1283 VP.n7 VP.t9 31.8125
R1284 VP.n60 VP.t2 31.8125
R1285 VP.n68 VP.t3 31.8125
R1286 VP.n75 VP.t7 31.8125
R1287 VP.n42 VP.t0 31.8125
R1288 VP.n35 VP.t6 31.8125
R1289 VP.n27 VP.t1 31.8125
R1290 VP.n17 VP.t8 31.8125
R1291 VP.n48 VP.n9 24.3439
R1292 VP.n50 VP.n49 24.3439
R1293 VP.n54 VP.n53 24.3439
R1294 VP.n59 VP.n5 24.3439
R1295 VP.n62 VP.n61 24.3439
R1296 VP.n67 VP.n66 24.3439
R1297 VP.n69 VP.n1 24.3439
R1298 VP.n74 VP.n73 24.3439
R1299 VP.n41 VP.n40 24.3439
R1300 VP.n34 VP.n33 24.3439
R1301 VP.n36 VP.n11 24.3439
R1302 VP.n26 VP.n15 24.3439
R1303 VP.n29 VP.n28 24.3439
R1304 VP.n21 VP.n20 24.3439
R1305 VP.n50 VP.n7 20.449
R1306 VP.n69 VP.n68 20.449
R1307 VP.n36 VP.n35 20.449
R1308 VP.n44 VP.n9 19.9621
R1309 VP.n75 VP.n74 19.9621
R1310 VP.n42 VP.n41 19.9621
R1311 VP.n19 VP.n18 13.3187
R1312 VP.n60 VP.n59 12.1722
R1313 VP.n61 VP.n60 12.1722
R1314 VP.n27 VP.n26 12.1722
R1315 VP.n28 VP.n27 12.1722
R1316 VP.n53 VP.n7 3.89545
R1317 VP.n68 VP.n67 3.89545
R1318 VP.n35 VP.n34 3.89545
R1319 VP.n20 VP.n17 3.89545
R1320 VP.n43 VP.n10 0.278398
R1321 VP.n46 VP.n45 0.278398
R1322 VP.n76 VP.n0 0.278398
R1323 VP.n19 VP.n16 0.189894
R1324 VP.n23 VP.n16 0.189894
R1325 VP.n24 VP.n23 0.189894
R1326 VP.n25 VP.n24 0.189894
R1327 VP.n25 VP.n14 0.189894
R1328 VP.n30 VP.n14 0.189894
R1329 VP.n31 VP.n30 0.189894
R1330 VP.n32 VP.n31 0.189894
R1331 VP.n32 VP.n12 0.189894
R1332 VP.n37 VP.n12 0.189894
R1333 VP.n38 VP.n37 0.189894
R1334 VP.n39 VP.n38 0.189894
R1335 VP.n39 VP.n10 0.189894
R1336 VP.n47 VP.n46 0.189894
R1337 VP.n47 VP.n8 0.189894
R1338 VP.n51 VP.n8 0.189894
R1339 VP.n52 VP.n51 0.189894
R1340 VP.n52 VP.n6 0.189894
R1341 VP.n56 VP.n6 0.189894
R1342 VP.n57 VP.n56 0.189894
R1343 VP.n58 VP.n57 0.189894
R1344 VP.n58 VP.n4 0.189894
R1345 VP.n63 VP.n4 0.189894
R1346 VP.n64 VP.n63 0.189894
R1347 VP.n65 VP.n64 0.189894
R1348 VP.n65 VP.n2 0.189894
R1349 VP.n70 VP.n2 0.189894
R1350 VP.n71 VP.n70 0.189894
R1351 VP.n72 VP.n71 0.189894
R1352 VP.n72 VP.n0 0.189894
R1353 VP VP.n76 0.153422
R1354 VTAIL.n56 VTAIL.n50 289.615
R1355 VTAIL.n8 VTAIL.n2 289.615
R1356 VTAIL.n44 VTAIL.n38 289.615
R1357 VTAIL.n28 VTAIL.n22 289.615
R1358 VTAIL.n55 VTAIL.n54 185
R1359 VTAIL.n57 VTAIL.n56 185
R1360 VTAIL.n7 VTAIL.n6 185
R1361 VTAIL.n9 VTAIL.n8 185
R1362 VTAIL.n45 VTAIL.n44 185
R1363 VTAIL.n43 VTAIL.n42 185
R1364 VTAIL.n29 VTAIL.n28 185
R1365 VTAIL.n27 VTAIL.n26 185
R1366 VTAIL.n53 VTAIL.t5 153.582
R1367 VTAIL.n5 VTAIL.t15 153.582
R1368 VTAIL.n41 VTAIL.t13 153.582
R1369 VTAIL.n25 VTAIL.t3 153.582
R1370 VTAIL.n56 VTAIL.n55 104.615
R1371 VTAIL.n8 VTAIL.n7 104.615
R1372 VTAIL.n44 VTAIL.n43 104.615
R1373 VTAIL.n28 VTAIL.n27 104.615
R1374 VTAIL.n63 VTAIL.n62 67.4121
R1375 VTAIL.n1 VTAIL.n0 67.4121
R1376 VTAIL.n15 VTAIL.n14 67.4121
R1377 VTAIL.n17 VTAIL.n16 67.4121
R1378 VTAIL.n37 VTAIL.n36 67.4121
R1379 VTAIL.n35 VTAIL.n34 67.4121
R1380 VTAIL.n21 VTAIL.n20 67.4121
R1381 VTAIL.n19 VTAIL.n18 67.4121
R1382 VTAIL.n55 VTAIL.t5 52.3082
R1383 VTAIL.n7 VTAIL.t15 52.3082
R1384 VTAIL.n43 VTAIL.t13 52.3082
R1385 VTAIL.n27 VTAIL.t3 52.3082
R1386 VTAIL.n61 VTAIL.n60 29.8581
R1387 VTAIL.n13 VTAIL.n12 29.8581
R1388 VTAIL.n49 VTAIL.n48 29.8581
R1389 VTAIL.n33 VTAIL.n32 29.8581
R1390 VTAIL.n19 VTAIL.n17 18.66
R1391 VTAIL.n61 VTAIL.n49 16.6514
R1392 VTAIL.n54 VTAIL.n53 10.1164
R1393 VTAIL.n6 VTAIL.n5 10.1164
R1394 VTAIL.n42 VTAIL.n41 10.1164
R1395 VTAIL.n26 VTAIL.n25 10.1164
R1396 VTAIL.n60 VTAIL.n59 9.45567
R1397 VTAIL.n12 VTAIL.n11 9.45567
R1398 VTAIL.n48 VTAIL.n47 9.45567
R1399 VTAIL.n32 VTAIL.n31 9.45567
R1400 VTAIL.n52 VTAIL.n51 9.3005
R1401 VTAIL.n59 VTAIL.n58 9.3005
R1402 VTAIL.n4 VTAIL.n3 9.3005
R1403 VTAIL.n11 VTAIL.n10 9.3005
R1404 VTAIL.n40 VTAIL.n39 9.3005
R1405 VTAIL.n47 VTAIL.n46 9.3005
R1406 VTAIL.n31 VTAIL.n30 9.3005
R1407 VTAIL.n24 VTAIL.n23 9.3005
R1408 VTAIL.n60 VTAIL.n50 8.92171
R1409 VTAIL.n12 VTAIL.n2 8.92171
R1410 VTAIL.n48 VTAIL.n38 8.92171
R1411 VTAIL.n32 VTAIL.n22 8.92171
R1412 VTAIL.n58 VTAIL.n57 8.14595
R1413 VTAIL.n10 VTAIL.n9 8.14595
R1414 VTAIL.n46 VTAIL.n45 8.14595
R1415 VTAIL.n30 VTAIL.n29 8.14595
R1416 VTAIL.n62 VTAIL.t4 7.5005
R1417 VTAIL.n62 VTAIL.t7 7.5005
R1418 VTAIL.n0 VTAIL.t2 7.5005
R1419 VTAIL.n0 VTAIL.t8 7.5005
R1420 VTAIL.n14 VTAIL.t14 7.5005
R1421 VTAIL.n14 VTAIL.t18 7.5005
R1422 VTAIL.n16 VTAIL.t12 7.5005
R1423 VTAIL.n16 VTAIL.t11 7.5005
R1424 VTAIL.n36 VTAIL.t10 7.5005
R1425 VTAIL.n36 VTAIL.t17 7.5005
R1426 VTAIL.n34 VTAIL.t19 7.5005
R1427 VTAIL.n34 VTAIL.t16 7.5005
R1428 VTAIL.n20 VTAIL.t0 7.5005
R1429 VTAIL.n20 VTAIL.t1 7.5005
R1430 VTAIL.n18 VTAIL.t6 7.5005
R1431 VTAIL.n18 VTAIL.t9 7.5005
R1432 VTAIL.n54 VTAIL.n52 7.3702
R1433 VTAIL.n6 VTAIL.n4 7.3702
R1434 VTAIL.n42 VTAIL.n40 7.3702
R1435 VTAIL.n26 VTAIL.n24 7.3702
R1436 VTAIL.n57 VTAIL.n52 5.81868
R1437 VTAIL.n9 VTAIL.n4 5.81868
R1438 VTAIL.n45 VTAIL.n40 5.81868
R1439 VTAIL.n29 VTAIL.n24 5.81868
R1440 VTAIL.n58 VTAIL.n50 5.04292
R1441 VTAIL.n10 VTAIL.n2 5.04292
R1442 VTAIL.n46 VTAIL.n38 5.04292
R1443 VTAIL.n30 VTAIL.n22 5.04292
R1444 VTAIL.n25 VTAIL.n23 3.00987
R1445 VTAIL.n53 VTAIL.n51 3.00987
R1446 VTAIL.n5 VTAIL.n3 3.00987
R1447 VTAIL.n41 VTAIL.n39 3.00987
R1448 VTAIL.n21 VTAIL.n19 2.00912
R1449 VTAIL.n33 VTAIL.n21 2.00912
R1450 VTAIL.n37 VTAIL.n35 2.00912
R1451 VTAIL.n49 VTAIL.n37 2.00912
R1452 VTAIL.n17 VTAIL.n15 2.00912
R1453 VTAIL.n15 VTAIL.n13 2.00912
R1454 VTAIL.n63 VTAIL.n61 2.00912
R1455 VTAIL VTAIL.n1 1.56516
R1456 VTAIL.n35 VTAIL.n33 1.47464
R1457 VTAIL.n13 VTAIL.n1 1.47464
R1458 VTAIL VTAIL.n63 0.444466
R1459 VTAIL.n59 VTAIL.n51 0.155672
R1460 VTAIL.n11 VTAIL.n3 0.155672
R1461 VTAIL.n47 VTAIL.n39 0.155672
R1462 VTAIL.n31 VTAIL.n23 0.155672
R1463 VDD1.n6 VDD1.n0 289.615
R1464 VDD1.n19 VDD1.n13 289.615
R1465 VDD1.n7 VDD1.n6 185
R1466 VDD1.n5 VDD1.n4 185
R1467 VDD1.n18 VDD1.n17 185
R1468 VDD1.n20 VDD1.n19 185
R1469 VDD1.n16 VDD1.t4 153.582
R1470 VDD1.n3 VDD1.t5 153.582
R1471 VDD1.n6 VDD1.n5 104.615
R1472 VDD1.n19 VDD1.n18 104.615
R1473 VDD1.n27 VDD1.n26 85.542
R1474 VDD1.n25 VDD1.n24 84.0909
R1475 VDD1.n29 VDD1.n28 84.0909
R1476 VDD1.n12 VDD1.n11 84.0909
R1477 VDD1.n5 VDD1.t5 52.3082
R1478 VDD1.n18 VDD1.t4 52.3082
R1479 VDD1.n12 VDD1.n10 48.5455
R1480 VDD1.n25 VDD1.n23 48.5455
R1481 VDD1.n29 VDD1.n27 37.1194
R1482 VDD1.n4 VDD1.n3 10.1164
R1483 VDD1.n17 VDD1.n16 10.1164
R1484 VDD1.n10 VDD1.n9 9.45567
R1485 VDD1.n23 VDD1.n22 9.45567
R1486 VDD1.n9 VDD1.n8 9.3005
R1487 VDD1.n2 VDD1.n1 9.3005
R1488 VDD1.n15 VDD1.n14 9.3005
R1489 VDD1.n22 VDD1.n21 9.3005
R1490 VDD1.n10 VDD1.n0 8.92171
R1491 VDD1.n23 VDD1.n13 8.92171
R1492 VDD1.n8 VDD1.n7 8.14595
R1493 VDD1.n21 VDD1.n20 8.14595
R1494 VDD1.n28 VDD1.t3 7.5005
R1495 VDD1.n28 VDD1.t9 7.5005
R1496 VDD1.n11 VDD1.t1 7.5005
R1497 VDD1.n11 VDD1.t8 7.5005
R1498 VDD1.n26 VDD1.t6 7.5005
R1499 VDD1.n26 VDD1.t2 7.5005
R1500 VDD1.n24 VDD1.t0 7.5005
R1501 VDD1.n24 VDD1.t7 7.5005
R1502 VDD1.n4 VDD1.n2 7.3702
R1503 VDD1.n17 VDD1.n15 7.3702
R1504 VDD1.n7 VDD1.n2 5.81868
R1505 VDD1.n20 VDD1.n15 5.81868
R1506 VDD1.n8 VDD1.n0 5.04292
R1507 VDD1.n21 VDD1.n13 5.04292
R1508 VDD1.n3 VDD1.n1 3.00987
R1509 VDD1.n16 VDD1.n14 3.00987
R1510 VDD1 VDD1.n29 1.44878
R1511 VDD1 VDD1.n12 0.560845
R1512 VDD1.n27 VDD1.n25 0.447309
R1513 VDD1.n9 VDD1.n1 0.155672
R1514 VDD1.n22 VDD1.n14 0.155672
R1515 VN.n65 VN.n34 161.3
R1516 VN.n64 VN.n63 161.3
R1517 VN.n62 VN.n35 161.3
R1518 VN.n61 VN.n60 161.3
R1519 VN.n58 VN.n36 161.3
R1520 VN.n57 VN.n56 161.3
R1521 VN.n55 VN.n37 161.3
R1522 VN.n54 VN.n53 161.3
R1523 VN.n52 VN.n38 161.3
R1524 VN.n50 VN.n49 161.3
R1525 VN.n48 VN.n39 161.3
R1526 VN.n47 VN.n46 161.3
R1527 VN.n45 VN.n40 161.3
R1528 VN.n44 VN.n43 161.3
R1529 VN.n31 VN.n0 161.3
R1530 VN.n30 VN.n29 161.3
R1531 VN.n28 VN.n1 161.3
R1532 VN.n27 VN.n26 161.3
R1533 VN.n24 VN.n2 161.3
R1534 VN.n23 VN.n22 161.3
R1535 VN.n21 VN.n3 161.3
R1536 VN.n20 VN.n19 161.3
R1537 VN.n18 VN.n4 161.3
R1538 VN.n16 VN.n15 161.3
R1539 VN.n14 VN.n5 161.3
R1540 VN.n13 VN.n12 161.3
R1541 VN.n11 VN.n6 161.3
R1542 VN.n10 VN.n9 161.3
R1543 VN.n33 VN.n32 90.6446
R1544 VN.n67 VN.n66 90.6446
R1545 VN.n8 VN.n7 65.7074
R1546 VN.n42 VN.n41 65.7074
R1547 VN.n8 VN.t9 62.1016
R1548 VN.n42 VN.t6 62.1016
R1549 VN.n30 VN.n1 56.4773
R1550 VN.n64 VN.n35 56.4773
R1551 VN.n12 VN.n5 48.6874
R1552 VN.n19 VN.n3 48.6874
R1553 VN.n46 VN.n39 48.6874
R1554 VN.n53 VN.n37 48.6874
R1555 VN VN.n67 43.0701
R1556 VN.n12 VN.n11 32.1338
R1557 VN.n23 VN.n3 32.1338
R1558 VN.n46 VN.n45 32.1338
R1559 VN.n57 VN.n37 32.1338
R1560 VN.n7 VN.t3 31.8125
R1561 VN.n17 VN.t2 31.8125
R1562 VN.n25 VN.t7 31.8125
R1563 VN.n32 VN.t8 31.8125
R1564 VN.n41 VN.t1 31.8125
R1565 VN.n51 VN.t5 31.8125
R1566 VN.n59 VN.t0 31.8125
R1567 VN.n66 VN.t4 31.8125
R1568 VN.n11 VN.n10 24.3439
R1569 VN.n16 VN.n5 24.3439
R1570 VN.n19 VN.n18 24.3439
R1571 VN.n24 VN.n23 24.3439
R1572 VN.n26 VN.n1 24.3439
R1573 VN.n31 VN.n30 24.3439
R1574 VN.n45 VN.n44 24.3439
R1575 VN.n53 VN.n52 24.3439
R1576 VN.n50 VN.n39 24.3439
R1577 VN.n60 VN.n35 24.3439
R1578 VN.n58 VN.n57 24.3439
R1579 VN.n65 VN.n64 24.3439
R1580 VN.n26 VN.n25 20.449
R1581 VN.n60 VN.n59 20.449
R1582 VN.n32 VN.n31 19.9621
R1583 VN.n66 VN.n65 19.9621
R1584 VN.n43 VN.n42 13.3187
R1585 VN.n9 VN.n8 13.3187
R1586 VN.n17 VN.n16 12.1722
R1587 VN.n18 VN.n17 12.1722
R1588 VN.n52 VN.n51 12.1722
R1589 VN.n51 VN.n50 12.1722
R1590 VN.n10 VN.n7 3.89545
R1591 VN.n25 VN.n24 3.89545
R1592 VN.n44 VN.n41 3.89545
R1593 VN.n59 VN.n58 3.89545
R1594 VN.n67 VN.n34 0.278398
R1595 VN.n33 VN.n0 0.278398
R1596 VN.n63 VN.n34 0.189894
R1597 VN.n63 VN.n62 0.189894
R1598 VN.n62 VN.n61 0.189894
R1599 VN.n61 VN.n36 0.189894
R1600 VN.n56 VN.n36 0.189894
R1601 VN.n56 VN.n55 0.189894
R1602 VN.n55 VN.n54 0.189894
R1603 VN.n54 VN.n38 0.189894
R1604 VN.n49 VN.n38 0.189894
R1605 VN.n49 VN.n48 0.189894
R1606 VN.n48 VN.n47 0.189894
R1607 VN.n47 VN.n40 0.189894
R1608 VN.n43 VN.n40 0.189894
R1609 VN.n9 VN.n6 0.189894
R1610 VN.n13 VN.n6 0.189894
R1611 VN.n14 VN.n13 0.189894
R1612 VN.n15 VN.n14 0.189894
R1613 VN.n15 VN.n4 0.189894
R1614 VN.n20 VN.n4 0.189894
R1615 VN.n21 VN.n20 0.189894
R1616 VN.n22 VN.n21 0.189894
R1617 VN.n22 VN.n2 0.189894
R1618 VN.n27 VN.n2 0.189894
R1619 VN.n28 VN.n27 0.189894
R1620 VN.n29 VN.n28 0.189894
R1621 VN.n29 VN.n0 0.189894
R1622 VN VN.n33 0.153422
R1623 VDD2.n21 VDD2.n15 289.615
R1624 VDD2.n6 VDD2.n0 289.615
R1625 VDD2.n22 VDD2.n21 185
R1626 VDD2.n20 VDD2.n19 185
R1627 VDD2.n5 VDD2.n4 185
R1628 VDD2.n7 VDD2.n6 185
R1629 VDD2.n3 VDD2.t0 153.582
R1630 VDD2.n18 VDD2.t5 153.582
R1631 VDD2.n21 VDD2.n20 104.615
R1632 VDD2.n6 VDD2.n5 104.615
R1633 VDD2.n14 VDD2.n13 85.542
R1634 VDD2 VDD2.n29 85.5391
R1635 VDD2.n12 VDD2.n11 84.0909
R1636 VDD2.n28 VDD2.n27 84.0909
R1637 VDD2.n20 VDD2.t5 52.3082
R1638 VDD2.n5 VDD2.t0 52.3082
R1639 VDD2.n12 VDD2.n10 48.5455
R1640 VDD2.n26 VDD2.n25 46.5369
R1641 VDD2.n26 VDD2.n14 35.5321
R1642 VDD2.n19 VDD2.n18 10.1164
R1643 VDD2.n4 VDD2.n3 10.1164
R1644 VDD2.n25 VDD2.n24 9.45567
R1645 VDD2.n10 VDD2.n9 9.45567
R1646 VDD2.n24 VDD2.n23 9.3005
R1647 VDD2.n17 VDD2.n16 9.3005
R1648 VDD2.n2 VDD2.n1 9.3005
R1649 VDD2.n9 VDD2.n8 9.3005
R1650 VDD2.n25 VDD2.n15 8.92171
R1651 VDD2.n10 VDD2.n0 8.92171
R1652 VDD2.n23 VDD2.n22 8.14595
R1653 VDD2.n8 VDD2.n7 8.14595
R1654 VDD2.n29 VDD2.t8 7.5005
R1655 VDD2.n29 VDD2.t3 7.5005
R1656 VDD2.n27 VDD2.t9 7.5005
R1657 VDD2.n27 VDD2.t4 7.5005
R1658 VDD2.n13 VDD2.t2 7.5005
R1659 VDD2.n13 VDD2.t1 7.5005
R1660 VDD2.n11 VDD2.t6 7.5005
R1661 VDD2.n11 VDD2.t7 7.5005
R1662 VDD2.n19 VDD2.n17 7.3702
R1663 VDD2.n4 VDD2.n2 7.3702
R1664 VDD2.n22 VDD2.n17 5.81868
R1665 VDD2.n7 VDD2.n2 5.81868
R1666 VDD2.n23 VDD2.n15 5.04292
R1667 VDD2.n8 VDD2.n0 5.04292
R1668 VDD2.n18 VDD2.n16 3.00987
R1669 VDD2.n3 VDD2.n1 3.00987
R1670 VDD2.n28 VDD2.n26 2.00912
R1671 VDD2 VDD2.n28 0.560845
R1672 VDD2.n14 VDD2.n12 0.447309
R1673 VDD2.n24 VDD2.n16 0.155672
R1674 VDD2.n9 VDD2.n1 0.155672
C0 VN VDD2 2.60093f
C1 VDD1 VN 0.157249f
C2 VDD1 VDD2 1.78268f
C3 VN VP 5.79487f
C4 VP VDD2 0.512349f
C5 VN VTAIL 3.62168f
C6 VDD1 VP 2.95296f
C7 VDD2 VTAIL 5.551f
C8 VDD1 VTAIL 5.50209f
C9 VP VTAIL 3.63584f
C10 VDD2 B 4.827616f
C11 VDD1 B 4.804292f
C12 VTAIL B 3.669198f
C13 VN B 14.440939f
C14 VP B 12.925384f
C15 VDD2.n0 B 0.033354f
C16 VDD2.n1 B 0.198977f
C17 VDD2.n2 B 0.012511f
C18 VDD2.t0 B 0.053437f
C19 VDD2.n3 B 0.08648f
C20 VDD2.n4 B 0.020247f
C21 VDD2.n5 B 0.022179f
C22 VDD2.n6 B 0.065129f
C23 VDD2.n7 B 0.013247f
C24 VDD2.n8 B 0.012511f
C25 VDD2.n9 B 0.05f
C26 VDD2.n10 B 0.060544f
C27 VDD2.t6 B 0.048572f
C28 VDD2.t7 B 0.048572f
C29 VDD2.n11 B 0.338218f
C30 VDD2.n12 B 0.553957f
C31 VDD2.t2 B 0.048572f
C32 VDD2.t1 B 0.048572f
C33 VDD2.n13 B 0.345895f
C34 VDD2.n14 B 1.88645f
C35 VDD2.n15 B 0.033354f
C36 VDD2.n16 B 0.198977f
C37 VDD2.n17 B 0.012511f
C38 VDD2.t5 B 0.053437f
C39 VDD2.n18 B 0.08648f
C40 VDD2.n19 B 0.020247f
C41 VDD2.n20 B 0.022179f
C42 VDD2.n21 B 0.065129f
C43 VDD2.n22 B 0.013247f
C44 VDD2.n23 B 0.012511f
C45 VDD2.n24 B 0.05f
C46 VDD2.n25 B 0.052544f
C47 VDD2.n26 B 1.78269f
C48 VDD2.t9 B 0.048572f
C49 VDD2.t4 B 0.048572f
C50 VDD2.n27 B 0.33822f
C51 VDD2.n28 B 0.375926f
C52 VDD2.t8 B 0.048572f
C53 VDD2.t3 B 0.048572f
C54 VDD2.n29 B 0.345871f
C55 VN.n0 B 0.040988f
C56 VN.t8 B 0.401923f
C57 VN.n1 B 0.045143f
C58 VN.n2 B 0.031088f
C59 VN.t7 B 0.401923f
C60 VN.n3 B 0.02819f
C61 VN.n4 B 0.031088f
C62 VN.t2 B 0.401923f
C63 VN.n5 B 0.05823f
C64 VN.n6 B 0.031088f
C65 VN.t3 B 0.401923f
C66 VN.n7 B 0.247794f
C67 VN.t9 B 0.565404f
C68 VN.n8 B 0.253012f
C69 VN.n9 B 0.232757f
C70 VN.n10 B 0.03408f
C71 VN.n11 B 0.062969f
C72 VN.n12 B 0.02819f
C73 VN.n13 B 0.031088f
C74 VN.n14 B 0.031088f
C75 VN.n15 B 0.031088f
C76 VN.n16 B 0.043855f
C77 VN.n17 B 0.182085f
C78 VN.n18 B 0.043855f
C79 VN.n19 B 0.05823f
C80 VN.n20 B 0.031088f
C81 VN.n21 B 0.031088f
C82 VN.n22 B 0.031088f
C83 VN.n23 B 0.062969f
C84 VN.n24 B 0.03408f
C85 VN.n25 B 0.182085f
C86 VN.n26 B 0.05363f
C87 VN.n27 B 0.031088f
C88 VN.n28 B 0.031088f
C89 VN.n29 B 0.031088f
C90 VN.n30 B 0.046016f
C91 VN.n31 B 0.053055f
C92 VN.n32 B 0.278427f
C93 VN.n33 B 0.037497f
C94 VN.n34 B 0.040988f
C95 VN.t4 B 0.401923f
C96 VN.n35 B 0.045143f
C97 VN.n36 B 0.031088f
C98 VN.t0 B 0.401923f
C99 VN.n37 B 0.02819f
C100 VN.n38 B 0.031088f
C101 VN.t5 B 0.401923f
C102 VN.n39 B 0.05823f
C103 VN.n40 B 0.031088f
C104 VN.t1 B 0.401923f
C105 VN.n41 B 0.247794f
C106 VN.t6 B 0.565404f
C107 VN.n42 B 0.253012f
C108 VN.n43 B 0.232757f
C109 VN.n44 B 0.03408f
C110 VN.n45 B 0.062969f
C111 VN.n46 B 0.02819f
C112 VN.n47 B 0.031088f
C113 VN.n48 B 0.031088f
C114 VN.n49 B 0.031088f
C115 VN.n50 B 0.043855f
C116 VN.n51 B 0.182085f
C117 VN.n52 B 0.043855f
C118 VN.n53 B 0.05823f
C119 VN.n54 B 0.031088f
C120 VN.n55 B 0.031088f
C121 VN.n56 B 0.031088f
C122 VN.n57 B 0.062969f
C123 VN.n58 B 0.03408f
C124 VN.n59 B 0.182085f
C125 VN.n60 B 0.05363f
C126 VN.n61 B 0.031088f
C127 VN.n62 B 0.031088f
C128 VN.n63 B 0.031088f
C129 VN.n64 B 0.046016f
C130 VN.n65 B 0.053055f
C131 VN.n66 B 0.278427f
C132 VN.n67 B 1.3665f
C133 VDD1.n0 B 0.034216f
C134 VDD1.n1 B 0.204116f
C135 VDD1.n2 B 0.012834f
C136 VDD1.t5 B 0.054817f
C137 VDD1.n3 B 0.088714f
C138 VDD1.n4 B 0.02077f
C139 VDD1.n5 B 0.022751f
C140 VDD1.n6 B 0.066811f
C141 VDD1.n7 B 0.013589f
C142 VDD1.n8 B 0.012834f
C143 VDD1.n9 B 0.051291f
C144 VDD1.n10 B 0.062108f
C145 VDD1.t1 B 0.049827f
C146 VDD1.t8 B 0.049827f
C147 VDD1.n11 B 0.346955f
C148 VDD1.n12 B 0.575761f
C149 VDD1.n13 B 0.034216f
C150 VDD1.n14 B 0.204116f
C151 VDD1.n15 B 0.012834f
C152 VDD1.t4 B 0.054817f
C153 VDD1.n16 B 0.088714f
C154 VDD1.n17 B 0.02077f
C155 VDD1.n18 B 0.022751f
C156 VDD1.n19 B 0.066811f
C157 VDD1.n20 B 0.013589f
C158 VDD1.n21 B 0.012834f
C159 VDD1.n22 B 0.051291f
C160 VDD1.n23 B 0.062108f
C161 VDD1.t0 B 0.049827f
C162 VDD1.t7 B 0.049827f
C163 VDD1.n24 B 0.346954f
C164 VDD1.n25 B 0.568264f
C165 VDD1.t6 B 0.049827f
C166 VDD1.t2 B 0.049827f
C167 VDD1.n26 B 0.354828f
C168 VDD1.n27 B 2.03227f
C169 VDD1.t3 B 0.049827f
C170 VDD1.t9 B 0.049827f
C171 VDD1.n28 B 0.346955f
C172 VDD1.n29 B 2.08511f
C173 VTAIL.t2 B 0.068959f
C174 VTAIL.t8 B 0.068959f
C175 VTAIL.n0 B 0.417381f
C176 VTAIL.n1 B 0.601618f
C177 VTAIL.n2 B 0.047353f
C178 VTAIL.n3 B 0.282491f
C179 VTAIL.n4 B 0.017762f
C180 VTAIL.t15 B 0.075865f
C181 VTAIL.n5 B 0.122777f
C182 VTAIL.n6 B 0.028746f
C183 VTAIL.n7 B 0.031487f
C184 VTAIL.n8 B 0.092464f
C185 VTAIL.n9 B 0.018807f
C186 VTAIL.n10 B 0.017762f
C187 VTAIL.n11 B 0.070986f
C188 VTAIL.n12 B 0.051727f
C189 VTAIL.n13 B 0.396127f
C190 VTAIL.t14 B 0.068959f
C191 VTAIL.t18 B 0.068959f
C192 VTAIL.n14 B 0.417381f
C193 VTAIL.n15 B 0.705832f
C194 VTAIL.t12 B 0.068959f
C195 VTAIL.t11 B 0.068959f
C196 VTAIL.n16 B 0.417381f
C197 VTAIL.n17 B 1.61118f
C198 VTAIL.t6 B 0.068959f
C199 VTAIL.t9 B 0.068959f
C200 VTAIL.n18 B 0.417383f
C201 VTAIL.n19 B 1.61118f
C202 VTAIL.t0 B 0.068959f
C203 VTAIL.t1 B 0.068959f
C204 VTAIL.n20 B 0.417383f
C205 VTAIL.n21 B 0.70583f
C206 VTAIL.n22 B 0.047353f
C207 VTAIL.n23 B 0.282491f
C208 VTAIL.n24 B 0.017762f
C209 VTAIL.t3 B 0.075865f
C210 VTAIL.n25 B 0.122777f
C211 VTAIL.n26 B 0.028746f
C212 VTAIL.n27 B 0.031487f
C213 VTAIL.n28 B 0.092464f
C214 VTAIL.n29 B 0.018807f
C215 VTAIL.n30 B 0.017762f
C216 VTAIL.n31 B 0.070986f
C217 VTAIL.n32 B 0.051727f
C218 VTAIL.n33 B 0.396127f
C219 VTAIL.t19 B 0.068959f
C220 VTAIL.t16 B 0.068959f
C221 VTAIL.n34 B 0.417383f
C222 VTAIL.n35 B 0.648902f
C223 VTAIL.t10 B 0.068959f
C224 VTAIL.t17 B 0.068959f
C225 VTAIL.n36 B 0.417383f
C226 VTAIL.n37 B 0.70583f
C227 VTAIL.n38 B 0.047353f
C228 VTAIL.n39 B 0.282491f
C229 VTAIL.n40 B 0.017762f
C230 VTAIL.t13 B 0.075865f
C231 VTAIL.n41 B 0.122777f
C232 VTAIL.n42 B 0.028746f
C233 VTAIL.n43 B 0.031487f
C234 VTAIL.n44 B 0.092464f
C235 VTAIL.n45 B 0.018807f
C236 VTAIL.n46 B 0.017762f
C237 VTAIL.n47 B 0.070986f
C238 VTAIL.n48 B 0.051727f
C239 VTAIL.n49 B 1.14447f
C240 VTAIL.n50 B 0.047353f
C241 VTAIL.n51 B 0.282491f
C242 VTAIL.n52 B 0.017762f
C243 VTAIL.t5 B 0.075865f
C244 VTAIL.n53 B 0.122777f
C245 VTAIL.n54 B 0.028746f
C246 VTAIL.n55 B 0.031487f
C247 VTAIL.n56 B 0.092464f
C248 VTAIL.n57 B 0.018807f
C249 VTAIL.n58 B 0.017762f
C250 VTAIL.n59 B 0.070986f
C251 VTAIL.n60 B 0.051727f
C252 VTAIL.n61 B 1.14447f
C253 VTAIL.t4 B 0.068959f
C254 VTAIL.t7 B 0.068959f
C255 VTAIL.n62 B 0.417381f
C256 VTAIL.n63 B 0.539181f
C257 VP.n0 B 0.042509f
C258 VP.t7 B 0.416838f
C259 VP.n1 B 0.046819f
C260 VP.n2 B 0.032241f
C261 VP.t3 B 0.416838f
C262 VP.n3 B 0.029236f
C263 VP.n4 B 0.032241f
C264 VP.t2 B 0.416838f
C265 VP.n5 B 0.060391f
C266 VP.n6 B 0.032241f
C267 VP.t9 B 0.416838f
C268 VP.n7 B 0.188842f
C269 VP.n8 B 0.032241f
C270 VP.n9 B 0.055024f
C271 VP.n10 B 0.042509f
C272 VP.t0 B 0.416838f
C273 VP.n11 B 0.046819f
C274 VP.n12 B 0.032241f
C275 VP.t6 B 0.416838f
C276 VP.n13 B 0.029236f
C277 VP.n14 B 0.032241f
C278 VP.t1 B 0.416838f
C279 VP.n15 B 0.060391f
C280 VP.n16 B 0.032241f
C281 VP.t8 B 0.416838f
C282 VP.n17 B 0.25699f
C283 VP.t4 B 0.586386f
C284 VP.n18 B 0.262401f
C285 VP.n19 B 0.241395f
C286 VP.n20 B 0.035344f
C287 VP.n21 B 0.065306f
C288 VP.n22 B 0.029236f
C289 VP.n23 B 0.032241f
C290 VP.n24 B 0.032241f
C291 VP.n25 B 0.032241f
C292 VP.n26 B 0.045482f
C293 VP.n27 B 0.188842f
C294 VP.n28 B 0.045482f
C295 VP.n29 B 0.060391f
C296 VP.n30 B 0.032241f
C297 VP.n31 B 0.032241f
C298 VP.n32 B 0.032241f
C299 VP.n33 B 0.065306f
C300 VP.n34 B 0.035344f
C301 VP.n35 B 0.188842f
C302 VP.n36 B 0.05562f
C303 VP.n37 B 0.032241f
C304 VP.n38 B 0.032241f
C305 VP.n39 B 0.032241f
C306 VP.n40 B 0.047724f
C307 VP.n41 B 0.055024f
C308 VP.n42 B 0.28876f
C309 VP.n43 B 1.39942f
C310 VP.t5 B 0.416838f
C311 VP.n44 B 0.28876f
C312 VP.n45 B 1.42643f
C313 VP.n46 B 0.042509f
C314 VP.n47 B 0.032241f
C315 VP.n48 B 0.047724f
C316 VP.n49 B 0.046819f
C317 VP.n50 B 0.05562f
C318 VP.n51 B 0.032241f
C319 VP.n52 B 0.032241f
C320 VP.n53 B 0.035344f
C321 VP.n54 B 0.065306f
C322 VP.n55 B 0.029236f
C323 VP.n56 B 0.032241f
C324 VP.n57 B 0.032241f
C325 VP.n58 B 0.032241f
C326 VP.n59 B 0.045482f
C327 VP.n60 B 0.188842f
C328 VP.n61 B 0.045482f
C329 VP.n62 B 0.060391f
C330 VP.n63 B 0.032241f
C331 VP.n64 B 0.032241f
C332 VP.n65 B 0.032241f
C333 VP.n66 B 0.065306f
C334 VP.n67 B 0.035344f
C335 VP.n68 B 0.188842f
C336 VP.n69 B 0.05562f
C337 VP.n70 B 0.032241f
C338 VP.n71 B 0.032241f
C339 VP.n72 B 0.032241f
C340 VP.n73 B 0.047724f
C341 VP.n74 B 0.055024f
C342 VP.n75 B 0.28876f
C343 VP.n76 B 0.038888f
.ends

