* NGSPICE file created from diff_pair_sample_1509.ext - technology: sky130A

.subckt diff_pair_sample_1509 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t1 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=2.32
X1 B.t11 B.t9 B.t10 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=2.32
X2 VTAIL.t10 VN.t1 VDD2.t0 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=2.32
X3 B.t8 B.t6 B.t7 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=2.32
X4 VTAIL.t5 VP.t0 VDD1.t5 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=2.32
X5 VDD2.t5 VN.t2 VTAIL.t9 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=2.32
X6 VDD2.t3 VN.t3 VTAIL.t8 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=2.32
X7 VDD1.t4 VP.t1 VTAIL.t2 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=2.32
X8 VDD2.t2 VN.t4 VTAIL.t7 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=2.32
X9 VTAIL.t1 VP.t2 VDD1.t3 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=3.08385 ps=19.02 w=18.69 l=2.32
X10 B.t5 B.t3 B.t4 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=2.32
X11 VDD1.t2 VP.t3 VTAIL.t3 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=3.08385 ps=19.02 w=18.69 l=2.32
X12 VDD1.t1 VP.t4 VTAIL.t0 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=2.32
X13 B.t2 B.t0 B.t1 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=7.2891 pd=38.16 as=0 ps=0 w=18.69 l=2.32
X14 VDD2.t4 VN.t5 VTAIL.t6 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=2.32
X15 VDD1.t0 VP.t5 VTAIL.t4 w_n3090_n4706# sky130_fd_pr__pfet_01v8 ad=3.08385 pd=19.02 as=7.2891 ps=38.16 w=18.69 l=2.32
R0 VN.n3 VN.t2 226.968
R1 VN.n17 VN.t4 226.968
R2 VN.n4 VN.t0 194.15
R3 VN.n12 VN.t5 194.15
R4 VN.n18 VN.t1 194.15
R5 VN.n26 VN.t3 194.15
R6 VN.n25 VN.n14 161.3
R7 VN.n24 VN.n23 161.3
R8 VN.n22 VN.n15 161.3
R9 VN.n21 VN.n20 161.3
R10 VN.n19 VN.n16 161.3
R11 VN.n11 VN.n0 161.3
R12 VN.n10 VN.n9 161.3
R13 VN.n8 VN.n1 161.3
R14 VN.n7 VN.n6 161.3
R15 VN.n5 VN.n2 161.3
R16 VN.n13 VN.n12 103.416
R17 VN.n27 VN.n26 103.416
R18 VN.n6 VN.n1 56.5193
R19 VN.n20 VN.n15 56.5193
R20 VN VN.n27 52.8353
R21 VN.n4 VN.n3 47.8187
R22 VN.n18 VN.n17 47.8187
R23 VN.n5 VN.n4 24.4675
R24 VN.n6 VN.n5 24.4675
R25 VN.n10 VN.n1 24.4675
R26 VN.n11 VN.n10 24.4675
R27 VN.n20 VN.n19 24.4675
R28 VN.n19 VN.n18 24.4675
R29 VN.n25 VN.n24 24.4675
R30 VN.n24 VN.n15 24.4675
R31 VN.n12 VN.n11 7.3406
R32 VN.n26 VN.n25 7.3406
R33 VN.n17 VN.n16 7.01727
R34 VN.n3 VN.n2 7.01727
R35 VN.n27 VN.n14 0.278367
R36 VN.n13 VN.n0 0.278367
R37 VN.n23 VN.n14 0.189894
R38 VN.n23 VN.n22 0.189894
R39 VN.n22 VN.n21 0.189894
R40 VN.n21 VN.n16 0.189894
R41 VN.n7 VN.n2 0.189894
R42 VN.n8 VN.n7 0.189894
R43 VN.n9 VN.n8 0.189894
R44 VN.n9 VN.n0 0.189894
R45 VN VN.n13 0.153454
R46 VDD2.n1 VDD2.t5 73.675
R47 VDD2.n2 VDD2.t3 72.0171
R48 VDD2.n1 VDD2.n0 70.7935
R49 VDD2 VDD2.n3 70.7907
R50 VDD2.n2 VDD2.n1 47.2519
R51 VDD2 VDD2.n2 1.77205
R52 VDD2.n3 VDD2.t0 1.73967
R53 VDD2.n3 VDD2.t2 1.73967
R54 VDD2.n0 VDD2.t1 1.73967
R55 VDD2.n0 VDD2.t4 1.73967
R56 VTAIL.n7 VTAIL.t7 55.3383
R57 VTAIL.n11 VTAIL.t6 55.3382
R58 VTAIL.n2 VTAIL.t0 55.3382
R59 VTAIL.n10 VTAIL.t4 55.3382
R60 VTAIL.n9 VTAIL.n8 53.5992
R61 VTAIL.n6 VTAIL.n5 53.5992
R62 VTAIL.n1 VTAIL.n0 53.599
R63 VTAIL.n4 VTAIL.n3 53.599
R64 VTAIL.n6 VTAIL.n4 33.0479
R65 VTAIL.n11 VTAIL.n10 30.7634
R66 VTAIL.n7 VTAIL.n6 2.28498
R67 VTAIL.n10 VTAIL.n9 2.28498
R68 VTAIL.n4 VTAIL.n2 2.28498
R69 VTAIL.n0 VTAIL.t9 1.73967
R70 VTAIL.n0 VTAIL.t11 1.73967
R71 VTAIL.n3 VTAIL.t2 1.73967
R72 VTAIL.n3 VTAIL.t1 1.73967
R73 VTAIL.n8 VTAIL.t3 1.73967
R74 VTAIL.n8 VTAIL.t5 1.73967
R75 VTAIL.n5 VTAIL.t8 1.73967
R76 VTAIL.n5 VTAIL.t10 1.73967
R77 VTAIL VTAIL.n11 1.65567
R78 VTAIL.n9 VTAIL.n7 1.61257
R79 VTAIL.n2 VTAIL.n1 1.61257
R80 VTAIL VTAIL.n1 0.62981
R81 B.n597 B.n596 585
R82 B.n598 B.n91 585
R83 B.n600 B.n599 585
R84 B.n601 B.n90 585
R85 B.n603 B.n602 585
R86 B.n604 B.n89 585
R87 B.n606 B.n605 585
R88 B.n607 B.n88 585
R89 B.n609 B.n608 585
R90 B.n610 B.n87 585
R91 B.n612 B.n611 585
R92 B.n613 B.n86 585
R93 B.n615 B.n614 585
R94 B.n616 B.n85 585
R95 B.n618 B.n617 585
R96 B.n619 B.n84 585
R97 B.n621 B.n620 585
R98 B.n622 B.n83 585
R99 B.n624 B.n623 585
R100 B.n625 B.n82 585
R101 B.n627 B.n626 585
R102 B.n628 B.n81 585
R103 B.n630 B.n629 585
R104 B.n631 B.n80 585
R105 B.n633 B.n632 585
R106 B.n634 B.n79 585
R107 B.n636 B.n635 585
R108 B.n637 B.n78 585
R109 B.n639 B.n638 585
R110 B.n640 B.n77 585
R111 B.n642 B.n641 585
R112 B.n643 B.n76 585
R113 B.n645 B.n644 585
R114 B.n646 B.n75 585
R115 B.n648 B.n647 585
R116 B.n649 B.n74 585
R117 B.n651 B.n650 585
R118 B.n652 B.n73 585
R119 B.n654 B.n653 585
R120 B.n655 B.n72 585
R121 B.n657 B.n656 585
R122 B.n658 B.n71 585
R123 B.n660 B.n659 585
R124 B.n661 B.n70 585
R125 B.n663 B.n662 585
R126 B.n664 B.n69 585
R127 B.n666 B.n665 585
R128 B.n667 B.n68 585
R129 B.n669 B.n668 585
R130 B.n670 B.n67 585
R131 B.n672 B.n671 585
R132 B.n673 B.n66 585
R133 B.n675 B.n674 585
R134 B.n676 B.n65 585
R135 B.n678 B.n677 585
R136 B.n679 B.n64 585
R137 B.n681 B.n680 585
R138 B.n682 B.n63 585
R139 B.n684 B.n683 585
R140 B.n685 B.n62 585
R141 B.n687 B.n686 585
R142 B.n689 B.n59 585
R143 B.n691 B.n690 585
R144 B.n692 B.n58 585
R145 B.n694 B.n693 585
R146 B.n695 B.n57 585
R147 B.n697 B.n696 585
R148 B.n698 B.n56 585
R149 B.n700 B.n699 585
R150 B.n701 B.n55 585
R151 B.n703 B.n702 585
R152 B.n705 B.n704 585
R153 B.n706 B.n51 585
R154 B.n708 B.n707 585
R155 B.n709 B.n50 585
R156 B.n711 B.n710 585
R157 B.n712 B.n49 585
R158 B.n714 B.n713 585
R159 B.n715 B.n48 585
R160 B.n717 B.n716 585
R161 B.n718 B.n47 585
R162 B.n720 B.n719 585
R163 B.n721 B.n46 585
R164 B.n723 B.n722 585
R165 B.n724 B.n45 585
R166 B.n726 B.n725 585
R167 B.n727 B.n44 585
R168 B.n729 B.n728 585
R169 B.n730 B.n43 585
R170 B.n732 B.n731 585
R171 B.n733 B.n42 585
R172 B.n735 B.n734 585
R173 B.n736 B.n41 585
R174 B.n738 B.n737 585
R175 B.n739 B.n40 585
R176 B.n741 B.n740 585
R177 B.n742 B.n39 585
R178 B.n744 B.n743 585
R179 B.n745 B.n38 585
R180 B.n747 B.n746 585
R181 B.n748 B.n37 585
R182 B.n750 B.n749 585
R183 B.n751 B.n36 585
R184 B.n753 B.n752 585
R185 B.n754 B.n35 585
R186 B.n756 B.n755 585
R187 B.n757 B.n34 585
R188 B.n759 B.n758 585
R189 B.n760 B.n33 585
R190 B.n762 B.n761 585
R191 B.n763 B.n32 585
R192 B.n765 B.n764 585
R193 B.n766 B.n31 585
R194 B.n768 B.n767 585
R195 B.n769 B.n30 585
R196 B.n771 B.n770 585
R197 B.n772 B.n29 585
R198 B.n774 B.n773 585
R199 B.n775 B.n28 585
R200 B.n777 B.n776 585
R201 B.n778 B.n27 585
R202 B.n780 B.n779 585
R203 B.n781 B.n26 585
R204 B.n783 B.n782 585
R205 B.n784 B.n25 585
R206 B.n786 B.n785 585
R207 B.n787 B.n24 585
R208 B.n789 B.n788 585
R209 B.n790 B.n23 585
R210 B.n792 B.n791 585
R211 B.n793 B.n22 585
R212 B.n795 B.n794 585
R213 B.n595 B.n92 585
R214 B.n594 B.n593 585
R215 B.n592 B.n93 585
R216 B.n591 B.n590 585
R217 B.n589 B.n94 585
R218 B.n588 B.n587 585
R219 B.n586 B.n95 585
R220 B.n585 B.n584 585
R221 B.n583 B.n96 585
R222 B.n582 B.n581 585
R223 B.n580 B.n97 585
R224 B.n579 B.n578 585
R225 B.n577 B.n98 585
R226 B.n576 B.n575 585
R227 B.n574 B.n99 585
R228 B.n573 B.n572 585
R229 B.n571 B.n100 585
R230 B.n570 B.n569 585
R231 B.n568 B.n101 585
R232 B.n567 B.n566 585
R233 B.n565 B.n102 585
R234 B.n564 B.n563 585
R235 B.n562 B.n103 585
R236 B.n561 B.n560 585
R237 B.n559 B.n104 585
R238 B.n558 B.n557 585
R239 B.n556 B.n105 585
R240 B.n555 B.n554 585
R241 B.n553 B.n106 585
R242 B.n552 B.n551 585
R243 B.n550 B.n107 585
R244 B.n549 B.n548 585
R245 B.n547 B.n108 585
R246 B.n546 B.n545 585
R247 B.n544 B.n109 585
R248 B.n543 B.n542 585
R249 B.n541 B.n110 585
R250 B.n540 B.n539 585
R251 B.n538 B.n111 585
R252 B.n537 B.n536 585
R253 B.n535 B.n112 585
R254 B.n534 B.n533 585
R255 B.n532 B.n113 585
R256 B.n531 B.n530 585
R257 B.n529 B.n114 585
R258 B.n528 B.n527 585
R259 B.n526 B.n115 585
R260 B.n525 B.n524 585
R261 B.n523 B.n116 585
R262 B.n522 B.n521 585
R263 B.n520 B.n117 585
R264 B.n519 B.n518 585
R265 B.n517 B.n118 585
R266 B.n516 B.n515 585
R267 B.n514 B.n119 585
R268 B.n513 B.n512 585
R269 B.n511 B.n120 585
R270 B.n510 B.n509 585
R271 B.n508 B.n121 585
R272 B.n507 B.n506 585
R273 B.n505 B.n122 585
R274 B.n504 B.n503 585
R275 B.n502 B.n123 585
R276 B.n501 B.n500 585
R277 B.n499 B.n124 585
R278 B.n498 B.n497 585
R279 B.n496 B.n125 585
R280 B.n495 B.n494 585
R281 B.n493 B.n126 585
R282 B.n492 B.n491 585
R283 B.n490 B.n127 585
R284 B.n489 B.n488 585
R285 B.n487 B.n128 585
R286 B.n486 B.n485 585
R287 B.n484 B.n129 585
R288 B.n483 B.n482 585
R289 B.n481 B.n130 585
R290 B.n480 B.n479 585
R291 B.n478 B.n131 585
R292 B.n279 B.n278 585
R293 B.n280 B.n201 585
R294 B.n282 B.n281 585
R295 B.n283 B.n200 585
R296 B.n285 B.n284 585
R297 B.n286 B.n199 585
R298 B.n288 B.n287 585
R299 B.n289 B.n198 585
R300 B.n291 B.n290 585
R301 B.n292 B.n197 585
R302 B.n294 B.n293 585
R303 B.n295 B.n196 585
R304 B.n297 B.n296 585
R305 B.n298 B.n195 585
R306 B.n300 B.n299 585
R307 B.n301 B.n194 585
R308 B.n303 B.n302 585
R309 B.n304 B.n193 585
R310 B.n306 B.n305 585
R311 B.n307 B.n192 585
R312 B.n309 B.n308 585
R313 B.n310 B.n191 585
R314 B.n312 B.n311 585
R315 B.n313 B.n190 585
R316 B.n315 B.n314 585
R317 B.n316 B.n189 585
R318 B.n318 B.n317 585
R319 B.n319 B.n188 585
R320 B.n321 B.n320 585
R321 B.n322 B.n187 585
R322 B.n324 B.n323 585
R323 B.n325 B.n186 585
R324 B.n327 B.n326 585
R325 B.n328 B.n185 585
R326 B.n330 B.n329 585
R327 B.n331 B.n184 585
R328 B.n333 B.n332 585
R329 B.n334 B.n183 585
R330 B.n336 B.n335 585
R331 B.n337 B.n182 585
R332 B.n339 B.n338 585
R333 B.n340 B.n181 585
R334 B.n342 B.n341 585
R335 B.n343 B.n180 585
R336 B.n345 B.n344 585
R337 B.n346 B.n179 585
R338 B.n348 B.n347 585
R339 B.n349 B.n178 585
R340 B.n351 B.n350 585
R341 B.n352 B.n177 585
R342 B.n354 B.n353 585
R343 B.n355 B.n176 585
R344 B.n357 B.n356 585
R345 B.n358 B.n175 585
R346 B.n360 B.n359 585
R347 B.n361 B.n174 585
R348 B.n363 B.n362 585
R349 B.n364 B.n173 585
R350 B.n366 B.n365 585
R351 B.n367 B.n172 585
R352 B.n369 B.n368 585
R353 B.n371 B.n169 585
R354 B.n373 B.n372 585
R355 B.n374 B.n168 585
R356 B.n376 B.n375 585
R357 B.n377 B.n167 585
R358 B.n379 B.n378 585
R359 B.n380 B.n166 585
R360 B.n382 B.n381 585
R361 B.n383 B.n165 585
R362 B.n385 B.n384 585
R363 B.n387 B.n386 585
R364 B.n388 B.n161 585
R365 B.n390 B.n389 585
R366 B.n391 B.n160 585
R367 B.n393 B.n392 585
R368 B.n394 B.n159 585
R369 B.n396 B.n395 585
R370 B.n397 B.n158 585
R371 B.n399 B.n398 585
R372 B.n400 B.n157 585
R373 B.n402 B.n401 585
R374 B.n403 B.n156 585
R375 B.n405 B.n404 585
R376 B.n406 B.n155 585
R377 B.n408 B.n407 585
R378 B.n409 B.n154 585
R379 B.n411 B.n410 585
R380 B.n412 B.n153 585
R381 B.n414 B.n413 585
R382 B.n415 B.n152 585
R383 B.n417 B.n416 585
R384 B.n418 B.n151 585
R385 B.n420 B.n419 585
R386 B.n421 B.n150 585
R387 B.n423 B.n422 585
R388 B.n424 B.n149 585
R389 B.n426 B.n425 585
R390 B.n427 B.n148 585
R391 B.n429 B.n428 585
R392 B.n430 B.n147 585
R393 B.n432 B.n431 585
R394 B.n433 B.n146 585
R395 B.n435 B.n434 585
R396 B.n436 B.n145 585
R397 B.n438 B.n437 585
R398 B.n439 B.n144 585
R399 B.n441 B.n440 585
R400 B.n442 B.n143 585
R401 B.n444 B.n443 585
R402 B.n445 B.n142 585
R403 B.n447 B.n446 585
R404 B.n448 B.n141 585
R405 B.n450 B.n449 585
R406 B.n451 B.n140 585
R407 B.n453 B.n452 585
R408 B.n454 B.n139 585
R409 B.n456 B.n455 585
R410 B.n457 B.n138 585
R411 B.n459 B.n458 585
R412 B.n460 B.n137 585
R413 B.n462 B.n461 585
R414 B.n463 B.n136 585
R415 B.n465 B.n464 585
R416 B.n466 B.n135 585
R417 B.n468 B.n467 585
R418 B.n469 B.n134 585
R419 B.n471 B.n470 585
R420 B.n472 B.n133 585
R421 B.n474 B.n473 585
R422 B.n475 B.n132 585
R423 B.n477 B.n476 585
R424 B.n277 B.n202 585
R425 B.n276 B.n275 585
R426 B.n274 B.n203 585
R427 B.n273 B.n272 585
R428 B.n271 B.n204 585
R429 B.n270 B.n269 585
R430 B.n268 B.n205 585
R431 B.n267 B.n266 585
R432 B.n265 B.n206 585
R433 B.n264 B.n263 585
R434 B.n262 B.n207 585
R435 B.n261 B.n260 585
R436 B.n259 B.n208 585
R437 B.n258 B.n257 585
R438 B.n256 B.n209 585
R439 B.n255 B.n254 585
R440 B.n253 B.n210 585
R441 B.n252 B.n251 585
R442 B.n250 B.n211 585
R443 B.n249 B.n248 585
R444 B.n247 B.n212 585
R445 B.n246 B.n245 585
R446 B.n244 B.n213 585
R447 B.n243 B.n242 585
R448 B.n241 B.n214 585
R449 B.n240 B.n239 585
R450 B.n238 B.n215 585
R451 B.n237 B.n236 585
R452 B.n235 B.n216 585
R453 B.n234 B.n233 585
R454 B.n232 B.n217 585
R455 B.n231 B.n230 585
R456 B.n229 B.n218 585
R457 B.n228 B.n227 585
R458 B.n226 B.n219 585
R459 B.n225 B.n224 585
R460 B.n223 B.n220 585
R461 B.n222 B.n221 585
R462 B.n2 B.n0 585
R463 B.n853 B.n1 585
R464 B.n852 B.n851 585
R465 B.n850 B.n3 585
R466 B.n849 B.n848 585
R467 B.n847 B.n4 585
R468 B.n846 B.n845 585
R469 B.n844 B.n5 585
R470 B.n843 B.n842 585
R471 B.n841 B.n6 585
R472 B.n840 B.n839 585
R473 B.n838 B.n7 585
R474 B.n837 B.n836 585
R475 B.n835 B.n8 585
R476 B.n834 B.n833 585
R477 B.n832 B.n9 585
R478 B.n831 B.n830 585
R479 B.n829 B.n10 585
R480 B.n828 B.n827 585
R481 B.n826 B.n11 585
R482 B.n825 B.n824 585
R483 B.n823 B.n12 585
R484 B.n822 B.n821 585
R485 B.n820 B.n13 585
R486 B.n819 B.n818 585
R487 B.n817 B.n14 585
R488 B.n816 B.n815 585
R489 B.n814 B.n15 585
R490 B.n813 B.n812 585
R491 B.n811 B.n16 585
R492 B.n810 B.n809 585
R493 B.n808 B.n17 585
R494 B.n807 B.n806 585
R495 B.n805 B.n18 585
R496 B.n804 B.n803 585
R497 B.n802 B.n19 585
R498 B.n801 B.n800 585
R499 B.n799 B.n20 585
R500 B.n798 B.n797 585
R501 B.n796 B.n21 585
R502 B.n855 B.n854 585
R503 B.n278 B.n277 559.769
R504 B.n794 B.n21 559.769
R505 B.n476 B.n131 559.769
R506 B.n596 B.n595 559.769
R507 B.n162 B.t9 401.731
R508 B.n170 B.t3 401.731
R509 B.n52 B.t6 401.731
R510 B.n60 B.t0 401.731
R511 B.n162 B.t11 163.933
R512 B.n60 B.t1 163.933
R513 B.n170 B.t5 163.909
R514 B.n52 B.t7 163.909
R515 B.n277 B.n276 163.367
R516 B.n276 B.n203 163.367
R517 B.n272 B.n203 163.367
R518 B.n272 B.n271 163.367
R519 B.n271 B.n270 163.367
R520 B.n270 B.n205 163.367
R521 B.n266 B.n205 163.367
R522 B.n266 B.n265 163.367
R523 B.n265 B.n264 163.367
R524 B.n264 B.n207 163.367
R525 B.n260 B.n207 163.367
R526 B.n260 B.n259 163.367
R527 B.n259 B.n258 163.367
R528 B.n258 B.n209 163.367
R529 B.n254 B.n209 163.367
R530 B.n254 B.n253 163.367
R531 B.n253 B.n252 163.367
R532 B.n252 B.n211 163.367
R533 B.n248 B.n211 163.367
R534 B.n248 B.n247 163.367
R535 B.n247 B.n246 163.367
R536 B.n246 B.n213 163.367
R537 B.n242 B.n213 163.367
R538 B.n242 B.n241 163.367
R539 B.n241 B.n240 163.367
R540 B.n240 B.n215 163.367
R541 B.n236 B.n215 163.367
R542 B.n236 B.n235 163.367
R543 B.n235 B.n234 163.367
R544 B.n234 B.n217 163.367
R545 B.n230 B.n217 163.367
R546 B.n230 B.n229 163.367
R547 B.n229 B.n228 163.367
R548 B.n228 B.n219 163.367
R549 B.n224 B.n219 163.367
R550 B.n224 B.n223 163.367
R551 B.n223 B.n222 163.367
R552 B.n222 B.n2 163.367
R553 B.n854 B.n2 163.367
R554 B.n854 B.n853 163.367
R555 B.n853 B.n852 163.367
R556 B.n852 B.n3 163.367
R557 B.n848 B.n3 163.367
R558 B.n848 B.n847 163.367
R559 B.n847 B.n846 163.367
R560 B.n846 B.n5 163.367
R561 B.n842 B.n5 163.367
R562 B.n842 B.n841 163.367
R563 B.n841 B.n840 163.367
R564 B.n840 B.n7 163.367
R565 B.n836 B.n7 163.367
R566 B.n836 B.n835 163.367
R567 B.n835 B.n834 163.367
R568 B.n834 B.n9 163.367
R569 B.n830 B.n9 163.367
R570 B.n830 B.n829 163.367
R571 B.n829 B.n828 163.367
R572 B.n828 B.n11 163.367
R573 B.n824 B.n11 163.367
R574 B.n824 B.n823 163.367
R575 B.n823 B.n822 163.367
R576 B.n822 B.n13 163.367
R577 B.n818 B.n13 163.367
R578 B.n818 B.n817 163.367
R579 B.n817 B.n816 163.367
R580 B.n816 B.n15 163.367
R581 B.n812 B.n15 163.367
R582 B.n812 B.n811 163.367
R583 B.n811 B.n810 163.367
R584 B.n810 B.n17 163.367
R585 B.n806 B.n17 163.367
R586 B.n806 B.n805 163.367
R587 B.n805 B.n804 163.367
R588 B.n804 B.n19 163.367
R589 B.n800 B.n19 163.367
R590 B.n800 B.n799 163.367
R591 B.n799 B.n798 163.367
R592 B.n798 B.n21 163.367
R593 B.n278 B.n201 163.367
R594 B.n282 B.n201 163.367
R595 B.n283 B.n282 163.367
R596 B.n284 B.n283 163.367
R597 B.n284 B.n199 163.367
R598 B.n288 B.n199 163.367
R599 B.n289 B.n288 163.367
R600 B.n290 B.n289 163.367
R601 B.n290 B.n197 163.367
R602 B.n294 B.n197 163.367
R603 B.n295 B.n294 163.367
R604 B.n296 B.n295 163.367
R605 B.n296 B.n195 163.367
R606 B.n300 B.n195 163.367
R607 B.n301 B.n300 163.367
R608 B.n302 B.n301 163.367
R609 B.n302 B.n193 163.367
R610 B.n306 B.n193 163.367
R611 B.n307 B.n306 163.367
R612 B.n308 B.n307 163.367
R613 B.n308 B.n191 163.367
R614 B.n312 B.n191 163.367
R615 B.n313 B.n312 163.367
R616 B.n314 B.n313 163.367
R617 B.n314 B.n189 163.367
R618 B.n318 B.n189 163.367
R619 B.n319 B.n318 163.367
R620 B.n320 B.n319 163.367
R621 B.n320 B.n187 163.367
R622 B.n324 B.n187 163.367
R623 B.n325 B.n324 163.367
R624 B.n326 B.n325 163.367
R625 B.n326 B.n185 163.367
R626 B.n330 B.n185 163.367
R627 B.n331 B.n330 163.367
R628 B.n332 B.n331 163.367
R629 B.n332 B.n183 163.367
R630 B.n336 B.n183 163.367
R631 B.n337 B.n336 163.367
R632 B.n338 B.n337 163.367
R633 B.n338 B.n181 163.367
R634 B.n342 B.n181 163.367
R635 B.n343 B.n342 163.367
R636 B.n344 B.n343 163.367
R637 B.n344 B.n179 163.367
R638 B.n348 B.n179 163.367
R639 B.n349 B.n348 163.367
R640 B.n350 B.n349 163.367
R641 B.n350 B.n177 163.367
R642 B.n354 B.n177 163.367
R643 B.n355 B.n354 163.367
R644 B.n356 B.n355 163.367
R645 B.n356 B.n175 163.367
R646 B.n360 B.n175 163.367
R647 B.n361 B.n360 163.367
R648 B.n362 B.n361 163.367
R649 B.n362 B.n173 163.367
R650 B.n366 B.n173 163.367
R651 B.n367 B.n366 163.367
R652 B.n368 B.n367 163.367
R653 B.n368 B.n169 163.367
R654 B.n373 B.n169 163.367
R655 B.n374 B.n373 163.367
R656 B.n375 B.n374 163.367
R657 B.n375 B.n167 163.367
R658 B.n379 B.n167 163.367
R659 B.n380 B.n379 163.367
R660 B.n381 B.n380 163.367
R661 B.n381 B.n165 163.367
R662 B.n385 B.n165 163.367
R663 B.n386 B.n385 163.367
R664 B.n386 B.n161 163.367
R665 B.n390 B.n161 163.367
R666 B.n391 B.n390 163.367
R667 B.n392 B.n391 163.367
R668 B.n392 B.n159 163.367
R669 B.n396 B.n159 163.367
R670 B.n397 B.n396 163.367
R671 B.n398 B.n397 163.367
R672 B.n398 B.n157 163.367
R673 B.n402 B.n157 163.367
R674 B.n403 B.n402 163.367
R675 B.n404 B.n403 163.367
R676 B.n404 B.n155 163.367
R677 B.n408 B.n155 163.367
R678 B.n409 B.n408 163.367
R679 B.n410 B.n409 163.367
R680 B.n410 B.n153 163.367
R681 B.n414 B.n153 163.367
R682 B.n415 B.n414 163.367
R683 B.n416 B.n415 163.367
R684 B.n416 B.n151 163.367
R685 B.n420 B.n151 163.367
R686 B.n421 B.n420 163.367
R687 B.n422 B.n421 163.367
R688 B.n422 B.n149 163.367
R689 B.n426 B.n149 163.367
R690 B.n427 B.n426 163.367
R691 B.n428 B.n427 163.367
R692 B.n428 B.n147 163.367
R693 B.n432 B.n147 163.367
R694 B.n433 B.n432 163.367
R695 B.n434 B.n433 163.367
R696 B.n434 B.n145 163.367
R697 B.n438 B.n145 163.367
R698 B.n439 B.n438 163.367
R699 B.n440 B.n439 163.367
R700 B.n440 B.n143 163.367
R701 B.n444 B.n143 163.367
R702 B.n445 B.n444 163.367
R703 B.n446 B.n445 163.367
R704 B.n446 B.n141 163.367
R705 B.n450 B.n141 163.367
R706 B.n451 B.n450 163.367
R707 B.n452 B.n451 163.367
R708 B.n452 B.n139 163.367
R709 B.n456 B.n139 163.367
R710 B.n457 B.n456 163.367
R711 B.n458 B.n457 163.367
R712 B.n458 B.n137 163.367
R713 B.n462 B.n137 163.367
R714 B.n463 B.n462 163.367
R715 B.n464 B.n463 163.367
R716 B.n464 B.n135 163.367
R717 B.n468 B.n135 163.367
R718 B.n469 B.n468 163.367
R719 B.n470 B.n469 163.367
R720 B.n470 B.n133 163.367
R721 B.n474 B.n133 163.367
R722 B.n475 B.n474 163.367
R723 B.n476 B.n475 163.367
R724 B.n480 B.n131 163.367
R725 B.n481 B.n480 163.367
R726 B.n482 B.n481 163.367
R727 B.n482 B.n129 163.367
R728 B.n486 B.n129 163.367
R729 B.n487 B.n486 163.367
R730 B.n488 B.n487 163.367
R731 B.n488 B.n127 163.367
R732 B.n492 B.n127 163.367
R733 B.n493 B.n492 163.367
R734 B.n494 B.n493 163.367
R735 B.n494 B.n125 163.367
R736 B.n498 B.n125 163.367
R737 B.n499 B.n498 163.367
R738 B.n500 B.n499 163.367
R739 B.n500 B.n123 163.367
R740 B.n504 B.n123 163.367
R741 B.n505 B.n504 163.367
R742 B.n506 B.n505 163.367
R743 B.n506 B.n121 163.367
R744 B.n510 B.n121 163.367
R745 B.n511 B.n510 163.367
R746 B.n512 B.n511 163.367
R747 B.n512 B.n119 163.367
R748 B.n516 B.n119 163.367
R749 B.n517 B.n516 163.367
R750 B.n518 B.n517 163.367
R751 B.n518 B.n117 163.367
R752 B.n522 B.n117 163.367
R753 B.n523 B.n522 163.367
R754 B.n524 B.n523 163.367
R755 B.n524 B.n115 163.367
R756 B.n528 B.n115 163.367
R757 B.n529 B.n528 163.367
R758 B.n530 B.n529 163.367
R759 B.n530 B.n113 163.367
R760 B.n534 B.n113 163.367
R761 B.n535 B.n534 163.367
R762 B.n536 B.n535 163.367
R763 B.n536 B.n111 163.367
R764 B.n540 B.n111 163.367
R765 B.n541 B.n540 163.367
R766 B.n542 B.n541 163.367
R767 B.n542 B.n109 163.367
R768 B.n546 B.n109 163.367
R769 B.n547 B.n546 163.367
R770 B.n548 B.n547 163.367
R771 B.n548 B.n107 163.367
R772 B.n552 B.n107 163.367
R773 B.n553 B.n552 163.367
R774 B.n554 B.n553 163.367
R775 B.n554 B.n105 163.367
R776 B.n558 B.n105 163.367
R777 B.n559 B.n558 163.367
R778 B.n560 B.n559 163.367
R779 B.n560 B.n103 163.367
R780 B.n564 B.n103 163.367
R781 B.n565 B.n564 163.367
R782 B.n566 B.n565 163.367
R783 B.n566 B.n101 163.367
R784 B.n570 B.n101 163.367
R785 B.n571 B.n570 163.367
R786 B.n572 B.n571 163.367
R787 B.n572 B.n99 163.367
R788 B.n576 B.n99 163.367
R789 B.n577 B.n576 163.367
R790 B.n578 B.n577 163.367
R791 B.n578 B.n97 163.367
R792 B.n582 B.n97 163.367
R793 B.n583 B.n582 163.367
R794 B.n584 B.n583 163.367
R795 B.n584 B.n95 163.367
R796 B.n588 B.n95 163.367
R797 B.n589 B.n588 163.367
R798 B.n590 B.n589 163.367
R799 B.n590 B.n93 163.367
R800 B.n594 B.n93 163.367
R801 B.n595 B.n594 163.367
R802 B.n794 B.n793 163.367
R803 B.n793 B.n792 163.367
R804 B.n792 B.n23 163.367
R805 B.n788 B.n23 163.367
R806 B.n788 B.n787 163.367
R807 B.n787 B.n786 163.367
R808 B.n786 B.n25 163.367
R809 B.n782 B.n25 163.367
R810 B.n782 B.n781 163.367
R811 B.n781 B.n780 163.367
R812 B.n780 B.n27 163.367
R813 B.n776 B.n27 163.367
R814 B.n776 B.n775 163.367
R815 B.n775 B.n774 163.367
R816 B.n774 B.n29 163.367
R817 B.n770 B.n29 163.367
R818 B.n770 B.n769 163.367
R819 B.n769 B.n768 163.367
R820 B.n768 B.n31 163.367
R821 B.n764 B.n31 163.367
R822 B.n764 B.n763 163.367
R823 B.n763 B.n762 163.367
R824 B.n762 B.n33 163.367
R825 B.n758 B.n33 163.367
R826 B.n758 B.n757 163.367
R827 B.n757 B.n756 163.367
R828 B.n756 B.n35 163.367
R829 B.n752 B.n35 163.367
R830 B.n752 B.n751 163.367
R831 B.n751 B.n750 163.367
R832 B.n750 B.n37 163.367
R833 B.n746 B.n37 163.367
R834 B.n746 B.n745 163.367
R835 B.n745 B.n744 163.367
R836 B.n744 B.n39 163.367
R837 B.n740 B.n39 163.367
R838 B.n740 B.n739 163.367
R839 B.n739 B.n738 163.367
R840 B.n738 B.n41 163.367
R841 B.n734 B.n41 163.367
R842 B.n734 B.n733 163.367
R843 B.n733 B.n732 163.367
R844 B.n732 B.n43 163.367
R845 B.n728 B.n43 163.367
R846 B.n728 B.n727 163.367
R847 B.n727 B.n726 163.367
R848 B.n726 B.n45 163.367
R849 B.n722 B.n45 163.367
R850 B.n722 B.n721 163.367
R851 B.n721 B.n720 163.367
R852 B.n720 B.n47 163.367
R853 B.n716 B.n47 163.367
R854 B.n716 B.n715 163.367
R855 B.n715 B.n714 163.367
R856 B.n714 B.n49 163.367
R857 B.n710 B.n49 163.367
R858 B.n710 B.n709 163.367
R859 B.n709 B.n708 163.367
R860 B.n708 B.n51 163.367
R861 B.n704 B.n51 163.367
R862 B.n704 B.n703 163.367
R863 B.n703 B.n55 163.367
R864 B.n699 B.n55 163.367
R865 B.n699 B.n698 163.367
R866 B.n698 B.n697 163.367
R867 B.n697 B.n57 163.367
R868 B.n693 B.n57 163.367
R869 B.n693 B.n692 163.367
R870 B.n692 B.n691 163.367
R871 B.n691 B.n59 163.367
R872 B.n686 B.n59 163.367
R873 B.n686 B.n685 163.367
R874 B.n685 B.n684 163.367
R875 B.n684 B.n63 163.367
R876 B.n680 B.n63 163.367
R877 B.n680 B.n679 163.367
R878 B.n679 B.n678 163.367
R879 B.n678 B.n65 163.367
R880 B.n674 B.n65 163.367
R881 B.n674 B.n673 163.367
R882 B.n673 B.n672 163.367
R883 B.n672 B.n67 163.367
R884 B.n668 B.n67 163.367
R885 B.n668 B.n667 163.367
R886 B.n667 B.n666 163.367
R887 B.n666 B.n69 163.367
R888 B.n662 B.n69 163.367
R889 B.n662 B.n661 163.367
R890 B.n661 B.n660 163.367
R891 B.n660 B.n71 163.367
R892 B.n656 B.n71 163.367
R893 B.n656 B.n655 163.367
R894 B.n655 B.n654 163.367
R895 B.n654 B.n73 163.367
R896 B.n650 B.n73 163.367
R897 B.n650 B.n649 163.367
R898 B.n649 B.n648 163.367
R899 B.n648 B.n75 163.367
R900 B.n644 B.n75 163.367
R901 B.n644 B.n643 163.367
R902 B.n643 B.n642 163.367
R903 B.n642 B.n77 163.367
R904 B.n638 B.n77 163.367
R905 B.n638 B.n637 163.367
R906 B.n637 B.n636 163.367
R907 B.n636 B.n79 163.367
R908 B.n632 B.n79 163.367
R909 B.n632 B.n631 163.367
R910 B.n631 B.n630 163.367
R911 B.n630 B.n81 163.367
R912 B.n626 B.n81 163.367
R913 B.n626 B.n625 163.367
R914 B.n625 B.n624 163.367
R915 B.n624 B.n83 163.367
R916 B.n620 B.n83 163.367
R917 B.n620 B.n619 163.367
R918 B.n619 B.n618 163.367
R919 B.n618 B.n85 163.367
R920 B.n614 B.n85 163.367
R921 B.n614 B.n613 163.367
R922 B.n613 B.n612 163.367
R923 B.n612 B.n87 163.367
R924 B.n608 B.n87 163.367
R925 B.n608 B.n607 163.367
R926 B.n607 B.n606 163.367
R927 B.n606 B.n89 163.367
R928 B.n602 B.n89 163.367
R929 B.n602 B.n601 163.367
R930 B.n601 B.n600 163.367
R931 B.n600 B.n91 163.367
R932 B.n596 B.n91 163.367
R933 B.n163 B.t10 112.538
R934 B.n61 B.t2 112.538
R935 B.n171 B.t4 112.514
R936 B.n53 B.t8 112.514
R937 B.n164 B.n163 59.5399
R938 B.n370 B.n171 59.5399
R939 B.n54 B.n53 59.5399
R940 B.n688 B.n61 59.5399
R941 B.n163 B.n162 51.3944
R942 B.n171 B.n170 51.3944
R943 B.n53 B.n52 51.3944
R944 B.n61 B.n60 51.3944
R945 B.n597 B.n92 36.3712
R946 B.n796 B.n795 36.3712
R947 B.n478 B.n477 36.3712
R948 B.n279 B.n202 36.3712
R949 B B.n855 18.0485
R950 B.n795 B.n22 10.6151
R951 B.n791 B.n22 10.6151
R952 B.n791 B.n790 10.6151
R953 B.n790 B.n789 10.6151
R954 B.n789 B.n24 10.6151
R955 B.n785 B.n24 10.6151
R956 B.n785 B.n784 10.6151
R957 B.n784 B.n783 10.6151
R958 B.n783 B.n26 10.6151
R959 B.n779 B.n26 10.6151
R960 B.n779 B.n778 10.6151
R961 B.n778 B.n777 10.6151
R962 B.n777 B.n28 10.6151
R963 B.n773 B.n28 10.6151
R964 B.n773 B.n772 10.6151
R965 B.n772 B.n771 10.6151
R966 B.n771 B.n30 10.6151
R967 B.n767 B.n30 10.6151
R968 B.n767 B.n766 10.6151
R969 B.n766 B.n765 10.6151
R970 B.n765 B.n32 10.6151
R971 B.n761 B.n32 10.6151
R972 B.n761 B.n760 10.6151
R973 B.n760 B.n759 10.6151
R974 B.n759 B.n34 10.6151
R975 B.n755 B.n34 10.6151
R976 B.n755 B.n754 10.6151
R977 B.n754 B.n753 10.6151
R978 B.n753 B.n36 10.6151
R979 B.n749 B.n36 10.6151
R980 B.n749 B.n748 10.6151
R981 B.n748 B.n747 10.6151
R982 B.n747 B.n38 10.6151
R983 B.n743 B.n38 10.6151
R984 B.n743 B.n742 10.6151
R985 B.n742 B.n741 10.6151
R986 B.n741 B.n40 10.6151
R987 B.n737 B.n40 10.6151
R988 B.n737 B.n736 10.6151
R989 B.n736 B.n735 10.6151
R990 B.n735 B.n42 10.6151
R991 B.n731 B.n42 10.6151
R992 B.n731 B.n730 10.6151
R993 B.n730 B.n729 10.6151
R994 B.n729 B.n44 10.6151
R995 B.n725 B.n44 10.6151
R996 B.n725 B.n724 10.6151
R997 B.n724 B.n723 10.6151
R998 B.n723 B.n46 10.6151
R999 B.n719 B.n46 10.6151
R1000 B.n719 B.n718 10.6151
R1001 B.n718 B.n717 10.6151
R1002 B.n717 B.n48 10.6151
R1003 B.n713 B.n48 10.6151
R1004 B.n713 B.n712 10.6151
R1005 B.n712 B.n711 10.6151
R1006 B.n711 B.n50 10.6151
R1007 B.n707 B.n50 10.6151
R1008 B.n707 B.n706 10.6151
R1009 B.n706 B.n705 10.6151
R1010 B.n702 B.n701 10.6151
R1011 B.n701 B.n700 10.6151
R1012 B.n700 B.n56 10.6151
R1013 B.n696 B.n56 10.6151
R1014 B.n696 B.n695 10.6151
R1015 B.n695 B.n694 10.6151
R1016 B.n694 B.n58 10.6151
R1017 B.n690 B.n58 10.6151
R1018 B.n690 B.n689 10.6151
R1019 B.n687 B.n62 10.6151
R1020 B.n683 B.n62 10.6151
R1021 B.n683 B.n682 10.6151
R1022 B.n682 B.n681 10.6151
R1023 B.n681 B.n64 10.6151
R1024 B.n677 B.n64 10.6151
R1025 B.n677 B.n676 10.6151
R1026 B.n676 B.n675 10.6151
R1027 B.n675 B.n66 10.6151
R1028 B.n671 B.n66 10.6151
R1029 B.n671 B.n670 10.6151
R1030 B.n670 B.n669 10.6151
R1031 B.n669 B.n68 10.6151
R1032 B.n665 B.n68 10.6151
R1033 B.n665 B.n664 10.6151
R1034 B.n664 B.n663 10.6151
R1035 B.n663 B.n70 10.6151
R1036 B.n659 B.n70 10.6151
R1037 B.n659 B.n658 10.6151
R1038 B.n658 B.n657 10.6151
R1039 B.n657 B.n72 10.6151
R1040 B.n653 B.n72 10.6151
R1041 B.n653 B.n652 10.6151
R1042 B.n652 B.n651 10.6151
R1043 B.n651 B.n74 10.6151
R1044 B.n647 B.n74 10.6151
R1045 B.n647 B.n646 10.6151
R1046 B.n646 B.n645 10.6151
R1047 B.n645 B.n76 10.6151
R1048 B.n641 B.n76 10.6151
R1049 B.n641 B.n640 10.6151
R1050 B.n640 B.n639 10.6151
R1051 B.n639 B.n78 10.6151
R1052 B.n635 B.n78 10.6151
R1053 B.n635 B.n634 10.6151
R1054 B.n634 B.n633 10.6151
R1055 B.n633 B.n80 10.6151
R1056 B.n629 B.n80 10.6151
R1057 B.n629 B.n628 10.6151
R1058 B.n628 B.n627 10.6151
R1059 B.n627 B.n82 10.6151
R1060 B.n623 B.n82 10.6151
R1061 B.n623 B.n622 10.6151
R1062 B.n622 B.n621 10.6151
R1063 B.n621 B.n84 10.6151
R1064 B.n617 B.n84 10.6151
R1065 B.n617 B.n616 10.6151
R1066 B.n616 B.n615 10.6151
R1067 B.n615 B.n86 10.6151
R1068 B.n611 B.n86 10.6151
R1069 B.n611 B.n610 10.6151
R1070 B.n610 B.n609 10.6151
R1071 B.n609 B.n88 10.6151
R1072 B.n605 B.n88 10.6151
R1073 B.n605 B.n604 10.6151
R1074 B.n604 B.n603 10.6151
R1075 B.n603 B.n90 10.6151
R1076 B.n599 B.n90 10.6151
R1077 B.n599 B.n598 10.6151
R1078 B.n598 B.n597 10.6151
R1079 B.n479 B.n478 10.6151
R1080 B.n479 B.n130 10.6151
R1081 B.n483 B.n130 10.6151
R1082 B.n484 B.n483 10.6151
R1083 B.n485 B.n484 10.6151
R1084 B.n485 B.n128 10.6151
R1085 B.n489 B.n128 10.6151
R1086 B.n490 B.n489 10.6151
R1087 B.n491 B.n490 10.6151
R1088 B.n491 B.n126 10.6151
R1089 B.n495 B.n126 10.6151
R1090 B.n496 B.n495 10.6151
R1091 B.n497 B.n496 10.6151
R1092 B.n497 B.n124 10.6151
R1093 B.n501 B.n124 10.6151
R1094 B.n502 B.n501 10.6151
R1095 B.n503 B.n502 10.6151
R1096 B.n503 B.n122 10.6151
R1097 B.n507 B.n122 10.6151
R1098 B.n508 B.n507 10.6151
R1099 B.n509 B.n508 10.6151
R1100 B.n509 B.n120 10.6151
R1101 B.n513 B.n120 10.6151
R1102 B.n514 B.n513 10.6151
R1103 B.n515 B.n514 10.6151
R1104 B.n515 B.n118 10.6151
R1105 B.n519 B.n118 10.6151
R1106 B.n520 B.n519 10.6151
R1107 B.n521 B.n520 10.6151
R1108 B.n521 B.n116 10.6151
R1109 B.n525 B.n116 10.6151
R1110 B.n526 B.n525 10.6151
R1111 B.n527 B.n526 10.6151
R1112 B.n527 B.n114 10.6151
R1113 B.n531 B.n114 10.6151
R1114 B.n532 B.n531 10.6151
R1115 B.n533 B.n532 10.6151
R1116 B.n533 B.n112 10.6151
R1117 B.n537 B.n112 10.6151
R1118 B.n538 B.n537 10.6151
R1119 B.n539 B.n538 10.6151
R1120 B.n539 B.n110 10.6151
R1121 B.n543 B.n110 10.6151
R1122 B.n544 B.n543 10.6151
R1123 B.n545 B.n544 10.6151
R1124 B.n545 B.n108 10.6151
R1125 B.n549 B.n108 10.6151
R1126 B.n550 B.n549 10.6151
R1127 B.n551 B.n550 10.6151
R1128 B.n551 B.n106 10.6151
R1129 B.n555 B.n106 10.6151
R1130 B.n556 B.n555 10.6151
R1131 B.n557 B.n556 10.6151
R1132 B.n557 B.n104 10.6151
R1133 B.n561 B.n104 10.6151
R1134 B.n562 B.n561 10.6151
R1135 B.n563 B.n562 10.6151
R1136 B.n563 B.n102 10.6151
R1137 B.n567 B.n102 10.6151
R1138 B.n568 B.n567 10.6151
R1139 B.n569 B.n568 10.6151
R1140 B.n569 B.n100 10.6151
R1141 B.n573 B.n100 10.6151
R1142 B.n574 B.n573 10.6151
R1143 B.n575 B.n574 10.6151
R1144 B.n575 B.n98 10.6151
R1145 B.n579 B.n98 10.6151
R1146 B.n580 B.n579 10.6151
R1147 B.n581 B.n580 10.6151
R1148 B.n581 B.n96 10.6151
R1149 B.n585 B.n96 10.6151
R1150 B.n586 B.n585 10.6151
R1151 B.n587 B.n586 10.6151
R1152 B.n587 B.n94 10.6151
R1153 B.n591 B.n94 10.6151
R1154 B.n592 B.n591 10.6151
R1155 B.n593 B.n592 10.6151
R1156 B.n593 B.n92 10.6151
R1157 B.n280 B.n279 10.6151
R1158 B.n281 B.n280 10.6151
R1159 B.n281 B.n200 10.6151
R1160 B.n285 B.n200 10.6151
R1161 B.n286 B.n285 10.6151
R1162 B.n287 B.n286 10.6151
R1163 B.n287 B.n198 10.6151
R1164 B.n291 B.n198 10.6151
R1165 B.n292 B.n291 10.6151
R1166 B.n293 B.n292 10.6151
R1167 B.n293 B.n196 10.6151
R1168 B.n297 B.n196 10.6151
R1169 B.n298 B.n297 10.6151
R1170 B.n299 B.n298 10.6151
R1171 B.n299 B.n194 10.6151
R1172 B.n303 B.n194 10.6151
R1173 B.n304 B.n303 10.6151
R1174 B.n305 B.n304 10.6151
R1175 B.n305 B.n192 10.6151
R1176 B.n309 B.n192 10.6151
R1177 B.n310 B.n309 10.6151
R1178 B.n311 B.n310 10.6151
R1179 B.n311 B.n190 10.6151
R1180 B.n315 B.n190 10.6151
R1181 B.n316 B.n315 10.6151
R1182 B.n317 B.n316 10.6151
R1183 B.n317 B.n188 10.6151
R1184 B.n321 B.n188 10.6151
R1185 B.n322 B.n321 10.6151
R1186 B.n323 B.n322 10.6151
R1187 B.n323 B.n186 10.6151
R1188 B.n327 B.n186 10.6151
R1189 B.n328 B.n327 10.6151
R1190 B.n329 B.n328 10.6151
R1191 B.n329 B.n184 10.6151
R1192 B.n333 B.n184 10.6151
R1193 B.n334 B.n333 10.6151
R1194 B.n335 B.n334 10.6151
R1195 B.n335 B.n182 10.6151
R1196 B.n339 B.n182 10.6151
R1197 B.n340 B.n339 10.6151
R1198 B.n341 B.n340 10.6151
R1199 B.n341 B.n180 10.6151
R1200 B.n345 B.n180 10.6151
R1201 B.n346 B.n345 10.6151
R1202 B.n347 B.n346 10.6151
R1203 B.n347 B.n178 10.6151
R1204 B.n351 B.n178 10.6151
R1205 B.n352 B.n351 10.6151
R1206 B.n353 B.n352 10.6151
R1207 B.n353 B.n176 10.6151
R1208 B.n357 B.n176 10.6151
R1209 B.n358 B.n357 10.6151
R1210 B.n359 B.n358 10.6151
R1211 B.n359 B.n174 10.6151
R1212 B.n363 B.n174 10.6151
R1213 B.n364 B.n363 10.6151
R1214 B.n365 B.n364 10.6151
R1215 B.n365 B.n172 10.6151
R1216 B.n369 B.n172 10.6151
R1217 B.n372 B.n371 10.6151
R1218 B.n372 B.n168 10.6151
R1219 B.n376 B.n168 10.6151
R1220 B.n377 B.n376 10.6151
R1221 B.n378 B.n377 10.6151
R1222 B.n378 B.n166 10.6151
R1223 B.n382 B.n166 10.6151
R1224 B.n383 B.n382 10.6151
R1225 B.n384 B.n383 10.6151
R1226 B.n388 B.n387 10.6151
R1227 B.n389 B.n388 10.6151
R1228 B.n389 B.n160 10.6151
R1229 B.n393 B.n160 10.6151
R1230 B.n394 B.n393 10.6151
R1231 B.n395 B.n394 10.6151
R1232 B.n395 B.n158 10.6151
R1233 B.n399 B.n158 10.6151
R1234 B.n400 B.n399 10.6151
R1235 B.n401 B.n400 10.6151
R1236 B.n401 B.n156 10.6151
R1237 B.n405 B.n156 10.6151
R1238 B.n406 B.n405 10.6151
R1239 B.n407 B.n406 10.6151
R1240 B.n407 B.n154 10.6151
R1241 B.n411 B.n154 10.6151
R1242 B.n412 B.n411 10.6151
R1243 B.n413 B.n412 10.6151
R1244 B.n413 B.n152 10.6151
R1245 B.n417 B.n152 10.6151
R1246 B.n418 B.n417 10.6151
R1247 B.n419 B.n418 10.6151
R1248 B.n419 B.n150 10.6151
R1249 B.n423 B.n150 10.6151
R1250 B.n424 B.n423 10.6151
R1251 B.n425 B.n424 10.6151
R1252 B.n425 B.n148 10.6151
R1253 B.n429 B.n148 10.6151
R1254 B.n430 B.n429 10.6151
R1255 B.n431 B.n430 10.6151
R1256 B.n431 B.n146 10.6151
R1257 B.n435 B.n146 10.6151
R1258 B.n436 B.n435 10.6151
R1259 B.n437 B.n436 10.6151
R1260 B.n437 B.n144 10.6151
R1261 B.n441 B.n144 10.6151
R1262 B.n442 B.n441 10.6151
R1263 B.n443 B.n442 10.6151
R1264 B.n443 B.n142 10.6151
R1265 B.n447 B.n142 10.6151
R1266 B.n448 B.n447 10.6151
R1267 B.n449 B.n448 10.6151
R1268 B.n449 B.n140 10.6151
R1269 B.n453 B.n140 10.6151
R1270 B.n454 B.n453 10.6151
R1271 B.n455 B.n454 10.6151
R1272 B.n455 B.n138 10.6151
R1273 B.n459 B.n138 10.6151
R1274 B.n460 B.n459 10.6151
R1275 B.n461 B.n460 10.6151
R1276 B.n461 B.n136 10.6151
R1277 B.n465 B.n136 10.6151
R1278 B.n466 B.n465 10.6151
R1279 B.n467 B.n466 10.6151
R1280 B.n467 B.n134 10.6151
R1281 B.n471 B.n134 10.6151
R1282 B.n472 B.n471 10.6151
R1283 B.n473 B.n472 10.6151
R1284 B.n473 B.n132 10.6151
R1285 B.n477 B.n132 10.6151
R1286 B.n275 B.n202 10.6151
R1287 B.n275 B.n274 10.6151
R1288 B.n274 B.n273 10.6151
R1289 B.n273 B.n204 10.6151
R1290 B.n269 B.n204 10.6151
R1291 B.n269 B.n268 10.6151
R1292 B.n268 B.n267 10.6151
R1293 B.n267 B.n206 10.6151
R1294 B.n263 B.n206 10.6151
R1295 B.n263 B.n262 10.6151
R1296 B.n262 B.n261 10.6151
R1297 B.n261 B.n208 10.6151
R1298 B.n257 B.n208 10.6151
R1299 B.n257 B.n256 10.6151
R1300 B.n256 B.n255 10.6151
R1301 B.n255 B.n210 10.6151
R1302 B.n251 B.n210 10.6151
R1303 B.n251 B.n250 10.6151
R1304 B.n250 B.n249 10.6151
R1305 B.n249 B.n212 10.6151
R1306 B.n245 B.n212 10.6151
R1307 B.n245 B.n244 10.6151
R1308 B.n244 B.n243 10.6151
R1309 B.n243 B.n214 10.6151
R1310 B.n239 B.n214 10.6151
R1311 B.n239 B.n238 10.6151
R1312 B.n238 B.n237 10.6151
R1313 B.n237 B.n216 10.6151
R1314 B.n233 B.n216 10.6151
R1315 B.n233 B.n232 10.6151
R1316 B.n232 B.n231 10.6151
R1317 B.n231 B.n218 10.6151
R1318 B.n227 B.n218 10.6151
R1319 B.n227 B.n226 10.6151
R1320 B.n226 B.n225 10.6151
R1321 B.n225 B.n220 10.6151
R1322 B.n221 B.n220 10.6151
R1323 B.n221 B.n0 10.6151
R1324 B.n851 B.n1 10.6151
R1325 B.n851 B.n850 10.6151
R1326 B.n850 B.n849 10.6151
R1327 B.n849 B.n4 10.6151
R1328 B.n845 B.n4 10.6151
R1329 B.n845 B.n844 10.6151
R1330 B.n844 B.n843 10.6151
R1331 B.n843 B.n6 10.6151
R1332 B.n839 B.n6 10.6151
R1333 B.n839 B.n838 10.6151
R1334 B.n838 B.n837 10.6151
R1335 B.n837 B.n8 10.6151
R1336 B.n833 B.n8 10.6151
R1337 B.n833 B.n832 10.6151
R1338 B.n832 B.n831 10.6151
R1339 B.n831 B.n10 10.6151
R1340 B.n827 B.n10 10.6151
R1341 B.n827 B.n826 10.6151
R1342 B.n826 B.n825 10.6151
R1343 B.n825 B.n12 10.6151
R1344 B.n821 B.n12 10.6151
R1345 B.n821 B.n820 10.6151
R1346 B.n820 B.n819 10.6151
R1347 B.n819 B.n14 10.6151
R1348 B.n815 B.n14 10.6151
R1349 B.n815 B.n814 10.6151
R1350 B.n814 B.n813 10.6151
R1351 B.n813 B.n16 10.6151
R1352 B.n809 B.n16 10.6151
R1353 B.n809 B.n808 10.6151
R1354 B.n808 B.n807 10.6151
R1355 B.n807 B.n18 10.6151
R1356 B.n803 B.n18 10.6151
R1357 B.n803 B.n802 10.6151
R1358 B.n802 B.n801 10.6151
R1359 B.n801 B.n20 10.6151
R1360 B.n797 B.n20 10.6151
R1361 B.n797 B.n796 10.6151
R1362 B.n705 B.n54 9.36635
R1363 B.n688 B.n687 9.36635
R1364 B.n370 B.n369 9.36635
R1365 B.n387 B.n164 9.36635
R1366 B.n855 B.n0 2.81026
R1367 B.n855 B.n1 2.81026
R1368 B.n702 B.n54 1.24928
R1369 B.n689 B.n688 1.24928
R1370 B.n371 B.n370 1.24928
R1371 B.n384 B.n164 1.24928
R1372 VP.n9 VP.t3 226.968
R1373 VP.n30 VP.t2 194.15
R1374 VP.n20 VP.t1 194.15
R1375 VP.n38 VP.t4 194.15
R1376 VP.n10 VP.t0 194.15
R1377 VP.n18 VP.t5 194.15
R1378 VP.n11 VP.n8 161.3
R1379 VP.n13 VP.n12 161.3
R1380 VP.n14 VP.n7 161.3
R1381 VP.n16 VP.n15 161.3
R1382 VP.n17 VP.n6 161.3
R1383 VP.n37 VP.n0 161.3
R1384 VP.n36 VP.n35 161.3
R1385 VP.n34 VP.n1 161.3
R1386 VP.n33 VP.n32 161.3
R1387 VP.n31 VP.n2 161.3
R1388 VP.n30 VP.n29 161.3
R1389 VP.n28 VP.n3 161.3
R1390 VP.n27 VP.n26 161.3
R1391 VP.n25 VP.n4 161.3
R1392 VP.n24 VP.n23 161.3
R1393 VP.n22 VP.n5 161.3
R1394 VP.n21 VP.n20 103.416
R1395 VP.n39 VP.n38 103.416
R1396 VP.n19 VP.n18 103.416
R1397 VP.n26 VP.n25 56.5193
R1398 VP.n32 VP.n1 56.5193
R1399 VP.n12 VP.n7 56.5193
R1400 VP.n21 VP.n19 52.5564
R1401 VP.n10 VP.n9 47.8187
R1402 VP.n24 VP.n5 24.4675
R1403 VP.n25 VP.n24 24.4675
R1404 VP.n26 VP.n3 24.4675
R1405 VP.n30 VP.n3 24.4675
R1406 VP.n31 VP.n30 24.4675
R1407 VP.n32 VP.n31 24.4675
R1408 VP.n36 VP.n1 24.4675
R1409 VP.n37 VP.n36 24.4675
R1410 VP.n16 VP.n7 24.4675
R1411 VP.n17 VP.n16 24.4675
R1412 VP.n11 VP.n10 24.4675
R1413 VP.n12 VP.n11 24.4675
R1414 VP.n20 VP.n5 7.3406
R1415 VP.n38 VP.n37 7.3406
R1416 VP.n18 VP.n17 7.3406
R1417 VP.n9 VP.n8 7.01727
R1418 VP.n19 VP.n6 0.278367
R1419 VP.n22 VP.n21 0.278367
R1420 VP.n39 VP.n0 0.278367
R1421 VP.n13 VP.n8 0.189894
R1422 VP.n14 VP.n13 0.189894
R1423 VP.n15 VP.n14 0.189894
R1424 VP.n15 VP.n6 0.189894
R1425 VP.n23 VP.n22 0.189894
R1426 VP.n23 VP.n4 0.189894
R1427 VP.n27 VP.n4 0.189894
R1428 VP.n28 VP.n27 0.189894
R1429 VP.n29 VP.n28 0.189894
R1430 VP.n29 VP.n2 0.189894
R1431 VP.n33 VP.n2 0.189894
R1432 VP.n34 VP.n33 0.189894
R1433 VP.n35 VP.n34 0.189894
R1434 VP.n35 VP.n0 0.189894
R1435 VP VP.n39 0.153454
R1436 VDD1 VDD1.t2 73.7886
R1437 VDD1.n1 VDD1.t4 73.675
R1438 VDD1.n1 VDD1.n0 70.7935
R1439 VDD1.n3 VDD1.n2 70.2778
R1440 VDD1.n3 VDD1.n1 48.9772
R1441 VDD1.n2 VDD1.t5 1.73967
R1442 VDD1.n2 VDD1.t0 1.73967
R1443 VDD1.n0 VDD1.t3 1.73967
R1444 VDD1.n0 VDD1.t1 1.73967
R1445 VDD1 VDD1.n3 0.513431
C0 VN w_n3090_n4706# 5.92111f
C1 VP w_n3090_n4706# 6.31982f
C2 VN VDD1 0.150434f
C3 VN VTAIL 9.82494f
C4 VP VDD1 10.304701f
C5 VP VTAIL 9.83937f
C6 VN VDD2 10.024401f
C7 B VN 1.18661f
C8 VP VDD2 0.435252f
C9 w_n3090_n4706# VDD1 2.69231f
C10 VP B 1.85089f
C11 VTAIL w_n3090_n4706# 3.89922f
C12 VDD2 w_n3090_n4706# 2.76847f
C13 VTAIL VDD1 10.2375f
C14 B w_n3090_n4706# 11.1648f
C15 VDD2 VDD1 1.29937f
C16 B VDD1 2.54439f
C17 VTAIL VDD2 10.2844f
C18 B VTAIL 5.04473f
C19 VP VN 7.89849f
C20 B VDD2 2.61177f
C21 VDD2 VSUBS 2.029451f
C22 VDD1 VSUBS 2.489794f
C23 VTAIL VSUBS 1.380813f
C24 VN VSUBS 5.875071f
C25 VP VSUBS 2.960472f
C26 B VSUBS 4.924554f
C27 w_n3090_n4706# VSUBS 0.177724p
C28 VDD1.t2 VSUBS 4.30612f
C29 VDD1.t4 VSUBS 4.30471f
C30 VDD1.t3 VSUBS 0.395237f
C31 VDD1.t1 VSUBS 0.395237f
C32 VDD1.n0 VSUBS 3.31136f
C33 VDD1.n1 VSUBS 4.1827f
C34 VDD1.t5 VSUBS 0.395237f
C35 VDD1.t0 VSUBS 0.395237f
C36 VDD1.n2 VSUBS 3.30569f
C37 VDD1.n3 VSUBS 3.74731f
C38 VP.n0 VSUBS 0.039052f
C39 VP.t4 VSUBS 3.53528f
C40 VP.n1 VSUBS 0.037054f
C41 VP.n2 VSUBS 0.029621f
C42 VP.t2 VSUBS 3.53528f
C43 VP.n3 VSUBS 0.055206f
C44 VP.n4 VSUBS 0.029621f
C45 VP.n5 VSUBS 0.036127f
C46 VP.n6 VSUBS 0.039052f
C47 VP.t5 VSUBS 3.53528f
C48 VP.n7 VSUBS 0.037054f
C49 VP.n8 VSUBS 0.277575f
C50 VP.t0 VSUBS 3.53528f
C51 VP.t3 VSUBS 3.73698f
C52 VP.n9 VSUBS 1.29046f
C53 VP.n10 VSUBS 1.32295f
C54 VP.n11 VSUBS 0.055206f
C55 VP.n12 VSUBS 0.049435f
C56 VP.n13 VSUBS 0.029621f
C57 VP.n14 VSUBS 0.029621f
C58 VP.n15 VSUBS 0.029621f
C59 VP.n16 VSUBS 0.055206f
C60 VP.n17 VSUBS 0.036127f
C61 VP.n18 VSUBS 1.31106f
C62 VP.n19 VSUBS 1.76935f
C63 VP.t1 VSUBS 3.53528f
C64 VP.n20 VSUBS 1.31106f
C65 VP.n21 VSUBS 1.78961f
C66 VP.n22 VSUBS 0.039052f
C67 VP.n23 VSUBS 0.029621f
C68 VP.n24 VSUBS 0.055206f
C69 VP.n25 VSUBS 0.037054f
C70 VP.n26 VSUBS 0.049435f
C71 VP.n27 VSUBS 0.029621f
C72 VP.n28 VSUBS 0.029621f
C73 VP.n29 VSUBS 0.029621f
C74 VP.n30 VSUBS 1.25503f
C75 VP.n31 VSUBS 0.055206f
C76 VP.n32 VSUBS 0.049435f
C77 VP.n33 VSUBS 0.029621f
C78 VP.n34 VSUBS 0.029621f
C79 VP.n35 VSUBS 0.029621f
C80 VP.n36 VSUBS 0.055206f
C81 VP.n37 VSUBS 0.036127f
C82 VP.n38 VSUBS 1.31106f
C83 VP.n39 VSUBS 0.047251f
C84 B.n0 VSUBS 0.004588f
C85 B.n1 VSUBS 0.004588f
C86 B.n2 VSUBS 0.007256f
C87 B.n3 VSUBS 0.007256f
C88 B.n4 VSUBS 0.007256f
C89 B.n5 VSUBS 0.007256f
C90 B.n6 VSUBS 0.007256f
C91 B.n7 VSUBS 0.007256f
C92 B.n8 VSUBS 0.007256f
C93 B.n9 VSUBS 0.007256f
C94 B.n10 VSUBS 0.007256f
C95 B.n11 VSUBS 0.007256f
C96 B.n12 VSUBS 0.007256f
C97 B.n13 VSUBS 0.007256f
C98 B.n14 VSUBS 0.007256f
C99 B.n15 VSUBS 0.007256f
C100 B.n16 VSUBS 0.007256f
C101 B.n17 VSUBS 0.007256f
C102 B.n18 VSUBS 0.007256f
C103 B.n19 VSUBS 0.007256f
C104 B.n20 VSUBS 0.007256f
C105 B.n21 VSUBS 0.017749f
C106 B.n22 VSUBS 0.007256f
C107 B.n23 VSUBS 0.007256f
C108 B.n24 VSUBS 0.007256f
C109 B.n25 VSUBS 0.007256f
C110 B.n26 VSUBS 0.007256f
C111 B.n27 VSUBS 0.007256f
C112 B.n28 VSUBS 0.007256f
C113 B.n29 VSUBS 0.007256f
C114 B.n30 VSUBS 0.007256f
C115 B.n31 VSUBS 0.007256f
C116 B.n32 VSUBS 0.007256f
C117 B.n33 VSUBS 0.007256f
C118 B.n34 VSUBS 0.007256f
C119 B.n35 VSUBS 0.007256f
C120 B.n36 VSUBS 0.007256f
C121 B.n37 VSUBS 0.007256f
C122 B.n38 VSUBS 0.007256f
C123 B.n39 VSUBS 0.007256f
C124 B.n40 VSUBS 0.007256f
C125 B.n41 VSUBS 0.007256f
C126 B.n42 VSUBS 0.007256f
C127 B.n43 VSUBS 0.007256f
C128 B.n44 VSUBS 0.007256f
C129 B.n45 VSUBS 0.007256f
C130 B.n46 VSUBS 0.007256f
C131 B.n47 VSUBS 0.007256f
C132 B.n48 VSUBS 0.007256f
C133 B.n49 VSUBS 0.007256f
C134 B.n50 VSUBS 0.007256f
C135 B.n51 VSUBS 0.007256f
C136 B.t8 VSUBS 0.655743f
C137 B.t7 VSUBS 0.675559f
C138 B.t6 VSUBS 1.97154f
C139 B.n52 VSUBS 0.357227f
C140 B.n53 VSUBS 0.073549f
C141 B.n54 VSUBS 0.016811f
C142 B.n55 VSUBS 0.007256f
C143 B.n56 VSUBS 0.007256f
C144 B.n57 VSUBS 0.007256f
C145 B.n58 VSUBS 0.007256f
C146 B.n59 VSUBS 0.007256f
C147 B.t2 VSUBS 0.655718f
C148 B.t1 VSUBS 0.675539f
C149 B.t0 VSUBS 1.97154f
C150 B.n60 VSUBS 0.357246f
C151 B.n61 VSUBS 0.073573f
C152 B.n62 VSUBS 0.007256f
C153 B.n63 VSUBS 0.007256f
C154 B.n64 VSUBS 0.007256f
C155 B.n65 VSUBS 0.007256f
C156 B.n66 VSUBS 0.007256f
C157 B.n67 VSUBS 0.007256f
C158 B.n68 VSUBS 0.007256f
C159 B.n69 VSUBS 0.007256f
C160 B.n70 VSUBS 0.007256f
C161 B.n71 VSUBS 0.007256f
C162 B.n72 VSUBS 0.007256f
C163 B.n73 VSUBS 0.007256f
C164 B.n74 VSUBS 0.007256f
C165 B.n75 VSUBS 0.007256f
C166 B.n76 VSUBS 0.007256f
C167 B.n77 VSUBS 0.007256f
C168 B.n78 VSUBS 0.007256f
C169 B.n79 VSUBS 0.007256f
C170 B.n80 VSUBS 0.007256f
C171 B.n81 VSUBS 0.007256f
C172 B.n82 VSUBS 0.007256f
C173 B.n83 VSUBS 0.007256f
C174 B.n84 VSUBS 0.007256f
C175 B.n85 VSUBS 0.007256f
C176 B.n86 VSUBS 0.007256f
C177 B.n87 VSUBS 0.007256f
C178 B.n88 VSUBS 0.007256f
C179 B.n89 VSUBS 0.007256f
C180 B.n90 VSUBS 0.007256f
C181 B.n91 VSUBS 0.007256f
C182 B.n92 VSUBS 0.018519f
C183 B.n93 VSUBS 0.007256f
C184 B.n94 VSUBS 0.007256f
C185 B.n95 VSUBS 0.007256f
C186 B.n96 VSUBS 0.007256f
C187 B.n97 VSUBS 0.007256f
C188 B.n98 VSUBS 0.007256f
C189 B.n99 VSUBS 0.007256f
C190 B.n100 VSUBS 0.007256f
C191 B.n101 VSUBS 0.007256f
C192 B.n102 VSUBS 0.007256f
C193 B.n103 VSUBS 0.007256f
C194 B.n104 VSUBS 0.007256f
C195 B.n105 VSUBS 0.007256f
C196 B.n106 VSUBS 0.007256f
C197 B.n107 VSUBS 0.007256f
C198 B.n108 VSUBS 0.007256f
C199 B.n109 VSUBS 0.007256f
C200 B.n110 VSUBS 0.007256f
C201 B.n111 VSUBS 0.007256f
C202 B.n112 VSUBS 0.007256f
C203 B.n113 VSUBS 0.007256f
C204 B.n114 VSUBS 0.007256f
C205 B.n115 VSUBS 0.007256f
C206 B.n116 VSUBS 0.007256f
C207 B.n117 VSUBS 0.007256f
C208 B.n118 VSUBS 0.007256f
C209 B.n119 VSUBS 0.007256f
C210 B.n120 VSUBS 0.007256f
C211 B.n121 VSUBS 0.007256f
C212 B.n122 VSUBS 0.007256f
C213 B.n123 VSUBS 0.007256f
C214 B.n124 VSUBS 0.007256f
C215 B.n125 VSUBS 0.007256f
C216 B.n126 VSUBS 0.007256f
C217 B.n127 VSUBS 0.007256f
C218 B.n128 VSUBS 0.007256f
C219 B.n129 VSUBS 0.007256f
C220 B.n130 VSUBS 0.007256f
C221 B.n131 VSUBS 0.017749f
C222 B.n132 VSUBS 0.007256f
C223 B.n133 VSUBS 0.007256f
C224 B.n134 VSUBS 0.007256f
C225 B.n135 VSUBS 0.007256f
C226 B.n136 VSUBS 0.007256f
C227 B.n137 VSUBS 0.007256f
C228 B.n138 VSUBS 0.007256f
C229 B.n139 VSUBS 0.007256f
C230 B.n140 VSUBS 0.007256f
C231 B.n141 VSUBS 0.007256f
C232 B.n142 VSUBS 0.007256f
C233 B.n143 VSUBS 0.007256f
C234 B.n144 VSUBS 0.007256f
C235 B.n145 VSUBS 0.007256f
C236 B.n146 VSUBS 0.007256f
C237 B.n147 VSUBS 0.007256f
C238 B.n148 VSUBS 0.007256f
C239 B.n149 VSUBS 0.007256f
C240 B.n150 VSUBS 0.007256f
C241 B.n151 VSUBS 0.007256f
C242 B.n152 VSUBS 0.007256f
C243 B.n153 VSUBS 0.007256f
C244 B.n154 VSUBS 0.007256f
C245 B.n155 VSUBS 0.007256f
C246 B.n156 VSUBS 0.007256f
C247 B.n157 VSUBS 0.007256f
C248 B.n158 VSUBS 0.007256f
C249 B.n159 VSUBS 0.007256f
C250 B.n160 VSUBS 0.007256f
C251 B.n161 VSUBS 0.007256f
C252 B.t10 VSUBS 0.655718f
C253 B.t11 VSUBS 0.675539f
C254 B.t9 VSUBS 1.97154f
C255 B.n162 VSUBS 0.357246f
C256 B.n163 VSUBS 0.073573f
C257 B.n164 VSUBS 0.016811f
C258 B.n165 VSUBS 0.007256f
C259 B.n166 VSUBS 0.007256f
C260 B.n167 VSUBS 0.007256f
C261 B.n168 VSUBS 0.007256f
C262 B.n169 VSUBS 0.007256f
C263 B.t4 VSUBS 0.655743f
C264 B.t5 VSUBS 0.675559f
C265 B.t3 VSUBS 1.97154f
C266 B.n170 VSUBS 0.357227f
C267 B.n171 VSUBS 0.073549f
C268 B.n172 VSUBS 0.007256f
C269 B.n173 VSUBS 0.007256f
C270 B.n174 VSUBS 0.007256f
C271 B.n175 VSUBS 0.007256f
C272 B.n176 VSUBS 0.007256f
C273 B.n177 VSUBS 0.007256f
C274 B.n178 VSUBS 0.007256f
C275 B.n179 VSUBS 0.007256f
C276 B.n180 VSUBS 0.007256f
C277 B.n181 VSUBS 0.007256f
C278 B.n182 VSUBS 0.007256f
C279 B.n183 VSUBS 0.007256f
C280 B.n184 VSUBS 0.007256f
C281 B.n185 VSUBS 0.007256f
C282 B.n186 VSUBS 0.007256f
C283 B.n187 VSUBS 0.007256f
C284 B.n188 VSUBS 0.007256f
C285 B.n189 VSUBS 0.007256f
C286 B.n190 VSUBS 0.007256f
C287 B.n191 VSUBS 0.007256f
C288 B.n192 VSUBS 0.007256f
C289 B.n193 VSUBS 0.007256f
C290 B.n194 VSUBS 0.007256f
C291 B.n195 VSUBS 0.007256f
C292 B.n196 VSUBS 0.007256f
C293 B.n197 VSUBS 0.007256f
C294 B.n198 VSUBS 0.007256f
C295 B.n199 VSUBS 0.007256f
C296 B.n200 VSUBS 0.007256f
C297 B.n201 VSUBS 0.007256f
C298 B.n202 VSUBS 0.017749f
C299 B.n203 VSUBS 0.007256f
C300 B.n204 VSUBS 0.007256f
C301 B.n205 VSUBS 0.007256f
C302 B.n206 VSUBS 0.007256f
C303 B.n207 VSUBS 0.007256f
C304 B.n208 VSUBS 0.007256f
C305 B.n209 VSUBS 0.007256f
C306 B.n210 VSUBS 0.007256f
C307 B.n211 VSUBS 0.007256f
C308 B.n212 VSUBS 0.007256f
C309 B.n213 VSUBS 0.007256f
C310 B.n214 VSUBS 0.007256f
C311 B.n215 VSUBS 0.007256f
C312 B.n216 VSUBS 0.007256f
C313 B.n217 VSUBS 0.007256f
C314 B.n218 VSUBS 0.007256f
C315 B.n219 VSUBS 0.007256f
C316 B.n220 VSUBS 0.007256f
C317 B.n221 VSUBS 0.007256f
C318 B.n222 VSUBS 0.007256f
C319 B.n223 VSUBS 0.007256f
C320 B.n224 VSUBS 0.007256f
C321 B.n225 VSUBS 0.007256f
C322 B.n226 VSUBS 0.007256f
C323 B.n227 VSUBS 0.007256f
C324 B.n228 VSUBS 0.007256f
C325 B.n229 VSUBS 0.007256f
C326 B.n230 VSUBS 0.007256f
C327 B.n231 VSUBS 0.007256f
C328 B.n232 VSUBS 0.007256f
C329 B.n233 VSUBS 0.007256f
C330 B.n234 VSUBS 0.007256f
C331 B.n235 VSUBS 0.007256f
C332 B.n236 VSUBS 0.007256f
C333 B.n237 VSUBS 0.007256f
C334 B.n238 VSUBS 0.007256f
C335 B.n239 VSUBS 0.007256f
C336 B.n240 VSUBS 0.007256f
C337 B.n241 VSUBS 0.007256f
C338 B.n242 VSUBS 0.007256f
C339 B.n243 VSUBS 0.007256f
C340 B.n244 VSUBS 0.007256f
C341 B.n245 VSUBS 0.007256f
C342 B.n246 VSUBS 0.007256f
C343 B.n247 VSUBS 0.007256f
C344 B.n248 VSUBS 0.007256f
C345 B.n249 VSUBS 0.007256f
C346 B.n250 VSUBS 0.007256f
C347 B.n251 VSUBS 0.007256f
C348 B.n252 VSUBS 0.007256f
C349 B.n253 VSUBS 0.007256f
C350 B.n254 VSUBS 0.007256f
C351 B.n255 VSUBS 0.007256f
C352 B.n256 VSUBS 0.007256f
C353 B.n257 VSUBS 0.007256f
C354 B.n258 VSUBS 0.007256f
C355 B.n259 VSUBS 0.007256f
C356 B.n260 VSUBS 0.007256f
C357 B.n261 VSUBS 0.007256f
C358 B.n262 VSUBS 0.007256f
C359 B.n263 VSUBS 0.007256f
C360 B.n264 VSUBS 0.007256f
C361 B.n265 VSUBS 0.007256f
C362 B.n266 VSUBS 0.007256f
C363 B.n267 VSUBS 0.007256f
C364 B.n268 VSUBS 0.007256f
C365 B.n269 VSUBS 0.007256f
C366 B.n270 VSUBS 0.007256f
C367 B.n271 VSUBS 0.007256f
C368 B.n272 VSUBS 0.007256f
C369 B.n273 VSUBS 0.007256f
C370 B.n274 VSUBS 0.007256f
C371 B.n275 VSUBS 0.007256f
C372 B.n276 VSUBS 0.007256f
C373 B.n277 VSUBS 0.017749f
C374 B.n278 VSUBS 0.018744f
C375 B.n279 VSUBS 0.018744f
C376 B.n280 VSUBS 0.007256f
C377 B.n281 VSUBS 0.007256f
C378 B.n282 VSUBS 0.007256f
C379 B.n283 VSUBS 0.007256f
C380 B.n284 VSUBS 0.007256f
C381 B.n285 VSUBS 0.007256f
C382 B.n286 VSUBS 0.007256f
C383 B.n287 VSUBS 0.007256f
C384 B.n288 VSUBS 0.007256f
C385 B.n289 VSUBS 0.007256f
C386 B.n290 VSUBS 0.007256f
C387 B.n291 VSUBS 0.007256f
C388 B.n292 VSUBS 0.007256f
C389 B.n293 VSUBS 0.007256f
C390 B.n294 VSUBS 0.007256f
C391 B.n295 VSUBS 0.007256f
C392 B.n296 VSUBS 0.007256f
C393 B.n297 VSUBS 0.007256f
C394 B.n298 VSUBS 0.007256f
C395 B.n299 VSUBS 0.007256f
C396 B.n300 VSUBS 0.007256f
C397 B.n301 VSUBS 0.007256f
C398 B.n302 VSUBS 0.007256f
C399 B.n303 VSUBS 0.007256f
C400 B.n304 VSUBS 0.007256f
C401 B.n305 VSUBS 0.007256f
C402 B.n306 VSUBS 0.007256f
C403 B.n307 VSUBS 0.007256f
C404 B.n308 VSUBS 0.007256f
C405 B.n309 VSUBS 0.007256f
C406 B.n310 VSUBS 0.007256f
C407 B.n311 VSUBS 0.007256f
C408 B.n312 VSUBS 0.007256f
C409 B.n313 VSUBS 0.007256f
C410 B.n314 VSUBS 0.007256f
C411 B.n315 VSUBS 0.007256f
C412 B.n316 VSUBS 0.007256f
C413 B.n317 VSUBS 0.007256f
C414 B.n318 VSUBS 0.007256f
C415 B.n319 VSUBS 0.007256f
C416 B.n320 VSUBS 0.007256f
C417 B.n321 VSUBS 0.007256f
C418 B.n322 VSUBS 0.007256f
C419 B.n323 VSUBS 0.007256f
C420 B.n324 VSUBS 0.007256f
C421 B.n325 VSUBS 0.007256f
C422 B.n326 VSUBS 0.007256f
C423 B.n327 VSUBS 0.007256f
C424 B.n328 VSUBS 0.007256f
C425 B.n329 VSUBS 0.007256f
C426 B.n330 VSUBS 0.007256f
C427 B.n331 VSUBS 0.007256f
C428 B.n332 VSUBS 0.007256f
C429 B.n333 VSUBS 0.007256f
C430 B.n334 VSUBS 0.007256f
C431 B.n335 VSUBS 0.007256f
C432 B.n336 VSUBS 0.007256f
C433 B.n337 VSUBS 0.007256f
C434 B.n338 VSUBS 0.007256f
C435 B.n339 VSUBS 0.007256f
C436 B.n340 VSUBS 0.007256f
C437 B.n341 VSUBS 0.007256f
C438 B.n342 VSUBS 0.007256f
C439 B.n343 VSUBS 0.007256f
C440 B.n344 VSUBS 0.007256f
C441 B.n345 VSUBS 0.007256f
C442 B.n346 VSUBS 0.007256f
C443 B.n347 VSUBS 0.007256f
C444 B.n348 VSUBS 0.007256f
C445 B.n349 VSUBS 0.007256f
C446 B.n350 VSUBS 0.007256f
C447 B.n351 VSUBS 0.007256f
C448 B.n352 VSUBS 0.007256f
C449 B.n353 VSUBS 0.007256f
C450 B.n354 VSUBS 0.007256f
C451 B.n355 VSUBS 0.007256f
C452 B.n356 VSUBS 0.007256f
C453 B.n357 VSUBS 0.007256f
C454 B.n358 VSUBS 0.007256f
C455 B.n359 VSUBS 0.007256f
C456 B.n360 VSUBS 0.007256f
C457 B.n361 VSUBS 0.007256f
C458 B.n362 VSUBS 0.007256f
C459 B.n363 VSUBS 0.007256f
C460 B.n364 VSUBS 0.007256f
C461 B.n365 VSUBS 0.007256f
C462 B.n366 VSUBS 0.007256f
C463 B.n367 VSUBS 0.007256f
C464 B.n368 VSUBS 0.007256f
C465 B.n369 VSUBS 0.006829f
C466 B.n370 VSUBS 0.016811f
C467 B.n371 VSUBS 0.004055f
C468 B.n372 VSUBS 0.007256f
C469 B.n373 VSUBS 0.007256f
C470 B.n374 VSUBS 0.007256f
C471 B.n375 VSUBS 0.007256f
C472 B.n376 VSUBS 0.007256f
C473 B.n377 VSUBS 0.007256f
C474 B.n378 VSUBS 0.007256f
C475 B.n379 VSUBS 0.007256f
C476 B.n380 VSUBS 0.007256f
C477 B.n381 VSUBS 0.007256f
C478 B.n382 VSUBS 0.007256f
C479 B.n383 VSUBS 0.007256f
C480 B.n384 VSUBS 0.004055f
C481 B.n385 VSUBS 0.007256f
C482 B.n386 VSUBS 0.007256f
C483 B.n387 VSUBS 0.006829f
C484 B.n388 VSUBS 0.007256f
C485 B.n389 VSUBS 0.007256f
C486 B.n390 VSUBS 0.007256f
C487 B.n391 VSUBS 0.007256f
C488 B.n392 VSUBS 0.007256f
C489 B.n393 VSUBS 0.007256f
C490 B.n394 VSUBS 0.007256f
C491 B.n395 VSUBS 0.007256f
C492 B.n396 VSUBS 0.007256f
C493 B.n397 VSUBS 0.007256f
C494 B.n398 VSUBS 0.007256f
C495 B.n399 VSUBS 0.007256f
C496 B.n400 VSUBS 0.007256f
C497 B.n401 VSUBS 0.007256f
C498 B.n402 VSUBS 0.007256f
C499 B.n403 VSUBS 0.007256f
C500 B.n404 VSUBS 0.007256f
C501 B.n405 VSUBS 0.007256f
C502 B.n406 VSUBS 0.007256f
C503 B.n407 VSUBS 0.007256f
C504 B.n408 VSUBS 0.007256f
C505 B.n409 VSUBS 0.007256f
C506 B.n410 VSUBS 0.007256f
C507 B.n411 VSUBS 0.007256f
C508 B.n412 VSUBS 0.007256f
C509 B.n413 VSUBS 0.007256f
C510 B.n414 VSUBS 0.007256f
C511 B.n415 VSUBS 0.007256f
C512 B.n416 VSUBS 0.007256f
C513 B.n417 VSUBS 0.007256f
C514 B.n418 VSUBS 0.007256f
C515 B.n419 VSUBS 0.007256f
C516 B.n420 VSUBS 0.007256f
C517 B.n421 VSUBS 0.007256f
C518 B.n422 VSUBS 0.007256f
C519 B.n423 VSUBS 0.007256f
C520 B.n424 VSUBS 0.007256f
C521 B.n425 VSUBS 0.007256f
C522 B.n426 VSUBS 0.007256f
C523 B.n427 VSUBS 0.007256f
C524 B.n428 VSUBS 0.007256f
C525 B.n429 VSUBS 0.007256f
C526 B.n430 VSUBS 0.007256f
C527 B.n431 VSUBS 0.007256f
C528 B.n432 VSUBS 0.007256f
C529 B.n433 VSUBS 0.007256f
C530 B.n434 VSUBS 0.007256f
C531 B.n435 VSUBS 0.007256f
C532 B.n436 VSUBS 0.007256f
C533 B.n437 VSUBS 0.007256f
C534 B.n438 VSUBS 0.007256f
C535 B.n439 VSUBS 0.007256f
C536 B.n440 VSUBS 0.007256f
C537 B.n441 VSUBS 0.007256f
C538 B.n442 VSUBS 0.007256f
C539 B.n443 VSUBS 0.007256f
C540 B.n444 VSUBS 0.007256f
C541 B.n445 VSUBS 0.007256f
C542 B.n446 VSUBS 0.007256f
C543 B.n447 VSUBS 0.007256f
C544 B.n448 VSUBS 0.007256f
C545 B.n449 VSUBS 0.007256f
C546 B.n450 VSUBS 0.007256f
C547 B.n451 VSUBS 0.007256f
C548 B.n452 VSUBS 0.007256f
C549 B.n453 VSUBS 0.007256f
C550 B.n454 VSUBS 0.007256f
C551 B.n455 VSUBS 0.007256f
C552 B.n456 VSUBS 0.007256f
C553 B.n457 VSUBS 0.007256f
C554 B.n458 VSUBS 0.007256f
C555 B.n459 VSUBS 0.007256f
C556 B.n460 VSUBS 0.007256f
C557 B.n461 VSUBS 0.007256f
C558 B.n462 VSUBS 0.007256f
C559 B.n463 VSUBS 0.007256f
C560 B.n464 VSUBS 0.007256f
C561 B.n465 VSUBS 0.007256f
C562 B.n466 VSUBS 0.007256f
C563 B.n467 VSUBS 0.007256f
C564 B.n468 VSUBS 0.007256f
C565 B.n469 VSUBS 0.007256f
C566 B.n470 VSUBS 0.007256f
C567 B.n471 VSUBS 0.007256f
C568 B.n472 VSUBS 0.007256f
C569 B.n473 VSUBS 0.007256f
C570 B.n474 VSUBS 0.007256f
C571 B.n475 VSUBS 0.007256f
C572 B.n476 VSUBS 0.018744f
C573 B.n477 VSUBS 0.018744f
C574 B.n478 VSUBS 0.017749f
C575 B.n479 VSUBS 0.007256f
C576 B.n480 VSUBS 0.007256f
C577 B.n481 VSUBS 0.007256f
C578 B.n482 VSUBS 0.007256f
C579 B.n483 VSUBS 0.007256f
C580 B.n484 VSUBS 0.007256f
C581 B.n485 VSUBS 0.007256f
C582 B.n486 VSUBS 0.007256f
C583 B.n487 VSUBS 0.007256f
C584 B.n488 VSUBS 0.007256f
C585 B.n489 VSUBS 0.007256f
C586 B.n490 VSUBS 0.007256f
C587 B.n491 VSUBS 0.007256f
C588 B.n492 VSUBS 0.007256f
C589 B.n493 VSUBS 0.007256f
C590 B.n494 VSUBS 0.007256f
C591 B.n495 VSUBS 0.007256f
C592 B.n496 VSUBS 0.007256f
C593 B.n497 VSUBS 0.007256f
C594 B.n498 VSUBS 0.007256f
C595 B.n499 VSUBS 0.007256f
C596 B.n500 VSUBS 0.007256f
C597 B.n501 VSUBS 0.007256f
C598 B.n502 VSUBS 0.007256f
C599 B.n503 VSUBS 0.007256f
C600 B.n504 VSUBS 0.007256f
C601 B.n505 VSUBS 0.007256f
C602 B.n506 VSUBS 0.007256f
C603 B.n507 VSUBS 0.007256f
C604 B.n508 VSUBS 0.007256f
C605 B.n509 VSUBS 0.007256f
C606 B.n510 VSUBS 0.007256f
C607 B.n511 VSUBS 0.007256f
C608 B.n512 VSUBS 0.007256f
C609 B.n513 VSUBS 0.007256f
C610 B.n514 VSUBS 0.007256f
C611 B.n515 VSUBS 0.007256f
C612 B.n516 VSUBS 0.007256f
C613 B.n517 VSUBS 0.007256f
C614 B.n518 VSUBS 0.007256f
C615 B.n519 VSUBS 0.007256f
C616 B.n520 VSUBS 0.007256f
C617 B.n521 VSUBS 0.007256f
C618 B.n522 VSUBS 0.007256f
C619 B.n523 VSUBS 0.007256f
C620 B.n524 VSUBS 0.007256f
C621 B.n525 VSUBS 0.007256f
C622 B.n526 VSUBS 0.007256f
C623 B.n527 VSUBS 0.007256f
C624 B.n528 VSUBS 0.007256f
C625 B.n529 VSUBS 0.007256f
C626 B.n530 VSUBS 0.007256f
C627 B.n531 VSUBS 0.007256f
C628 B.n532 VSUBS 0.007256f
C629 B.n533 VSUBS 0.007256f
C630 B.n534 VSUBS 0.007256f
C631 B.n535 VSUBS 0.007256f
C632 B.n536 VSUBS 0.007256f
C633 B.n537 VSUBS 0.007256f
C634 B.n538 VSUBS 0.007256f
C635 B.n539 VSUBS 0.007256f
C636 B.n540 VSUBS 0.007256f
C637 B.n541 VSUBS 0.007256f
C638 B.n542 VSUBS 0.007256f
C639 B.n543 VSUBS 0.007256f
C640 B.n544 VSUBS 0.007256f
C641 B.n545 VSUBS 0.007256f
C642 B.n546 VSUBS 0.007256f
C643 B.n547 VSUBS 0.007256f
C644 B.n548 VSUBS 0.007256f
C645 B.n549 VSUBS 0.007256f
C646 B.n550 VSUBS 0.007256f
C647 B.n551 VSUBS 0.007256f
C648 B.n552 VSUBS 0.007256f
C649 B.n553 VSUBS 0.007256f
C650 B.n554 VSUBS 0.007256f
C651 B.n555 VSUBS 0.007256f
C652 B.n556 VSUBS 0.007256f
C653 B.n557 VSUBS 0.007256f
C654 B.n558 VSUBS 0.007256f
C655 B.n559 VSUBS 0.007256f
C656 B.n560 VSUBS 0.007256f
C657 B.n561 VSUBS 0.007256f
C658 B.n562 VSUBS 0.007256f
C659 B.n563 VSUBS 0.007256f
C660 B.n564 VSUBS 0.007256f
C661 B.n565 VSUBS 0.007256f
C662 B.n566 VSUBS 0.007256f
C663 B.n567 VSUBS 0.007256f
C664 B.n568 VSUBS 0.007256f
C665 B.n569 VSUBS 0.007256f
C666 B.n570 VSUBS 0.007256f
C667 B.n571 VSUBS 0.007256f
C668 B.n572 VSUBS 0.007256f
C669 B.n573 VSUBS 0.007256f
C670 B.n574 VSUBS 0.007256f
C671 B.n575 VSUBS 0.007256f
C672 B.n576 VSUBS 0.007256f
C673 B.n577 VSUBS 0.007256f
C674 B.n578 VSUBS 0.007256f
C675 B.n579 VSUBS 0.007256f
C676 B.n580 VSUBS 0.007256f
C677 B.n581 VSUBS 0.007256f
C678 B.n582 VSUBS 0.007256f
C679 B.n583 VSUBS 0.007256f
C680 B.n584 VSUBS 0.007256f
C681 B.n585 VSUBS 0.007256f
C682 B.n586 VSUBS 0.007256f
C683 B.n587 VSUBS 0.007256f
C684 B.n588 VSUBS 0.007256f
C685 B.n589 VSUBS 0.007256f
C686 B.n590 VSUBS 0.007256f
C687 B.n591 VSUBS 0.007256f
C688 B.n592 VSUBS 0.007256f
C689 B.n593 VSUBS 0.007256f
C690 B.n594 VSUBS 0.007256f
C691 B.n595 VSUBS 0.017749f
C692 B.n596 VSUBS 0.018744f
C693 B.n597 VSUBS 0.017974f
C694 B.n598 VSUBS 0.007256f
C695 B.n599 VSUBS 0.007256f
C696 B.n600 VSUBS 0.007256f
C697 B.n601 VSUBS 0.007256f
C698 B.n602 VSUBS 0.007256f
C699 B.n603 VSUBS 0.007256f
C700 B.n604 VSUBS 0.007256f
C701 B.n605 VSUBS 0.007256f
C702 B.n606 VSUBS 0.007256f
C703 B.n607 VSUBS 0.007256f
C704 B.n608 VSUBS 0.007256f
C705 B.n609 VSUBS 0.007256f
C706 B.n610 VSUBS 0.007256f
C707 B.n611 VSUBS 0.007256f
C708 B.n612 VSUBS 0.007256f
C709 B.n613 VSUBS 0.007256f
C710 B.n614 VSUBS 0.007256f
C711 B.n615 VSUBS 0.007256f
C712 B.n616 VSUBS 0.007256f
C713 B.n617 VSUBS 0.007256f
C714 B.n618 VSUBS 0.007256f
C715 B.n619 VSUBS 0.007256f
C716 B.n620 VSUBS 0.007256f
C717 B.n621 VSUBS 0.007256f
C718 B.n622 VSUBS 0.007256f
C719 B.n623 VSUBS 0.007256f
C720 B.n624 VSUBS 0.007256f
C721 B.n625 VSUBS 0.007256f
C722 B.n626 VSUBS 0.007256f
C723 B.n627 VSUBS 0.007256f
C724 B.n628 VSUBS 0.007256f
C725 B.n629 VSUBS 0.007256f
C726 B.n630 VSUBS 0.007256f
C727 B.n631 VSUBS 0.007256f
C728 B.n632 VSUBS 0.007256f
C729 B.n633 VSUBS 0.007256f
C730 B.n634 VSUBS 0.007256f
C731 B.n635 VSUBS 0.007256f
C732 B.n636 VSUBS 0.007256f
C733 B.n637 VSUBS 0.007256f
C734 B.n638 VSUBS 0.007256f
C735 B.n639 VSUBS 0.007256f
C736 B.n640 VSUBS 0.007256f
C737 B.n641 VSUBS 0.007256f
C738 B.n642 VSUBS 0.007256f
C739 B.n643 VSUBS 0.007256f
C740 B.n644 VSUBS 0.007256f
C741 B.n645 VSUBS 0.007256f
C742 B.n646 VSUBS 0.007256f
C743 B.n647 VSUBS 0.007256f
C744 B.n648 VSUBS 0.007256f
C745 B.n649 VSUBS 0.007256f
C746 B.n650 VSUBS 0.007256f
C747 B.n651 VSUBS 0.007256f
C748 B.n652 VSUBS 0.007256f
C749 B.n653 VSUBS 0.007256f
C750 B.n654 VSUBS 0.007256f
C751 B.n655 VSUBS 0.007256f
C752 B.n656 VSUBS 0.007256f
C753 B.n657 VSUBS 0.007256f
C754 B.n658 VSUBS 0.007256f
C755 B.n659 VSUBS 0.007256f
C756 B.n660 VSUBS 0.007256f
C757 B.n661 VSUBS 0.007256f
C758 B.n662 VSUBS 0.007256f
C759 B.n663 VSUBS 0.007256f
C760 B.n664 VSUBS 0.007256f
C761 B.n665 VSUBS 0.007256f
C762 B.n666 VSUBS 0.007256f
C763 B.n667 VSUBS 0.007256f
C764 B.n668 VSUBS 0.007256f
C765 B.n669 VSUBS 0.007256f
C766 B.n670 VSUBS 0.007256f
C767 B.n671 VSUBS 0.007256f
C768 B.n672 VSUBS 0.007256f
C769 B.n673 VSUBS 0.007256f
C770 B.n674 VSUBS 0.007256f
C771 B.n675 VSUBS 0.007256f
C772 B.n676 VSUBS 0.007256f
C773 B.n677 VSUBS 0.007256f
C774 B.n678 VSUBS 0.007256f
C775 B.n679 VSUBS 0.007256f
C776 B.n680 VSUBS 0.007256f
C777 B.n681 VSUBS 0.007256f
C778 B.n682 VSUBS 0.007256f
C779 B.n683 VSUBS 0.007256f
C780 B.n684 VSUBS 0.007256f
C781 B.n685 VSUBS 0.007256f
C782 B.n686 VSUBS 0.007256f
C783 B.n687 VSUBS 0.006829f
C784 B.n688 VSUBS 0.016811f
C785 B.n689 VSUBS 0.004055f
C786 B.n690 VSUBS 0.007256f
C787 B.n691 VSUBS 0.007256f
C788 B.n692 VSUBS 0.007256f
C789 B.n693 VSUBS 0.007256f
C790 B.n694 VSUBS 0.007256f
C791 B.n695 VSUBS 0.007256f
C792 B.n696 VSUBS 0.007256f
C793 B.n697 VSUBS 0.007256f
C794 B.n698 VSUBS 0.007256f
C795 B.n699 VSUBS 0.007256f
C796 B.n700 VSUBS 0.007256f
C797 B.n701 VSUBS 0.007256f
C798 B.n702 VSUBS 0.004055f
C799 B.n703 VSUBS 0.007256f
C800 B.n704 VSUBS 0.007256f
C801 B.n705 VSUBS 0.006829f
C802 B.n706 VSUBS 0.007256f
C803 B.n707 VSUBS 0.007256f
C804 B.n708 VSUBS 0.007256f
C805 B.n709 VSUBS 0.007256f
C806 B.n710 VSUBS 0.007256f
C807 B.n711 VSUBS 0.007256f
C808 B.n712 VSUBS 0.007256f
C809 B.n713 VSUBS 0.007256f
C810 B.n714 VSUBS 0.007256f
C811 B.n715 VSUBS 0.007256f
C812 B.n716 VSUBS 0.007256f
C813 B.n717 VSUBS 0.007256f
C814 B.n718 VSUBS 0.007256f
C815 B.n719 VSUBS 0.007256f
C816 B.n720 VSUBS 0.007256f
C817 B.n721 VSUBS 0.007256f
C818 B.n722 VSUBS 0.007256f
C819 B.n723 VSUBS 0.007256f
C820 B.n724 VSUBS 0.007256f
C821 B.n725 VSUBS 0.007256f
C822 B.n726 VSUBS 0.007256f
C823 B.n727 VSUBS 0.007256f
C824 B.n728 VSUBS 0.007256f
C825 B.n729 VSUBS 0.007256f
C826 B.n730 VSUBS 0.007256f
C827 B.n731 VSUBS 0.007256f
C828 B.n732 VSUBS 0.007256f
C829 B.n733 VSUBS 0.007256f
C830 B.n734 VSUBS 0.007256f
C831 B.n735 VSUBS 0.007256f
C832 B.n736 VSUBS 0.007256f
C833 B.n737 VSUBS 0.007256f
C834 B.n738 VSUBS 0.007256f
C835 B.n739 VSUBS 0.007256f
C836 B.n740 VSUBS 0.007256f
C837 B.n741 VSUBS 0.007256f
C838 B.n742 VSUBS 0.007256f
C839 B.n743 VSUBS 0.007256f
C840 B.n744 VSUBS 0.007256f
C841 B.n745 VSUBS 0.007256f
C842 B.n746 VSUBS 0.007256f
C843 B.n747 VSUBS 0.007256f
C844 B.n748 VSUBS 0.007256f
C845 B.n749 VSUBS 0.007256f
C846 B.n750 VSUBS 0.007256f
C847 B.n751 VSUBS 0.007256f
C848 B.n752 VSUBS 0.007256f
C849 B.n753 VSUBS 0.007256f
C850 B.n754 VSUBS 0.007256f
C851 B.n755 VSUBS 0.007256f
C852 B.n756 VSUBS 0.007256f
C853 B.n757 VSUBS 0.007256f
C854 B.n758 VSUBS 0.007256f
C855 B.n759 VSUBS 0.007256f
C856 B.n760 VSUBS 0.007256f
C857 B.n761 VSUBS 0.007256f
C858 B.n762 VSUBS 0.007256f
C859 B.n763 VSUBS 0.007256f
C860 B.n764 VSUBS 0.007256f
C861 B.n765 VSUBS 0.007256f
C862 B.n766 VSUBS 0.007256f
C863 B.n767 VSUBS 0.007256f
C864 B.n768 VSUBS 0.007256f
C865 B.n769 VSUBS 0.007256f
C866 B.n770 VSUBS 0.007256f
C867 B.n771 VSUBS 0.007256f
C868 B.n772 VSUBS 0.007256f
C869 B.n773 VSUBS 0.007256f
C870 B.n774 VSUBS 0.007256f
C871 B.n775 VSUBS 0.007256f
C872 B.n776 VSUBS 0.007256f
C873 B.n777 VSUBS 0.007256f
C874 B.n778 VSUBS 0.007256f
C875 B.n779 VSUBS 0.007256f
C876 B.n780 VSUBS 0.007256f
C877 B.n781 VSUBS 0.007256f
C878 B.n782 VSUBS 0.007256f
C879 B.n783 VSUBS 0.007256f
C880 B.n784 VSUBS 0.007256f
C881 B.n785 VSUBS 0.007256f
C882 B.n786 VSUBS 0.007256f
C883 B.n787 VSUBS 0.007256f
C884 B.n788 VSUBS 0.007256f
C885 B.n789 VSUBS 0.007256f
C886 B.n790 VSUBS 0.007256f
C887 B.n791 VSUBS 0.007256f
C888 B.n792 VSUBS 0.007256f
C889 B.n793 VSUBS 0.007256f
C890 B.n794 VSUBS 0.018744f
C891 B.n795 VSUBS 0.018744f
C892 B.n796 VSUBS 0.017749f
C893 B.n797 VSUBS 0.007256f
C894 B.n798 VSUBS 0.007256f
C895 B.n799 VSUBS 0.007256f
C896 B.n800 VSUBS 0.007256f
C897 B.n801 VSUBS 0.007256f
C898 B.n802 VSUBS 0.007256f
C899 B.n803 VSUBS 0.007256f
C900 B.n804 VSUBS 0.007256f
C901 B.n805 VSUBS 0.007256f
C902 B.n806 VSUBS 0.007256f
C903 B.n807 VSUBS 0.007256f
C904 B.n808 VSUBS 0.007256f
C905 B.n809 VSUBS 0.007256f
C906 B.n810 VSUBS 0.007256f
C907 B.n811 VSUBS 0.007256f
C908 B.n812 VSUBS 0.007256f
C909 B.n813 VSUBS 0.007256f
C910 B.n814 VSUBS 0.007256f
C911 B.n815 VSUBS 0.007256f
C912 B.n816 VSUBS 0.007256f
C913 B.n817 VSUBS 0.007256f
C914 B.n818 VSUBS 0.007256f
C915 B.n819 VSUBS 0.007256f
C916 B.n820 VSUBS 0.007256f
C917 B.n821 VSUBS 0.007256f
C918 B.n822 VSUBS 0.007256f
C919 B.n823 VSUBS 0.007256f
C920 B.n824 VSUBS 0.007256f
C921 B.n825 VSUBS 0.007256f
C922 B.n826 VSUBS 0.007256f
C923 B.n827 VSUBS 0.007256f
C924 B.n828 VSUBS 0.007256f
C925 B.n829 VSUBS 0.007256f
C926 B.n830 VSUBS 0.007256f
C927 B.n831 VSUBS 0.007256f
C928 B.n832 VSUBS 0.007256f
C929 B.n833 VSUBS 0.007256f
C930 B.n834 VSUBS 0.007256f
C931 B.n835 VSUBS 0.007256f
C932 B.n836 VSUBS 0.007256f
C933 B.n837 VSUBS 0.007256f
C934 B.n838 VSUBS 0.007256f
C935 B.n839 VSUBS 0.007256f
C936 B.n840 VSUBS 0.007256f
C937 B.n841 VSUBS 0.007256f
C938 B.n842 VSUBS 0.007256f
C939 B.n843 VSUBS 0.007256f
C940 B.n844 VSUBS 0.007256f
C941 B.n845 VSUBS 0.007256f
C942 B.n846 VSUBS 0.007256f
C943 B.n847 VSUBS 0.007256f
C944 B.n848 VSUBS 0.007256f
C945 B.n849 VSUBS 0.007256f
C946 B.n850 VSUBS 0.007256f
C947 B.n851 VSUBS 0.007256f
C948 B.n852 VSUBS 0.007256f
C949 B.n853 VSUBS 0.007256f
C950 B.n854 VSUBS 0.007256f
C951 B.n855 VSUBS 0.01643f
C952 VTAIL.t9 VSUBS 0.402311f
C953 VTAIL.t11 VSUBS 0.402311f
C954 VTAIL.n0 VSUBS 3.20078f
C955 VTAIL.n1 VSUBS 0.856291f
C956 VTAIL.t0 VSUBS 4.17554f
C957 VTAIL.n2 VSUBS 1.12401f
C958 VTAIL.t2 VSUBS 0.402311f
C959 VTAIL.t1 VSUBS 0.402311f
C960 VTAIL.n3 VSUBS 3.20078f
C961 VTAIL.n4 VSUBS 3.0453f
C962 VTAIL.t8 VSUBS 0.402311f
C963 VTAIL.t10 VSUBS 0.402311f
C964 VTAIL.n5 VSUBS 3.20078f
C965 VTAIL.n6 VSUBS 3.04529f
C966 VTAIL.t7 VSUBS 4.17557f
C967 VTAIL.n7 VSUBS 1.12398f
C968 VTAIL.t3 VSUBS 0.402311f
C969 VTAIL.t5 VSUBS 0.402311f
C970 VTAIL.n8 VSUBS 3.20078f
C971 VTAIL.n9 VSUBS 1.00156f
C972 VTAIL.t4 VSUBS 4.17554f
C973 VTAIL.n10 VSUBS 2.96723f
C974 VTAIL.t6 VSUBS 4.17554f
C975 VTAIL.n11 VSUBS 2.912f
C976 VDD2.t5 VSUBS 4.32133f
C977 VDD2.t1 VSUBS 0.396763f
C978 VDD2.t4 VSUBS 0.396763f
C979 VDD2.n0 VSUBS 3.32415f
C980 VDD2.n1 VSUBS 4.0689f
C981 VDD2.t3 VSUBS 4.30387f
C982 VDD2.n2 VSUBS 3.80036f
C983 VDD2.t0 VSUBS 0.396763f
C984 VDD2.t2 VSUBS 0.396763f
C985 VDD2.n3 VSUBS 3.3241f
C986 VN.n0 VSUBS 0.038209f
C987 VN.t5 VSUBS 3.45893f
C988 VN.n1 VSUBS 0.036254f
C989 VN.n2 VSUBS 0.271581f
C990 VN.t0 VSUBS 3.45893f
C991 VN.t2 VSUBS 3.65628f
C992 VN.n3 VSUBS 1.26259f
C993 VN.n4 VSUBS 1.29438f
C994 VN.n5 VSUBS 0.054014f
C995 VN.n6 VSUBS 0.048367f
C996 VN.n7 VSUBS 0.028981f
C997 VN.n8 VSUBS 0.028981f
C998 VN.n9 VSUBS 0.028981f
C999 VN.n10 VSUBS 0.054014f
C1000 VN.n11 VSUBS 0.035347f
C1001 VN.n12 VSUBS 1.28274f
C1002 VN.n13 VSUBS 0.046231f
C1003 VN.n14 VSUBS 0.038209f
C1004 VN.t3 VSUBS 3.45893f
C1005 VN.n15 VSUBS 0.036254f
C1006 VN.n16 VSUBS 0.271581f
C1007 VN.t1 VSUBS 3.45893f
C1008 VN.t4 VSUBS 3.65628f
C1009 VN.n17 VSUBS 1.26259f
C1010 VN.n18 VSUBS 1.29438f
C1011 VN.n19 VSUBS 0.054014f
C1012 VN.n20 VSUBS 0.048367f
C1013 VN.n21 VSUBS 0.028981f
C1014 VN.n22 VSUBS 0.028981f
C1015 VN.n23 VSUBS 0.028981f
C1016 VN.n24 VSUBS 0.054014f
C1017 VN.n25 VSUBS 0.035347f
C1018 VN.n26 VSUBS 1.28274f
C1019 VN.n27 VSUBS 1.74659f
.ends

