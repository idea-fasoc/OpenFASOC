* NGSPICE file created from diff_pair_sample_0308.ext - technology: sky130A

.subckt diff_pair_sample_0308 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t16 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=0.31
X1 VTAIL.t3 VN.t0 VDD2.t9 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X2 B.t11 B.t9 B.t10 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=0.31
X3 VDD2.t8 VN.t1 VTAIL.t4 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=0.31
X4 VDD2.t7 VN.t2 VTAIL.t7 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=0.31
X5 B.t8 B.t6 B.t7 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=0.31
X6 VTAIL.t9 VP.t1 VDD1.t8 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X7 VDD1.t7 VP.t2 VTAIL.t10 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=0.31
X8 VTAIL.t12 VP.t3 VDD1.t6 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X9 VDD1.t5 VP.t4 VTAIL.t15 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X10 VDD1.t4 VP.t5 VTAIL.t11 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=3.0591 ps=18.87 w=18.54 l=0.31
X11 VDD2.t6 VN.t3 VTAIL.t2 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=0.31
X12 VTAIL.t18 VN.t4 VDD2.t5 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X13 VTAIL.t14 VP.t6 VDD1.t3 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X14 B.t5 B.t3 B.t4 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=0.31
X15 B.t2 B.t0 B.t1 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=7.2306 pd=37.86 as=0 ps=0 w=18.54 l=0.31
X16 VDD1.t2 VP.t7 VTAIL.t8 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=0.31
X17 VDD1.t1 VP.t8 VTAIL.t17 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X18 VDD2.t4 VN.t5 VTAIL.t19 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X19 VTAIL.t6 VN.t6 VDD2.t3 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X20 VDD2.t2 VN.t7 VTAIL.t0 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=7.2306 ps=37.86 w=18.54 l=0.31
X21 VTAIL.t5 VN.t8 VDD2.t1 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X22 VDD2.t0 VN.t9 VTAIL.t1 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
X23 VTAIL.t13 VP.t9 VDD1.t0 w_n1738_n4676# sky130_fd_pr__pfet_01v8 ad=3.0591 pd=18.87 as=3.0591 ps=18.87 w=18.54 l=0.31
R0 VP.n21 VP.t7 1583.3
R1 VP.n14 VP.t2 1583.3
R2 VP.n5 VP.t5 1583.3
R3 VP.n11 VP.t0 1583.3
R4 VP.n18 VP.t4 1542.4
R5 VP.n20 VP.t3 1542.4
R6 VP.n13 VP.t6 1542.4
R7 VP.n8 VP.t8 1542.4
R8 VP.n4 VP.t9 1542.4
R9 VP.n10 VP.t1 1542.4
R10 VP.n6 VP.n5 161.489
R11 VP.n22 VP.n21 161.3
R12 VP.n6 VP.n3 161.3
R13 VP.n8 VP.n7 161.3
R14 VP.n9 VP.n2 161.3
R15 VP.n12 VP.n11 161.3
R16 VP.n19 VP.n0 161.3
R17 VP.n18 VP.n17 161.3
R18 VP.n16 VP.n1 161.3
R19 VP.n15 VP.n14 161.3
R20 VP.n18 VP.n1 73.0308
R21 VP.n19 VP.n18 73.0308
R22 VP.n8 VP.n3 73.0308
R23 VP.n9 VP.n8 73.0308
R24 VP.n14 VP.n13 52.5823
R25 VP.n21 VP.n20 52.5823
R26 VP.n5 VP.n4 52.5823
R27 VP.n11 VP.n10 52.5823
R28 VP.n15 VP.n12 45.6899
R29 VP.n13 VP.n1 20.449
R30 VP.n20 VP.n19 20.449
R31 VP.n4 VP.n3 20.449
R32 VP.n10 VP.n9 20.449
R33 VP.n7 VP.n6 0.189894
R34 VP.n7 VP.n2 0.189894
R35 VP.n12 VP.n2 0.189894
R36 VP.n16 VP.n15 0.189894
R37 VP.n17 VP.n16 0.189894
R38 VP.n17 VP.n0 0.189894
R39 VP.n22 VP.n0 0.189894
R40 VP VP.n22 0.0516364
R41 VTAIL.n11 VTAIL.t2 52.4433
R42 VTAIL.n17 VTAIL.t0 52.4431
R43 VTAIL.n2 VTAIL.t8 52.4431
R44 VTAIL.n16 VTAIL.t16 52.4431
R45 VTAIL.n15 VTAIL.n14 50.6901
R46 VTAIL.n13 VTAIL.n12 50.6901
R47 VTAIL.n10 VTAIL.n9 50.6901
R48 VTAIL.n8 VTAIL.n7 50.6901
R49 VTAIL.n19 VTAIL.n18 50.6899
R50 VTAIL.n1 VTAIL.n0 50.6899
R51 VTAIL.n4 VTAIL.n3 50.6899
R52 VTAIL.n6 VTAIL.n5 50.6899
R53 VTAIL.n8 VTAIL.n6 29.4531
R54 VTAIL.n17 VTAIL.n16 28.9014
R55 VTAIL.n18 VTAIL.t1 1.75374
R56 VTAIL.n18 VTAIL.t6 1.75374
R57 VTAIL.n0 VTAIL.t7 1.75374
R58 VTAIL.n0 VTAIL.t5 1.75374
R59 VTAIL.n3 VTAIL.t15 1.75374
R60 VTAIL.n3 VTAIL.t12 1.75374
R61 VTAIL.n5 VTAIL.t10 1.75374
R62 VTAIL.n5 VTAIL.t14 1.75374
R63 VTAIL.n14 VTAIL.t17 1.75374
R64 VTAIL.n14 VTAIL.t9 1.75374
R65 VTAIL.n12 VTAIL.t11 1.75374
R66 VTAIL.n12 VTAIL.t13 1.75374
R67 VTAIL.n9 VTAIL.t19 1.75374
R68 VTAIL.n9 VTAIL.t3 1.75374
R69 VTAIL.n7 VTAIL.t4 1.75374
R70 VTAIL.n7 VTAIL.t18 1.75374
R71 VTAIL.n13 VTAIL.n11 0.74619
R72 VTAIL.n2 VTAIL.n1 0.74619
R73 VTAIL.n10 VTAIL.n8 0.552224
R74 VTAIL.n11 VTAIL.n10 0.552224
R75 VTAIL.n15 VTAIL.n13 0.552224
R76 VTAIL.n16 VTAIL.n15 0.552224
R77 VTAIL.n6 VTAIL.n4 0.552224
R78 VTAIL.n4 VTAIL.n2 0.552224
R79 VTAIL.n19 VTAIL.n17 0.552224
R80 VTAIL VTAIL.n1 0.472483
R81 VTAIL VTAIL.n19 0.0802414
R82 VDD1.n1 VDD1.t4 69.6738
R83 VDD1.n3 VDD1.t7 69.6737
R84 VDD1.n5 VDD1.n4 67.7271
R85 VDD1.n1 VDD1.n0 67.3689
R86 VDD1.n7 VDD1.n6 67.3687
R87 VDD1.n3 VDD1.n2 67.3686
R88 VDD1.n7 VDD1.n5 43.1776
R89 VDD1.n6 VDD1.t8 1.75374
R90 VDD1.n6 VDD1.t9 1.75374
R91 VDD1.n0 VDD1.t0 1.75374
R92 VDD1.n0 VDD1.t1 1.75374
R93 VDD1.n4 VDD1.t6 1.75374
R94 VDD1.n4 VDD1.t2 1.75374
R95 VDD1.n2 VDD1.t3 1.75374
R96 VDD1.n2 VDD1.t5 1.75374
R97 VDD1 VDD1.n7 0.356103
R98 VDD1 VDD1.n1 0.196621
R99 VDD1.n5 VDD1.n3 0.083085
R100 VN.n9 VN.t7 1583.3
R101 VN.n3 VN.t2 1583.3
R102 VN.n20 VN.t1 1583.3
R103 VN.n14 VN.t3 1583.3
R104 VN.n6 VN.t9 1542.4
R105 VN.n8 VN.t6 1542.4
R106 VN.n2 VN.t8 1542.4
R107 VN.n17 VN.t5 1542.4
R108 VN.n19 VN.t4 1542.4
R109 VN.n13 VN.t0 1542.4
R110 VN.n15 VN.n14 161.489
R111 VN.n4 VN.n3 161.489
R112 VN.n10 VN.n9 161.3
R113 VN.n21 VN.n20 161.3
R114 VN.n18 VN.n11 161.3
R115 VN.n17 VN.n16 161.3
R116 VN.n15 VN.n12 161.3
R117 VN.n7 VN.n0 161.3
R118 VN.n6 VN.n5 161.3
R119 VN.n4 VN.n1 161.3
R120 VN.n6 VN.n1 73.0308
R121 VN.n7 VN.n6 73.0308
R122 VN.n18 VN.n17 73.0308
R123 VN.n17 VN.n12 73.0308
R124 VN.n3 VN.n2 52.5823
R125 VN.n9 VN.n8 52.5823
R126 VN.n20 VN.n19 52.5823
R127 VN.n14 VN.n13 52.5823
R128 VN VN.n21 46.0706
R129 VN.n2 VN.n1 20.449
R130 VN.n8 VN.n7 20.449
R131 VN.n19 VN.n18 20.449
R132 VN.n13 VN.n12 20.449
R133 VN.n21 VN.n11 0.189894
R134 VN.n16 VN.n11 0.189894
R135 VN.n16 VN.n15 0.189894
R136 VN.n5 VN.n4 0.189894
R137 VN.n5 VN.n0 0.189894
R138 VN.n10 VN.n0 0.189894
R139 VN VN.n10 0.0516364
R140 VDD2.n1 VDD2.t7 69.6737
R141 VDD2.n4 VDD2.t8 69.1221
R142 VDD2.n3 VDD2.n2 67.7271
R143 VDD2 VDD2.n7 67.7243
R144 VDD2.n6 VDD2.n5 67.3689
R145 VDD2.n1 VDD2.n0 67.3686
R146 VDD2.n4 VDD2.n3 42.3187
R147 VDD2.n7 VDD2.t9 1.75374
R148 VDD2.n7 VDD2.t6 1.75374
R149 VDD2.n5 VDD2.t5 1.75374
R150 VDD2.n5 VDD2.t4 1.75374
R151 VDD2.n2 VDD2.t3 1.75374
R152 VDD2.n2 VDD2.t2 1.75374
R153 VDD2.n0 VDD2.t1 1.75374
R154 VDD2.n0 VDD2.t0 1.75374
R155 VDD2.n6 VDD2.n4 0.552224
R156 VDD2 VDD2.n6 0.196621
R157 VDD2.n3 VDD2.n1 0.083085
R158 B.n140 B.t9 1656.31
R159 B.n132 B.t0 1656.31
R160 B.n50 B.t6 1656.31
R161 B.n42 B.t3 1656.31
R162 B.n405 B.n404 585
R163 B.n403 B.n102 585
R164 B.n402 B.n401 585
R165 B.n400 B.n103 585
R166 B.n399 B.n398 585
R167 B.n397 B.n104 585
R168 B.n396 B.n395 585
R169 B.n394 B.n105 585
R170 B.n393 B.n392 585
R171 B.n391 B.n106 585
R172 B.n390 B.n389 585
R173 B.n388 B.n107 585
R174 B.n387 B.n386 585
R175 B.n385 B.n108 585
R176 B.n384 B.n383 585
R177 B.n382 B.n109 585
R178 B.n381 B.n380 585
R179 B.n379 B.n110 585
R180 B.n378 B.n377 585
R181 B.n376 B.n111 585
R182 B.n375 B.n374 585
R183 B.n373 B.n112 585
R184 B.n372 B.n371 585
R185 B.n370 B.n113 585
R186 B.n369 B.n368 585
R187 B.n367 B.n114 585
R188 B.n366 B.n365 585
R189 B.n364 B.n115 585
R190 B.n363 B.n362 585
R191 B.n361 B.n116 585
R192 B.n360 B.n359 585
R193 B.n358 B.n117 585
R194 B.n357 B.n356 585
R195 B.n355 B.n118 585
R196 B.n354 B.n353 585
R197 B.n352 B.n119 585
R198 B.n351 B.n350 585
R199 B.n349 B.n120 585
R200 B.n348 B.n347 585
R201 B.n346 B.n121 585
R202 B.n345 B.n344 585
R203 B.n343 B.n122 585
R204 B.n342 B.n341 585
R205 B.n340 B.n123 585
R206 B.n339 B.n338 585
R207 B.n337 B.n124 585
R208 B.n336 B.n335 585
R209 B.n334 B.n125 585
R210 B.n333 B.n332 585
R211 B.n331 B.n126 585
R212 B.n330 B.n329 585
R213 B.n328 B.n127 585
R214 B.n327 B.n326 585
R215 B.n325 B.n128 585
R216 B.n324 B.n323 585
R217 B.n322 B.n129 585
R218 B.n321 B.n320 585
R219 B.n319 B.n130 585
R220 B.n318 B.n317 585
R221 B.n316 B.n131 585
R222 B.n315 B.n314 585
R223 B.n313 B.n312 585
R224 B.n311 B.n135 585
R225 B.n310 B.n309 585
R226 B.n308 B.n136 585
R227 B.n307 B.n306 585
R228 B.n305 B.n137 585
R229 B.n304 B.n303 585
R230 B.n302 B.n138 585
R231 B.n301 B.n300 585
R232 B.n298 B.n139 585
R233 B.n297 B.n296 585
R234 B.n295 B.n142 585
R235 B.n294 B.n293 585
R236 B.n292 B.n143 585
R237 B.n291 B.n290 585
R238 B.n289 B.n144 585
R239 B.n288 B.n287 585
R240 B.n286 B.n145 585
R241 B.n285 B.n284 585
R242 B.n283 B.n146 585
R243 B.n282 B.n281 585
R244 B.n280 B.n147 585
R245 B.n279 B.n278 585
R246 B.n277 B.n148 585
R247 B.n276 B.n275 585
R248 B.n274 B.n149 585
R249 B.n273 B.n272 585
R250 B.n271 B.n150 585
R251 B.n270 B.n269 585
R252 B.n268 B.n151 585
R253 B.n267 B.n266 585
R254 B.n265 B.n152 585
R255 B.n264 B.n263 585
R256 B.n262 B.n153 585
R257 B.n261 B.n260 585
R258 B.n259 B.n154 585
R259 B.n258 B.n257 585
R260 B.n256 B.n155 585
R261 B.n255 B.n254 585
R262 B.n253 B.n156 585
R263 B.n252 B.n251 585
R264 B.n250 B.n157 585
R265 B.n249 B.n248 585
R266 B.n247 B.n158 585
R267 B.n246 B.n245 585
R268 B.n244 B.n159 585
R269 B.n243 B.n242 585
R270 B.n241 B.n160 585
R271 B.n240 B.n239 585
R272 B.n238 B.n161 585
R273 B.n237 B.n236 585
R274 B.n235 B.n162 585
R275 B.n234 B.n233 585
R276 B.n232 B.n163 585
R277 B.n231 B.n230 585
R278 B.n229 B.n164 585
R279 B.n228 B.n227 585
R280 B.n226 B.n165 585
R281 B.n225 B.n224 585
R282 B.n223 B.n166 585
R283 B.n222 B.n221 585
R284 B.n220 B.n167 585
R285 B.n219 B.n218 585
R286 B.n217 B.n168 585
R287 B.n216 B.n215 585
R288 B.n214 B.n169 585
R289 B.n213 B.n212 585
R290 B.n211 B.n170 585
R291 B.n210 B.n209 585
R292 B.n208 B.n171 585
R293 B.n406 B.n101 585
R294 B.n408 B.n407 585
R295 B.n409 B.n100 585
R296 B.n411 B.n410 585
R297 B.n412 B.n99 585
R298 B.n414 B.n413 585
R299 B.n415 B.n98 585
R300 B.n417 B.n416 585
R301 B.n418 B.n97 585
R302 B.n420 B.n419 585
R303 B.n421 B.n96 585
R304 B.n423 B.n422 585
R305 B.n424 B.n95 585
R306 B.n426 B.n425 585
R307 B.n427 B.n94 585
R308 B.n429 B.n428 585
R309 B.n430 B.n93 585
R310 B.n432 B.n431 585
R311 B.n433 B.n92 585
R312 B.n435 B.n434 585
R313 B.n436 B.n91 585
R314 B.n438 B.n437 585
R315 B.n439 B.n90 585
R316 B.n441 B.n440 585
R317 B.n442 B.n89 585
R318 B.n444 B.n443 585
R319 B.n445 B.n88 585
R320 B.n447 B.n446 585
R321 B.n448 B.n87 585
R322 B.n450 B.n449 585
R323 B.n451 B.n86 585
R324 B.n453 B.n452 585
R325 B.n454 B.n85 585
R326 B.n456 B.n455 585
R327 B.n457 B.n84 585
R328 B.n459 B.n458 585
R329 B.n460 B.n83 585
R330 B.n462 B.n461 585
R331 B.n463 B.n82 585
R332 B.n465 B.n464 585
R333 B.n663 B.n662 585
R334 B.n661 B.n12 585
R335 B.n660 B.n659 585
R336 B.n658 B.n13 585
R337 B.n657 B.n656 585
R338 B.n655 B.n14 585
R339 B.n654 B.n653 585
R340 B.n652 B.n15 585
R341 B.n651 B.n650 585
R342 B.n649 B.n16 585
R343 B.n648 B.n647 585
R344 B.n646 B.n17 585
R345 B.n645 B.n644 585
R346 B.n643 B.n18 585
R347 B.n642 B.n641 585
R348 B.n640 B.n19 585
R349 B.n639 B.n638 585
R350 B.n637 B.n20 585
R351 B.n636 B.n635 585
R352 B.n634 B.n21 585
R353 B.n633 B.n632 585
R354 B.n631 B.n22 585
R355 B.n630 B.n629 585
R356 B.n628 B.n23 585
R357 B.n627 B.n626 585
R358 B.n625 B.n24 585
R359 B.n624 B.n623 585
R360 B.n622 B.n25 585
R361 B.n621 B.n620 585
R362 B.n619 B.n26 585
R363 B.n618 B.n617 585
R364 B.n616 B.n27 585
R365 B.n615 B.n614 585
R366 B.n613 B.n28 585
R367 B.n612 B.n611 585
R368 B.n610 B.n29 585
R369 B.n609 B.n608 585
R370 B.n607 B.n30 585
R371 B.n606 B.n605 585
R372 B.n604 B.n31 585
R373 B.n603 B.n602 585
R374 B.n601 B.n32 585
R375 B.n600 B.n599 585
R376 B.n598 B.n33 585
R377 B.n597 B.n596 585
R378 B.n595 B.n34 585
R379 B.n594 B.n593 585
R380 B.n592 B.n35 585
R381 B.n591 B.n590 585
R382 B.n589 B.n36 585
R383 B.n588 B.n587 585
R384 B.n586 B.n37 585
R385 B.n585 B.n584 585
R386 B.n583 B.n38 585
R387 B.n582 B.n581 585
R388 B.n580 B.n39 585
R389 B.n579 B.n578 585
R390 B.n577 B.n40 585
R391 B.n576 B.n575 585
R392 B.n574 B.n41 585
R393 B.n573 B.n572 585
R394 B.n571 B.n570 585
R395 B.n569 B.n45 585
R396 B.n568 B.n567 585
R397 B.n566 B.n46 585
R398 B.n565 B.n564 585
R399 B.n563 B.n47 585
R400 B.n562 B.n561 585
R401 B.n560 B.n48 585
R402 B.n559 B.n558 585
R403 B.n556 B.n49 585
R404 B.n555 B.n554 585
R405 B.n553 B.n52 585
R406 B.n552 B.n551 585
R407 B.n550 B.n53 585
R408 B.n549 B.n548 585
R409 B.n547 B.n54 585
R410 B.n546 B.n545 585
R411 B.n544 B.n55 585
R412 B.n543 B.n542 585
R413 B.n541 B.n56 585
R414 B.n540 B.n539 585
R415 B.n538 B.n57 585
R416 B.n537 B.n536 585
R417 B.n535 B.n58 585
R418 B.n534 B.n533 585
R419 B.n532 B.n59 585
R420 B.n531 B.n530 585
R421 B.n529 B.n60 585
R422 B.n528 B.n527 585
R423 B.n526 B.n61 585
R424 B.n525 B.n524 585
R425 B.n523 B.n62 585
R426 B.n522 B.n521 585
R427 B.n520 B.n63 585
R428 B.n519 B.n518 585
R429 B.n517 B.n64 585
R430 B.n516 B.n515 585
R431 B.n514 B.n65 585
R432 B.n513 B.n512 585
R433 B.n511 B.n66 585
R434 B.n510 B.n509 585
R435 B.n508 B.n67 585
R436 B.n507 B.n506 585
R437 B.n505 B.n68 585
R438 B.n504 B.n503 585
R439 B.n502 B.n69 585
R440 B.n501 B.n500 585
R441 B.n499 B.n70 585
R442 B.n498 B.n497 585
R443 B.n496 B.n71 585
R444 B.n495 B.n494 585
R445 B.n493 B.n72 585
R446 B.n492 B.n491 585
R447 B.n490 B.n73 585
R448 B.n489 B.n488 585
R449 B.n487 B.n74 585
R450 B.n486 B.n485 585
R451 B.n484 B.n75 585
R452 B.n483 B.n482 585
R453 B.n481 B.n76 585
R454 B.n480 B.n479 585
R455 B.n478 B.n77 585
R456 B.n477 B.n476 585
R457 B.n475 B.n78 585
R458 B.n474 B.n473 585
R459 B.n472 B.n79 585
R460 B.n471 B.n470 585
R461 B.n469 B.n80 585
R462 B.n468 B.n467 585
R463 B.n466 B.n81 585
R464 B.n664 B.n11 585
R465 B.n666 B.n665 585
R466 B.n667 B.n10 585
R467 B.n669 B.n668 585
R468 B.n670 B.n9 585
R469 B.n672 B.n671 585
R470 B.n673 B.n8 585
R471 B.n675 B.n674 585
R472 B.n676 B.n7 585
R473 B.n678 B.n677 585
R474 B.n679 B.n6 585
R475 B.n681 B.n680 585
R476 B.n682 B.n5 585
R477 B.n684 B.n683 585
R478 B.n685 B.n4 585
R479 B.n687 B.n686 585
R480 B.n688 B.n3 585
R481 B.n690 B.n689 585
R482 B.n691 B.n0 585
R483 B.n2 B.n1 585
R484 B.n181 B.n180 585
R485 B.n183 B.n182 585
R486 B.n184 B.n179 585
R487 B.n186 B.n185 585
R488 B.n187 B.n178 585
R489 B.n189 B.n188 585
R490 B.n190 B.n177 585
R491 B.n192 B.n191 585
R492 B.n193 B.n176 585
R493 B.n195 B.n194 585
R494 B.n196 B.n175 585
R495 B.n198 B.n197 585
R496 B.n199 B.n174 585
R497 B.n201 B.n200 585
R498 B.n202 B.n173 585
R499 B.n204 B.n203 585
R500 B.n205 B.n172 585
R501 B.n207 B.n206 585
R502 B.n206 B.n171 506.916
R503 B.n404 B.n101 506.916
R504 B.n464 B.n81 506.916
R505 B.n662 B.n11 506.916
R506 B.n693 B.n692 256.663
R507 B.n692 B.n691 235.042
R508 B.n692 B.n2 235.042
R509 B.n210 B.n171 163.367
R510 B.n211 B.n210 163.367
R511 B.n212 B.n211 163.367
R512 B.n212 B.n169 163.367
R513 B.n216 B.n169 163.367
R514 B.n217 B.n216 163.367
R515 B.n218 B.n217 163.367
R516 B.n218 B.n167 163.367
R517 B.n222 B.n167 163.367
R518 B.n223 B.n222 163.367
R519 B.n224 B.n223 163.367
R520 B.n224 B.n165 163.367
R521 B.n228 B.n165 163.367
R522 B.n229 B.n228 163.367
R523 B.n230 B.n229 163.367
R524 B.n230 B.n163 163.367
R525 B.n234 B.n163 163.367
R526 B.n235 B.n234 163.367
R527 B.n236 B.n235 163.367
R528 B.n236 B.n161 163.367
R529 B.n240 B.n161 163.367
R530 B.n241 B.n240 163.367
R531 B.n242 B.n241 163.367
R532 B.n242 B.n159 163.367
R533 B.n246 B.n159 163.367
R534 B.n247 B.n246 163.367
R535 B.n248 B.n247 163.367
R536 B.n248 B.n157 163.367
R537 B.n252 B.n157 163.367
R538 B.n253 B.n252 163.367
R539 B.n254 B.n253 163.367
R540 B.n254 B.n155 163.367
R541 B.n258 B.n155 163.367
R542 B.n259 B.n258 163.367
R543 B.n260 B.n259 163.367
R544 B.n260 B.n153 163.367
R545 B.n264 B.n153 163.367
R546 B.n265 B.n264 163.367
R547 B.n266 B.n265 163.367
R548 B.n266 B.n151 163.367
R549 B.n270 B.n151 163.367
R550 B.n271 B.n270 163.367
R551 B.n272 B.n271 163.367
R552 B.n272 B.n149 163.367
R553 B.n276 B.n149 163.367
R554 B.n277 B.n276 163.367
R555 B.n278 B.n277 163.367
R556 B.n278 B.n147 163.367
R557 B.n282 B.n147 163.367
R558 B.n283 B.n282 163.367
R559 B.n284 B.n283 163.367
R560 B.n284 B.n145 163.367
R561 B.n288 B.n145 163.367
R562 B.n289 B.n288 163.367
R563 B.n290 B.n289 163.367
R564 B.n290 B.n143 163.367
R565 B.n294 B.n143 163.367
R566 B.n295 B.n294 163.367
R567 B.n296 B.n295 163.367
R568 B.n296 B.n139 163.367
R569 B.n301 B.n139 163.367
R570 B.n302 B.n301 163.367
R571 B.n303 B.n302 163.367
R572 B.n303 B.n137 163.367
R573 B.n307 B.n137 163.367
R574 B.n308 B.n307 163.367
R575 B.n309 B.n308 163.367
R576 B.n309 B.n135 163.367
R577 B.n313 B.n135 163.367
R578 B.n314 B.n313 163.367
R579 B.n314 B.n131 163.367
R580 B.n318 B.n131 163.367
R581 B.n319 B.n318 163.367
R582 B.n320 B.n319 163.367
R583 B.n320 B.n129 163.367
R584 B.n324 B.n129 163.367
R585 B.n325 B.n324 163.367
R586 B.n326 B.n325 163.367
R587 B.n326 B.n127 163.367
R588 B.n330 B.n127 163.367
R589 B.n331 B.n330 163.367
R590 B.n332 B.n331 163.367
R591 B.n332 B.n125 163.367
R592 B.n336 B.n125 163.367
R593 B.n337 B.n336 163.367
R594 B.n338 B.n337 163.367
R595 B.n338 B.n123 163.367
R596 B.n342 B.n123 163.367
R597 B.n343 B.n342 163.367
R598 B.n344 B.n343 163.367
R599 B.n344 B.n121 163.367
R600 B.n348 B.n121 163.367
R601 B.n349 B.n348 163.367
R602 B.n350 B.n349 163.367
R603 B.n350 B.n119 163.367
R604 B.n354 B.n119 163.367
R605 B.n355 B.n354 163.367
R606 B.n356 B.n355 163.367
R607 B.n356 B.n117 163.367
R608 B.n360 B.n117 163.367
R609 B.n361 B.n360 163.367
R610 B.n362 B.n361 163.367
R611 B.n362 B.n115 163.367
R612 B.n366 B.n115 163.367
R613 B.n367 B.n366 163.367
R614 B.n368 B.n367 163.367
R615 B.n368 B.n113 163.367
R616 B.n372 B.n113 163.367
R617 B.n373 B.n372 163.367
R618 B.n374 B.n373 163.367
R619 B.n374 B.n111 163.367
R620 B.n378 B.n111 163.367
R621 B.n379 B.n378 163.367
R622 B.n380 B.n379 163.367
R623 B.n380 B.n109 163.367
R624 B.n384 B.n109 163.367
R625 B.n385 B.n384 163.367
R626 B.n386 B.n385 163.367
R627 B.n386 B.n107 163.367
R628 B.n390 B.n107 163.367
R629 B.n391 B.n390 163.367
R630 B.n392 B.n391 163.367
R631 B.n392 B.n105 163.367
R632 B.n396 B.n105 163.367
R633 B.n397 B.n396 163.367
R634 B.n398 B.n397 163.367
R635 B.n398 B.n103 163.367
R636 B.n402 B.n103 163.367
R637 B.n403 B.n402 163.367
R638 B.n404 B.n403 163.367
R639 B.n464 B.n463 163.367
R640 B.n463 B.n462 163.367
R641 B.n462 B.n83 163.367
R642 B.n458 B.n83 163.367
R643 B.n458 B.n457 163.367
R644 B.n457 B.n456 163.367
R645 B.n456 B.n85 163.367
R646 B.n452 B.n85 163.367
R647 B.n452 B.n451 163.367
R648 B.n451 B.n450 163.367
R649 B.n450 B.n87 163.367
R650 B.n446 B.n87 163.367
R651 B.n446 B.n445 163.367
R652 B.n445 B.n444 163.367
R653 B.n444 B.n89 163.367
R654 B.n440 B.n89 163.367
R655 B.n440 B.n439 163.367
R656 B.n439 B.n438 163.367
R657 B.n438 B.n91 163.367
R658 B.n434 B.n91 163.367
R659 B.n434 B.n433 163.367
R660 B.n433 B.n432 163.367
R661 B.n432 B.n93 163.367
R662 B.n428 B.n93 163.367
R663 B.n428 B.n427 163.367
R664 B.n427 B.n426 163.367
R665 B.n426 B.n95 163.367
R666 B.n422 B.n95 163.367
R667 B.n422 B.n421 163.367
R668 B.n421 B.n420 163.367
R669 B.n420 B.n97 163.367
R670 B.n416 B.n97 163.367
R671 B.n416 B.n415 163.367
R672 B.n415 B.n414 163.367
R673 B.n414 B.n99 163.367
R674 B.n410 B.n99 163.367
R675 B.n410 B.n409 163.367
R676 B.n409 B.n408 163.367
R677 B.n408 B.n101 163.367
R678 B.n662 B.n661 163.367
R679 B.n661 B.n660 163.367
R680 B.n660 B.n13 163.367
R681 B.n656 B.n13 163.367
R682 B.n656 B.n655 163.367
R683 B.n655 B.n654 163.367
R684 B.n654 B.n15 163.367
R685 B.n650 B.n15 163.367
R686 B.n650 B.n649 163.367
R687 B.n649 B.n648 163.367
R688 B.n648 B.n17 163.367
R689 B.n644 B.n17 163.367
R690 B.n644 B.n643 163.367
R691 B.n643 B.n642 163.367
R692 B.n642 B.n19 163.367
R693 B.n638 B.n19 163.367
R694 B.n638 B.n637 163.367
R695 B.n637 B.n636 163.367
R696 B.n636 B.n21 163.367
R697 B.n632 B.n21 163.367
R698 B.n632 B.n631 163.367
R699 B.n631 B.n630 163.367
R700 B.n630 B.n23 163.367
R701 B.n626 B.n23 163.367
R702 B.n626 B.n625 163.367
R703 B.n625 B.n624 163.367
R704 B.n624 B.n25 163.367
R705 B.n620 B.n25 163.367
R706 B.n620 B.n619 163.367
R707 B.n619 B.n618 163.367
R708 B.n618 B.n27 163.367
R709 B.n614 B.n27 163.367
R710 B.n614 B.n613 163.367
R711 B.n613 B.n612 163.367
R712 B.n612 B.n29 163.367
R713 B.n608 B.n29 163.367
R714 B.n608 B.n607 163.367
R715 B.n607 B.n606 163.367
R716 B.n606 B.n31 163.367
R717 B.n602 B.n31 163.367
R718 B.n602 B.n601 163.367
R719 B.n601 B.n600 163.367
R720 B.n600 B.n33 163.367
R721 B.n596 B.n33 163.367
R722 B.n596 B.n595 163.367
R723 B.n595 B.n594 163.367
R724 B.n594 B.n35 163.367
R725 B.n590 B.n35 163.367
R726 B.n590 B.n589 163.367
R727 B.n589 B.n588 163.367
R728 B.n588 B.n37 163.367
R729 B.n584 B.n37 163.367
R730 B.n584 B.n583 163.367
R731 B.n583 B.n582 163.367
R732 B.n582 B.n39 163.367
R733 B.n578 B.n39 163.367
R734 B.n578 B.n577 163.367
R735 B.n577 B.n576 163.367
R736 B.n576 B.n41 163.367
R737 B.n572 B.n41 163.367
R738 B.n572 B.n571 163.367
R739 B.n571 B.n45 163.367
R740 B.n567 B.n45 163.367
R741 B.n567 B.n566 163.367
R742 B.n566 B.n565 163.367
R743 B.n565 B.n47 163.367
R744 B.n561 B.n47 163.367
R745 B.n561 B.n560 163.367
R746 B.n560 B.n559 163.367
R747 B.n559 B.n49 163.367
R748 B.n554 B.n49 163.367
R749 B.n554 B.n553 163.367
R750 B.n553 B.n552 163.367
R751 B.n552 B.n53 163.367
R752 B.n548 B.n53 163.367
R753 B.n548 B.n547 163.367
R754 B.n547 B.n546 163.367
R755 B.n546 B.n55 163.367
R756 B.n542 B.n55 163.367
R757 B.n542 B.n541 163.367
R758 B.n541 B.n540 163.367
R759 B.n540 B.n57 163.367
R760 B.n536 B.n57 163.367
R761 B.n536 B.n535 163.367
R762 B.n535 B.n534 163.367
R763 B.n534 B.n59 163.367
R764 B.n530 B.n59 163.367
R765 B.n530 B.n529 163.367
R766 B.n529 B.n528 163.367
R767 B.n528 B.n61 163.367
R768 B.n524 B.n61 163.367
R769 B.n524 B.n523 163.367
R770 B.n523 B.n522 163.367
R771 B.n522 B.n63 163.367
R772 B.n518 B.n63 163.367
R773 B.n518 B.n517 163.367
R774 B.n517 B.n516 163.367
R775 B.n516 B.n65 163.367
R776 B.n512 B.n65 163.367
R777 B.n512 B.n511 163.367
R778 B.n511 B.n510 163.367
R779 B.n510 B.n67 163.367
R780 B.n506 B.n67 163.367
R781 B.n506 B.n505 163.367
R782 B.n505 B.n504 163.367
R783 B.n504 B.n69 163.367
R784 B.n500 B.n69 163.367
R785 B.n500 B.n499 163.367
R786 B.n499 B.n498 163.367
R787 B.n498 B.n71 163.367
R788 B.n494 B.n71 163.367
R789 B.n494 B.n493 163.367
R790 B.n493 B.n492 163.367
R791 B.n492 B.n73 163.367
R792 B.n488 B.n73 163.367
R793 B.n488 B.n487 163.367
R794 B.n487 B.n486 163.367
R795 B.n486 B.n75 163.367
R796 B.n482 B.n75 163.367
R797 B.n482 B.n481 163.367
R798 B.n481 B.n480 163.367
R799 B.n480 B.n77 163.367
R800 B.n476 B.n77 163.367
R801 B.n476 B.n475 163.367
R802 B.n475 B.n474 163.367
R803 B.n474 B.n79 163.367
R804 B.n470 B.n79 163.367
R805 B.n470 B.n469 163.367
R806 B.n469 B.n468 163.367
R807 B.n468 B.n81 163.367
R808 B.n666 B.n11 163.367
R809 B.n667 B.n666 163.367
R810 B.n668 B.n667 163.367
R811 B.n668 B.n9 163.367
R812 B.n672 B.n9 163.367
R813 B.n673 B.n672 163.367
R814 B.n674 B.n673 163.367
R815 B.n674 B.n7 163.367
R816 B.n678 B.n7 163.367
R817 B.n679 B.n678 163.367
R818 B.n680 B.n679 163.367
R819 B.n680 B.n5 163.367
R820 B.n684 B.n5 163.367
R821 B.n685 B.n684 163.367
R822 B.n686 B.n685 163.367
R823 B.n686 B.n3 163.367
R824 B.n690 B.n3 163.367
R825 B.n691 B.n690 163.367
R826 B.n181 B.n2 163.367
R827 B.n182 B.n181 163.367
R828 B.n182 B.n179 163.367
R829 B.n186 B.n179 163.367
R830 B.n187 B.n186 163.367
R831 B.n188 B.n187 163.367
R832 B.n188 B.n177 163.367
R833 B.n192 B.n177 163.367
R834 B.n193 B.n192 163.367
R835 B.n194 B.n193 163.367
R836 B.n194 B.n175 163.367
R837 B.n198 B.n175 163.367
R838 B.n199 B.n198 163.367
R839 B.n200 B.n199 163.367
R840 B.n200 B.n173 163.367
R841 B.n204 B.n173 163.367
R842 B.n205 B.n204 163.367
R843 B.n206 B.n205 163.367
R844 B.n132 B.t1 122.055
R845 B.n50 B.t8 122.055
R846 B.n140 B.t10 122.031
R847 B.n42 B.t5 122.031
R848 B.n133 B.t2 109.644
R849 B.n51 B.t7 109.644
R850 B.n141 B.t11 109.62
R851 B.n43 B.t4 109.62
R852 B.n299 B.n141 59.5399
R853 B.n134 B.n133 59.5399
R854 B.n557 B.n51 59.5399
R855 B.n44 B.n43 59.5399
R856 B.n664 B.n663 32.9371
R857 B.n466 B.n465 32.9371
R858 B.n406 B.n405 32.9371
R859 B.n208 B.n207 32.9371
R860 B B.n693 18.0485
R861 B.n141 B.n140 12.4126
R862 B.n133 B.n132 12.4126
R863 B.n51 B.n50 12.4126
R864 B.n43 B.n42 12.4126
R865 B.n665 B.n664 10.6151
R866 B.n665 B.n10 10.6151
R867 B.n669 B.n10 10.6151
R868 B.n670 B.n669 10.6151
R869 B.n671 B.n670 10.6151
R870 B.n671 B.n8 10.6151
R871 B.n675 B.n8 10.6151
R872 B.n676 B.n675 10.6151
R873 B.n677 B.n676 10.6151
R874 B.n677 B.n6 10.6151
R875 B.n681 B.n6 10.6151
R876 B.n682 B.n681 10.6151
R877 B.n683 B.n682 10.6151
R878 B.n683 B.n4 10.6151
R879 B.n687 B.n4 10.6151
R880 B.n688 B.n687 10.6151
R881 B.n689 B.n688 10.6151
R882 B.n689 B.n0 10.6151
R883 B.n663 B.n12 10.6151
R884 B.n659 B.n12 10.6151
R885 B.n659 B.n658 10.6151
R886 B.n658 B.n657 10.6151
R887 B.n657 B.n14 10.6151
R888 B.n653 B.n14 10.6151
R889 B.n653 B.n652 10.6151
R890 B.n652 B.n651 10.6151
R891 B.n651 B.n16 10.6151
R892 B.n647 B.n16 10.6151
R893 B.n647 B.n646 10.6151
R894 B.n646 B.n645 10.6151
R895 B.n645 B.n18 10.6151
R896 B.n641 B.n18 10.6151
R897 B.n641 B.n640 10.6151
R898 B.n640 B.n639 10.6151
R899 B.n639 B.n20 10.6151
R900 B.n635 B.n20 10.6151
R901 B.n635 B.n634 10.6151
R902 B.n634 B.n633 10.6151
R903 B.n633 B.n22 10.6151
R904 B.n629 B.n22 10.6151
R905 B.n629 B.n628 10.6151
R906 B.n628 B.n627 10.6151
R907 B.n627 B.n24 10.6151
R908 B.n623 B.n24 10.6151
R909 B.n623 B.n622 10.6151
R910 B.n622 B.n621 10.6151
R911 B.n621 B.n26 10.6151
R912 B.n617 B.n26 10.6151
R913 B.n617 B.n616 10.6151
R914 B.n616 B.n615 10.6151
R915 B.n615 B.n28 10.6151
R916 B.n611 B.n28 10.6151
R917 B.n611 B.n610 10.6151
R918 B.n610 B.n609 10.6151
R919 B.n609 B.n30 10.6151
R920 B.n605 B.n30 10.6151
R921 B.n605 B.n604 10.6151
R922 B.n604 B.n603 10.6151
R923 B.n603 B.n32 10.6151
R924 B.n599 B.n32 10.6151
R925 B.n599 B.n598 10.6151
R926 B.n598 B.n597 10.6151
R927 B.n597 B.n34 10.6151
R928 B.n593 B.n34 10.6151
R929 B.n593 B.n592 10.6151
R930 B.n592 B.n591 10.6151
R931 B.n591 B.n36 10.6151
R932 B.n587 B.n36 10.6151
R933 B.n587 B.n586 10.6151
R934 B.n586 B.n585 10.6151
R935 B.n585 B.n38 10.6151
R936 B.n581 B.n38 10.6151
R937 B.n581 B.n580 10.6151
R938 B.n580 B.n579 10.6151
R939 B.n579 B.n40 10.6151
R940 B.n575 B.n40 10.6151
R941 B.n575 B.n574 10.6151
R942 B.n574 B.n573 10.6151
R943 B.n570 B.n569 10.6151
R944 B.n569 B.n568 10.6151
R945 B.n568 B.n46 10.6151
R946 B.n564 B.n46 10.6151
R947 B.n564 B.n563 10.6151
R948 B.n563 B.n562 10.6151
R949 B.n562 B.n48 10.6151
R950 B.n558 B.n48 10.6151
R951 B.n556 B.n555 10.6151
R952 B.n555 B.n52 10.6151
R953 B.n551 B.n52 10.6151
R954 B.n551 B.n550 10.6151
R955 B.n550 B.n549 10.6151
R956 B.n549 B.n54 10.6151
R957 B.n545 B.n54 10.6151
R958 B.n545 B.n544 10.6151
R959 B.n544 B.n543 10.6151
R960 B.n543 B.n56 10.6151
R961 B.n539 B.n56 10.6151
R962 B.n539 B.n538 10.6151
R963 B.n538 B.n537 10.6151
R964 B.n537 B.n58 10.6151
R965 B.n533 B.n58 10.6151
R966 B.n533 B.n532 10.6151
R967 B.n532 B.n531 10.6151
R968 B.n531 B.n60 10.6151
R969 B.n527 B.n60 10.6151
R970 B.n527 B.n526 10.6151
R971 B.n526 B.n525 10.6151
R972 B.n525 B.n62 10.6151
R973 B.n521 B.n62 10.6151
R974 B.n521 B.n520 10.6151
R975 B.n520 B.n519 10.6151
R976 B.n519 B.n64 10.6151
R977 B.n515 B.n64 10.6151
R978 B.n515 B.n514 10.6151
R979 B.n514 B.n513 10.6151
R980 B.n513 B.n66 10.6151
R981 B.n509 B.n66 10.6151
R982 B.n509 B.n508 10.6151
R983 B.n508 B.n507 10.6151
R984 B.n507 B.n68 10.6151
R985 B.n503 B.n68 10.6151
R986 B.n503 B.n502 10.6151
R987 B.n502 B.n501 10.6151
R988 B.n501 B.n70 10.6151
R989 B.n497 B.n70 10.6151
R990 B.n497 B.n496 10.6151
R991 B.n496 B.n495 10.6151
R992 B.n495 B.n72 10.6151
R993 B.n491 B.n72 10.6151
R994 B.n491 B.n490 10.6151
R995 B.n490 B.n489 10.6151
R996 B.n489 B.n74 10.6151
R997 B.n485 B.n74 10.6151
R998 B.n485 B.n484 10.6151
R999 B.n484 B.n483 10.6151
R1000 B.n483 B.n76 10.6151
R1001 B.n479 B.n76 10.6151
R1002 B.n479 B.n478 10.6151
R1003 B.n478 B.n477 10.6151
R1004 B.n477 B.n78 10.6151
R1005 B.n473 B.n78 10.6151
R1006 B.n473 B.n472 10.6151
R1007 B.n472 B.n471 10.6151
R1008 B.n471 B.n80 10.6151
R1009 B.n467 B.n80 10.6151
R1010 B.n467 B.n466 10.6151
R1011 B.n465 B.n82 10.6151
R1012 B.n461 B.n82 10.6151
R1013 B.n461 B.n460 10.6151
R1014 B.n460 B.n459 10.6151
R1015 B.n459 B.n84 10.6151
R1016 B.n455 B.n84 10.6151
R1017 B.n455 B.n454 10.6151
R1018 B.n454 B.n453 10.6151
R1019 B.n453 B.n86 10.6151
R1020 B.n449 B.n86 10.6151
R1021 B.n449 B.n448 10.6151
R1022 B.n448 B.n447 10.6151
R1023 B.n447 B.n88 10.6151
R1024 B.n443 B.n88 10.6151
R1025 B.n443 B.n442 10.6151
R1026 B.n442 B.n441 10.6151
R1027 B.n441 B.n90 10.6151
R1028 B.n437 B.n90 10.6151
R1029 B.n437 B.n436 10.6151
R1030 B.n436 B.n435 10.6151
R1031 B.n435 B.n92 10.6151
R1032 B.n431 B.n92 10.6151
R1033 B.n431 B.n430 10.6151
R1034 B.n430 B.n429 10.6151
R1035 B.n429 B.n94 10.6151
R1036 B.n425 B.n94 10.6151
R1037 B.n425 B.n424 10.6151
R1038 B.n424 B.n423 10.6151
R1039 B.n423 B.n96 10.6151
R1040 B.n419 B.n96 10.6151
R1041 B.n419 B.n418 10.6151
R1042 B.n418 B.n417 10.6151
R1043 B.n417 B.n98 10.6151
R1044 B.n413 B.n98 10.6151
R1045 B.n413 B.n412 10.6151
R1046 B.n412 B.n411 10.6151
R1047 B.n411 B.n100 10.6151
R1048 B.n407 B.n100 10.6151
R1049 B.n407 B.n406 10.6151
R1050 B.n180 B.n1 10.6151
R1051 B.n183 B.n180 10.6151
R1052 B.n184 B.n183 10.6151
R1053 B.n185 B.n184 10.6151
R1054 B.n185 B.n178 10.6151
R1055 B.n189 B.n178 10.6151
R1056 B.n190 B.n189 10.6151
R1057 B.n191 B.n190 10.6151
R1058 B.n191 B.n176 10.6151
R1059 B.n195 B.n176 10.6151
R1060 B.n196 B.n195 10.6151
R1061 B.n197 B.n196 10.6151
R1062 B.n197 B.n174 10.6151
R1063 B.n201 B.n174 10.6151
R1064 B.n202 B.n201 10.6151
R1065 B.n203 B.n202 10.6151
R1066 B.n203 B.n172 10.6151
R1067 B.n207 B.n172 10.6151
R1068 B.n209 B.n208 10.6151
R1069 B.n209 B.n170 10.6151
R1070 B.n213 B.n170 10.6151
R1071 B.n214 B.n213 10.6151
R1072 B.n215 B.n214 10.6151
R1073 B.n215 B.n168 10.6151
R1074 B.n219 B.n168 10.6151
R1075 B.n220 B.n219 10.6151
R1076 B.n221 B.n220 10.6151
R1077 B.n221 B.n166 10.6151
R1078 B.n225 B.n166 10.6151
R1079 B.n226 B.n225 10.6151
R1080 B.n227 B.n226 10.6151
R1081 B.n227 B.n164 10.6151
R1082 B.n231 B.n164 10.6151
R1083 B.n232 B.n231 10.6151
R1084 B.n233 B.n232 10.6151
R1085 B.n233 B.n162 10.6151
R1086 B.n237 B.n162 10.6151
R1087 B.n238 B.n237 10.6151
R1088 B.n239 B.n238 10.6151
R1089 B.n239 B.n160 10.6151
R1090 B.n243 B.n160 10.6151
R1091 B.n244 B.n243 10.6151
R1092 B.n245 B.n244 10.6151
R1093 B.n245 B.n158 10.6151
R1094 B.n249 B.n158 10.6151
R1095 B.n250 B.n249 10.6151
R1096 B.n251 B.n250 10.6151
R1097 B.n251 B.n156 10.6151
R1098 B.n255 B.n156 10.6151
R1099 B.n256 B.n255 10.6151
R1100 B.n257 B.n256 10.6151
R1101 B.n257 B.n154 10.6151
R1102 B.n261 B.n154 10.6151
R1103 B.n262 B.n261 10.6151
R1104 B.n263 B.n262 10.6151
R1105 B.n263 B.n152 10.6151
R1106 B.n267 B.n152 10.6151
R1107 B.n268 B.n267 10.6151
R1108 B.n269 B.n268 10.6151
R1109 B.n269 B.n150 10.6151
R1110 B.n273 B.n150 10.6151
R1111 B.n274 B.n273 10.6151
R1112 B.n275 B.n274 10.6151
R1113 B.n275 B.n148 10.6151
R1114 B.n279 B.n148 10.6151
R1115 B.n280 B.n279 10.6151
R1116 B.n281 B.n280 10.6151
R1117 B.n281 B.n146 10.6151
R1118 B.n285 B.n146 10.6151
R1119 B.n286 B.n285 10.6151
R1120 B.n287 B.n286 10.6151
R1121 B.n287 B.n144 10.6151
R1122 B.n291 B.n144 10.6151
R1123 B.n292 B.n291 10.6151
R1124 B.n293 B.n292 10.6151
R1125 B.n293 B.n142 10.6151
R1126 B.n297 B.n142 10.6151
R1127 B.n298 B.n297 10.6151
R1128 B.n300 B.n138 10.6151
R1129 B.n304 B.n138 10.6151
R1130 B.n305 B.n304 10.6151
R1131 B.n306 B.n305 10.6151
R1132 B.n306 B.n136 10.6151
R1133 B.n310 B.n136 10.6151
R1134 B.n311 B.n310 10.6151
R1135 B.n312 B.n311 10.6151
R1136 B.n316 B.n315 10.6151
R1137 B.n317 B.n316 10.6151
R1138 B.n317 B.n130 10.6151
R1139 B.n321 B.n130 10.6151
R1140 B.n322 B.n321 10.6151
R1141 B.n323 B.n322 10.6151
R1142 B.n323 B.n128 10.6151
R1143 B.n327 B.n128 10.6151
R1144 B.n328 B.n327 10.6151
R1145 B.n329 B.n328 10.6151
R1146 B.n329 B.n126 10.6151
R1147 B.n333 B.n126 10.6151
R1148 B.n334 B.n333 10.6151
R1149 B.n335 B.n334 10.6151
R1150 B.n335 B.n124 10.6151
R1151 B.n339 B.n124 10.6151
R1152 B.n340 B.n339 10.6151
R1153 B.n341 B.n340 10.6151
R1154 B.n341 B.n122 10.6151
R1155 B.n345 B.n122 10.6151
R1156 B.n346 B.n345 10.6151
R1157 B.n347 B.n346 10.6151
R1158 B.n347 B.n120 10.6151
R1159 B.n351 B.n120 10.6151
R1160 B.n352 B.n351 10.6151
R1161 B.n353 B.n352 10.6151
R1162 B.n353 B.n118 10.6151
R1163 B.n357 B.n118 10.6151
R1164 B.n358 B.n357 10.6151
R1165 B.n359 B.n358 10.6151
R1166 B.n359 B.n116 10.6151
R1167 B.n363 B.n116 10.6151
R1168 B.n364 B.n363 10.6151
R1169 B.n365 B.n364 10.6151
R1170 B.n365 B.n114 10.6151
R1171 B.n369 B.n114 10.6151
R1172 B.n370 B.n369 10.6151
R1173 B.n371 B.n370 10.6151
R1174 B.n371 B.n112 10.6151
R1175 B.n375 B.n112 10.6151
R1176 B.n376 B.n375 10.6151
R1177 B.n377 B.n376 10.6151
R1178 B.n377 B.n110 10.6151
R1179 B.n381 B.n110 10.6151
R1180 B.n382 B.n381 10.6151
R1181 B.n383 B.n382 10.6151
R1182 B.n383 B.n108 10.6151
R1183 B.n387 B.n108 10.6151
R1184 B.n388 B.n387 10.6151
R1185 B.n389 B.n388 10.6151
R1186 B.n389 B.n106 10.6151
R1187 B.n393 B.n106 10.6151
R1188 B.n394 B.n393 10.6151
R1189 B.n395 B.n394 10.6151
R1190 B.n395 B.n104 10.6151
R1191 B.n399 B.n104 10.6151
R1192 B.n400 B.n399 10.6151
R1193 B.n401 B.n400 10.6151
R1194 B.n401 B.n102 10.6151
R1195 B.n405 B.n102 10.6151
R1196 B.n693 B.n0 8.11757
R1197 B.n693 B.n1 8.11757
R1198 B.n570 B.n44 6.5566
R1199 B.n558 B.n557 6.5566
R1200 B.n300 B.n299 6.5566
R1201 B.n312 B.n134 6.5566
R1202 B.n573 B.n44 4.05904
R1203 B.n557 B.n556 4.05904
R1204 B.n299 B.n298 4.05904
R1205 B.n315 B.n134 4.05904
C0 VN VDD1 0.148351f
C1 VN VTAIL 5.41749f
C2 VN B 0.775418f
C3 VTAIL VDD1 30.6713f
C4 VDD2 VN 6.07716f
C5 VN VP 6.23039f
C6 VDD1 B 1.9892f
C7 VTAIL B 3.51814f
C8 VN w_n1738_n4676# 3.13821f
C9 VDD2 VDD1 0.733759f
C10 VDD1 VP 6.21439f
C11 VDD2 VTAIL 30.6965f
C12 VTAIL VP 5.4326f
C13 VDD1 w_n1738_n4676# 2.3529f
C14 VDD2 B 2.01857f
C15 VP B 1.1314f
C16 VTAIL w_n1738_n4676# 4.11224f
C17 B w_n1738_n4676# 8.54523f
C18 VDD2 VP 0.293443f
C19 VDD2 w_n1738_n4676# 2.37752f
C20 VP w_n1738_n4676# 3.35742f
C21 VDD2 VSUBS 1.758379f
C22 VDD1 VSUBS 1.234287f
C23 VTAIL VSUBS 0.698912f
C24 VN VSUBS 5.24545f
C25 VP VSUBS 1.578381f
C26 B VSUBS 3.073959f
C27 w_n1738_n4676# VSUBS 99.337105f
C28 B.n0 VSUBS 0.007404f
C29 B.n1 VSUBS 0.007404f
C30 B.n2 VSUBS 0.01095f
C31 B.n3 VSUBS 0.008391f
C32 B.n4 VSUBS 0.008391f
C33 B.n5 VSUBS 0.008391f
C34 B.n6 VSUBS 0.008391f
C35 B.n7 VSUBS 0.008391f
C36 B.n8 VSUBS 0.008391f
C37 B.n9 VSUBS 0.008391f
C38 B.n10 VSUBS 0.008391f
C39 B.n11 VSUBS 0.019468f
C40 B.n12 VSUBS 0.008391f
C41 B.n13 VSUBS 0.008391f
C42 B.n14 VSUBS 0.008391f
C43 B.n15 VSUBS 0.008391f
C44 B.n16 VSUBS 0.008391f
C45 B.n17 VSUBS 0.008391f
C46 B.n18 VSUBS 0.008391f
C47 B.n19 VSUBS 0.008391f
C48 B.n20 VSUBS 0.008391f
C49 B.n21 VSUBS 0.008391f
C50 B.n22 VSUBS 0.008391f
C51 B.n23 VSUBS 0.008391f
C52 B.n24 VSUBS 0.008391f
C53 B.n25 VSUBS 0.008391f
C54 B.n26 VSUBS 0.008391f
C55 B.n27 VSUBS 0.008391f
C56 B.n28 VSUBS 0.008391f
C57 B.n29 VSUBS 0.008391f
C58 B.n30 VSUBS 0.008391f
C59 B.n31 VSUBS 0.008391f
C60 B.n32 VSUBS 0.008391f
C61 B.n33 VSUBS 0.008391f
C62 B.n34 VSUBS 0.008391f
C63 B.n35 VSUBS 0.008391f
C64 B.n36 VSUBS 0.008391f
C65 B.n37 VSUBS 0.008391f
C66 B.n38 VSUBS 0.008391f
C67 B.n39 VSUBS 0.008391f
C68 B.n40 VSUBS 0.008391f
C69 B.n41 VSUBS 0.008391f
C70 B.t4 VSUBS 0.751823f
C71 B.t5 VSUBS 0.758242f
C72 B.t3 VSUBS 0.267206f
C73 B.n42 VSUBS 0.148361f
C74 B.n43 VSUBS 0.075084f
C75 B.n44 VSUBS 0.019441f
C76 B.n45 VSUBS 0.008391f
C77 B.n46 VSUBS 0.008391f
C78 B.n47 VSUBS 0.008391f
C79 B.n48 VSUBS 0.008391f
C80 B.n49 VSUBS 0.008391f
C81 B.t7 VSUBS 0.751794f
C82 B.t8 VSUBS 0.758215f
C83 B.t6 VSUBS 0.267206f
C84 B.n50 VSUBS 0.148388f
C85 B.n51 VSUBS 0.075113f
C86 B.n52 VSUBS 0.008391f
C87 B.n53 VSUBS 0.008391f
C88 B.n54 VSUBS 0.008391f
C89 B.n55 VSUBS 0.008391f
C90 B.n56 VSUBS 0.008391f
C91 B.n57 VSUBS 0.008391f
C92 B.n58 VSUBS 0.008391f
C93 B.n59 VSUBS 0.008391f
C94 B.n60 VSUBS 0.008391f
C95 B.n61 VSUBS 0.008391f
C96 B.n62 VSUBS 0.008391f
C97 B.n63 VSUBS 0.008391f
C98 B.n64 VSUBS 0.008391f
C99 B.n65 VSUBS 0.008391f
C100 B.n66 VSUBS 0.008391f
C101 B.n67 VSUBS 0.008391f
C102 B.n68 VSUBS 0.008391f
C103 B.n69 VSUBS 0.008391f
C104 B.n70 VSUBS 0.008391f
C105 B.n71 VSUBS 0.008391f
C106 B.n72 VSUBS 0.008391f
C107 B.n73 VSUBS 0.008391f
C108 B.n74 VSUBS 0.008391f
C109 B.n75 VSUBS 0.008391f
C110 B.n76 VSUBS 0.008391f
C111 B.n77 VSUBS 0.008391f
C112 B.n78 VSUBS 0.008391f
C113 B.n79 VSUBS 0.008391f
C114 B.n80 VSUBS 0.008391f
C115 B.n81 VSUBS 0.020019f
C116 B.n82 VSUBS 0.008391f
C117 B.n83 VSUBS 0.008391f
C118 B.n84 VSUBS 0.008391f
C119 B.n85 VSUBS 0.008391f
C120 B.n86 VSUBS 0.008391f
C121 B.n87 VSUBS 0.008391f
C122 B.n88 VSUBS 0.008391f
C123 B.n89 VSUBS 0.008391f
C124 B.n90 VSUBS 0.008391f
C125 B.n91 VSUBS 0.008391f
C126 B.n92 VSUBS 0.008391f
C127 B.n93 VSUBS 0.008391f
C128 B.n94 VSUBS 0.008391f
C129 B.n95 VSUBS 0.008391f
C130 B.n96 VSUBS 0.008391f
C131 B.n97 VSUBS 0.008391f
C132 B.n98 VSUBS 0.008391f
C133 B.n99 VSUBS 0.008391f
C134 B.n100 VSUBS 0.008391f
C135 B.n101 VSUBS 0.019468f
C136 B.n102 VSUBS 0.008391f
C137 B.n103 VSUBS 0.008391f
C138 B.n104 VSUBS 0.008391f
C139 B.n105 VSUBS 0.008391f
C140 B.n106 VSUBS 0.008391f
C141 B.n107 VSUBS 0.008391f
C142 B.n108 VSUBS 0.008391f
C143 B.n109 VSUBS 0.008391f
C144 B.n110 VSUBS 0.008391f
C145 B.n111 VSUBS 0.008391f
C146 B.n112 VSUBS 0.008391f
C147 B.n113 VSUBS 0.008391f
C148 B.n114 VSUBS 0.008391f
C149 B.n115 VSUBS 0.008391f
C150 B.n116 VSUBS 0.008391f
C151 B.n117 VSUBS 0.008391f
C152 B.n118 VSUBS 0.008391f
C153 B.n119 VSUBS 0.008391f
C154 B.n120 VSUBS 0.008391f
C155 B.n121 VSUBS 0.008391f
C156 B.n122 VSUBS 0.008391f
C157 B.n123 VSUBS 0.008391f
C158 B.n124 VSUBS 0.008391f
C159 B.n125 VSUBS 0.008391f
C160 B.n126 VSUBS 0.008391f
C161 B.n127 VSUBS 0.008391f
C162 B.n128 VSUBS 0.008391f
C163 B.n129 VSUBS 0.008391f
C164 B.n130 VSUBS 0.008391f
C165 B.n131 VSUBS 0.008391f
C166 B.t2 VSUBS 0.751794f
C167 B.t1 VSUBS 0.758215f
C168 B.t0 VSUBS 0.267206f
C169 B.n132 VSUBS 0.148388f
C170 B.n133 VSUBS 0.075113f
C171 B.n134 VSUBS 0.019441f
C172 B.n135 VSUBS 0.008391f
C173 B.n136 VSUBS 0.008391f
C174 B.n137 VSUBS 0.008391f
C175 B.n138 VSUBS 0.008391f
C176 B.n139 VSUBS 0.008391f
C177 B.t11 VSUBS 0.751823f
C178 B.t10 VSUBS 0.758242f
C179 B.t9 VSUBS 0.267206f
C180 B.n140 VSUBS 0.148361f
C181 B.n141 VSUBS 0.075084f
C182 B.n142 VSUBS 0.008391f
C183 B.n143 VSUBS 0.008391f
C184 B.n144 VSUBS 0.008391f
C185 B.n145 VSUBS 0.008391f
C186 B.n146 VSUBS 0.008391f
C187 B.n147 VSUBS 0.008391f
C188 B.n148 VSUBS 0.008391f
C189 B.n149 VSUBS 0.008391f
C190 B.n150 VSUBS 0.008391f
C191 B.n151 VSUBS 0.008391f
C192 B.n152 VSUBS 0.008391f
C193 B.n153 VSUBS 0.008391f
C194 B.n154 VSUBS 0.008391f
C195 B.n155 VSUBS 0.008391f
C196 B.n156 VSUBS 0.008391f
C197 B.n157 VSUBS 0.008391f
C198 B.n158 VSUBS 0.008391f
C199 B.n159 VSUBS 0.008391f
C200 B.n160 VSUBS 0.008391f
C201 B.n161 VSUBS 0.008391f
C202 B.n162 VSUBS 0.008391f
C203 B.n163 VSUBS 0.008391f
C204 B.n164 VSUBS 0.008391f
C205 B.n165 VSUBS 0.008391f
C206 B.n166 VSUBS 0.008391f
C207 B.n167 VSUBS 0.008391f
C208 B.n168 VSUBS 0.008391f
C209 B.n169 VSUBS 0.008391f
C210 B.n170 VSUBS 0.008391f
C211 B.n171 VSUBS 0.020019f
C212 B.n172 VSUBS 0.008391f
C213 B.n173 VSUBS 0.008391f
C214 B.n174 VSUBS 0.008391f
C215 B.n175 VSUBS 0.008391f
C216 B.n176 VSUBS 0.008391f
C217 B.n177 VSUBS 0.008391f
C218 B.n178 VSUBS 0.008391f
C219 B.n179 VSUBS 0.008391f
C220 B.n180 VSUBS 0.008391f
C221 B.n181 VSUBS 0.008391f
C222 B.n182 VSUBS 0.008391f
C223 B.n183 VSUBS 0.008391f
C224 B.n184 VSUBS 0.008391f
C225 B.n185 VSUBS 0.008391f
C226 B.n186 VSUBS 0.008391f
C227 B.n187 VSUBS 0.008391f
C228 B.n188 VSUBS 0.008391f
C229 B.n189 VSUBS 0.008391f
C230 B.n190 VSUBS 0.008391f
C231 B.n191 VSUBS 0.008391f
C232 B.n192 VSUBS 0.008391f
C233 B.n193 VSUBS 0.008391f
C234 B.n194 VSUBS 0.008391f
C235 B.n195 VSUBS 0.008391f
C236 B.n196 VSUBS 0.008391f
C237 B.n197 VSUBS 0.008391f
C238 B.n198 VSUBS 0.008391f
C239 B.n199 VSUBS 0.008391f
C240 B.n200 VSUBS 0.008391f
C241 B.n201 VSUBS 0.008391f
C242 B.n202 VSUBS 0.008391f
C243 B.n203 VSUBS 0.008391f
C244 B.n204 VSUBS 0.008391f
C245 B.n205 VSUBS 0.008391f
C246 B.n206 VSUBS 0.019468f
C247 B.n207 VSUBS 0.019468f
C248 B.n208 VSUBS 0.020019f
C249 B.n209 VSUBS 0.008391f
C250 B.n210 VSUBS 0.008391f
C251 B.n211 VSUBS 0.008391f
C252 B.n212 VSUBS 0.008391f
C253 B.n213 VSUBS 0.008391f
C254 B.n214 VSUBS 0.008391f
C255 B.n215 VSUBS 0.008391f
C256 B.n216 VSUBS 0.008391f
C257 B.n217 VSUBS 0.008391f
C258 B.n218 VSUBS 0.008391f
C259 B.n219 VSUBS 0.008391f
C260 B.n220 VSUBS 0.008391f
C261 B.n221 VSUBS 0.008391f
C262 B.n222 VSUBS 0.008391f
C263 B.n223 VSUBS 0.008391f
C264 B.n224 VSUBS 0.008391f
C265 B.n225 VSUBS 0.008391f
C266 B.n226 VSUBS 0.008391f
C267 B.n227 VSUBS 0.008391f
C268 B.n228 VSUBS 0.008391f
C269 B.n229 VSUBS 0.008391f
C270 B.n230 VSUBS 0.008391f
C271 B.n231 VSUBS 0.008391f
C272 B.n232 VSUBS 0.008391f
C273 B.n233 VSUBS 0.008391f
C274 B.n234 VSUBS 0.008391f
C275 B.n235 VSUBS 0.008391f
C276 B.n236 VSUBS 0.008391f
C277 B.n237 VSUBS 0.008391f
C278 B.n238 VSUBS 0.008391f
C279 B.n239 VSUBS 0.008391f
C280 B.n240 VSUBS 0.008391f
C281 B.n241 VSUBS 0.008391f
C282 B.n242 VSUBS 0.008391f
C283 B.n243 VSUBS 0.008391f
C284 B.n244 VSUBS 0.008391f
C285 B.n245 VSUBS 0.008391f
C286 B.n246 VSUBS 0.008391f
C287 B.n247 VSUBS 0.008391f
C288 B.n248 VSUBS 0.008391f
C289 B.n249 VSUBS 0.008391f
C290 B.n250 VSUBS 0.008391f
C291 B.n251 VSUBS 0.008391f
C292 B.n252 VSUBS 0.008391f
C293 B.n253 VSUBS 0.008391f
C294 B.n254 VSUBS 0.008391f
C295 B.n255 VSUBS 0.008391f
C296 B.n256 VSUBS 0.008391f
C297 B.n257 VSUBS 0.008391f
C298 B.n258 VSUBS 0.008391f
C299 B.n259 VSUBS 0.008391f
C300 B.n260 VSUBS 0.008391f
C301 B.n261 VSUBS 0.008391f
C302 B.n262 VSUBS 0.008391f
C303 B.n263 VSUBS 0.008391f
C304 B.n264 VSUBS 0.008391f
C305 B.n265 VSUBS 0.008391f
C306 B.n266 VSUBS 0.008391f
C307 B.n267 VSUBS 0.008391f
C308 B.n268 VSUBS 0.008391f
C309 B.n269 VSUBS 0.008391f
C310 B.n270 VSUBS 0.008391f
C311 B.n271 VSUBS 0.008391f
C312 B.n272 VSUBS 0.008391f
C313 B.n273 VSUBS 0.008391f
C314 B.n274 VSUBS 0.008391f
C315 B.n275 VSUBS 0.008391f
C316 B.n276 VSUBS 0.008391f
C317 B.n277 VSUBS 0.008391f
C318 B.n278 VSUBS 0.008391f
C319 B.n279 VSUBS 0.008391f
C320 B.n280 VSUBS 0.008391f
C321 B.n281 VSUBS 0.008391f
C322 B.n282 VSUBS 0.008391f
C323 B.n283 VSUBS 0.008391f
C324 B.n284 VSUBS 0.008391f
C325 B.n285 VSUBS 0.008391f
C326 B.n286 VSUBS 0.008391f
C327 B.n287 VSUBS 0.008391f
C328 B.n288 VSUBS 0.008391f
C329 B.n289 VSUBS 0.008391f
C330 B.n290 VSUBS 0.008391f
C331 B.n291 VSUBS 0.008391f
C332 B.n292 VSUBS 0.008391f
C333 B.n293 VSUBS 0.008391f
C334 B.n294 VSUBS 0.008391f
C335 B.n295 VSUBS 0.008391f
C336 B.n296 VSUBS 0.008391f
C337 B.n297 VSUBS 0.008391f
C338 B.n298 VSUBS 0.0058f
C339 B.n299 VSUBS 0.019441f
C340 B.n300 VSUBS 0.006787f
C341 B.n301 VSUBS 0.008391f
C342 B.n302 VSUBS 0.008391f
C343 B.n303 VSUBS 0.008391f
C344 B.n304 VSUBS 0.008391f
C345 B.n305 VSUBS 0.008391f
C346 B.n306 VSUBS 0.008391f
C347 B.n307 VSUBS 0.008391f
C348 B.n308 VSUBS 0.008391f
C349 B.n309 VSUBS 0.008391f
C350 B.n310 VSUBS 0.008391f
C351 B.n311 VSUBS 0.008391f
C352 B.n312 VSUBS 0.006787f
C353 B.n313 VSUBS 0.008391f
C354 B.n314 VSUBS 0.008391f
C355 B.n315 VSUBS 0.0058f
C356 B.n316 VSUBS 0.008391f
C357 B.n317 VSUBS 0.008391f
C358 B.n318 VSUBS 0.008391f
C359 B.n319 VSUBS 0.008391f
C360 B.n320 VSUBS 0.008391f
C361 B.n321 VSUBS 0.008391f
C362 B.n322 VSUBS 0.008391f
C363 B.n323 VSUBS 0.008391f
C364 B.n324 VSUBS 0.008391f
C365 B.n325 VSUBS 0.008391f
C366 B.n326 VSUBS 0.008391f
C367 B.n327 VSUBS 0.008391f
C368 B.n328 VSUBS 0.008391f
C369 B.n329 VSUBS 0.008391f
C370 B.n330 VSUBS 0.008391f
C371 B.n331 VSUBS 0.008391f
C372 B.n332 VSUBS 0.008391f
C373 B.n333 VSUBS 0.008391f
C374 B.n334 VSUBS 0.008391f
C375 B.n335 VSUBS 0.008391f
C376 B.n336 VSUBS 0.008391f
C377 B.n337 VSUBS 0.008391f
C378 B.n338 VSUBS 0.008391f
C379 B.n339 VSUBS 0.008391f
C380 B.n340 VSUBS 0.008391f
C381 B.n341 VSUBS 0.008391f
C382 B.n342 VSUBS 0.008391f
C383 B.n343 VSUBS 0.008391f
C384 B.n344 VSUBS 0.008391f
C385 B.n345 VSUBS 0.008391f
C386 B.n346 VSUBS 0.008391f
C387 B.n347 VSUBS 0.008391f
C388 B.n348 VSUBS 0.008391f
C389 B.n349 VSUBS 0.008391f
C390 B.n350 VSUBS 0.008391f
C391 B.n351 VSUBS 0.008391f
C392 B.n352 VSUBS 0.008391f
C393 B.n353 VSUBS 0.008391f
C394 B.n354 VSUBS 0.008391f
C395 B.n355 VSUBS 0.008391f
C396 B.n356 VSUBS 0.008391f
C397 B.n357 VSUBS 0.008391f
C398 B.n358 VSUBS 0.008391f
C399 B.n359 VSUBS 0.008391f
C400 B.n360 VSUBS 0.008391f
C401 B.n361 VSUBS 0.008391f
C402 B.n362 VSUBS 0.008391f
C403 B.n363 VSUBS 0.008391f
C404 B.n364 VSUBS 0.008391f
C405 B.n365 VSUBS 0.008391f
C406 B.n366 VSUBS 0.008391f
C407 B.n367 VSUBS 0.008391f
C408 B.n368 VSUBS 0.008391f
C409 B.n369 VSUBS 0.008391f
C410 B.n370 VSUBS 0.008391f
C411 B.n371 VSUBS 0.008391f
C412 B.n372 VSUBS 0.008391f
C413 B.n373 VSUBS 0.008391f
C414 B.n374 VSUBS 0.008391f
C415 B.n375 VSUBS 0.008391f
C416 B.n376 VSUBS 0.008391f
C417 B.n377 VSUBS 0.008391f
C418 B.n378 VSUBS 0.008391f
C419 B.n379 VSUBS 0.008391f
C420 B.n380 VSUBS 0.008391f
C421 B.n381 VSUBS 0.008391f
C422 B.n382 VSUBS 0.008391f
C423 B.n383 VSUBS 0.008391f
C424 B.n384 VSUBS 0.008391f
C425 B.n385 VSUBS 0.008391f
C426 B.n386 VSUBS 0.008391f
C427 B.n387 VSUBS 0.008391f
C428 B.n388 VSUBS 0.008391f
C429 B.n389 VSUBS 0.008391f
C430 B.n390 VSUBS 0.008391f
C431 B.n391 VSUBS 0.008391f
C432 B.n392 VSUBS 0.008391f
C433 B.n393 VSUBS 0.008391f
C434 B.n394 VSUBS 0.008391f
C435 B.n395 VSUBS 0.008391f
C436 B.n396 VSUBS 0.008391f
C437 B.n397 VSUBS 0.008391f
C438 B.n398 VSUBS 0.008391f
C439 B.n399 VSUBS 0.008391f
C440 B.n400 VSUBS 0.008391f
C441 B.n401 VSUBS 0.008391f
C442 B.n402 VSUBS 0.008391f
C443 B.n403 VSUBS 0.008391f
C444 B.n404 VSUBS 0.020019f
C445 B.n405 VSUBS 0.019036f
C446 B.n406 VSUBS 0.020451f
C447 B.n407 VSUBS 0.008391f
C448 B.n408 VSUBS 0.008391f
C449 B.n409 VSUBS 0.008391f
C450 B.n410 VSUBS 0.008391f
C451 B.n411 VSUBS 0.008391f
C452 B.n412 VSUBS 0.008391f
C453 B.n413 VSUBS 0.008391f
C454 B.n414 VSUBS 0.008391f
C455 B.n415 VSUBS 0.008391f
C456 B.n416 VSUBS 0.008391f
C457 B.n417 VSUBS 0.008391f
C458 B.n418 VSUBS 0.008391f
C459 B.n419 VSUBS 0.008391f
C460 B.n420 VSUBS 0.008391f
C461 B.n421 VSUBS 0.008391f
C462 B.n422 VSUBS 0.008391f
C463 B.n423 VSUBS 0.008391f
C464 B.n424 VSUBS 0.008391f
C465 B.n425 VSUBS 0.008391f
C466 B.n426 VSUBS 0.008391f
C467 B.n427 VSUBS 0.008391f
C468 B.n428 VSUBS 0.008391f
C469 B.n429 VSUBS 0.008391f
C470 B.n430 VSUBS 0.008391f
C471 B.n431 VSUBS 0.008391f
C472 B.n432 VSUBS 0.008391f
C473 B.n433 VSUBS 0.008391f
C474 B.n434 VSUBS 0.008391f
C475 B.n435 VSUBS 0.008391f
C476 B.n436 VSUBS 0.008391f
C477 B.n437 VSUBS 0.008391f
C478 B.n438 VSUBS 0.008391f
C479 B.n439 VSUBS 0.008391f
C480 B.n440 VSUBS 0.008391f
C481 B.n441 VSUBS 0.008391f
C482 B.n442 VSUBS 0.008391f
C483 B.n443 VSUBS 0.008391f
C484 B.n444 VSUBS 0.008391f
C485 B.n445 VSUBS 0.008391f
C486 B.n446 VSUBS 0.008391f
C487 B.n447 VSUBS 0.008391f
C488 B.n448 VSUBS 0.008391f
C489 B.n449 VSUBS 0.008391f
C490 B.n450 VSUBS 0.008391f
C491 B.n451 VSUBS 0.008391f
C492 B.n452 VSUBS 0.008391f
C493 B.n453 VSUBS 0.008391f
C494 B.n454 VSUBS 0.008391f
C495 B.n455 VSUBS 0.008391f
C496 B.n456 VSUBS 0.008391f
C497 B.n457 VSUBS 0.008391f
C498 B.n458 VSUBS 0.008391f
C499 B.n459 VSUBS 0.008391f
C500 B.n460 VSUBS 0.008391f
C501 B.n461 VSUBS 0.008391f
C502 B.n462 VSUBS 0.008391f
C503 B.n463 VSUBS 0.008391f
C504 B.n464 VSUBS 0.019468f
C505 B.n465 VSUBS 0.019468f
C506 B.n466 VSUBS 0.020019f
C507 B.n467 VSUBS 0.008391f
C508 B.n468 VSUBS 0.008391f
C509 B.n469 VSUBS 0.008391f
C510 B.n470 VSUBS 0.008391f
C511 B.n471 VSUBS 0.008391f
C512 B.n472 VSUBS 0.008391f
C513 B.n473 VSUBS 0.008391f
C514 B.n474 VSUBS 0.008391f
C515 B.n475 VSUBS 0.008391f
C516 B.n476 VSUBS 0.008391f
C517 B.n477 VSUBS 0.008391f
C518 B.n478 VSUBS 0.008391f
C519 B.n479 VSUBS 0.008391f
C520 B.n480 VSUBS 0.008391f
C521 B.n481 VSUBS 0.008391f
C522 B.n482 VSUBS 0.008391f
C523 B.n483 VSUBS 0.008391f
C524 B.n484 VSUBS 0.008391f
C525 B.n485 VSUBS 0.008391f
C526 B.n486 VSUBS 0.008391f
C527 B.n487 VSUBS 0.008391f
C528 B.n488 VSUBS 0.008391f
C529 B.n489 VSUBS 0.008391f
C530 B.n490 VSUBS 0.008391f
C531 B.n491 VSUBS 0.008391f
C532 B.n492 VSUBS 0.008391f
C533 B.n493 VSUBS 0.008391f
C534 B.n494 VSUBS 0.008391f
C535 B.n495 VSUBS 0.008391f
C536 B.n496 VSUBS 0.008391f
C537 B.n497 VSUBS 0.008391f
C538 B.n498 VSUBS 0.008391f
C539 B.n499 VSUBS 0.008391f
C540 B.n500 VSUBS 0.008391f
C541 B.n501 VSUBS 0.008391f
C542 B.n502 VSUBS 0.008391f
C543 B.n503 VSUBS 0.008391f
C544 B.n504 VSUBS 0.008391f
C545 B.n505 VSUBS 0.008391f
C546 B.n506 VSUBS 0.008391f
C547 B.n507 VSUBS 0.008391f
C548 B.n508 VSUBS 0.008391f
C549 B.n509 VSUBS 0.008391f
C550 B.n510 VSUBS 0.008391f
C551 B.n511 VSUBS 0.008391f
C552 B.n512 VSUBS 0.008391f
C553 B.n513 VSUBS 0.008391f
C554 B.n514 VSUBS 0.008391f
C555 B.n515 VSUBS 0.008391f
C556 B.n516 VSUBS 0.008391f
C557 B.n517 VSUBS 0.008391f
C558 B.n518 VSUBS 0.008391f
C559 B.n519 VSUBS 0.008391f
C560 B.n520 VSUBS 0.008391f
C561 B.n521 VSUBS 0.008391f
C562 B.n522 VSUBS 0.008391f
C563 B.n523 VSUBS 0.008391f
C564 B.n524 VSUBS 0.008391f
C565 B.n525 VSUBS 0.008391f
C566 B.n526 VSUBS 0.008391f
C567 B.n527 VSUBS 0.008391f
C568 B.n528 VSUBS 0.008391f
C569 B.n529 VSUBS 0.008391f
C570 B.n530 VSUBS 0.008391f
C571 B.n531 VSUBS 0.008391f
C572 B.n532 VSUBS 0.008391f
C573 B.n533 VSUBS 0.008391f
C574 B.n534 VSUBS 0.008391f
C575 B.n535 VSUBS 0.008391f
C576 B.n536 VSUBS 0.008391f
C577 B.n537 VSUBS 0.008391f
C578 B.n538 VSUBS 0.008391f
C579 B.n539 VSUBS 0.008391f
C580 B.n540 VSUBS 0.008391f
C581 B.n541 VSUBS 0.008391f
C582 B.n542 VSUBS 0.008391f
C583 B.n543 VSUBS 0.008391f
C584 B.n544 VSUBS 0.008391f
C585 B.n545 VSUBS 0.008391f
C586 B.n546 VSUBS 0.008391f
C587 B.n547 VSUBS 0.008391f
C588 B.n548 VSUBS 0.008391f
C589 B.n549 VSUBS 0.008391f
C590 B.n550 VSUBS 0.008391f
C591 B.n551 VSUBS 0.008391f
C592 B.n552 VSUBS 0.008391f
C593 B.n553 VSUBS 0.008391f
C594 B.n554 VSUBS 0.008391f
C595 B.n555 VSUBS 0.008391f
C596 B.n556 VSUBS 0.0058f
C597 B.n557 VSUBS 0.019441f
C598 B.n558 VSUBS 0.006787f
C599 B.n559 VSUBS 0.008391f
C600 B.n560 VSUBS 0.008391f
C601 B.n561 VSUBS 0.008391f
C602 B.n562 VSUBS 0.008391f
C603 B.n563 VSUBS 0.008391f
C604 B.n564 VSUBS 0.008391f
C605 B.n565 VSUBS 0.008391f
C606 B.n566 VSUBS 0.008391f
C607 B.n567 VSUBS 0.008391f
C608 B.n568 VSUBS 0.008391f
C609 B.n569 VSUBS 0.008391f
C610 B.n570 VSUBS 0.006787f
C611 B.n571 VSUBS 0.008391f
C612 B.n572 VSUBS 0.008391f
C613 B.n573 VSUBS 0.0058f
C614 B.n574 VSUBS 0.008391f
C615 B.n575 VSUBS 0.008391f
C616 B.n576 VSUBS 0.008391f
C617 B.n577 VSUBS 0.008391f
C618 B.n578 VSUBS 0.008391f
C619 B.n579 VSUBS 0.008391f
C620 B.n580 VSUBS 0.008391f
C621 B.n581 VSUBS 0.008391f
C622 B.n582 VSUBS 0.008391f
C623 B.n583 VSUBS 0.008391f
C624 B.n584 VSUBS 0.008391f
C625 B.n585 VSUBS 0.008391f
C626 B.n586 VSUBS 0.008391f
C627 B.n587 VSUBS 0.008391f
C628 B.n588 VSUBS 0.008391f
C629 B.n589 VSUBS 0.008391f
C630 B.n590 VSUBS 0.008391f
C631 B.n591 VSUBS 0.008391f
C632 B.n592 VSUBS 0.008391f
C633 B.n593 VSUBS 0.008391f
C634 B.n594 VSUBS 0.008391f
C635 B.n595 VSUBS 0.008391f
C636 B.n596 VSUBS 0.008391f
C637 B.n597 VSUBS 0.008391f
C638 B.n598 VSUBS 0.008391f
C639 B.n599 VSUBS 0.008391f
C640 B.n600 VSUBS 0.008391f
C641 B.n601 VSUBS 0.008391f
C642 B.n602 VSUBS 0.008391f
C643 B.n603 VSUBS 0.008391f
C644 B.n604 VSUBS 0.008391f
C645 B.n605 VSUBS 0.008391f
C646 B.n606 VSUBS 0.008391f
C647 B.n607 VSUBS 0.008391f
C648 B.n608 VSUBS 0.008391f
C649 B.n609 VSUBS 0.008391f
C650 B.n610 VSUBS 0.008391f
C651 B.n611 VSUBS 0.008391f
C652 B.n612 VSUBS 0.008391f
C653 B.n613 VSUBS 0.008391f
C654 B.n614 VSUBS 0.008391f
C655 B.n615 VSUBS 0.008391f
C656 B.n616 VSUBS 0.008391f
C657 B.n617 VSUBS 0.008391f
C658 B.n618 VSUBS 0.008391f
C659 B.n619 VSUBS 0.008391f
C660 B.n620 VSUBS 0.008391f
C661 B.n621 VSUBS 0.008391f
C662 B.n622 VSUBS 0.008391f
C663 B.n623 VSUBS 0.008391f
C664 B.n624 VSUBS 0.008391f
C665 B.n625 VSUBS 0.008391f
C666 B.n626 VSUBS 0.008391f
C667 B.n627 VSUBS 0.008391f
C668 B.n628 VSUBS 0.008391f
C669 B.n629 VSUBS 0.008391f
C670 B.n630 VSUBS 0.008391f
C671 B.n631 VSUBS 0.008391f
C672 B.n632 VSUBS 0.008391f
C673 B.n633 VSUBS 0.008391f
C674 B.n634 VSUBS 0.008391f
C675 B.n635 VSUBS 0.008391f
C676 B.n636 VSUBS 0.008391f
C677 B.n637 VSUBS 0.008391f
C678 B.n638 VSUBS 0.008391f
C679 B.n639 VSUBS 0.008391f
C680 B.n640 VSUBS 0.008391f
C681 B.n641 VSUBS 0.008391f
C682 B.n642 VSUBS 0.008391f
C683 B.n643 VSUBS 0.008391f
C684 B.n644 VSUBS 0.008391f
C685 B.n645 VSUBS 0.008391f
C686 B.n646 VSUBS 0.008391f
C687 B.n647 VSUBS 0.008391f
C688 B.n648 VSUBS 0.008391f
C689 B.n649 VSUBS 0.008391f
C690 B.n650 VSUBS 0.008391f
C691 B.n651 VSUBS 0.008391f
C692 B.n652 VSUBS 0.008391f
C693 B.n653 VSUBS 0.008391f
C694 B.n654 VSUBS 0.008391f
C695 B.n655 VSUBS 0.008391f
C696 B.n656 VSUBS 0.008391f
C697 B.n657 VSUBS 0.008391f
C698 B.n658 VSUBS 0.008391f
C699 B.n659 VSUBS 0.008391f
C700 B.n660 VSUBS 0.008391f
C701 B.n661 VSUBS 0.008391f
C702 B.n662 VSUBS 0.020019f
C703 B.n663 VSUBS 0.020019f
C704 B.n664 VSUBS 0.019468f
C705 B.n665 VSUBS 0.008391f
C706 B.n666 VSUBS 0.008391f
C707 B.n667 VSUBS 0.008391f
C708 B.n668 VSUBS 0.008391f
C709 B.n669 VSUBS 0.008391f
C710 B.n670 VSUBS 0.008391f
C711 B.n671 VSUBS 0.008391f
C712 B.n672 VSUBS 0.008391f
C713 B.n673 VSUBS 0.008391f
C714 B.n674 VSUBS 0.008391f
C715 B.n675 VSUBS 0.008391f
C716 B.n676 VSUBS 0.008391f
C717 B.n677 VSUBS 0.008391f
C718 B.n678 VSUBS 0.008391f
C719 B.n679 VSUBS 0.008391f
C720 B.n680 VSUBS 0.008391f
C721 B.n681 VSUBS 0.008391f
C722 B.n682 VSUBS 0.008391f
C723 B.n683 VSUBS 0.008391f
C724 B.n684 VSUBS 0.008391f
C725 B.n685 VSUBS 0.008391f
C726 B.n686 VSUBS 0.008391f
C727 B.n687 VSUBS 0.008391f
C728 B.n688 VSUBS 0.008391f
C729 B.n689 VSUBS 0.008391f
C730 B.n690 VSUBS 0.008391f
C731 B.n691 VSUBS 0.01095f
C732 B.n692 VSUBS 0.011664f
C733 B.n693 VSUBS 0.023196f
C734 VDD2.t7 VSUBS 5.27985f
C735 VDD2.t1 VSUBS 0.488613f
C736 VDD2.t0 VSUBS 0.488613f
C737 VDD2.n0 VSUBS 4.06494f
C738 VDD2.n1 VSUBS 1.60622f
C739 VDD2.t3 VSUBS 0.488613f
C740 VDD2.t2 VSUBS 0.488613f
C741 VDD2.n2 VSUBS 4.06908f
C742 VDD2.n3 VSUBS 3.18921f
C743 VDD2.t8 VSUBS 5.27302f
C744 VDD2.n4 VSUBS 4.09f
C745 VDD2.t5 VSUBS 0.488613f
C746 VDD2.t4 VSUBS 0.488613f
C747 VDD2.n5 VSUBS 4.06494f
C748 VDD2.n6 VSUBS 0.749514f
C749 VDD2.t9 VSUBS 0.488613f
C750 VDD2.t6 VSUBS 0.488613f
C751 VDD2.n7 VSUBS 4.06902f
C752 VN.n0 VSUBS 0.062653f
C753 VN.t6 VSUBS 1.01459f
C754 VN.t9 VSUBS 1.01459f
C755 VN.n1 VSUBS 0.026192f
C756 VN.t2 VSUBS 1.02447f
C757 VN.t8 VSUBS 1.01459f
C758 VN.n2 VSUBS 0.379282f
C759 VN.n3 VSUBS 0.399154f
C760 VN.n4 VSUBS 0.139508f
C761 VN.n5 VSUBS 0.062653f
C762 VN.n6 VSUBS 0.400066f
C763 VN.n7 VSUBS 0.026192f
C764 VN.n8 VSUBS 0.379282f
C765 VN.t7 VSUBS 1.02447f
C766 VN.n9 VSUBS 0.399063f
C767 VN.n10 VSUBS 0.048554f
C768 VN.n11 VSUBS 0.062653f
C769 VN.t1 VSUBS 1.02447f
C770 VN.t4 VSUBS 1.01459f
C771 VN.t5 VSUBS 1.01459f
C772 VN.n12 VSUBS 0.026192f
C773 VN.t0 VSUBS 1.01459f
C774 VN.n13 VSUBS 0.379282f
C775 VN.t3 VSUBS 1.02447f
C776 VN.n14 VSUBS 0.399154f
C777 VN.n15 VSUBS 0.139508f
C778 VN.n16 VSUBS 0.062653f
C779 VN.n17 VSUBS 0.400066f
C780 VN.n18 VSUBS 0.026192f
C781 VN.n19 VSUBS 0.379282f
C782 VN.n20 VSUBS 0.399063f
C783 VN.n21 VSUBS 3.00543f
C784 VDD1.t4 VSUBS 5.02138f
C785 VDD1.t0 VSUBS 0.464691f
C786 VDD1.t1 VSUBS 0.464691f
C787 VDD1.n0 VSUBS 3.86592f
C788 VDD1.n1 VSUBS 1.53025f
C789 VDD1.t7 VSUBS 5.02135f
C790 VDD1.t3 VSUBS 0.464691f
C791 VDD1.t5 VSUBS 0.464691f
C792 VDD1.n2 VSUBS 3.86592f
C793 VDD1.n3 VSUBS 1.52758f
C794 VDD1.t6 VSUBS 0.464691f
C795 VDD1.t2 VSUBS 0.464691f
C796 VDD1.n4 VSUBS 3.86985f
C797 VDD1.n5 VSUBS 3.12059f
C798 VDD1.t8 VSUBS 0.464691f
C799 VDD1.t9 VSUBS 0.464691f
C800 VDD1.n6 VSUBS 3.86591f
C801 VDD1.n7 VSUBS 3.83734f
C802 VTAIL.t7 VSUBS 0.489101f
C803 VTAIL.t5 VSUBS 0.489101f
C804 VTAIL.n0 VSUBS 3.85068f
C805 VTAIL.n1 VSUBS 0.973737f
C806 VTAIL.t8 VSUBS 5.0276f
C807 VTAIL.n2 VSUBS 1.13931f
C808 VTAIL.t15 VSUBS 0.489101f
C809 VTAIL.t12 VSUBS 0.489101f
C810 VTAIL.n3 VSUBS 3.85068f
C811 VTAIL.n4 VSUBS 0.96145f
C812 VTAIL.t10 VSUBS 0.489101f
C813 VTAIL.t14 VSUBS 0.489101f
C814 VTAIL.n5 VSUBS 3.85068f
C815 VTAIL.n6 VSUBS 3.19354f
C816 VTAIL.t4 VSUBS 0.489101f
C817 VTAIL.t18 VSUBS 0.489101f
C818 VTAIL.n7 VSUBS 3.85069f
C819 VTAIL.n8 VSUBS 3.19353f
C820 VTAIL.t19 VSUBS 0.489101f
C821 VTAIL.t3 VSUBS 0.489101f
C822 VTAIL.n9 VSUBS 3.85069f
C823 VTAIL.n10 VSUBS 0.961442f
C824 VTAIL.t2 VSUBS 5.02764f
C825 VTAIL.n11 VSUBS 1.13927f
C826 VTAIL.t11 VSUBS 0.489101f
C827 VTAIL.t13 VSUBS 0.489101f
C828 VTAIL.n12 VSUBS 3.85069f
C829 VTAIL.n13 VSUBS 0.982307f
C830 VTAIL.t17 VSUBS 0.489101f
C831 VTAIL.t9 VSUBS 0.489101f
C832 VTAIL.n14 VSUBS 3.85069f
C833 VTAIL.n15 VSUBS 0.961442f
C834 VTAIL.t16 VSUBS 5.0276f
C835 VTAIL.n16 VSUBS 3.29118f
C836 VTAIL.t0 VSUBS 5.0276f
C837 VTAIL.n17 VSUBS 3.29118f
C838 VTAIL.t1 VSUBS 0.489101f
C839 VTAIL.t6 VSUBS 0.489101f
C840 VTAIL.n18 VSUBS 3.85068f
C841 VTAIL.n19 VSUBS 0.910679f
C842 VP.n0 VSUBS 0.064129f
C843 VP.t3 VSUBS 1.03849f
C844 VP.t4 VSUBS 1.03849f
C845 VP.n1 VSUBS 0.026809f
C846 VP.n2 VSUBS 0.064129f
C847 VP.t1 VSUBS 1.03849f
C848 VP.t8 VSUBS 1.03849f
C849 VP.n3 VSUBS 0.026809f
C850 VP.t5 VSUBS 1.04861f
C851 VP.t9 VSUBS 1.03849f
C852 VP.n4 VSUBS 0.388219f
C853 VP.n5 VSUBS 0.40856f
C854 VP.n6 VSUBS 0.142795f
C855 VP.n7 VSUBS 0.064129f
C856 VP.n8 VSUBS 0.409493f
C857 VP.n9 VSUBS 0.026809f
C858 VP.n10 VSUBS 0.388219f
C859 VP.t0 VSUBS 1.04861f
C860 VP.n11 VSUBS 0.408467f
C861 VP.n12 VSUBS 3.03436f
C862 VP.t2 VSUBS 1.04861f
C863 VP.t6 VSUBS 1.03849f
C864 VP.n13 VSUBS 0.388219f
C865 VP.n14 VSUBS 0.408467f
C866 VP.n15 VSUBS 3.08496f
C867 VP.n16 VSUBS 0.064129f
C868 VP.n17 VSUBS 0.064129f
C869 VP.n18 VSUBS 0.409493f
C870 VP.n19 VSUBS 0.026809f
C871 VP.n20 VSUBS 0.388219f
C872 VP.t7 VSUBS 1.04861f
C873 VP.n21 VSUBS 0.408467f
C874 VP.n22 VSUBS 0.049698f
.ends

