* NGSPICE file created from diff_pair_sample_0382.ext - technology: sky130A

.subckt diff_pair_sample_0382 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t14 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.35
X1 B.t11 B.t9 B.t10 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.35
X2 VTAIL.t13 VP.t1 VDD1.t6 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.35
X3 VTAIL.t15 VP.t2 VDD1.t5 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
X4 VTAIL.t8 VP.t3 VDD1.t4 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.35
X5 B.t8 B.t6 B.t7 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.35
X6 VDD2.t7 VN.t0 VTAIL.t4 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.35
X7 B.t5 B.t3 B.t4 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.35
X8 VDD2.t6 VN.t1 VTAIL.t6 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
X9 VDD2.t5 VN.t2 VTAIL.t1 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.35
X10 VDD1.t3 VP.t4 VTAIL.t10 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
X11 VDD1.t2 VP.t5 VTAIL.t9 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=1.4196 ps=8.06 w=3.64 l=1.35
X12 VDD1.t1 VP.t6 VTAIL.t11 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
X13 VTAIL.t3 VN.t3 VDD2.t4 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.35
X14 B.t2 B.t0 B.t1 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0 ps=0 w=3.64 l=1.35
X15 VTAIL.t0 VN.t4 VDD2.t3 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
X16 VTAIL.t12 VP.t7 VDD1.t0 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
X17 VTAIL.t5 VN.t5 VDD2.t2 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=1.4196 pd=8.06 as=0.6006 ps=3.97 w=3.64 l=1.35
X18 VTAIL.t7 VN.t6 VDD2.t1 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
X19 VDD2.t0 VN.t7 VTAIL.t2 w_n2650_n1696# sky130_fd_pr__pfet_01v8 ad=0.6006 pd=3.97 as=0.6006 ps=3.97 w=3.64 l=1.35
R0 VP.n25 VP.n5 172.499
R1 VP.n44 VP.n43 172.499
R2 VP.n24 VP.n23 172.499
R3 VP.n12 VP.n9 161.3
R4 VP.n14 VP.n13 161.3
R5 VP.n15 VP.n8 161.3
R6 VP.n18 VP.n17 161.3
R7 VP.n19 VP.n7 161.3
R8 VP.n21 VP.n20 161.3
R9 VP.n22 VP.n6 161.3
R10 VP.n42 VP.n0 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n39 VP.n1 161.3
R13 VP.n38 VP.n37 161.3
R14 VP.n35 VP.n2 161.3
R15 VP.n34 VP.n33 161.3
R16 VP.n32 VP.n3 161.3
R17 VP.n31 VP.n30 161.3
R18 VP.n28 VP.n4 161.3
R19 VP.n27 VP.n26 161.3
R20 VP.n11 VP.t1 94.5391
R21 VP.n5 VP.t3 64.9812
R22 VP.n29 VP.t4 64.9812
R23 VP.n36 VP.t2 64.9812
R24 VP.n43 VP.t0 64.9812
R25 VP.n23 VP.t5 64.9812
R26 VP.n16 VP.t7 64.9812
R27 VP.n10 VP.t6 64.9812
R28 VP.n11 VP.n10 60.6301
R29 VP.n35 VP.n34 56.4773
R30 VP.n15 VP.n14 56.4773
R31 VP.n30 VP.n28 47.2268
R32 VP.n41 VP.n1 47.2268
R33 VP.n21 VP.n7 47.2268
R34 VP.n25 VP.n24 38.652
R35 VP.n28 VP.n27 33.5944
R36 VP.n42 VP.n41 33.5944
R37 VP.n22 VP.n21 33.5944
R38 VP.n12 VP.n11 27.0891
R39 VP.n34 VP.n3 24.3439
R40 VP.n37 VP.n35 24.3439
R41 VP.n17 VP.n15 24.3439
R42 VP.n14 VP.n9 24.3439
R43 VP.n30 VP.n29 19.9621
R44 VP.n36 VP.n1 19.9621
R45 VP.n16 VP.n7 19.9621
R46 VP.n27 VP.n5 13.146
R47 VP.n43 VP.n42 13.146
R48 VP.n23 VP.n22 13.146
R49 VP.n29 VP.n3 4.38232
R50 VP.n37 VP.n36 4.38232
R51 VP.n17 VP.n16 4.38232
R52 VP.n10 VP.n9 4.38232
R53 VP.n13 VP.n12 0.189894
R54 VP.n13 VP.n8 0.189894
R55 VP.n18 VP.n8 0.189894
R56 VP.n19 VP.n18 0.189894
R57 VP.n20 VP.n19 0.189894
R58 VP.n20 VP.n6 0.189894
R59 VP.n24 VP.n6 0.189894
R60 VP.n26 VP.n25 0.189894
R61 VP.n26 VP.n4 0.189894
R62 VP.n31 VP.n4 0.189894
R63 VP.n32 VP.n31 0.189894
R64 VP.n33 VP.n32 0.189894
R65 VP.n33 VP.n2 0.189894
R66 VP.n38 VP.n2 0.189894
R67 VP.n39 VP.n38 0.189894
R68 VP.n40 VP.n39 0.189894
R69 VP.n40 VP.n0 0.189894
R70 VP.n44 VP.n0 0.189894
R71 VP VP.n44 0.0516364
R72 VTAIL.n11 VTAIL.t13 115.263
R73 VTAIL.n10 VTAIL.t4 115.263
R74 VTAIL.n7 VTAIL.t5 115.263
R75 VTAIL.n15 VTAIL.t1 115.263
R76 VTAIL.n2 VTAIL.t3 115.263
R77 VTAIL.n3 VTAIL.t14 115.263
R78 VTAIL.n6 VTAIL.t8 115.263
R79 VTAIL.n14 VTAIL.t9 115.263
R80 VTAIL.n13 VTAIL.n12 106.332
R81 VTAIL.n9 VTAIL.n8 106.332
R82 VTAIL.n1 VTAIL.n0 106.332
R83 VTAIL.n5 VTAIL.n4 106.332
R84 VTAIL.n15 VTAIL.n14 16.9531
R85 VTAIL.n7 VTAIL.n6 16.9531
R86 VTAIL.n0 VTAIL.t2 8.93044
R87 VTAIL.n0 VTAIL.t7 8.93044
R88 VTAIL.n4 VTAIL.t10 8.93044
R89 VTAIL.n4 VTAIL.t15 8.93044
R90 VTAIL.n12 VTAIL.t11 8.93044
R91 VTAIL.n12 VTAIL.t12 8.93044
R92 VTAIL.n8 VTAIL.t6 8.93044
R93 VTAIL.n8 VTAIL.t0 8.93044
R94 VTAIL.n9 VTAIL.n7 1.44878
R95 VTAIL.n10 VTAIL.n9 1.44878
R96 VTAIL.n13 VTAIL.n11 1.44878
R97 VTAIL.n14 VTAIL.n13 1.44878
R98 VTAIL.n6 VTAIL.n5 1.44878
R99 VTAIL.n5 VTAIL.n3 1.44878
R100 VTAIL.n2 VTAIL.n1 1.44878
R101 VTAIL VTAIL.n15 1.39059
R102 VTAIL.n11 VTAIL.n10 0.470328
R103 VTAIL.n3 VTAIL.n2 0.470328
R104 VTAIL VTAIL.n1 0.0586897
R105 VDD1 VDD1.n0 123.793
R106 VDD1.n3 VDD1.n2 123.68
R107 VDD1.n3 VDD1.n1 123.68
R108 VDD1.n5 VDD1.n4 123.011
R109 VDD1.n5 VDD1.n3 33.9535
R110 VDD1.n4 VDD1.t0 8.93044
R111 VDD1.n4 VDD1.t2 8.93044
R112 VDD1.n0 VDD1.t6 8.93044
R113 VDD1.n0 VDD1.t1 8.93044
R114 VDD1.n2 VDD1.t5 8.93044
R115 VDD1.n2 VDD1.t7 8.93044
R116 VDD1.n1 VDD1.t4 8.93044
R117 VDD1.n1 VDD1.t3 8.93044
R118 VDD1 VDD1.n5 0.666448
R119 B.n338 B.n337 585
R120 B.n339 B.n44 585
R121 B.n341 B.n340 585
R122 B.n342 B.n43 585
R123 B.n344 B.n343 585
R124 B.n345 B.n42 585
R125 B.n347 B.n346 585
R126 B.n348 B.n41 585
R127 B.n350 B.n349 585
R128 B.n351 B.n40 585
R129 B.n353 B.n352 585
R130 B.n354 B.n39 585
R131 B.n356 B.n355 585
R132 B.n357 B.n38 585
R133 B.n359 B.n358 585
R134 B.n360 B.n37 585
R135 B.n362 B.n361 585
R136 B.n364 B.n363 585
R137 B.n365 B.n33 585
R138 B.n367 B.n366 585
R139 B.n368 B.n32 585
R140 B.n370 B.n369 585
R141 B.n371 B.n31 585
R142 B.n373 B.n372 585
R143 B.n374 B.n30 585
R144 B.n376 B.n375 585
R145 B.n377 B.n27 585
R146 B.n380 B.n379 585
R147 B.n381 B.n26 585
R148 B.n383 B.n382 585
R149 B.n384 B.n25 585
R150 B.n386 B.n385 585
R151 B.n387 B.n24 585
R152 B.n389 B.n388 585
R153 B.n390 B.n23 585
R154 B.n392 B.n391 585
R155 B.n393 B.n22 585
R156 B.n395 B.n394 585
R157 B.n396 B.n21 585
R158 B.n398 B.n397 585
R159 B.n399 B.n20 585
R160 B.n401 B.n400 585
R161 B.n402 B.n19 585
R162 B.n404 B.n403 585
R163 B.n336 B.n45 585
R164 B.n335 B.n334 585
R165 B.n333 B.n46 585
R166 B.n332 B.n331 585
R167 B.n330 B.n47 585
R168 B.n329 B.n328 585
R169 B.n327 B.n48 585
R170 B.n326 B.n325 585
R171 B.n324 B.n49 585
R172 B.n323 B.n322 585
R173 B.n321 B.n50 585
R174 B.n320 B.n319 585
R175 B.n318 B.n51 585
R176 B.n317 B.n316 585
R177 B.n315 B.n52 585
R178 B.n314 B.n313 585
R179 B.n312 B.n53 585
R180 B.n311 B.n310 585
R181 B.n309 B.n54 585
R182 B.n308 B.n307 585
R183 B.n306 B.n55 585
R184 B.n305 B.n304 585
R185 B.n303 B.n56 585
R186 B.n302 B.n301 585
R187 B.n300 B.n57 585
R188 B.n299 B.n298 585
R189 B.n297 B.n58 585
R190 B.n296 B.n295 585
R191 B.n294 B.n59 585
R192 B.n293 B.n292 585
R193 B.n291 B.n60 585
R194 B.n290 B.n289 585
R195 B.n288 B.n61 585
R196 B.n287 B.n286 585
R197 B.n285 B.n62 585
R198 B.n284 B.n283 585
R199 B.n282 B.n63 585
R200 B.n281 B.n280 585
R201 B.n279 B.n64 585
R202 B.n278 B.n277 585
R203 B.n276 B.n65 585
R204 B.n275 B.n274 585
R205 B.n273 B.n66 585
R206 B.n272 B.n271 585
R207 B.n270 B.n67 585
R208 B.n269 B.n268 585
R209 B.n267 B.n68 585
R210 B.n266 B.n265 585
R211 B.n264 B.n69 585
R212 B.n263 B.n262 585
R213 B.n261 B.n70 585
R214 B.n260 B.n259 585
R215 B.n258 B.n71 585
R216 B.n257 B.n256 585
R217 B.n255 B.n72 585
R218 B.n254 B.n253 585
R219 B.n252 B.n73 585
R220 B.n251 B.n250 585
R221 B.n249 B.n74 585
R222 B.n248 B.n247 585
R223 B.n246 B.n75 585
R224 B.n245 B.n244 585
R225 B.n243 B.n76 585
R226 B.n242 B.n241 585
R227 B.n240 B.n77 585
R228 B.n239 B.n238 585
R229 B.n237 B.n78 585
R230 B.n170 B.n169 585
R231 B.n171 B.n104 585
R232 B.n173 B.n172 585
R233 B.n174 B.n103 585
R234 B.n176 B.n175 585
R235 B.n177 B.n102 585
R236 B.n179 B.n178 585
R237 B.n180 B.n101 585
R238 B.n182 B.n181 585
R239 B.n183 B.n100 585
R240 B.n185 B.n184 585
R241 B.n186 B.n99 585
R242 B.n188 B.n187 585
R243 B.n189 B.n98 585
R244 B.n191 B.n190 585
R245 B.n192 B.n97 585
R246 B.n194 B.n193 585
R247 B.n196 B.n195 585
R248 B.n197 B.n93 585
R249 B.n199 B.n198 585
R250 B.n200 B.n92 585
R251 B.n202 B.n201 585
R252 B.n203 B.n91 585
R253 B.n205 B.n204 585
R254 B.n206 B.n90 585
R255 B.n208 B.n207 585
R256 B.n209 B.n87 585
R257 B.n212 B.n211 585
R258 B.n213 B.n86 585
R259 B.n215 B.n214 585
R260 B.n216 B.n85 585
R261 B.n218 B.n217 585
R262 B.n219 B.n84 585
R263 B.n221 B.n220 585
R264 B.n222 B.n83 585
R265 B.n224 B.n223 585
R266 B.n225 B.n82 585
R267 B.n227 B.n226 585
R268 B.n228 B.n81 585
R269 B.n230 B.n229 585
R270 B.n231 B.n80 585
R271 B.n233 B.n232 585
R272 B.n234 B.n79 585
R273 B.n236 B.n235 585
R274 B.n168 B.n105 585
R275 B.n167 B.n166 585
R276 B.n165 B.n106 585
R277 B.n164 B.n163 585
R278 B.n162 B.n107 585
R279 B.n161 B.n160 585
R280 B.n159 B.n108 585
R281 B.n158 B.n157 585
R282 B.n156 B.n109 585
R283 B.n155 B.n154 585
R284 B.n153 B.n110 585
R285 B.n152 B.n151 585
R286 B.n150 B.n111 585
R287 B.n149 B.n148 585
R288 B.n147 B.n112 585
R289 B.n146 B.n145 585
R290 B.n144 B.n113 585
R291 B.n143 B.n142 585
R292 B.n141 B.n114 585
R293 B.n140 B.n139 585
R294 B.n138 B.n115 585
R295 B.n137 B.n136 585
R296 B.n135 B.n116 585
R297 B.n134 B.n133 585
R298 B.n132 B.n117 585
R299 B.n131 B.n130 585
R300 B.n129 B.n118 585
R301 B.n128 B.n127 585
R302 B.n126 B.n119 585
R303 B.n125 B.n124 585
R304 B.n123 B.n120 585
R305 B.n122 B.n121 585
R306 B.n2 B.n0 585
R307 B.n453 B.n1 585
R308 B.n452 B.n451 585
R309 B.n450 B.n3 585
R310 B.n449 B.n448 585
R311 B.n447 B.n4 585
R312 B.n446 B.n445 585
R313 B.n444 B.n5 585
R314 B.n443 B.n442 585
R315 B.n441 B.n6 585
R316 B.n440 B.n439 585
R317 B.n438 B.n7 585
R318 B.n437 B.n436 585
R319 B.n435 B.n8 585
R320 B.n434 B.n433 585
R321 B.n432 B.n9 585
R322 B.n431 B.n430 585
R323 B.n429 B.n10 585
R324 B.n428 B.n427 585
R325 B.n426 B.n11 585
R326 B.n425 B.n424 585
R327 B.n423 B.n12 585
R328 B.n422 B.n421 585
R329 B.n420 B.n13 585
R330 B.n419 B.n418 585
R331 B.n417 B.n14 585
R332 B.n416 B.n415 585
R333 B.n414 B.n15 585
R334 B.n413 B.n412 585
R335 B.n411 B.n16 585
R336 B.n410 B.n409 585
R337 B.n408 B.n17 585
R338 B.n407 B.n406 585
R339 B.n405 B.n18 585
R340 B.n455 B.n454 585
R341 B.n170 B.n105 439.647
R342 B.n405 B.n404 439.647
R343 B.n237 B.n236 439.647
R344 B.n338 B.n45 439.647
R345 B.n88 B.t0 270.457
R346 B.n34 B.t6 270.457
R347 B.n94 B.t9 269.959
R348 B.n28 B.t3 269.959
R349 B.n88 B.t2 163.429
R350 B.n34 B.t7 163.429
R351 B.n94 B.t11 163.427
R352 B.n28 B.t4 163.427
R353 B.n166 B.n105 163.367
R354 B.n166 B.n165 163.367
R355 B.n165 B.n164 163.367
R356 B.n164 B.n107 163.367
R357 B.n160 B.n107 163.367
R358 B.n160 B.n159 163.367
R359 B.n159 B.n158 163.367
R360 B.n158 B.n109 163.367
R361 B.n154 B.n109 163.367
R362 B.n154 B.n153 163.367
R363 B.n153 B.n152 163.367
R364 B.n152 B.n111 163.367
R365 B.n148 B.n111 163.367
R366 B.n148 B.n147 163.367
R367 B.n147 B.n146 163.367
R368 B.n146 B.n113 163.367
R369 B.n142 B.n113 163.367
R370 B.n142 B.n141 163.367
R371 B.n141 B.n140 163.367
R372 B.n140 B.n115 163.367
R373 B.n136 B.n115 163.367
R374 B.n136 B.n135 163.367
R375 B.n135 B.n134 163.367
R376 B.n134 B.n117 163.367
R377 B.n130 B.n117 163.367
R378 B.n130 B.n129 163.367
R379 B.n129 B.n128 163.367
R380 B.n128 B.n119 163.367
R381 B.n124 B.n119 163.367
R382 B.n124 B.n123 163.367
R383 B.n123 B.n122 163.367
R384 B.n122 B.n2 163.367
R385 B.n454 B.n2 163.367
R386 B.n454 B.n453 163.367
R387 B.n453 B.n452 163.367
R388 B.n452 B.n3 163.367
R389 B.n448 B.n3 163.367
R390 B.n448 B.n447 163.367
R391 B.n447 B.n446 163.367
R392 B.n446 B.n5 163.367
R393 B.n442 B.n5 163.367
R394 B.n442 B.n441 163.367
R395 B.n441 B.n440 163.367
R396 B.n440 B.n7 163.367
R397 B.n436 B.n7 163.367
R398 B.n436 B.n435 163.367
R399 B.n435 B.n434 163.367
R400 B.n434 B.n9 163.367
R401 B.n430 B.n9 163.367
R402 B.n430 B.n429 163.367
R403 B.n429 B.n428 163.367
R404 B.n428 B.n11 163.367
R405 B.n424 B.n11 163.367
R406 B.n424 B.n423 163.367
R407 B.n423 B.n422 163.367
R408 B.n422 B.n13 163.367
R409 B.n418 B.n13 163.367
R410 B.n418 B.n417 163.367
R411 B.n417 B.n416 163.367
R412 B.n416 B.n15 163.367
R413 B.n412 B.n15 163.367
R414 B.n412 B.n411 163.367
R415 B.n411 B.n410 163.367
R416 B.n410 B.n17 163.367
R417 B.n406 B.n17 163.367
R418 B.n406 B.n405 163.367
R419 B.n171 B.n170 163.367
R420 B.n172 B.n171 163.367
R421 B.n172 B.n103 163.367
R422 B.n176 B.n103 163.367
R423 B.n177 B.n176 163.367
R424 B.n178 B.n177 163.367
R425 B.n178 B.n101 163.367
R426 B.n182 B.n101 163.367
R427 B.n183 B.n182 163.367
R428 B.n184 B.n183 163.367
R429 B.n184 B.n99 163.367
R430 B.n188 B.n99 163.367
R431 B.n189 B.n188 163.367
R432 B.n190 B.n189 163.367
R433 B.n190 B.n97 163.367
R434 B.n194 B.n97 163.367
R435 B.n195 B.n194 163.367
R436 B.n195 B.n93 163.367
R437 B.n199 B.n93 163.367
R438 B.n200 B.n199 163.367
R439 B.n201 B.n200 163.367
R440 B.n201 B.n91 163.367
R441 B.n205 B.n91 163.367
R442 B.n206 B.n205 163.367
R443 B.n207 B.n206 163.367
R444 B.n207 B.n87 163.367
R445 B.n212 B.n87 163.367
R446 B.n213 B.n212 163.367
R447 B.n214 B.n213 163.367
R448 B.n214 B.n85 163.367
R449 B.n218 B.n85 163.367
R450 B.n219 B.n218 163.367
R451 B.n220 B.n219 163.367
R452 B.n220 B.n83 163.367
R453 B.n224 B.n83 163.367
R454 B.n225 B.n224 163.367
R455 B.n226 B.n225 163.367
R456 B.n226 B.n81 163.367
R457 B.n230 B.n81 163.367
R458 B.n231 B.n230 163.367
R459 B.n232 B.n231 163.367
R460 B.n232 B.n79 163.367
R461 B.n236 B.n79 163.367
R462 B.n238 B.n237 163.367
R463 B.n238 B.n77 163.367
R464 B.n242 B.n77 163.367
R465 B.n243 B.n242 163.367
R466 B.n244 B.n243 163.367
R467 B.n244 B.n75 163.367
R468 B.n248 B.n75 163.367
R469 B.n249 B.n248 163.367
R470 B.n250 B.n249 163.367
R471 B.n250 B.n73 163.367
R472 B.n254 B.n73 163.367
R473 B.n255 B.n254 163.367
R474 B.n256 B.n255 163.367
R475 B.n256 B.n71 163.367
R476 B.n260 B.n71 163.367
R477 B.n261 B.n260 163.367
R478 B.n262 B.n261 163.367
R479 B.n262 B.n69 163.367
R480 B.n266 B.n69 163.367
R481 B.n267 B.n266 163.367
R482 B.n268 B.n267 163.367
R483 B.n268 B.n67 163.367
R484 B.n272 B.n67 163.367
R485 B.n273 B.n272 163.367
R486 B.n274 B.n273 163.367
R487 B.n274 B.n65 163.367
R488 B.n278 B.n65 163.367
R489 B.n279 B.n278 163.367
R490 B.n280 B.n279 163.367
R491 B.n280 B.n63 163.367
R492 B.n284 B.n63 163.367
R493 B.n285 B.n284 163.367
R494 B.n286 B.n285 163.367
R495 B.n286 B.n61 163.367
R496 B.n290 B.n61 163.367
R497 B.n291 B.n290 163.367
R498 B.n292 B.n291 163.367
R499 B.n292 B.n59 163.367
R500 B.n296 B.n59 163.367
R501 B.n297 B.n296 163.367
R502 B.n298 B.n297 163.367
R503 B.n298 B.n57 163.367
R504 B.n302 B.n57 163.367
R505 B.n303 B.n302 163.367
R506 B.n304 B.n303 163.367
R507 B.n304 B.n55 163.367
R508 B.n308 B.n55 163.367
R509 B.n309 B.n308 163.367
R510 B.n310 B.n309 163.367
R511 B.n310 B.n53 163.367
R512 B.n314 B.n53 163.367
R513 B.n315 B.n314 163.367
R514 B.n316 B.n315 163.367
R515 B.n316 B.n51 163.367
R516 B.n320 B.n51 163.367
R517 B.n321 B.n320 163.367
R518 B.n322 B.n321 163.367
R519 B.n322 B.n49 163.367
R520 B.n326 B.n49 163.367
R521 B.n327 B.n326 163.367
R522 B.n328 B.n327 163.367
R523 B.n328 B.n47 163.367
R524 B.n332 B.n47 163.367
R525 B.n333 B.n332 163.367
R526 B.n334 B.n333 163.367
R527 B.n334 B.n45 163.367
R528 B.n404 B.n19 163.367
R529 B.n400 B.n19 163.367
R530 B.n400 B.n399 163.367
R531 B.n399 B.n398 163.367
R532 B.n398 B.n21 163.367
R533 B.n394 B.n21 163.367
R534 B.n394 B.n393 163.367
R535 B.n393 B.n392 163.367
R536 B.n392 B.n23 163.367
R537 B.n388 B.n23 163.367
R538 B.n388 B.n387 163.367
R539 B.n387 B.n386 163.367
R540 B.n386 B.n25 163.367
R541 B.n382 B.n25 163.367
R542 B.n382 B.n381 163.367
R543 B.n381 B.n380 163.367
R544 B.n380 B.n27 163.367
R545 B.n375 B.n27 163.367
R546 B.n375 B.n374 163.367
R547 B.n374 B.n373 163.367
R548 B.n373 B.n31 163.367
R549 B.n369 B.n31 163.367
R550 B.n369 B.n368 163.367
R551 B.n368 B.n367 163.367
R552 B.n367 B.n33 163.367
R553 B.n363 B.n33 163.367
R554 B.n363 B.n362 163.367
R555 B.n362 B.n37 163.367
R556 B.n358 B.n37 163.367
R557 B.n358 B.n357 163.367
R558 B.n357 B.n356 163.367
R559 B.n356 B.n39 163.367
R560 B.n352 B.n39 163.367
R561 B.n352 B.n351 163.367
R562 B.n351 B.n350 163.367
R563 B.n350 B.n41 163.367
R564 B.n346 B.n41 163.367
R565 B.n346 B.n345 163.367
R566 B.n345 B.n344 163.367
R567 B.n344 B.n43 163.367
R568 B.n340 B.n43 163.367
R569 B.n340 B.n339 163.367
R570 B.n339 B.n338 163.367
R571 B.n89 B.t1 130.847
R572 B.n35 B.t8 130.847
R573 B.n95 B.t10 130.845
R574 B.n29 B.t5 130.845
R575 B.n210 B.n89 59.5399
R576 B.n96 B.n95 59.5399
R577 B.n378 B.n29 59.5399
R578 B.n36 B.n35 59.5399
R579 B.n89 B.n88 32.5823
R580 B.n95 B.n94 32.5823
R581 B.n29 B.n28 32.5823
R582 B.n35 B.n34 32.5823
R583 B.n403 B.n18 28.5664
R584 B.n235 B.n78 28.5664
R585 B.n169 B.n168 28.5664
R586 B.n337 B.n336 28.5664
R587 B B.n455 18.0485
R588 B.n403 B.n402 10.6151
R589 B.n402 B.n401 10.6151
R590 B.n401 B.n20 10.6151
R591 B.n397 B.n20 10.6151
R592 B.n397 B.n396 10.6151
R593 B.n396 B.n395 10.6151
R594 B.n395 B.n22 10.6151
R595 B.n391 B.n22 10.6151
R596 B.n391 B.n390 10.6151
R597 B.n390 B.n389 10.6151
R598 B.n389 B.n24 10.6151
R599 B.n385 B.n24 10.6151
R600 B.n385 B.n384 10.6151
R601 B.n384 B.n383 10.6151
R602 B.n383 B.n26 10.6151
R603 B.n379 B.n26 10.6151
R604 B.n377 B.n376 10.6151
R605 B.n376 B.n30 10.6151
R606 B.n372 B.n30 10.6151
R607 B.n372 B.n371 10.6151
R608 B.n371 B.n370 10.6151
R609 B.n370 B.n32 10.6151
R610 B.n366 B.n32 10.6151
R611 B.n366 B.n365 10.6151
R612 B.n365 B.n364 10.6151
R613 B.n361 B.n360 10.6151
R614 B.n360 B.n359 10.6151
R615 B.n359 B.n38 10.6151
R616 B.n355 B.n38 10.6151
R617 B.n355 B.n354 10.6151
R618 B.n354 B.n353 10.6151
R619 B.n353 B.n40 10.6151
R620 B.n349 B.n40 10.6151
R621 B.n349 B.n348 10.6151
R622 B.n348 B.n347 10.6151
R623 B.n347 B.n42 10.6151
R624 B.n343 B.n42 10.6151
R625 B.n343 B.n342 10.6151
R626 B.n342 B.n341 10.6151
R627 B.n341 B.n44 10.6151
R628 B.n337 B.n44 10.6151
R629 B.n239 B.n78 10.6151
R630 B.n240 B.n239 10.6151
R631 B.n241 B.n240 10.6151
R632 B.n241 B.n76 10.6151
R633 B.n245 B.n76 10.6151
R634 B.n246 B.n245 10.6151
R635 B.n247 B.n246 10.6151
R636 B.n247 B.n74 10.6151
R637 B.n251 B.n74 10.6151
R638 B.n252 B.n251 10.6151
R639 B.n253 B.n252 10.6151
R640 B.n253 B.n72 10.6151
R641 B.n257 B.n72 10.6151
R642 B.n258 B.n257 10.6151
R643 B.n259 B.n258 10.6151
R644 B.n259 B.n70 10.6151
R645 B.n263 B.n70 10.6151
R646 B.n264 B.n263 10.6151
R647 B.n265 B.n264 10.6151
R648 B.n265 B.n68 10.6151
R649 B.n269 B.n68 10.6151
R650 B.n270 B.n269 10.6151
R651 B.n271 B.n270 10.6151
R652 B.n271 B.n66 10.6151
R653 B.n275 B.n66 10.6151
R654 B.n276 B.n275 10.6151
R655 B.n277 B.n276 10.6151
R656 B.n277 B.n64 10.6151
R657 B.n281 B.n64 10.6151
R658 B.n282 B.n281 10.6151
R659 B.n283 B.n282 10.6151
R660 B.n283 B.n62 10.6151
R661 B.n287 B.n62 10.6151
R662 B.n288 B.n287 10.6151
R663 B.n289 B.n288 10.6151
R664 B.n289 B.n60 10.6151
R665 B.n293 B.n60 10.6151
R666 B.n294 B.n293 10.6151
R667 B.n295 B.n294 10.6151
R668 B.n295 B.n58 10.6151
R669 B.n299 B.n58 10.6151
R670 B.n300 B.n299 10.6151
R671 B.n301 B.n300 10.6151
R672 B.n301 B.n56 10.6151
R673 B.n305 B.n56 10.6151
R674 B.n306 B.n305 10.6151
R675 B.n307 B.n306 10.6151
R676 B.n307 B.n54 10.6151
R677 B.n311 B.n54 10.6151
R678 B.n312 B.n311 10.6151
R679 B.n313 B.n312 10.6151
R680 B.n313 B.n52 10.6151
R681 B.n317 B.n52 10.6151
R682 B.n318 B.n317 10.6151
R683 B.n319 B.n318 10.6151
R684 B.n319 B.n50 10.6151
R685 B.n323 B.n50 10.6151
R686 B.n324 B.n323 10.6151
R687 B.n325 B.n324 10.6151
R688 B.n325 B.n48 10.6151
R689 B.n329 B.n48 10.6151
R690 B.n330 B.n329 10.6151
R691 B.n331 B.n330 10.6151
R692 B.n331 B.n46 10.6151
R693 B.n335 B.n46 10.6151
R694 B.n336 B.n335 10.6151
R695 B.n169 B.n104 10.6151
R696 B.n173 B.n104 10.6151
R697 B.n174 B.n173 10.6151
R698 B.n175 B.n174 10.6151
R699 B.n175 B.n102 10.6151
R700 B.n179 B.n102 10.6151
R701 B.n180 B.n179 10.6151
R702 B.n181 B.n180 10.6151
R703 B.n181 B.n100 10.6151
R704 B.n185 B.n100 10.6151
R705 B.n186 B.n185 10.6151
R706 B.n187 B.n186 10.6151
R707 B.n187 B.n98 10.6151
R708 B.n191 B.n98 10.6151
R709 B.n192 B.n191 10.6151
R710 B.n193 B.n192 10.6151
R711 B.n197 B.n196 10.6151
R712 B.n198 B.n197 10.6151
R713 B.n198 B.n92 10.6151
R714 B.n202 B.n92 10.6151
R715 B.n203 B.n202 10.6151
R716 B.n204 B.n203 10.6151
R717 B.n204 B.n90 10.6151
R718 B.n208 B.n90 10.6151
R719 B.n209 B.n208 10.6151
R720 B.n211 B.n86 10.6151
R721 B.n215 B.n86 10.6151
R722 B.n216 B.n215 10.6151
R723 B.n217 B.n216 10.6151
R724 B.n217 B.n84 10.6151
R725 B.n221 B.n84 10.6151
R726 B.n222 B.n221 10.6151
R727 B.n223 B.n222 10.6151
R728 B.n223 B.n82 10.6151
R729 B.n227 B.n82 10.6151
R730 B.n228 B.n227 10.6151
R731 B.n229 B.n228 10.6151
R732 B.n229 B.n80 10.6151
R733 B.n233 B.n80 10.6151
R734 B.n234 B.n233 10.6151
R735 B.n235 B.n234 10.6151
R736 B.n168 B.n167 10.6151
R737 B.n167 B.n106 10.6151
R738 B.n163 B.n106 10.6151
R739 B.n163 B.n162 10.6151
R740 B.n162 B.n161 10.6151
R741 B.n161 B.n108 10.6151
R742 B.n157 B.n108 10.6151
R743 B.n157 B.n156 10.6151
R744 B.n156 B.n155 10.6151
R745 B.n155 B.n110 10.6151
R746 B.n151 B.n110 10.6151
R747 B.n151 B.n150 10.6151
R748 B.n150 B.n149 10.6151
R749 B.n149 B.n112 10.6151
R750 B.n145 B.n112 10.6151
R751 B.n145 B.n144 10.6151
R752 B.n144 B.n143 10.6151
R753 B.n143 B.n114 10.6151
R754 B.n139 B.n114 10.6151
R755 B.n139 B.n138 10.6151
R756 B.n138 B.n137 10.6151
R757 B.n137 B.n116 10.6151
R758 B.n133 B.n116 10.6151
R759 B.n133 B.n132 10.6151
R760 B.n132 B.n131 10.6151
R761 B.n131 B.n118 10.6151
R762 B.n127 B.n118 10.6151
R763 B.n127 B.n126 10.6151
R764 B.n126 B.n125 10.6151
R765 B.n125 B.n120 10.6151
R766 B.n121 B.n120 10.6151
R767 B.n121 B.n0 10.6151
R768 B.n451 B.n1 10.6151
R769 B.n451 B.n450 10.6151
R770 B.n450 B.n449 10.6151
R771 B.n449 B.n4 10.6151
R772 B.n445 B.n4 10.6151
R773 B.n445 B.n444 10.6151
R774 B.n444 B.n443 10.6151
R775 B.n443 B.n6 10.6151
R776 B.n439 B.n6 10.6151
R777 B.n439 B.n438 10.6151
R778 B.n438 B.n437 10.6151
R779 B.n437 B.n8 10.6151
R780 B.n433 B.n8 10.6151
R781 B.n433 B.n432 10.6151
R782 B.n432 B.n431 10.6151
R783 B.n431 B.n10 10.6151
R784 B.n427 B.n10 10.6151
R785 B.n427 B.n426 10.6151
R786 B.n426 B.n425 10.6151
R787 B.n425 B.n12 10.6151
R788 B.n421 B.n12 10.6151
R789 B.n421 B.n420 10.6151
R790 B.n420 B.n419 10.6151
R791 B.n419 B.n14 10.6151
R792 B.n415 B.n14 10.6151
R793 B.n415 B.n414 10.6151
R794 B.n414 B.n413 10.6151
R795 B.n413 B.n16 10.6151
R796 B.n409 B.n16 10.6151
R797 B.n409 B.n408 10.6151
R798 B.n408 B.n407 10.6151
R799 B.n407 B.n18 10.6151
R800 B.n379 B.n378 9.52245
R801 B.n361 B.n36 9.52245
R802 B.n193 B.n96 9.52245
R803 B.n211 B.n210 9.52245
R804 B.n455 B.n0 2.81026
R805 B.n455 B.n1 2.81026
R806 B.n378 B.n377 1.09318
R807 B.n364 B.n36 1.09318
R808 B.n196 B.n96 1.09318
R809 B.n210 B.n209 1.09318
R810 VN.n18 VN.n17 172.499
R811 VN.n37 VN.n36 172.499
R812 VN.n35 VN.n19 161.3
R813 VN.n34 VN.n33 161.3
R814 VN.n32 VN.n20 161.3
R815 VN.n31 VN.n30 161.3
R816 VN.n29 VN.n21 161.3
R817 VN.n28 VN.n27 161.3
R818 VN.n26 VN.n23 161.3
R819 VN.n16 VN.n0 161.3
R820 VN.n15 VN.n14 161.3
R821 VN.n13 VN.n1 161.3
R822 VN.n12 VN.n11 161.3
R823 VN.n9 VN.n2 161.3
R824 VN.n8 VN.n7 161.3
R825 VN.n6 VN.n3 161.3
R826 VN.n5 VN.t3 94.5391
R827 VN.n25 VN.t0 94.5391
R828 VN.n4 VN.t7 64.9812
R829 VN.n10 VN.t6 64.9812
R830 VN.n17 VN.t2 64.9812
R831 VN.n24 VN.t4 64.9812
R832 VN.n22 VN.t1 64.9812
R833 VN.n36 VN.t5 64.9812
R834 VN.n5 VN.n4 60.6301
R835 VN.n25 VN.n24 60.6301
R836 VN.n9 VN.n8 56.4773
R837 VN.n29 VN.n28 56.4773
R838 VN.n15 VN.n1 47.2268
R839 VN.n34 VN.n20 47.2268
R840 VN VN.n37 39.0327
R841 VN.n16 VN.n15 33.5944
R842 VN.n35 VN.n34 33.5944
R843 VN.n26 VN.n25 27.0891
R844 VN.n6 VN.n5 27.0891
R845 VN.n8 VN.n3 24.3439
R846 VN.n11 VN.n9 24.3439
R847 VN.n28 VN.n23 24.3439
R848 VN.n30 VN.n29 24.3439
R849 VN.n10 VN.n1 19.9621
R850 VN.n22 VN.n20 19.9621
R851 VN.n17 VN.n16 13.146
R852 VN.n36 VN.n35 13.146
R853 VN.n4 VN.n3 4.38232
R854 VN.n11 VN.n10 4.38232
R855 VN.n24 VN.n23 4.38232
R856 VN.n30 VN.n22 4.38232
R857 VN.n37 VN.n19 0.189894
R858 VN.n33 VN.n19 0.189894
R859 VN.n33 VN.n32 0.189894
R860 VN.n32 VN.n31 0.189894
R861 VN.n31 VN.n21 0.189894
R862 VN.n27 VN.n21 0.189894
R863 VN.n27 VN.n26 0.189894
R864 VN.n7 VN.n6 0.189894
R865 VN.n7 VN.n2 0.189894
R866 VN.n12 VN.n2 0.189894
R867 VN.n13 VN.n12 0.189894
R868 VN.n14 VN.n13 0.189894
R869 VN.n14 VN.n0 0.189894
R870 VN.n18 VN.n0 0.189894
R871 VN VN.n18 0.0516364
R872 VDD2.n2 VDD2.n1 123.68
R873 VDD2.n2 VDD2.n0 123.68
R874 VDD2 VDD2.n5 123.677
R875 VDD2.n4 VDD2.n3 123.011
R876 VDD2.n4 VDD2.n2 33.3705
R877 VDD2.n5 VDD2.t3 8.93044
R878 VDD2.n5 VDD2.t7 8.93044
R879 VDD2.n3 VDD2.t2 8.93044
R880 VDD2.n3 VDD2.t6 8.93044
R881 VDD2.n1 VDD2.t1 8.93044
R882 VDD2.n1 VDD2.t5 8.93044
R883 VDD2.n0 VDD2.t4 8.93044
R884 VDD2.n0 VDD2.t0 8.93044
R885 VDD2 VDD2.n4 0.782828
C0 VDD1 VTAIL 4.56211f
C1 VDD1 B 1.04297f
C2 VP w_n2650_n1696# 5.23699f
C3 VN VP 4.595799f
C4 VTAIL w_n2650_n1696# 2.14334f
C5 VN VTAIL 2.96115f
C6 VDD2 VDD1 1.15064f
C7 B w_n2650_n1696# 5.87279f
C8 VN B 0.845047f
C9 VDD2 w_n2650_n1696# 1.37f
C10 VN VDD2 2.51246f
C11 VP VTAIL 2.97526f
C12 VP B 1.40864f
C13 B VTAIL 1.80952f
C14 VDD1 w_n2650_n1696# 1.3082f
C15 VN VDD1 0.153374f
C16 VDD2 VP 0.391069f
C17 VDD2 VTAIL 4.60815f
C18 VN w_n2650_n1696# 4.89801f
C19 VDD2 B 1.09989f
C20 VDD1 VP 2.74882f
C21 VDD2 VSUBS 1.115773f
C22 VDD1 VSUBS 1.544475f
C23 VTAIL VSUBS 0.4865f
C24 VN VSUBS 4.84672f
C25 VP VSUBS 1.82528f
C26 B VSUBS 2.750167f
C27 w_n2650_n1696# VSUBS 56.699398f
C28 VDD2.t4 VSUBS 0.071299f
C29 VDD2.t0 VSUBS 0.071299f
C30 VDD2.n0 VSUBS 0.405666f
C31 VDD2.t1 VSUBS 0.071299f
C32 VDD2.t5 VSUBS 0.071299f
C33 VDD2.n1 VSUBS 0.405666f
C34 VDD2.n2 VSUBS 2.30397f
C35 VDD2.t2 VSUBS 0.071299f
C36 VDD2.t6 VSUBS 0.071299f
C37 VDD2.n3 VSUBS 0.402863f
C38 VDD2.n4 VSUBS 1.97542f
C39 VDD2.t3 VSUBS 0.071299f
C40 VDD2.t7 VSUBS 0.071299f
C41 VDD2.n5 VSUBS 0.405647f
C42 VN.n0 VSUBS 0.054356f
C43 VN.t2 VSUBS 0.678637f
C44 VN.n1 VSUBS 0.094227f
C45 VN.n2 VSUBS 0.054356f
C46 VN.n3 VSUBS 0.060593f
C47 VN.t3 VSUBS 0.82891f
C48 VN.t7 VSUBS 0.678637f
C49 VN.n4 VSUBS 0.376288f
C50 VN.n5 VSUBS 0.411324f
C51 VN.n6 VSUBS 0.289453f
C52 VN.n7 VSUBS 0.054356f
C53 VN.n8 VSUBS 0.079696f
C54 VN.n9 VSUBS 0.079696f
C55 VN.t6 VSUBS 0.678637f
C56 VN.n10 VSUBS 0.299788f
C57 VN.n11 VSUBS 0.060593f
C58 VN.n12 VSUBS 0.054356f
C59 VN.n13 VSUBS 0.054356f
C60 VN.n14 VSUBS 0.054356f
C61 VN.n15 VSUBS 0.047533f
C62 VN.n16 VSUBS 0.087272f
C63 VN.n17 VSUBS 0.406274f
C64 VN.n18 VSUBS 0.049517f
C65 VN.n19 VSUBS 0.054356f
C66 VN.t5 VSUBS 0.678637f
C67 VN.n20 VSUBS 0.094227f
C68 VN.n21 VSUBS 0.054356f
C69 VN.t1 VSUBS 0.678637f
C70 VN.n22 VSUBS 0.299788f
C71 VN.n23 VSUBS 0.060593f
C72 VN.t0 VSUBS 0.82891f
C73 VN.t4 VSUBS 0.678637f
C74 VN.n24 VSUBS 0.376288f
C75 VN.n25 VSUBS 0.411324f
C76 VN.n26 VSUBS 0.289453f
C77 VN.n27 VSUBS 0.054356f
C78 VN.n28 VSUBS 0.079696f
C79 VN.n29 VSUBS 0.079696f
C80 VN.n30 VSUBS 0.060593f
C81 VN.n31 VSUBS 0.054356f
C82 VN.n32 VSUBS 0.054356f
C83 VN.n33 VSUBS 0.054356f
C84 VN.n34 VSUBS 0.047533f
C85 VN.n35 VSUBS 0.087272f
C86 VN.n36 VSUBS 0.406274f
C87 VN.n37 VSUBS 1.98877f
C88 B.n0 VSUBS 0.00469f
C89 B.n1 VSUBS 0.00469f
C90 B.n2 VSUBS 0.007417f
C91 B.n3 VSUBS 0.007417f
C92 B.n4 VSUBS 0.007417f
C93 B.n5 VSUBS 0.007417f
C94 B.n6 VSUBS 0.007417f
C95 B.n7 VSUBS 0.007417f
C96 B.n8 VSUBS 0.007417f
C97 B.n9 VSUBS 0.007417f
C98 B.n10 VSUBS 0.007417f
C99 B.n11 VSUBS 0.007417f
C100 B.n12 VSUBS 0.007417f
C101 B.n13 VSUBS 0.007417f
C102 B.n14 VSUBS 0.007417f
C103 B.n15 VSUBS 0.007417f
C104 B.n16 VSUBS 0.007417f
C105 B.n17 VSUBS 0.007417f
C106 B.n18 VSUBS 0.015447f
C107 B.n19 VSUBS 0.007417f
C108 B.n20 VSUBS 0.007417f
C109 B.n21 VSUBS 0.007417f
C110 B.n22 VSUBS 0.007417f
C111 B.n23 VSUBS 0.007417f
C112 B.n24 VSUBS 0.007417f
C113 B.n25 VSUBS 0.007417f
C114 B.n26 VSUBS 0.007417f
C115 B.n27 VSUBS 0.007417f
C116 B.t5 VSUBS 0.098369f
C117 B.t4 VSUBS 0.109497f
C118 B.t3 VSUBS 0.24435f
C119 B.n28 VSUBS 0.08232f
C120 B.n29 VSUBS 0.066393f
C121 B.n30 VSUBS 0.007417f
C122 B.n31 VSUBS 0.007417f
C123 B.n32 VSUBS 0.007417f
C124 B.n33 VSUBS 0.007417f
C125 B.t8 VSUBS 0.098369f
C126 B.t7 VSUBS 0.109497f
C127 B.t6 VSUBS 0.244379f
C128 B.n34 VSUBS 0.08229f
C129 B.n35 VSUBS 0.066393f
C130 B.n36 VSUBS 0.017184f
C131 B.n37 VSUBS 0.007417f
C132 B.n38 VSUBS 0.007417f
C133 B.n39 VSUBS 0.007417f
C134 B.n40 VSUBS 0.007417f
C135 B.n41 VSUBS 0.007417f
C136 B.n42 VSUBS 0.007417f
C137 B.n43 VSUBS 0.007417f
C138 B.n44 VSUBS 0.007417f
C139 B.n45 VSUBS 0.015447f
C140 B.n46 VSUBS 0.007417f
C141 B.n47 VSUBS 0.007417f
C142 B.n48 VSUBS 0.007417f
C143 B.n49 VSUBS 0.007417f
C144 B.n50 VSUBS 0.007417f
C145 B.n51 VSUBS 0.007417f
C146 B.n52 VSUBS 0.007417f
C147 B.n53 VSUBS 0.007417f
C148 B.n54 VSUBS 0.007417f
C149 B.n55 VSUBS 0.007417f
C150 B.n56 VSUBS 0.007417f
C151 B.n57 VSUBS 0.007417f
C152 B.n58 VSUBS 0.007417f
C153 B.n59 VSUBS 0.007417f
C154 B.n60 VSUBS 0.007417f
C155 B.n61 VSUBS 0.007417f
C156 B.n62 VSUBS 0.007417f
C157 B.n63 VSUBS 0.007417f
C158 B.n64 VSUBS 0.007417f
C159 B.n65 VSUBS 0.007417f
C160 B.n66 VSUBS 0.007417f
C161 B.n67 VSUBS 0.007417f
C162 B.n68 VSUBS 0.007417f
C163 B.n69 VSUBS 0.007417f
C164 B.n70 VSUBS 0.007417f
C165 B.n71 VSUBS 0.007417f
C166 B.n72 VSUBS 0.007417f
C167 B.n73 VSUBS 0.007417f
C168 B.n74 VSUBS 0.007417f
C169 B.n75 VSUBS 0.007417f
C170 B.n76 VSUBS 0.007417f
C171 B.n77 VSUBS 0.007417f
C172 B.n78 VSUBS 0.015447f
C173 B.n79 VSUBS 0.007417f
C174 B.n80 VSUBS 0.007417f
C175 B.n81 VSUBS 0.007417f
C176 B.n82 VSUBS 0.007417f
C177 B.n83 VSUBS 0.007417f
C178 B.n84 VSUBS 0.007417f
C179 B.n85 VSUBS 0.007417f
C180 B.n86 VSUBS 0.007417f
C181 B.n87 VSUBS 0.007417f
C182 B.t1 VSUBS 0.098369f
C183 B.t2 VSUBS 0.109497f
C184 B.t0 VSUBS 0.244379f
C185 B.n88 VSUBS 0.08229f
C186 B.n89 VSUBS 0.066393f
C187 B.n90 VSUBS 0.007417f
C188 B.n91 VSUBS 0.007417f
C189 B.n92 VSUBS 0.007417f
C190 B.n93 VSUBS 0.007417f
C191 B.t10 VSUBS 0.098369f
C192 B.t11 VSUBS 0.109497f
C193 B.t9 VSUBS 0.24435f
C194 B.n94 VSUBS 0.08232f
C195 B.n95 VSUBS 0.066393f
C196 B.n96 VSUBS 0.017184f
C197 B.n97 VSUBS 0.007417f
C198 B.n98 VSUBS 0.007417f
C199 B.n99 VSUBS 0.007417f
C200 B.n100 VSUBS 0.007417f
C201 B.n101 VSUBS 0.007417f
C202 B.n102 VSUBS 0.007417f
C203 B.n103 VSUBS 0.007417f
C204 B.n104 VSUBS 0.007417f
C205 B.n105 VSUBS 0.015447f
C206 B.n106 VSUBS 0.007417f
C207 B.n107 VSUBS 0.007417f
C208 B.n108 VSUBS 0.007417f
C209 B.n109 VSUBS 0.007417f
C210 B.n110 VSUBS 0.007417f
C211 B.n111 VSUBS 0.007417f
C212 B.n112 VSUBS 0.007417f
C213 B.n113 VSUBS 0.007417f
C214 B.n114 VSUBS 0.007417f
C215 B.n115 VSUBS 0.007417f
C216 B.n116 VSUBS 0.007417f
C217 B.n117 VSUBS 0.007417f
C218 B.n118 VSUBS 0.007417f
C219 B.n119 VSUBS 0.007417f
C220 B.n120 VSUBS 0.007417f
C221 B.n121 VSUBS 0.007417f
C222 B.n122 VSUBS 0.007417f
C223 B.n123 VSUBS 0.007417f
C224 B.n124 VSUBS 0.007417f
C225 B.n125 VSUBS 0.007417f
C226 B.n126 VSUBS 0.007417f
C227 B.n127 VSUBS 0.007417f
C228 B.n128 VSUBS 0.007417f
C229 B.n129 VSUBS 0.007417f
C230 B.n130 VSUBS 0.007417f
C231 B.n131 VSUBS 0.007417f
C232 B.n132 VSUBS 0.007417f
C233 B.n133 VSUBS 0.007417f
C234 B.n134 VSUBS 0.007417f
C235 B.n135 VSUBS 0.007417f
C236 B.n136 VSUBS 0.007417f
C237 B.n137 VSUBS 0.007417f
C238 B.n138 VSUBS 0.007417f
C239 B.n139 VSUBS 0.007417f
C240 B.n140 VSUBS 0.007417f
C241 B.n141 VSUBS 0.007417f
C242 B.n142 VSUBS 0.007417f
C243 B.n143 VSUBS 0.007417f
C244 B.n144 VSUBS 0.007417f
C245 B.n145 VSUBS 0.007417f
C246 B.n146 VSUBS 0.007417f
C247 B.n147 VSUBS 0.007417f
C248 B.n148 VSUBS 0.007417f
C249 B.n149 VSUBS 0.007417f
C250 B.n150 VSUBS 0.007417f
C251 B.n151 VSUBS 0.007417f
C252 B.n152 VSUBS 0.007417f
C253 B.n153 VSUBS 0.007417f
C254 B.n154 VSUBS 0.007417f
C255 B.n155 VSUBS 0.007417f
C256 B.n156 VSUBS 0.007417f
C257 B.n157 VSUBS 0.007417f
C258 B.n158 VSUBS 0.007417f
C259 B.n159 VSUBS 0.007417f
C260 B.n160 VSUBS 0.007417f
C261 B.n161 VSUBS 0.007417f
C262 B.n162 VSUBS 0.007417f
C263 B.n163 VSUBS 0.007417f
C264 B.n164 VSUBS 0.007417f
C265 B.n165 VSUBS 0.007417f
C266 B.n166 VSUBS 0.007417f
C267 B.n167 VSUBS 0.007417f
C268 B.n168 VSUBS 0.015447f
C269 B.n169 VSUBS 0.0164f
C270 B.n170 VSUBS 0.0164f
C271 B.n171 VSUBS 0.007417f
C272 B.n172 VSUBS 0.007417f
C273 B.n173 VSUBS 0.007417f
C274 B.n174 VSUBS 0.007417f
C275 B.n175 VSUBS 0.007417f
C276 B.n176 VSUBS 0.007417f
C277 B.n177 VSUBS 0.007417f
C278 B.n178 VSUBS 0.007417f
C279 B.n179 VSUBS 0.007417f
C280 B.n180 VSUBS 0.007417f
C281 B.n181 VSUBS 0.007417f
C282 B.n182 VSUBS 0.007417f
C283 B.n183 VSUBS 0.007417f
C284 B.n184 VSUBS 0.007417f
C285 B.n185 VSUBS 0.007417f
C286 B.n186 VSUBS 0.007417f
C287 B.n187 VSUBS 0.007417f
C288 B.n188 VSUBS 0.007417f
C289 B.n189 VSUBS 0.007417f
C290 B.n190 VSUBS 0.007417f
C291 B.n191 VSUBS 0.007417f
C292 B.n192 VSUBS 0.007417f
C293 B.n193 VSUBS 0.007035f
C294 B.n194 VSUBS 0.007417f
C295 B.n195 VSUBS 0.007417f
C296 B.n196 VSUBS 0.00409f
C297 B.n197 VSUBS 0.007417f
C298 B.n198 VSUBS 0.007417f
C299 B.n199 VSUBS 0.007417f
C300 B.n200 VSUBS 0.007417f
C301 B.n201 VSUBS 0.007417f
C302 B.n202 VSUBS 0.007417f
C303 B.n203 VSUBS 0.007417f
C304 B.n204 VSUBS 0.007417f
C305 B.n205 VSUBS 0.007417f
C306 B.n206 VSUBS 0.007417f
C307 B.n207 VSUBS 0.007417f
C308 B.n208 VSUBS 0.007417f
C309 B.n209 VSUBS 0.00409f
C310 B.n210 VSUBS 0.017184f
C311 B.n211 VSUBS 0.007035f
C312 B.n212 VSUBS 0.007417f
C313 B.n213 VSUBS 0.007417f
C314 B.n214 VSUBS 0.007417f
C315 B.n215 VSUBS 0.007417f
C316 B.n216 VSUBS 0.007417f
C317 B.n217 VSUBS 0.007417f
C318 B.n218 VSUBS 0.007417f
C319 B.n219 VSUBS 0.007417f
C320 B.n220 VSUBS 0.007417f
C321 B.n221 VSUBS 0.007417f
C322 B.n222 VSUBS 0.007417f
C323 B.n223 VSUBS 0.007417f
C324 B.n224 VSUBS 0.007417f
C325 B.n225 VSUBS 0.007417f
C326 B.n226 VSUBS 0.007417f
C327 B.n227 VSUBS 0.007417f
C328 B.n228 VSUBS 0.007417f
C329 B.n229 VSUBS 0.007417f
C330 B.n230 VSUBS 0.007417f
C331 B.n231 VSUBS 0.007417f
C332 B.n232 VSUBS 0.007417f
C333 B.n233 VSUBS 0.007417f
C334 B.n234 VSUBS 0.007417f
C335 B.n235 VSUBS 0.0164f
C336 B.n236 VSUBS 0.0164f
C337 B.n237 VSUBS 0.015447f
C338 B.n238 VSUBS 0.007417f
C339 B.n239 VSUBS 0.007417f
C340 B.n240 VSUBS 0.007417f
C341 B.n241 VSUBS 0.007417f
C342 B.n242 VSUBS 0.007417f
C343 B.n243 VSUBS 0.007417f
C344 B.n244 VSUBS 0.007417f
C345 B.n245 VSUBS 0.007417f
C346 B.n246 VSUBS 0.007417f
C347 B.n247 VSUBS 0.007417f
C348 B.n248 VSUBS 0.007417f
C349 B.n249 VSUBS 0.007417f
C350 B.n250 VSUBS 0.007417f
C351 B.n251 VSUBS 0.007417f
C352 B.n252 VSUBS 0.007417f
C353 B.n253 VSUBS 0.007417f
C354 B.n254 VSUBS 0.007417f
C355 B.n255 VSUBS 0.007417f
C356 B.n256 VSUBS 0.007417f
C357 B.n257 VSUBS 0.007417f
C358 B.n258 VSUBS 0.007417f
C359 B.n259 VSUBS 0.007417f
C360 B.n260 VSUBS 0.007417f
C361 B.n261 VSUBS 0.007417f
C362 B.n262 VSUBS 0.007417f
C363 B.n263 VSUBS 0.007417f
C364 B.n264 VSUBS 0.007417f
C365 B.n265 VSUBS 0.007417f
C366 B.n266 VSUBS 0.007417f
C367 B.n267 VSUBS 0.007417f
C368 B.n268 VSUBS 0.007417f
C369 B.n269 VSUBS 0.007417f
C370 B.n270 VSUBS 0.007417f
C371 B.n271 VSUBS 0.007417f
C372 B.n272 VSUBS 0.007417f
C373 B.n273 VSUBS 0.007417f
C374 B.n274 VSUBS 0.007417f
C375 B.n275 VSUBS 0.007417f
C376 B.n276 VSUBS 0.007417f
C377 B.n277 VSUBS 0.007417f
C378 B.n278 VSUBS 0.007417f
C379 B.n279 VSUBS 0.007417f
C380 B.n280 VSUBS 0.007417f
C381 B.n281 VSUBS 0.007417f
C382 B.n282 VSUBS 0.007417f
C383 B.n283 VSUBS 0.007417f
C384 B.n284 VSUBS 0.007417f
C385 B.n285 VSUBS 0.007417f
C386 B.n286 VSUBS 0.007417f
C387 B.n287 VSUBS 0.007417f
C388 B.n288 VSUBS 0.007417f
C389 B.n289 VSUBS 0.007417f
C390 B.n290 VSUBS 0.007417f
C391 B.n291 VSUBS 0.007417f
C392 B.n292 VSUBS 0.007417f
C393 B.n293 VSUBS 0.007417f
C394 B.n294 VSUBS 0.007417f
C395 B.n295 VSUBS 0.007417f
C396 B.n296 VSUBS 0.007417f
C397 B.n297 VSUBS 0.007417f
C398 B.n298 VSUBS 0.007417f
C399 B.n299 VSUBS 0.007417f
C400 B.n300 VSUBS 0.007417f
C401 B.n301 VSUBS 0.007417f
C402 B.n302 VSUBS 0.007417f
C403 B.n303 VSUBS 0.007417f
C404 B.n304 VSUBS 0.007417f
C405 B.n305 VSUBS 0.007417f
C406 B.n306 VSUBS 0.007417f
C407 B.n307 VSUBS 0.007417f
C408 B.n308 VSUBS 0.007417f
C409 B.n309 VSUBS 0.007417f
C410 B.n310 VSUBS 0.007417f
C411 B.n311 VSUBS 0.007417f
C412 B.n312 VSUBS 0.007417f
C413 B.n313 VSUBS 0.007417f
C414 B.n314 VSUBS 0.007417f
C415 B.n315 VSUBS 0.007417f
C416 B.n316 VSUBS 0.007417f
C417 B.n317 VSUBS 0.007417f
C418 B.n318 VSUBS 0.007417f
C419 B.n319 VSUBS 0.007417f
C420 B.n320 VSUBS 0.007417f
C421 B.n321 VSUBS 0.007417f
C422 B.n322 VSUBS 0.007417f
C423 B.n323 VSUBS 0.007417f
C424 B.n324 VSUBS 0.007417f
C425 B.n325 VSUBS 0.007417f
C426 B.n326 VSUBS 0.007417f
C427 B.n327 VSUBS 0.007417f
C428 B.n328 VSUBS 0.007417f
C429 B.n329 VSUBS 0.007417f
C430 B.n330 VSUBS 0.007417f
C431 B.n331 VSUBS 0.007417f
C432 B.n332 VSUBS 0.007417f
C433 B.n333 VSUBS 0.007417f
C434 B.n334 VSUBS 0.007417f
C435 B.n335 VSUBS 0.007417f
C436 B.n336 VSUBS 0.016449f
C437 B.n337 VSUBS 0.015398f
C438 B.n338 VSUBS 0.0164f
C439 B.n339 VSUBS 0.007417f
C440 B.n340 VSUBS 0.007417f
C441 B.n341 VSUBS 0.007417f
C442 B.n342 VSUBS 0.007417f
C443 B.n343 VSUBS 0.007417f
C444 B.n344 VSUBS 0.007417f
C445 B.n345 VSUBS 0.007417f
C446 B.n346 VSUBS 0.007417f
C447 B.n347 VSUBS 0.007417f
C448 B.n348 VSUBS 0.007417f
C449 B.n349 VSUBS 0.007417f
C450 B.n350 VSUBS 0.007417f
C451 B.n351 VSUBS 0.007417f
C452 B.n352 VSUBS 0.007417f
C453 B.n353 VSUBS 0.007417f
C454 B.n354 VSUBS 0.007417f
C455 B.n355 VSUBS 0.007417f
C456 B.n356 VSUBS 0.007417f
C457 B.n357 VSUBS 0.007417f
C458 B.n358 VSUBS 0.007417f
C459 B.n359 VSUBS 0.007417f
C460 B.n360 VSUBS 0.007417f
C461 B.n361 VSUBS 0.007035f
C462 B.n362 VSUBS 0.007417f
C463 B.n363 VSUBS 0.007417f
C464 B.n364 VSUBS 0.00409f
C465 B.n365 VSUBS 0.007417f
C466 B.n366 VSUBS 0.007417f
C467 B.n367 VSUBS 0.007417f
C468 B.n368 VSUBS 0.007417f
C469 B.n369 VSUBS 0.007417f
C470 B.n370 VSUBS 0.007417f
C471 B.n371 VSUBS 0.007417f
C472 B.n372 VSUBS 0.007417f
C473 B.n373 VSUBS 0.007417f
C474 B.n374 VSUBS 0.007417f
C475 B.n375 VSUBS 0.007417f
C476 B.n376 VSUBS 0.007417f
C477 B.n377 VSUBS 0.00409f
C478 B.n378 VSUBS 0.017184f
C479 B.n379 VSUBS 0.007035f
C480 B.n380 VSUBS 0.007417f
C481 B.n381 VSUBS 0.007417f
C482 B.n382 VSUBS 0.007417f
C483 B.n383 VSUBS 0.007417f
C484 B.n384 VSUBS 0.007417f
C485 B.n385 VSUBS 0.007417f
C486 B.n386 VSUBS 0.007417f
C487 B.n387 VSUBS 0.007417f
C488 B.n388 VSUBS 0.007417f
C489 B.n389 VSUBS 0.007417f
C490 B.n390 VSUBS 0.007417f
C491 B.n391 VSUBS 0.007417f
C492 B.n392 VSUBS 0.007417f
C493 B.n393 VSUBS 0.007417f
C494 B.n394 VSUBS 0.007417f
C495 B.n395 VSUBS 0.007417f
C496 B.n396 VSUBS 0.007417f
C497 B.n397 VSUBS 0.007417f
C498 B.n398 VSUBS 0.007417f
C499 B.n399 VSUBS 0.007417f
C500 B.n400 VSUBS 0.007417f
C501 B.n401 VSUBS 0.007417f
C502 B.n402 VSUBS 0.007417f
C503 B.n403 VSUBS 0.0164f
C504 B.n404 VSUBS 0.0164f
C505 B.n405 VSUBS 0.015447f
C506 B.n406 VSUBS 0.007417f
C507 B.n407 VSUBS 0.007417f
C508 B.n408 VSUBS 0.007417f
C509 B.n409 VSUBS 0.007417f
C510 B.n410 VSUBS 0.007417f
C511 B.n411 VSUBS 0.007417f
C512 B.n412 VSUBS 0.007417f
C513 B.n413 VSUBS 0.007417f
C514 B.n414 VSUBS 0.007417f
C515 B.n415 VSUBS 0.007417f
C516 B.n416 VSUBS 0.007417f
C517 B.n417 VSUBS 0.007417f
C518 B.n418 VSUBS 0.007417f
C519 B.n419 VSUBS 0.007417f
C520 B.n420 VSUBS 0.007417f
C521 B.n421 VSUBS 0.007417f
C522 B.n422 VSUBS 0.007417f
C523 B.n423 VSUBS 0.007417f
C524 B.n424 VSUBS 0.007417f
C525 B.n425 VSUBS 0.007417f
C526 B.n426 VSUBS 0.007417f
C527 B.n427 VSUBS 0.007417f
C528 B.n428 VSUBS 0.007417f
C529 B.n429 VSUBS 0.007417f
C530 B.n430 VSUBS 0.007417f
C531 B.n431 VSUBS 0.007417f
C532 B.n432 VSUBS 0.007417f
C533 B.n433 VSUBS 0.007417f
C534 B.n434 VSUBS 0.007417f
C535 B.n435 VSUBS 0.007417f
C536 B.n436 VSUBS 0.007417f
C537 B.n437 VSUBS 0.007417f
C538 B.n438 VSUBS 0.007417f
C539 B.n439 VSUBS 0.007417f
C540 B.n440 VSUBS 0.007417f
C541 B.n441 VSUBS 0.007417f
C542 B.n442 VSUBS 0.007417f
C543 B.n443 VSUBS 0.007417f
C544 B.n444 VSUBS 0.007417f
C545 B.n445 VSUBS 0.007417f
C546 B.n446 VSUBS 0.007417f
C547 B.n447 VSUBS 0.007417f
C548 B.n448 VSUBS 0.007417f
C549 B.n449 VSUBS 0.007417f
C550 B.n450 VSUBS 0.007417f
C551 B.n451 VSUBS 0.007417f
C552 B.n452 VSUBS 0.007417f
C553 B.n453 VSUBS 0.007417f
C554 B.n454 VSUBS 0.007417f
C555 B.n455 VSUBS 0.016794f
C556 VDD1.t6 VSUBS 0.072374f
C557 VDD1.t1 VSUBS 0.072374f
C558 VDD1.n0 VSUBS 0.412317f
C559 VDD1.t4 VSUBS 0.072374f
C560 VDD1.t3 VSUBS 0.072374f
C561 VDD1.n1 VSUBS 0.411783f
C562 VDD1.t5 VSUBS 0.072374f
C563 VDD1.t7 VSUBS 0.072374f
C564 VDD1.n2 VSUBS 0.411783f
C565 VDD1.n3 VSUBS 2.39216f
C566 VDD1.t0 VSUBS 0.072374f
C567 VDD1.t2 VSUBS 0.072374f
C568 VDD1.n4 VSUBS 0.408936f
C569 VDD1.n5 VSUBS 2.03527f
C570 VTAIL.t2 VSUBS 0.079927f
C571 VTAIL.t7 VSUBS 0.079927f
C572 VTAIL.n0 VSUBS 0.392896f
C573 VTAIL.n1 VSUBS 0.535438f
C574 VTAIL.t3 VSUBS 0.569742f
C575 VTAIL.n2 VSUBS 0.61343f
C576 VTAIL.t14 VSUBS 0.569742f
C577 VTAIL.n3 VSUBS 0.61343f
C578 VTAIL.t10 VSUBS 0.079927f
C579 VTAIL.t15 VSUBS 0.079927f
C580 VTAIL.n4 VSUBS 0.392896f
C581 VTAIL.n5 VSUBS 0.659899f
C582 VTAIL.t8 VSUBS 0.569742f
C583 VTAIL.n6 VSUBS 1.35944f
C584 VTAIL.t5 VSUBS 0.569744f
C585 VTAIL.n7 VSUBS 1.35944f
C586 VTAIL.t6 VSUBS 0.079927f
C587 VTAIL.t0 VSUBS 0.079927f
C588 VTAIL.n8 VSUBS 0.392898f
C589 VTAIL.n9 VSUBS 0.659897f
C590 VTAIL.t4 VSUBS 0.569744f
C591 VTAIL.n10 VSUBS 0.613427f
C592 VTAIL.t13 VSUBS 0.569744f
C593 VTAIL.n11 VSUBS 0.613427f
C594 VTAIL.t11 VSUBS 0.079927f
C595 VTAIL.t12 VSUBS 0.079927f
C596 VTAIL.n12 VSUBS 0.392898f
C597 VTAIL.n13 VSUBS 0.659897f
C598 VTAIL.t9 VSUBS 0.569742f
C599 VTAIL.n14 VSUBS 1.35944f
C600 VTAIL.t1 VSUBS 0.569742f
C601 VTAIL.n15 VSUBS 1.35423f
C602 VP.n0 VSUBS 0.056456f
C603 VP.t0 VSUBS 0.704848f
C604 VP.n1 VSUBS 0.097866f
C605 VP.n2 VSUBS 0.056456f
C606 VP.n3 VSUBS 0.062933f
C607 VP.n4 VSUBS 0.056456f
C608 VP.t3 VSUBS 0.704848f
C609 VP.n5 VSUBS 0.421966f
C610 VP.n6 VSUBS 0.056456f
C611 VP.t5 VSUBS 0.704848f
C612 VP.n7 VSUBS 0.097866f
C613 VP.n8 VSUBS 0.056456f
C614 VP.n9 VSUBS 0.062933f
C615 VP.t1 VSUBS 0.860926f
C616 VP.t6 VSUBS 0.704848f
C617 VP.n10 VSUBS 0.390822f
C618 VP.n11 VSUBS 0.427211f
C619 VP.n12 VSUBS 0.300633f
C620 VP.n13 VSUBS 0.056456f
C621 VP.n14 VSUBS 0.082774f
C622 VP.n15 VSUBS 0.082774f
C623 VP.t7 VSUBS 0.704848f
C624 VP.n16 VSUBS 0.311367f
C625 VP.n17 VSUBS 0.062933f
C626 VP.n18 VSUBS 0.056456f
C627 VP.n19 VSUBS 0.056456f
C628 VP.n20 VSUBS 0.056456f
C629 VP.n21 VSUBS 0.049369f
C630 VP.n22 VSUBS 0.090643f
C631 VP.n23 VSUBS 0.421966f
C632 VP.n24 VSUBS 2.02832f
C633 VP.n25 VSUBS 2.08068f
C634 VP.n26 VSUBS 0.056456f
C635 VP.n27 VSUBS 0.090643f
C636 VP.n28 VSUBS 0.049369f
C637 VP.t4 VSUBS 0.704848f
C638 VP.n29 VSUBS 0.311367f
C639 VP.n30 VSUBS 0.097866f
C640 VP.n31 VSUBS 0.056456f
C641 VP.n32 VSUBS 0.056456f
C642 VP.n33 VSUBS 0.056456f
C643 VP.n34 VSUBS 0.082774f
C644 VP.n35 VSUBS 0.082774f
C645 VP.t2 VSUBS 0.704848f
C646 VP.n36 VSUBS 0.311367f
C647 VP.n37 VSUBS 0.062933f
C648 VP.n38 VSUBS 0.056456f
C649 VP.n39 VSUBS 0.056456f
C650 VP.n40 VSUBS 0.056456f
C651 VP.n41 VSUBS 0.049369f
C652 VP.n42 VSUBS 0.090643f
C653 VP.n43 VSUBS 0.421966f
C654 VP.n44 VSUBS 0.051429f
.ends

