* NGSPICE file created from diff_pair_sample_0918.ext - technology: sky130A

.subckt diff_pair_sample_0918 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=0.43
X1 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=7.0707 ps=37.04 w=18.13 l=0.43
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=7.0707 ps=37.04 w=18.13 l=0.43
X3 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=7.0707 ps=37.04 w=18.13 l=0.43
X4 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=0.43
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=0.43
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=0 ps=0 w=18.13 l=0.43
X7 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.0707 pd=37.04 as=7.0707 ps=37.04 w=18.13 l=0.43
R0 B.n95 B.t6 1224.49
R1 B.n93 B.t13 1224.49
R2 B.n405 B.t10 1224.49
R3 B.n411 B.t2 1224.49
R4 B.n757 B.n756 585
R5 B.n758 B.n757 585
R6 B.n351 B.n92 585
R7 B.n350 B.n349 585
R8 B.n348 B.n347 585
R9 B.n346 B.n345 585
R10 B.n344 B.n343 585
R11 B.n342 B.n341 585
R12 B.n340 B.n339 585
R13 B.n338 B.n337 585
R14 B.n336 B.n335 585
R15 B.n334 B.n333 585
R16 B.n332 B.n331 585
R17 B.n330 B.n329 585
R18 B.n328 B.n327 585
R19 B.n326 B.n325 585
R20 B.n324 B.n323 585
R21 B.n322 B.n321 585
R22 B.n320 B.n319 585
R23 B.n318 B.n317 585
R24 B.n316 B.n315 585
R25 B.n314 B.n313 585
R26 B.n312 B.n311 585
R27 B.n310 B.n309 585
R28 B.n308 B.n307 585
R29 B.n306 B.n305 585
R30 B.n304 B.n303 585
R31 B.n302 B.n301 585
R32 B.n300 B.n299 585
R33 B.n298 B.n297 585
R34 B.n296 B.n295 585
R35 B.n294 B.n293 585
R36 B.n292 B.n291 585
R37 B.n290 B.n289 585
R38 B.n288 B.n287 585
R39 B.n286 B.n285 585
R40 B.n284 B.n283 585
R41 B.n282 B.n281 585
R42 B.n280 B.n279 585
R43 B.n278 B.n277 585
R44 B.n276 B.n275 585
R45 B.n274 B.n273 585
R46 B.n272 B.n271 585
R47 B.n270 B.n269 585
R48 B.n268 B.n267 585
R49 B.n266 B.n265 585
R50 B.n264 B.n263 585
R51 B.n262 B.n261 585
R52 B.n260 B.n259 585
R53 B.n258 B.n257 585
R54 B.n256 B.n255 585
R55 B.n254 B.n253 585
R56 B.n252 B.n251 585
R57 B.n250 B.n249 585
R58 B.n248 B.n247 585
R59 B.n246 B.n245 585
R60 B.n244 B.n243 585
R61 B.n242 B.n241 585
R62 B.n240 B.n239 585
R63 B.n238 B.n237 585
R64 B.n236 B.n235 585
R65 B.n233 B.n232 585
R66 B.n231 B.n230 585
R67 B.n229 B.n228 585
R68 B.n227 B.n226 585
R69 B.n225 B.n224 585
R70 B.n223 B.n222 585
R71 B.n221 B.n220 585
R72 B.n219 B.n218 585
R73 B.n217 B.n216 585
R74 B.n215 B.n214 585
R75 B.n213 B.n212 585
R76 B.n211 B.n210 585
R77 B.n209 B.n208 585
R78 B.n207 B.n206 585
R79 B.n205 B.n204 585
R80 B.n203 B.n202 585
R81 B.n201 B.n200 585
R82 B.n199 B.n198 585
R83 B.n197 B.n196 585
R84 B.n195 B.n194 585
R85 B.n193 B.n192 585
R86 B.n191 B.n190 585
R87 B.n189 B.n188 585
R88 B.n187 B.n186 585
R89 B.n185 B.n184 585
R90 B.n183 B.n182 585
R91 B.n181 B.n180 585
R92 B.n179 B.n178 585
R93 B.n177 B.n176 585
R94 B.n175 B.n174 585
R95 B.n173 B.n172 585
R96 B.n171 B.n170 585
R97 B.n169 B.n168 585
R98 B.n167 B.n166 585
R99 B.n165 B.n164 585
R100 B.n163 B.n162 585
R101 B.n161 B.n160 585
R102 B.n159 B.n158 585
R103 B.n157 B.n156 585
R104 B.n155 B.n154 585
R105 B.n153 B.n152 585
R106 B.n151 B.n150 585
R107 B.n149 B.n148 585
R108 B.n147 B.n146 585
R109 B.n145 B.n144 585
R110 B.n143 B.n142 585
R111 B.n141 B.n140 585
R112 B.n139 B.n138 585
R113 B.n137 B.n136 585
R114 B.n135 B.n134 585
R115 B.n133 B.n132 585
R116 B.n131 B.n130 585
R117 B.n129 B.n128 585
R118 B.n127 B.n126 585
R119 B.n125 B.n124 585
R120 B.n123 B.n122 585
R121 B.n121 B.n120 585
R122 B.n119 B.n118 585
R123 B.n117 B.n116 585
R124 B.n115 B.n114 585
R125 B.n113 B.n112 585
R126 B.n111 B.n110 585
R127 B.n109 B.n108 585
R128 B.n107 B.n106 585
R129 B.n105 B.n104 585
R130 B.n103 B.n102 585
R131 B.n101 B.n100 585
R132 B.n99 B.n98 585
R133 B.n26 B.n25 585
R134 B.n755 B.n27 585
R135 B.n759 B.n27 585
R136 B.n754 B.n753 585
R137 B.n753 B.n23 585
R138 B.n752 B.n22 585
R139 B.n765 B.n22 585
R140 B.n751 B.n21 585
R141 B.n766 B.n21 585
R142 B.n750 B.n20 585
R143 B.n767 B.n20 585
R144 B.n749 B.n748 585
R145 B.n748 B.n16 585
R146 B.n747 B.n15 585
R147 B.n773 B.n15 585
R148 B.n746 B.n14 585
R149 B.n774 B.n14 585
R150 B.n745 B.n13 585
R151 B.n775 B.n13 585
R152 B.n744 B.n743 585
R153 B.n743 B.n12 585
R154 B.n742 B.n741 585
R155 B.n742 B.n8 585
R156 B.n740 B.n7 585
R157 B.n782 B.n7 585
R158 B.n739 B.n6 585
R159 B.n783 B.n6 585
R160 B.n738 B.n5 585
R161 B.n784 B.n5 585
R162 B.n737 B.n736 585
R163 B.n736 B.n4 585
R164 B.n735 B.n352 585
R165 B.n735 B.n734 585
R166 B.n724 B.n353 585
R167 B.n727 B.n353 585
R168 B.n726 B.n725 585
R169 B.n728 B.n726 585
R170 B.n723 B.n358 585
R171 B.n358 B.n357 585
R172 B.n722 B.n721 585
R173 B.n721 B.n720 585
R174 B.n360 B.n359 585
R175 B.n361 B.n360 585
R176 B.n713 B.n712 585
R177 B.n714 B.n713 585
R178 B.n711 B.n366 585
R179 B.n366 B.n365 585
R180 B.n710 B.n709 585
R181 B.n709 B.n708 585
R182 B.n368 B.n367 585
R183 B.n369 B.n368 585
R184 B.n701 B.n700 585
R185 B.n702 B.n701 585
R186 B.n372 B.n371 585
R187 B.n444 B.n442 585
R188 B.n445 B.n441 585
R189 B.n445 B.n373 585
R190 B.n448 B.n447 585
R191 B.n449 B.n440 585
R192 B.n451 B.n450 585
R193 B.n453 B.n439 585
R194 B.n456 B.n455 585
R195 B.n457 B.n438 585
R196 B.n459 B.n458 585
R197 B.n461 B.n437 585
R198 B.n464 B.n463 585
R199 B.n465 B.n436 585
R200 B.n467 B.n466 585
R201 B.n469 B.n435 585
R202 B.n472 B.n471 585
R203 B.n473 B.n434 585
R204 B.n475 B.n474 585
R205 B.n477 B.n433 585
R206 B.n480 B.n479 585
R207 B.n481 B.n432 585
R208 B.n483 B.n482 585
R209 B.n485 B.n431 585
R210 B.n488 B.n487 585
R211 B.n489 B.n430 585
R212 B.n491 B.n490 585
R213 B.n493 B.n429 585
R214 B.n496 B.n495 585
R215 B.n497 B.n428 585
R216 B.n499 B.n498 585
R217 B.n501 B.n427 585
R218 B.n504 B.n503 585
R219 B.n505 B.n426 585
R220 B.n507 B.n506 585
R221 B.n509 B.n425 585
R222 B.n512 B.n511 585
R223 B.n513 B.n424 585
R224 B.n515 B.n514 585
R225 B.n517 B.n423 585
R226 B.n520 B.n519 585
R227 B.n521 B.n422 585
R228 B.n523 B.n522 585
R229 B.n525 B.n421 585
R230 B.n528 B.n527 585
R231 B.n529 B.n420 585
R232 B.n531 B.n530 585
R233 B.n533 B.n419 585
R234 B.n536 B.n535 585
R235 B.n537 B.n418 585
R236 B.n539 B.n538 585
R237 B.n541 B.n417 585
R238 B.n544 B.n543 585
R239 B.n545 B.n416 585
R240 B.n547 B.n546 585
R241 B.n549 B.n415 585
R242 B.n552 B.n551 585
R243 B.n553 B.n414 585
R244 B.n555 B.n554 585
R245 B.n557 B.n413 585
R246 B.n560 B.n559 585
R247 B.n562 B.n410 585
R248 B.n564 B.n563 585
R249 B.n566 B.n409 585
R250 B.n569 B.n568 585
R251 B.n570 B.n408 585
R252 B.n572 B.n571 585
R253 B.n574 B.n407 585
R254 B.n577 B.n576 585
R255 B.n578 B.n404 585
R256 B.n581 B.n580 585
R257 B.n583 B.n403 585
R258 B.n586 B.n585 585
R259 B.n587 B.n402 585
R260 B.n589 B.n588 585
R261 B.n591 B.n401 585
R262 B.n594 B.n593 585
R263 B.n595 B.n400 585
R264 B.n597 B.n596 585
R265 B.n599 B.n399 585
R266 B.n602 B.n601 585
R267 B.n603 B.n398 585
R268 B.n605 B.n604 585
R269 B.n607 B.n397 585
R270 B.n610 B.n609 585
R271 B.n611 B.n396 585
R272 B.n613 B.n612 585
R273 B.n615 B.n395 585
R274 B.n618 B.n617 585
R275 B.n619 B.n394 585
R276 B.n621 B.n620 585
R277 B.n623 B.n393 585
R278 B.n626 B.n625 585
R279 B.n627 B.n392 585
R280 B.n629 B.n628 585
R281 B.n631 B.n391 585
R282 B.n634 B.n633 585
R283 B.n635 B.n390 585
R284 B.n637 B.n636 585
R285 B.n639 B.n389 585
R286 B.n642 B.n641 585
R287 B.n643 B.n388 585
R288 B.n645 B.n644 585
R289 B.n647 B.n387 585
R290 B.n650 B.n649 585
R291 B.n651 B.n386 585
R292 B.n653 B.n652 585
R293 B.n655 B.n385 585
R294 B.n658 B.n657 585
R295 B.n659 B.n384 585
R296 B.n661 B.n660 585
R297 B.n663 B.n383 585
R298 B.n666 B.n665 585
R299 B.n667 B.n382 585
R300 B.n669 B.n668 585
R301 B.n671 B.n381 585
R302 B.n674 B.n673 585
R303 B.n675 B.n380 585
R304 B.n677 B.n676 585
R305 B.n679 B.n379 585
R306 B.n682 B.n681 585
R307 B.n683 B.n378 585
R308 B.n685 B.n684 585
R309 B.n687 B.n377 585
R310 B.n690 B.n689 585
R311 B.n691 B.n376 585
R312 B.n693 B.n692 585
R313 B.n695 B.n375 585
R314 B.n698 B.n697 585
R315 B.n699 B.n374 585
R316 B.n704 B.n703 585
R317 B.n703 B.n702 585
R318 B.n705 B.n370 585
R319 B.n370 B.n369 585
R320 B.n707 B.n706 585
R321 B.n708 B.n707 585
R322 B.n364 B.n363 585
R323 B.n365 B.n364 585
R324 B.n716 B.n715 585
R325 B.n715 B.n714 585
R326 B.n717 B.n362 585
R327 B.n362 B.n361 585
R328 B.n719 B.n718 585
R329 B.n720 B.n719 585
R330 B.n356 B.n355 585
R331 B.n357 B.n356 585
R332 B.n730 B.n729 585
R333 B.n729 B.n728 585
R334 B.n731 B.n354 585
R335 B.n727 B.n354 585
R336 B.n733 B.n732 585
R337 B.n734 B.n733 585
R338 B.n3 B.n0 585
R339 B.n4 B.n3 585
R340 B.n781 B.n1 585
R341 B.n782 B.n781 585
R342 B.n780 B.n779 585
R343 B.n780 B.n8 585
R344 B.n778 B.n9 585
R345 B.n12 B.n9 585
R346 B.n777 B.n776 585
R347 B.n776 B.n775 585
R348 B.n11 B.n10 585
R349 B.n774 B.n11 585
R350 B.n772 B.n771 585
R351 B.n773 B.n772 585
R352 B.n770 B.n17 585
R353 B.n17 B.n16 585
R354 B.n769 B.n768 585
R355 B.n768 B.n767 585
R356 B.n19 B.n18 585
R357 B.n766 B.n19 585
R358 B.n764 B.n763 585
R359 B.n765 B.n764 585
R360 B.n762 B.n24 585
R361 B.n24 B.n23 585
R362 B.n761 B.n760 585
R363 B.n760 B.n759 585
R364 B.n785 B.n784 585
R365 B.n783 B.n2 585
R366 B.n760 B.n26 511.721
R367 B.n757 B.n27 511.721
R368 B.n701 B.n374 511.721
R369 B.n703 B.n372 511.721
R370 B.n93 B.t14 402.353
R371 B.n405 B.t12 402.353
R372 B.n95 B.t8 402.353
R373 B.n411 B.t5 402.353
R374 B.n94 B.t15 387.613
R375 B.n406 B.t11 387.613
R376 B.n96 B.t9 387.613
R377 B.n412 B.t4 387.613
R378 B.n758 B.n91 256.663
R379 B.n758 B.n90 256.663
R380 B.n758 B.n89 256.663
R381 B.n758 B.n88 256.663
R382 B.n758 B.n87 256.663
R383 B.n758 B.n86 256.663
R384 B.n758 B.n85 256.663
R385 B.n758 B.n84 256.663
R386 B.n758 B.n83 256.663
R387 B.n758 B.n82 256.663
R388 B.n758 B.n81 256.663
R389 B.n758 B.n80 256.663
R390 B.n758 B.n79 256.663
R391 B.n758 B.n78 256.663
R392 B.n758 B.n77 256.663
R393 B.n758 B.n76 256.663
R394 B.n758 B.n75 256.663
R395 B.n758 B.n74 256.663
R396 B.n758 B.n73 256.663
R397 B.n758 B.n72 256.663
R398 B.n758 B.n71 256.663
R399 B.n758 B.n70 256.663
R400 B.n758 B.n69 256.663
R401 B.n758 B.n68 256.663
R402 B.n758 B.n67 256.663
R403 B.n758 B.n66 256.663
R404 B.n758 B.n65 256.663
R405 B.n758 B.n64 256.663
R406 B.n758 B.n63 256.663
R407 B.n758 B.n62 256.663
R408 B.n758 B.n61 256.663
R409 B.n758 B.n60 256.663
R410 B.n758 B.n59 256.663
R411 B.n758 B.n58 256.663
R412 B.n758 B.n57 256.663
R413 B.n758 B.n56 256.663
R414 B.n758 B.n55 256.663
R415 B.n758 B.n54 256.663
R416 B.n758 B.n53 256.663
R417 B.n758 B.n52 256.663
R418 B.n758 B.n51 256.663
R419 B.n758 B.n50 256.663
R420 B.n758 B.n49 256.663
R421 B.n758 B.n48 256.663
R422 B.n758 B.n47 256.663
R423 B.n758 B.n46 256.663
R424 B.n758 B.n45 256.663
R425 B.n758 B.n44 256.663
R426 B.n758 B.n43 256.663
R427 B.n758 B.n42 256.663
R428 B.n758 B.n41 256.663
R429 B.n758 B.n40 256.663
R430 B.n758 B.n39 256.663
R431 B.n758 B.n38 256.663
R432 B.n758 B.n37 256.663
R433 B.n758 B.n36 256.663
R434 B.n758 B.n35 256.663
R435 B.n758 B.n34 256.663
R436 B.n758 B.n33 256.663
R437 B.n758 B.n32 256.663
R438 B.n758 B.n31 256.663
R439 B.n758 B.n30 256.663
R440 B.n758 B.n29 256.663
R441 B.n758 B.n28 256.663
R442 B.n443 B.n373 256.663
R443 B.n446 B.n373 256.663
R444 B.n452 B.n373 256.663
R445 B.n454 B.n373 256.663
R446 B.n460 B.n373 256.663
R447 B.n462 B.n373 256.663
R448 B.n468 B.n373 256.663
R449 B.n470 B.n373 256.663
R450 B.n476 B.n373 256.663
R451 B.n478 B.n373 256.663
R452 B.n484 B.n373 256.663
R453 B.n486 B.n373 256.663
R454 B.n492 B.n373 256.663
R455 B.n494 B.n373 256.663
R456 B.n500 B.n373 256.663
R457 B.n502 B.n373 256.663
R458 B.n508 B.n373 256.663
R459 B.n510 B.n373 256.663
R460 B.n516 B.n373 256.663
R461 B.n518 B.n373 256.663
R462 B.n524 B.n373 256.663
R463 B.n526 B.n373 256.663
R464 B.n532 B.n373 256.663
R465 B.n534 B.n373 256.663
R466 B.n540 B.n373 256.663
R467 B.n542 B.n373 256.663
R468 B.n548 B.n373 256.663
R469 B.n550 B.n373 256.663
R470 B.n556 B.n373 256.663
R471 B.n558 B.n373 256.663
R472 B.n565 B.n373 256.663
R473 B.n567 B.n373 256.663
R474 B.n573 B.n373 256.663
R475 B.n575 B.n373 256.663
R476 B.n582 B.n373 256.663
R477 B.n584 B.n373 256.663
R478 B.n590 B.n373 256.663
R479 B.n592 B.n373 256.663
R480 B.n598 B.n373 256.663
R481 B.n600 B.n373 256.663
R482 B.n606 B.n373 256.663
R483 B.n608 B.n373 256.663
R484 B.n614 B.n373 256.663
R485 B.n616 B.n373 256.663
R486 B.n622 B.n373 256.663
R487 B.n624 B.n373 256.663
R488 B.n630 B.n373 256.663
R489 B.n632 B.n373 256.663
R490 B.n638 B.n373 256.663
R491 B.n640 B.n373 256.663
R492 B.n646 B.n373 256.663
R493 B.n648 B.n373 256.663
R494 B.n654 B.n373 256.663
R495 B.n656 B.n373 256.663
R496 B.n662 B.n373 256.663
R497 B.n664 B.n373 256.663
R498 B.n670 B.n373 256.663
R499 B.n672 B.n373 256.663
R500 B.n678 B.n373 256.663
R501 B.n680 B.n373 256.663
R502 B.n686 B.n373 256.663
R503 B.n688 B.n373 256.663
R504 B.n694 B.n373 256.663
R505 B.n696 B.n373 256.663
R506 B.n787 B.n786 256.663
R507 B.n100 B.n99 163.367
R508 B.n104 B.n103 163.367
R509 B.n108 B.n107 163.367
R510 B.n112 B.n111 163.367
R511 B.n116 B.n115 163.367
R512 B.n120 B.n119 163.367
R513 B.n124 B.n123 163.367
R514 B.n128 B.n127 163.367
R515 B.n132 B.n131 163.367
R516 B.n136 B.n135 163.367
R517 B.n140 B.n139 163.367
R518 B.n144 B.n143 163.367
R519 B.n148 B.n147 163.367
R520 B.n152 B.n151 163.367
R521 B.n156 B.n155 163.367
R522 B.n160 B.n159 163.367
R523 B.n164 B.n163 163.367
R524 B.n168 B.n167 163.367
R525 B.n172 B.n171 163.367
R526 B.n176 B.n175 163.367
R527 B.n180 B.n179 163.367
R528 B.n184 B.n183 163.367
R529 B.n188 B.n187 163.367
R530 B.n192 B.n191 163.367
R531 B.n196 B.n195 163.367
R532 B.n200 B.n199 163.367
R533 B.n204 B.n203 163.367
R534 B.n208 B.n207 163.367
R535 B.n212 B.n211 163.367
R536 B.n216 B.n215 163.367
R537 B.n220 B.n219 163.367
R538 B.n224 B.n223 163.367
R539 B.n228 B.n227 163.367
R540 B.n232 B.n231 163.367
R541 B.n237 B.n236 163.367
R542 B.n241 B.n240 163.367
R543 B.n245 B.n244 163.367
R544 B.n249 B.n248 163.367
R545 B.n253 B.n252 163.367
R546 B.n257 B.n256 163.367
R547 B.n261 B.n260 163.367
R548 B.n265 B.n264 163.367
R549 B.n269 B.n268 163.367
R550 B.n273 B.n272 163.367
R551 B.n277 B.n276 163.367
R552 B.n281 B.n280 163.367
R553 B.n285 B.n284 163.367
R554 B.n289 B.n288 163.367
R555 B.n293 B.n292 163.367
R556 B.n297 B.n296 163.367
R557 B.n301 B.n300 163.367
R558 B.n305 B.n304 163.367
R559 B.n309 B.n308 163.367
R560 B.n313 B.n312 163.367
R561 B.n317 B.n316 163.367
R562 B.n321 B.n320 163.367
R563 B.n325 B.n324 163.367
R564 B.n329 B.n328 163.367
R565 B.n333 B.n332 163.367
R566 B.n337 B.n336 163.367
R567 B.n341 B.n340 163.367
R568 B.n345 B.n344 163.367
R569 B.n349 B.n348 163.367
R570 B.n757 B.n92 163.367
R571 B.n701 B.n368 163.367
R572 B.n709 B.n368 163.367
R573 B.n709 B.n366 163.367
R574 B.n713 B.n366 163.367
R575 B.n713 B.n360 163.367
R576 B.n721 B.n360 163.367
R577 B.n721 B.n358 163.367
R578 B.n726 B.n358 163.367
R579 B.n726 B.n353 163.367
R580 B.n735 B.n353 163.367
R581 B.n736 B.n735 163.367
R582 B.n736 B.n5 163.367
R583 B.n6 B.n5 163.367
R584 B.n7 B.n6 163.367
R585 B.n742 B.n7 163.367
R586 B.n743 B.n742 163.367
R587 B.n743 B.n13 163.367
R588 B.n14 B.n13 163.367
R589 B.n15 B.n14 163.367
R590 B.n748 B.n15 163.367
R591 B.n748 B.n20 163.367
R592 B.n21 B.n20 163.367
R593 B.n22 B.n21 163.367
R594 B.n753 B.n22 163.367
R595 B.n753 B.n27 163.367
R596 B.n445 B.n444 163.367
R597 B.n447 B.n445 163.367
R598 B.n451 B.n440 163.367
R599 B.n455 B.n453 163.367
R600 B.n459 B.n438 163.367
R601 B.n463 B.n461 163.367
R602 B.n467 B.n436 163.367
R603 B.n471 B.n469 163.367
R604 B.n475 B.n434 163.367
R605 B.n479 B.n477 163.367
R606 B.n483 B.n432 163.367
R607 B.n487 B.n485 163.367
R608 B.n491 B.n430 163.367
R609 B.n495 B.n493 163.367
R610 B.n499 B.n428 163.367
R611 B.n503 B.n501 163.367
R612 B.n507 B.n426 163.367
R613 B.n511 B.n509 163.367
R614 B.n515 B.n424 163.367
R615 B.n519 B.n517 163.367
R616 B.n523 B.n422 163.367
R617 B.n527 B.n525 163.367
R618 B.n531 B.n420 163.367
R619 B.n535 B.n533 163.367
R620 B.n539 B.n418 163.367
R621 B.n543 B.n541 163.367
R622 B.n547 B.n416 163.367
R623 B.n551 B.n549 163.367
R624 B.n555 B.n414 163.367
R625 B.n559 B.n557 163.367
R626 B.n564 B.n410 163.367
R627 B.n568 B.n566 163.367
R628 B.n572 B.n408 163.367
R629 B.n576 B.n574 163.367
R630 B.n581 B.n404 163.367
R631 B.n585 B.n583 163.367
R632 B.n589 B.n402 163.367
R633 B.n593 B.n591 163.367
R634 B.n597 B.n400 163.367
R635 B.n601 B.n599 163.367
R636 B.n605 B.n398 163.367
R637 B.n609 B.n607 163.367
R638 B.n613 B.n396 163.367
R639 B.n617 B.n615 163.367
R640 B.n621 B.n394 163.367
R641 B.n625 B.n623 163.367
R642 B.n629 B.n392 163.367
R643 B.n633 B.n631 163.367
R644 B.n637 B.n390 163.367
R645 B.n641 B.n639 163.367
R646 B.n645 B.n388 163.367
R647 B.n649 B.n647 163.367
R648 B.n653 B.n386 163.367
R649 B.n657 B.n655 163.367
R650 B.n661 B.n384 163.367
R651 B.n665 B.n663 163.367
R652 B.n669 B.n382 163.367
R653 B.n673 B.n671 163.367
R654 B.n677 B.n380 163.367
R655 B.n681 B.n679 163.367
R656 B.n685 B.n378 163.367
R657 B.n689 B.n687 163.367
R658 B.n693 B.n376 163.367
R659 B.n697 B.n695 163.367
R660 B.n703 B.n370 163.367
R661 B.n707 B.n370 163.367
R662 B.n707 B.n364 163.367
R663 B.n715 B.n364 163.367
R664 B.n715 B.n362 163.367
R665 B.n719 B.n362 163.367
R666 B.n719 B.n356 163.367
R667 B.n729 B.n356 163.367
R668 B.n729 B.n354 163.367
R669 B.n733 B.n354 163.367
R670 B.n733 B.n3 163.367
R671 B.n785 B.n3 163.367
R672 B.n781 B.n2 163.367
R673 B.n781 B.n780 163.367
R674 B.n780 B.n9 163.367
R675 B.n776 B.n9 163.367
R676 B.n776 B.n11 163.367
R677 B.n772 B.n11 163.367
R678 B.n772 B.n17 163.367
R679 B.n768 B.n17 163.367
R680 B.n768 B.n19 163.367
R681 B.n764 B.n19 163.367
R682 B.n764 B.n24 163.367
R683 B.n760 B.n24 163.367
R684 B.n28 B.n26 71.676
R685 B.n100 B.n29 71.676
R686 B.n104 B.n30 71.676
R687 B.n108 B.n31 71.676
R688 B.n112 B.n32 71.676
R689 B.n116 B.n33 71.676
R690 B.n120 B.n34 71.676
R691 B.n124 B.n35 71.676
R692 B.n128 B.n36 71.676
R693 B.n132 B.n37 71.676
R694 B.n136 B.n38 71.676
R695 B.n140 B.n39 71.676
R696 B.n144 B.n40 71.676
R697 B.n148 B.n41 71.676
R698 B.n152 B.n42 71.676
R699 B.n156 B.n43 71.676
R700 B.n160 B.n44 71.676
R701 B.n164 B.n45 71.676
R702 B.n168 B.n46 71.676
R703 B.n172 B.n47 71.676
R704 B.n176 B.n48 71.676
R705 B.n180 B.n49 71.676
R706 B.n184 B.n50 71.676
R707 B.n188 B.n51 71.676
R708 B.n192 B.n52 71.676
R709 B.n196 B.n53 71.676
R710 B.n200 B.n54 71.676
R711 B.n204 B.n55 71.676
R712 B.n208 B.n56 71.676
R713 B.n212 B.n57 71.676
R714 B.n216 B.n58 71.676
R715 B.n220 B.n59 71.676
R716 B.n224 B.n60 71.676
R717 B.n228 B.n61 71.676
R718 B.n232 B.n62 71.676
R719 B.n237 B.n63 71.676
R720 B.n241 B.n64 71.676
R721 B.n245 B.n65 71.676
R722 B.n249 B.n66 71.676
R723 B.n253 B.n67 71.676
R724 B.n257 B.n68 71.676
R725 B.n261 B.n69 71.676
R726 B.n265 B.n70 71.676
R727 B.n269 B.n71 71.676
R728 B.n273 B.n72 71.676
R729 B.n277 B.n73 71.676
R730 B.n281 B.n74 71.676
R731 B.n285 B.n75 71.676
R732 B.n289 B.n76 71.676
R733 B.n293 B.n77 71.676
R734 B.n297 B.n78 71.676
R735 B.n301 B.n79 71.676
R736 B.n305 B.n80 71.676
R737 B.n309 B.n81 71.676
R738 B.n313 B.n82 71.676
R739 B.n317 B.n83 71.676
R740 B.n321 B.n84 71.676
R741 B.n325 B.n85 71.676
R742 B.n329 B.n86 71.676
R743 B.n333 B.n87 71.676
R744 B.n337 B.n88 71.676
R745 B.n341 B.n89 71.676
R746 B.n345 B.n90 71.676
R747 B.n349 B.n91 71.676
R748 B.n92 B.n91 71.676
R749 B.n348 B.n90 71.676
R750 B.n344 B.n89 71.676
R751 B.n340 B.n88 71.676
R752 B.n336 B.n87 71.676
R753 B.n332 B.n86 71.676
R754 B.n328 B.n85 71.676
R755 B.n324 B.n84 71.676
R756 B.n320 B.n83 71.676
R757 B.n316 B.n82 71.676
R758 B.n312 B.n81 71.676
R759 B.n308 B.n80 71.676
R760 B.n304 B.n79 71.676
R761 B.n300 B.n78 71.676
R762 B.n296 B.n77 71.676
R763 B.n292 B.n76 71.676
R764 B.n288 B.n75 71.676
R765 B.n284 B.n74 71.676
R766 B.n280 B.n73 71.676
R767 B.n276 B.n72 71.676
R768 B.n272 B.n71 71.676
R769 B.n268 B.n70 71.676
R770 B.n264 B.n69 71.676
R771 B.n260 B.n68 71.676
R772 B.n256 B.n67 71.676
R773 B.n252 B.n66 71.676
R774 B.n248 B.n65 71.676
R775 B.n244 B.n64 71.676
R776 B.n240 B.n63 71.676
R777 B.n236 B.n62 71.676
R778 B.n231 B.n61 71.676
R779 B.n227 B.n60 71.676
R780 B.n223 B.n59 71.676
R781 B.n219 B.n58 71.676
R782 B.n215 B.n57 71.676
R783 B.n211 B.n56 71.676
R784 B.n207 B.n55 71.676
R785 B.n203 B.n54 71.676
R786 B.n199 B.n53 71.676
R787 B.n195 B.n52 71.676
R788 B.n191 B.n51 71.676
R789 B.n187 B.n50 71.676
R790 B.n183 B.n49 71.676
R791 B.n179 B.n48 71.676
R792 B.n175 B.n47 71.676
R793 B.n171 B.n46 71.676
R794 B.n167 B.n45 71.676
R795 B.n163 B.n44 71.676
R796 B.n159 B.n43 71.676
R797 B.n155 B.n42 71.676
R798 B.n151 B.n41 71.676
R799 B.n147 B.n40 71.676
R800 B.n143 B.n39 71.676
R801 B.n139 B.n38 71.676
R802 B.n135 B.n37 71.676
R803 B.n131 B.n36 71.676
R804 B.n127 B.n35 71.676
R805 B.n123 B.n34 71.676
R806 B.n119 B.n33 71.676
R807 B.n115 B.n32 71.676
R808 B.n111 B.n31 71.676
R809 B.n107 B.n30 71.676
R810 B.n103 B.n29 71.676
R811 B.n99 B.n28 71.676
R812 B.n443 B.n372 71.676
R813 B.n447 B.n446 71.676
R814 B.n452 B.n451 71.676
R815 B.n455 B.n454 71.676
R816 B.n460 B.n459 71.676
R817 B.n463 B.n462 71.676
R818 B.n468 B.n467 71.676
R819 B.n471 B.n470 71.676
R820 B.n476 B.n475 71.676
R821 B.n479 B.n478 71.676
R822 B.n484 B.n483 71.676
R823 B.n487 B.n486 71.676
R824 B.n492 B.n491 71.676
R825 B.n495 B.n494 71.676
R826 B.n500 B.n499 71.676
R827 B.n503 B.n502 71.676
R828 B.n508 B.n507 71.676
R829 B.n511 B.n510 71.676
R830 B.n516 B.n515 71.676
R831 B.n519 B.n518 71.676
R832 B.n524 B.n523 71.676
R833 B.n527 B.n526 71.676
R834 B.n532 B.n531 71.676
R835 B.n535 B.n534 71.676
R836 B.n540 B.n539 71.676
R837 B.n543 B.n542 71.676
R838 B.n548 B.n547 71.676
R839 B.n551 B.n550 71.676
R840 B.n556 B.n555 71.676
R841 B.n559 B.n558 71.676
R842 B.n565 B.n564 71.676
R843 B.n568 B.n567 71.676
R844 B.n573 B.n572 71.676
R845 B.n576 B.n575 71.676
R846 B.n582 B.n581 71.676
R847 B.n585 B.n584 71.676
R848 B.n590 B.n589 71.676
R849 B.n593 B.n592 71.676
R850 B.n598 B.n597 71.676
R851 B.n601 B.n600 71.676
R852 B.n606 B.n605 71.676
R853 B.n609 B.n608 71.676
R854 B.n614 B.n613 71.676
R855 B.n617 B.n616 71.676
R856 B.n622 B.n621 71.676
R857 B.n625 B.n624 71.676
R858 B.n630 B.n629 71.676
R859 B.n633 B.n632 71.676
R860 B.n638 B.n637 71.676
R861 B.n641 B.n640 71.676
R862 B.n646 B.n645 71.676
R863 B.n649 B.n648 71.676
R864 B.n654 B.n653 71.676
R865 B.n657 B.n656 71.676
R866 B.n662 B.n661 71.676
R867 B.n665 B.n664 71.676
R868 B.n670 B.n669 71.676
R869 B.n673 B.n672 71.676
R870 B.n678 B.n677 71.676
R871 B.n681 B.n680 71.676
R872 B.n686 B.n685 71.676
R873 B.n689 B.n688 71.676
R874 B.n694 B.n693 71.676
R875 B.n697 B.n696 71.676
R876 B.n444 B.n443 71.676
R877 B.n446 B.n440 71.676
R878 B.n453 B.n452 71.676
R879 B.n454 B.n438 71.676
R880 B.n461 B.n460 71.676
R881 B.n462 B.n436 71.676
R882 B.n469 B.n468 71.676
R883 B.n470 B.n434 71.676
R884 B.n477 B.n476 71.676
R885 B.n478 B.n432 71.676
R886 B.n485 B.n484 71.676
R887 B.n486 B.n430 71.676
R888 B.n493 B.n492 71.676
R889 B.n494 B.n428 71.676
R890 B.n501 B.n500 71.676
R891 B.n502 B.n426 71.676
R892 B.n509 B.n508 71.676
R893 B.n510 B.n424 71.676
R894 B.n517 B.n516 71.676
R895 B.n518 B.n422 71.676
R896 B.n525 B.n524 71.676
R897 B.n526 B.n420 71.676
R898 B.n533 B.n532 71.676
R899 B.n534 B.n418 71.676
R900 B.n541 B.n540 71.676
R901 B.n542 B.n416 71.676
R902 B.n549 B.n548 71.676
R903 B.n550 B.n414 71.676
R904 B.n557 B.n556 71.676
R905 B.n558 B.n410 71.676
R906 B.n566 B.n565 71.676
R907 B.n567 B.n408 71.676
R908 B.n574 B.n573 71.676
R909 B.n575 B.n404 71.676
R910 B.n583 B.n582 71.676
R911 B.n584 B.n402 71.676
R912 B.n591 B.n590 71.676
R913 B.n592 B.n400 71.676
R914 B.n599 B.n598 71.676
R915 B.n600 B.n398 71.676
R916 B.n607 B.n606 71.676
R917 B.n608 B.n396 71.676
R918 B.n615 B.n614 71.676
R919 B.n616 B.n394 71.676
R920 B.n623 B.n622 71.676
R921 B.n624 B.n392 71.676
R922 B.n631 B.n630 71.676
R923 B.n632 B.n390 71.676
R924 B.n639 B.n638 71.676
R925 B.n640 B.n388 71.676
R926 B.n647 B.n646 71.676
R927 B.n648 B.n386 71.676
R928 B.n655 B.n654 71.676
R929 B.n656 B.n384 71.676
R930 B.n663 B.n662 71.676
R931 B.n664 B.n382 71.676
R932 B.n671 B.n670 71.676
R933 B.n672 B.n380 71.676
R934 B.n679 B.n678 71.676
R935 B.n680 B.n378 71.676
R936 B.n687 B.n686 71.676
R937 B.n688 B.n376 71.676
R938 B.n695 B.n694 71.676
R939 B.n696 B.n374 71.676
R940 B.n786 B.n785 71.676
R941 B.n786 B.n2 71.676
R942 B.n702 B.n373 60.5768
R943 B.n759 B.n758 60.5768
R944 B.n97 B.n96 59.5399
R945 B.n234 B.n94 59.5399
R946 B.n579 B.n406 59.5399
R947 B.n561 B.n412 59.5399
R948 B.n704 B.n371 33.2493
R949 B.n700 B.n699 33.2493
R950 B.n756 B.n755 33.2493
R951 B.n761 B.n25 33.2493
R952 B.n702 B.n369 31.9322
R953 B.n708 B.n369 31.9322
R954 B.n708 B.n365 31.9322
R955 B.n714 B.n365 31.9322
R956 B.n720 B.n361 31.9322
R957 B.n720 B.n357 31.9322
R958 B.n728 B.n357 31.9322
R959 B.n728 B.n727 31.9322
R960 B.n734 B.n4 31.9322
R961 B.n784 B.n4 31.9322
R962 B.n784 B.n783 31.9322
R963 B.n783 B.n782 31.9322
R964 B.n782 B.n8 31.9322
R965 B.n775 B.n12 31.9322
R966 B.n775 B.n774 31.9322
R967 B.n774 B.n773 31.9322
R968 B.n773 B.n16 31.9322
R969 B.n767 B.n766 31.9322
R970 B.n766 B.n765 31.9322
R971 B.n765 B.n23 31.9322
R972 B.n759 B.n23 31.9322
R973 B.n727 B.t1 24.8884
R974 B.n12 B.t0 24.8884
R975 B.t3 B.n361 21.1318
R976 B.t7 B.n16 21.1318
R977 B B.n787 18.0485
R978 B.n96 B.n95 14.7399
R979 B.n94 B.n93 14.7399
R980 B.n406 B.n405 14.7399
R981 B.n412 B.n411 14.7399
R982 B.n714 B.t3 10.8009
R983 B.n767 B.t7 10.8009
R984 B.n705 B.n704 10.6151
R985 B.n706 B.n705 10.6151
R986 B.n706 B.n363 10.6151
R987 B.n716 B.n363 10.6151
R988 B.n717 B.n716 10.6151
R989 B.n718 B.n717 10.6151
R990 B.n718 B.n355 10.6151
R991 B.n730 B.n355 10.6151
R992 B.n731 B.n730 10.6151
R993 B.n732 B.n731 10.6151
R994 B.n732 B.n0 10.6151
R995 B.n442 B.n371 10.6151
R996 B.n442 B.n441 10.6151
R997 B.n448 B.n441 10.6151
R998 B.n449 B.n448 10.6151
R999 B.n450 B.n449 10.6151
R1000 B.n450 B.n439 10.6151
R1001 B.n456 B.n439 10.6151
R1002 B.n457 B.n456 10.6151
R1003 B.n458 B.n457 10.6151
R1004 B.n458 B.n437 10.6151
R1005 B.n464 B.n437 10.6151
R1006 B.n465 B.n464 10.6151
R1007 B.n466 B.n465 10.6151
R1008 B.n466 B.n435 10.6151
R1009 B.n472 B.n435 10.6151
R1010 B.n473 B.n472 10.6151
R1011 B.n474 B.n473 10.6151
R1012 B.n474 B.n433 10.6151
R1013 B.n480 B.n433 10.6151
R1014 B.n481 B.n480 10.6151
R1015 B.n482 B.n481 10.6151
R1016 B.n482 B.n431 10.6151
R1017 B.n488 B.n431 10.6151
R1018 B.n489 B.n488 10.6151
R1019 B.n490 B.n489 10.6151
R1020 B.n490 B.n429 10.6151
R1021 B.n496 B.n429 10.6151
R1022 B.n497 B.n496 10.6151
R1023 B.n498 B.n497 10.6151
R1024 B.n498 B.n427 10.6151
R1025 B.n504 B.n427 10.6151
R1026 B.n505 B.n504 10.6151
R1027 B.n506 B.n505 10.6151
R1028 B.n506 B.n425 10.6151
R1029 B.n512 B.n425 10.6151
R1030 B.n513 B.n512 10.6151
R1031 B.n514 B.n513 10.6151
R1032 B.n514 B.n423 10.6151
R1033 B.n520 B.n423 10.6151
R1034 B.n521 B.n520 10.6151
R1035 B.n522 B.n521 10.6151
R1036 B.n522 B.n421 10.6151
R1037 B.n528 B.n421 10.6151
R1038 B.n529 B.n528 10.6151
R1039 B.n530 B.n529 10.6151
R1040 B.n530 B.n419 10.6151
R1041 B.n536 B.n419 10.6151
R1042 B.n537 B.n536 10.6151
R1043 B.n538 B.n537 10.6151
R1044 B.n538 B.n417 10.6151
R1045 B.n544 B.n417 10.6151
R1046 B.n545 B.n544 10.6151
R1047 B.n546 B.n545 10.6151
R1048 B.n546 B.n415 10.6151
R1049 B.n552 B.n415 10.6151
R1050 B.n553 B.n552 10.6151
R1051 B.n554 B.n553 10.6151
R1052 B.n554 B.n413 10.6151
R1053 B.n560 B.n413 10.6151
R1054 B.n563 B.n562 10.6151
R1055 B.n563 B.n409 10.6151
R1056 B.n569 B.n409 10.6151
R1057 B.n570 B.n569 10.6151
R1058 B.n571 B.n570 10.6151
R1059 B.n571 B.n407 10.6151
R1060 B.n577 B.n407 10.6151
R1061 B.n578 B.n577 10.6151
R1062 B.n580 B.n403 10.6151
R1063 B.n586 B.n403 10.6151
R1064 B.n587 B.n586 10.6151
R1065 B.n588 B.n587 10.6151
R1066 B.n588 B.n401 10.6151
R1067 B.n594 B.n401 10.6151
R1068 B.n595 B.n594 10.6151
R1069 B.n596 B.n595 10.6151
R1070 B.n596 B.n399 10.6151
R1071 B.n602 B.n399 10.6151
R1072 B.n603 B.n602 10.6151
R1073 B.n604 B.n603 10.6151
R1074 B.n604 B.n397 10.6151
R1075 B.n610 B.n397 10.6151
R1076 B.n611 B.n610 10.6151
R1077 B.n612 B.n611 10.6151
R1078 B.n612 B.n395 10.6151
R1079 B.n618 B.n395 10.6151
R1080 B.n619 B.n618 10.6151
R1081 B.n620 B.n619 10.6151
R1082 B.n620 B.n393 10.6151
R1083 B.n626 B.n393 10.6151
R1084 B.n627 B.n626 10.6151
R1085 B.n628 B.n627 10.6151
R1086 B.n628 B.n391 10.6151
R1087 B.n634 B.n391 10.6151
R1088 B.n635 B.n634 10.6151
R1089 B.n636 B.n635 10.6151
R1090 B.n636 B.n389 10.6151
R1091 B.n642 B.n389 10.6151
R1092 B.n643 B.n642 10.6151
R1093 B.n644 B.n643 10.6151
R1094 B.n644 B.n387 10.6151
R1095 B.n650 B.n387 10.6151
R1096 B.n651 B.n650 10.6151
R1097 B.n652 B.n651 10.6151
R1098 B.n652 B.n385 10.6151
R1099 B.n658 B.n385 10.6151
R1100 B.n659 B.n658 10.6151
R1101 B.n660 B.n659 10.6151
R1102 B.n660 B.n383 10.6151
R1103 B.n666 B.n383 10.6151
R1104 B.n667 B.n666 10.6151
R1105 B.n668 B.n667 10.6151
R1106 B.n668 B.n381 10.6151
R1107 B.n674 B.n381 10.6151
R1108 B.n675 B.n674 10.6151
R1109 B.n676 B.n675 10.6151
R1110 B.n676 B.n379 10.6151
R1111 B.n682 B.n379 10.6151
R1112 B.n683 B.n682 10.6151
R1113 B.n684 B.n683 10.6151
R1114 B.n684 B.n377 10.6151
R1115 B.n690 B.n377 10.6151
R1116 B.n691 B.n690 10.6151
R1117 B.n692 B.n691 10.6151
R1118 B.n692 B.n375 10.6151
R1119 B.n698 B.n375 10.6151
R1120 B.n699 B.n698 10.6151
R1121 B.n700 B.n367 10.6151
R1122 B.n710 B.n367 10.6151
R1123 B.n711 B.n710 10.6151
R1124 B.n712 B.n711 10.6151
R1125 B.n712 B.n359 10.6151
R1126 B.n722 B.n359 10.6151
R1127 B.n723 B.n722 10.6151
R1128 B.n725 B.n723 10.6151
R1129 B.n725 B.n724 10.6151
R1130 B.n724 B.n352 10.6151
R1131 B.n737 B.n352 10.6151
R1132 B.n738 B.n737 10.6151
R1133 B.n739 B.n738 10.6151
R1134 B.n740 B.n739 10.6151
R1135 B.n741 B.n740 10.6151
R1136 B.n744 B.n741 10.6151
R1137 B.n745 B.n744 10.6151
R1138 B.n746 B.n745 10.6151
R1139 B.n747 B.n746 10.6151
R1140 B.n749 B.n747 10.6151
R1141 B.n750 B.n749 10.6151
R1142 B.n751 B.n750 10.6151
R1143 B.n752 B.n751 10.6151
R1144 B.n754 B.n752 10.6151
R1145 B.n755 B.n754 10.6151
R1146 B.n779 B.n1 10.6151
R1147 B.n779 B.n778 10.6151
R1148 B.n778 B.n777 10.6151
R1149 B.n777 B.n10 10.6151
R1150 B.n771 B.n10 10.6151
R1151 B.n771 B.n770 10.6151
R1152 B.n770 B.n769 10.6151
R1153 B.n769 B.n18 10.6151
R1154 B.n763 B.n18 10.6151
R1155 B.n763 B.n762 10.6151
R1156 B.n762 B.n761 10.6151
R1157 B.n98 B.n25 10.6151
R1158 B.n101 B.n98 10.6151
R1159 B.n102 B.n101 10.6151
R1160 B.n105 B.n102 10.6151
R1161 B.n106 B.n105 10.6151
R1162 B.n109 B.n106 10.6151
R1163 B.n110 B.n109 10.6151
R1164 B.n113 B.n110 10.6151
R1165 B.n114 B.n113 10.6151
R1166 B.n117 B.n114 10.6151
R1167 B.n118 B.n117 10.6151
R1168 B.n121 B.n118 10.6151
R1169 B.n122 B.n121 10.6151
R1170 B.n125 B.n122 10.6151
R1171 B.n126 B.n125 10.6151
R1172 B.n129 B.n126 10.6151
R1173 B.n130 B.n129 10.6151
R1174 B.n133 B.n130 10.6151
R1175 B.n134 B.n133 10.6151
R1176 B.n137 B.n134 10.6151
R1177 B.n138 B.n137 10.6151
R1178 B.n141 B.n138 10.6151
R1179 B.n142 B.n141 10.6151
R1180 B.n145 B.n142 10.6151
R1181 B.n146 B.n145 10.6151
R1182 B.n149 B.n146 10.6151
R1183 B.n150 B.n149 10.6151
R1184 B.n153 B.n150 10.6151
R1185 B.n154 B.n153 10.6151
R1186 B.n157 B.n154 10.6151
R1187 B.n158 B.n157 10.6151
R1188 B.n161 B.n158 10.6151
R1189 B.n162 B.n161 10.6151
R1190 B.n165 B.n162 10.6151
R1191 B.n166 B.n165 10.6151
R1192 B.n169 B.n166 10.6151
R1193 B.n170 B.n169 10.6151
R1194 B.n173 B.n170 10.6151
R1195 B.n174 B.n173 10.6151
R1196 B.n177 B.n174 10.6151
R1197 B.n178 B.n177 10.6151
R1198 B.n181 B.n178 10.6151
R1199 B.n182 B.n181 10.6151
R1200 B.n185 B.n182 10.6151
R1201 B.n186 B.n185 10.6151
R1202 B.n189 B.n186 10.6151
R1203 B.n190 B.n189 10.6151
R1204 B.n193 B.n190 10.6151
R1205 B.n194 B.n193 10.6151
R1206 B.n197 B.n194 10.6151
R1207 B.n198 B.n197 10.6151
R1208 B.n201 B.n198 10.6151
R1209 B.n202 B.n201 10.6151
R1210 B.n205 B.n202 10.6151
R1211 B.n206 B.n205 10.6151
R1212 B.n209 B.n206 10.6151
R1213 B.n210 B.n209 10.6151
R1214 B.n213 B.n210 10.6151
R1215 B.n214 B.n213 10.6151
R1216 B.n218 B.n217 10.6151
R1217 B.n221 B.n218 10.6151
R1218 B.n222 B.n221 10.6151
R1219 B.n225 B.n222 10.6151
R1220 B.n226 B.n225 10.6151
R1221 B.n229 B.n226 10.6151
R1222 B.n230 B.n229 10.6151
R1223 B.n233 B.n230 10.6151
R1224 B.n238 B.n235 10.6151
R1225 B.n239 B.n238 10.6151
R1226 B.n242 B.n239 10.6151
R1227 B.n243 B.n242 10.6151
R1228 B.n246 B.n243 10.6151
R1229 B.n247 B.n246 10.6151
R1230 B.n250 B.n247 10.6151
R1231 B.n251 B.n250 10.6151
R1232 B.n254 B.n251 10.6151
R1233 B.n255 B.n254 10.6151
R1234 B.n258 B.n255 10.6151
R1235 B.n259 B.n258 10.6151
R1236 B.n262 B.n259 10.6151
R1237 B.n263 B.n262 10.6151
R1238 B.n266 B.n263 10.6151
R1239 B.n267 B.n266 10.6151
R1240 B.n270 B.n267 10.6151
R1241 B.n271 B.n270 10.6151
R1242 B.n274 B.n271 10.6151
R1243 B.n275 B.n274 10.6151
R1244 B.n278 B.n275 10.6151
R1245 B.n279 B.n278 10.6151
R1246 B.n282 B.n279 10.6151
R1247 B.n283 B.n282 10.6151
R1248 B.n286 B.n283 10.6151
R1249 B.n287 B.n286 10.6151
R1250 B.n290 B.n287 10.6151
R1251 B.n291 B.n290 10.6151
R1252 B.n294 B.n291 10.6151
R1253 B.n295 B.n294 10.6151
R1254 B.n298 B.n295 10.6151
R1255 B.n299 B.n298 10.6151
R1256 B.n302 B.n299 10.6151
R1257 B.n303 B.n302 10.6151
R1258 B.n306 B.n303 10.6151
R1259 B.n307 B.n306 10.6151
R1260 B.n310 B.n307 10.6151
R1261 B.n311 B.n310 10.6151
R1262 B.n314 B.n311 10.6151
R1263 B.n315 B.n314 10.6151
R1264 B.n318 B.n315 10.6151
R1265 B.n319 B.n318 10.6151
R1266 B.n322 B.n319 10.6151
R1267 B.n323 B.n322 10.6151
R1268 B.n326 B.n323 10.6151
R1269 B.n327 B.n326 10.6151
R1270 B.n330 B.n327 10.6151
R1271 B.n331 B.n330 10.6151
R1272 B.n334 B.n331 10.6151
R1273 B.n335 B.n334 10.6151
R1274 B.n338 B.n335 10.6151
R1275 B.n339 B.n338 10.6151
R1276 B.n342 B.n339 10.6151
R1277 B.n343 B.n342 10.6151
R1278 B.n346 B.n343 10.6151
R1279 B.n347 B.n346 10.6151
R1280 B.n350 B.n347 10.6151
R1281 B.n351 B.n350 10.6151
R1282 B.n756 B.n351 10.6151
R1283 B.n787 B.n0 8.11757
R1284 B.n787 B.n1 8.11757
R1285 B.n562 B.n561 7.18099
R1286 B.n579 B.n578 7.18099
R1287 B.n217 B.n97 7.18099
R1288 B.n234 B.n233 7.18099
R1289 B.n734 B.t1 7.04426
R1290 B.t0 B.n8 7.04426
R1291 B.n561 B.n560 3.43465
R1292 B.n580 B.n579 3.43465
R1293 B.n214 B.n97 3.43465
R1294 B.n235 B.n234 3.43465
R1295 VN VN.t0 1313.28
R1296 VN VN.t1 1269.39
R1297 VTAIL.n402 VTAIL.n306 289.615
R1298 VTAIL.n96 VTAIL.n0 289.615
R1299 VTAIL.n300 VTAIL.n204 289.615
R1300 VTAIL.n198 VTAIL.n102 289.615
R1301 VTAIL.n338 VTAIL.n337 185
R1302 VTAIL.n343 VTAIL.n342 185
R1303 VTAIL.n345 VTAIL.n344 185
R1304 VTAIL.n334 VTAIL.n333 185
R1305 VTAIL.n351 VTAIL.n350 185
R1306 VTAIL.n353 VTAIL.n352 185
R1307 VTAIL.n330 VTAIL.n329 185
R1308 VTAIL.n359 VTAIL.n358 185
R1309 VTAIL.n361 VTAIL.n360 185
R1310 VTAIL.n326 VTAIL.n325 185
R1311 VTAIL.n367 VTAIL.n366 185
R1312 VTAIL.n369 VTAIL.n368 185
R1313 VTAIL.n322 VTAIL.n321 185
R1314 VTAIL.n375 VTAIL.n374 185
R1315 VTAIL.n377 VTAIL.n376 185
R1316 VTAIL.n318 VTAIL.n317 185
R1317 VTAIL.n384 VTAIL.n383 185
R1318 VTAIL.n385 VTAIL.n316 185
R1319 VTAIL.n387 VTAIL.n386 185
R1320 VTAIL.n314 VTAIL.n313 185
R1321 VTAIL.n393 VTAIL.n392 185
R1322 VTAIL.n395 VTAIL.n394 185
R1323 VTAIL.n310 VTAIL.n309 185
R1324 VTAIL.n401 VTAIL.n400 185
R1325 VTAIL.n403 VTAIL.n402 185
R1326 VTAIL.n32 VTAIL.n31 185
R1327 VTAIL.n37 VTAIL.n36 185
R1328 VTAIL.n39 VTAIL.n38 185
R1329 VTAIL.n28 VTAIL.n27 185
R1330 VTAIL.n45 VTAIL.n44 185
R1331 VTAIL.n47 VTAIL.n46 185
R1332 VTAIL.n24 VTAIL.n23 185
R1333 VTAIL.n53 VTAIL.n52 185
R1334 VTAIL.n55 VTAIL.n54 185
R1335 VTAIL.n20 VTAIL.n19 185
R1336 VTAIL.n61 VTAIL.n60 185
R1337 VTAIL.n63 VTAIL.n62 185
R1338 VTAIL.n16 VTAIL.n15 185
R1339 VTAIL.n69 VTAIL.n68 185
R1340 VTAIL.n71 VTAIL.n70 185
R1341 VTAIL.n12 VTAIL.n11 185
R1342 VTAIL.n78 VTAIL.n77 185
R1343 VTAIL.n79 VTAIL.n10 185
R1344 VTAIL.n81 VTAIL.n80 185
R1345 VTAIL.n8 VTAIL.n7 185
R1346 VTAIL.n87 VTAIL.n86 185
R1347 VTAIL.n89 VTAIL.n88 185
R1348 VTAIL.n4 VTAIL.n3 185
R1349 VTAIL.n95 VTAIL.n94 185
R1350 VTAIL.n97 VTAIL.n96 185
R1351 VTAIL.n301 VTAIL.n300 185
R1352 VTAIL.n299 VTAIL.n298 185
R1353 VTAIL.n208 VTAIL.n207 185
R1354 VTAIL.n293 VTAIL.n292 185
R1355 VTAIL.n291 VTAIL.n290 185
R1356 VTAIL.n212 VTAIL.n211 185
R1357 VTAIL.n285 VTAIL.n284 185
R1358 VTAIL.n283 VTAIL.n214 185
R1359 VTAIL.n282 VTAIL.n281 185
R1360 VTAIL.n217 VTAIL.n215 185
R1361 VTAIL.n276 VTAIL.n275 185
R1362 VTAIL.n274 VTAIL.n273 185
R1363 VTAIL.n221 VTAIL.n220 185
R1364 VTAIL.n268 VTAIL.n267 185
R1365 VTAIL.n266 VTAIL.n265 185
R1366 VTAIL.n225 VTAIL.n224 185
R1367 VTAIL.n260 VTAIL.n259 185
R1368 VTAIL.n258 VTAIL.n257 185
R1369 VTAIL.n229 VTAIL.n228 185
R1370 VTAIL.n252 VTAIL.n251 185
R1371 VTAIL.n250 VTAIL.n249 185
R1372 VTAIL.n233 VTAIL.n232 185
R1373 VTAIL.n244 VTAIL.n243 185
R1374 VTAIL.n242 VTAIL.n241 185
R1375 VTAIL.n237 VTAIL.n236 185
R1376 VTAIL.n199 VTAIL.n198 185
R1377 VTAIL.n197 VTAIL.n196 185
R1378 VTAIL.n106 VTAIL.n105 185
R1379 VTAIL.n191 VTAIL.n190 185
R1380 VTAIL.n189 VTAIL.n188 185
R1381 VTAIL.n110 VTAIL.n109 185
R1382 VTAIL.n183 VTAIL.n182 185
R1383 VTAIL.n181 VTAIL.n112 185
R1384 VTAIL.n180 VTAIL.n179 185
R1385 VTAIL.n115 VTAIL.n113 185
R1386 VTAIL.n174 VTAIL.n173 185
R1387 VTAIL.n172 VTAIL.n171 185
R1388 VTAIL.n119 VTAIL.n118 185
R1389 VTAIL.n166 VTAIL.n165 185
R1390 VTAIL.n164 VTAIL.n163 185
R1391 VTAIL.n123 VTAIL.n122 185
R1392 VTAIL.n158 VTAIL.n157 185
R1393 VTAIL.n156 VTAIL.n155 185
R1394 VTAIL.n127 VTAIL.n126 185
R1395 VTAIL.n150 VTAIL.n149 185
R1396 VTAIL.n148 VTAIL.n147 185
R1397 VTAIL.n131 VTAIL.n130 185
R1398 VTAIL.n142 VTAIL.n141 185
R1399 VTAIL.n140 VTAIL.n139 185
R1400 VTAIL.n135 VTAIL.n134 185
R1401 VTAIL.n339 VTAIL.t3 147.659
R1402 VTAIL.n33 VTAIL.t1 147.659
R1403 VTAIL.n238 VTAIL.t0 147.659
R1404 VTAIL.n136 VTAIL.t2 147.659
R1405 VTAIL.n343 VTAIL.n337 104.615
R1406 VTAIL.n344 VTAIL.n343 104.615
R1407 VTAIL.n344 VTAIL.n333 104.615
R1408 VTAIL.n351 VTAIL.n333 104.615
R1409 VTAIL.n352 VTAIL.n351 104.615
R1410 VTAIL.n352 VTAIL.n329 104.615
R1411 VTAIL.n359 VTAIL.n329 104.615
R1412 VTAIL.n360 VTAIL.n359 104.615
R1413 VTAIL.n360 VTAIL.n325 104.615
R1414 VTAIL.n367 VTAIL.n325 104.615
R1415 VTAIL.n368 VTAIL.n367 104.615
R1416 VTAIL.n368 VTAIL.n321 104.615
R1417 VTAIL.n375 VTAIL.n321 104.615
R1418 VTAIL.n376 VTAIL.n375 104.615
R1419 VTAIL.n376 VTAIL.n317 104.615
R1420 VTAIL.n384 VTAIL.n317 104.615
R1421 VTAIL.n385 VTAIL.n384 104.615
R1422 VTAIL.n386 VTAIL.n385 104.615
R1423 VTAIL.n386 VTAIL.n313 104.615
R1424 VTAIL.n393 VTAIL.n313 104.615
R1425 VTAIL.n394 VTAIL.n393 104.615
R1426 VTAIL.n394 VTAIL.n309 104.615
R1427 VTAIL.n401 VTAIL.n309 104.615
R1428 VTAIL.n402 VTAIL.n401 104.615
R1429 VTAIL.n37 VTAIL.n31 104.615
R1430 VTAIL.n38 VTAIL.n37 104.615
R1431 VTAIL.n38 VTAIL.n27 104.615
R1432 VTAIL.n45 VTAIL.n27 104.615
R1433 VTAIL.n46 VTAIL.n45 104.615
R1434 VTAIL.n46 VTAIL.n23 104.615
R1435 VTAIL.n53 VTAIL.n23 104.615
R1436 VTAIL.n54 VTAIL.n53 104.615
R1437 VTAIL.n54 VTAIL.n19 104.615
R1438 VTAIL.n61 VTAIL.n19 104.615
R1439 VTAIL.n62 VTAIL.n61 104.615
R1440 VTAIL.n62 VTAIL.n15 104.615
R1441 VTAIL.n69 VTAIL.n15 104.615
R1442 VTAIL.n70 VTAIL.n69 104.615
R1443 VTAIL.n70 VTAIL.n11 104.615
R1444 VTAIL.n78 VTAIL.n11 104.615
R1445 VTAIL.n79 VTAIL.n78 104.615
R1446 VTAIL.n80 VTAIL.n79 104.615
R1447 VTAIL.n80 VTAIL.n7 104.615
R1448 VTAIL.n87 VTAIL.n7 104.615
R1449 VTAIL.n88 VTAIL.n87 104.615
R1450 VTAIL.n88 VTAIL.n3 104.615
R1451 VTAIL.n95 VTAIL.n3 104.615
R1452 VTAIL.n96 VTAIL.n95 104.615
R1453 VTAIL.n300 VTAIL.n299 104.615
R1454 VTAIL.n299 VTAIL.n207 104.615
R1455 VTAIL.n292 VTAIL.n207 104.615
R1456 VTAIL.n292 VTAIL.n291 104.615
R1457 VTAIL.n291 VTAIL.n211 104.615
R1458 VTAIL.n284 VTAIL.n211 104.615
R1459 VTAIL.n284 VTAIL.n283 104.615
R1460 VTAIL.n283 VTAIL.n282 104.615
R1461 VTAIL.n282 VTAIL.n215 104.615
R1462 VTAIL.n275 VTAIL.n215 104.615
R1463 VTAIL.n275 VTAIL.n274 104.615
R1464 VTAIL.n274 VTAIL.n220 104.615
R1465 VTAIL.n267 VTAIL.n220 104.615
R1466 VTAIL.n267 VTAIL.n266 104.615
R1467 VTAIL.n266 VTAIL.n224 104.615
R1468 VTAIL.n259 VTAIL.n224 104.615
R1469 VTAIL.n259 VTAIL.n258 104.615
R1470 VTAIL.n258 VTAIL.n228 104.615
R1471 VTAIL.n251 VTAIL.n228 104.615
R1472 VTAIL.n251 VTAIL.n250 104.615
R1473 VTAIL.n250 VTAIL.n232 104.615
R1474 VTAIL.n243 VTAIL.n232 104.615
R1475 VTAIL.n243 VTAIL.n242 104.615
R1476 VTAIL.n242 VTAIL.n236 104.615
R1477 VTAIL.n198 VTAIL.n197 104.615
R1478 VTAIL.n197 VTAIL.n105 104.615
R1479 VTAIL.n190 VTAIL.n105 104.615
R1480 VTAIL.n190 VTAIL.n189 104.615
R1481 VTAIL.n189 VTAIL.n109 104.615
R1482 VTAIL.n182 VTAIL.n109 104.615
R1483 VTAIL.n182 VTAIL.n181 104.615
R1484 VTAIL.n181 VTAIL.n180 104.615
R1485 VTAIL.n180 VTAIL.n113 104.615
R1486 VTAIL.n173 VTAIL.n113 104.615
R1487 VTAIL.n173 VTAIL.n172 104.615
R1488 VTAIL.n172 VTAIL.n118 104.615
R1489 VTAIL.n165 VTAIL.n118 104.615
R1490 VTAIL.n165 VTAIL.n164 104.615
R1491 VTAIL.n164 VTAIL.n122 104.615
R1492 VTAIL.n157 VTAIL.n122 104.615
R1493 VTAIL.n157 VTAIL.n156 104.615
R1494 VTAIL.n156 VTAIL.n126 104.615
R1495 VTAIL.n149 VTAIL.n126 104.615
R1496 VTAIL.n149 VTAIL.n148 104.615
R1497 VTAIL.n148 VTAIL.n130 104.615
R1498 VTAIL.n141 VTAIL.n130 104.615
R1499 VTAIL.n141 VTAIL.n140 104.615
R1500 VTAIL.n140 VTAIL.n134 104.615
R1501 VTAIL.t3 VTAIL.n337 52.3082
R1502 VTAIL.t1 VTAIL.n31 52.3082
R1503 VTAIL.t0 VTAIL.n236 52.3082
R1504 VTAIL.t2 VTAIL.n134 52.3082
R1505 VTAIL.n407 VTAIL.n406 30.052
R1506 VTAIL.n101 VTAIL.n100 30.052
R1507 VTAIL.n305 VTAIL.n304 30.052
R1508 VTAIL.n203 VTAIL.n202 30.052
R1509 VTAIL.n203 VTAIL.n101 29.3238
R1510 VTAIL.n407 VTAIL.n305 28.6686
R1511 VTAIL.n339 VTAIL.n338 15.6677
R1512 VTAIL.n33 VTAIL.n32 15.6677
R1513 VTAIL.n238 VTAIL.n237 15.6677
R1514 VTAIL.n136 VTAIL.n135 15.6677
R1515 VTAIL.n387 VTAIL.n316 13.1884
R1516 VTAIL.n81 VTAIL.n10 13.1884
R1517 VTAIL.n285 VTAIL.n214 13.1884
R1518 VTAIL.n183 VTAIL.n112 13.1884
R1519 VTAIL.n342 VTAIL.n341 12.8005
R1520 VTAIL.n383 VTAIL.n382 12.8005
R1521 VTAIL.n388 VTAIL.n314 12.8005
R1522 VTAIL.n36 VTAIL.n35 12.8005
R1523 VTAIL.n77 VTAIL.n76 12.8005
R1524 VTAIL.n82 VTAIL.n8 12.8005
R1525 VTAIL.n286 VTAIL.n212 12.8005
R1526 VTAIL.n281 VTAIL.n216 12.8005
R1527 VTAIL.n241 VTAIL.n240 12.8005
R1528 VTAIL.n184 VTAIL.n110 12.8005
R1529 VTAIL.n179 VTAIL.n114 12.8005
R1530 VTAIL.n139 VTAIL.n138 12.8005
R1531 VTAIL.n345 VTAIL.n336 12.0247
R1532 VTAIL.n381 VTAIL.n318 12.0247
R1533 VTAIL.n392 VTAIL.n391 12.0247
R1534 VTAIL.n39 VTAIL.n30 12.0247
R1535 VTAIL.n75 VTAIL.n12 12.0247
R1536 VTAIL.n86 VTAIL.n85 12.0247
R1537 VTAIL.n290 VTAIL.n289 12.0247
R1538 VTAIL.n280 VTAIL.n217 12.0247
R1539 VTAIL.n244 VTAIL.n235 12.0247
R1540 VTAIL.n188 VTAIL.n187 12.0247
R1541 VTAIL.n178 VTAIL.n115 12.0247
R1542 VTAIL.n142 VTAIL.n133 12.0247
R1543 VTAIL.n346 VTAIL.n334 11.249
R1544 VTAIL.n378 VTAIL.n377 11.249
R1545 VTAIL.n395 VTAIL.n312 11.249
R1546 VTAIL.n40 VTAIL.n28 11.249
R1547 VTAIL.n72 VTAIL.n71 11.249
R1548 VTAIL.n89 VTAIL.n6 11.249
R1549 VTAIL.n293 VTAIL.n210 11.249
R1550 VTAIL.n277 VTAIL.n276 11.249
R1551 VTAIL.n245 VTAIL.n233 11.249
R1552 VTAIL.n191 VTAIL.n108 11.249
R1553 VTAIL.n175 VTAIL.n174 11.249
R1554 VTAIL.n143 VTAIL.n131 11.249
R1555 VTAIL.n350 VTAIL.n349 10.4732
R1556 VTAIL.n374 VTAIL.n320 10.4732
R1557 VTAIL.n396 VTAIL.n310 10.4732
R1558 VTAIL.n44 VTAIL.n43 10.4732
R1559 VTAIL.n68 VTAIL.n14 10.4732
R1560 VTAIL.n90 VTAIL.n4 10.4732
R1561 VTAIL.n294 VTAIL.n208 10.4732
R1562 VTAIL.n273 VTAIL.n219 10.4732
R1563 VTAIL.n249 VTAIL.n248 10.4732
R1564 VTAIL.n192 VTAIL.n106 10.4732
R1565 VTAIL.n171 VTAIL.n117 10.4732
R1566 VTAIL.n147 VTAIL.n146 10.4732
R1567 VTAIL.n353 VTAIL.n332 9.69747
R1568 VTAIL.n373 VTAIL.n322 9.69747
R1569 VTAIL.n400 VTAIL.n399 9.69747
R1570 VTAIL.n47 VTAIL.n26 9.69747
R1571 VTAIL.n67 VTAIL.n16 9.69747
R1572 VTAIL.n94 VTAIL.n93 9.69747
R1573 VTAIL.n298 VTAIL.n297 9.69747
R1574 VTAIL.n272 VTAIL.n221 9.69747
R1575 VTAIL.n252 VTAIL.n231 9.69747
R1576 VTAIL.n196 VTAIL.n195 9.69747
R1577 VTAIL.n170 VTAIL.n119 9.69747
R1578 VTAIL.n150 VTAIL.n129 9.69747
R1579 VTAIL.n406 VTAIL.n405 9.45567
R1580 VTAIL.n100 VTAIL.n99 9.45567
R1581 VTAIL.n304 VTAIL.n303 9.45567
R1582 VTAIL.n202 VTAIL.n201 9.45567
R1583 VTAIL.n405 VTAIL.n404 9.3005
R1584 VTAIL.n308 VTAIL.n307 9.3005
R1585 VTAIL.n399 VTAIL.n398 9.3005
R1586 VTAIL.n397 VTAIL.n396 9.3005
R1587 VTAIL.n312 VTAIL.n311 9.3005
R1588 VTAIL.n391 VTAIL.n390 9.3005
R1589 VTAIL.n389 VTAIL.n388 9.3005
R1590 VTAIL.n328 VTAIL.n327 9.3005
R1591 VTAIL.n357 VTAIL.n356 9.3005
R1592 VTAIL.n355 VTAIL.n354 9.3005
R1593 VTAIL.n332 VTAIL.n331 9.3005
R1594 VTAIL.n349 VTAIL.n348 9.3005
R1595 VTAIL.n347 VTAIL.n346 9.3005
R1596 VTAIL.n336 VTAIL.n335 9.3005
R1597 VTAIL.n341 VTAIL.n340 9.3005
R1598 VTAIL.n363 VTAIL.n362 9.3005
R1599 VTAIL.n365 VTAIL.n364 9.3005
R1600 VTAIL.n324 VTAIL.n323 9.3005
R1601 VTAIL.n371 VTAIL.n370 9.3005
R1602 VTAIL.n373 VTAIL.n372 9.3005
R1603 VTAIL.n320 VTAIL.n319 9.3005
R1604 VTAIL.n379 VTAIL.n378 9.3005
R1605 VTAIL.n381 VTAIL.n380 9.3005
R1606 VTAIL.n382 VTAIL.n315 9.3005
R1607 VTAIL.n99 VTAIL.n98 9.3005
R1608 VTAIL.n2 VTAIL.n1 9.3005
R1609 VTAIL.n93 VTAIL.n92 9.3005
R1610 VTAIL.n91 VTAIL.n90 9.3005
R1611 VTAIL.n6 VTAIL.n5 9.3005
R1612 VTAIL.n85 VTAIL.n84 9.3005
R1613 VTAIL.n83 VTAIL.n82 9.3005
R1614 VTAIL.n22 VTAIL.n21 9.3005
R1615 VTAIL.n51 VTAIL.n50 9.3005
R1616 VTAIL.n49 VTAIL.n48 9.3005
R1617 VTAIL.n26 VTAIL.n25 9.3005
R1618 VTAIL.n43 VTAIL.n42 9.3005
R1619 VTAIL.n41 VTAIL.n40 9.3005
R1620 VTAIL.n30 VTAIL.n29 9.3005
R1621 VTAIL.n35 VTAIL.n34 9.3005
R1622 VTAIL.n57 VTAIL.n56 9.3005
R1623 VTAIL.n59 VTAIL.n58 9.3005
R1624 VTAIL.n18 VTAIL.n17 9.3005
R1625 VTAIL.n65 VTAIL.n64 9.3005
R1626 VTAIL.n67 VTAIL.n66 9.3005
R1627 VTAIL.n14 VTAIL.n13 9.3005
R1628 VTAIL.n73 VTAIL.n72 9.3005
R1629 VTAIL.n75 VTAIL.n74 9.3005
R1630 VTAIL.n76 VTAIL.n9 9.3005
R1631 VTAIL.n264 VTAIL.n263 9.3005
R1632 VTAIL.n223 VTAIL.n222 9.3005
R1633 VTAIL.n270 VTAIL.n269 9.3005
R1634 VTAIL.n272 VTAIL.n271 9.3005
R1635 VTAIL.n219 VTAIL.n218 9.3005
R1636 VTAIL.n278 VTAIL.n277 9.3005
R1637 VTAIL.n280 VTAIL.n279 9.3005
R1638 VTAIL.n216 VTAIL.n213 9.3005
R1639 VTAIL.n303 VTAIL.n302 9.3005
R1640 VTAIL.n206 VTAIL.n205 9.3005
R1641 VTAIL.n297 VTAIL.n296 9.3005
R1642 VTAIL.n295 VTAIL.n294 9.3005
R1643 VTAIL.n210 VTAIL.n209 9.3005
R1644 VTAIL.n289 VTAIL.n288 9.3005
R1645 VTAIL.n287 VTAIL.n286 9.3005
R1646 VTAIL.n262 VTAIL.n261 9.3005
R1647 VTAIL.n227 VTAIL.n226 9.3005
R1648 VTAIL.n256 VTAIL.n255 9.3005
R1649 VTAIL.n254 VTAIL.n253 9.3005
R1650 VTAIL.n231 VTAIL.n230 9.3005
R1651 VTAIL.n248 VTAIL.n247 9.3005
R1652 VTAIL.n246 VTAIL.n245 9.3005
R1653 VTAIL.n235 VTAIL.n234 9.3005
R1654 VTAIL.n240 VTAIL.n239 9.3005
R1655 VTAIL.n162 VTAIL.n161 9.3005
R1656 VTAIL.n121 VTAIL.n120 9.3005
R1657 VTAIL.n168 VTAIL.n167 9.3005
R1658 VTAIL.n170 VTAIL.n169 9.3005
R1659 VTAIL.n117 VTAIL.n116 9.3005
R1660 VTAIL.n176 VTAIL.n175 9.3005
R1661 VTAIL.n178 VTAIL.n177 9.3005
R1662 VTAIL.n114 VTAIL.n111 9.3005
R1663 VTAIL.n201 VTAIL.n200 9.3005
R1664 VTAIL.n104 VTAIL.n103 9.3005
R1665 VTAIL.n195 VTAIL.n194 9.3005
R1666 VTAIL.n193 VTAIL.n192 9.3005
R1667 VTAIL.n108 VTAIL.n107 9.3005
R1668 VTAIL.n187 VTAIL.n186 9.3005
R1669 VTAIL.n185 VTAIL.n184 9.3005
R1670 VTAIL.n160 VTAIL.n159 9.3005
R1671 VTAIL.n125 VTAIL.n124 9.3005
R1672 VTAIL.n154 VTAIL.n153 9.3005
R1673 VTAIL.n152 VTAIL.n151 9.3005
R1674 VTAIL.n129 VTAIL.n128 9.3005
R1675 VTAIL.n146 VTAIL.n145 9.3005
R1676 VTAIL.n144 VTAIL.n143 9.3005
R1677 VTAIL.n133 VTAIL.n132 9.3005
R1678 VTAIL.n138 VTAIL.n137 9.3005
R1679 VTAIL.n354 VTAIL.n330 8.92171
R1680 VTAIL.n370 VTAIL.n369 8.92171
R1681 VTAIL.n403 VTAIL.n308 8.92171
R1682 VTAIL.n48 VTAIL.n24 8.92171
R1683 VTAIL.n64 VTAIL.n63 8.92171
R1684 VTAIL.n97 VTAIL.n2 8.92171
R1685 VTAIL.n301 VTAIL.n206 8.92171
R1686 VTAIL.n269 VTAIL.n268 8.92171
R1687 VTAIL.n253 VTAIL.n229 8.92171
R1688 VTAIL.n199 VTAIL.n104 8.92171
R1689 VTAIL.n167 VTAIL.n166 8.92171
R1690 VTAIL.n151 VTAIL.n127 8.92171
R1691 VTAIL.n358 VTAIL.n357 8.14595
R1692 VTAIL.n366 VTAIL.n324 8.14595
R1693 VTAIL.n404 VTAIL.n306 8.14595
R1694 VTAIL.n52 VTAIL.n51 8.14595
R1695 VTAIL.n60 VTAIL.n18 8.14595
R1696 VTAIL.n98 VTAIL.n0 8.14595
R1697 VTAIL.n302 VTAIL.n204 8.14595
R1698 VTAIL.n265 VTAIL.n223 8.14595
R1699 VTAIL.n257 VTAIL.n256 8.14595
R1700 VTAIL.n200 VTAIL.n102 8.14595
R1701 VTAIL.n163 VTAIL.n121 8.14595
R1702 VTAIL.n155 VTAIL.n154 8.14595
R1703 VTAIL.n361 VTAIL.n328 7.3702
R1704 VTAIL.n365 VTAIL.n326 7.3702
R1705 VTAIL.n55 VTAIL.n22 7.3702
R1706 VTAIL.n59 VTAIL.n20 7.3702
R1707 VTAIL.n264 VTAIL.n225 7.3702
R1708 VTAIL.n260 VTAIL.n227 7.3702
R1709 VTAIL.n162 VTAIL.n123 7.3702
R1710 VTAIL.n158 VTAIL.n125 7.3702
R1711 VTAIL.n362 VTAIL.n361 6.59444
R1712 VTAIL.n362 VTAIL.n326 6.59444
R1713 VTAIL.n56 VTAIL.n55 6.59444
R1714 VTAIL.n56 VTAIL.n20 6.59444
R1715 VTAIL.n261 VTAIL.n225 6.59444
R1716 VTAIL.n261 VTAIL.n260 6.59444
R1717 VTAIL.n159 VTAIL.n123 6.59444
R1718 VTAIL.n159 VTAIL.n158 6.59444
R1719 VTAIL.n358 VTAIL.n328 5.81868
R1720 VTAIL.n366 VTAIL.n365 5.81868
R1721 VTAIL.n406 VTAIL.n306 5.81868
R1722 VTAIL.n52 VTAIL.n22 5.81868
R1723 VTAIL.n60 VTAIL.n59 5.81868
R1724 VTAIL.n100 VTAIL.n0 5.81868
R1725 VTAIL.n304 VTAIL.n204 5.81868
R1726 VTAIL.n265 VTAIL.n264 5.81868
R1727 VTAIL.n257 VTAIL.n227 5.81868
R1728 VTAIL.n202 VTAIL.n102 5.81868
R1729 VTAIL.n163 VTAIL.n162 5.81868
R1730 VTAIL.n155 VTAIL.n125 5.81868
R1731 VTAIL.n357 VTAIL.n330 5.04292
R1732 VTAIL.n369 VTAIL.n324 5.04292
R1733 VTAIL.n404 VTAIL.n403 5.04292
R1734 VTAIL.n51 VTAIL.n24 5.04292
R1735 VTAIL.n63 VTAIL.n18 5.04292
R1736 VTAIL.n98 VTAIL.n97 5.04292
R1737 VTAIL.n302 VTAIL.n301 5.04292
R1738 VTAIL.n268 VTAIL.n223 5.04292
R1739 VTAIL.n256 VTAIL.n229 5.04292
R1740 VTAIL.n200 VTAIL.n199 5.04292
R1741 VTAIL.n166 VTAIL.n121 5.04292
R1742 VTAIL.n154 VTAIL.n127 5.04292
R1743 VTAIL.n340 VTAIL.n339 4.38563
R1744 VTAIL.n34 VTAIL.n33 4.38563
R1745 VTAIL.n239 VTAIL.n238 4.38563
R1746 VTAIL.n137 VTAIL.n136 4.38563
R1747 VTAIL.n354 VTAIL.n353 4.26717
R1748 VTAIL.n370 VTAIL.n322 4.26717
R1749 VTAIL.n400 VTAIL.n308 4.26717
R1750 VTAIL.n48 VTAIL.n47 4.26717
R1751 VTAIL.n64 VTAIL.n16 4.26717
R1752 VTAIL.n94 VTAIL.n2 4.26717
R1753 VTAIL.n298 VTAIL.n206 4.26717
R1754 VTAIL.n269 VTAIL.n221 4.26717
R1755 VTAIL.n253 VTAIL.n252 4.26717
R1756 VTAIL.n196 VTAIL.n104 4.26717
R1757 VTAIL.n167 VTAIL.n119 4.26717
R1758 VTAIL.n151 VTAIL.n150 4.26717
R1759 VTAIL.n350 VTAIL.n332 3.49141
R1760 VTAIL.n374 VTAIL.n373 3.49141
R1761 VTAIL.n399 VTAIL.n310 3.49141
R1762 VTAIL.n44 VTAIL.n26 3.49141
R1763 VTAIL.n68 VTAIL.n67 3.49141
R1764 VTAIL.n93 VTAIL.n4 3.49141
R1765 VTAIL.n297 VTAIL.n208 3.49141
R1766 VTAIL.n273 VTAIL.n272 3.49141
R1767 VTAIL.n249 VTAIL.n231 3.49141
R1768 VTAIL.n195 VTAIL.n106 3.49141
R1769 VTAIL.n171 VTAIL.n170 3.49141
R1770 VTAIL.n147 VTAIL.n129 3.49141
R1771 VTAIL.n349 VTAIL.n334 2.71565
R1772 VTAIL.n377 VTAIL.n320 2.71565
R1773 VTAIL.n396 VTAIL.n395 2.71565
R1774 VTAIL.n43 VTAIL.n28 2.71565
R1775 VTAIL.n71 VTAIL.n14 2.71565
R1776 VTAIL.n90 VTAIL.n89 2.71565
R1777 VTAIL.n294 VTAIL.n293 2.71565
R1778 VTAIL.n276 VTAIL.n219 2.71565
R1779 VTAIL.n248 VTAIL.n233 2.71565
R1780 VTAIL.n192 VTAIL.n191 2.71565
R1781 VTAIL.n174 VTAIL.n117 2.71565
R1782 VTAIL.n146 VTAIL.n131 2.71565
R1783 VTAIL.n346 VTAIL.n345 1.93989
R1784 VTAIL.n378 VTAIL.n318 1.93989
R1785 VTAIL.n392 VTAIL.n312 1.93989
R1786 VTAIL.n40 VTAIL.n39 1.93989
R1787 VTAIL.n72 VTAIL.n12 1.93989
R1788 VTAIL.n86 VTAIL.n6 1.93989
R1789 VTAIL.n290 VTAIL.n210 1.93989
R1790 VTAIL.n277 VTAIL.n217 1.93989
R1791 VTAIL.n245 VTAIL.n244 1.93989
R1792 VTAIL.n188 VTAIL.n108 1.93989
R1793 VTAIL.n175 VTAIL.n115 1.93989
R1794 VTAIL.n143 VTAIL.n142 1.93989
R1795 VTAIL.n342 VTAIL.n336 1.16414
R1796 VTAIL.n383 VTAIL.n381 1.16414
R1797 VTAIL.n391 VTAIL.n314 1.16414
R1798 VTAIL.n36 VTAIL.n30 1.16414
R1799 VTAIL.n77 VTAIL.n75 1.16414
R1800 VTAIL.n85 VTAIL.n8 1.16414
R1801 VTAIL.n289 VTAIL.n212 1.16414
R1802 VTAIL.n281 VTAIL.n280 1.16414
R1803 VTAIL.n241 VTAIL.n235 1.16414
R1804 VTAIL.n187 VTAIL.n110 1.16414
R1805 VTAIL.n179 VTAIL.n178 1.16414
R1806 VTAIL.n139 VTAIL.n133 1.16414
R1807 VTAIL.n305 VTAIL.n203 0.797914
R1808 VTAIL VTAIL.n101 0.69231
R1809 VTAIL.n341 VTAIL.n338 0.388379
R1810 VTAIL.n382 VTAIL.n316 0.388379
R1811 VTAIL.n388 VTAIL.n387 0.388379
R1812 VTAIL.n35 VTAIL.n32 0.388379
R1813 VTAIL.n76 VTAIL.n10 0.388379
R1814 VTAIL.n82 VTAIL.n81 0.388379
R1815 VTAIL.n286 VTAIL.n285 0.388379
R1816 VTAIL.n216 VTAIL.n214 0.388379
R1817 VTAIL.n240 VTAIL.n237 0.388379
R1818 VTAIL.n184 VTAIL.n183 0.388379
R1819 VTAIL.n114 VTAIL.n112 0.388379
R1820 VTAIL.n138 VTAIL.n135 0.388379
R1821 VTAIL.n340 VTAIL.n335 0.155672
R1822 VTAIL.n347 VTAIL.n335 0.155672
R1823 VTAIL.n348 VTAIL.n347 0.155672
R1824 VTAIL.n348 VTAIL.n331 0.155672
R1825 VTAIL.n355 VTAIL.n331 0.155672
R1826 VTAIL.n356 VTAIL.n355 0.155672
R1827 VTAIL.n356 VTAIL.n327 0.155672
R1828 VTAIL.n363 VTAIL.n327 0.155672
R1829 VTAIL.n364 VTAIL.n363 0.155672
R1830 VTAIL.n364 VTAIL.n323 0.155672
R1831 VTAIL.n371 VTAIL.n323 0.155672
R1832 VTAIL.n372 VTAIL.n371 0.155672
R1833 VTAIL.n372 VTAIL.n319 0.155672
R1834 VTAIL.n379 VTAIL.n319 0.155672
R1835 VTAIL.n380 VTAIL.n379 0.155672
R1836 VTAIL.n380 VTAIL.n315 0.155672
R1837 VTAIL.n389 VTAIL.n315 0.155672
R1838 VTAIL.n390 VTAIL.n389 0.155672
R1839 VTAIL.n390 VTAIL.n311 0.155672
R1840 VTAIL.n397 VTAIL.n311 0.155672
R1841 VTAIL.n398 VTAIL.n397 0.155672
R1842 VTAIL.n398 VTAIL.n307 0.155672
R1843 VTAIL.n405 VTAIL.n307 0.155672
R1844 VTAIL.n34 VTAIL.n29 0.155672
R1845 VTAIL.n41 VTAIL.n29 0.155672
R1846 VTAIL.n42 VTAIL.n41 0.155672
R1847 VTAIL.n42 VTAIL.n25 0.155672
R1848 VTAIL.n49 VTAIL.n25 0.155672
R1849 VTAIL.n50 VTAIL.n49 0.155672
R1850 VTAIL.n50 VTAIL.n21 0.155672
R1851 VTAIL.n57 VTAIL.n21 0.155672
R1852 VTAIL.n58 VTAIL.n57 0.155672
R1853 VTAIL.n58 VTAIL.n17 0.155672
R1854 VTAIL.n65 VTAIL.n17 0.155672
R1855 VTAIL.n66 VTAIL.n65 0.155672
R1856 VTAIL.n66 VTAIL.n13 0.155672
R1857 VTAIL.n73 VTAIL.n13 0.155672
R1858 VTAIL.n74 VTAIL.n73 0.155672
R1859 VTAIL.n74 VTAIL.n9 0.155672
R1860 VTAIL.n83 VTAIL.n9 0.155672
R1861 VTAIL.n84 VTAIL.n83 0.155672
R1862 VTAIL.n84 VTAIL.n5 0.155672
R1863 VTAIL.n91 VTAIL.n5 0.155672
R1864 VTAIL.n92 VTAIL.n91 0.155672
R1865 VTAIL.n92 VTAIL.n1 0.155672
R1866 VTAIL.n99 VTAIL.n1 0.155672
R1867 VTAIL.n303 VTAIL.n205 0.155672
R1868 VTAIL.n296 VTAIL.n205 0.155672
R1869 VTAIL.n296 VTAIL.n295 0.155672
R1870 VTAIL.n295 VTAIL.n209 0.155672
R1871 VTAIL.n288 VTAIL.n209 0.155672
R1872 VTAIL.n288 VTAIL.n287 0.155672
R1873 VTAIL.n287 VTAIL.n213 0.155672
R1874 VTAIL.n279 VTAIL.n213 0.155672
R1875 VTAIL.n279 VTAIL.n278 0.155672
R1876 VTAIL.n278 VTAIL.n218 0.155672
R1877 VTAIL.n271 VTAIL.n218 0.155672
R1878 VTAIL.n271 VTAIL.n270 0.155672
R1879 VTAIL.n270 VTAIL.n222 0.155672
R1880 VTAIL.n263 VTAIL.n222 0.155672
R1881 VTAIL.n263 VTAIL.n262 0.155672
R1882 VTAIL.n262 VTAIL.n226 0.155672
R1883 VTAIL.n255 VTAIL.n226 0.155672
R1884 VTAIL.n255 VTAIL.n254 0.155672
R1885 VTAIL.n254 VTAIL.n230 0.155672
R1886 VTAIL.n247 VTAIL.n230 0.155672
R1887 VTAIL.n247 VTAIL.n246 0.155672
R1888 VTAIL.n246 VTAIL.n234 0.155672
R1889 VTAIL.n239 VTAIL.n234 0.155672
R1890 VTAIL.n201 VTAIL.n103 0.155672
R1891 VTAIL.n194 VTAIL.n103 0.155672
R1892 VTAIL.n194 VTAIL.n193 0.155672
R1893 VTAIL.n193 VTAIL.n107 0.155672
R1894 VTAIL.n186 VTAIL.n107 0.155672
R1895 VTAIL.n186 VTAIL.n185 0.155672
R1896 VTAIL.n185 VTAIL.n111 0.155672
R1897 VTAIL.n177 VTAIL.n111 0.155672
R1898 VTAIL.n177 VTAIL.n176 0.155672
R1899 VTAIL.n176 VTAIL.n116 0.155672
R1900 VTAIL.n169 VTAIL.n116 0.155672
R1901 VTAIL.n169 VTAIL.n168 0.155672
R1902 VTAIL.n168 VTAIL.n120 0.155672
R1903 VTAIL.n161 VTAIL.n120 0.155672
R1904 VTAIL.n161 VTAIL.n160 0.155672
R1905 VTAIL.n160 VTAIL.n124 0.155672
R1906 VTAIL.n153 VTAIL.n124 0.155672
R1907 VTAIL.n153 VTAIL.n152 0.155672
R1908 VTAIL.n152 VTAIL.n128 0.155672
R1909 VTAIL.n145 VTAIL.n128 0.155672
R1910 VTAIL.n145 VTAIL.n144 0.155672
R1911 VTAIL.n144 VTAIL.n132 0.155672
R1912 VTAIL.n137 VTAIL.n132 0.155672
R1913 VTAIL VTAIL.n407 0.106103
R1914 VDD2.n197 VDD2.n101 289.615
R1915 VDD2.n96 VDD2.n0 289.615
R1916 VDD2.n198 VDD2.n197 185
R1917 VDD2.n196 VDD2.n195 185
R1918 VDD2.n105 VDD2.n104 185
R1919 VDD2.n190 VDD2.n189 185
R1920 VDD2.n188 VDD2.n187 185
R1921 VDD2.n109 VDD2.n108 185
R1922 VDD2.n182 VDD2.n181 185
R1923 VDD2.n180 VDD2.n111 185
R1924 VDD2.n179 VDD2.n178 185
R1925 VDD2.n114 VDD2.n112 185
R1926 VDD2.n173 VDD2.n172 185
R1927 VDD2.n171 VDD2.n170 185
R1928 VDD2.n118 VDD2.n117 185
R1929 VDD2.n165 VDD2.n164 185
R1930 VDD2.n163 VDD2.n162 185
R1931 VDD2.n122 VDD2.n121 185
R1932 VDD2.n157 VDD2.n156 185
R1933 VDD2.n155 VDD2.n154 185
R1934 VDD2.n126 VDD2.n125 185
R1935 VDD2.n149 VDD2.n148 185
R1936 VDD2.n147 VDD2.n146 185
R1937 VDD2.n130 VDD2.n129 185
R1938 VDD2.n141 VDD2.n140 185
R1939 VDD2.n139 VDD2.n138 185
R1940 VDD2.n134 VDD2.n133 185
R1941 VDD2.n32 VDD2.n31 185
R1942 VDD2.n37 VDD2.n36 185
R1943 VDD2.n39 VDD2.n38 185
R1944 VDD2.n28 VDD2.n27 185
R1945 VDD2.n45 VDD2.n44 185
R1946 VDD2.n47 VDD2.n46 185
R1947 VDD2.n24 VDD2.n23 185
R1948 VDD2.n53 VDD2.n52 185
R1949 VDD2.n55 VDD2.n54 185
R1950 VDD2.n20 VDD2.n19 185
R1951 VDD2.n61 VDD2.n60 185
R1952 VDD2.n63 VDD2.n62 185
R1953 VDD2.n16 VDD2.n15 185
R1954 VDD2.n69 VDD2.n68 185
R1955 VDD2.n71 VDD2.n70 185
R1956 VDD2.n12 VDD2.n11 185
R1957 VDD2.n78 VDD2.n77 185
R1958 VDD2.n79 VDD2.n10 185
R1959 VDD2.n81 VDD2.n80 185
R1960 VDD2.n8 VDD2.n7 185
R1961 VDD2.n87 VDD2.n86 185
R1962 VDD2.n89 VDD2.n88 185
R1963 VDD2.n4 VDD2.n3 185
R1964 VDD2.n95 VDD2.n94 185
R1965 VDD2.n97 VDD2.n96 185
R1966 VDD2.n135 VDD2.t1 147.659
R1967 VDD2.n33 VDD2.t0 147.659
R1968 VDD2.n197 VDD2.n196 104.615
R1969 VDD2.n196 VDD2.n104 104.615
R1970 VDD2.n189 VDD2.n104 104.615
R1971 VDD2.n189 VDD2.n188 104.615
R1972 VDD2.n188 VDD2.n108 104.615
R1973 VDD2.n181 VDD2.n108 104.615
R1974 VDD2.n181 VDD2.n180 104.615
R1975 VDD2.n180 VDD2.n179 104.615
R1976 VDD2.n179 VDD2.n112 104.615
R1977 VDD2.n172 VDD2.n112 104.615
R1978 VDD2.n172 VDD2.n171 104.615
R1979 VDD2.n171 VDD2.n117 104.615
R1980 VDD2.n164 VDD2.n117 104.615
R1981 VDD2.n164 VDD2.n163 104.615
R1982 VDD2.n163 VDD2.n121 104.615
R1983 VDD2.n156 VDD2.n121 104.615
R1984 VDD2.n156 VDD2.n155 104.615
R1985 VDD2.n155 VDD2.n125 104.615
R1986 VDD2.n148 VDD2.n125 104.615
R1987 VDD2.n148 VDD2.n147 104.615
R1988 VDD2.n147 VDD2.n129 104.615
R1989 VDD2.n140 VDD2.n129 104.615
R1990 VDD2.n140 VDD2.n139 104.615
R1991 VDD2.n139 VDD2.n133 104.615
R1992 VDD2.n37 VDD2.n31 104.615
R1993 VDD2.n38 VDD2.n37 104.615
R1994 VDD2.n38 VDD2.n27 104.615
R1995 VDD2.n45 VDD2.n27 104.615
R1996 VDD2.n46 VDD2.n45 104.615
R1997 VDD2.n46 VDD2.n23 104.615
R1998 VDD2.n53 VDD2.n23 104.615
R1999 VDD2.n54 VDD2.n53 104.615
R2000 VDD2.n54 VDD2.n19 104.615
R2001 VDD2.n61 VDD2.n19 104.615
R2002 VDD2.n62 VDD2.n61 104.615
R2003 VDD2.n62 VDD2.n15 104.615
R2004 VDD2.n69 VDD2.n15 104.615
R2005 VDD2.n70 VDD2.n69 104.615
R2006 VDD2.n70 VDD2.n11 104.615
R2007 VDD2.n78 VDD2.n11 104.615
R2008 VDD2.n79 VDD2.n78 104.615
R2009 VDD2.n80 VDD2.n79 104.615
R2010 VDD2.n80 VDD2.n7 104.615
R2011 VDD2.n87 VDD2.n7 104.615
R2012 VDD2.n88 VDD2.n87 104.615
R2013 VDD2.n88 VDD2.n3 104.615
R2014 VDD2.n95 VDD2.n3 104.615
R2015 VDD2.n96 VDD2.n95 104.615
R2016 VDD2.n202 VDD2.n100 87.3471
R2017 VDD2.t1 VDD2.n133 52.3082
R2018 VDD2.t0 VDD2.n31 52.3082
R2019 VDD2.n202 VDD2.n201 46.7308
R2020 VDD2.n135 VDD2.n134 15.6677
R2021 VDD2.n33 VDD2.n32 15.6677
R2022 VDD2.n182 VDD2.n111 13.1884
R2023 VDD2.n81 VDD2.n10 13.1884
R2024 VDD2.n183 VDD2.n109 12.8005
R2025 VDD2.n178 VDD2.n113 12.8005
R2026 VDD2.n138 VDD2.n137 12.8005
R2027 VDD2.n36 VDD2.n35 12.8005
R2028 VDD2.n77 VDD2.n76 12.8005
R2029 VDD2.n82 VDD2.n8 12.8005
R2030 VDD2.n187 VDD2.n186 12.0247
R2031 VDD2.n177 VDD2.n114 12.0247
R2032 VDD2.n141 VDD2.n132 12.0247
R2033 VDD2.n39 VDD2.n30 12.0247
R2034 VDD2.n75 VDD2.n12 12.0247
R2035 VDD2.n86 VDD2.n85 12.0247
R2036 VDD2.n190 VDD2.n107 11.249
R2037 VDD2.n174 VDD2.n173 11.249
R2038 VDD2.n142 VDD2.n130 11.249
R2039 VDD2.n40 VDD2.n28 11.249
R2040 VDD2.n72 VDD2.n71 11.249
R2041 VDD2.n89 VDD2.n6 11.249
R2042 VDD2.n191 VDD2.n105 10.4732
R2043 VDD2.n170 VDD2.n116 10.4732
R2044 VDD2.n146 VDD2.n145 10.4732
R2045 VDD2.n44 VDD2.n43 10.4732
R2046 VDD2.n68 VDD2.n14 10.4732
R2047 VDD2.n90 VDD2.n4 10.4732
R2048 VDD2.n195 VDD2.n194 9.69747
R2049 VDD2.n169 VDD2.n118 9.69747
R2050 VDD2.n149 VDD2.n128 9.69747
R2051 VDD2.n47 VDD2.n26 9.69747
R2052 VDD2.n67 VDD2.n16 9.69747
R2053 VDD2.n94 VDD2.n93 9.69747
R2054 VDD2.n201 VDD2.n200 9.45567
R2055 VDD2.n100 VDD2.n99 9.45567
R2056 VDD2.n161 VDD2.n160 9.3005
R2057 VDD2.n120 VDD2.n119 9.3005
R2058 VDD2.n167 VDD2.n166 9.3005
R2059 VDD2.n169 VDD2.n168 9.3005
R2060 VDD2.n116 VDD2.n115 9.3005
R2061 VDD2.n175 VDD2.n174 9.3005
R2062 VDD2.n177 VDD2.n176 9.3005
R2063 VDD2.n113 VDD2.n110 9.3005
R2064 VDD2.n200 VDD2.n199 9.3005
R2065 VDD2.n103 VDD2.n102 9.3005
R2066 VDD2.n194 VDD2.n193 9.3005
R2067 VDD2.n192 VDD2.n191 9.3005
R2068 VDD2.n107 VDD2.n106 9.3005
R2069 VDD2.n186 VDD2.n185 9.3005
R2070 VDD2.n184 VDD2.n183 9.3005
R2071 VDD2.n159 VDD2.n158 9.3005
R2072 VDD2.n124 VDD2.n123 9.3005
R2073 VDD2.n153 VDD2.n152 9.3005
R2074 VDD2.n151 VDD2.n150 9.3005
R2075 VDD2.n128 VDD2.n127 9.3005
R2076 VDD2.n145 VDD2.n144 9.3005
R2077 VDD2.n143 VDD2.n142 9.3005
R2078 VDD2.n132 VDD2.n131 9.3005
R2079 VDD2.n137 VDD2.n136 9.3005
R2080 VDD2.n99 VDD2.n98 9.3005
R2081 VDD2.n2 VDD2.n1 9.3005
R2082 VDD2.n93 VDD2.n92 9.3005
R2083 VDD2.n91 VDD2.n90 9.3005
R2084 VDD2.n6 VDD2.n5 9.3005
R2085 VDD2.n85 VDD2.n84 9.3005
R2086 VDD2.n83 VDD2.n82 9.3005
R2087 VDD2.n22 VDD2.n21 9.3005
R2088 VDD2.n51 VDD2.n50 9.3005
R2089 VDD2.n49 VDD2.n48 9.3005
R2090 VDD2.n26 VDD2.n25 9.3005
R2091 VDD2.n43 VDD2.n42 9.3005
R2092 VDD2.n41 VDD2.n40 9.3005
R2093 VDD2.n30 VDD2.n29 9.3005
R2094 VDD2.n35 VDD2.n34 9.3005
R2095 VDD2.n57 VDD2.n56 9.3005
R2096 VDD2.n59 VDD2.n58 9.3005
R2097 VDD2.n18 VDD2.n17 9.3005
R2098 VDD2.n65 VDD2.n64 9.3005
R2099 VDD2.n67 VDD2.n66 9.3005
R2100 VDD2.n14 VDD2.n13 9.3005
R2101 VDD2.n73 VDD2.n72 9.3005
R2102 VDD2.n75 VDD2.n74 9.3005
R2103 VDD2.n76 VDD2.n9 9.3005
R2104 VDD2.n198 VDD2.n103 8.92171
R2105 VDD2.n166 VDD2.n165 8.92171
R2106 VDD2.n150 VDD2.n126 8.92171
R2107 VDD2.n48 VDD2.n24 8.92171
R2108 VDD2.n64 VDD2.n63 8.92171
R2109 VDD2.n97 VDD2.n2 8.92171
R2110 VDD2.n199 VDD2.n101 8.14595
R2111 VDD2.n162 VDD2.n120 8.14595
R2112 VDD2.n154 VDD2.n153 8.14595
R2113 VDD2.n52 VDD2.n51 8.14595
R2114 VDD2.n60 VDD2.n18 8.14595
R2115 VDD2.n98 VDD2.n0 8.14595
R2116 VDD2.n161 VDD2.n122 7.3702
R2117 VDD2.n157 VDD2.n124 7.3702
R2118 VDD2.n55 VDD2.n22 7.3702
R2119 VDD2.n59 VDD2.n20 7.3702
R2120 VDD2.n158 VDD2.n122 6.59444
R2121 VDD2.n158 VDD2.n157 6.59444
R2122 VDD2.n56 VDD2.n55 6.59444
R2123 VDD2.n56 VDD2.n20 6.59444
R2124 VDD2.n201 VDD2.n101 5.81868
R2125 VDD2.n162 VDD2.n161 5.81868
R2126 VDD2.n154 VDD2.n124 5.81868
R2127 VDD2.n52 VDD2.n22 5.81868
R2128 VDD2.n60 VDD2.n59 5.81868
R2129 VDD2.n100 VDD2.n0 5.81868
R2130 VDD2.n199 VDD2.n198 5.04292
R2131 VDD2.n165 VDD2.n120 5.04292
R2132 VDD2.n153 VDD2.n126 5.04292
R2133 VDD2.n51 VDD2.n24 5.04292
R2134 VDD2.n63 VDD2.n18 5.04292
R2135 VDD2.n98 VDD2.n97 5.04292
R2136 VDD2.n136 VDD2.n135 4.38563
R2137 VDD2.n34 VDD2.n33 4.38563
R2138 VDD2.n195 VDD2.n103 4.26717
R2139 VDD2.n166 VDD2.n118 4.26717
R2140 VDD2.n150 VDD2.n149 4.26717
R2141 VDD2.n48 VDD2.n47 4.26717
R2142 VDD2.n64 VDD2.n16 4.26717
R2143 VDD2.n94 VDD2.n2 4.26717
R2144 VDD2.n194 VDD2.n105 3.49141
R2145 VDD2.n170 VDD2.n169 3.49141
R2146 VDD2.n146 VDD2.n128 3.49141
R2147 VDD2.n44 VDD2.n26 3.49141
R2148 VDD2.n68 VDD2.n67 3.49141
R2149 VDD2.n93 VDD2.n4 3.49141
R2150 VDD2.n191 VDD2.n190 2.71565
R2151 VDD2.n173 VDD2.n116 2.71565
R2152 VDD2.n145 VDD2.n130 2.71565
R2153 VDD2.n43 VDD2.n28 2.71565
R2154 VDD2.n71 VDD2.n14 2.71565
R2155 VDD2.n90 VDD2.n89 2.71565
R2156 VDD2.n187 VDD2.n107 1.93989
R2157 VDD2.n174 VDD2.n114 1.93989
R2158 VDD2.n142 VDD2.n141 1.93989
R2159 VDD2.n40 VDD2.n39 1.93989
R2160 VDD2.n72 VDD2.n12 1.93989
R2161 VDD2.n86 VDD2.n6 1.93989
R2162 VDD2.n186 VDD2.n109 1.16414
R2163 VDD2.n178 VDD2.n177 1.16414
R2164 VDD2.n138 VDD2.n132 1.16414
R2165 VDD2.n36 VDD2.n30 1.16414
R2166 VDD2.n77 VDD2.n75 1.16414
R2167 VDD2.n85 VDD2.n8 1.16414
R2168 VDD2.n183 VDD2.n182 0.388379
R2169 VDD2.n113 VDD2.n111 0.388379
R2170 VDD2.n137 VDD2.n134 0.388379
R2171 VDD2.n35 VDD2.n32 0.388379
R2172 VDD2.n76 VDD2.n10 0.388379
R2173 VDD2.n82 VDD2.n81 0.388379
R2174 VDD2 VDD2.n202 0.222483
R2175 VDD2.n200 VDD2.n102 0.155672
R2176 VDD2.n193 VDD2.n102 0.155672
R2177 VDD2.n193 VDD2.n192 0.155672
R2178 VDD2.n192 VDD2.n106 0.155672
R2179 VDD2.n185 VDD2.n106 0.155672
R2180 VDD2.n185 VDD2.n184 0.155672
R2181 VDD2.n184 VDD2.n110 0.155672
R2182 VDD2.n176 VDD2.n110 0.155672
R2183 VDD2.n176 VDD2.n175 0.155672
R2184 VDD2.n175 VDD2.n115 0.155672
R2185 VDD2.n168 VDD2.n115 0.155672
R2186 VDD2.n168 VDD2.n167 0.155672
R2187 VDD2.n167 VDD2.n119 0.155672
R2188 VDD2.n160 VDD2.n119 0.155672
R2189 VDD2.n160 VDD2.n159 0.155672
R2190 VDD2.n159 VDD2.n123 0.155672
R2191 VDD2.n152 VDD2.n123 0.155672
R2192 VDD2.n152 VDD2.n151 0.155672
R2193 VDD2.n151 VDD2.n127 0.155672
R2194 VDD2.n144 VDD2.n127 0.155672
R2195 VDD2.n144 VDD2.n143 0.155672
R2196 VDD2.n143 VDD2.n131 0.155672
R2197 VDD2.n136 VDD2.n131 0.155672
R2198 VDD2.n34 VDD2.n29 0.155672
R2199 VDD2.n41 VDD2.n29 0.155672
R2200 VDD2.n42 VDD2.n41 0.155672
R2201 VDD2.n42 VDD2.n25 0.155672
R2202 VDD2.n49 VDD2.n25 0.155672
R2203 VDD2.n50 VDD2.n49 0.155672
R2204 VDD2.n50 VDD2.n21 0.155672
R2205 VDD2.n57 VDD2.n21 0.155672
R2206 VDD2.n58 VDD2.n57 0.155672
R2207 VDD2.n58 VDD2.n17 0.155672
R2208 VDD2.n65 VDD2.n17 0.155672
R2209 VDD2.n66 VDD2.n65 0.155672
R2210 VDD2.n66 VDD2.n13 0.155672
R2211 VDD2.n73 VDD2.n13 0.155672
R2212 VDD2.n74 VDD2.n73 0.155672
R2213 VDD2.n74 VDD2.n9 0.155672
R2214 VDD2.n83 VDD2.n9 0.155672
R2215 VDD2.n84 VDD2.n83 0.155672
R2216 VDD2.n84 VDD2.n5 0.155672
R2217 VDD2.n91 VDD2.n5 0.155672
R2218 VDD2.n92 VDD2.n91 0.155672
R2219 VDD2.n92 VDD2.n1 0.155672
R2220 VDD2.n99 VDD2.n1 0.155672
R2221 VP.n0 VP.t1 1312.9
R2222 VP.n0 VP.t0 1269.34
R2223 VP VP.n0 0.0516364
R2224 VDD1.n96 VDD1.n0 289.615
R2225 VDD1.n197 VDD1.n101 289.615
R2226 VDD1.n97 VDD1.n96 185
R2227 VDD1.n95 VDD1.n94 185
R2228 VDD1.n4 VDD1.n3 185
R2229 VDD1.n89 VDD1.n88 185
R2230 VDD1.n87 VDD1.n86 185
R2231 VDD1.n8 VDD1.n7 185
R2232 VDD1.n81 VDD1.n80 185
R2233 VDD1.n79 VDD1.n10 185
R2234 VDD1.n78 VDD1.n77 185
R2235 VDD1.n13 VDD1.n11 185
R2236 VDD1.n72 VDD1.n71 185
R2237 VDD1.n70 VDD1.n69 185
R2238 VDD1.n17 VDD1.n16 185
R2239 VDD1.n64 VDD1.n63 185
R2240 VDD1.n62 VDD1.n61 185
R2241 VDD1.n21 VDD1.n20 185
R2242 VDD1.n56 VDD1.n55 185
R2243 VDD1.n54 VDD1.n53 185
R2244 VDD1.n25 VDD1.n24 185
R2245 VDD1.n48 VDD1.n47 185
R2246 VDD1.n46 VDD1.n45 185
R2247 VDD1.n29 VDD1.n28 185
R2248 VDD1.n40 VDD1.n39 185
R2249 VDD1.n38 VDD1.n37 185
R2250 VDD1.n33 VDD1.n32 185
R2251 VDD1.n133 VDD1.n132 185
R2252 VDD1.n138 VDD1.n137 185
R2253 VDD1.n140 VDD1.n139 185
R2254 VDD1.n129 VDD1.n128 185
R2255 VDD1.n146 VDD1.n145 185
R2256 VDD1.n148 VDD1.n147 185
R2257 VDD1.n125 VDD1.n124 185
R2258 VDD1.n154 VDD1.n153 185
R2259 VDD1.n156 VDD1.n155 185
R2260 VDD1.n121 VDD1.n120 185
R2261 VDD1.n162 VDD1.n161 185
R2262 VDD1.n164 VDD1.n163 185
R2263 VDD1.n117 VDD1.n116 185
R2264 VDD1.n170 VDD1.n169 185
R2265 VDD1.n172 VDD1.n171 185
R2266 VDD1.n113 VDD1.n112 185
R2267 VDD1.n179 VDD1.n178 185
R2268 VDD1.n180 VDD1.n111 185
R2269 VDD1.n182 VDD1.n181 185
R2270 VDD1.n109 VDD1.n108 185
R2271 VDD1.n188 VDD1.n187 185
R2272 VDD1.n190 VDD1.n189 185
R2273 VDD1.n105 VDD1.n104 185
R2274 VDD1.n196 VDD1.n195 185
R2275 VDD1.n198 VDD1.n197 185
R2276 VDD1.n34 VDD1.t0 147.659
R2277 VDD1.n134 VDD1.t1 147.659
R2278 VDD1.n96 VDD1.n95 104.615
R2279 VDD1.n95 VDD1.n3 104.615
R2280 VDD1.n88 VDD1.n3 104.615
R2281 VDD1.n88 VDD1.n87 104.615
R2282 VDD1.n87 VDD1.n7 104.615
R2283 VDD1.n80 VDD1.n7 104.615
R2284 VDD1.n80 VDD1.n79 104.615
R2285 VDD1.n79 VDD1.n78 104.615
R2286 VDD1.n78 VDD1.n11 104.615
R2287 VDD1.n71 VDD1.n11 104.615
R2288 VDD1.n71 VDD1.n70 104.615
R2289 VDD1.n70 VDD1.n16 104.615
R2290 VDD1.n63 VDD1.n16 104.615
R2291 VDD1.n63 VDD1.n62 104.615
R2292 VDD1.n62 VDD1.n20 104.615
R2293 VDD1.n55 VDD1.n20 104.615
R2294 VDD1.n55 VDD1.n54 104.615
R2295 VDD1.n54 VDD1.n24 104.615
R2296 VDD1.n47 VDD1.n24 104.615
R2297 VDD1.n47 VDD1.n46 104.615
R2298 VDD1.n46 VDD1.n28 104.615
R2299 VDD1.n39 VDD1.n28 104.615
R2300 VDD1.n39 VDD1.n38 104.615
R2301 VDD1.n38 VDD1.n32 104.615
R2302 VDD1.n138 VDD1.n132 104.615
R2303 VDD1.n139 VDD1.n138 104.615
R2304 VDD1.n139 VDD1.n128 104.615
R2305 VDD1.n146 VDD1.n128 104.615
R2306 VDD1.n147 VDD1.n146 104.615
R2307 VDD1.n147 VDD1.n124 104.615
R2308 VDD1.n154 VDD1.n124 104.615
R2309 VDD1.n155 VDD1.n154 104.615
R2310 VDD1.n155 VDD1.n120 104.615
R2311 VDD1.n162 VDD1.n120 104.615
R2312 VDD1.n163 VDD1.n162 104.615
R2313 VDD1.n163 VDD1.n116 104.615
R2314 VDD1.n170 VDD1.n116 104.615
R2315 VDD1.n171 VDD1.n170 104.615
R2316 VDD1.n171 VDD1.n112 104.615
R2317 VDD1.n179 VDD1.n112 104.615
R2318 VDD1.n180 VDD1.n179 104.615
R2319 VDD1.n181 VDD1.n180 104.615
R2320 VDD1.n181 VDD1.n108 104.615
R2321 VDD1.n188 VDD1.n108 104.615
R2322 VDD1.n189 VDD1.n188 104.615
R2323 VDD1.n189 VDD1.n104 104.615
R2324 VDD1.n196 VDD1.n104 104.615
R2325 VDD1.n197 VDD1.n196 104.615
R2326 VDD1 VDD1.n201 88.0358
R2327 VDD1.t0 VDD1.n32 52.3082
R2328 VDD1.t1 VDD1.n132 52.3082
R2329 VDD1 VDD1.n100 46.9528
R2330 VDD1.n34 VDD1.n33 15.6677
R2331 VDD1.n134 VDD1.n133 15.6677
R2332 VDD1.n81 VDD1.n10 13.1884
R2333 VDD1.n182 VDD1.n111 13.1884
R2334 VDD1.n82 VDD1.n8 12.8005
R2335 VDD1.n77 VDD1.n12 12.8005
R2336 VDD1.n37 VDD1.n36 12.8005
R2337 VDD1.n137 VDD1.n136 12.8005
R2338 VDD1.n178 VDD1.n177 12.8005
R2339 VDD1.n183 VDD1.n109 12.8005
R2340 VDD1.n86 VDD1.n85 12.0247
R2341 VDD1.n76 VDD1.n13 12.0247
R2342 VDD1.n40 VDD1.n31 12.0247
R2343 VDD1.n140 VDD1.n131 12.0247
R2344 VDD1.n176 VDD1.n113 12.0247
R2345 VDD1.n187 VDD1.n186 12.0247
R2346 VDD1.n89 VDD1.n6 11.249
R2347 VDD1.n73 VDD1.n72 11.249
R2348 VDD1.n41 VDD1.n29 11.249
R2349 VDD1.n141 VDD1.n129 11.249
R2350 VDD1.n173 VDD1.n172 11.249
R2351 VDD1.n190 VDD1.n107 11.249
R2352 VDD1.n90 VDD1.n4 10.4732
R2353 VDD1.n69 VDD1.n15 10.4732
R2354 VDD1.n45 VDD1.n44 10.4732
R2355 VDD1.n145 VDD1.n144 10.4732
R2356 VDD1.n169 VDD1.n115 10.4732
R2357 VDD1.n191 VDD1.n105 10.4732
R2358 VDD1.n94 VDD1.n93 9.69747
R2359 VDD1.n68 VDD1.n17 9.69747
R2360 VDD1.n48 VDD1.n27 9.69747
R2361 VDD1.n148 VDD1.n127 9.69747
R2362 VDD1.n168 VDD1.n117 9.69747
R2363 VDD1.n195 VDD1.n194 9.69747
R2364 VDD1.n100 VDD1.n99 9.45567
R2365 VDD1.n201 VDD1.n200 9.45567
R2366 VDD1.n60 VDD1.n59 9.3005
R2367 VDD1.n19 VDD1.n18 9.3005
R2368 VDD1.n66 VDD1.n65 9.3005
R2369 VDD1.n68 VDD1.n67 9.3005
R2370 VDD1.n15 VDD1.n14 9.3005
R2371 VDD1.n74 VDD1.n73 9.3005
R2372 VDD1.n76 VDD1.n75 9.3005
R2373 VDD1.n12 VDD1.n9 9.3005
R2374 VDD1.n99 VDD1.n98 9.3005
R2375 VDD1.n2 VDD1.n1 9.3005
R2376 VDD1.n93 VDD1.n92 9.3005
R2377 VDD1.n91 VDD1.n90 9.3005
R2378 VDD1.n6 VDD1.n5 9.3005
R2379 VDD1.n85 VDD1.n84 9.3005
R2380 VDD1.n83 VDD1.n82 9.3005
R2381 VDD1.n58 VDD1.n57 9.3005
R2382 VDD1.n23 VDD1.n22 9.3005
R2383 VDD1.n52 VDD1.n51 9.3005
R2384 VDD1.n50 VDD1.n49 9.3005
R2385 VDD1.n27 VDD1.n26 9.3005
R2386 VDD1.n44 VDD1.n43 9.3005
R2387 VDD1.n42 VDD1.n41 9.3005
R2388 VDD1.n31 VDD1.n30 9.3005
R2389 VDD1.n36 VDD1.n35 9.3005
R2390 VDD1.n200 VDD1.n199 9.3005
R2391 VDD1.n103 VDD1.n102 9.3005
R2392 VDD1.n194 VDD1.n193 9.3005
R2393 VDD1.n192 VDD1.n191 9.3005
R2394 VDD1.n107 VDD1.n106 9.3005
R2395 VDD1.n186 VDD1.n185 9.3005
R2396 VDD1.n184 VDD1.n183 9.3005
R2397 VDD1.n123 VDD1.n122 9.3005
R2398 VDD1.n152 VDD1.n151 9.3005
R2399 VDD1.n150 VDD1.n149 9.3005
R2400 VDD1.n127 VDD1.n126 9.3005
R2401 VDD1.n144 VDD1.n143 9.3005
R2402 VDD1.n142 VDD1.n141 9.3005
R2403 VDD1.n131 VDD1.n130 9.3005
R2404 VDD1.n136 VDD1.n135 9.3005
R2405 VDD1.n158 VDD1.n157 9.3005
R2406 VDD1.n160 VDD1.n159 9.3005
R2407 VDD1.n119 VDD1.n118 9.3005
R2408 VDD1.n166 VDD1.n165 9.3005
R2409 VDD1.n168 VDD1.n167 9.3005
R2410 VDD1.n115 VDD1.n114 9.3005
R2411 VDD1.n174 VDD1.n173 9.3005
R2412 VDD1.n176 VDD1.n175 9.3005
R2413 VDD1.n177 VDD1.n110 9.3005
R2414 VDD1.n97 VDD1.n2 8.92171
R2415 VDD1.n65 VDD1.n64 8.92171
R2416 VDD1.n49 VDD1.n25 8.92171
R2417 VDD1.n149 VDD1.n125 8.92171
R2418 VDD1.n165 VDD1.n164 8.92171
R2419 VDD1.n198 VDD1.n103 8.92171
R2420 VDD1.n98 VDD1.n0 8.14595
R2421 VDD1.n61 VDD1.n19 8.14595
R2422 VDD1.n53 VDD1.n52 8.14595
R2423 VDD1.n153 VDD1.n152 8.14595
R2424 VDD1.n161 VDD1.n119 8.14595
R2425 VDD1.n199 VDD1.n101 8.14595
R2426 VDD1.n60 VDD1.n21 7.3702
R2427 VDD1.n56 VDD1.n23 7.3702
R2428 VDD1.n156 VDD1.n123 7.3702
R2429 VDD1.n160 VDD1.n121 7.3702
R2430 VDD1.n57 VDD1.n21 6.59444
R2431 VDD1.n57 VDD1.n56 6.59444
R2432 VDD1.n157 VDD1.n156 6.59444
R2433 VDD1.n157 VDD1.n121 6.59444
R2434 VDD1.n100 VDD1.n0 5.81868
R2435 VDD1.n61 VDD1.n60 5.81868
R2436 VDD1.n53 VDD1.n23 5.81868
R2437 VDD1.n153 VDD1.n123 5.81868
R2438 VDD1.n161 VDD1.n160 5.81868
R2439 VDD1.n201 VDD1.n101 5.81868
R2440 VDD1.n98 VDD1.n97 5.04292
R2441 VDD1.n64 VDD1.n19 5.04292
R2442 VDD1.n52 VDD1.n25 5.04292
R2443 VDD1.n152 VDD1.n125 5.04292
R2444 VDD1.n164 VDD1.n119 5.04292
R2445 VDD1.n199 VDD1.n198 5.04292
R2446 VDD1.n35 VDD1.n34 4.38563
R2447 VDD1.n135 VDD1.n134 4.38563
R2448 VDD1.n94 VDD1.n2 4.26717
R2449 VDD1.n65 VDD1.n17 4.26717
R2450 VDD1.n49 VDD1.n48 4.26717
R2451 VDD1.n149 VDD1.n148 4.26717
R2452 VDD1.n165 VDD1.n117 4.26717
R2453 VDD1.n195 VDD1.n103 4.26717
R2454 VDD1.n93 VDD1.n4 3.49141
R2455 VDD1.n69 VDD1.n68 3.49141
R2456 VDD1.n45 VDD1.n27 3.49141
R2457 VDD1.n145 VDD1.n127 3.49141
R2458 VDD1.n169 VDD1.n168 3.49141
R2459 VDD1.n194 VDD1.n105 3.49141
R2460 VDD1.n90 VDD1.n89 2.71565
R2461 VDD1.n72 VDD1.n15 2.71565
R2462 VDD1.n44 VDD1.n29 2.71565
R2463 VDD1.n144 VDD1.n129 2.71565
R2464 VDD1.n172 VDD1.n115 2.71565
R2465 VDD1.n191 VDD1.n190 2.71565
R2466 VDD1.n86 VDD1.n6 1.93989
R2467 VDD1.n73 VDD1.n13 1.93989
R2468 VDD1.n41 VDD1.n40 1.93989
R2469 VDD1.n141 VDD1.n140 1.93989
R2470 VDD1.n173 VDD1.n113 1.93989
R2471 VDD1.n187 VDD1.n107 1.93989
R2472 VDD1.n85 VDD1.n8 1.16414
R2473 VDD1.n77 VDD1.n76 1.16414
R2474 VDD1.n37 VDD1.n31 1.16414
R2475 VDD1.n137 VDD1.n131 1.16414
R2476 VDD1.n178 VDD1.n176 1.16414
R2477 VDD1.n186 VDD1.n109 1.16414
R2478 VDD1.n82 VDD1.n81 0.388379
R2479 VDD1.n12 VDD1.n10 0.388379
R2480 VDD1.n36 VDD1.n33 0.388379
R2481 VDD1.n136 VDD1.n133 0.388379
R2482 VDD1.n177 VDD1.n111 0.388379
R2483 VDD1.n183 VDD1.n182 0.388379
R2484 VDD1.n99 VDD1.n1 0.155672
R2485 VDD1.n92 VDD1.n1 0.155672
R2486 VDD1.n92 VDD1.n91 0.155672
R2487 VDD1.n91 VDD1.n5 0.155672
R2488 VDD1.n84 VDD1.n5 0.155672
R2489 VDD1.n84 VDD1.n83 0.155672
R2490 VDD1.n83 VDD1.n9 0.155672
R2491 VDD1.n75 VDD1.n9 0.155672
R2492 VDD1.n75 VDD1.n74 0.155672
R2493 VDD1.n74 VDD1.n14 0.155672
R2494 VDD1.n67 VDD1.n14 0.155672
R2495 VDD1.n67 VDD1.n66 0.155672
R2496 VDD1.n66 VDD1.n18 0.155672
R2497 VDD1.n59 VDD1.n18 0.155672
R2498 VDD1.n59 VDD1.n58 0.155672
R2499 VDD1.n58 VDD1.n22 0.155672
R2500 VDD1.n51 VDD1.n22 0.155672
R2501 VDD1.n51 VDD1.n50 0.155672
R2502 VDD1.n50 VDD1.n26 0.155672
R2503 VDD1.n43 VDD1.n26 0.155672
R2504 VDD1.n43 VDD1.n42 0.155672
R2505 VDD1.n42 VDD1.n30 0.155672
R2506 VDD1.n35 VDD1.n30 0.155672
R2507 VDD1.n135 VDD1.n130 0.155672
R2508 VDD1.n142 VDD1.n130 0.155672
R2509 VDD1.n143 VDD1.n142 0.155672
R2510 VDD1.n143 VDD1.n126 0.155672
R2511 VDD1.n150 VDD1.n126 0.155672
R2512 VDD1.n151 VDD1.n150 0.155672
R2513 VDD1.n151 VDD1.n122 0.155672
R2514 VDD1.n158 VDD1.n122 0.155672
R2515 VDD1.n159 VDD1.n158 0.155672
R2516 VDD1.n159 VDD1.n118 0.155672
R2517 VDD1.n166 VDD1.n118 0.155672
R2518 VDD1.n167 VDD1.n166 0.155672
R2519 VDD1.n167 VDD1.n114 0.155672
R2520 VDD1.n174 VDD1.n114 0.155672
R2521 VDD1.n175 VDD1.n174 0.155672
R2522 VDD1.n175 VDD1.n110 0.155672
R2523 VDD1.n184 VDD1.n110 0.155672
R2524 VDD1.n185 VDD1.n184 0.155672
R2525 VDD1.n185 VDD1.n106 0.155672
R2526 VDD1.n192 VDD1.n106 0.155672
R2527 VDD1.n193 VDD1.n192 0.155672
R2528 VDD1.n193 VDD1.n102 0.155672
R2529 VDD1.n200 VDD1.n102 0.155672
C0 VDD2 VN 2.38288f
C1 VDD1 VTAIL 8.99365f
C2 VDD2 VTAIL 9.020451f
C3 VDD1 VDD2 0.439602f
C4 VP VN 5.57477f
C5 VP VTAIL 1.55597f
C6 VN VTAIL 1.54096f
C7 VDD1 VP 2.47204f
C8 VDD1 VN 0.148466f
C9 VDD2 VP 0.244848f
C10 VDD2 B 4.759857f
C11 VDD1 B 7.80527f
C12 VTAIL B 7.880941f
C13 VN B 9.650929f
C14 VP B 4.120632f
C15 VDD1.n0 B 0.029491f
C16 VDD1.n1 B 0.02215f
C17 VDD1.n2 B 0.011903f
C18 VDD1.n3 B 0.028134f
C19 VDD1.n4 B 0.012603f
C20 VDD1.n5 B 0.02215f
C21 VDD1.n6 B 0.011903f
C22 VDD1.n7 B 0.028134f
C23 VDD1.n8 B 0.012603f
C24 VDD1.n9 B 0.02215f
C25 VDD1.n10 B 0.012253f
C26 VDD1.n11 B 0.028134f
C27 VDD1.n12 B 0.011903f
C28 VDD1.n13 B 0.012603f
C29 VDD1.n14 B 0.02215f
C30 VDD1.n15 B 0.011903f
C31 VDD1.n16 B 0.028134f
C32 VDD1.n17 B 0.012603f
C33 VDD1.n18 B 0.02215f
C34 VDD1.n19 B 0.011903f
C35 VDD1.n20 B 0.028134f
C36 VDD1.n21 B 0.012603f
C37 VDD1.n22 B 0.02215f
C38 VDD1.n23 B 0.011903f
C39 VDD1.n24 B 0.028134f
C40 VDD1.n25 B 0.012603f
C41 VDD1.n26 B 0.02215f
C42 VDD1.n27 B 0.011903f
C43 VDD1.n28 B 0.028134f
C44 VDD1.n29 B 0.012603f
C45 VDD1.n30 B 0.02215f
C46 VDD1.n31 B 0.011903f
C47 VDD1.n32 B 0.0211f
C48 VDD1.n33 B 0.016619f
C49 VDD1.t0 B 0.046627f
C50 VDD1.n34 B 0.161853f
C51 VDD1.n35 B 1.75889f
C52 VDD1.n36 B 0.011903f
C53 VDD1.n37 B 0.012603f
C54 VDD1.n38 B 0.028134f
C55 VDD1.n39 B 0.028134f
C56 VDD1.n40 B 0.012603f
C57 VDD1.n41 B 0.011903f
C58 VDD1.n42 B 0.02215f
C59 VDD1.n43 B 0.02215f
C60 VDD1.n44 B 0.011903f
C61 VDD1.n45 B 0.012603f
C62 VDD1.n46 B 0.028134f
C63 VDD1.n47 B 0.028134f
C64 VDD1.n48 B 0.012603f
C65 VDD1.n49 B 0.011903f
C66 VDD1.n50 B 0.02215f
C67 VDD1.n51 B 0.02215f
C68 VDD1.n52 B 0.011903f
C69 VDD1.n53 B 0.012603f
C70 VDD1.n54 B 0.028134f
C71 VDD1.n55 B 0.028134f
C72 VDD1.n56 B 0.012603f
C73 VDD1.n57 B 0.011903f
C74 VDD1.n58 B 0.02215f
C75 VDD1.n59 B 0.02215f
C76 VDD1.n60 B 0.011903f
C77 VDD1.n61 B 0.012603f
C78 VDD1.n62 B 0.028134f
C79 VDD1.n63 B 0.028134f
C80 VDD1.n64 B 0.012603f
C81 VDD1.n65 B 0.011903f
C82 VDD1.n66 B 0.02215f
C83 VDD1.n67 B 0.02215f
C84 VDD1.n68 B 0.011903f
C85 VDD1.n69 B 0.012603f
C86 VDD1.n70 B 0.028134f
C87 VDD1.n71 B 0.028134f
C88 VDD1.n72 B 0.012603f
C89 VDD1.n73 B 0.011903f
C90 VDD1.n74 B 0.02215f
C91 VDD1.n75 B 0.02215f
C92 VDD1.n76 B 0.011903f
C93 VDD1.n77 B 0.012603f
C94 VDD1.n78 B 0.028134f
C95 VDD1.n79 B 0.028134f
C96 VDD1.n80 B 0.028134f
C97 VDD1.n81 B 0.012253f
C98 VDD1.n82 B 0.011903f
C99 VDD1.n83 B 0.02215f
C100 VDD1.n84 B 0.02215f
C101 VDD1.n85 B 0.011903f
C102 VDD1.n86 B 0.012603f
C103 VDD1.n87 B 0.028134f
C104 VDD1.n88 B 0.028134f
C105 VDD1.n89 B 0.012603f
C106 VDD1.n90 B 0.011903f
C107 VDD1.n91 B 0.02215f
C108 VDD1.n92 B 0.02215f
C109 VDD1.n93 B 0.011903f
C110 VDD1.n94 B 0.012603f
C111 VDD1.n95 B 0.028134f
C112 VDD1.n96 B 0.057998f
C113 VDD1.n97 B 0.012603f
C114 VDD1.n98 B 0.011903f
C115 VDD1.n99 B 0.047871f
C116 VDD1.n100 B 0.047638f
C117 VDD1.n101 B 0.029491f
C118 VDD1.n102 B 0.02215f
C119 VDD1.n103 B 0.011903f
C120 VDD1.n104 B 0.028134f
C121 VDD1.n105 B 0.012603f
C122 VDD1.n106 B 0.02215f
C123 VDD1.n107 B 0.011903f
C124 VDD1.n108 B 0.028134f
C125 VDD1.n109 B 0.012603f
C126 VDD1.n110 B 0.02215f
C127 VDD1.n111 B 0.012253f
C128 VDD1.n112 B 0.028134f
C129 VDD1.n113 B 0.012603f
C130 VDD1.n114 B 0.02215f
C131 VDD1.n115 B 0.011903f
C132 VDD1.n116 B 0.028134f
C133 VDD1.n117 B 0.012603f
C134 VDD1.n118 B 0.02215f
C135 VDD1.n119 B 0.011903f
C136 VDD1.n120 B 0.028134f
C137 VDD1.n121 B 0.012603f
C138 VDD1.n122 B 0.02215f
C139 VDD1.n123 B 0.011903f
C140 VDD1.n124 B 0.028134f
C141 VDD1.n125 B 0.012603f
C142 VDD1.n126 B 0.02215f
C143 VDD1.n127 B 0.011903f
C144 VDD1.n128 B 0.028134f
C145 VDD1.n129 B 0.012603f
C146 VDD1.n130 B 0.02215f
C147 VDD1.n131 B 0.011903f
C148 VDD1.n132 B 0.0211f
C149 VDD1.n133 B 0.016619f
C150 VDD1.t1 B 0.046627f
C151 VDD1.n134 B 0.161853f
C152 VDD1.n135 B 1.75889f
C153 VDD1.n136 B 0.011903f
C154 VDD1.n137 B 0.012603f
C155 VDD1.n138 B 0.028134f
C156 VDD1.n139 B 0.028134f
C157 VDD1.n140 B 0.012603f
C158 VDD1.n141 B 0.011903f
C159 VDD1.n142 B 0.02215f
C160 VDD1.n143 B 0.02215f
C161 VDD1.n144 B 0.011903f
C162 VDD1.n145 B 0.012603f
C163 VDD1.n146 B 0.028134f
C164 VDD1.n147 B 0.028134f
C165 VDD1.n148 B 0.012603f
C166 VDD1.n149 B 0.011903f
C167 VDD1.n150 B 0.02215f
C168 VDD1.n151 B 0.02215f
C169 VDD1.n152 B 0.011903f
C170 VDD1.n153 B 0.012603f
C171 VDD1.n154 B 0.028134f
C172 VDD1.n155 B 0.028134f
C173 VDD1.n156 B 0.012603f
C174 VDD1.n157 B 0.011903f
C175 VDD1.n158 B 0.02215f
C176 VDD1.n159 B 0.02215f
C177 VDD1.n160 B 0.011903f
C178 VDD1.n161 B 0.012603f
C179 VDD1.n162 B 0.028134f
C180 VDD1.n163 B 0.028134f
C181 VDD1.n164 B 0.012603f
C182 VDD1.n165 B 0.011903f
C183 VDD1.n166 B 0.02215f
C184 VDD1.n167 B 0.02215f
C185 VDD1.n168 B 0.011903f
C186 VDD1.n169 B 0.012603f
C187 VDD1.n170 B 0.028134f
C188 VDD1.n171 B 0.028134f
C189 VDD1.n172 B 0.012603f
C190 VDD1.n173 B 0.011903f
C191 VDD1.n174 B 0.02215f
C192 VDD1.n175 B 0.02215f
C193 VDD1.n176 B 0.011903f
C194 VDD1.n177 B 0.011903f
C195 VDD1.n178 B 0.012603f
C196 VDD1.n179 B 0.028134f
C197 VDD1.n180 B 0.028134f
C198 VDD1.n181 B 0.028134f
C199 VDD1.n182 B 0.012253f
C200 VDD1.n183 B 0.011903f
C201 VDD1.n184 B 0.02215f
C202 VDD1.n185 B 0.02215f
C203 VDD1.n186 B 0.011903f
C204 VDD1.n187 B 0.012603f
C205 VDD1.n188 B 0.028134f
C206 VDD1.n189 B 0.028134f
C207 VDD1.n190 B 0.012603f
C208 VDD1.n191 B 0.011903f
C209 VDD1.n192 B 0.02215f
C210 VDD1.n193 B 0.02215f
C211 VDD1.n194 B 0.011903f
C212 VDD1.n195 B 0.012603f
C213 VDD1.n196 B 0.028134f
C214 VDD1.n197 B 0.057998f
C215 VDD1.n198 B 0.012603f
C216 VDD1.n199 B 0.011903f
C217 VDD1.n200 B 0.047871f
C218 VDD1.n201 B 0.765124f
C219 VP.t1 B 1.34978f
C220 VP.t0 B 1.25789f
C221 VP.n0 B 5.48244f
C222 VDD2.n0 B 0.029444f
C223 VDD2.n1 B 0.022115f
C224 VDD2.n2 B 0.011884f
C225 VDD2.n3 B 0.028089f
C226 VDD2.n4 B 0.012583f
C227 VDD2.n5 B 0.022115f
C228 VDD2.n6 B 0.011884f
C229 VDD2.n7 B 0.028089f
C230 VDD2.n8 B 0.012583f
C231 VDD2.n9 B 0.022115f
C232 VDD2.n10 B 0.012233f
C233 VDD2.n11 B 0.028089f
C234 VDD2.n12 B 0.012583f
C235 VDD2.n13 B 0.022115f
C236 VDD2.n14 B 0.011884f
C237 VDD2.n15 B 0.028089f
C238 VDD2.n16 B 0.012583f
C239 VDD2.n17 B 0.022115f
C240 VDD2.n18 B 0.011884f
C241 VDD2.n19 B 0.028089f
C242 VDD2.n20 B 0.012583f
C243 VDD2.n21 B 0.022115f
C244 VDD2.n22 B 0.011884f
C245 VDD2.n23 B 0.028089f
C246 VDD2.n24 B 0.012583f
C247 VDD2.n25 B 0.022115f
C248 VDD2.n26 B 0.011884f
C249 VDD2.n27 B 0.028089f
C250 VDD2.n28 B 0.012583f
C251 VDD2.n29 B 0.022115f
C252 VDD2.n30 B 0.011884f
C253 VDD2.n31 B 0.021067f
C254 VDD2.n32 B 0.016593f
C255 VDD2.t0 B 0.046553f
C256 VDD2.n33 B 0.161595f
C257 VDD2.n34 B 1.75609f
C258 VDD2.n35 B 0.011884f
C259 VDD2.n36 B 0.012583f
C260 VDD2.n37 B 0.028089f
C261 VDD2.n38 B 0.028089f
C262 VDD2.n39 B 0.012583f
C263 VDD2.n40 B 0.011884f
C264 VDD2.n41 B 0.022115f
C265 VDD2.n42 B 0.022115f
C266 VDD2.n43 B 0.011884f
C267 VDD2.n44 B 0.012583f
C268 VDD2.n45 B 0.028089f
C269 VDD2.n46 B 0.028089f
C270 VDD2.n47 B 0.012583f
C271 VDD2.n48 B 0.011884f
C272 VDD2.n49 B 0.022115f
C273 VDD2.n50 B 0.022115f
C274 VDD2.n51 B 0.011884f
C275 VDD2.n52 B 0.012583f
C276 VDD2.n53 B 0.028089f
C277 VDD2.n54 B 0.028089f
C278 VDD2.n55 B 0.012583f
C279 VDD2.n56 B 0.011884f
C280 VDD2.n57 B 0.022115f
C281 VDD2.n58 B 0.022115f
C282 VDD2.n59 B 0.011884f
C283 VDD2.n60 B 0.012583f
C284 VDD2.n61 B 0.028089f
C285 VDD2.n62 B 0.028089f
C286 VDD2.n63 B 0.012583f
C287 VDD2.n64 B 0.011884f
C288 VDD2.n65 B 0.022115f
C289 VDD2.n66 B 0.022115f
C290 VDD2.n67 B 0.011884f
C291 VDD2.n68 B 0.012583f
C292 VDD2.n69 B 0.028089f
C293 VDD2.n70 B 0.028089f
C294 VDD2.n71 B 0.012583f
C295 VDD2.n72 B 0.011884f
C296 VDD2.n73 B 0.022115f
C297 VDD2.n74 B 0.022115f
C298 VDD2.n75 B 0.011884f
C299 VDD2.n76 B 0.011884f
C300 VDD2.n77 B 0.012583f
C301 VDD2.n78 B 0.028089f
C302 VDD2.n79 B 0.028089f
C303 VDD2.n80 B 0.028089f
C304 VDD2.n81 B 0.012233f
C305 VDD2.n82 B 0.011884f
C306 VDD2.n83 B 0.022115f
C307 VDD2.n84 B 0.022115f
C308 VDD2.n85 B 0.011884f
C309 VDD2.n86 B 0.012583f
C310 VDD2.n87 B 0.028089f
C311 VDD2.n88 B 0.028089f
C312 VDD2.n89 B 0.012583f
C313 VDD2.n90 B 0.011884f
C314 VDD2.n91 B 0.022115f
C315 VDD2.n92 B 0.022115f
C316 VDD2.n93 B 0.011884f
C317 VDD2.n94 B 0.012583f
C318 VDD2.n95 B 0.028089f
C319 VDD2.n96 B 0.057905f
C320 VDD2.n97 B 0.012583f
C321 VDD2.n98 B 0.011884f
C322 VDD2.n99 B 0.047795f
C323 VDD2.n100 B 0.733041f
C324 VDD2.n101 B 0.029444f
C325 VDD2.n102 B 0.022115f
C326 VDD2.n103 B 0.011884f
C327 VDD2.n104 B 0.028089f
C328 VDD2.n105 B 0.012583f
C329 VDD2.n106 B 0.022115f
C330 VDD2.n107 B 0.011884f
C331 VDD2.n108 B 0.028089f
C332 VDD2.n109 B 0.012583f
C333 VDD2.n110 B 0.022115f
C334 VDD2.n111 B 0.012233f
C335 VDD2.n112 B 0.028089f
C336 VDD2.n113 B 0.011884f
C337 VDD2.n114 B 0.012583f
C338 VDD2.n115 B 0.022115f
C339 VDD2.n116 B 0.011884f
C340 VDD2.n117 B 0.028089f
C341 VDD2.n118 B 0.012583f
C342 VDD2.n119 B 0.022115f
C343 VDD2.n120 B 0.011884f
C344 VDD2.n121 B 0.028089f
C345 VDD2.n122 B 0.012583f
C346 VDD2.n123 B 0.022115f
C347 VDD2.n124 B 0.011884f
C348 VDD2.n125 B 0.028089f
C349 VDD2.n126 B 0.012583f
C350 VDD2.n127 B 0.022115f
C351 VDD2.n128 B 0.011884f
C352 VDD2.n129 B 0.028089f
C353 VDD2.n130 B 0.012583f
C354 VDD2.n131 B 0.022115f
C355 VDD2.n132 B 0.011884f
C356 VDD2.n133 B 0.021067f
C357 VDD2.n134 B 0.016593f
C358 VDD2.t1 B 0.046553f
C359 VDD2.n135 B 0.161595f
C360 VDD2.n136 B 1.75609f
C361 VDD2.n137 B 0.011884f
C362 VDD2.n138 B 0.012583f
C363 VDD2.n139 B 0.028089f
C364 VDD2.n140 B 0.028089f
C365 VDD2.n141 B 0.012583f
C366 VDD2.n142 B 0.011884f
C367 VDD2.n143 B 0.022115f
C368 VDD2.n144 B 0.022115f
C369 VDD2.n145 B 0.011884f
C370 VDD2.n146 B 0.012583f
C371 VDD2.n147 B 0.028089f
C372 VDD2.n148 B 0.028089f
C373 VDD2.n149 B 0.012583f
C374 VDD2.n150 B 0.011884f
C375 VDD2.n151 B 0.022115f
C376 VDD2.n152 B 0.022115f
C377 VDD2.n153 B 0.011884f
C378 VDD2.n154 B 0.012583f
C379 VDD2.n155 B 0.028089f
C380 VDD2.n156 B 0.028089f
C381 VDD2.n157 B 0.012583f
C382 VDD2.n158 B 0.011884f
C383 VDD2.n159 B 0.022115f
C384 VDD2.n160 B 0.022115f
C385 VDD2.n161 B 0.011884f
C386 VDD2.n162 B 0.012583f
C387 VDD2.n163 B 0.028089f
C388 VDD2.n164 B 0.028089f
C389 VDD2.n165 B 0.012583f
C390 VDD2.n166 B 0.011884f
C391 VDD2.n167 B 0.022115f
C392 VDD2.n168 B 0.022115f
C393 VDD2.n169 B 0.011884f
C394 VDD2.n170 B 0.012583f
C395 VDD2.n171 B 0.028089f
C396 VDD2.n172 B 0.028089f
C397 VDD2.n173 B 0.012583f
C398 VDD2.n174 B 0.011884f
C399 VDD2.n175 B 0.022115f
C400 VDD2.n176 B 0.022115f
C401 VDD2.n177 B 0.011884f
C402 VDD2.n178 B 0.012583f
C403 VDD2.n179 B 0.028089f
C404 VDD2.n180 B 0.028089f
C405 VDD2.n181 B 0.028089f
C406 VDD2.n182 B 0.012233f
C407 VDD2.n183 B 0.011884f
C408 VDD2.n184 B 0.022115f
C409 VDD2.n185 B 0.022115f
C410 VDD2.n186 B 0.011884f
C411 VDD2.n187 B 0.012583f
C412 VDD2.n188 B 0.028089f
C413 VDD2.n189 B 0.028089f
C414 VDD2.n190 B 0.012583f
C415 VDD2.n191 B 0.011884f
C416 VDD2.n192 B 0.022115f
C417 VDD2.n193 B 0.022115f
C418 VDD2.n194 B 0.011884f
C419 VDD2.n195 B 0.012583f
C420 VDD2.n196 B 0.028089f
C421 VDD2.n197 B 0.057905f
C422 VDD2.n198 B 0.012583f
C423 VDD2.n199 B 0.011884f
C424 VDD2.n200 B 0.047795f
C425 VDD2.n201 B 0.047295f
C426 VDD2.n202 B 2.86765f
C427 VTAIL.n0 B 0.024323f
C428 VTAIL.n1 B 0.018269f
C429 VTAIL.n2 B 0.009817f
C430 VTAIL.n3 B 0.023204f
C431 VTAIL.n4 B 0.010394f
C432 VTAIL.n5 B 0.018269f
C433 VTAIL.n6 B 0.009817f
C434 VTAIL.n7 B 0.023204f
C435 VTAIL.n8 B 0.010394f
C436 VTAIL.n9 B 0.018269f
C437 VTAIL.n10 B 0.010106f
C438 VTAIL.n11 B 0.023204f
C439 VTAIL.n12 B 0.010394f
C440 VTAIL.n13 B 0.018269f
C441 VTAIL.n14 B 0.009817f
C442 VTAIL.n15 B 0.023204f
C443 VTAIL.n16 B 0.010394f
C444 VTAIL.n17 B 0.018269f
C445 VTAIL.n18 B 0.009817f
C446 VTAIL.n19 B 0.023204f
C447 VTAIL.n20 B 0.010394f
C448 VTAIL.n21 B 0.018269f
C449 VTAIL.n22 B 0.009817f
C450 VTAIL.n23 B 0.023204f
C451 VTAIL.n24 B 0.010394f
C452 VTAIL.n25 B 0.018269f
C453 VTAIL.n26 B 0.009817f
C454 VTAIL.n27 B 0.023204f
C455 VTAIL.n28 B 0.010394f
C456 VTAIL.n29 B 0.018269f
C457 VTAIL.n30 B 0.009817f
C458 VTAIL.n31 B 0.017403f
C459 VTAIL.n32 B 0.013707f
C460 VTAIL.t1 B 0.038457f
C461 VTAIL.n33 B 0.133492f
C462 VTAIL.n34 B 1.45068f
C463 VTAIL.n35 B 0.009817f
C464 VTAIL.n36 B 0.010394f
C465 VTAIL.n37 B 0.023204f
C466 VTAIL.n38 B 0.023204f
C467 VTAIL.n39 B 0.010394f
C468 VTAIL.n40 B 0.009817f
C469 VTAIL.n41 B 0.018269f
C470 VTAIL.n42 B 0.018269f
C471 VTAIL.n43 B 0.009817f
C472 VTAIL.n44 B 0.010394f
C473 VTAIL.n45 B 0.023204f
C474 VTAIL.n46 B 0.023204f
C475 VTAIL.n47 B 0.010394f
C476 VTAIL.n48 B 0.009817f
C477 VTAIL.n49 B 0.018269f
C478 VTAIL.n50 B 0.018269f
C479 VTAIL.n51 B 0.009817f
C480 VTAIL.n52 B 0.010394f
C481 VTAIL.n53 B 0.023204f
C482 VTAIL.n54 B 0.023204f
C483 VTAIL.n55 B 0.010394f
C484 VTAIL.n56 B 0.009817f
C485 VTAIL.n57 B 0.018269f
C486 VTAIL.n58 B 0.018269f
C487 VTAIL.n59 B 0.009817f
C488 VTAIL.n60 B 0.010394f
C489 VTAIL.n61 B 0.023204f
C490 VTAIL.n62 B 0.023204f
C491 VTAIL.n63 B 0.010394f
C492 VTAIL.n64 B 0.009817f
C493 VTAIL.n65 B 0.018269f
C494 VTAIL.n66 B 0.018269f
C495 VTAIL.n67 B 0.009817f
C496 VTAIL.n68 B 0.010394f
C497 VTAIL.n69 B 0.023204f
C498 VTAIL.n70 B 0.023204f
C499 VTAIL.n71 B 0.010394f
C500 VTAIL.n72 B 0.009817f
C501 VTAIL.n73 B 0.018269f
C502 VTAIL.n74 B 0.018269f
C503 VTAIL.n75 B 0.009817f
C504 VTAIL.n76 B 0.009817f
C505 VTAIL.n77 B 0.010394f
C506 VTAIL.n78 B 0.023204f
C507 VTAIL.n79 B 0.023204f
C508 VTAIL.n80 B 0.023204f
C509 VTAIL.n81 B 0.010106f
C510 VTAIL.n82 B 0.009817f
C511 VTAIL.n83 B 0.018269f
C512 VTAIL.n84 B 0.018269f
C513 VTAIL.n85 B 0.009817f
C514 VTAIL.n86 B 0.010394f
C515 VTAIL.n87 B 0.023204f
C516 VTAIL.n88 B 0.023204f
C517 VTAIL.n89 B 0.010394f
C518 VTAIL.n90 B 0.009817f
C519 VTAIL.n91 B 0.018269f
C520 VTAIL.n92 B 0.018269f
C521 VTAIL.n93 B 0.009817f
C522 VTAIL.n94 B 0.010394f
C523 VTAIL.n95 B 0.023204f
C524 VTAIL.n96 B 0.047835f
C525 VTAIL.n97 B 0.010394f
C526 VTAIL.n98 B 0.009817f
C527 VTAIL.n99 B 0.039483f
C528 VTAIL.n100 B 0.026432f
C529 VTAIL.n101 B 1.30115f
C530 VTAIL.n102 B 0.024323f
C531 VTAIL.n103 B 0.018269f
C532 VTAIL.n104 B 0.009817f
C533 VTAIL.n105 B 0.023204f
C534 VTAIL.n106 B 0.010394f
C535 VTAIL.n107 B 0.018269f
C536 VTAIL.n108 B 0.009817f
C537 VTAIL.n109 B 0.023204f
C538 VTAIL.n110 B 0.010394f
C539 VTAIL.n111 B 0.018269f
C540 VTAIL.n112 B 0.010106f
C541 VTAIL.n113 B 0.023204f
C542 VTAIL.n114 B 0.009817f
C543 VTAIL.n115 B 0.010394f
C544 VTAIL.n116 B 0.018269f
C545 VTAIL.n117 B 0.009817f
C546 VTAIL.n118 B 0.023204f
C547 VTAIL.n119 B 0.010394f
C548 VTAIL.n120 B 0.018269f
C549 VTAIL.n121 B 0.009817f
C550 VTAIL.n122 B 0.023204f
C551 VTAIL.n123 B 0.010394f
C552 VTAIL.n124 B 0.018269f
C553 VTAIL.n125 B 0.009817f
C554 VTAIL.n126 B 0.023204f
C555 VTAIL.n127 B 0.010394f
C556 VTAIL.n128 B 0.018269f
C557 VTAIL.n129 B 0.009817f
C558 VTAIL.n130 B 0.023204f
C559 VTAIL.n131 B 0.010394f
C560 VTAIL.n132 B 0.018269f
C561 VTAIL.n133 B 0.009817f
C562 VTAIL.n134 B 0.017403f
C563 VTAIL.n135 B 0.013707f
C564 VTAIL.t2 B 0.038457f
C565 VTAIL.n136 B 0.133492f
C566 VTAIL.n137 B 1.45068f
C567 VTAIL.n138 B 0.009817f
C568 VTAIL.n139 B 0.010394f
C569 VTAIL.n140 B 0.023204f
C570 VTAIL.n141 B 0.023204f
C571 VTAIL.n142 B 0.010394f
C572 VTAIL.n143 B 0.009817f
C573 VTAIL.n144 B 0.018269f
C574 VTAIL.n145 B 0.018269f
C575 VTAIL.n146 B 0.009817f
C576 VTAIL.n147 B 0.010394f
C577 VTAIL.n148 B 0.023204f
C578 VTAIL.n149 B 0.023204f
C579 VTAIL.n150 B 0.010394f
C580 VTAIL.n151 B 0.009817f
C581 VTAIL.n152 B 0.018269f
C582 VTAIL.n153 B 0.018269f
C583 VTAIL.n154 B 0.009817f
C584 VTAIL.n155 B 0.010394f
C585 VTAIL.n156 B 0.023204f
C586 VTAIL.n157 B 0.023204f
C587 VTAIL.n158 B 0.010394f
C588 VTAIL.n159 B 0.009817f
C589 VTAIL.n160 B 0.018269f
C590 VTAIL.n161 B 0.018269f
C591 VTAIL.n162 B 0.009817f
C592 VTAIL.n163 B 0.010394f
C593 VTAIL.n164 B 0.023204f
C594 VTAIL.n165 B 0.023204f
C595 VTAIL.n166 B 0.010394f
C596 VTAIL.n167 B 0.009817f
C597 VTAIL.n168 B 0.018269f
C598 VTAIL.n169 B 0.018269f
C599 VTAIL.n170 B 0.009817f
C600 VTAIL.n171 B 0.010394f
C601 VTAIL.n172 B 0.023204f
C602 VTAIL.n173 B 0.023204f
C603 VTAIL.n174 B 0.010394f
C604 VTAIL.n175 B 0.009817f
C605 VTAIL.n176 B 0.018269f
C606 VTAIL.n177 B 0.018269f
C607 VTAIL.n178 B 0.009817f
C608 VTAIL.n179 B 0.010394f
C609 VTAIL.n180 B 0.023204f
C610 VTAIL.n181 B 0.023204f
C611 VTAIL.n182 B 0.023204f
C612 VTAIL.n183 B 0.010106f
C613 VTAIL.n184 B 0.009817f
C614 VTAIL.n185 B 0.018269f
C615 VTAIL.n186 B 0.018269f
C616 VTAIL.n187 B 0.009817f
C617 VTAIL.n188 B 0.010394f
C618 VTAIL.n189 B 0.023204f
C619 VTAIL.n190 B 0.023204f
C620 VTAIL.n191 B 0.010394f
C621 VTAIL.n192 B 0.009817f
C622 VTAIL.n193 B 0.018269f
C623 VTAIL.n194 B 0.018269f
C624 VTAIL.n195 B 0.009817f
C625 VTAIL.n196 B 0.010394f
C626 VTAIL.n197 B 0.023204f
C627 VTAIL.n198 B 0.047835f
C628 VTAIL.n199 B 0.010394f
C629 VTAIL.n200 B 0.009817f
C630 VTAIL.n201 B 0.039483f
C631 VTAIL.n202 B 0.026432f
C632 VTAIL.n203 B 1.30737f
C633 VTAIL.n204 B 0.024323f
C634 VTAIL.n205 B 0.018269f
C635 VTAIL.n206 B 0.009817f
C636 VTAIL.n207 B 0.023204f
C637 VTAIL.n208 B 0.010394f
C638 VTAIL.n209 B 0.018269f
C639 VTAIL.n210 B 0.009817f
C640 VTAIL.n211 B 0.023204f
C641 VTAIL.n212 B 0.010394f
C642 VTAIL.n213 B 0.018269f
C643 VTAIL.n214 B 0.010106f
C644 VTAIL.n215 B 0.023204f
C645 VTAIL.n216 B 0.009817f
C646 VTAIL.n217 B 0.010394f
C647 VTAIL.n218 B 0.018269f
C648 VTAIL.n219 B 0.009817f
C649 VTAIL.n220 B 0.023204f
C650 VTAIL.n221 B 0.010394f
C651 VTAIL.n222 B 0.018269f
C652 VTAIL.n223 B 0.009817f
C653 VTAIL.n224 B 0.023204f
C654 VTAIL.n225 B 0.010394f
C655 VTAIL.n226 B 0.018269f
C656 VTAIL.n227 B 0.009817f
C657 VTAIL.n228 B 0.023204f
C658 VTAIL.n229 B 0.010394f
C659 VTAIL.n230 B 0.018269f
C660 VTAIL.n231 B 0.009817f
C661 VTAIL.n232 B 0.023204f
C662 VTAIL.n233 B 0.010394f
C663 VTAIL.n234 B 0.018269f
C664 VTAIL.n235 B 0.009817f
C665 VTAIL.n236 B 0.017403f
C666 VTAIL.n237 B 0.013707f
C667 VTAIL.t0 B 0.038457f
C668 VTAIL.n238 B 0.133492f
C669 VTAIL.n239 B 1.45068f
C670 VTAIL.n240 B 0.009817f
C671 VTAIL.n241 B 0.010394f
C672 VTAIL.n242 B 0.023204f
C673 VTAIL.n243 B 0.023204f
C674 VTAIL.n244 B 0.010394f
C675 VTAIL.n245 B 0.009817f
C676 VTAIL.n246 B 0.018269f
C677 VTAIL.n247 B 0.018269f
C678 VTAIL.n248 B 0.009817f
C679 VTAIL.n249 B 0.010394f
C680 VTAIL.n250 B 0.023204f
C681 VTAIL.n251 B 0.023204f
C682 VTAIL.n252 B 0.010394f
C683 VTAIL.n253 B 0.009817f
C684 VTAIL.n254 B 0.018269f
C685 VTAIL.n255 B 0.018269f
C686 VTAIL.n256 B 0.009817f
C687 VTAIL.n257 B 0.010394f
C688 VTAIL.n258 B 0.023204f
C689 VTAIL.n259 B 0.023204f
C690 VTAIL.n260 B 0.010394f
C691 VTAIL.n261 B 0.009817f
C692 VTAIL.n262 B 0.018269f
C693 VTAIL.n263 B 0.018269f
C694 VTAIL.n264 B 0.009817f
C695 VTAIL.n265 B 0.010394f
C696 VTAIL.n266 B 0.023204f
C697 VTAIL.n267 B 0.023204f
C698 VTAIL.n268 B 0.010394f
C699 VTAIL.n269 B 0.009817f
C700 VTAIL.n270 B 0.018269f
C701 VTAIL.n271 B 0.018269f
C702 VTAIL.n272 B 0.009817f
C703 VTAIL.n273 B 0.010394f
C704 VTAIL.n274 B 0.023204f
C705 VTAIL.n275 B 0.023204f
C706 VTAIL.n276 B 0.010394f
C707 VTAIL.n277 B 0.009817f
C708 VTAIL.n278 B 0.018269f
C709 VTAIL.n279 B 0.018269f
C710 VTAIL.n280 B 0.009817f
C711 VTAIL.n281 B 0.010394f
C712 VTAIL.n282 B 0.023204f
C713 VTAIL.n283 B 0.023204f
C714 VTAIL.n284 B 0.023204f
C715 VTAIL.n285 B 0.010106f
C716 VTAIL.n286 B 0.009817f
C717 VTAIL.n287 B 0.018269f
C718 VTAIL.n288 B 0.018269f
C719 VTAIL.n289 B 0.009817f
C720 VTAIL.n290 B 0.010394f
C721 VTAIL.n291 B 0.023204f
C722 VTAIL.n292 B 0.023204f
C723 VTAIL.n293 B 0.010394f
C724 VTAIL.n294 B 0.009817f
C725 VTAIL.n295 B 0.018269f
C726 VTAIL.n296 B 0.018269f
C727 VTAIL.n297 B 0.009817f
C728 VTAIL.n298 B 0.010394f
C729 VTAIL.n299 B 0.023204f
C730 VTAIL.n300 B 0.047835f
C731 VTAIL.n301 B 0.010394f
C732 VTAIL.n302 B 0.009817f
C733 VTAIL.n303 B 0.039483f
C734 VTAIL.n304 B 0.026432f
C735 VTAIL.n305 B 1.2688f
C736 VTAIL.n306 B 0.024323f
C737 VTAIL.n307 B 0.018269f
C738 VTAIL.n308 B 0.009817f
C739 VTAIL.n309 B 0.023204f
C740 VTAIL.n310 B 0.010394f
C741 VTAIL.n311 B 0.018269f
C742 VTAIL.n312 B 0.009817f
C743 VTAIL.n313 B 0.023204f
C744 VTAIL.n314 B 0.010394f
C745 VTAIL.n315 B 0.018269f
C746 VTAIL.n316 B 0.010106f
C747 VTAIL.n317 B 0.023204f
C748 VTAIL.n318 B 0.010394f
C749 VTAIL.n319 B 0.018269f
C750 VTAIL.n320 B 0.009817f
C751 VTAIL.n321 B 0.023204f
C752 VTAIL.n322 B 0.010394f
C753 VTAIL.n323 B 0.018269f
C754 VTAIL.n324 B 0.009817f
C755 VTAIL.n325 B 0.023204f
C756 VTAIL.n326 B 0.010394f
C757 VTAIL.n327 B 0.018269f
C758 VTAIL.n328 B 0.009817f
C759 VTAIL.n329 B 0.023204f
C760 VTAIL.n330 B 0.010394f
C761 VTAIL.n331 B 0.018269f
C762 VTAIL.n332 B 0.009817f
C763 VTAIL.n333 B 0.023204f
C764 VTAIL.n334 B 0.010394f
C765 VTAIL.n335 B 0.018269f
C766 VTAIL.n336 B 0.009817f
C767 VTAIL.n337 B 0.017403f
C768 VTAIL.n338 B 0.013707f
C769 VTAIL.t3 B 0.038457f
C770 VTAIL.n339 B 0.133492f
C771 VTAIL.n340 B 1.45068f
C772 VTAIL.n341 B 0.009817f
C773 VTAIL.n342 B 0.010394f
C774 VTAIL.n343 B 0.023204f
C775 VTAIL.n344 B 0.023204f
C776 VTAIL.n345 B 0.010394f
C777 VTAIL.n346 B 0.009817f
C778 VTAIL.n347 B 0.018269f
C779 VTAIL.n348 B 0.018269f
C780 VTAIL.n349 B 0.009817f
C781 VTAIL.n350 B 0.010394f
C782 VTAIL.n351 B 0.023204f
C783 VTAIL.n352 B 0.023204f
C784 VTAIL.n353 B 0.010394f
C785 VTAIL.n354 B 0.009817f
C786 VTAIL.n355 B 0.018269f
C787 VTAIL.n356 B 0.018269f
C788 VTAIL.n357 B 0.009817f
C789 VTAIL.n358 B 0.010394f
C790 VTAIL.n359 B 0.023204f
C791 VTAIL.n360 B 0.023204f
C792 VTAIL.n361 B 0.010394f
C793 VTAIL.n362 B 0.009817f
C794 VTAIL.n363 B 0.018269f
C795 VTAIL.n364 B 0.018269f
C796 VTAIL.n365 B 0.009817f
C797 VTAIL.n366 B 0.010394f
C798 VTAIL.n367 B 0.023204f
C799 VTAIL.n368 B 0.023204f
C800 VTAIL.n369 B 0.010394f
C801 VTAIL.n370 B 0.009817f
C802 VTAIL.n371 B 0.018269f
C803 VTAIL.n372 B 0.018269f
C804 VTAIL.n373 B 0.009817f
C805 VTAIL.n374 B 0.010394f
C806 VTAIL.n375 B 0.023204f
C807 VTAIL.n376 B 0.023204f
C808 VTAIL.n377 B 0.010394f
C809 VTAIL.n378 B 0.009817f
C810 VTAIL.n379 B 0.018269f
C811 VTAIL.n380 B 0.018269f
C812 VTAIL.n381 B 0.009817f
C813 VTAIL.n382 B 0.009817f
C814 VTAIL.n383 B 0.010394f
C815 VTAIL.n384 B 0.023204f
C816 VTAIL.n385 B 0.023204f
C817 VTAIL.n386 B 0.023204f
C818 VTAIL.n387 B 0.010106f
C819 VTAIL.n388 B 0.009817f
C820 VTAIL.n389 B 0.018269f
C821 VTAIL.n390 B 0.018269f
C822 VTAIL.n391 B 0.009817f
C823 VTAIL.n392 B 0.010394f
C824 VTAIL.n393 B 0.023204f
C825 VTAIL.n394 B 0.023204f
C826 VTAIL.n395 B 0.010394f
C827 VTAIL.n396 B 0.009817f
C828 VTAIL.n397 B 0.018269f
C829 VTAIL.n398 B 0.018269f
C830 VTAIL.n399 B 0.009817f
C831 VTAIL.n400 B 0.010394f
C832 VTAIL.n401 B 0.023204f
C833 VTAIL.n402 B 0.047835f
C834 VTAIL.n403 B 0.010394f
C835 VTAIL.n404 B 0.009817f
C836 VTAIL.n405 B 0.039483f
C837 VTAIL.n406 B 0.026432f
C838 VTAIL.n407 B 1.22807f
C839 VN.t1 B 1.23078f
C840 VN.t0 B 1.32259f
.ends

