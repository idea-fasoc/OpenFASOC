* NGSPICE file created from diff_pair_sample_0148.ext - technology: sky130A

.subckt diff_pair_sample_0148 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=2.6832 ps=14.54 w=6.88 l=0.25
X1 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=0 ps=0 w=6.88 l=0.25
X2 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=0 ps=0 w=6.88 l=0.25
X3 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=2.6832 ps=14.54 w=6.88 l=0.25
X4 VDD2.t0 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=2.6832 ps=14.54 w=6.88 l=0.25
X5 VDD1.t0 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=2.6832 ps=14.54 w=6.88 l=0.25
X6 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=0 ps=0 w=6.88 l=0.25
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6832 pd=14.54 as=0 ps=0 w=6.88 l=0.25
R0 VN VN.t0 1008.89
R1 VN VN.t1 974.004
R2 VTAIL.n1 VTAIL.t3 54.3221
R3 VTAIL.n3 VTAIL.t2 54.322
R4 VTAIL.n0 VTAIL.t1 54.322
R5 VTAIL.n2 VTAIL.t0 54.322
R6 VTAIL.n1 VTAIL.n0 19.3152
R7 VTAIL.n3 VTAIL.n2 18.8152
R8 VTAIL.n2 VTAIL.n1 0.720328
R9 VTAIL VTAIL.n0 0.653517
R10 VTAIL VTAIL.n3 0.0673103
R11 VDD2.n0 VDD2.t0 101.609
R12 VDD2.n0 VDD2.t1 71.0008
R13 VDD2 VDD2.n0 0.18369
R14 B.n62 B.t2 887.533
R15 B.n59 B.t6 887.533
R16 B.n243 B.t9 887.533
R17 B.n240 B.t13 887.533
R18 B.n420 B.n419 585
R19 B.n421 B.n420 585
R20 B.n187 B.n58 585
R21 B.n186 B.n185 585
R22 B.n184 B.n183 585
R23 B.n182 B.n181 585
R24 B.n180 B.n179 585
R25 B.n178 B.n177 585
R26 B.n176 B.n175 585
R27 B.n174 B.n173 585
R28 B.n172 B.n171 585
R29 B.n170 B.n169 585
R30 B.n168 B.n167 585
R31 B.n166 B.n165 585
R32 B.n164 B.n163 585
R33 B.n162 B.n161 585
R34 B.n160 B.n159 585
R35 B.n158 B.n157 585
R36 B.n156 B.n155 585
R37 B.n154 B.n153 585
R38 B.n152 B.n151 585
R39 B.n150 B.n149 585
R40 B.n148 B.n147 585
R41 B.n146 B.n145 585
R42 B.n144 B.n143 585
R43 B.n142 B.n141 585
R44 B.n140 B.n139 585
R45 B.n138 B.n137 585
R46 B.n136 B.n135 585
R47 B.n134 B.n133 585
R48 B.n132 B.n131 585
R49 B.n130 B.n129 585
R50 B.n128 B.n127 585
R51 B.n126 B.n125 585
R52 B.n124 B.n123 585
R53 B.n122 B.n121 585
R54 B.n120 B.n119 585
R55 B.n117 B.n116 585
R56 B.n115 B.n114 585
R57 B.n113 B.n112 585
R58 B.n111 B.n110 585
R59 B.n109 B.n108 585
R60 B.n107 B.n106 585
R61 B.n105 B.n104 585
R62 B.n103 B.n102 585
R63 B.n101 B.n100 585
R64 B.n99 B.n98 585
R65 B.n97 B.n96 585
R66 B.n95 B.n94 585
R67 B.n93 B.n92 585
R68 B.n91 B.n90 585
R69 B.n89 B.n88 585
R70 B.n87 B.n86 585
R71 B.n85 B.n84 585
R72 B.n83 B.n82 585
R73 B.n81 B.n80 585
R74 B.n79 B.n78 585
R75 B.n77 B.n76 585
R76 B.n75 B.n74 585
R77 B.n73 B.n72 585
R78 B.n71 B.n70 585
R79 B.n69 B.n68 585
R80 B.n67 B.n66 585
R81 B.n65 B.n64 585
R82 B.n418 B.n26 585
R83 B.n422 B.n26 585
R84 B.n417 B.n25 585
R85 B.n423 B.n25 585
R86 B.n416 B.n415 585
R87 B.n415 B.n21 585
R88 B.n414 B.n20 585
R89 B.n429 B.n20 585
R90 B.n413 B.n19 585
R91 B.n430 B.n19 585
R92 B.n412 B.n18 585
R93 B.n431 B.n18 585
R94 B.n411 B.n410 585
R95 B.n410 B.n13 585
R96 B.n409 B.n12 585
R97 B.n437 B.n12 585
R98 B.n408 B.n11 585
R99 B.n438 B.n11 585
R100 B.n407 B.n10 585
R101 B.n439 B.n10 585
R102 B.n406 B.n7 585
R103 B.n442 B.n7 585
R104 B.n405 B.n6 585
R105 B.n443 B.n6 585
R106 B.n404 B.n5 585
R107 B.n444 B.n5 585
R108 B.n403 B.n402 585
R109 B.n402 B.n4 585
R110 B.n401 B.n188 585
R111 B.n401 B.n400 585
R112 B.n391 B.n189 585
R113 B.n190 B.n189 585
R114 B.n393 B.n392 585
R115 B.n394 B.n393 585
R116 B.n390 B.n195 585
R117 B.n195 B.n194 585
R118 B.n389 B.n388 585
R119 B.n388 B.n387 585
R120 B.n197 B.n196 585
R121 B.n380 B.n197 585
R122 B.n379 B.n378 585
R123 B.n381 B.n379 585
R124 B.n377 B.n202 585
R125 B.n202 B.n201 585
R126 B.n376 B.n375 585
R127 B.n375 B.n374 585
R128 B.n204 B.n203 585
R129 B.n205 B.n204 585
R130 B.n370 B.n369 585
R131 B.n208 B.n207 585
R132 B.n366 B.n365 585
R133 B.n367 B.n366 585
R134 B.n364 B.n239 585
R135 B.n363 B.n362 585
R136 B.n361 B.n360 585
R137 B.n359 B.n358 585
R138 B.n357 B.n356 585
R139 B.n355 B.n354 585
R140 B.n353 B.n352 585
R141 B.n351 B.n350 585
R142 B.n349 B.n348 585
R143 B.n347 B.n346 585
R144 B.n345 B.n344 585
R145 B.n343 B.n342 585
R146 B.n341 B.n340 585
R147 B.n339 B.n338 585
R148 B.n337 B.n336 585
R149 B.n335 B.n334 585
R150 B.n333 B.n332 585
R151 B.n331 B.n330 585
R152 B.n329 B.n328 585
R153 B.n327 B.n326 585
R154 B.n325 B.n324 585
R155 B.n323 B.n322 585
R156 B.n321 B.n320 585
R157 B.n319 B.n318 585
R158 B.n317 B.n316 585
R159 B.n315 B.n314 585
R160 B.n313 B.n312 585
R161 B.n311 B.n310 585
R162 B.n309 B.n308 585
R163 B.n307 B.n306 585
R164 B.n305 B.n304 585
R165 B.n303 B.n302 585
R166 B.n301 B.n300 585
R167 B.n298 B.n297 585
R168 B.n296 B.n295 585
R169 B.n294 B.n293 585
R170 B.n292 B.n291 585
R171 B.n290 B.n289 585
R172 B.n288 B.n287 585
R173 B.n286 B.n285 585
R174 B.n284 B.n283 585
R175 B.n282 B.n281 585
R176 B.n280 B.n279 585
R177 B.n278 B.n277 585
R178 B.n276 B.n275 585
R179 B.n274 B.n273 585
R180 B.n272 B.n271 585
R181 B.n270 B.n269 585
R182 B.n268 B.n267 585
R183 B.n266 B.n265 585
R184 B.n264 B.n263 585
R185 B.n262 B.n261 585
R186 B.n260 B.n259 585
R187 B.n258 B.n257 585
R188 B.n256 B.n255 585
R189 B.n254 B.n253 585
R190 B.n252 B.n251 585
R191 B.n250 B.n249 585
R192 B.n248 B.n247 585
R193 B.n246 B.n245 585
R194 B.n371 B.n206 585
R195 B.n206 B.n205 585
R196 B.n373 B.n372 585
R197 B.n374 B.n373 585
R198 B.n200 B.n199 585
R199 B.n201 B.n200 585
R200 B.n383 B.n382 585
R201 B.n382 B.n381 585
R202 B.n384 B.n198 585
R203 B.n380 B.n198 585
R204 B.n386 B.n385 585
R205 B.n387 B.n386 585
R206 B.n193 B.n192 585
R207 B.n194 B.n193 585
R208 B.n396 B.n395 585
R209 B.n395 B.n394 585
R210 B.n397 B.n191 585
R211 B.n191 B.n190 585
R212 B.n399 B.n398 585
R213 B.n400 B.n399 585
R214 B.n3 B.n0 585
R215 B.n4 B.n3 585
R216 B.n441 B.n1 585
R217 B.n442 B.n441 585
R218 B.n440 B.n9 585
R219 B.n440 B.n439 585
R220 B.n15 B.n8 585
R221 B.n438 B.n8 585
R222 B.n436 B.n435 585
R223 B.n437 B.n436 585
R224 B.n434 B.n14 585
R225 B.n14 B.n13 585
R226 B.n433 B.n432 585
R227 B.n432 B.n431 585
R228 B.n17 B.n16 585
R229 B.n430 B.n17 585
R230 B.n428 B.n427 585
R231 B.n429 B.n428 585
R232 B.n426 B.n22 585
R233 B.n22 B.n21 585
R234 B.n425 B.n424 585
R235 B.n424 B.n423 585
R236 B.n24 B.n23 585
R237 B.n422 B.n24 585
R238 B.n445 B.n444 585
R239 B.n443 B.n2 585
R240 B.n64 B.n24 487.695
R241 B.n420 B.n26 487.695
R242 B.n245 B.n204 487.695
R243 B.n369 B.n206 487.695
R244 B.n421 B.n57 256.663
R245 B.n421 B.n56 256.663
R246 B.n421 B.n55 256.663
R247 B.n421 B.n54 256.663
R248 B.n421 B.n53 256.663
R249 B.n421 B.n52 256.663
R250 B.n421 B.n51 256.663
R251 B.n421 B.n50 256.663
R252 B.n421 B.n49 256.663
R253 B.n421 B.n48 256.663
R254 B.n421 B.n47 256.663
R255 B.n421 B.n46 256.663
R256 B.n421 B.n45 256.663
R257 B.n421 B.n44 256.663
R258 B.n421 B.n43 256.663
R259 B.n421 B.n42 256.663
R260 B.n421 B.n41 256.663
R261 B.n421 B.n40 256.663
R262 B.n421 B.n39 256.663
R263 B.n421 B.n38 256.663
R264 B.n421 B.n37 256.663
R265 B.n421 B.n36 256.663
R266 B.n421 B.n35 256.663
R267 B.n421 B.n34 256.663
R268 B.n421 B.n33 256.663
R269 B.n421 B.n32 256.663
R270 B.n421 B.n31 256.663
R271 B.n421 B.n30 256.663
R272 B.n421 B.n29 256.663
R273 B.n421 B.n28 256.663
R274 B.n421 B.n27 256.663
R275 B.n368 B.n367 256.663
R276 B.n367 B.n209 256.663
R277 B.n367 B.n210 256.663
R278 B.n367 B.n211 256.663
R279 B.n367 B.n212 256.663
R280 B.n367 B.n213 256.663
R281 B.n367 B.n214 256.663
R282 B.n367 B.n215 256.663
R283 B.n367 B.n216 256.663
R284 B.n367 B.n217 256.663
R285 B.n367 B.n218 256.663
R286 B.n367 B.n219 256.663
R287 B.n367 B.n220 256.663
R288 B.n367 B.n221 256.663
R289 B.n367 B.n222 256.663
R290 B.n367 B.n223 256.663
R291 B.n367 B.n224 256.663
R292 B.n367 B.n225 256.663
R293 B.n367 B.n226 256.663
R294 B.n367 B.n227 256.663
R295 B.n367 B.n228 256.663
R296 B.n367 B.n229 256.663
R297 B.n367 B.n230 256.663
R298 B.n367 B.n231 256.663
R299 B.n367 B.n232 256.663
R300 B.n367 B.n233 256.663
R301 B.n367 B.n234 256.663
R302 B.n367 B.n235 256.663
R303 B.n367 B.n236 256.663
R304 B.n367 B.n237 256.663
R305 B.n367 B.n238 256.663
R306 B.n447 B.n446 256.663
R307 B.n68 B.n67 163.367
R308 B.n72 B.n71 163.367
R309 B.n76 B.n75 163.367
R310 B.n80 B.n79 163.367
R311 B.n84 B.n83 163.367
R312 B.n88 B.n87 163.367
R313 B.n92 B.n91 163.367
R314 B.n96 B.n95 163.367
R315 B.n100 B.n99 163.367
R316 B.n104 B.n103 163.367
R317 B.n108 B.n107 163.367
R318 B.n112 B.n111 163.367
R319 B.n116 B.n115 163.367
R320 B.n121 B.n120 163.367
R321 B.n125 B.n124 163.367
R322 B.n129 B.n128 163.367
R323 B.n133 B.n132 163.367
R324 B.n137 B.n136 163.367
R325 B.n141 B.n140 163.367
R326 B.n145 B.n144 163.367
R327 B.n149 B.n148 163.367
R328 B.n153 B.n152 163.367
R329 B.n157 B.n156 163.367
R330 B.n161 B.n160 163.367
R331 B.n165 B.n164 163.367
R332 B.n169 B.n168 163.367
R333 B.n173 B.n172 163.367
R334 B.n177 B.n176 163.367
R335 B.n181 B.n180 163.367
R336 B.n185 B.n184 163.367
R337 B.n420 B.n58 163.367
R338 B.n375 B.n204 163.367
R339 B.n375 B.n202 163.367
R340 B.n379 B.n202 163.367
R341 B.n379 B.n197 163.367
R342 B.n388 B.n197 163.367
R343 B.n388 B.n195 163.367
R344 B.n393 B.n195 163.367
R345 B.n393 B.n189 163.367
R346 B.n401 B.n189 163.367
R347 B.n402 B.n401 163.367
R348 B.n402 B.n5 163.367
R349 B.n6 B.n5 163.367
R350 B.n7 B.n6 163.367
R351 B.n10 B.n7 163.367
R352 B.n11 B.n10 163.367
R353 B.n12 B.n11 163.367
R354 B.n410 B.n12 163.367
R355 B.n410 B.n18 163.367
R356 B.n19 B.n18 163.367
R357 B.n20 B.n19 163.367
R358 B.n415 B.n20 163.367
R359 B.n415 B.n25 163.367
R360 B.n26 B.n25 163.367
R361 B.n366 B.n208 163.367
R362 B.n366 B.n239 163.367
R363 B.n362 B.n361 163.367
R364 B.n358 B.n357 163.367
R365 B.n354 B.n353 163.367
R366 B.n350 B.n349 163.367
R367 B.n346 B.n345 163.367
R368 B.n342 B.n341 163.367
R369 B.n338 B.n337 163.367
R370 B.n334 B.n333 163.367
R371 B.n330 B.n329 163.367
R372 B.n326 B.n325 163.367
R373 B.n322 B.n321 163.367
R374 B.n318 B.n317 163.367
R375 B.n314 B.n313 163.367
R376 B.n310 B.n309 163.367
R377 B.n306 B.n305 163.367
R378 B.n302 B.n301 163.367
R379 B.n297 B.n296 163.367
R380 B.n293 B.n292 163.367
R381 B.n289 B.n288 163.367
R382 B.n285 B.n284 163.367
R383 B.n281 B.n280 163.367
R384 B.n277 B.n276 163.367
R385 B.n273 B.n272 163.367
R386 B.n269 B.n268 163.367
R387 B.n265 B.n264 163.367
R388 B.n261 B.n260 163.367
R389 B.n257 B.n256 163.367
R390 B.n253 B.n252 163.367
R391 B.n249 B.n248 163.367
R392 B.n373 B.n206 163.367
R393 B.n373 B.n200 163.367
R394 B.n382 B.n200 163.367
R395 B.n382 B.n198 163.367
R396 B.n386 B.n198 163.367
R397 B.n386 B.n193 163.367
R398 B.n395 B.n193 163.367
R399 B.n395 B.n191 163.367
R400 B.n399 B.n191 163.367
R401 B.n399 B.n3 163.367
R402 B.n445 B.n3 163.367
R403 B.n441 B.n2 163.367
R404 B.n441 B.n440 163.367
R405 B.n440 B.n8 163.367
R406 B.n436 B.n8 163.367
R407 B.n436 B.n14 163.367
R408 B.n432 B.n14 163.367
R409 B.n432 B.n17 163.367
R410 B.n428 B.n17 163.367
R411 B.n428 B.n22 163.367
R412 B.n424 B.n22 163.367
R413 B.n424 B.n24 163.367
R414 B.n367 B.n205 112.936
R415 B.n422 B.n421 112.936
R416 B.n59 B.t7 81.8144
R417 B.n243 B.t12 81.8144
R418 B.n62 B.t4 81.8066
R419 B.n240 B.t15 81.8066
R420 B.n64 B.n27 71.676
R421 B.n68 B.n28 71.676
R422 B.n72 B.n29 71.676
R423 B.n76 B.n30 71.676
R424 B.n80 B.n31 71.676
R425 B.n84 B.n32 71.676
R426 B.n88 B.n33 71.676
R427 B.n92 B.n34 71.676
R428 B.n96 B.n35 71.676
R429 B.n100 B.n36 71.676
R430 B.n104 B.n37 71.676
R431 B.n108 B.n38 71.676
R432 B.n112 B.n39 71.676
R433 B.n116 B.n40 71.676
R434 B.n121 B.n41 71.676
R435 B.n125 B.n42 71.676
R436 B.n129 B.n43 71.676
R437 B.n133 B.n44 71.676
R438 B.n137 B.n45 71.676
R439 B.n141 B.n46 71.676
R440 B.n145 B.n47 71.676
R441 B.n149 B.n48 71.676
R442 B.n153 B.n49 71.676
R443 B.n157 B.n50 71.676
R444 B.n161 B.n51 71.676
R445 B.n165 B.n52 71.676
R446 B.n169 B.n53 71.676
R447 B.n173 B.n54 71.676
R448 B.n177 B.n55 71.676
R449 B.n181 B.n56 71.676
R450 B.n185 B.n57 71.676
R451 B.n58 B.n57 71.676
R452 B.n184 B.n56 71.676
R453 B.n180 B.n55 71.676
R454 B.n176 B.n54 71.676
R455 B.n172 B.n53 71.676
R456 B.n168 B.n52 71.676
R457 B.n164 B.n51 71.676
R458 B.n160 B.n50 71.676
R459 B.n156 B.n49 71.676
R460 B.n152 B.n48 71.676
R461 B.n148 B.n47 71.676
R462 B.n144 B.n46 71.676
R463 B.n140 B.n45 71.676
R464 B.n136 B.n44 71.676
R465 B.n132 B.n43 71.676
R466 B.n128 B.n42 71.676
R467 B.n124 B.n41 71.676
R468 B.n120 B.n40 71.676
R469 B.n115 B.n39 71.676
R470 B.n111 B.n38 71.676
R471 B.n107 B.n37 71.676
R472 B.n103 B.n36 71.676
R473 B.n99 B.n35 71.676
R474 B.n95 B.n34 71.676
R475 B.n91 B.n33 71.676
R476 B.n87 B.n32 71.676
R477 B.n83 B.n31 71.676
R478 B.n79 B.n30 71.676
R479 B.n75 B.n29 71.676
R480 B.n71 B.n28 71.676
R481 B.n67 B.n27 71.676
R482 B.n369 B.n368 71.676
R483 B.n239 B.n209 71.676
R484 B.n361 B.n210 71.676
R485 B.n357 B.n211 71.676
R486 B.n353 B.n212 71.676
R487 B.n349 B.n213 71.676
R488 B.n345 B.n214 71.676
R489 B.n341 B.n215 71.676
R490 B.n337 B.n216 71.676
R491 B.n333 B.n217 71.676
R492 B.n329 B.n218 71.676
R493 B.n325 B.n219 71.676
R494 B.n321 B.n220 71.676
R495 B.n317 B.n221 71.676
R496 B.n313 B.n222 71.676
R497 B.n309 B.n223 71.676
R498 B.n305 B.n224 71.676
R499 B.n301 B.n225 71.676
R500 B.n296 B.n226 71.676
R501 B.n292 B.n227 71.676
R502 B.n288 B.n228 71.676
R503 B.n284 B.n229 71.676
R504 B.n280 B.n230 71.676
R505 B.n276 B.n231 71.676
R506 B.n272 B.n232 71.676
R507 B.n268 B.n233 71.676
R508 B.n264 B.n234 71.676
R509 B.n260 B.n235 71.676
R510 B.n256 B.n236 71.676
R511 B.n252 B.n237 71.676
R512 B.n248 B.n238 71.676
R513 B.n368 B.n208 71.676
R514 B.n362 B.n209 71.676
R515 B.n358 B.n210 71.676
R516 B.n354 B.n211 71.676
R517 B.n350 B.n212 71.676
R518 B.n346 B.n213 71.676
R519 B.n342 B.n214 71.676
R520 B.n338 B.n215 71.676
R521 B.n334 B.n216 71.676
R522 B.n330 B.n217 71.676
R523 B.n326 B.n218 71.676
R524 B.n322 B.n219 71.676
R525 B.n318 B.n220 71.676
R526 B.n314 B.n221 71.676
R527 B.n310 B.n222 71.676
R528 B.n306 B.n223 71.676
R529 B.n302 B.n224 71.676
R530 B.n297 B.n225 71.676
R531 B.n293 B.n226 71.676
R532 B.n289 B.n227 71.676
R533 B.n285 B.n228 71.676
R534 B.n281 B.n229 71.676
R535 B.n277 B.n230 71.676
R536 B.n273 B.n231 71.676
R537 B.n269 B.n232 71.676
R538 B.n265 B.n233 71.676
R539 B.n261 B.n234 71.676
R540 B.n257 B.n235 71.676
R541 B.n253 B.n236 71.676
R542 B.n249 B.n237 71.676
R543 B.n245 B.n238 71.676
R544 B.n446 B.n445 71.676
R545 B.n446 B.n2 71.676
R546 B.n60 B.t8 70.5659
R547 B.n244 B.t11 70.5659
R548 B.n63 B.t5 70.5581
R549 B.n241 B.t14 70.5581
R550 B.n374 B.n205 61.4379
R551 B.n374 B.n201 61.4379
R552 B.n381 B.n201 61.4379
R553 B.n381 B.n380 61.4379
R554 B.n387 B.n194 61.4379
R555 B.n394 B.n194 61.4379
R556 B.n394 B.n190 61.4379
R557 B.n400 B.n190 61.4379
R558 B.n444 B.n4 61.4379
R559 B.n444 B.n443 61.4379
R560 B.n443 B.n442 61.4379
R561 B.n439 B.n438 61.4379
R562 B.n438 B.n437 61.4379
R563 B.n437 B.n13 61.4379
R564 B.n431 B.n13 61.4379
R565 B.n430 B.n429 61.4379
R566 B.n429 B.n21 61.4379
R567 B.n423 B.n21 61.4379
R568 B.n423 B.n422 61.4379
R569 B.n118 B.n63 59.5399
R570 B.n61 B.n60 59.5399
R571 B.n299 B.n244 59.5399
R572 B.n242 B.n241 59.5399
R573 B.t1 B.n4 58.7274
R574 B.n442 B.t0 58.7274
R575 B.n387 B.t10 53.3065
R576 B.n431 B.t3 53.3065
R577 B.n371 B.n370 31.6883
R578 B.n246 B.n203 31.6883
R579 B.n419 B.n418 31.6883
R580 B.n65 B.n23 31.6883
R581 B B.n447 18.0485
R582 B.n63 B.n62 11.249
R583 B.n60 B.n59 11.249
R584 B.n244 B.n243 11.249
R585 B.n241 B.n240 11.249
R586 B.n372 B.n371 10.6151
R587 B.n372 B.n199 10.6151
R588 B.n383 B.n199 10.6151
R589 B.n384 B.n383 10.6151
R590 B.n385 B.n384 10.6151
R591 B.n385 B.n192 10.6151
R592 B.n396 B.n192 10.6151
R593 B.n397 B.n396 10.6151
R594 B.n398 B.n397 10.6151
R595 B.n398 B.n0 10.6151
R596 B.n370 B.n207 10.6151
R597 B.n365 B.n207 10.6151
R598 B.n365 B.n364 10.6151
R599 B.n364 B.n363 10.6151
R600 B.n363 B.n360 10.6151
R601 B.n360 B.n359 10.6151
R602 B.n359 B.n356 10.6151
R603 B.n356 B.n355 10.6151
R604 B.n355 B.n352 10.6151
R605 B.n352 B.n351 10.6151
R606 B.n351 B.n348 10.6151
R607 B.n348 B.n347 10.6151
R608 B.n347 B.n344 10.6151
R609 B.n344 B.n343 10.6151
R610 B.n343 B.n340 10.6151
R611 B.n340 B.n339 10.6151
R612 B.n339 B.n336 10.6151
R613 B.n336 B.n335 10.6151
R614 B.n335 B.n332 10.6151
R615 B.n332 B.n331 10.6151
R616 B.n331 B.n328 10.6151
R617 B.n328 B.n327 10.6151
R618 B.n327 B.n324 10.6151
R619 B.n324 B.n323 10.6151
R620 B.n323 B.n320 10.6151
R621 B.n320 B.n319 10.6151
R622 B.n316 B.n315 10.6151
R623 B.n315 B.n312 10.6151
R624 B.n312 B.n311 10.6151
R625 B.n311 B.n308 10.6151
R626 B.n308 B.n307 10.6151
R627 B.n307 B.n304 10.6151
R628 B.n304 B.n303 10.6151
R629 B.n303 B.n300 10.6151
R630 B.n298 B.n295 10.6151
R631 B.n295 B.n294 10.6151
R632 B.n294 B.n291 10.6151
R633 B.n291 B.n290 10.6151
R634 B.n290 B.n287 10.6151
R635 B.n287 B.n286 10.6151
R636 B.n286 B.n283 10.6151
R637 B.n283 B.n282 10.6151
R638 B.n282 B.n279 10.6151
R639 B.n279 B.n278 10.6151
R640 B.n278 B.n275 10.6151
R641 B.n275 B.n274 10.6151
R642 B.n274 B.n271 10.6151
R643 B.n271 B.n270 10.6151
R644 B.n270 B.n267 10.6151
R645 B.n267 B.n266 10.6151
R646 B.n266 B.n263 10.6151
R647 B.n263 B.n262 10.6151
R648 B.n262 B.n259 10.6151
R649 B.n259 B.n258 10.6151
R650 B.n258 B.n255 10.6151
R651 B.n255 B.n254 10.6151
R652 B.n254 B.n251 10.6151
R653 B.n251 B.n250 10.6151
R654 B.n250 B.n247 10.6151
R655 B.n247 B.n246 10.6151
R656 B.n376 B.n203 10.6151
R657 B.n377 B.n376 10.6151
R658 B.n378 B.n377 10.6151
R659 B.n378 B.n196 10.6151
R660 B.n389 B.n196 10.6151
R661 B.n390 B.n389 10.6151
R662 B.n392 B.n390 10.6151
R663 B.n392 B.n391 10.6151
R664 B.n391 B.n188 10.6151
R665 B.n403 B.n188 10.6151
R666 B.n404 B.n403 10.6151
R667 B.n405 B.n404 10.6151
R668 B.n406 B.n405 10.6151
R669 B.n407 B.n406 10.6151
R670 B.n408 B.n407 10.6151
R671 B.n409 B.n408 10.6151
R672 B.n411 B.n409 10.6151
R673 B.n412 B.n411 10.6151
R674 B.n413 B.n412 10.6151
R675 B.n414 B.n413 10.6151
R676 B.n416 B.n414 10.6151
R677 B.n417 B.n416 10.6151
R678 B.n418 B.n417 10.6151
R679 B.n9 B.n1 10.6151
R680 B.n15 B.n9 10.6151
R681 B.n435 B.n15 10.6151
R682 B.n435 B.n434 10.6151
R683 B.n434 B.n433 10.6151
R684 B.n433 B.n16 10.6151
R685 B.n427 B.n16 10.6151
R686 B.n427 B.n426 10.6151
R687 B.n426 B.n425 10.6151
R688 B.n425 B.n23 10.6151
R689 B.n66 B.n65 10.6151
R690 B.n69 B.n66 10.6151
R691 B.n70 B.n69 10.6151
R692 B.n73 B.n70 10.6151
R693 B.n74 B.n73 10.6151
R694 B.n77 B.n74 10.6151
R695 B.n78 B.n77 10.6151
R696 B.n81 B.n78 10.6151
R697 B.n82 B.n81 10.6151
R698 B.n85 B.n82 10.6151
R699 B.n86 B.n85 10.6151
R700 B.n89 B.n86 10.6151
R701 B.n90 B.n89 10.6151
R702 B.n93 B.n90 10.6151
R703 B.n94 B.n93 10.6151
R704 B.n97 B.n94 10.6151
R705 B.n98 B.n97 10.6151
R706 B.n101 B.n98 10.6151
R707 B.n102 B.n101 10.6151
R708 B.n105 B.n102 10.6151
R709 B.n106 B.n105 10.6151
R710 B.n109 B.n106 10.6151
R711 B.n110 B.n109 10.6151
R712 B.n113 B.n110 10.6151
R713 B.n114 B.n113 10.6151
R714 B.n117 B.n114 10.6151
R715 B.n122 B.n119 10.6151
R716 B.n123 B.n122 10.6151
R717 B.n126 B.n123 10.6151
R718 B.n127 B.n126 10.6151
R719 B.n130 B.n127 10.6151
R720 B.n131 B.n130 10.6151
R721 B.n134 B.n131 10.6151
R722 B.n135 B.n134 10.6151
R723 B.n139 B.n138 10.6151
R724 B.n142 B.n139 10.6151
R725 B.n143 B.n142 10.6151
R726 B.n146 B.n143 10.6151
R727 B.n147 B.n146 10.6151
R728 B.n150 B.n147 10.6151
R729 B.n151 B.n150 10.6151
R730 B.n154 B.n151 10.6151
R731 B.n155 B.n154 10.6151
R732 B.n158 B.n155 10.6151
R733 B.n159 B.n158 10.6151
R734 B.n162 B.n159 10.6151
R735 B.n163 B.n162 10.6151
R736 B.n166 B.n163 10.6151
R737 B.n167 B.n166 10.6151
R738 B.n170 B.n167 10.6151
R739 B.n171 B.n170 10.6151
R740 B.n174 B.n171 10.6151
R741 B.n175 B.n174 10.6151
R742 B.n178 B.n175 10.6151
R743 B.n179 B.n178 10.6151
R744 B.n182 B.n179 10.6151
R745 B.n183 B.n182 10.6151
R746 B.n186 B.n183 10.6151
R747 B.n187 B.n186 10.6151
R748 B.n419 B.n187 10.6151
R749 B.n380 B.t10 8.13192
R750 B.t3 B.n430 8.13192
R751 B.n447 B.n0 8.11757
R752 B.n447 B.n1 8.11757
R753 B.n316 B.n242 7.18099
R754 B.n300 B.n299 7.18099
R755 B.n119 B.n118 7.18099
R756 B.n135 B.n61 7.18099
R757 B.n319 B.n242 3.43465
R758 B.n299 B.n298 3.43465
R759 B.n118 B.n117 3.43465
R760 B.n138 B.n61 3.43465
R761 B.n400 B.t1 2.71097
R762 B.n439 B.t0 2.71097
R763 VP.n0 VP.t1 1008.51
R764 VP.n0 VP.t0 973.952
R765 VP VP.n0 0.0516364
R766 VDD1 VDD1.t1 102.258
R767 VDD1 VDD1.t0 71.1839
C0 VN VDD2 0.872326f
C1 VTAIL VN 0.556889f
C2 VN VP 3.41268f
C3 VN VDD1 0.148705f
C4 VTAIL VDD2 4.68437f
C5 VP VDD2 0.235747f
C6 VDD1 VDD2 0.420497f
C7 VTAIL VP 0.571383f
C8 VTAIL VDD1 4.65187f
C9 VP VDD1 0.956408f
C10 VDD2 B 2.659269f
C11 VDD1 B 4.80176f
C12 VTAIL B 3.824967f
C13 VN B 6.08262f
C14 VP B 3.130516f
C15 VDD1.t0 B 1.17248f
C16 VDD1.t1 B 1.47281f
C17 VP.t1 B 0.295603f
C18 VP.t0 B 0.246635f
C19 VP.n0 B 2.8522f
C20 VDD2.t0 B 1.47778f
C21 VDD2.t1 B 1.19048f
C22 VDD2.n0 B 2.00302f
C23 VTAIL.t1 B 1.25055f
C24 VTAIL.n0 B 1.11263f
C25 VTAIL.t3 B 1.25056f
C26 VTAIL.n1 B 1.11743f
C27 VTAIL.t0 B 1.25055f
C28 VTAIL.n2 B 1.08146f
C29 VTAIL.t2 B 1.25055f
C30 VTAIL.n3 B 1.03447f
C31 VN.t1 B 0.242009f
C32 VN.t0 B 0.29161f
.ends

