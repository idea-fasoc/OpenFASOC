* NGSPICE file created from diff_pair_sample_1712.ext - technology: sky130A

.subckt diff_pair_sample_1712 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=0 ps=0 w=19.62 l=2.19
X1 VDD1.t7 VP.t0 VTAIL.t9 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=7.6518 ps=40.02 w=19.62 l=2.19
X2 VTAIL.t10 VP.t1 VDD1.t6 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X3 VTAIL.t2 VN.t0 VDD2.t7 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=3.2373 ps=19.95 w=19.62 l=2.19
X4 VDD2.t6 VN.t1 VTAIL.t0 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=7.6518 ps=40.02 w=19.62 l=2.19
X5 VTAIL.t1 VN.t2 VDD2.t5 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X6 VDD1.t5 VP.t2 VTAIL.t13 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X7 VTAIL.t12 VP.t3 VDD1.t4 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X8 VDD2.t4 VN.t3 VTAIL.t6 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=7.6518 ps=40.02 w=19.62 l=2.19
X9 VTAIL.t15 VP.t4 VDD1.t3 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=3.2373 ps=19.95 w=19.62 l=2.19
X10 VTAIL.t4 VN.t4 VDD2.t3 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X11 B.t8 B.t6 B.t7 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=0 ps=0 w=19.62 l=2.19
X12 B.t5 B.t3 B.t4 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=0 ps=0 w=19.62 l=2.19
X13 VTAIL.t7 VN.t5 VDD2.t2 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=3.2373 ps=19.95 w=19.62 l=2.19
X14 B.t2 B.t0 B.t1 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=0 ps=0 w=19.62 l=2.19
X15 VTAIL.t8 VP.t5 VDD1.t2 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=7.6518 pd=40.02 as=3.2373 ps=19.95 w=19.62 l=2.19
X16 VDD2.t1 VN.t6 VTAIL.t3 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X17 VDD1.t1 VP.t6 VTAIL.t14 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X18 VDD2.t0 VN.t7 VTAIL.t5 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=3.2373 ps=19.95 w=19.62 l=2.19
X19 VDD1.t0 VP.t7 VTAIL.t11 w_n3490_n4892# sky130_fd_pr__pfet_01v8 ad=3.2373 pd=19.95 as=7.6518 ps=40.02 w=19.62 l=2.19
R0 B.n651 B.n98 585
R1 B.n653 B.n652 585
R2 B.n654 B.n97 585
R3 B.n656 B.n655 585
R4 B.n657 B.n96 585
R5 B.n659 B.n658 585
R6 B.n660 B.n95 585
R7 B.n662 B.n661 585
R8 B.n663 B.n94 585
R9 B.n665 B.n664 585
R10 B.n666 B.n93 585
R11 B.n668 B.n667 585
R12 B.n669 B.n92 585
R13 B.n671 B.n670 585
R14 B.n672 B.n91 585
R15 B.n674 B.n673 585
R16 B.n675 B.n90 585
R17 B.n677 B.n676 585
R18 B.n678 B.n89 585
R19 B.n680 B.n679 585
R20 B.n681 B.n88 585
R21 B.n683 B.n682 585
R22 B.n684 B.n87 585
R23 B.n686 B.n685 585
R24 B.n687 B.n86 585
R25 B.n689 B.n688 585
R26 B.n690 B.n85 585
R27 B.n692 B.n691 585
R28 B.n693 B.n84 585
R29 B.n695 B.n694 585
R30 B.n696 B.n83 585
R31 B.n698 B.n697 585
R32 B.n699 B.n82 585
R33 B.n701 B.n700 585
R34 B.n702 B.n81 585
R35 B.n704 B.n703 585
R36 B.n705 B.n80 585
R37 B.n707 B.n706 585
R38 B.n708 B.n79 585
R39 B.n710 B.n709 585
R40 B.n711 B.n78 585
R41 B.n713 B.n712 585
R42 B.n714 B.n77 585
R43 B.n716 B.n715 585
R44 B.n717 B.n76 585
R45 B.n719 B.n718 585
R46 B.n720 B.n75 585
R47 B.n722 B.n721 585
R48 B.n723 B.n74 585
R49 B.n725 B.n724 585
R50 B.n726 B.n73 585
R51 B.n728 B.n727 585
R52 B.n729 B.n72 585
R53 B.n731 B.n730 585
R54 B.n732 B.n71 585
R55 B.n734 B.n733 585
R56 B.n735 B.n70 585
R57 B.n737 B.n736 585
R58 B.n738 B.n69 585
R59 B.n740 B.n739 585
R60 B.n741 B.n68 585
R61 B.n743 B.n742 585
R62 B.n744 B.n67 585
R63 B.n746 B.n745 585
R64 B.n748 B.n64 585
R65 B.n750 B.n749 585
R66 B.n751 B.n63 585
R67 B.n753 B.n752 585
R68 B.n754 B.n62 585
R69 B.n756 B.n755 585
R70 B.n757 B.n61 585
R71 B.n759 B.n758 585
R72 B.n760 B.n57 585
R73 B.n762 B.n761 585
R74 B.n763 B.n56 585
R75 B.n765 B.n764 585
R76 B.n766 B.n55 585
R77 B.n768 B.n767 585
R78 B.n769 B.n54 585
R79 B.n771 B.n770 585
R80 B.n772 B.n53 585
R81 B.n774 B.n773 585
R82 B.n775 B.n52 585
R83 B.n777 B.n776 585
R84 B.n778 B.n51 585
R85 B.n780 B.n779 585
R86 B.n781 B.n50 585
R87 B.n783 B.n782 585
R88 B.n784 B.n49 585
R89 B.n786 B.n785 585
R90 B.n787 B.n48 585
R91 B.n789 B.n788 585
R92 B.n790 B.n47 585
R93 B.n792 B.n791 585
R94 B.n793 B.n46 585
R95 B.n795 B.n794 585
R96 B.n796 B.n45 585
R97 B.n798 B.n797 585
R98 B.n799 B.n44 585
R99 B.n801 B.n800 585
R100 B.n802 B.n43 585
R101 B.n804 B.n803 585
R102 B.n805 B.n42 585
R103 B.n807 B.n806 585
R104 B.n808 B.n41 585
R105 B.n810 B.n809 585
R106 B.n811 B.n40 585
R107 B.n813 B.n812 585
R108 B.n814 B.n39 585
R109 B.n816 B.n815 585
R110 B.n817 B.n38 585
R111 B.n819 B.n818 585
R112 B.n820 B.n37 585
R113 B.n822 B.n821 585
R114 B.n823 B.n36 585
R115 B.n825 B.n824 585
R116 B.n826 B.n35 585
R117 B.n828 B.n827 585
R118 B.n829 B.n34 585
R119 B.n831 B.n830 585
R120 B.n832 B.n33 585
R121 B.n834 B.n833 585
R122 B.n835 B.n32 585
R123 B.n837 B.n836 585
R124 B.n838 B.n31 585
R125 B.n840 B.n839 585
R126 B.n841 B.n30 585
R127 B.n843 B.n842 585
R128 B.n844 B.n29 585
R129 B.n846 B.n845 585
R130 B.n847 B.n28 585
R131 B.n849 B.n848 585
R132 B.n850 B.n27 585
R133 B.n852 B.n851 585
R134 B.n853 B.n26 585
R135 B.n855 B.n854 585
R136 B.n856 B.n25 585
R137 B.n858 B.n857 585
R138 B.n650 B.n649 585
R139 B.n648 B.n99 585
R140 B.n647 B.n646 585
R141 B.n645 B.n100 585
R142 B.n644 B.n643 585
R143 B.n642 B.n101 585
R144 B.n641 B.n640 585
R145 B.n639 B.n102 585
R146 B.n638 B.n637 585
R147 B.n636 B.n103 585
R148 B.n635 B.n634 585
R149 B.n633 B.n104 585
R150 B.n632 B.n631 585
R151 B.n630 B.n105 585
R152 B.n629 B.n628 585
R153 B.n627 B.n106 585
R154 B.n626 B.n625 585
R155 B.n624 B.n107 585
R156 B.n623 B.n622 585
R157 B.n621 B.n108 585
R158 B.n620 B.n619 585
R159 B.n618 B.n109 585
R160 B.n617 B.n616 585
R161 B.n615 B.n110 585
R162 B.n614 B.n613 585
R163 B.n612 B.n111 585
R164 B.n611 B.n610 585
R165 B.n609 B.n112 585
R166 B.n608 B.n607 585
R167 B.n606 B.n113 585
R168 B.n605 B.n604 585
R169 B.n603 B.n114 585
R170 B.n602 B.n601 585
R171 B.n600 B.n115 585
R172 B.n599 B.n598 585
R173 B.n597 B.n116 585
R174 B.n596 B.n595 585
R175 B.n594 B.n117 585
R176 B.n593 B.n592 585
R177 B.n591 B.n118 585
R178 B.n590 B.n589 585
R179 B.n588 B.n119 585
R180 B.n587 B.n586 585
R181 B.n585 B.n120 585
R182 B.n584 B.n583 585
R183 B.n582 B.n121 585
R184 B.n581 B.n580 585
R185 B.n579 B.n122 585
R186 B.n578 B.n577 585
R187 B.n576 B.n123 585
R188 B.n575 B.n574 585
R189 B.n573 B.n124 585
R190 B.n572 B.n571 585
R191 B.n570 B.n125 585
R192 B.n569 B.n568 585
R193 B.n567 B.n126 585
R194 B.n566 B.n565 585
R195 B.n564 B.n127 585
R196 B.n563 B.n562 585
R197 B.n561 B.n128 585
R198 B.n560 B.n559 585
R199 B.n558 B.n129 585
R200 B.n557 B.n556 585
R201 B.n555 B.n130 585
R202 B.n554 B.n553 585
R203 B.n552 B.n131 585
R204 B.n551 B.n550 585
R205 B.n549 B.n132 585
R206 B.n548 B.n547 585
R207 B.n546 B.n133 585
R208 B.n545 B.n544 585
R209 B.n543 B.n134 585
R210 B.n542 B.n541 585
R211 B.n540 B.n135 585
R212 B.n539 B.n538 585
R213 B.n537 B.n136 585
R214 B.n536 B.n535 585
R215 B.n534 B.n137 585
R216 B.n533 B.n532 585
R217 B.n531 B.n138 585
R218 B.n530 B.n529 585
R219 B.n528 B.n139 585
R220 B.n527 B.n526 585
R221 B.n525 B.n140 585
R222 B.n524 B.n523 585
R223 B.n522 B.n141 585
R224 B.n521 B.n520 585
R225 B.n519 B.n142 585
R226 B.n518 B.n517 585
R227 B.n516 B.n143 585
R228 B.n515 B.n514 585
R229 B.n306 B.n217 585
R230 B.n308 B.n307 585
R231 B.n309 B.n216 585
R232 B.n311 B.n310 585
R233 B.n312 B.n215 585
R234 B.n314 B.n313 585
R235 B.n315 B.n214 585
R236 B.n317 B.n316 585
R237 B.n318 B.n213 585
R238 B.n320 B.n319 585
R239 B.n321 B.n212 585
R240 B.n323 B.n322 585
R241 B.n324 B.n211 585
R242 B.n326 B.n325 585
R243 B.n327 B.n210 585
R244 B.n329 B.n328 585
R245 B.n330 B.n209 585
R246 B.n332 B.n331 585
R247 B.n333 B.n208 585
R248 B.n335 B.n334 585
R249 B.n336 B.n207 585
R250 B.n338 B.n337 585
R251 B.n339 B.n206 585
R252 B.n341 B.n340 585
R253 B.n342 B.n205 585
R254 B.n344 B.n343 585
R255 B.n345 B.n204 585
R256 B.n347 B.n346 585
R257 B.n348 B.n203 585
R258 B.n350 B.n349 585
R259 B.n351 B.n202 585
R260 B.n353 B.n352 585
R261 B.n354 B.n201 585
R262 B.n356 B.n355 585
R263 B.n357 B.n200 585
R264 B.n359 B.n358 585
R265 B.n360 B.n199 585
R266 B.n362 B.n361 585
R267 B.n363 B.n198 585
R268 B.n365 B.n364 585
R269 B.n366 B.n197 585
R270 B.n368 B.n367 585
R271 B.n369 B.n196 585
R272 B.n371 B.n370 585
R273 B.n372 B.n195 585
R274 B.n374 B.n373 585
R275 B.n375 B.n194 585
R276 B.n377 B.n376 585
R277 B.n378 B.n193 585
R278 B.n380 B.n379 585
R279 B.n381 B.n192 585
R280 B.n383 B.n382 585
R281 B.n384 B.n191 585
R282 B.n386 B.n385 585
R283 B.n387 B.n190 585
R284 B.n389 B.n388 585
R285 B.n390 B.n189 585
R286 B.n392 B.n391 585
R287 B.n393 B.n188 585
R288 B.n395 B.n394 585
R289 B.n396 B.n187 585
R290 B.n398 B.n397 585
R291 B.n399 B.n186 585
R292 B.n401 B.n400 585
R293 B.n403 B.n402 585
R294 B.n404 B.n182 585
R295 B.n406 B.n405 585
R296 B.n407 B.n181 585
R297 B.n409 B.n408 585
R298 B.n410 B.n180 585
R299 B.n412 B.n411 585
R300 B.n413 B.n179 585
R301 B.n415 B.n414 585
R302 B.n416 B.n176 585
R303 B.n419 B.n418 585
R304 B.n420 B.n175 585
R305 B.n422 B.n421 585
R306 B.n423 B.n174 585
R307 B.n425 B.n424 585
R308 B.n426 B.n173 585
R309 B.n428 B.n427 585
R310 B.n429 B.n172 585
R311 B.n431 B.n430 585
R312 B.n432 B.n171 585
R313 B.n434 B.n433 585
R314 B.n435 B.n170 585
R315 B.n437 B.n436 585
R316 B.n438 B.n169 585
R317 B.n440 B.n439 585
R318 B.n441 B.n168 585
R319 B.n443 B.n442 585
R320 B.n444 B.n167 585
R321 B.n446 B.n445 585
R322 B.n447 B.n166 585
R323 B.n449 B.n448 585
R324 B.n450 B.n165 585
R325 B.n452 B.n451 585
R326 B.n453 B.n164 585
R327 B.n455 B.n454 585
R328 B.n456 B.n163 585
R329 B.n458 B.n457 585
R330 B.n459 B.n162 585
R331 B.n461 B.n460 585
R332 B.n462 B.n161 585
R333 B.n464 B.n463 585
R334 B.n465 B.n160 585
R335 B.n467 B.n466 585
R336 B.n468 B.n159 585
R337 B.n470 B.n469 585
R338 B.n471 B.n158 585
R339 B.n473 B.n472 585
R340 B.n474 B.n157 585
R341 B.n476 B.n475 585
R342 B.n477 B.n156 585
R343 B.n479 B.n478 585
R344 B.n480 B.n155 585
R345 B.n482 B.n481 585
R346 B.n483 B.n154 585
R347 B.n485 B.n484 585
R348 B.n486 B.n153 585
R349 B.n488 B.n487 585
R350 B.n489 B.n152 585
R351 B.n491 B.n490 585
R352 B.n492 B.n151 585
R353 B.n494 B.n493 585
R354 B.n495 B.n150 585
R355 B.n497 B.n496 585
R356 B.n498 B.n149 585
R357 B.n500 B.n499 585
R358 B.n501 B.n148 585
R359 B.n503 B.n502 585
R360 B.n504 B.n147 585
R361 B.n506 B.n505 585
R362 B.n507 B.n146 585
R363 B.n509 B.n508 585
R364 B.n510 B.n145 585
R365 B.n512 B.n511 585
R366 B.n513 B.n144 585
R367 B.n305 B.n304 585
R368 B.n303 B.n218 585
R369 B.n302 B.n301 585
R370 B.n300 B.n219 585
R371 B.n299 B.n298 585
R372 B.n297 B.n220 585
R373 B.n296 B.n295 585
R374 B.n294 B.n221 585
R375 B.n293 B.n292 585
R376 B.n291 B.n222 585
R377 B.n290 B.n289 585
R378 B.n288 B.n223 585
R379 B.n287 B.n286 585
R380 B.n285 B.n224 585
R381 B.n284 B.n283 585
R382 B.n282 B.n225 585
R383 B.n281 B.n280 585
R384 B.n279 B.n226 585
R385 B.n278 B.n277 585
R386 B.n276 B.n227 585
R387 B.n275 B.n274 585
R388 B.n273 B.n228 585
R389 B.n272 B.n271 585
R390 B.n270 B.n229 585
R391 B.n269 B.n268 585
R392 B.n267 B.n230 585
R393 B.n266 B.n265 585
R394 B.n264 B.n231 585
R395 B.n263 B.n262 585
R396 B.n261 B.n232 585
R397 B.n260 B.n259 585
R398 B.n258 B.n233 585
R399 B.n257 B.n256 585
R400 B.n255 B.n234 585
R401 B.n254 B.n253 585
R402 B.n252 B.n235 585
R403 B.n251 B.n250 585
R404 B.n249 B.n236 585
R405 B.n248 B.n247 585
R406 B.n246 B.n237 585
R407 B.n245 B.n244 585
R408 B.n243 B.n238 585
R409 B.n242 B.n241 585
R410 B.n240 B.n239 585
R411 B.n2 B.n0 585
R412 B.n925 B.n1 585
R413 B.n924 B.n923 585
R414 B.n922 B.n3 585
R415 B.n921 B.n920 585
R416 B.n919 B.n4 585
R417 B.n918 B.n917 585
R418 B.n916 B.n5 585
R419 B.n915 B.n914 585
R420 B.n913 B.n6 585
R421 B.n912 B.n911 585
R422 B.n910 B.n7 585
R423 B.n909 B.n908 585
R424 B.n907 B.n8 585
R425 B.n906 B.n905 585
R426 B.n904 B.n9 585
R427 B.n903 B.n902 585
R428 B.n901 B.n10 585
R429 B.n900 B.n899 585
R430 B.n898 B.n11 585
R431 B.n897 B.n896 585
R432 B.n895 B.n12 585
R433 B.n894 B.n893 585
R434 B.n892 B.n13 585
R435 B.n891 B.n890 585
R436 B.n889 B.n14 585
R437 B.n888 B.n887 585
R438 B.n886 B.n15 585
R439 B.n885 B.n884 585
R440 B.n883 B.n16 585
R441 B.n882 B.n881 585
R442 B.n880 B.n17 585
R443 B.n879 B.n878 585
R444 B.n877 B.n18 585
R445 B.n876 B.n875 585
R446 B.n874 B.n19 585
R447 B.n873 B.n872 585
R448 B.n871 B.n20 585
R449 B.n870 B.n869 585
R450 B.n868 B.n21 585
R451 B.n867 B.n866 585
R452 B.n865 B.n22 585
R453 B.n864 B.n863 585
R454 B.n862 B.n23 585
R455 B.n861 B.n860 585
R456 B.n859 B.n24 585
R457 B.n927 B.n926 585
R458 B.n177 B.t5 561.846
R459 B.n65 B.t1 561.846
R460 B.n183 B.t8 561.846
R461 B.n58 B.t10 561.846
R462 B.n178 B.t4 512.973
R463 B.n66 B.t2 512.973
R464 B.n184 B.t7 512.973
R465 B.n59 B.t11 512.973
R466 B.n306 B.n305 497.305
R467 B.n859 B.n858 497.305
R468 B.n515 B.n144 497.305
R469 B.n649 B.n98 497.305
R470 B.n177 B.t3 423.241
R471 B.n183 B.t6 423.241
R472 B.n58 B.t9 423.241
R473 B.n65 B.t0 423.241
R474 B.n305 B.n218 163.367
R475 B.n301 B.n218 163.367
R476 B.n301 B.n300 163.367
R477 B.n300 B.n299 163.367
R478 B.n299 B.n220 163.367
R479 B.n295 B.n220 163.367
R480 B.n295 B.n294 163.367
R481 B.n294 B.n293 163.367
R482 B.n293 B.n222 163.367
R483 B.n289 B.n222 163.367
R484 B.n289 B.n288 163.367
R485 B.n288 B.n287 163.367
R486 B.n287 B.n224 163.367
R487 B.n283 B.n224 163.367
R488 B.n283 B.n282 163.367
R489 B.n282 B.n281 163.367
R490 B.n281 B.n226 163.367
R491 B.n277 B.n226 163.367
R492 B.n277 B.n276 163.367
R493 B.n276 B.n275 163.367
R494 B.n275 B.n228 163.367
R495 B.n271 B.n228 163.367
R496 B.n271 B.n270 163.367
R497 B.n270 B.n269 163.367
R498 B.n269 B.n230 163.367
R499 B.n265 B.n230 163.367
R500 B.n265 B.n264 163.367
R501 B.n264 B.n263 163.367
R502 B.n263 B.n232 163.367
R503 B.n259 B.n232 163.367
R504 B.n259 B.n258 163.367
R505 B.n258 B.n257 163.367
R506 B.n257 B.n234 163.367
R507 B.n253 B.n234 163.367
R508 B.n253 B.n252 163.367
R509 B.n252 B.n251 163.367
R510 B.n251 B.n236 163.367
R511 B.n247 B.n236 163.367
R512 B.n247 B.n246 163.367
R513 B.n246 B.n245 163.367
R514 B.n245 B.n238 163.367
R515 B.n241 B.n238 163.367
R516 B.n241 B.n240 163.367
R517 B.n240 B.n2 163.367
R518 B.n926 B.n2 163.367
R519 B.n926 B.n925 163.367
R520 B.n925 B.n924 163.367
R521 B.n924 B.n3 163.367
R522 B.n920 B.n3 163.367
R523 B.n920 B.n919 163.367
R524 B.n919 B.n918 163.367
R525 B.n918 B.n5 163.367
R526 B.n914 B.n5 163.367
R527 B.n914 B.n913 163.367
R528 B.n913 B.n912 163.367
R529 B.n912 B.n7 163.367
R530 B.n908 B.n7 163.367
R531 B.n908 B.n907 163.367
R532 B.n907 B.n906 163.367
R533 B.n906 B.n9 163.367
R534 B.n902 B.n9 163.367
R535 B.n902 B.n901 163.367
R536 B.n901 B.n900 163.367
R537 B.n900 B.n11 163.367
R538 B.n896 B.n11 163.367
R539 B.n896 B.n895 163.367
R540 B.n895 B.n894 163.367
R541 B.n894 B.n13 163.367
R542 B.n890 B.n13 163.367
R543 B.n890 B.n889 163.367
R544 B.n889 B.n888 163.367
R545 B.n888 B.n15 163.367
R546 B.n884 B.n15 163.367
R547 B.n884 B.n883 163.367
R548 B.n883 B.n882 163.367
R549 B.n882 B.n17 163.367
R550 B.n878 B.n17 163.367
R551 B.n878 B.n877 163.367
R552 B.n877 B.n876 163.367
R553 B.n876 B.n19 163.367
R554 B.n872 B.n19 163.367
R555 B.n872 B.n871 163.367
R556 B.n871 B.n870 163.367
R557 B.n870 B.n21 163.367
R558 B.n866 B.n21 163.367
R559 B.n866 B.n865 163.367
R560 B.n865 B.n864 163.367
R561 B.n864 B.n23 163.367
R562 B.n860 B.n23 163.367
R563 B.n860 B.n859 163.367
R564 B.n307 B.n306 163.367
R565 B.n307 B.n216 163.367
R566 B.n311 B.n216 163.367
R567 B.n312 B.n311 163.367
R568 B.n313 B.n312 163.367
R569 B.n313 B.n214 163.367
R570 B.n317 B.n214 163.367
R571 B.n318 B.n317 163.367
R572 B.n319 B.n318 163.367
R573 B.n319 B.n212 163.367
R574 B.n323 B.n212 163.367
R575 B.n324 B.n323 163.367
R576 B.n325 B.n324 163.367
R577 B.n325 B.n210 163.367
R578 B.n329 B.n210 163.367
R579 B.n330 B.n329 163.367
R580 B.n331 B.n330 163.367
R581 B.n331 B.n208 163.367
R582 B.n335 B.n208 163.367
R583 B.n336 B.n335 163.367
R584 B.n337 B.n336 163.367
R585 B.n337 B.n206 163.367
R586 B.n341 B.n206 163.367
R587 B.n342 B.n341 163.367
R588 B.n343 B.n342 163.367
R589 B.n343 B.n204 163.367
R590 B.n347 B.n204 163.367
R591 B.n348 B.n347 163.367
R592 B.n349 B.n348 163.367
R593 B.n349 B.n202 163.367
R594 B.n353 B.n202 163.367
R595 B.n354 B.n353 163.367
R596 B.n355 B.n354 163.367
R597 B.n355 B.n200 163.367
R598 B.n359 B.n200 163.367
R599 B.n360 B.n359 163.367
R600 B.n361 B.n360 163.367
R601 B.n361 B.n198 163.367
R602 B.n365 B.n198 163.367
R603 B.n366 B.n365 163.367
R604 B.n367 B.n366 163.367
R605 B.n367 B.n196 163.367
R606 B.n371 B.n196 163.367
R607 B.n372 B.n371 163.367
R608 B.n373 B.n372 163.367
R609 B.n373 B.n194 163.367
R610 B.n377 B.n194 163.367
R611 B.n378 B.n377 163.367
R612 B.n379 B.n378 163.367
R613 B.n379 B.n192 163.367
R614 B.n383 B.n192 163.367
R615 B.n384 B.n383 163.367
R616 B.n385 B.n384 163.367
R617 B.n385 B.n190 163.367
R618 B.n389 B.n190 163.367
R619 B.n390 B.n389 163.367
R620 B.n391 B.n390 163.367
R621 B.n391 B.n188 163.367
R622 B.n395 B.n188 163.367
R623 B.n396 B.n395 163.367
R624 B.n397 B.n396 163.367
R625 B.n397 B.n186 163.367
R626 B.n401 B.n186 163.367
R627 B.n402 B.n401 163.367
R628 B.n402 B.n182 163.367
R629 B.n406 B.n182 163.367
R630 B.n407 B.n406 163.367
R631 B.n408 B.n407 163.367
R632 B.n408 B.n180 163.367
R633 B.n412 B.n180 163.367
R634 B.n413 B.n412 163.367
R635 B.n414 B.n413 163.367
R636 B.n414 B.n176 163.367
R637 B.n419 B.n176 163.367
R638 B.n420 B.n419 163.367
R639 B.n421 B.n420 163.367
R640 B.n421 B.n174 163.367
R641 B.n425 B.n174 163.367
R642 B.n426 B.n425 163.367
R643 B.n427 B.n426 163.367
R644 B.n427 B.n172 163.367
R645 B.n431 B.n172 163.367
R646 B.n432 B.n431 163.367
R647 B.n433 B.n432 163.367
R648 B.n433 B.n170 163.367
R649 B.n437 B.n170 163.367
R650 B.n438 B.n437 163.367
R651 B.n439 B.n438 163.367
R652 B.n439 B.n168 163.367
R653 B.n443 B.n168 163.367
R654 B.n444 B.n443 163.367
R655 B.n445 B.n444 163.367
R656 B.n445 B.n166 163.367
R657 B.n449 B.n166 163.367
R658 B.n450 B.n449 163.367
R659 B.n451 B.n450 163.367
R660 B.n451 B.n164 163.367
R661 B.n455 B.n164 163.367
R662 B.n456 B.n455 163.367
R663 B.n457 B.n456 163.367
R664 B.n457 B.n162 163.367
R665 B.n461 B.n162 163.367
R666 B.n462 B.n461 163.367
R667 B.n463 B.n462 163.367
R668 B.n463 B.n160 163.367
R669 B.n467 B.n160 163.367
R670 B.n468 B.n467 163.367
R671 B.n469 B.n468 163.367
R672 B.n469 B.n158 163.367
R673 B.n473 B.n158 163.367
R674 B.n474 B.n473 163.367
R675 B.n475 B.n474 163.367
R676 B.n475 B.n156 163.367
R677 B.n479 B.n156 163.367
R678 B.n480 B.n479 163.367
R679 B.n481 B.n480 163.367
R680 B.n481 B.n154 163.367
R681 B.n485 B.n154 163.367
R682 B.n486 B.n485 163.367
R683 B.n487 B.n486 163.367
R684 B.n487 B.n152 163.367
R685 B.n491 B.n152 163.367
R686 B.n492 B.n491 163.367
R687 B.n493 B.n492 163.367
R688 B.n493 B.n150 163.367
R689 B.n497 B.n150 163.367
R690 B.n498 B.n497 163.367
R691 B.n499 B.n498 163.367
R692 B.n499 B.n148 163.367
R693 B.n503 B.n148 163.367
R694 B.n504 B.n503 163.367
R695 B.n505 B.n504 163.367
R696 B.n505 B.n146 163.367
R697 B.n509 B.n146 163.367
R698 B.n510 B.n509 163.367
R699 B.n511 B.n510 163.367
R700 B.n511 B.n144 163.367
R701 B.n516 B.n515 163.367
R702 B.n517 B.n516 163.367
R703 B.n517 B.n142 163.367
R704 B.n521 B.n142 163.367
R705 B.n522 B.n521 163.367
R706 B.n523 B.n522 163.367
R707 B.n523 B.n140 163.367
R708 B.n527 B.n140 163.367
R709 B.n528 B.n527 163.367
R710 B.n529 B.n528 163.367
R711 B.n529 B.n138 163.367
R712 B.n533 B.n138 163.367
R713 B.n534 B.n533 163.367
R714 B.n535 B.n534 163.367
R715 B.n535 B.n136 163.367
R716 B.n539 B.n136 163.367
R717 B.n540 B.n539 163.367
R718 B.n541 B.n540 163.367
R719 B.n541 B.n134 163.367
R720 B.n545 B.n134 163.367
R721 B.n546 B.n545 163.367
R722 B.n547 B.n546 163.367
R723 B.n547 B.n132 163.367
R724 B.n551 B.n132 163.367
R725 B.n552 B.n551 163.367
R726 B.n553 B.n552 163.367
R727 B.n553 B.n130 163.367
R728 B.n557 B.n130 163.367
R729 B.n558 B.n557 163.367
R730 B.n559 B.n558 163.367
R731 B.n559 B.n128 163.367
R732 B.n563 B.n128 163.367
R733 B.n564 B.n563 163.367
R734 B.n565 B.n564 163.367
R735 B.n565 B.n126 163.367
R736 B.n569 B.n126 163.367
R737 B.n570 B.n569 163.367
R738 B.n571 B.n570 163.367
R739 B.n571 B.n124 163.367
R740 B.n575 B.n124 163.367
R741 B.n576 B.n575 163.367
R742 B.n577 B.n576 163.367
R743 B.n577 B.n122 163.367
R744 B.n581 B.n122 163.367
R745 B.n582 B.n581 163.367
R746 B.n583 B.n582 163.367
R747 B.n583 B.n120 163.367
R748 B.n587 B.n120 163.367
R749 B.n588 B.n587 163.367
R750 B.n589 B.n588 163.367
R751 B.n589 B.n118 163.367
R752 B.n593 B.n118 163.367
R753 B.n594 B.n593 163.367
R754 B.n595 B.n594 163.367
R755 B.n595 B.n116 163.367
R756 B.n599 B.n116 163.367
R757 B.n600 B.n599 163.367
R758 B.n601 B.n600 163.367
R759 B.n601 B.n114 163.367
R760 B.n605 B.n114 163.367
R761 B.n606 B.n605 163.367
R762 B.n607 B.n606 163.367
R763 B.n607 B.n112 163.367
R764 B.n611 B.n112 163.367
R765 B.n612 B.n611 163.367
R766 B.n613 B.n612 163.367
R767 B.n613 B.n110 163.367
R768 B.n617 B.n110 163.367
R769 B.n618 B.n617 163.367
R770 B.n619 B.n618 163.367
R771 B.n619 B.n108 163.367
R772 B.n623 B.n108 163.367
R773 B.n624 B.n623 163.367
R774 B.n625 B.n624 163.367
R775 B.n625 B.n106 163.367
R776 B.n629 B.n106 163.367
R777 B.n630 B.n629 163.367
R778 B.n631 B.n630 163.367
R779 B.n631 B.n104 163.367
R780 B.n635 B.n104 163.367
R781 B.n636 B.n635 163.367
R782 B.n637 B.n636 163.367
R783 B.n637 B.n102 163.367
R784 B.n641 B.n102 163.367
R785 B.n642 B.n641 163.367
R786 B.n643 B.n642 163.367
R787 B.n643 B.n100 163.367
R788 B.n647 B.n100 163.367
R789 B.n648 B.n647 163.367
R790 B.n649 B.n648 163.367
R791 B.n858 B.n25 163.367
R792 B.n854 B.n25 163.367
R793 B.n854 B.n853 163.367
R794 B.n853 B.n852 163.367
R795 B.n852 B.n27 163.367
R796 B.n848 B.n27 163.367
R797 B.n848 B.n847 163.367
R798 B.n847 B.n846 163.367
R799 B.n846 B.n29 163.367
R800 B.n842 B.n29 163.367
R801 B.n842 B.n841 163.367
R802 B.n841 B.n840 163.367
R803 B.n840 B.n31 163.367
R804 B.n836 B.n31 163.367
R805 B.n836 B.n835 163.367
R806 B.n835 B.n834 163.367
R807 B.n834 B.n33 163.367
R808 B.n830 B.n33 163.367
R809 B.n830 B.n829 163.367
R810 B.n829 B.n828 163.367
R811 B.n828 B.n35 163.367
R812 B.n824 B.n35 163.367
R813 B.n824 B.n823 163.367
R814 B.n823 B.n822 163.367
R815 B.n822 B.n37 163.367
R816 B.n818 B.n37 163.367
R817 B.n818 B.n817 163.367
R818 B.n817 B.n816 163.367
R819 B.n816 B.n39 163.367
R820 B.n812 B.n39 163.367
R821 B.n812 B.n811 163.367
R822 B.n811 B.n810 163.367
R823 B.n810 B.n41 163.367
R824 B.n806 B.n41 163.367
R825 B.n806 B.n805 163.367
R826 B.n805 B.n804 163.367
R827 B.n804 B.n43 163.367
R828 B.n800 B.n43 163.367
R829 B.n800 B.n799 163.367
R830 B.n799 B.n798 163.367
R831 B.n798 B.n45 163.367
R832 B.n794 B.n45 163.367
R833 B.n794 B.n793 163.367
R834 B.n793 B.n792 163.367
R835 B.n792 B.n47 163.367
R836 B.n788 B.n47 163.367
R837 B.n788 B.n787 163.367
R838 B.n787 B.n786 163.367
R839 B.n786 B.n49 163.367
R840 B.n782 B.n49 163.367
R841 B.n782 B.n781 163.367
R842 B.n781 B.n780 163.367
R843 B.n780 B.n51 163.367
R844 B.n776 B.n51 163.367
R845 B.n776 B.n775 163.367
R846 B.n775 B.n774 163.367
R847 B.n774 B.n53 163.367
R848 B.n770 B.n53 163.367
R849 B.n770 B.n769 163.367
R850 B.n769 B.n768 163.367
R851 B.n768 B.n55 163.367
R852 B.n764 B.n55 163.367
R853 B.n764 B.n763 163.367
R854 B.n763 B.n762 163.367
R855 B.n762 B.n57 163.367
R856 B.n758 B.n57 163.367
R857 B.n758 B.n757 163.367
R858 B.n757 B.n756 163.367
R859 B.n756 B.n62 163.367
R860 B.n752 B.n62 163.367
R861 B.n752 B.n751 163.367
R862 B.n751 B.n750 163.367
R863 B.n750 B.n64 163.367
R864 B.n745 B.n64 163.367
R865 B.n745 B.n744 163.367
R866 B.n744 B.n743 163.367
R867 B.n743 B.n68 163.367
R868 B.n739 B.n68 163.367
R869 B.n739 B.n738 163.367
R870 B.n738 B.n737 163.367
R871 B.n737 B.n70 163.367
R872 B.n733 B.n70 163.367
R873 B.n733 B.n732 163.367
R874 B.n732 B.n731 163.367
R875 B.n731 B.n72 163.367
R876 B.n727 B.n72 163.367
R877 B.n727 B.n726 163.367
R878 B.n726 B.n725 163.367
R879 B.n725 B.n74 163.367
R880 B.n721 B.n74 163.367
R881 B.n721 B.n720 163.367
R882 B.n720 B.n719 163.367
R883 B.n719 B.n76 163.367
R884 B.n715 B.n76 163.367
R885 B.n715 B.n714 163.367
R886 B.n714 B.n713 163.367
R887 B.n713 B.n78 163.367
R888 B.n709 B.n78 163.367
R889 B.n709 B.n708 163.367
R890 B.n708 B.n707 163.367
R891 B.n707 B.n80 163.367
R892 B.n703 B.n80 163.367
R893 B.n703 B.n702 163.367
R894 B.n702 B.n701 163.367
R895 B.n701 B.n82 163.367
R896 B.n697 B.n82 163.367
R897 B.n697 B.n696 163.367
R898 B.n696 B.n695 163.367
R899 B.n695 B.n84 163.367
R900 B.n691 B.n84 163.367
R901 B.n691 B.n690 163.367
R902 B.n690 B.n689 163.367
R903 B.n689 B.n86 163.367
R904 B.n685 B.n86 163.367
R905 B.n685 B.n684 163.367
R906 B.n684 B.n683 163.367
R907 B.n683 B.n88 163.367
R908 B.n679 B.n88 163.367
R909 B.n679 B.n678 163.367
R910 B.n678 B.n677 163.367
R911 B.n677 B.n90 163.367
R912 B.n673 B.n90 163.367
R913 B.n673 B.n672 163.367
R914 B.n672 B.n671 163.367
R915 B.n671 B.n92 163.367
R916 B.n667 B.n92 163.367
R917 B.n667 B.n666 163.367
R918 B.n666 B.n665 163.367
R919 B.n665 B.n94 163.367
R920 B.n661 B.n94 163.367
R921 B.n661 B.n660 163.367
R922 B.n660 B.n659 163.367
R923 B.n659 B.n96 163.367
R924 B.n655 B.n96 163.367
R925 B.n655 B.n654 163.367
R926 B.n654 B.n653 163.367
R927 B.n653 B.n98 163.367
R928 B.n417 B.n178 59.5399
R929 B.n185 B.n184 59.5399
R930 B.n60 B.n59 59.5399
R931 B.n747 B.n66 59.5399
R932 B.n178 B.n177 48.8732
R933 B.n184 B.n183 48.8732
R934 B.n59 B.n58 48.8732
R935 B.n66 B.n65 48.8732
R936 B.n857 B.n24 32.3127
R937 B.n651 B.n650 32.3127
R938 B.n514 B.n513 32.3127
R939 B.n304 B.n217 32.3127
R940 B B.n927 18.0485
R941 B.n857 B.n856 10.6151
R942 B.n856 B.n855 10.6151
R943 B.n855 B.n26 10.6151
R944 B.n851 B.n26 10.6151
R945 B.n851 B.n850 10.6151
R946 B.n850 B.n849 10.6151
R947 B.n849 B.n28 10.6151
R948 B.n845 B.n28 10.6151
R949 B.n845 B.n844 10.6151
R950 B.n844 B.n843 10.6151
R951 B.n843 B.n30 10.6151
R952 B.n839 B.n30 10.6151
R953 B.n839 B.n838 10.6151
R954 B.n838 B.n837 10.6151
R955 B.n837 B.n32 10.6151
R956 B.n833 B.n32 10.6151
R957 B.n833 B.n832 10.6151
R958 B.n832 B.n831 10.6151
R959 B.n831 B.n34 10.6151
R960 B.n827 B.n34 10.6151
R961 B.n827 B.n826 10.6151
R962 B.n826 B.n825 10.6151
R963 B.n825 B.n36 10.6151
R964 B.n821 B.n36 10.6151
R965 B.n821 B.n820 10.6151
R966 B.n820 B.n819 10.6151
R967 B.n819 B.n38 10.6151
R968 B.n815 B.n38 10.6151
R969 B.n815 B.n814 10.6151
R970 B.n814 B.n813 10.6151
R971 B.n813 B.n40 10.6151
R972 B.n809 B.n40 10.6151
R973 B.n809 B.n808 10.6151
R974 B.n808 B.n807 10.6151
R975 B.n807 B.n42 10.6151
R976 B.n803 B.n42 10.6151
R977 B.n803 B.n802 10.6151
R978 B.n802 B.n801 10.6151
R979 B.n801 B.n44 10.6151
R980 B.n797 B.n44 10.6151
R981 B.n797 B.n796 10.6151
R982 B.n796 B.n795 10.6151
R983 B.n795 B.n46 10.6151
R984 B.n791 B.n46 10.6151
R985 B.n791 B.n790 10.6151
R986 B.n790 B.n789 10.6151
R987 B.n789 B.n48 10.6151
R988 B.n785 B.n48 10.6151
R989 B.n785 B.n784 10.6151
R990 B.n784 B.n783 10.6151
R991 B.n783 B.n50 10.6151
R992 B.n779 B.n50 10.6151
R993 B.n779 B.n778 10.6151
R994 B.n778 B.n777 10.6151
R995 B.n777 B.n52 10.6151
R996 B.n773 B.n52 10.6151
R997 B.n773 B.n772 10.6151
R998 B.n772 B.n771 10.6151
R999 B.n771 B.n54 10.6151
R1000 B.n767 B.n54 10.6151
R1001 B.n767 B.n766 10.6151
R1002 B.n766 B.n765 10.6151
R1003 B.n765 B.n56 10.6151
R1004 B.n761 B.n760 10.6151
R1005 B.n760 B.n759 10.6151
R1006 B.n759 B.n61 10.6151
R1007 B.n755 B.n61 10.6151
R1008 B.n755 B.n754 10.6151
R1009 B.n754 B.n753 10.6151
R1010 B.n753 B.n63 10.6151
R1011 B.n749 B.n63 10.6151
R1012 B.n749 B.n748 10.6151
R1013 B.n746 B.n67 10.6151
R1014 B.n742 B.n67 10.6151
R1015 B.n742 B.n741 10.6151
R1016 B.n741 B.n740 10.6151
R1017 B.n740 B.n69 10.6151
R1018 B.n736 B.n69 10.6151
R1019 B.n736 B.n735 10.6151
R1020 B.n735 B.n734 10.6151
R1021 B.n734 B.n71 10.6151
R1022 B.n730 B.n71 10.6151
R1023 B.n730 B.n729 10.6151
R1024 B.n729 B.n728 10.6151
R1025 B.n728 B.n73 10.6151
R1026 B.n724 B.n73 10.6151
R1027 B.n724 B.n723 10.6151
R1028 B.n723 B.n722 10.6151
R1029 B.n722 B.n75 10.6151
R1030 B.n718 B.n75 10.6151
R1031 B.n718 B.n717 10.6151
R1032 B.n717 B.n716 10.6151
R1033 B.n716 B.n77 10.6151
R1034 B.n712 B.n77 10.6151
R1035 B.n712 B.n711 10.6151
R1036 B.n711 B.n710 10.6151
R1037 B.n710 B.n79 10.6151
R1038 B.n706 B.n79 10.6151
R1039 B.n706 B.n705 10.6151
R1040 B.n705 B.n704 10.6151
R1041 B.n704 B.n81 10.6151
R1042 B.n700 B.n81 10.6151
R1043 B.n700 B.n699 10.6151
R1044 B.n699 B.n698 10.6151
R1045 B.n698 B.n83 10.6151
R1046 B.n694 B.n83 10.6151
R1047 B.n694 B.n693 10.6151
R1048 B.n693 B.n692 10.6151
R1049 B.n692 B.n85 10.6151
R1050 B.n688 B.n85 10.6151
R1051 B.n688 B.n687 10.6151
R1052 B.n687 B.n686 10.6151
R1053 B.n686 B.n87 10.6151
R1054 B.n682 B.n87 10.6151
R1055 B.n682 B.n681 10.6151
R1056 B.n681 B.n680 10.6151
R1057 B.n680 B.n89 10.6151
R1058 B.n676 B.n89 10.6151
R1059 B.n676 B.n675 10.6151
R1060 B.n675 B.n674 10.6151
R1061 B.n674 B.n91 10.6151
R1062 B.n670 B.n91 10.6151
R1063 B.n670 B.n669 10.6151
R1064 B.n669 B.n668 10.6151
R1065 B.n668 B.n93 10.6151
R1066 B.n664 B.n93 10.6151
R1067 B.n664 B.n663 10.6151
R1068 B.n663 B.n662 10.6151
R1069 B.n662 B.n95 10.6151
R1070 B.n658 B.n95 10.6151
R1071 B.n658 B.n657 10.6151
R1072 B.n657 B.n656 10.6151
R1073 B.n656 B.n97 10.6151
R1074 B.n652 B.n97 10.6151
R1075 B.n652 B.n651 10.6151
R1076 B.n514 B.n143 10.6151
R1077 B.n518 B.n143 10.6151
R1078 B.n519 B.n518 10.6151
R1079 B.n520 B.n519 10.6151
R1080 B.n520 B.n141 10.6151
R1081 B.n524 B.n141 10.6151
R1082 B.n525 B.n524 10.6151
R1083 B.n526 B.n525 10.6151
R1084 B.n526 B.n139 10.6151
R1085 B.n530 B.n139 10.6151
R1086 B.n531 B.n530 10.6151
R1087 B.n532 B.n531 10.6151
R1088 B.n532 B.n137 10.6151
R1089 B.n536 B.n137 10.6151
R1090 B.n537 B.n536 10.6151
R1091 B.n538 B.n537 10.6151
R1092 B.n538 B.n135 10.6151
R1093 B.n542 B.n135 10.6151
R1094 B.n543 B.n542 10.6151
R1095 B.n544 B.n543 10.6151
R1096 B.n544 B.n133 10.6151
R1097 B.n548 B.n133 10.6151
R1098 B.n549 B.n548 10.6151
R1099 B.n550 B.n549 10.6151
R1100 B.n550 B.n131 10.6151
R1101 B.n554 B.n131 10.6151
R1102 B.n555 B.n554 10.6151
R1103 B.n556 B.n555 10.6151
R1104 B.n556 B.n129 10.6151
R1105 B.n560 B.n129 10.6151
R1106 B.n561 B.n560 10.6151
R1107 B.n562 B.n561 10.6151
R1108 B.n562 B.n127 10.6151
R1109 B.n566 B.n127 10.6151
R1110 B.n567 B.n566 10.6151
R1111 B.n568 B.n567 10.6151
R1112 B.n568 B.n125 10.6151
R1113 B.n572 B.n125 10.6151
R1114 B.n573 B.n572 10.6151
R1115 B.n574 B.n573 10.6151
R1116 B.n574 B.n123 10.6151
R1117 B.n578 B.n123 10.6151
R1118 B.n579 B.n578 10.6151
R1119 B.n580 B.n579 10.6151
R1120 B.n580 B.n121 10.6151
R1121 B.n584 B.n121 10.6151
R1122 B.n585 B.n584 10.6151
R1123 B.n586 B.n585 10.6151
R1124 B.n586 B.n119 10.6151
R1125 B.n590 B.n119 10.6151
R1126 B.n591 B.n590 10.6151
R1127 B.n592 B.n591 10.6151
R1128 B.n592 B.n117 10.6151
R1129 B.n596 B.n117 10.6151
R1130 B.n597 B.n596 10.6151
R1131 B.n598 B.n597 10.6151
R1132 B.n598 B.n115 10.6151
R1133 B.n602 B.n115 10.6151
R1134 B.n603 B.n602 10.6151
R1135 B.n604 B.n603 10.6151
R1136 B.n604 B.n113 10.6151
R1137 B.n608 B.n113 10.6151
R1138 B.n609 B.n608 10.6151
R1139 B.n610 B.n609 10.6151
R1140 B.n610 B.n111 10.6151
R1141 B.n614 B.n111 10.6151
R1142 B.n615 B.n614 10.6151
R1143 B.n616 B.n615 10.6151
R1144 B.n616 B.n109 10.6151
R1145 B.n620 B.n109 10.6151
R1146 B.n621 B.n620 10.6151
R1147 B.n622 B.n621 10.6151
R1148 B.n622 B.n107 10.6151
R1149 B.n626 B.n107 10.6151
R1150 B.n627 B.n626 10.6151
R1151 B.n628 B.n627 10.6151
R1152 B.n628 B.n105 10.6151
R1153 B.n632 B.n105 10.6151
R1154 B.n633 B.n632 10.6151
R1155 B.n634 B.n633 10.6151
R1156 B.n634 B.n103 10.6151
R1157 B.n638 B.n103 10.6151
R1158 B.n639 B.n638 10.6151
R1159 B.n640 B.n639 10.6151
R1160 B.n640 B.n101 10.6151
R1161 B.n644 B.n101 10.6151
R1162 B.n645 B.n644 10.6151
R1163 B.n646 B.n645 10.6151
R1164 B.n646 B.n99 10.6151
R1165 B.n650 B.n99 10.6151
R1166 B.n308 B.n217 10.6151
R1167 B.n309 B.n308 10.6151
R1168 B.n310 B.n309 10.6151
R1169 B.n310 B.n215 10.6151
R1170 B.n314 B.n215 10.6151
R1171 B.n315 B.n314 10.6151
R1172 B.n316 B.n315 10.6151
R1173 B.n316 B.n213 10.6151
R1174 B.n320 B.n213 10.6151
R1175 B.n321 B.n320 10.6151
R1176 B.n322 B.n321 10.6151
R1177 B.n322 B.n211 10.6151
R1178 B.n326 B.n211 10.6151
R1179 B.n327 B.n326 10.6151
R1180 B.n328 B.n327 10.6151
R1181 B.n328 B.n209 10.6151
R1182 B.n332 B.n209 10.6151
R1183 B.n333 B.n332 10.6151
R1184 B.n334 B.n333 10.6151
R1185 B.n334 B.n207 10.6151
R1186 B.n338 B.n207 10.6151
R1187 B.n339 B.n338 10.6151
R1188 B.n340 B.n339 10.6151
R1189 B.n340 B.n205 10.6151
R1190 B.n344 B.n205 10.6151
R1191 B.n345 B.n344 10.6151
R1192 B.n346 B.n345 10.6151
R1193 B.n346 B.n203 10.6151
R1194 B.n350 B.n203 10.6151
R1195 B.n351 B.n350 10.6151
R1196 B.n352 B.n351 10.6151
R1197 B.n352 B.n201 10.6151
R1198 B.n356 B.n201 10.6151
R1199 B.n357 B.n356 10.6151
R1200 B.n358 B.n357 10.6151
R1201 B.n358 B.n199 10.6151
R1202 B.n362 B.n199 10.6151
R1203 B.n363 B.n362 10.6151
R1204 B.n364 B.n363 10.6151
R1205 B.n364 B.n197 10.6151
R1206 B.n368 B.n197 10.6151
R1207 B.n369 B.n368 10.6151
R1208 B.n370 B.n369 10.6151
R1209 B.n370 B.n195 10.6151
R1210 B.n374 B.n195 10.6151
R1211 B.n375 B.n374 10.6151
R1212 B.n376 B.n375 10.6151
R1213 B.n376 B.n193 10.6151
R1214 B.n380 B.n193 10.6151
R1215 B.n381 B.n380 10.6151
R1216 B.n382 B.n381 10.6151
R1217 B.n382 B.n191 10.6151
R1218 B.n386 B.n191 10.6151
R1219 B.n387 B.n386 10.6151
R1220 B.n388 B.n387 10.6151
R1221 B.n388 B.n189 10.6151
R1222 B.n392 B.n189 10.6151
R1223 B.n393 B.n392 10.6151
R1224 B.n394 B.n393 10.6151
R1225 B.n394 B.n187 10.6151
R1226 B.n398 B.n187 10.6151
R1227 B.n399 B.n398 10.6151
R1228 B.n400 B.n399 10.6151
R1229 B.n404 B.n403 10.6151
R1230 B.n405 B.n404 10.6151
R1231 B.n405 B.n181 10.6151
R1232 B.n409 B.n181 10.6151
R1233 B.n410 B.n409 10.6151
R1234 B.n411 B.n410 10.6151
R1235 B.n411 B.n179 10.6151
R1236 B.n415 B.n179 10.6151
R1237 B.n416 B.n415 10.6151
R1238 B.n418 B.n175 10.6151
R1239 B.n422 B.n175 10.6151
R1240 B.n423 B.n422 10.6151
R1241 B.n424 B.n423 10.6151
R1242 B.n424 B.n173 10.6151
R1243 B.n428 B.n173 10.6151
R1244 B.n429 B.n428 10.6151
R1245 B.n430 B.n429 10.6151
R1246 B.n430 B.n171 10.6151
R1247 B.n434 B.n171 10.6151
R1248 B.n435 B.n434 10.6151
R1249 B.n436 B.n435 10.6151
R1250 B.n436 B.n169 10.6151
R1251 B.n440 B.n169 10.6151
R1252 B.n441 B.n440 10.6151
R1253 B.n442 B.n441 10.6151
R1254 B.n442 B.n167 10.6151
R1255 B.n446 B.n167 10.6151
R1256 B.n447 B.n446 10.6151
R1257 B.n448 B.n447 10.6151
R1258 B.n448 B.n165 10.6151
R1259 B.n452 B.n165 10.6151
R1260 B.n453 B.n452 10.6151
R1261 B.n454 B.n453 10.6151
R1262 B.n454 B.n163 10.6151
R1263 B.n458 B.n163 10.6151
R1264 B.n459 B.n458 10.6151
R1265 B.n460 B.n459 10.6151
R1266 B.n460 B.n161 10.6151
R1267 B.n464 B.n161 10.6151
R1268 B.n465 B.n464 10.6151
R1269 B.n466 B.n465 10.6151
R1270 B.n466 B.n159 10.6151
R1271 B.n470 B.n159 10.6151
R1272 B.n471 B.n470 10.6151
R1273 B.n472 B.n471 10.6151
R1274 B.n472 B.n157 10.6151
R1275 B.n476 B.n157 10.6151
R1276 B.n477 B.n476 10.6151
R1277 B.n478 B.n477 10.6151
R1278 B.n478 B.n155 10.6151
R1279 B.n482 B.n155 10.6151
R1280 B.n483 B.n482 10.6151
R1281 B.n484 B.n483 10.6151
R1282 B.n484 B.n153 10.6151
R1283 B.n488 B.n153 10.6151
R1284 B.n489 B.n488 10.6151
R1285 B.n490 B.n489 10.6151
R1286 B.n490 B.n151 10.6151
R1287 B.n494 B.n151 10.6151
R1288 B.n495 B.n494 10.6151
R1289 B.n496 B.n495 10.6151
R1290 B.n496 B.n149 10.6151
R1291 B.n500 B.n149 10.6151
R1292 B.n501 B.n500 10.6151
R1293 B.n502 B.n501 10.6151
R1294 B.n502 B.n147 10.6151
R1295 B.n506 B.n147 10.6151
R1296 B.n507 B.n506 10.6151
R1297 B.n508 B.n507 10.6151
R1298 B.n508 B.n145 10.6151
R1299 B.n512 B.n145 10.6151
R1300 B.n513 B.n512 10.6151
R1301 B.n304 B.n303 10.6151
R1302 B.n303 B.n302 10.6151
R1303 B.n302 B.n219 10.6151
R1304 B.n298 B.n219 10.6151
R1305 B.n298 B.n297 10.6151
R1306 B.n297 B.n296 10.6151
R1307 B.n296 B.n221 10.6151
R1308 B.n292 B.n221 10.6151
R1309 B.n292 B.n291 10.6151
R1310 B.n291 B.n290 10.6151
R1311 B.n290 B.n223 10.6151
R1312 B.n286 B.n223 10.6151
R1313 B.n286 B.n285 10.6151
R1314 B.n285 B.n284 10.6151
R1315 B.n284 B.n225 10.6151
R1316 B.n280 B.n225 10.6151
R1317 B.n280 B.n279 10.6151
R1318 B.n279 B.n278 10.6151
R1319 B.n278 B.n227 10.6151
R1320 B.n274 B.n227 10.6151
R1321 B.n274 B.n273 10.6151
R1322 B.n273 B.n272 10.6151
R1323 B.n272 B.n229 10.6151
R1324 B.n268 B.n229 10.6151
R1325 B.n268 B.n267 10.6151
R1326 B.n267 B.n266 10.6151
R1327 B.n266 B.n231 10.6151
R1328 B.n262 B.n231 10.6151
R1329 B.n262 B.n261 10.6151
R1330 B.n261 B.n260 10.6151
R1331 B.n260 B.n233 10.6151
R1332 B.n256 B.n233 10.6151
R1333 B.n256 B.n255 10.6151
R1334 B.n255 B.n254 10.6151
R1335 B.n254 B.n235 10.6151
R1336 B.n250 B.n235 10.6151
R1337 B.n250 B.n249 10.6151
R1338 B.n249 B.n248 10.6151
R1339 B.n248 B.n237 10.6151
R1340 B.n244 B.n237 10.6151
R1341 B.n244 B.n243 10.6151
R1342 B.n243 B.n242 10.6151
R1343 B.n242 B.n239 10.6151
R1344 B.n239 B.n0 10.6151
R1345 B.n923 B.n1 10.6151
R1346 B.n923 B.n922 10.6151
R1347 B.n922 B.n921 10.6151
R1348 B.n921 B.n4 10.6151
R1349 B.n917 B.n4 10.6151
R1350 B.n917 B.n916 10.6151
R1351 B.n916 B.n915 10.6151
R1352 B.n915 B.n6 10.6151
R1353 B.n911 B.n6 10.6151
R1354 B.n911 B.n910 10.6151
R1355 B.n910 B.n909 10.6151
R1356 B.n909 B.n8 10.6151
R1357 B.n905 B.n8 10.6151
R1358 B.n905 B.n904 10.6151
R1359 B.n904 B.n903 10.6151
R1360 B.n903 B.n10 10.6151
R1361 B.n899 B.n10 10.6151
R1362 B.n899 B.n898 10.6151
R1363 B.n898 B.n897 10.6151
R1364 B.n897 B.n12 10.6151
R1365 B.n893 B.n12 10.6151
R1366 B.n893 B.n892 10.6151
R1367 B.n892 B.n891 10.6151
R1368 B.n891 B.n14 10.6151
R1369 B.n887 B.n14 10.6151
R1370 B.n887 B.n886 10.6151
R1371 B.n886 B.n885 10.6151
R1372 B.n885 B.n16 10.6151
R1373 B.n881 B.n16 10.6151
R1374 B.n881 B.n880 10.6151
R1375 B.n880 B.n879 10.6151
R1376 B.n879 B.n18 10.6151
R1377 B.n875 B.n18 10.6151
R1378 B.n875 B.n874 10.6151
R1379 B.n874 B.n873 10.6151
R1380 B.n873 B.n20 10.6151
R1381 B.n869 B.n20 10.6151
R1382 B.n869 B.n868 10.6151
R1383 B.n868 B.n867 10.6151
R1384 B.n867 B.n22 10.6151
R1385 B.n863 B.n22 10.6151
R1386 B.n863 B.n862 10.6151
R1387 B.n862 B.n861 10.6151
R1388 B.n861 B.n24 10.6151
R1389 B.n60 B.n56 9.36635
R1390 B.n747 B.n746 9.36635
R1391 B.n400 B.n185 9.36635
R1392 B.n418 B.n417 9.36635
R1393 B.n927 B.n0 2.81026
R1394 B.n927 B.n1 2.81026
R1395 B.n761 B.n60 1.24928
R1396 B.n748 B.n747 1.24928
R1397 B.n403 B.n185 1.24928
R1398 B.n417 B.n416 1.24928
R1399 VP.n14 VP.t5 248.438
R1400 VP.n34 VP.t4 215.911
R1401 VP.n5 VP.t2 215.911
R1402 VP.n51 VP.t3 215.911
R1403 VP.n59 VP.t7 215.911
R1404 VP.n31 VP.t0 215.911
R1405 VP.n23 VP.t1 215.911
R1406 VP.n13 VP.t6 215.911
R1407 VP.n16 VP.n15 161.3
R1408 VP.n17 VP.n12 161.3
R1409 VP.n19 VP.n18 161.3
R1410 VP.n20 VP.n11 161.3
R1411 VP.n22 VP.n21 161.3
R1412 VP.n24 VP.n10 161.3
R1413 VP.n26 VP.n25 161.3
R1414 VP.n27 VP.n9 161.3
R1415 VP.n29 VP.n28 161.3
R1416 VP.n30 VP.n8 161.3
R1417 VP.n58 VP.n0 161.3
R1418 VP.n57 VP.n56 161.3
R1419 VP.n55 VP.n1 161.3
R1420 VP.n54 VP.n53 161.3
R1421 VP.n52 VP.n2 161.3
R1422 VP.n50 VP.n49 161.3
R1423 VP.n48 VP.n3 161.3
R1424 VP.n47 VP.n46 161.3
R1425 VP.n45 VP.n4 161.3
R1426 VP.n44 VP.n43 161.3
R1427 VP.n42 VP.n41 161.3
R1428 VP.n40 VP.n6 161.3
R1429 VP.n39 VP.n38 161.3
R1430 VP.n37 VP.n7 161.3
R1431 VP.n36 VP.n35 161.3
R1432 VP.n34 VP.n33 97.1368
R1433 VP.n60 VP.n59 97.1368
R1434 VP.n32 VP.n31 97.1368
R1435 VP.n14 VP.n13 58.8804
R1436 VP.n33 VP.n32 54.7269
R1437 VP.n39 VP.n7 42.5146
R1438 VP.n57 VP.n1 42.5146
R1439 VP.n29 VP.n9 42.5146
R1440 VP.n46 VP.n45 40.577
R1441 VP.n46 VP.n3 40.577
R1442 VP.n18 VP.n11 40.577
R1443 VP.n18 VP.n17 40.577
R1444 VP.n40 VP.n39 38.6395
R1445 VP.n53 VP.n1 38.6395
R1446 VP.n25 VP.n9 38.6395
R1447 VP.n35 VP.n7 24.5923
R1448 VP.n41 VP.n40 24.5923
R1449 VP.n45 VP.n44 24.5923
R1450 VP.n50 VP.n3 24.5923
R1451 VP.n53 VP.n52 24.5923
R1452 VP.n58 VP.n57 24.5923
R1453 VP.n30 VP.n29 24.5923
R1454 VP.n22 VP.n11 24.5923
R1455 VP.n25 VP.n24 24.5923
R1456 VP.n17 VP.n16 24.5923
R1457 VP.n35 VP.n34 13.7719
R1458 VP.n59 VP.n58 13.7719
R1459 VP.n31 VP.n30 13.7719
R1460 VP.n44 VP.n5 12.7883
R1461 VP.n51 VP.n50 12.7883
R1462 VP.n23 VP.n22 12.7883
R1463 VP.n16 VP.n13 12.7883
R1464 VP.n41 VP.n5 11.8046
R1465 VP.n52 VP.n51 11.8046
R1466 VP.n24 VP.n23 11.8046
R1467 VP.n15 VP.n14 9.55925
R1468 VP.n32 VP.n8 0.278335
R1469 VP.n36 VP.n33 0.278335
R1470 VP.n60 VP.n0 0.278335
R1471 VP.n15 VP.n12 0.189894
R1472 VP.n19 VP.n12 0.189894
R1473 VP.n20 VP.n19 0.189894
R1474 VP.n21 VP.n20 0.189894
R1475 VP.n21 VP.n10 0.189894
R1476 VP.n26 VP.n10 0.189894
R1477 VP.n27 VP.n26 0.189894
R1478 VP.n28 VP.n27 0.189894
R1479 VP.n28 VP.n8 0.189894
R1480 VP.n37 VP.n36 0.189894
R1481 VP.n38 VP.n37 0.189894
R1482 VP.n38 VP.n6 0.189894
R1483 VP.n42 VP.n6 0.189894
R1484 VP.n43 VP.n42 0.189894
R1485 VP.n43 VP.n4 0.189894
R1486 VP.n47 VP.n4 0.189894
R1487 VP.n48 VP.n47 0.189894
R1488 VP.n49 VP.n48 0.189894
R1489 VP.n49 VP.n2 0.189894
R1490 VP.n54 VP.n2 0.189894
R1491 VP.n55 VP.n54 0.189894
R1492 VP.n56 VP.n55 0.189894
R1493 VP.n56 VP.n0 0.189894
R1494 VP VP.n60 0.153485
R1495 VTAIL.n882 VTAIL.n778 756.745
R1496 VTAIL.n106 VTAIL.n2 756.745
R1497 VTAIL.n216 VTAIL.n112 756.745
R1498 VTAIL.n328 VTAIL.n224 756.745
R1499 VTAIL.n772 VTAIL.n668 756.745
R1500 VTAIL.n660 VTAIL.n556 756.745
R1501 VTAIL.n550 VTAIL.n446 756.745
R1502 VTAIL.n438 VTAIL.n334 756.745
R1503 VTAIL.n815 VTAIL.n814 585
R1504 VTAIL.n817 VTAIL.n816 585
R1505 VTAIL.n810 VTAIL.n809 585
R1506 VTAIL.n823 VTAIL.n822 585
R1507 VTAIL.n825 VTAIL.n824 585
R1508 VTAIL.n806 VTAIL.n805 585
R1509 VTAIL.n831 VTAIL.n830 585
R1510 VTAIL.n833 VTAIL.n832 585
R1511 VTAIL.n802 VTAIL.n801 585
R1512 VTAIL.n839 VTAIL.n838 585
R1513 VTAIL.n841 VTAIL.n840 585
R1514 VTAIL.n798 VTAIL.n797 585
R1515 VTAIL.n847 VTAIL.n846 585
R1516 VTAIL.n849 VTAIL.n848 585
R1517 VTAIL.n794 VTAIL.n793 585
R1518 VTAIL.n856 VTAIL.n855 585
R1519 VTAIL.n857 VTAIL.n792 585
R1520 VTAIL.n859 VTAIL.n858 585
R1521 VTAIL.n790 VTAIL.n789 585
R1522 VTAIL.n865 VTAIL.n864 585
R1523 VTAIL.n867 VTAIL.n866 585
R1524 VTAIL.n786 VTAIL.n785 585
R1525 VTAIL.n873 VTAIL.n872 585
R1526 VTAIL.n875 VTAIL.n874 585
R1527 VTAIL.n782 VTAIL.n781 585
R1528 VTAIL.n881 VTAIL.n880 585
R1529 VTAIL.n883 VTAIL.n882 585
R1530 VTAIL.n39 VTAIL.n38 585
R1531 VTAIL.n41 VTAIL.n40 585
R1532 VTAIL.n34 VTAIL.n33 585
R1533 VTAIL.n47 VTAIL.n46 585
R1534 VTAIL.n49 VTAIL.n48 585
R1535 VTAIL.n30 VTAIL.n29 585
R1536 VTAIL.n55 VTAIL.n54 585
R1537 VTAIL.n57 VTAIL.n56 585
R1538 VTAIL.n26 VTAIL.n25 585
R1539 VTAIL.n63 VTAIL.n62 585
R1540 VTAIL.n65 VTAIL.n64 585
R1541 VTAIL.n22 VTAIL.n21 585
R1542 VTAIL.n71 VTAIL.n70 585
R1543 VTAIL.n73 VTAIL.n72 585
R1544 VTAIL.n18 VTAIL.n17 585
R1545 VTAIL.n80 VTAIL.n79 585
R1546 VTAIL.n81 VTAIL.n16 585
R1547 VTAIL.n83 VTAIL.n82 585
R1548 VTAIL.n14 VTAIL.n13 585
R1549 VTAIL.n89 VTAIL.n88 585
R1550 VTAIL.n91 VTAIL.n90 585
R1551 VTAIL.n10 VTAIL.n9 585
R1552 VTAIL.n97 VTAIL.n96 585
R1553 VTAIL.n99 VTAIL.n98 585
R1554 VTAIL.n6 VTAIL.n5 585
R1555 VTAIL.n105 VTAIL.n104 585
R1556 VTAIL.n107 VTAIL.n106 585
R1557 VTAIL.n149 VTAIL.n148 585
R1558 VTAIL.n151 VTAIL.n150 585
R1559 VTAIL.n144 VTAIL.n143 585
R1560 VTAIL.n157 VTAIL.n156 585
R1561 VTAIL.n159 VTAIL.n158 585
R1562 VTAIL.n140 VTAIL.n139 585
R1563 VTAIL.n165 VTAIL.n164 585
R1564 VTAIL.n167 VTAIL.n166 585
R1565 VTAIL.n136 VTAIL.n135 585
R1566 VTAIL.n173 VTAIL.n172 585
R1567 VTAIL.n175 VTAIL.n174 585
R1568 VTAIL.n132 VTAIL.n131 585
R1569 VTAIL.n181 VTAIL.n180 585
R1570 VTAIL.n183 VTAIL.n182 585
R1571 VTAIL.n128 VTAIL.n127 585
R1572 VTAIL.n190 VTAIL.n189 585
R1573 VTAIL.n191 VTAIL.n126 585
R1574 VTAIL.n193 VTAIL.n192 585
R1575 VTAIL.n124 VTAIL.n123 585
R1576 VTAIL.n199 VTAIL.n198 585
R1577 VTAIL.n201 VTAIL.n200 585
R1578 VTAIL.n120 VTAIL.n119 585
R1579 VTAIL.n207 VTAIL.n206 585
R1580 VTAIL.n209 VTAIL.n208 585
R1581 VTAIL.n116 VTAIL.n115 585
R1582 VTAIL.n215 VTAIL.n214 585
R1583 VTAIL.n217 VTAIL.n216 585
R1584 VTAIL.n261 VTAIL.n260 585
R1585 VTAIL.n263 VTAIL.n262 585
R1586 VTAIL.n256 VTAIL.n255 585
R1587 VTAIL.n269 VTAIL.n268 585
R1588 VTAIL.n271 VTAIL.n270 585
R1589 VTAIL.n252 VTAIL.n251 585
R1590 VTAIL.n277 VTAIL.n276 585
R1591 VTAIL.n279 VTAIL.n278 585
R1592 VTAIL.n248 VTAIL.n247 585
R1593 VTAIL.n285 VTAIL.n284 585
R1594 VTAIL.n287 VTAIL.n286 585
R1595 VTAIL.n244 VTAIL.n243 585
R1596 VTAIL.n293 VTAIL.n292 585
R1597 VTAIL.n295 VTAIL.n294 585
R1598 VTAIL.n240 VTAIL.n239 585
R1599 VTAIL.n302 VTAIL.n301 585
R1600 VTAIL.n303 VTAIL.n238 585
R1601 VTAIL.n305 VTAIL.n304 585
R1602 VTAIL.n236 VTAIL.n235 585
R1603 VTAIL.n311 VTAIL.n310 585
R1604 VTAIL.n313 VTAIL.n312 585
R1605 VTAIL.n232 VTAIL.n231 585
R1606 VTAIL.n319 VTAIL.n318 585
R1607 VTAIL.n321 VTAIL.n320 585
R1608 VTAIL.n228 VTAIL.n227 585
R1609 VTAIL.n327 VTAIL.n326 585
R1610 VTAIL.n329 VTAIL.n328 585
R1611 VTAIL.n773 VTAIL.n772 585
R1612 VTAIL.n771 VTAIL.n770 585
R1613 VTAIL.n672 VTAIL.n671 585
R1614 VTAIL.n765 VTAIL.n764 585
R1615 VTAIL.n763 VTAIL.n762 585
R1616 VTAIL.n676 VTAIL.n675 585
R1617 VTAIL.n757 VTAIL.n756 585
R1618 VTAIL.n755 VTAIL.n754 585
R1619 VTAIL.n680 VTAIL.n679 585
R1620 VTAIL.n684 VTAIL.n682 585
R1621 VTAIL.n749 VTAIL.n748 585
R1622 VTAIL.n747 VTAIL.n746 585
R1623 VTAIL.n686 VTAIL.n685 585
R1624 VTAIL.n741 VTAIL.n740 585
R1625 VTAIL.n739 VTAIL.n738 585
R1626 VTAIL.n690 VTAIL.n689 585
R1627 VTAIL.n733 VTAIL.n732 585
R1628 VTAIL.n731 VTAIL.n730 585
R1629 VTAIL.n694 VTAIL.n693 585
R1630 VTAIL.n725 VTAIL.n724 585
R1631 VTAIL.n723 VTAIL.n722 585
R1632 VTAIL.n698 VTAIL.n697 585
R1633 VTAIL.n717 VTAIL.n716 585
R1634 VTAIL.n715 VTAIL.n714 585
R1635 VTAIL.n702 VTAIL.n701 585
R1636 VTAIL.n709 VTAIL.n708 585
R1637 VTAIL.n707 VTAIL.n706 585
R1638 VTAIL.n661 VTAIL.n660 585
R1639 VTAIL.n659 VTAIL.n658 585
R1640 VTAIL.n560 VTAIL.n559 585
R1641 VTAIL.n653 VTAIL.n652 585
R1642 VTAIL.n651 VTAIL.n650 585
R1643 VTAIL.n564 VTAIL.n563 585
R1644 VTAIL.n645 VTAIL.n644 585
R1645 VTAIL.n643 VTAIL.n642 585
R1646 VTAIL.n568 VTAIL.n567 585
R1647 VTAIL.n572 VTAIL.n570 585
R1648 VTAIL.n637 VTAIL.n636 585
R1649 VTAIL.n635 VTAIL.n634 585
R1650 VTAIL.n574 VTAIL.n573 585
R1651 VTAIL.n629 VTAIL.n628 585
R1652 VTAIL.n627 VTAIL.n626 585
R1653 VTAIL.n578 VTAIL.n577 585
R1654 VTAIL.n621 VTAIL.n620 585
R1655 VTAIL.n619 VTAIL.n618 585
R1656 VTAIL.n582 VTAIL.n581 585
R1657 VTAIL.n613 VTAIL.n612 585
R1658 VTAIL.n611 VTAIL.n610 585
R1659 VTAIL.n586 VTAIL.n585 585
R1660 VTAIL.n605 VTAIL.n604 585
R1661 VTAIL.n603 VTAIL.n602 585
R1662 VTAIL.n590 VTAIL.n589 585
R1663 VTAIL.n597 VTAIL.n596 585
R1664 VTAIL.n595 VTAIL.n594 585
R1665 VTAIL.n551 VTAIL.n550 585
R1666 VTAIL.n549 VTAIL.n548 585
R1667 VTAIL.n450 VTAIL.n449 585
R1668 VTAIL.n543 VTAIL.n542 585
R1669 VTAIL.n541 VTAIL.n540 585
R1670 VTAIL.n454 VTAIL.n453 585
R1671 VTAIL.n535 VTAIL.n534 585
R1672 VTAIL.n533 VTAIL.n532 585
R1673 VTAIL.n458 VTAIL.n457 585
R1674 VTAIL.n462 VTAIL.n460 585
R1675 VTAIL.n527 VTAIL.n526 585
R1676 VTAIL.n525 VTAIL.n524 585
R1677 VTAIL.n464 VTAIL.n463 585
R1678 VTAIL.n519 VTAIL.n518 585
R1679 VTAIL.n517 VTAIL.n516 585
R1680 VTAIL.n468 VTAIL.n467 585
R1681 VTAIL.n511 VTAIL.n510 585
R1682 VTAIL.n509 VTAIL.n508 585
R1683 VTAIL.n472 VTAIL.n471 585
R1684 VTAIL.n503 VTAIL.n502 585
R1685 VTAIL.n501 VTAIL.n500 585
R1686 VTAIL.n476 VTAIL.n475 585
R1687 VTAIL.n495 VTAIL.n494 585
R1688 VTAIL.n493 VTAIL.n492 585
R1689 VTAIL.n480 VTAIL.n479 585
R1690 VTAIL.n487 VTAIL.n486 585
R1691 VTAIL.n485 VTAIL.n484 585
R1692 VTAIL.n439 VTAIL.n438 585
R1693 VTAIL.n437 VTAIL.n436 585
R1694 VTAIL.n338 VTAIL.n337 585
R1695 VTAIL.n431 VTAIL.n430 585
R1696 VTAIL.n429 VTAIL.n428 585
R1697 VTAIL.n342 VTAIL.n341 585
R1698 VTAIL.n423 VTAIL.n422 585
R1699 VTAIL.n421 VTAIL.n420 585
R1700 VTAIL.n346 VTAIL.n345 585
R1701 VTAIL.n350 VTAIL.n348 585
R1702 VTAIL.n415 VTAIL.n414 585
R1703 VTAIL.n413 VTAIL.n412 585
R1704 VTAIL.n352 VTAIL.n351 585
R1705 VTAIL.n407 VTAIL.n406 585
R1706 VTAIL.n405 VTAIL.n404 585
R1707 VTAIL.n356 VTAIL.n355 585
R1708 VTAIL.n399 VTAIL.n398 585
R1709 VTAIL.n397 VTAIL.n396 585
R1710 VTAIL.n360 VTAIL.n359 585
R1711 VTAIL.n391 VTAIL.n390 585
R1712 VTAIL.n389 VTAIL.n388 585
R1713 VTAIL.n364 VTAIL.n363 585
R1714 VTAIL.n383 VTAIL.n382 585
R1715 VTAIL.n381 VTAIL.n380 585
R1716 VTAIL.n368 VTAIL.n367 585
R1717 VTAIL.n375 VTAIL.n374 585
R1718 VTAIL.n373 VTAIL.n372 585
R1719 VTAIL.n813 VTAIL.t0 327.466
R1720 VTAIL.n37 VTAIL.t7 327.466
R1721 VTAIL.n147 VTAIL.t11 327.466
R1722 VTAIL.n259 VTAIL.t15 327.466
R1723 VTAIL.n705 VTAIL.t9 327.466
R1724 VTAIL.n593 VTAIL.t8 327.466
R1725 VTAIL.n483 VTAIL.t6 327.466
R1726 VTAIL.n371 VTAIL.t2 327.466
R1727 VTAIL.n816 VTAIL.n815 171.744
R1728 VTAIL.n816 VTAIL.n809 171.744
R1729 VTAIL.n823 VTAIL.n809 171.744
R1730 VTAIL.n824 VTAIL.n823 171.744
R1731 VTAIL.n824 VTAIL.n805 171.744
R1732 VTAIL.n831 VTAIL.n805 171.744
R1733 VTAIL.n832 VTAIL.n831 171.744
R1734 VTAIL.n832 VTAIL.n801 171.744
R1735 VTAIL.n839 VTAIL.n801 171.744
R1736 VTAIL.n840 VTAIL.n839 171.744
R1737 VTAIL.n840 VTAIL.n797 171.744
R1738 VTAIL.n847 VTAIL.n797 171.744
R1739 VTAIL.n848 VTAIL.n847 171.744
R1740 VTAIL.n848 VTAIL.n793 171.744
R1741 VTAIL.n856 VTAIL.n793 171.744
R1742 VTAIL.n857 VTAIL.n856 171.744
R1743 VTAIL.n858 VTAIL.n857 171.744
R1744 VTAIL.n858 VTAIL.n789 171.744
R1745 VTAIL.n865 VTAIL.n789 171.744
R1746 VTAIL.n866 VTAIL.n865 171.744
R1747 VTAIL.n866 VTAIL.n785 171.744
R1748 VTAIL.n873 VTAIL.n785 171.744
R1749 VTAIL.n874 VTAIL.n873 171.744
R1750 VTAIL.n874 VTAIL.n781 171.744
R1751 VTAIL.n881 VTAIL.n781 171.744
R1752 VTAIL.n882 VTAIL.n881 171.744
R1753 VTAIL.n40 VTAIL.n39 171.744
R1754 VTAIL.n40 VTAIL.n33 171.744
R1755 VTAIL.n47 VTAIL.n33 171.744
R1756 VTAIL.n48 VTAIL.n47 171.744
R1757 VTAIL.n48 VTAIL.n29 171.744
R1758 VTAIL.n55 VTAIL.n29 171.744
R1759 VTAIL.n56 VTAIL.n55 171.744
R1760 VTAIL.n56 VTAIL.n25 171.744
R1761 VTAIL.n63 VTAIL.n25 171.744
R1762 VTAIL.n64 VTAIL.n63 171.744
R1763 VTAIL.n64 VTAIL.n21 171.744
R1764 VTAIL.n71 VTAIL.n21 171.744
R1765 VTAIL.n72 VTAIL.n71 171.744
R1766 VTAIL.n72 VTAIL.n17 171.744
R1767 VTAIL.n80 VTAIL.n17 171.744
R1768 VTAIL.n81 VTAIL.n80 171.744
R1769 VTAIL.n82 VTAIL.n81 171.744
R1770 VTAIL.n82 VTAIL.n13 171.744
R1771 VTAIL.n89 VTAIL.n13 171.744
R1772 VTAIL.n90 VTAIL.n89 171.744
R1773 VTAIL.n90 VTAIL.n9 171.744
R1774 VTAIL.n97 VTAIL.n9 171.744
R1775 VTAIL.n98 VTAIL.n97 171.744
R1776 VTAIL.n98 VTAIL.n5 171.744
R1777 VTAIL.n105 VTAIL.n5 171.744
R1778 VTAIL.n106 VTAIL.n105 171.744
R1779 VTAIL.n150 VTAIL.n149 171.744
R1780 VTAIL.n150 VTAIL.n143 171.744
R1781 VTAIL.n157 VTAIL.n143 171.744
R1782 VTAIL.n158 VTAIL.n157 171.744
R1783 VTAIL.n158 VTAIL.n139 171.744
R1784 VTAIL.n165 VTAIL.n139 171.744
R1785 VTAIL.n166 VTAIL.n165 171.744
R1786 VTAIL.n166 VTAIL.n135 171.744
R1787 VTAIL.n173 VTAIL.n135 171.744
R1788 VTAIL.n174 VTAIL.n173 171.744
R1789 VTAIL.n174 VTAIL.n131 171.744
R1790 VTAIL.n181 VTAIL.n131 171.744
R1791 VTAIL.n182 VTAIL.n181 171.744
R1792 VTAIL.n182 VTAIL.n127 171.744
R1793 VTAIL.n190 VTAIL.n127 171.744
R1794 VTAIL.n191 VTAIL.n190 171.744
R1795 VTAIL.n192 VTAIL.n191 171.744
R1796 VTAIL.n192 VTAIL.n123 171.744
R1797 VTAIL.n199 VTAIL.n123 171.744
R1798 VTAIL.n200 VTAIL.n199 171.744
R1799 VTAIL.n200 VTAIL.n119 171.744
R1800 VTAIL.n207 VTAIL.n119 171.744
R1801 VTAIL.n208 VTAIL.n207 171.744
R1802 VTAIL.n208 VTAIL.n115 171.744
R1803 VTAIL.n215 VTAIL.n115 171.744
R1804 VTAIL.n216 VTAIL.n215 171.744
R1805 VTAIL.n262 VTAIL.n261 171.744
R1806 VTAIL.n262 VTAIL.n255 171.744
R1807 VTAIL.n269 VTAIL.n255 171.744
R1808 VTAIL.n270 VTAIL.n269 171.744
R1809 VTAIL.n270 VTAIL.n251 171.744
R1810 VTAIL.n277 VTAIL.n251 171.744
R1811 VTAIL.n278 VTAIL.n277 171.744
R1812 VTAIL.n278 VTAIL.n247 171.744
R1813 VTAIL.n285 VTAIL.n247 171.744
R1814 VTAIL.n286 VTAIL.n285 171.744
R1815 VTAIL.n286 VTAIL.n243 171.744
R1816 VTAIL.n293 VTAIL.n243 171.744
R1817 VTAIL.n294 VTAIL.n293 171.744
R1818 VTAIL.n294 VTAIL.n239 171.744
R1819 VTAIL.n302 VTAIL.n239 171.744
R1820 VTAIL.n303 VTAIL.n302 171.744
R1821 VTAIL.n304 VTAIL.n303 171.744
R1822 VTAIL.n304 VTAIL.n235 171.744
R1823 VTAIL.n311 VTAIL.n235 171.744
R1824 VTAIL.n312 VTAIL.n311 171.744
R1825 VTAIL.n312 VTAIL.n231 171.744
R1826 VTAIL.n319 VTAIL.n231 171.744
R1827 VTAIL.n320 VTAIL.n319 171.744
R1828 VTAIL.n320 VTAIL.n227 171.744
R1829 VTAIL.n327 VTAIL.n227 171.744
R1830 VTAIL.n328 VTAIL.n327 171.744
R1831 VTAIL.n772 VTAIL.n771 171.744
R1832 VTAIL.n771 VTAIL.n671 171.744
R1833 VTAIL.n764 VTAIL.n671 171.744
R1834 VTAIL.n764 VTAIL.n763 171.744
R1835 VTAIL.n763 VTAIL.n675 171.744
R1836 VTAIL.n756 VTAIL.n675 171.744
R1837 VTAIL.n756 VTAIL.n755 171.744
R1838 VTAIL.n755 VTAIL.n679 171.744
R1839 VTAIL.n684 VTAIL.n679 171.744
R1840 VTAIL.n748 VTAIL.n684 171.744
R1841 VTAIL.n748 VTAIL.n747 171.744
R1842 VTAIL.n747 VTAIL.n685 171.744
R1843 VTAIL.n740 VTAIL.n685 171.744
R1844 VTAIL.n740 VTAIL.n739 171.744
R1845 VTAIL.n739 VTAIL.n689 171.744
R1846 VTAIL.n732 VTAIL.n689 171.744
R1847 VTAIL.n732 VTAIL.n731 171.744
R1848 VTAIL.n731 VTAIL.n693 171.744
R1849 VTAIL.n724 VTAIL.n693 171.744
R1850 VTAIL.n724 VTAIL.n723 171.744
R1851 VTAIL.n723 VTAIL.n697 171.744
R1852 VTAIL.n716 VTAIL.n697 171.744
R1853 VTAIL.n716 VTAIL.n715 171.744
R1854 VTAIL.n715 VTAIL.n701 171.744
R1855 VTAIL.n708 VTAIL.n701 171.744
R1856 VTAIL.n708 VTAIL.n707 171.744
R1857 VTAIL.n660 VTAIL.n659 171.744
R1858 VTAIL.n659 VTAIL.n559 171.744
R1859 VTAIL.n652 VTAIL.n559 171.744
R1860 VTAIL.n652 VTAIL.n651 171.744
R1861 VTAIL.n651 VTAIL.n563 171.744
R1862 VTAIL.n644 VTAIL.n563 171.744
R1863 VTAIL.n644 VTAIL.n643 171.744
R1864 VTAIL.n643 VTAIL.n567 171.744
R1865 VTAIL.n572 VTAIL.n567 171.744
R1866 VTAIL.n636 VTAIL.n572 171.744
R1867 VTAIL.n636 VTAIL.n635 171.744
R1868 VTAIL.n635 VTAIL.n573 171.744
R1869 VTAIL.n628 VTAIL.n573 171.744
R1870 VTAIL.n628 VTAIL.n627 171.744
R1871 VTAIL.n627 VTAIL.n577 171.744
R1872 VTAIL.n620 VTAIL.n577 171.744
R1873 VTAIL.n620 VTAIL.n619 171.744
R1874 VTAIL.n619 VTAIL.n581 171.744
R1875 VTAIL.n612 VTAIL.n581 171.744
R1876 VTAIL.n612 VTAIL.n611 171.744
R1877 VTAIL.n611 VTAIL.n585 171.744
R1878 VTAIL.n604 VTAIL.n585 171.744
R1879 VTAIL.n604 VTAIL.n603 171.744
R1880 VTAIL.n603 VTAIL.n589 171.744
R1881 VTAIL.n596 VTAIL.n589 171.744
R1882 VTAIL.n596 VTAIL.n595 171.744
R1883 VTAIL.n550 VTAIL.n549 171.744
R1884 VTAIL.n549 VTAIL.n449 171.744
R1885 VTAIL.n542 VTAIL.n449 171.744
R1886 VTAIL.n542 VTAIL.n541 171.744
R1887 VTAIL.n541 VTAIL.n453 171.744
R1888 VTAIL.n534 VTAIL.n453 171.744
R1889 VTAIL.n534 VTAIL.n533 171.744
R1890 VTAIL.n533 VTAIL.n457 171.744
R1891 VTAIL.n462 VTAIL.n457 171.744
R1892 VTAIL.n526 VTAIL.n462 171.744
R1893 VTAIL.n526 VTAIL.n525 171.744
R1894 VTAIL.n525 VTAIL.n463 171.744
R1895 VTAIL.n518 VTAIL.n463 171.744
R1896 VTAIL.n518 VTAIL.n517 171.744
R1897 VTAIL.n517 VTAIL.n467 171.744
R1898 VTAIL.n510 VTAIL.n467 171.744
R1899 VTAIL.n510 VTAIL.n509 171.744
R1900 VTAIL.n509 VTAIL.n471 171.744
R1901 VTAIL.n502 VTAIL.n471 171.744
R1902 VTAIL.n502 VTAIL.n501 171.744
R1903 VTAIL.n501 VTAIL.n475 171.744
R1904 VTAIL.n494 VTAIL.n475 171.744
R1905 VTAIL.n494 VTAIL.n493 171.744
R1906 VTAIL.n493 VTAIL.n479 171.744
R1907 VTAIL.n486 VTAIL.n479 171.744
R1908 VTAIL.n486 VTAIL.n485 171.744
R1909 VTAIL.n438 VTAIL.n437 171.744
R1910 VTAIL.n437 VTAIL.n337 171.744
R1911 VTAIL.n430 VTAIL.n337 171.744
R1912 VTAIL.n430 VTAIL.n429 171.744
R1913 VTAIL.n429 VTAIL.n341 171.744
R1914 VTAIL.n422 VTAIL.n341 171.744
R1915 VTAIL.n422 VTAIL.n421 171.744
R1916 VTAIL.n421 VTAIL.n345 171.744
R1917 VTAIL.n350 VTAIL.n345 171.744
R1918 VTAIL.n414 VTAIL.n350 171.744
R1919 VTAIL.n414 VTAIL.n413 171.744
R1920 VTAIL.n413 VTAIL.n351 171.744
R1921 VTAIL.n406 VTAIL.n351 171.744
R1922 VTAIL.n406 VTAIL.n405 171.744
R1923 VTAIL.n405 VTAIL.n355 171.744
R1924 VTAIL.n398 VTAIL.n355 171.744
R1925 VTAIL.n398 VTAIL.n397 171.744
R1926 VTAIL.n397 VTAIL.n359 171.744
R1927 VTAIL.n390 VTAIL.n359 171.744
R1928 VTAIL.n390 VTAIL.n389 171.744
R1929 VTAIL.n389 VTAIL.n363 171.744
R1930 VTAIL.n382 VTAIL.n363 171.744
R1931 VTAIL.n382 VTAIL.n381 171.744
R1932 VTAIL.n381 VTAIL.n367 171.744
R1933 VTAIL.n374 VTAIL.n367 171.744
R1934 VTAIL.n374 VTAIL.n373 171.744
R1935 VTAIL.n815 VTAIL.t0 85.8723
R1936 VTAIL.n39 VTAIL.t7 85.8723
R1937 VTAIL.n149 VTAIL.t11 85.8723
R1938 VTAIL.n261 VTAIL.t15 85.8723
R1939 VTAIL.n707 VTAIL.t9 85.8723
R1940 VTAIL.n595 VTAIL.t8 85.8723
R1941 VTAIL.n485 VTAIL.t6 85.8723
R1942 VTAIL.n373 VTAIL.t2 85.8723
R1943 VTAIL.n667 VTAIL.n666 50.2674
R1944 VTAIL.n445 VTAIL.n444 50.2674
R1945 VTAIL.n1 VTAIL.n0 50.2672
R1946 VTAIL.n223 VTAIL.n222 50.2672
R1947 VTAIL.n887 VTAIL.n777 31.4531
R1948 VTAIL.n443 VTAIL.n333 31.4531
R1949 VTAIL.n887 VTAIL.n886 31.0217
R1950 VTAIL.n111 VTAIL.n110 31.0217
R1951 VTAIL.n221 VTAIL.n220 31.0217
R1952 VTAIL.n333 VTAIL.n332 31.0217
R1953 VTAIL.n777 VTAIL.n776 31.0217
R1954 VTAIL.n665 VTAIL.n664 31.0217
R1955 VTAIL.n555 VTAIL.n554 31.0217
R1956 VTAIL.n443 VTAIL.n442 31.0217
R1957 VTAIL.n814 VTAIL.n813 16.3895
R1958 VTAIL.n38 VTAIL.n37 16.3895
R1959 VTAIL.n148 VTAIL.n147 16.3895
R1960 VTAIL.n260 VTAIL.n259 16.3895
R1961 VTAIL.n706 VTAIL.n705 16.3895
R1962 VTAIL.n594 VTAIL.n593 16.3895
R1963 VTAIL.n484 VTAIL.n483 16.3895
R1964 VTAIL.n372 VTAIL.n371 16.3895
R1965 VTAIL.n859 VTAIL.n790 13.1884
R1966 VTAIL.n83 VTAIL.n14 13.1884
R1967 VTAIL.n193 VTAIL.n124 13.1884
R1968 VTAIL.n305 VTAIL.n236 13.1884
R1969 VTAIL.n682 VTAIL.n680 13.1884
R1970 VTAIL.n570 VTAIL.n568 13.1884
R1971 VTAIL.n460 VTAIL.n458 13.1884
R1972 VTAIL.n348 VTAIL.n346 13.1884
R1973 VTAIL.n817 VTAIL.n812 12.8005
R1974 VTAIL.n860 VTAIL.n792 12.8005
R1975 VTAIL.n864 VTAIL.n863 12.8005
R1976 VTAIL.n41 VTAIL.n36 12.8005
R1977 VTAIL.n84 VTAIL.n16 12.8005
R1978 VTAIL.n88 VTAIL.n87 12.8005
R1979 VTAIL.n151 VTAIL.n146 12.8005
R1980 VTAIL.n194 VTAIL.n126 12.8005
R1981 VTAIL.n198 VTAIL.n197 12.8005
R1982 VTAIL.n263 VTAIL.n258 12.8005
R1983 VTAIL.n306 VTAIL.n238 12.8005
R1984 VTAIL.n310 VTAIL.n309 12.8005
R1985 VTAIL.n754 VTAIL.n753 12.8005
R1986 VTAIL.n750 VTAIL.n749 12.8005
R1987 VTAIL.n709 VTAIL.n704 12.8005
R1988 VTAIL.n642 VTAIL.n641 12.8005
R1989 VTAIL.n638 VTAIL.n637 12.8005
R1990 VTAIL.n597 VTAIL.n592 12.8005
R1991 VTAIL.n532 VTAIL.n531 12.8005
R1992 VTAIL.n528 VTAIL.n527 12.8005
R1993 VTAIL.n487 VTAIL.n482 12.8005
R1994 VTAIL.n420 VTAIL.n419 12.8005
R1995 VTAIL.n416 VTAIL.n415 12.8005
R1996 VTAIL.n375 VTAIL.n370 12.8005
R1997 VTAIL.n818 VTAIL.n810 12.0247
R1998 VTAIL.n855 VTAIL.n854 12.0247
R1999 VTAIL.n867 VTAIL.n788 12.0247
R2000 VTAIL.n42 VTAIL.n34 12.0247
R2001 VTAIL.n79 VTAIL.n78 12.0247
R2002 VTAIL.n91 VTAIL.n12 12.0247
R2003 VTAIL.n152 VTAIL.n144 12.0247
R2004 VTAIL.n189 VTAIL.n188 12.0247
R2005 VTAIL.n201 VTAIL.n122 12.0247
R2006 VTAIL.n264 VTAIL.n256 12.0247
R2007 VTAIL.n301 VTAIL.n300 12.0247
R2008 VTAIL.n313 VTAIL.n234 12.0247
R2009 VTAIL.n757 VTAIL.n678 12.0247
R2010 VTAIL.n746 VTAIL.n683 12.0247
R2011 VTAIL.n710 VTAIL.n702 12.0247
R2012 VTAIL.n645 VTAIL.n566 12.0247
R2013 VTAIL.n634 VTAIL.n571 12.0247
R2014 VTAIL.n598 VTAIL.n590 12.0247
R2015 VTAIL.n535 VTAIL.n456 12.0247
R2016 VTAIL.n524 VTAIL.n461 12.0247
R2017 VTAIL.n488 VTAIL.n480 12.0247
R2018 VTAIL.n423 VTAIL.n344 12.0247
R2019 VTAIL.n412 VTAIL.n349 12.0247
R2020 VTAIL.n376 VTAIL.n368 12.0247
R2021 VTAIL.n822 VTAIL.n821 11.249
R2022 VTAIL.n853 VTAIL.n794 11.249
R2023 VTAIL.n868 VTAIL.n786 11.249
R2024 VTAIL.n46 VTAIL.n45 11.249
R2025 VTAIL.n77 VTAIL.n18 11.249
R2026 VTAIL.n92 VTAIL.n10 11.249
R2027 VTAIL.n156 VTAIL.n155 11.249
R2028 VTAIL.n187 VTAIL.n128 11.249
R2029 VTAIL.n202 VTAIL.n120 11.249
R2030 VTAIL.n268 VTAIL.n267 11.249
R2031 VTAIL.n299 VTAIL.n240 11.249
R2032 VTAIL.n314 VTAIL.n232 11.249
R2033 VTAIL.n758 VTAIL.n676 11.249
R2034 VTAIL.n745 VTAIL.n686 11.249
R2035 VTAIL.n714 VTAIL.n713 11.249
R2036 VTAIL.n646 VTAIL.n564 11.249
R2037 VTAIL.n633 VTAIL.n574 11.249
R2038 VTAIL.n602 VTAIL.n601 11.249
R2039 VTAIL.n536 VTAIL.n454 11.249
R2040 VTAIL.n523 VTAIL.n464 11.249
R2041 VTAIL.n492 VTAIL.n491 11.249
R2042 VTAIL.n424 VTAIL.n342 11.249
R2043 VTAIL.n411 VTAIL.n352 11.249
R2044 VTAIL.n380 VTAIL.n379 11.249
R2045 VTAIL.n825 VTAIL.n808 10.4732
R2046 VTAIL.n850 VTAIL.n849 10.4732
R2047 VTAIL.n872 VTAIL.n871 10.4732
R2048 VTAIL.n49 VTAIL.n32 10.4732
R2049 VTAIL.n74 VTAIL.n73 10.4732
R2050 VTAIL.n96 VTAIL.n95 10.4732
R2051 VTAIL.n159 VTAIL.n142 10.4732
R2052 VTAIL.n184 VTAIL.n183 10.4732
R2053 VTAIL.n206 VTAIL.n205 10.4732
R2054 VTAIL.n271 VTAIL.n254 10.4732
R2055 VTAIL.n296 VTAIL.n295 10.4732
R2056 VTAIL.n318 VTAIL.n317 10.4732
R2057 VTAIL.n762 VTAIL.n761 10.4732
R2058 VTAIL.n742 VTAIL.n741 10.4732
R2059 VTAIL.n717 VTAIL.n700 10.4732
R2060 VTAIL.n650 VTAIL.n649 10.4732
R2061 VTAIL.n630 VTAIL.n629 10.4732
R2062 VTAIL.n605 VTAIL.n588 10.4732
R2063 VTAIL.n540 VTAIL.n539 10.4732
R2064 VTAIL.n520 VTAIL.n519 10.4732
R2065 VTAIL.n495 VTAIL.n478 10.4732
R2066 VTAIL.n428 VTAIL.n427 10.4732
R2067 VTAIL.n408 VTAIL.n407 10.4732
R2068 VTAIL.n383 VTAIL.n366 10.4732
R2069 VTAIL.n826 VTAIL.n806 9.69747
R2070 VTAIL.n846 VTAIL.n796 9.69747
R2071 VTAIL.n875 VTAIL.n784 9.69747
R2072 VTAIL.n50 VTAIL.n30 9.69747
R2073 VTAIL.n70 VTAIL.n20 9.69747
R2074 VTAIL.n99 VTAIL.n8 9.69747
R2075 VTAIL.n160 VTAIL.n140 9.69747
R2076 VTAIL.n180 VTAIL.n130 9.69747
R2077 VTAIL.n209 VTAIL.n118 9.69747
R2078 VTAIL.n272 VTAIL.n252 9.69747
R2079 VTAIL.n292 VTAIL.n242 9.69747
R2080 VTAIL.n321 VTAIL.n230 9.69747
R2081 VTAIL.n765 VTAIL.n674 9.69747
R2082 VTAIL.n738 VTAIL.n688 9.69747
R2083 VTAIL.n718 VTAIL.n698 9.69747
R2084 VTAIL.n653 VTAIL.n562 9.69747
R2085 VTAIL.n626 VTAIL.n576 9.69747
R2086 VTAIL.n606 VTAIL.n586 9.69747
R2087 VTAIL.n543 VTAIL.n452 9.69747
R2088 VTAIL.n516 VTAIL.n466 9.69747
R2089 VTAIL.n496 VTAIL.n476 9.69747
R2090 VTAIL.n431 VTAIL.n340 9.69747
R2091 VTAIL.n404 VTAIL.n354 9.69747
R2092 VTAIL.n384 VTAIL.n364 9.69747
R2093 VTAIL.n886 VTAIL.n885 9.45567
R2094 VTAIL.n110 VTAIL.n109 9.45567
R2095 VTAIL.n220 VTAIL.n219 9.45567
R2096 VTAIL.n332 VTAIL.n331 9.45567
R2097 VTAIL.n776 VTAIL.n775 9.45567
R2098 VTAIL.n664 VTAIL.n663 9.45567
R2099 VTAIL.n554 VTAIL.n553 9.45567
R2100 VTAIL.n442 VTAIL.n441 9.45567
R2101 VTAIL.n885 VTAIL.n884 9.3005
R2102 VTAIL.n879 VTAIL.n878 9.3005
R2103 VTAIL.n877 VTAIL.n876 9.3005
R2104 VTAIL.n784 VTAIL.n783 9.3005
R2105 VTAIL.n871 VTAIL.n870 9.3005
R2106 VTAIL.n869 VTAIL.n868 9.3005
R2107 VTAIL.n788 VTAIL.n787 9.3005
R2108 VTAIL.n863 VTAIL.n862 9.3005
R2109 VTAIL.n835 VTAIL.n834 9.3005
R2110 VTAIL.n804 VTAIL.n803 9.3005
R2111 VTAIL.n829 VTAIL.n828 9.3005
R2112 VTAIL.n827 VTAIL.n826 9.3005
R2113 VTAIL.n808 VTAIL.n807 9.3005
R2114 VTAIL.n821 VTAIL.n820 9.3005
R2115 VTAIL.n819 VTAIL.n818 9.3005
R2116 VTAIL.n812 VTAIL.n811 9.3005
R2117 VTAIL.n837 VTAIL.n836 9.3005
R2118 VTAIL.n800 VTAIL.n799 9.3005
R2119 VTAIL.n843 VTAIL.n842 9.3005
R2120 VTAIL.n845 VTAIL.n844 9.3005
R2121 VTAIL.n796 VTAIL.n795 9.3005
R2122 VTAIL.n851 VTAIL.n850 9.3005
R2123 VTAIL.n853 VTAIL.n852 9.3005
R2124 VTAIL.n854 VTAIL.n791 9.3005
R2125 VTAIL.n861 VTAIL.n860 9.3005
R2126 VTAIL.n780 VTAIL.n779 9.3005
R2127 VTAIL.n109 VTAIL.n108 9.3005
R2128 VTAIL.n103 VTAIL.n102 9.3005
R2129 VTAIL.n101 VTAIL.n100 9.3005
R2130 VTAIL.n8 VTAIL.n7 9.3005
R2131 VTAIL.n95 VTAIL.n94 9.3005
R2132 VTAIL.n93 VTAIL.n92 9.3005
R2133 VTAIL.n12 VTAIL.n11 9.3005
R2134 VTAIL.n87 VTAIL.n86 9.3005
R2135 VTAIL.n59 VTAIL.n58 9.3005
R2136 VTAIL.n28 VTAIL.n27 9.3005
R2137 VTAIL.n53 VTAIL.n52 9.3005
R2138 VTAIL.n51 VTAIL.n50 9.3005
R2139 VTAIL.n32 VTAIL.n31 9.3005
R2140 VTAIL.n45 VTAIL.n44 9.3005
R2141 VTAIL.n43 VTAIL.n42 9.3005
R2142 VTAIL.n36 VTAIL.n35 9.3005
R2143 VTAIL.n61 VTAIL.n60 9.3005
R2144 VTAIL.n24 VTAIL.n23 9.3005
R2145 VTAIL.n67 VTAIL.n66 9.3005
R2146 VTAIL.n69 VTAIL.n68 9.3005
R2147 VTAIL.n20 VTAIL.n19 9.3005
R2148 VTAIL.n75 VTAIL.n74 9.3005
R2149 VTAIL.n77 VTAIL.n76 9.3005
R2150 VTAIL.n78 VTAIL.n15 9.3005
R2151 VTAIL.n85 VTAIL.n84 9.3005
R2152 VTAIL.n4 VTAIL.n3 9.3005
R2153 VTAIL.n219 VTAIL.n218 9.3005
R2154 VTAIL.n213 VTAIL.n212 9.3005
R2155 VTAIL.n211 VTAIL.n210 9.3005
R2156 VTAIL.n118 VTAIL.n117 9.3005
R2157 VTAIL.n205 VTAIL.n204 9.3005
R2158 VTAIL.n203 VTAIL.n202 9.3005
R2159 VTAIL.n122 VTAIL.n121 9.3005
R2160 VTAIL.n197 VTAIL.n196 9.3005
R2161 VTAIL.n169 VTAIL.n168 9.3005
R2162 VTAIL.n138 VTAIL.n137 9.3005
R2163 VTAIL.n163 VTAIL.n162 9.3005
R2164 VTAIL.n161 VTAIL.n160 9.3005
R2165 VTAIL.n142 VTAIL.n141 9.3005
R2166 VTAIL.n155 VTAIL.n154 9.3005
R2167 VTAIL.n153 VTAIL.n152 9.3005
R2168 VTAIL.n146 VTAIL.n145 9.3005
R2169 VTAIL.n171 VTAIL.n170 9.3005
R2170 VTAIL.n134 VTAIL.n133 9.3005
R2171 VTAIL.n177 VTAIL.n176 9.3005
R2172 VTAIL.n179 VTAIL.n178 9.3005
R2173 VTAIL.n130 VTAIL.n129 9.3005
R2174 VTAIL.n185 VTAIL.n184 9.3005
R2175 VTAIL.n187 VTAIL.n186 9.3005
R2176 VTAIL.n188 VTAIL.n125 9.3005
R2177 VTAIL.n195 VTAIL.n194 9.3005
R2178 VTAIL.n114 VTAIL.n113 9.3005
R2179 VTAIL.n331 VTAIL.n330 9.3005
R2180 VTAIL.n325 VTAIL.n324 9.3005
R2181 VTAIL.n323 VTAIL.n322 9.3005
R2182 VTAIL.n230 VTAIL.n229 9.3005
R2183 VTAIL.n317 VTAIL.n316 9.3005
R2184 VTAIL.n315 VTAIL.n314 9.3005
R2185 VTAIL.n234 VTAIL.n233 9.3005
R2186 VTAIL.n309 VTAIL.n308 9.3005
R2187 VTAIL.n281 VTAIL.n280 9.3005
R2188 VTAIL.n250 VTAIL.n249 9.3005
R2189 VTAIL.n275 VTAIL.n274 9.3005
R2190 VTAIL.n273 VTAIL.n272 9.3005
R2191 VTAIL.n254 VTAIL.n253 9.3005
R2192 VTAIL.n267 VTAIL.n266 9.3005
R2193 VTAIL.n265 VTAIL.n264 9.3005
R2194 VTAIL.n258 VTAIL.n257 9.3005
R2195 VTAIL.n283 VTAIL.n282 9.3005
R2196 VTAIL.n246 VTAIL.n245 9.3005
R2197 VTAIL.n289 VTAIL.n288 9.3005
R2198 VTAIL.n291 VTAIL.n290 9.3005
R2199 VTAIL.n242 VTAIL.n241 9.3005
R2200 VTAIL.n297 VTAIL.n296 9.3005
R2201 VTAIL.n299 VTAIL.n298 9.3005
R2202 VTAIL.n300 VTAIL.n237 9.3005
R2203 VTAIL.n307 VTAIL.n306 9.3005
R2204 VTAIL.n226 VTAIL.n225 9.3005
R2205 VTAIL.n692 VTAIL.n691 9.3005
R2206 VTAIL.n735 VTAIL.n734 9.3005
R2207 VTAIL.n737 VTAIL.n736 9.3005
R2208 VTAIL.n688 VTAIL.n687 9.3005
R2209 VTAIL.n743 VTAIL.n742 9.3005
R2210 VTAIL.n745 VTAIL.n744 9.3005
R2211 VTAIL.n683 VTAIL.n681 9.3005
R2212 VTAIL.n751 VTAIL.n750 9.3005
R2213 VTAIL.n775 VTAIL.n774 9.3005
R2214 VTAIL.n670 VTAIL.n669 9.3005
R2215 VTAIL.n769 VTAIL.n768 9.3005
R2216 VTAIL.n767 VTAIL.n766 9.3005
R2217 VTAIL.n674 VTAIL.n673 9.3005
R2218 VTAIL.n761 VTAIL.n760 9.3005
R2219 VTAIL.n759 VTAIL.n758 9.3005
R2220 VTAIL.n678 VTAIL.n677 9.3005
R2221 VTAIL.n753 VTAIL.n752 9.3005
R2222 VTAIL.n729 VTAIL.n728 9.3005
R2223 VTAIL.n727 VTAIL.n726 9.3005
R2224 VTAIL.n696 VTAIL.n695 9.3005
R2225 VTAIL.n721 VTAIL.n720 9.3005
R2226 VTAIL.n719 VTAIL.n718 9.3005
R2227 VTAIL.n700 VTAIL.n699 9.3005
R2228 VTAIL.n713 VTAIL.n712 9.3005
R2229 VTAIL.n711 VTAIL.n710 9.3005
R2230 VTAIL.n704 VTAIL.n703 9.3005
R2231 VTAIL.n580 VTAIL.n579 9.3005
R2232 VTAIL.n623 VTAIL.n622 9.3005
R2233 VTAIL.n625 VTAIL.n624 9.3005
R2234 VTAIL.n576 VTAIL.n575 9.3005
R2235 VTAIL.n631 VTAIL.n630 9.3005
R2236 VTAIL.n633 VTAIL.n632 9.3005
R2237 VTAIL.n571 VTAIL.n569 9.3005
R2238 VTAIL.n639 VTAIL.n638 9.3005
R2239 VTAIL.n663 VTAIL.n662 9.3005
R2240 VTAIL.n558 VTAIL.n557 9.3005
R2241 VTAIL.n657 VTAIL.n656 9.3005
R2242 VTAIL.n655 VTAIL.n654 9.3005
R2243 VTAIL.n562 VTAIL.n561 9.3005
R2244 VTAIL.n649 VTAIL.n648 9.3005
R2245 VTAIL.n647 VTAIL.n646 9.3005
R2246 VTAIL.n566 VTAIL.n565 9.3005
R2247 VTAIL.n641 VTAIL.n640 9.3005
R2248 VTAIL.n617 VTAIL.n616 9.3005
R2249 VTAIL.n615 VTAIL.n614 9.3005
R2250 VTAIL.n584 VTAIL.n583 9.3005
R2251 VTAIL.n609 VTAIL.n608 9.3005
R2252 VTAIL.n607 VTAIL.n606 9.3005
R2253 VTAIL.n588 VTAIL.n587 9.3005
R2254 VTAIL.n601 VTAIL.n600 9.3005
R2255 VTAIL.n599 VTAIL.n598 9.3005
R2256 VTAIL.n592 VTAIL.n591 9.3005
R2257 VTAIL.n470 VTAIL.n469 9.3005
R2258 VTAIL.n513 VTAIL.n512 9.3005
R2259 VTAIL.n515 VTAIL.n514 9.3005
R2260 VTAIL.n466 VTAIL.n465 9.3005
R2261 VTAIL.n521 VTAIL.n520 9.3005
R2262 VTAIL.n523 VTAIL.n522 9.3005
R2263 VTAIL.n461 VTAIL.n459 9.3005
R2264 VTAIL.n529 VTAIL.n528 9.3005
R2265 VTAIL.n553 VTAIL.n552 9.3005
R2266 VTAIL.n448 VTAIL.n447 9.3005
R2267 VTAIL.n547 VTAIL.n546 9.3005
R2268 VTAIL.n545 VTAIL.n544 9.3005
R2269 VTAIL.n452 VTAIL.n451 9.3005
R2270 VTAIL.n539 VTAIL.n538 9.3005
R2271 VTAIL.n537 VTAIL.n536 9.3005
R2272 VTAIL.n456 VTAIL.n455 9.3005
R2273 VTAIL.n531 VTAIL.n530 9.3005
R2274 VTAIL.n507 VTAIL.n506 9.3005
R2275 VTAIL.n505 VTAIL.n504 9.3005
R2276 VTAIL.n474 VTAIL.n473 9.3005
R2277 VTAIL.n499 VTAIL.n498 9.3005
R2278 VTAIL.n497 VTAIL.n496 9.3005
R2279 VTAIL.n478 VTAIL.n477 9.3005
R2280 VTAIL.n491 VTAIL.n490 9.3005
R2281 VTAIL.n489 VTAIL.n488 9.3005
R2282 VTAIL.n482 VTAIL.n481 9.3005
R2283 VTAIL.n358 VTAIL.n357 9.3005
R2284 VTAIL.n401 VTAIL.n400 9.3005
R2285 VTAIL.n403 VTAIL.n402 9.3005
R2286 VTAIL.n354 VTAIL.n353 9.3005
R2287 VTAIL.n409 VTAIL.n408 9.3005
R2288 VTAIL.n411 VTAIL.n410 9.3005
R2289 VTAIL.n349 VTAIL.n347 9.3005
R2290 VTAIL.n417 VTAIL.n416 9.3005
R2291 VTAIL.n441 VTAIL.n440 9.3005
R2292 VTAIL.n336 VTAIL.n335 9.3005
R2293 VTAIL.n435 VTAIL.n434 9.3005
R2294 VTAIL.n433 VTAIL.n432 9.3005
R2295 VTAIL.n340 VTAIL.n339 9.3005
R2296 VTAIL.n427 VTAIL.n426 9.3005
R2297 VTAIL.n425 VTAIL.n424 9.3005
R2298 VTAIL.n344 VTAIL.n343 9.3005
R2299 VTAIL.n419 VTAIL.n418 9.3005
R2300 VTAIL.n395 VTAIL.n394 9.3005
R2301 VTAIL.n393 VTAIL.n392 9.3005
R2302 VTAIL.n362 VTAIL.n361 9.3005
R2303 VTAIL.n387 VTAIL.n386 9.3005
R2304 VTAIL.n385 VTAIL.n384 9.3005
R2305 VTAIL.n366 VTAIL.n365 9.3005
R2306 VTAIL.n379 VTAIL.n378 9.3005
R2307 VTAIL.n377 VTAIL.n376 9.3005
R2308 VTAIL.n370 VTAIL.n369 9.3005
R2309 VTAIL.n830 VTAIL.n829 8.92171
R2310 VTAIL.n845 VTAIL.n798 8.92171
R2311 VTAIL.n876 VTAIL.n782 8.92171
R2312 VTAIL.n54 VTAIL.n53 8.92171
R2313 VTAIL.n69 VTAIL.n22 8.92171
R2314 VTAIL.n100 VTAIL.n6 8.92171
R2315 VTAIL.n164 VTAIL.n163 8.92171
R2316 VTAIL.n179 VTAIL.n132 8.92171
R2317 VTAIL.n210 VTAIL.n116 8.92171
R2318 VTAIL.n276 VTAIL.n275 8.92171
R2319 VTAIL.n291 VTAIL.n244 8.92171
R2320 VTAIL.n322 VTAIL.n228 8.92171
R2321 VTAIL.n766 VTAIL.n672 8.92171
R2322 VTAIL.n737 VTAIL.n690 8.92171
R2323 VTAIL.n722 VTAIL.n721 8.92171
R2324 VTAIL.n654 VTAIL.n560 8.92171
R2325 VTAIL.n625 VTAIL.n578 8.92171
R2326 VTAIL.n610 VTAIL.n609 8.92171
R2327 VTAIL.n544 VTAIL.n450 8.92171
R2328 VTAIL.n515 VTAIL.n468 8.92171
R2329 VTAIL.n500 VTAIL.n499 8.92171
R2330 VTAIL.n432 VTAIL.n338 8.92171
R2331 VTAIL.n403 VTAIL.n356 8.92171
R2332 VTAIL.n388 VTAIL.n387 8.92171
R2333 VTAIL.n833 VTAIL.n804 8.14595
R2334 VTAIL.n842 VTAIL.n841 8.14595
R2335 VTAIL.n880 VTAIL.n879 8.14595
R2336 VTAIL.n57 VTAIL.n28 8.14595
R2337 VTAIL.n66 VTAIL.n65 8.14595
R2338 VTAIL.n104 VTAIL.n103 8.14595
R2339 VTAIL.n167 VTAIL.n138 8.14595
R2340 VTAIL.n176 VTAIL.n175 8.14595
R2341 VTAIL.n214 VTAIL.n213 8.14595
R2342 VTAIL.n279 VTAIL.n250 8.14595
R2343 VTAIL.n288 VTAIL.n287 8.14595
R2344 VTAIL.n326 VTAIL.n325 8.14595
R2345 VTAIL.n770 VTAIL.n769 8.14595
R2346 VTAIL.n734 VTAIL.n733 8.14595
R2347 VTAIL.n725 VTAIL.n696 8.14595
R2348 VTAIL.n658 VTAIL.n657 8.14595
R2349 VTAIL.n622 VTAIL.n621 8.14595
R2350 VTAIL.n613 VTAIL.n584 8.14595
R2351 VTAIL.n548 VTAIL.n547 8.14595
R2352 VTAIL.n512 VTAIL.n511 8.14595
R2353 VTAIL.n503 VTAIL.n474 8.14595
R2354 VTAIL.n436 VTAIL.n435 8.14595
R2355 VTAIL.n400 VTAIL.n399 8.14595
R2356 VTAIL.n391 VTAIL.n362 8.14595
R2357 VTAIL.n834 VTAIL.n802 7.3702
R2358 VTAIL.n838 VTAIL.n800 7.3702
R2359 VTAIL.n883 VTAIL.n780 7.3702
R2360 VTAIL.n886 VTAIL.n778 7.3702
R2361 VTAIL.n58 VTAIL.n26 7.3702
R2362 VTAIL.n62 VTAIL.n24 7.3702
R2363 VTAIL.n107 VTAIL.n4 7.3702
R2364 VTAIL.n110 VTAIL.n2 7.3702
R2365 VTAIL.n168 VTAIL.n136 7.3702
R2366 VTAIL.n172 VTAIL.n134 7.3702
R2367 VTAIL.n217 VTAIL.n114 7.3702
R2368 VTAIL.n220 VTAIL.n112 7.3702
R2369 VTAIL.n280 VTAIL.n248 7.3702
R2370 VTAIL.n284 VTAIL.n246 7.3702
R2371 VTAIL.n329 VTAIL.n226 7.3702
R2372 VTAIL.n332 VTAIL.n224 7.3702
R2373 VTAIL.n776 VTAIL.n668 7.3702
R2374 VTAIL.n773 VTAIL.n670 7.3702
R2375 VTAIL.n730 VTAIL.n692 7.3702
R2376 VTAIL.n726 VTAIL.n694 7.3702
R2377 VTAIL.n664 VTAIL.n556 7.3702
R2378 VTAIL.n661 VTAIL.n558 7.3702
R2379 VTAIL.n618 VTAIL.n580 7.3702
R2380 VTAIL.n614 VTAIL.n582 7.3702
R2381 VTAIL.n554 VTAIL.n446 7.3702
R2382 VTAIL.n551 VTAIL.n448 7.3702
R2383 VTAIL.n508 VTAIL.n470 7.3702
R2384 VTAIL.n504 VTAIL.n472 7.3702
R2385 VTAIL.n442 VTAIL.n334 7.3702
R2386 VTAIL.n439 VTAIL.n336 7.3702
R2387 VTAIL.n396 VTAIL.n358 7.3702
R2388 VTAIL.n392 VTAIL.n360 7.3702
R2389 VTAIL.n837 VTAIL.n802 6.59444
R2390 VTAIL.n838 VTAIL.n837 6.59444
R2391 VTAIL.n884 VTAIL.n883 6.59444
R2392 VTAIL.n884 VTAIL.n778 6.59444
R2393 VTAIL.n61 VTAIL.n26 6.59444
R2394 VTAIL.n62 VTAIL.n61 6.59444
R2395 VTAIL.n108 VTAIL.n107 6.59444
R2396 VTAIL.n108 VTAIL.n2 6.59444
R2397 VTAIL.n171 VTAIL.n136 6.59444
R2398 VTAIL.n172 VTAIL.n171 6.59444
R2399 VTAIL.n218 VTAIL.n217 6.59444
R2400 VTAIL.n218 VTAIL.n112 6.59444
R2401 VTAIL.n283 VTAIL.n248 6.59444
R2402 VTAIL.n284 VTAIL.n283 6.59444
R2403 VTAIL.n330 VTAIL.n329 6.59444
R2404 VTAIL.n330 VTAIL.n224 6.59444
R2405 VTAIL.n774 VTAIL.n668 6.59444
R2406 VTAIL.n774 VTAIL.n773 6.59444
R2407 VTAIL.n730 VTAIL.n729 6.59444
R2408 VTAIL.n729 VTAIL.n694 6.59444
R2409 VTAIL.n662 VTAIL.n556 6.59444
R2410 VTAIL.n662 VTAIL.n661 6.59444
R2411 VTAIL.n618 VTAIL.n617 6.59444
R2412 VTAIL.n617 VTAIL.n582 6.59444
R2413 VTAIL.n552 VTAIL.n446 6.59444
R2414 VTAIL.n552 VTAIL.n551 6.59444
R2415 VTAIL.n508 VTAIL.n507 6.59444
R2416 VTAIL.n507 VTAIL.n472 6.59444
R2417 VTAIL.n440 VTAIL.n334 6.59444
R2418 VTAIL.n440 VTAIL.n439 6.59444
R2419 VTAIL.n396 VTAIL.n395 6.59444
R2420 VTAIL.n395 VTAIL.n360 6.59444
R2421 VTAIL.n834 VTAIL.n833 5.81868
R2422 VTAIL.n841 VTAIL.n800 5.81868
R2423 VTAIL.n880 VTAIL.n780 5.81868
R2424 VTAIL.n58 VTAIL.n57 5.81868
R2425 VTAIL.n65 VTAIL.n24 5.81868
R2426 VTAIL.n104 VTAIL.n4 5.81868
R2427 VTAIL.n168 VTAIL.n167 5.81868
R2428 VTAIL.n175 VTAIL.n134 5.81868
R2429 VTAIL.n214 VTAIL.n114 5.81868
R2430 VTAIL.n280 VTAIL.n279 5.81868
R2431 VTAIL.n287 VTAIL.n246 5.81868
R2432 VTAIL.n326 VTAIL.n226 5.81868
R2433 VTAIL.n770 VTAIL.n670 5.81868
R2434 VTAIL.n733 VTAIL.n692 5.81868
R2435 VTAIL.n726 VTAIL.n725 5.81868
R2436 VTAIL.n658 VTAIL.n558 5.81868
R2437 VTAIL.n621 VTAIL.n580 5.81868
R2438 VTAIL.n614 VTAIL.n613 5.81868
R2439 VTAIL.n548 VTAIL.n448 5.81868
R2440 VTAIL.n511 VTAIL.n470 5.81868
R2441 VTAIL.n504 VTAIL.n503 5.81868
R2442 VTAIL.n436 VTAIL.n336 5.81868
R2443 VTAIL.n399 VTAIL.n358 5.81868
R2444 VTAIL.n392 VTAIL.n391 5.81868
R2445 VTAIL.n830 VTAIL.n804 5.04292
R2446 VTAIL.n842 VTAIL.n798 5.04292
R2447 VTAIL.n879 VTAIL.n782 5.04292
R2448 VTAIL.n54 VTAIL.n28 5.04292
R2449 VTAIL.n66 VTAIL.n22 5.04292
R2450 VTAIL.n103 VTAIL.n6 5.04292
R2451 VTAIL.n164 VTAIL.n138 5.04292
R2452 VTAIL.n176 VTAIL.n132 5.04292
R2453 VTAIL.n213 VTAIL.n116 5.04292
R2454 VTAIL.n276 VTAIL.n250 5.04292
R2455 VTAIL.n288 VTAIL.n244 5.04292
R2456 VTAIL.n325 VTAIL.n228 5.04292
R2457 VTAIL.n769 VTAIL.n672 5.04292
R2458 VTAIL.n734 VTAIL.n690 5.04292
R2459 VTAIL.n722 VTAIL.n696 5.04292
R2460 VTAIL.n657 VTAIL.n560 5.04292
R2461 VTAIL.n622 VTAIL.n578 5.04292
R2462 VTAIL.n610 VTAIL.n584 5.04292
R2463 VTAIL.n547 VTAIL.n450 5.04292
R2464 VTAIL.n512 VTAIL.n468 5.04292
R2465 VTAIL.n500 VTAIL.n474 5.04292
R2466 VTAIL.n435 VTAIL.n338 5.04292
R2467 VTAIL.n400 VTAIL.n356 5.04292
R2468 VTAIL.n388 VTAIL.n362 5.04292
R2469 VTAIL.n829 VTAIL.n806 4.26717
R2470 VTAIL.n846 VTAIL.n845 4.26717
R2471 VTAIL.n876 VTAIL.n875 4.26717
R2472 VTAIL.n53 VTAIL.n30 4.26717
R2473 VTAIL.n70 VTAIL.n69 4.26717
R2474 VTAIL.n100 VTAIL.n99 4.26717
R2475 VTAIL.n163 VTAIL.n140 4.26717
R2476 VTAIL.n180 VTAIL.n179 4.26717
R2477 VTAIL.n210 VTAIL.n209 4.26717
R2478 VTAIL.n275 VTAIL.n252 4.26717
R2479 VTAIL.n292 VTAIL.n291 4.26717
R2480 VTAIL.n322 VTAIL.n321 4.26717
R2481 VTAIL.n766 VTAIL.n765 4.26717
R2482 VTAIL.n738 VTAIL.n737 4.26717
R2483 VTAIL.n721 VTAIL.n698 4.26717
R2484 VTAIL.n654 VTAIL.n653 4.26717
R2485 VTAIL.n626 VTAIL.n625 4.26717
R2486 VTAIL.n609 VTAIL.n586 4.26717
R2487 VTAIL.n544 VTAIL.n543 4.26717
R2488 VTAIL.n516 VTAIL.n515 4.26717
R2489 VTAIL.n499 VTAIL.n476 4.26717
R2490 VTAIL.n432 VTAIL.n431 4.26717
R2491 VTAIL.n404 VTAIL.n403 4.26717
R2492 VTAIL.n387 VTAIL.n364 4.26717
R2493 VTAIL.n813 VTAIL.n811 3.70982
R2494 VTAIL.n37 VTAIL.n35 3.70982
R2495 VTAIL.n147 VTAIL.n145 3.70982
R2496 VTAIL.n259 VTAIL.n257 3.70982
R2497 VTAIL.n705 VTAIL.n703 3.70982
R2498 VTAIL.n593 VTAIL.n591 3.70982
R2499 VTAIL.n483 VTAIL.n481 3.70982
R2500 VTAIL.n371 VTAIL.n369 3.70982
R2501 VTAIL.n826 VTAIL.n825 3.49141
R2502 VTAIL.n849 VTAIL.n796 3.49141
R2503 VTAIL.n872 VTAIL.n784 3.49141
R2504 VTAIL.n50 VTAIL.n49 3.49141
R2505 VTAIL.n73 VTAIL.n20 3.49141
R2506 VTAIL.n96 VTAIL.n8 3.49141
R2507 VTAIL.n160 VTAIL.n159 3.49141
R2508 VTAIL.n183 VTAIL.n130 3.49141
R2509 VTAIL.n206 VTAIL.n118 3.49141
R2510 VTAIL.n272 VTAIL.n271 3.49141
R2511 VTAIL.n295 VTAIL.n242 3.49141
R2512 VTAIL.n318 VTAIL.n230 3.49141
R2513 VTAIL.n762 VTAIL.n674 3.49141
R2514 VTAIL.n741 VTAIL.n688 3.49141
R2515 VTAIL.n718 VTAIL.n717 3.49141
R2516 VTAIL.n650 VTAIL.n562 3.49141
R2517 VTAIL.n629 VTAIL.n576 3.49141
R2518 VTAIL.n606 VTAIL.n605 3.49141
R2519 VTAIL.n540 VTAIL.n452 3.49141
R2520 VTAIL.n519 VTAIL.n466 3.49141
R2521 VTAIL.n496 VTAIL.n495 3.49141
R2522 VTAIL.n428 VTAIL.n340 3.49141
R2523 VTAIL.n407 VTAIL.n354 3.49141
R2524 VTAIL.n384 VTAIL.n383 3.49141
R2525 VTAIL.n822 VTAIL.n808 2.71565
R2526 VTAIL.n850 VTAIL.n794 2.71565
R2527 VTAIL.n871 VTAIL.n786 2.71565
R2528 VTAIL.n46 VTAIL.n32 2.71565
R2529 VTAIL.n74 VTAIL.n18 2.71565
R2530 VTAIL.n95 VTAIL.n10 2.71565
R2531 VTAIL.n156 VTAIL.n142 2.71565
R2532 VTAIL.n184 VTAIL.n128 2.71565
R2533 VTAIL.n205 VTAIL.n120 2.71565
R2534 VTAIL.n268 VTAIL.n254 2.71565
R2535 VTAIL.n296 VTAIL.n240 2.71565
R2536 VTAIL.n317 VTAIL.n232 2.71565
R2537 VTAIL.n761 VTAIL.n676 2.71565
R2538 VTAIL.n742 VTAIL.n686 2.71565
R2539 VTAIL.n714 VTAIL.n700 2.71565
R2540 VTAIL.n649 VTAIL.n564 2.71565
R2541 VTAIL.n630 VTAIL.n574 2.71565
R2542 VTAIL.n602 VTAIL.n588 2.71565
R2543 VTAIL.n539 VTAIL.n454 2.71565
R2544 VTAIL.n520 VTAIL.n464 2.71565
R2545 VTAIL.n492 VTAIL.n478 2.71565
R2546 VTAIL.n427 VTAIL.n342 2.71565
R2547 VTAIL.n408 VTAIL.n352 2.71565
R2548 VTAIL.n380 VTAIL.n366 2.71565
R2549 VTAIL.n445 VTAIL.n443 2.17291
R2550 VTAIL.n555 VTAIL.n445 2.17291
R2551 VTAIL.n667 VTAIL.n665 2.17291
R2552 VTAIL.n777 VTAIL.n667 2.17291
R2553 VTAIL.n333 VTAIL.n223 2.17291
R2554 VTAIL.n223 VTAIL.n221 2.17291
R2555 VTAIL.n111 VTAIL.n1 2.17291
R2556 VTAIL VTAIL.n887 2.11472
R2557 VTAIL.n821 VTAIL.n810 1.93989
R2558 VTAIL.n855 VTAIL.n853 1.93989
R2559 VTAIL.n868 VTAIL.n867 1.93989
R2560 VTAIL.n45 VTAIL.n34 1.93989
R2561 VTAIL.n79 VTAIL.n77 1.93989
R2562 VTAIL.n92 VTAIL.n91 1.93989
R2563 VTAIL.n155 VTAIL.n144 1.93989
R2564 VTAIL.n189 VTAIL.n187 1.93989
R2565 VTAIL.n202 VTAIL.n201 1.93989
R2566 VTAIL.n267 VTAIL.n256 1.93989
R2567 VTAIL.n301 VTAIL.n299 1.93989
R2568 VTAIL.n314 VTAIL.n313 1.93989
R2569 VTAIL.n758 VTAIL.n757 1.93989
R2570 VTAIL.n746 VTAIL.n745 1.93989
R2571 VTAIL.n713 VTAIL.n702 1.93989
R2572 VTAIL.n646 VTAIL.n645 1.93989
R2573 VTAIL.n634 VTAIL.n633 1.93989
R2574 VTAIL.n601 VTAIL.n590 1.93989
R2575 VTAIL.n536 VTAIL.n535 1.93989
R2576 VTAIL.n524 VTAIL.n523 1.93989
R2577 VTAIL.n491 VTAIL.n480 1.93989
R2578 VTAIL.n424 VTAIL.n423 1.93989
R2579 VTAIL.n412 VTAIL.n411 1.93989
R2580 VTAIL.n379 VTAIL.n368 1.93989
R2581 VTAIL.n0 VTAIL.t3 1.65723
R2582 VTAIL.n0 VTAIL.t1 1.65723
R2583 VTAIL.n222 VTAIL.t13 1.65723
R2584 VTAIL.n222 VTAIL.t12 1.65723
R2585 VTAIL.n666 VTAIL.t14 1.65723
R2586 VTAIL.n666 VTAIL.t10 1.65723
R2587 VTAIL.n444 VTAIL.t5 1.65723
R2588 VTAIL.n444 VTAIL.t4 1.65723
R2589 VTAIL.n818 VTAIL.n817 1.16414
R2590 VTAIL.n854 VTAIL.n792 1.16414
R2591 VTAIL.n864 VTAIL.n788 1.16414
R2592 VTAIL.n42 VTAIL.n41 1.16414
R2593 VTAIL.n78 VTAIL.n16 1.16414
R2594 VTAIL.n88 VTAIL.n12 1.16414
R2595 VTAIL.n152 VTAIL.n151 1.16414
R2596 VTAIL.n188 VTAIL.n126 1.16414
R2597 VTAIL.n198 VTAIL.n122 1.16414
R2598 VTAIL.n264 VTAIL.n263 1.16414
R2599 VTAIL.n300 VTAIL.n238 1.16414
R2600 VTAIL.n310 VTAIL.n234 1.16414
R2601 VTAIL.n754 VTAIL.n678 1.16414
R2602 VTAIL.n749 VTAIL.n683 1.16414
R2603 VTAIL.n710 VTAIL.n709 1.16414
R2604 VTAIL.n642 VTAIL.n566 1.16414
R2605 VTAIL.n637 VTAIL.n571 1.16414
R2606 VTAIL.n598 VTAIL.n597 1.16414
R2607 VTAIL.n532 VTAIL.n456 1.16414
R2608 VTAIL.n527 VTAIL.n461 1.16414
R2609 VTAIL.n488 VTAIL.n487 1.16414
R2610 VTAIL.n420 VTAIL.n344 1.16414
R2611 VTAIL.n415 VTAIL.n349 1.16414
R2612 VTAIL.n376 VTAIL.n375 1.16414
R2613 VTAIL.n665 VTAIL.n555 0.470328
R2614 VTAIL.n221 VTAIL.n111 0.470328
R2615 VTAIL.n814 VTAIL.n812 0.388379
R2616 VTAIL.n860 VTAIL.n859 0.388379
R2617 VTAIL.n863 VTAIL.n790 0.388379
R2618 VTAIL.n38 VTAIL.n36 0.388379
R2619 VTAIL.n84 VTAIL.n83 0.388379
R2620 VTAIL.n87 VTAIL.n14 0.388379
R2621 VTAIL.n148 VTAIL.n146 0.388379
R2622 VTAIL.n194 VTAIL.n193 0.388379
R2623 VTAIL.n197 VTAIL.n124 0.388379
R2624 VTAIL.n260 VTAIL.n258 0.388379
R2625 VTAIL.n306 VTAIL.n305 0.388379
R2626 VTAIL.n309 VTAIL.n236 0.388379
R2627 VTAIL.n753 VTAIL.n680 0.388379
R2628 VTAIL.n750 VTAIL.n682 0.388379
R2629 VTAIL.n706 VTAIL.n704 0.388379
R2630 VTAIL.n641 VTAIL.n568 0.388379
R2631 VTAIL.n638 VTAIL.n570 0.388379
R2632 VTAIL.n594 VTAIL.n592 0.388379
R2633 VTAIL.n531 VTAIL.n458 0.388379
R2634 VTAIL.n528 VTAIL.n460 0.388379
R2635 VTAIL.n484 VTAIL.n482 0.388379
R2636 VTAIL.n419 VTAIL.n346 0.388379
R2637 VTAIL.n416 VTAIL.n348 0.388379
R2638 VTAIL.n372 VTAIL.n370 0.388379
R2639 VTAIL.n819 VTAIL.n811 0.155672
R2640 VTAIL.n820 VTAIL.n819 0.155672
R2641 VTAIL.n820 VTAIL.n807 0.155672
R2642 VTAIL.n827 VTAIL.n807 0.155672
R2643 VTAIL.n828 VTAIL.n827 0.155672
R2644 VTAIL.n828 VTAIL.n803 0.155672
R2645 VTAIL.n835 VTAIL.n803 0.155672
R2646 VTAIL.n836 VTAIL.n835 0.155672
R2647 VTAIL.n836 VTAIL.n799 0.155672
R2648 VTAIL.n843 VTAIL.n799 0.155672
R2649 VTAIL.n844 VTAIL.n843 0.155672
R2650 VTAIL.n844 VTAIL.n795 0.155672
R2651 VTAIL.n851 VTAIL.n795 0.155672
R2652 VTAIL.n852 VTAIL.n851 0.155672
R2653 VTAIL.n852 VTAIL.n791 0.155672
R2654 VTAIL.n861 VTAIL.n791 0.155672
R2655 VTAIL.n862 VTAIL.n861 0.155672
R2656 VTAIL.n862 VTAIL.n787 0.155672
R2657 VTAIL.n869 VTAIL.n787 0.155672
R2658 VTAIL.n870 VTAIL.n869 0.155672
R2659 VTAIL.n870 VTAIL.n783 0.155672
R2660 VTAIL.n877 VTAIL.n783 0.155672
R2661 VTAIL.n878 VTAIL.n877 0.155672
R2662 VTAIL.n878 VTAIL.n779 0.155672
R2663 VTAIL.n885 VTAIL.n779 0.155672
R2664 VTAIL.n43 VTAIL.n35 0.155672
R2665 VTAIL.n44 VTAIL.n43 0.155672
R2666 VTAIL.n44 VTAIL.n31 0.155672
R2667 VTAIL.n51 VTAIL.n31 0.155672
R2668 VTAIL.n52 VTAIL.n51 0.155672
R2669 VTAIL.n52 VTAIL.n27 0.155672
R2670 VTAIL.n59 VTAIL.n27 0.155672
R2671 VTAIL.n60 VTAIL.n59 0.155672
R2672 VTAIL.n60 VTAIL.n23 0.155672
R2673 VTAIL.n67 VTAIL.n23 0.155672
R2674 VTAIL.n68 VTAIL.n67 0.155672
R2675 VTAIL.n68 VTAIL.n19 0.155672
R2676 VTAIL.n75 VTAIL.n19 0.155672
R2677 VTAIL.n76 VTAIL.n75 0.155672
R2678 VTAIL.n76 VTAIL.n15 0.155672
R2679 VTAIL.n85 VTAIL.n15 0.155672
R2680 VTAIL.n86 VTAIL.n85 0.155672
R2681 VTAIL.n86 VTAIL.n11 0.155672
R2682 VTAIL.n93 VTAIL.n11 0.155672
R2683 VTAIL.n94 VTAIL.n93 0.155672
R2684 VTAIL.n94 VTAIL.n7 0.155672
R2685 VTAIL.n101 VTAIL.n7 0.155672
R2686 VTAIL.n102 VTAIL.n101 0.155672
R2687 VTAIL.n102 VTAIL.n3 0.155672
R2688 VTAIL.n109 VTAIL.n3 0.155672
R2689 VTAIL.n153 VTAIL.n145 0.155672
R2690 VTAIL.n154 VTAIL.n153 0.155672
R2691 VTAIL.n154 VTAIL.n141 0.155672
R2692 VTAIL.n161 VTAIL.n141 0.155672
R2693 VTAIL.n162 VTAIL.n161 0.155672
R2694 VTAIL.n162 VTAIL.n137 0.155672
R2695 VTAIL.n169 VTAIL.n137 0.155672
R2696 VTAIL.n170 VTAIL.n169 0.155672
R2697 VTAIL.n170 VTAIL.n133 0.155672
R2698 VTAIL.n177 VTAIL.n133 0.155672
R2699 VTAIL.n178 VTAIL.n177 0.155672
R2700 VTAIL.n178 VTAIL.n129 0.155672
R2701 VTAIL.n185 VTAIL.n129 0.155672
R2702 VTAIL.n186 VTAIL.n185 0.155672
R2703 VTAIL.n186 VTAIL.n125 0.155672
R2704 VTAIL.n195 VTAIL.n125 0.155672
R2705 VTAIL.n196 VTAIL.n195 0.155672
R2706 VTAIL.n196 VTAIL.n121 0.155672
R2707 VTAIL.n203 VTAIL.n121 0.155672
R2708 VTAIL.n204 VTAIL.n203 0.155672
R2709 VTAIL.n204 VTAIL.n117 0.155672
R2710 VTAIL.n211 VTAIL.n117 0.155672
R2711 VTAIL.n212 VTAIL.n211 0.155672
R2712 VTAIL.n212 VTAIL.n113 0.155672
R2713 VTAIL.n219 VTAIL.n113 0.155672
R2714 VTAIL.n265 VTAIL.n257 0.155672
R2715 VTAIL.n266 VTAIL.n265 0.155672
R2716 VTAIL.n266 VTAIL.n253 0.155672
R2717 VTAIL.n273 VTAIL.n253 0.155672
R2718 VTAIL.n274 VTAIL.n273 0.155672
R2719 VTAIL.n274 VTAIL.n249 0.155672
R2720 VTAIL.n281 VTAIL.n249 0.155672
R2721 VTAIL.n282 VTAIL.n281 0.155672
R2722 VTAIL.n282 VTAIL.n245 0.155672
R2723 VTAIL.n289 VTAIL.n245 0.155672
R2724 VTAIL.n290 VTAIL.n289 0.155672
R2725 VTAIL.n290 VTAIL.n241 0.155672
R2726 VTAIL.n297 VTAIL.n241 0.155672
R2727 VTAIL.n298 VTAIL.n297 0.155672
R2728 VTAIL.n298 VTAIL.n237 0.155672
R2729 VTAIL.n307 VTAIL.n237 0.155672
R2730 VTAIL.n308 VTAIL.n307 0.155672
R2731 VTAIL.n308 VTAIL.n233 0.155672
R2732 VTAIL.n315 VTAIL.n233 0.155672
R2733 VTAIL.n316 VTAIL.n315 0.155672
R2734 VTAIL.n316 VTAIL.n229 0.155672
R2735 VTAIL.n323 VTAIL.n229 0.155672
R2736 VTAIL.n324 VTAIL.n323 0.155672
R2737 VTAIL.n324 VTAIL.n225 0.155672
R2738 VTAIL.n331 VTAIL.n225 0.155672
R2739 VTAIL.n775 VTAIL.n669 0.155672
R2740 VTAIL.n768 VTAIL.n669 0.155672
R2741 VTAIL.n768 VTAIL.n767 0.155672
R2742 VTAIL.n767 VTAIL.n673 0.155672
R2743 VTAIL.n760 VTAIL.n673 0.155672
R2744 VTAIL.n760 VTAIL.n759 0.155672
R2745 VTAIL.n759 VTAIL.n677 0.155672
R2746 VTAIL.n752 VTAIL.n677 0.155672
R2747 VTAIL.n752 VTAIL.n751 0.155672
R2748 VTAIL.n751 VTAIL.n681 0.155672
R2749 VTAIL.n744 VTAIL.n681 0.155672
R2750 VTAIL.n744 VTAIL.n743 0.155672
R2751 VTAIL.n743 VTAIL.n687 0.155672
R2752 VTAIL.n736 VTAIL.n687 0.155672
R2753 VTAIL.n736 VTAIL.n735 0.155672
R2754 VTAIL.n735 VTAIL.n691 0.155672
R2755 VTAIL.n728 VTAIL.n691 0.155672
R2756 VTAIL.n728 VTAIL.n727 0.155672
R2757 VTAIL.n727 VTAIL.n695 0.155672
R2758 VTAIL.n720 VTAIL.n695 0.155672
R2759 VTAIL.n720 VTAIL.n719 0.155672
R2760 VTAIL.n719 VTAIL.n699 0.155672
R2761 VTAIL.n712 VTAIL.n699 0.155672
R2762 VTAIL.n712 VTAIL.n711 0.155672
R2763 VTAIL.n711 VTAIL.n703 0.155672
R2764 VTAIL.n663 VTAIL.n557 0.155672
R2765 VTAIL.n656 VTAIL.n557 0.155672
R2766 VTAIL.n656 VTAIL.n655 0.155672
R2767 VTAIL.n655 VTAIL.n561 0.155672
R2768 VTAIL.n648 VTAIL.n561 0.155672
R2769 VTAIL.n648 VTAIL.n647 0.155672
R2770 VTAIL.n647 VTAIL.n565 0.155672
R2771 VTAIL.n640 VTAIL.n565 0.155672
R2772 VTAIL.n640 VTAIL.n639 0.155672
R2773 VTAIL.n639 VTAIL.n569 0.155672
R2774 VTAIL.n632 VTAIL.n569 0.155672
R2775 VTAIL.n632 VTAIL.n631 0.155672
R2776 VTAIL.n631 VTAIL.n575 0.155672
R2777 VTAIL.n624 VTAIL.n575 0.155672
R2778 VTAIL.n624 VTAIL.n623 0.155672
R2779 VTAIL.n623 VTAIL.n579 0.155672
R2780 VTAIL.n616 VTAIL.n579 0.155672
R2781 VTAIL.n616 VTAIL.n615 0.155672
R2782 VTAIL.n615 VTAIL.n583 0.155672
R2783 VTAIL.n608 VTAIL.n583 0.155672
R2784 VTAIL.n608 VTAIL.n607 0.155672
R2785 VTAIL.n607 VTAIL.n587 0.155672
R2786 VTAIL.n600 VTAIL.n587 0.155672
R2787 VTAIL.n600 VTAIL.n599 0.155672
R2788 VTAIL.n599 VTAIL.n591 0.155672
R2789 VTAIL.n553 VTAIL.n447 0.155672
R2790 VTAIL.n546 VTAIL.n447 0.155672
R2791 VTAIL.n546 VTAIL.n545 0.155672
R2792 VTAIL.n545 VTAIL.n451 0.155672
R2793 VTAIL.n538 VTAIL.n451 0.155672
R2794 VTAIL.n538 VTAIL.n537 0.155672
R2795 VTAIL.n537 VTAIL.n455 0.155672
R2796 VTAIL.n530 VTAIL.n455 0.155672
R2797 VTAIL.n530 VTAIL.n529 0.155672
R2798 VTAIL.n529 VTAIL.n459 0.155672
R2799 VTAIL.n522 VTAIL.n459 0.155672
R2800 VTAIL.n522 VTAIL.n521 0.155672
R2801 VTAIL.n521 VTAIL.n465 0.155672
R2802 VTAIL.n514 VTAIL.n465 0.155672
R2803 VTAIL.n514 VTAIL.n513 0.155672
R2804 VTAIL.n513 VTAIL.n469 0.155672
R2805 VTAIL.n506 VTAIL.n469 0.155672
R2806 VTAIL.n506 VTAIL.n505 0.155672
R2807 VTAIL.n505 VTAIL.n473 0.155672
R2808 VTAIL.n498 VTAIL.n473 0.155672
R2809 VTAIL.n498 VTAIL.n497 0.155672
R2810 VTAIL.n497 VTAIL.n477 0.155672
R2811 VTAIL.n490 VTAIL.n477 0.155672
R2812 VTAIL.n490 VTAIL.n489 0.155672
R2813 VTAIL.n489 VTAIL.n481 0.155672
R2814 VTAIL.n441 VTAIL.n335 0.155672
R2815 VTAIL.n434 VTAIL.n335 0.155672
R2816 VTAIL.n434 VTAIL.n433 0.155672
R2817 VTAIL.n433 VTAIL.n339 0.155672
R2818 VTAIL.n426 VTAIL.n339 0.155672
R2819 VTAIL.n426 VTAIL.n425 0.155672
R2820 VTAIL.n425 VTAIL.n343 0.155672
R2821 VTAIL.n418 VTAIL.n343 0.155672
R2822 VTAIL.n418 VTAIL.n417 0.155672
R2823 VTAIL.n417 VTAIL.n347 0.155672
R2824 VTAIL.n410 VTAIL.n347 0.155672
R2825 VTAIL.n410 VTAIL.n409 0.155672
R2826 VTAIL.n409 VTAIL.n353 0.155672
R2827 VTAIL.n402 VTAIL.n353 0.155672
R2828 VTAIL.n402 VTAIL.n401 0.155672
R2829 VTAIL.n401 VTAIL.n357 0.155672
R2830 VTAIL.n394 VTAIL.n357 0.155672
R2831 VTAIL.n394 VTAIL.n393 0.155672
R2832 VTAIL.n393 VTAIL.n361 0.155672
R2833 VTAIL.n386 VTAIL.n361 0.155672
R2834 VTAIL.n386 VTAIL.n385 0.155672
R2835 VTAIL.n385 VTAIL.n365 0.155672
R2836 VTAIL.n378 VTAIL.n365 0.155672
R2837 VTAIL.n378 VTAIL.n377 0.155672
R2838 VTAIL.n377 VTAIL.n369 0.155672
R2839 VTAIL VTAIL.n1 0.0586897
R2840 VDD1 VDD1.n0 68.0905
R2841 VDD1.n3 VDD1.n2 67.9768
R2842 VDD1.n3 VDD1.n1 67.9768
R2843 VDD1.n5 VDD1.n4 66.9459
R2844 VDD1.n5 VDD1.n3 50.988
R2845 VDD1.n4 VDD1.t6 1.65723
R2846 VDD1.n4 VDD1.t7 1.65723
R2847 VDD1.n0 VDD1.t2 1.65723
R2848 VDD1.n0 VDD1.t1 1.65723
R2849 VDD1.n2 VDD1.t4 1.65723
R2850 VDD1.n2 VDD1.t0 1.65723
R2851 VDD1.n1 VDD1.t3 1.65723
R2852 VDD1.n1 VDD1.t5 1.65723
R2853 VDD1 VDD1.n5 1.02852
R2854 VN.n6 VN.t5 248.438
R2855 VN.n31 VN.t3 248.438
R2856 VN.n5 VN.t6 215.911
R2857 VN.n15 VN.t2 215.911
R2858 VN.n23 VN.t1 215.911
R2859 VN.n30 VN.t4 215.911
R2860 VN.n40 VN.t7 215.911
R2861 VN.n48 VN.t0 215.911
R2862 VN.n47 VN.n25 161.3
R2863 VN.n46 VN.n45 161.3
R2864 VN.n44 VN.n26 161.3
R2865 VN.n43 VN.n42 161.3
R2866 VN.n41 VN.n27 161.3
R2867 VN.n39 VN.n38 161.3
R2868 VN.n37 VN.n28 161.3
R2869 VN.n36 VN.n35 161.3
R2870 VN.n34 VN.n29 161.3
R2871 VN.n33 VN.n32 161.3
R2872 VN.n22 VN.n0 161.3
R2873 VN.n21 VN.n20 161.3
R2874 VN.n19 VN.n1 161.3
R2875 VN.n18 VN.n17 161.3
R2876 VN.n16 VN.n2 161.3
R2877 VN.n14 VN.n13 161.3
R2878 VN.n12 VN.n3 161.3
R2879 VN.n11 VN.n10 161.3
R2880 VN.n9 VN.n4 161.3
R2881 VN.n8 VN.n7 161.3
R2882 VN.n24 VN.n23 97.1368
R2883 VN.n49 VN.n48 97.1368
R2884 VN.n6 VN.n5 58.8804
R2885 VN.n31 VN.n30 58.8804
R2886 VN VN.n49 55.0058
R2887 VN.n21 VN.n1 42.5146
R2888 VN.n46 VN.n26 42.5146
R2889 VN.n10 VN.n9 40.577
R2890 VN.n10 VN.n3 40.577
R2891 VN.n35 VN.n34 40.577
R2892 VN.n35 VN.n28 40.577
R2893 VN.n17 VN.n1 38.6395
R2894 VN.n42 VN.n26 38.6395
R2895 VN.n9 VN.n8 24.5923
R2896 VN.n14 VN.n3 24.5923
R2897 VN.n17 VN.n16 24.5923
R2898 VN.n22 VN.n21 24.5923
R2899 VN.n34 VN.n33 24.5923
R2900 VN.n42 VN.n41 24.5923
R2901 VN.n39 VN.n28 24.5923
R2902 VN.n47 VN.n46 24.5923
R2903 VN.n23 VN.n22 13.7719
R2904 VN.n48 VN.n47 13.7719
R2905 VN.n8 VN.n5 12.7883
R2906 VN.n15 VN.n14 12.7883
R2907 VN.n33 VN.n30 12.7883
R2908 VN.n40 VN.n39 12.7883
R2909 VN.n16 VN.n15 11.8046
R2910 VN.n41 VN.n40 11.8046
R2911 VN.n32 VN.n31 9.55925
R2912 VN.n7 VN.n6 9.55925
R2913 VN.n49 VN.n25 0.278335
R2914 VN.n24 VN.n0 0.278335
R2915 VN.n45 VN.n25 0.189894
R2916 VN.n45 VN.n44 0.189894
R2917 VN.n44 VN.n43 0.189894
R2918 VN.n43 VN.n27 0.189894
R2919 VN.n38 VN.n27 0.189894
R2920 VN.n38 VN.n37 0.189894
R2921 VN.n37 VN.n36 0.189894
R2922 VN.n36 VN.n29 0.189894
R2923 VN.n32 VN.n29 0.189894
R2924 VN.n7 VN.n4 0.189894
R2925 VN.n11 VN.n4 0.189894
R2926 VN.n12 VN.n11 0.189894
R2927 VN.n13 VN.n12 0.189894
R2928 VN.n13 VN.n2 0.189894
R2929 VN.n18 VN.n2 0.189894
R2930 VN.n19 VN.n18 0.189894
R2931 VN.n20 VN.n19 0.189894
R2932 VN.n20 VN.n0 0.189894
R2933 VN VN.n24 0.153485
R2934 VDD2.n2 VDD2.n1 67.9768
R2935 VDD2.n2 VDD2.n0 67.9768
R2936 VDD2 VDD2.n5 67.974
R2937 VDD2.n4 VDD2.n3 66.9461
R2938 VDD2.n4 VDD2.n2 50.4049
R2939 VDD2.n5 VDD2.t3 1.65723
R2940 VDD2.n5 VDD2.t4 1.65723
R2941 VDD2.n3 VDD2.t7 1.65723
R2942 VDD2.n3 VDD2.t0 1.65723
R2943 VDD2.n1 VDD2.t5 1.65723
R2944 VDD2.n1 VDD2.t6 1.65723
R2945 VDD2.n0 VDD2.t2 1.65723
R2946 VDD2.n0 VDD2.t1 1.65723
R2947 VDD2 VDD2.n4 1.1449
C0 VDD1 w_n3490_n4892# 2.01891f
C1 B w_n3490_n4892# 11.6243f
C2 VDD2 w_n3490_n4892# 2.11642f
C3 VN w_n3490_n4892# 7.1354f
C4 VP w_n3490_n4892# 7.58727f
C5 VDD1 B 1.73073f
C6 VDD1 VDD2 1.56095f
C7 VTAIL w_n3490_n4892# 5.91488f
C8 VDD1 VN 0.150882f
C9 VDD2 B 1.81386f
C10 VDD1 VP 13.761201f
C11 B VN 1.22276f
C12 B VP 1.97806f
C13 VDD2 VN 13.4374f
C14 VDD1 VTAIL 10.8799f
C15 VDD2 VP 0.475938f
C16 VP VN 8.56975f
C17 B VTAIL 7.22173f
C18 VDD2 VTAIL 10.9316f
C19 VN VTAIL 13.3701f
C20 VP VTAIL 13.3842f
C21 VDD2 VSUBS 1.971573f
C22 VDD1 VSUBS 2.54613f
C23 VTAIL VSUBS 1.621269f
C24 VN VSUBS 6.57792f
C25 VP VSUBS 3.443894f
C26 B VSUBS 5.185984f
C27 w_n3490_n4892# VSUBS 0.208521p
C28 VDD2.t2 VSUBS 0.411704f
C29 VDD2.t1 VSUBS 0.411704f
C30 VDD2.n0 VSUBS 3.46025f
C31 VDD2.t5 VSUBS 0.411704f
C32 VDD2.t6 VSUBS 0.411704f
C33 VDD2.n1 VSUBS 3.46025f
C34 VDD2.n2 VSUBS 4.36928f
C35 VDD2.t7 VSUBS 0.411704f
C36 VDD2.t0 VSUBS 0.411704f
C37 VDD2.n3 VSUBS 3.44779f
C38 VDD2.n4 VSUBS 3.91341f
C39 VDD2.t3 VSUBS 0.411704f
C40 VDD2.t4 VSUBS 0.411704f
C41 VDD2.n5 VSUBS 3.4602f
C42 VN.n0 VSUBS 0.037416f
C43 VN.t1 VSUBS 3.35953f
C44 VN.n1 VSUBS 0.023068f
C45 VN.n2 VSUBS 0.028382f
C46 VN.t2 VSUBS 3.35953f
C47 VN.n3 VSUBS 0.056111f
C48 VN.n4 VSUBS 0.028382f
C49 VN.t6 VSUBS 3.35953f
C50 VN.n5 VSUBS 1.23823f
C51 VN.t5 VSUBS 3.5318f
C52 VN.n6 VSUBS 1.22917f
C53 VN.n7 VSUBS 0.241275f
C54 VN.n8 VSUBS 0.040159f
C55 VN.n9 VSUBS 0.056111f
C56 VN.n10 VSUBS 0.022923f
C57 VN.n11 VSUBS 0.028382f
C58 VN.n12 VSUBS 0.028382f
C59 VN.n13 VSUBS 0.028382f
C60 VN.n14 VSUBS 0.040159f
C61 VN.n15 VSUBS 1.16518f
C62 VN.n16 VSUBS 0.03912f
C63 VN.n17 VSUBS 0.056598f
C64 VN.n18 VSUBS 0.028382f
C65 VN.n19 VSUBS 0.028382f
C66 VN.n20 VSUBS 0.028382f
C67 VN.n21 VSUBS 0.055479f
C68 VN.n22 VSUBS 0.041199f
C69 VN.n23 VSUBS 1.24962f
C70 VN.n24 VSUBS 0.040185f
C71 VN.n25 VSUBS 0.037416f
C72 VN.t0 VSUBS 3.35953f
C73 VN.n26 VSUBS 0.023068f
C74 VN.n27 VSUBS 0.028382f
C75 VN.t7 VSUBS 3.35953f
C76 VN.n28 VSUBS 0.056111f
C77 VN.n29 VSUBS 0.028382f
C78 VN.t4 VSUBS 3.35953f
C79 VN.n30 VSUBS 1.23823f
C80 VN.t3 VSUBS 3.5318f
C81 VN.n31 VSUBS 1.22917f
C82 VN.n32 VSUBS 0.241275f
C83 VN.n33 VSUBS 0.040159f
C84 VN.n34 VSUBS 0.056111f
C85 VN.n35 VSUBS 0.022923f
C86 VN.n36 VSUBS 0.028382f
C87 VN.n37 VSUBS 0.028382f
C88 VN.n38 VSUBS 0.028382f
C89 VN.n39 VSUBS 0.040159f
C90 VN.n40 VSUBS 1.16518f
C91 VN.n41 VSUBS 0.03912f
C92 VN.n42 VSUBS 0.056598f
C93 VN.n43 VSUBS 0.028382f
C94 VN.n44 VSUBS 0.028382f
C95 VN.n45 VSUBS 0.028382f
C96 VN.n46 VSUBS 0.055479f
C97 VN.n47 VSUBS 0.041199f
C98 VN.n48 VSUBS 1.24962f
C99 VN.n49 VSUBS 1.80648f
C100 VDD1.t2 VSUBS 0.414841f
C101 VDD1.t1 VSUBS 0.414841f
C102 VDD1.n0 VSUBS 3.48814f
C103 VDD1.t3 VSUBS 0.414841f
C104 VDD1.t5 VSUBS 0.414841f
C105 VDD1.n1 VSUBS 3.48661f
C106 VDD1.t4 VSUBS 0.414841f
C107 VDD1.t0 VSUBS 0.414841f
C108 VDD1.n2 VSUBS 3.48661f
C109 VDD1.n3 VSUBS 4.45819f
C110 VDD1.t6 VSUBS 0.414841f
C111 VDD1.t7 VSUBS 0.414841f
C112 VDD1.n4 VSUBS 3.47404f
C113 VDD1.n5 VSUBS 3.97642f
C114 VTAIL.t3 VSUBS 0.358924f
C115 VTAIL.t1 VSUBS 0.358924f
C116 VTAIL.n0 VSUBS 2.85183f
C117 VTAIL.n1 VSUBS 0.75721f
C118 VTAIL.n2 VSUBS 0.025536f
C119 VTAIL.n3 VSUBS 0.02315f
C120 VTAIL.n4 VSUBS 0.01244f
C121 VTAIL.n5 VSUBS 0.029403f
C122 VTAIL.n6 VSUBS 0.013172f
C123 VTAIL.n7 VSUBS 0.02315f
C124 VTAIL.n8 VSUBS 0.01244f
C125 VTAIL.n9 VSUBS 0.029403f
C126 VTAIL.n10 VSUBS 0.013172f
C127 VTAIL.n11 VSUBS 0.02315f
C128 VTAIL.n12 VSUBS 0.01244f
C129 VTAIL.n13 VSUBS 0.029403f
C130 VTAIL.n14 VSUBS 0.012806f
C131 VTAIL.n15 VSUBS 0.02315f
C132 VTAIL.n16 VSUBS 0.013172f
C133 VTAIL.n17 VSUBS 0.029403f
C134 VTAIL.n18 VSUBS 0.013172f
C135 VTAIL.n19 VSUBS 0.02315f
C136 VTAIL.n20 VSUBS 0.01244f
C137 VTAIL.n21 VSUBS 0.029403f
C138 VTAIL.n22 VSUBS 0.013172f
C139 VTAIL.n23 VSUBS 0.02315f
C140 VTAIL.n24 VSUBS 0.01244f
C141 VTAIL.n25 VSUBS 0.029403f
C142 VTAIL.n26 VSUBS 0.013172f
C143 VTAIL.n27 VSUBS 0.02315f
C144 VTAIL.n28 VSUBS 0.01244f
C145 VTAIL.n29 VSUBS 0.029403f
C146 VTAIL.n30 VSUBS 0.013172f
C147 VTAIL.n31 VSUBS 0.02315f
C148 VTAIL.n32 VSUBS 0.01244f
C149 VTAIL.n33 VSUBS 0.029403f
C150 VTAIL.n34 VSUBS 0.013172f
C151 VTAIL.n35 VSUBS 1.9637f
C152 VTAIL.n36 VSUBS 0.01244f
C153 VTAIL.t7 VSUBS 0.063212f
C154 VTAIL.n37 VSUBS 0.194733f
C155 VTAIL.n38 VSUBS 0.018705f
C156 VTAIL.n39 VSUBS 0.022052f
C157 VTAIL.n40 VSUBS 0.029403f
C158 VTAIL.n41 VSUBS 0.013172f
C159 VTAIL.n42 VSUBS 0.01244f
C160 VTAIL.n43 VSUBS 0.02315f
C161 VTAIL.n44 VSUBS 0.02315f
C162 VTAIL.n45 VSUBS 0.01244f
C163 VTAIL.n46 VSUBS 0.013172f
C164 VTAIL.n47 VSUBS 0.029403f
C165 VTAIL.n48 VSUBS 0.029403f
C166 VTAIL.n49 VSUBS 0.013172f
C167 VTAIL.n50 VSUBS 0.01244f
C168 VTAIL.n51 VSUBS 0.02315f
C169 VTAIL.n52 VSUBS 0.02315f
C170 VTAIL.n53 VSUBS 0.01244f
C171 VTAIL.n54 VSUBS 0.013172f
C172 VTAIL.n55 VSUBS 0.029403f
C173 VTAIL.n56 VSUBS 0.029403f
C174 VTAIL.n57 VSUBS 0.013172f
C175 VTAIL.n58 VSUBS 0.01244f
C176 VTAIL.n59 VSUBS 0.02315f
C177 VTAIL.n60 VSUBS 0.02315f
C178 VTAIL.n61 VSUBS 0.01244f
C179 VTAIL.n62 VSUBS 0.013172f
C180 VTAIL.n63 VSUBS 0.029403f
C181 VTAIL.n64 VSUBS 0.029403f
C182 VTAIL.n65 VSUBS 0.013172f
C183 VTAIL.n66 VSUBS 0.01244f
C184 VTAIL.n67 VSUBS 0.02315f
C185 VTAIL.n68 VSUBS 0.02315f
C186 VTAIL.n69 VSUBS 0.01244f
C187 VTAIL.n70 VSUBS 0.013172f
C188 VTAIL.n71 VSUBS 0.029403f
C189 VTAIL.n72 VSUBS 0.029403f
C190 VTAIL.n73 VSUBS 0.013172f
C191 VTAIL.n74 VSUBS 0.01244f
C192 VTAIL.n75 VSUBS 0.02315f
C193 VTAIL.n76 VSUBS 0.02315f
C194 VTAIL.n77 VSUBS 0.01244f
C195 VTAIL.n78 VSUBS 0.01244f
C196 VTAIL.n79 VSUBS 0.013172f
C197 VTAIL.n80 VSUBS 0.029403f
C198 VTAIL.n81 VSUBS 0.029403f
C199 VTAIL.n82 VSUBS 0.029403f
C200 VTAIL.n83 VSUBS 0.012806f
C201 VTAIL.n84 VSUBS 0.01244f
C202 VTAIL.n85 VSUBS 0.02315f
C203 VTAIL.n86 VSUBS 0.02315f
C204 VTAIL.n87 VSUBS 0.01244f
C205 VTAIL.n88 VSUBS 0.013172f
C206 VTAIL.n89 VSUBS 0.029403f
C207 VTAIL.n90 VSUBS 0.029403f
C208 VTAIL.n91 VSUBS 0.013172f
C209 VTAIL.n92 VSUBS 0.01244f
C210 VTAIL.n93 VSUBS 0.02315f
C211 VTAIL.n94 VSUBS 0.02315f
C212 VTAIL.n95 VSUBS 0.01244f
C213 VTAIL.n96 VSUBS 0.013172f
C214 VTAIL.n97 VSUBS 0.029403f
C215 VTAIL.n98 VSUBS 0.029403f
C216 VTAIL.n99 VSUBS 0.013172f
C217 VTAIL.n100 VSUBS 0.01244f
C218 VTAIL.n101 VSUBS 0.02315f
C219 VTAIL.n102 VSUBS 0.02315f
C220 VTAIL.n103 VSUBS 0.01244f
C221 VTAIL.n104 VSUBS 0.013172f
C222 VTAIL.n105 VSUBS 0.029403f
C223 VTAIL.n106 VSUBS 0.07152f
C224 VTAIL.n107 VSUBS 0.013172f
C225 VTAIL.n108 VSUBS 0.01244f
C226 VTAIL.n109 VSUBS 0.051612f
C227 VTAIL.n110 VSUBS 0.035923f
C228 VTAIL.n111 VSUBS 0.215798f
C229 VTAIL.n112 VSUBS 0.025536f
C230 VTAIL.n113 VSUBS 0.02315f
C231 VTAIL.n114 VSUBS 0.01244f
C232 VTAIL.n115 VSUBS 0.029403f
C233 VTAIL.n116 VSUBS 0.013172f
C234 VTAIL.n117 VSUBS 0.02315f
C235 VTAIL.n118 VSUBS 0.01244f
C236 VTAIL.n119 VSUBS 0.029403f
C237 VTAIL.n120 VSUBS 0.013172f
C238 VTAIL.n121 VSUBS 0.02315f
C239 VTAIL.n122 VSUBS 0.01244f
C240 VTAIL.n123 VSUBS 0.029403f
C241 VTAIL.n124 VSUBS 0.012806f
C242 VTAIL.n125 VSUBS 0.02315f
C243 VTAIL.n126 VSUBS 0.013172f
C244 VTAIL.n127 VSUBS 0.029403f
C245 VTAIL.n128 VSUBS 0.013172f
C246 VTAIL.n129 VSUBS 0.02315f
C247 VTAIL.n130 VSUBS 0.01244f
C248 VTAIL.n131 VSUBS 0.029403f
C249 VTAIL.n132 VSUBS 0.013172f
C250 VTAIL.n133 VSUBS 0.02315f
C251 VTAIL.n134 VSUBS 0.01244f
C252 VTAIL.n135 VSUBS 0.029403f
C253 VTAIL.n136 VSUBS 0.013172f
C254 VTAIL.n137 VSUBS 0.02315f
C255 VTAIL.n138 VSUBS 0.01244f
C256 VTAIL.n139 VSUBS 0.029403f
C257 VTAIL.n140 VSUBS 0.013172f
C258 VTAIL.n141 VSUBS 0.02315f
C259 VTAIL.n142 VSUBS 0.01244f
C260 VTAIL.n143 VSUBS 0.029403f
C261 VTAIL.n144 VSUBS 0.013172f
C262 VTAIL.n145 VSUBS 1.9637f
C263 VTAIL.n146 VSUBS 0.01244f
C264 VTAIL.t11 VSUBS 0.063212f
C265 VTAIL.n147 VSUBS 0.194733f
C266 VTAIL.n148 VSUBS 0.018705f
C267 VTAIL.n149 VSUBS 0.022052f
C268 VTAIL.n150 VSUBS 0.029403f
C269 VTAIL.n151 VSUBS 0.013172f
C270 VTAIL.n152 VSUBS 0.01244f
C271 VTAIL.n153 VSUBS 0.02315f
C272 VTAIL.n154 VSUBS 0.02315f
C273 VTAIL.n155 VSUBS 0.01244f
C274 VTAIL.n156 VSUBS 0.013172f
C275 VTAIL.n157 VSUBS 0.029403f
C276 VTAIL.n158 VSUBS 0.029403f
C277 VTAIL.n159 VSUBS 0.013172f
C278 VTAIL.n160 VSUBS 0.01244f
C279 VTAIL.n161 VSUBS 0.02315f
C280 VTAIL.n162 VSUBS 0.02315f
C281 VTAIL.n163 VSUBS 0.01244f
C282 VTAIL.n164 VSUBS 0.013172f
C283 VTAIL.n165 VSUBS 0.029403f
C284 VTAIL.n166 VSUBS 0.029403f
C285 VTAIL.n167 VSUBS 0.013172f
C286 VTAIL.n168 VSUBS 0.01244f
C287 VTAIL.n169 VSUBS 0.02315f
C288 VTAIL.n170 VSUBS 0.02315f
C289 VTAIL.n171 VSUBS 0.01244f
C290 VTAIL.n172 VSUBS 0.013172f
C291 VTAIL.n173 VSUBS 0.029403f
C292 VTAIL.n174 VSUBS 0.029403f
C293 VTAIL.n175 VSUBS 0.013172f
C294 VTAIL.n176 VSUBS 0.01244f
C295 VTAIL.n177 VSUBS 0.02315f
C296 VTAIL.n178 VSUBS 0.02315f
C297 VTAIL.n179 VSUBS 0.01244f
C298 VTAIL.n180 VSUBS 0.013172f
C299 VTAIL.n181 VSUBS 0.029403f
C300 VTAIL.n182 VSUBS 0.029403f
C301 VTAIL.n183 VSUBS 0.013172f
C302 VTAIL.n184 VSUBS 0.01244f
C303 VTAIL.n185 VSUBS 0.02315f
C304 VTAIL.n186 VSUBS 0.02315f
C305 VTAIL.n187 VSUBS 0.01244f
C306 VTAIL.n188 VSUBS 0.01244f
C307 VTAIL.n189 VSUBS 0.013172f
C308 VTAIL.n190 VSUBS 0.029403f
C309 VTAIL.n191 VSUBS 0.029403f
C310 VTAIL.n192 VSUBS 0.029403f
C311 VTAIL.n193 VSUBS 0.012806f
C312 VTAIL.n194 VSUBS 0.01244f
C313 VTAIL.n195 VSUBS 0.02315f
C314 VTAIL.n196 VSUBS 0.02315f
C315 VTAIL.n197 VSUBS 0.01244f
C316 VTAIL.n198 VSUBS 0.013172f
C317 VTAIL.n199 VSUBS 0.029403f
C318 VTAIL.n200 VSUBS 0.029403f
C319 VTAIL.n201 VSUBS 0.013172f
C320 VTAIL.n202 VSUBS 0.01244f
C321 VTAIL.n203 VSUBS 0.02315f
C322 VTAIL.n204 VSUBS 0.02315f
C323 VTAIL.n205 VSUBS 0.01244f
C324 VTAIL.n206 VSUBS 0.013172f
C325 VTAIL.n207 VSUBS 0.029403f
C326 VTAIL.n208 VSUBS 0.029403f
C327 VTAIL.n209 VSUBS 0.013172f
C328 VTAIL.n210 VSUBS 0.01244f
C329 VTAIL.n211 VSUBS 0.02315f
C330 VTAIL.n212 VSUBS 0.02315f
C331 VTAIL.n213 VSUBS 0.01244f
C332 VTAIL.n214 VSUBS 0.013172f
C333 VTAIL.n215 VSUBS 0.029403f
C334 VTAIL.n216 VSUBS 0.07152f
C335 VTAIL.n217 VSUBS 0.013172f
C336 VTAIL.n218 VSUBS 0.01244f
C337 VTAIL.n219 VSUBS 0.051612f
C338 VTAIL.n220 VSUBS 0.035923f
C339 VTAIL.n221 VSUBS 0.215798f
C340 VTAIL.t13 VSUBS 0.358924f
C341 VTAIL.t12 VSUBS 0.358924f
C342 VTAIL.n222 VSUBS 2.85183f
C343 VTAIL.n223 VSUBS 0.914919f
C344 VTAIL.n224 VSUBS 0.025536f
C345 VTAIL.n225 VSUBS 0.02315f
C346 VTAIL.n226 VSUBS 0.01244f
C347 VTAIL.n227 VSUBS 0.029403f
C348 VTAIL.n228 VSUBS 0.013172f
C349 VTAIL.n229 VSUBS 0.02315f
C350 VTAIL.n230 VSUBS 0.01244f
C351 VTAIL.n231 VSUBS 0.029403f
C352 VTAIL.n232 VSUBS 0.013172f
C353 VTAIL.n233 VSUBS 0.02315f
C354 VTAIL.n234 VSUBS 0.01244f
C355 VTAIL.n235 VSUBS 0.029403f
C356 VTAIL.n236 VSUBS 0.012806f
C357 VTAIL.n237 VSUBS 0.02315f
C358 VTAIL.n238 VSUBS 0.013172f
C359 VTAIL.n239 VSUBS 0.029403f
C360 VTAIL.n240 VSUBS 0.013172f
C361 VTAIL.n241 VSUBS 0.02315f
C362 VTAIL.n242 VSUBS 0.01244f
C363 VTAIL.n243 VSUBS 0.029403f
C364 VTAIL.n244 VSUBS 0.013172f
C365 VTAIL.n245 VSUBS 0.02315f
C366 VTAIL.n246 VSUBS 0.01244f
C367 VTAIL.n247 VSUBS 0.029403f
C368 VTAIL.n248 VSUBS 0.013172f
C369 VTAIL.n249 VSUBS 0.02315f
C370 VTAIL.n250 VSUBS 0.01244f
C371 VTAIL.n251 VSUBS 0.029403f
C372 VTAIL.n252 VSUBS 0.013172f
C373 VTAIL.n253 VSUBS 0.02315f
C374 VTAIL.n254 VSUBS 0.01244f
C375 VTAIL.n255 VSUBS 0.029403f
C376 VTAIL.n256 VSUBS 0.013172f
C377 VTAIL.n257 VSUBS 1.9637f
C378 VTAIL.n258 VSUBS 0.01244f
C379 VTAIL.t15 VSUBS 0.063212f
C380 VTAIL.n259 VSUBS 0.194733f
C381 VTAIL.n260 VSUBS 0.018705f
C382 VTAIL.n261 VSUBS 0.022052f
C383 VTAIL.n262 VSUBS 0.029403f
C384 VTAIL.n263 VSUBS 0.013172f
C385 VTAIL.n264 VSUBS 0.01244f
C386 VTAIL.n265 VSUBS 0.02315f
C387 VTAIL.n266 VSUBS 0.02315f
C388 VTAIL.n267 VSUBS 0.01244f
C389 VTAIL.n268 VSUBS 0.013172f
C390 VTAIL.n269 VSUBS 0.029403f
C391 VTAIL.n270 VSUBS 0.029403f
C392 VTAIL.n271 VSUBS 0.013172f
C393 VTAIL.n272 VSUBS 0.01244f
C394 VTAIL.n273 VSUBS 0.02315f
C395 VTAIL.n274 VSUBS 0.02315f
C396 VTAIL.n275 VSUBS 0.01244f
C397 VTAIL.n276 VSUBS 0.013172f
C398 VTAIL.n277 VSUBS 0.029403f
C399 VTAIL.n278 VSUBS 0.029403f
C400 VTAIL.n279 VSUBS 0.013172f
C401 VTAIL.n280 VSUBS 0.01244f
C402 VTAIL.n281 VSUBS 0.02315f
C403 VTAIL.n282 VSUBS 0.02315f
C404 VTAIL.n283 VSUBS 0.01244f
C405 VTAIL.n284 VSUBS 0.013172f
C406 VTAIL.n285 VSUBS 0.029403f
C407 VTAIL.n286 VSUBS 0.029403f
C408 VTAIL.n287 VSUBS 0.013172f
C409 VTAIL.n288 VSUBS 0.01244f
C410 VTAIL.n289 VSUBS 0.02315f
C411 VTAIL.n290 VSUBS 0.02315f
C412 VTAIL.n291 VSUBS 0.01244f
C413 VTAIL.n292 VSUBS 0.013172f
C414 VTAIL.n293 VSUBS 0.029403f
C415 VTAIL.n294 VSUBS 0.029403f
C416 VTAIL.n295 VSUBS 0.013172f
C417 VTAIL.n296 VSUBS 0.01244f
C418 VTAIL.n297 VSUBS 0.02315f
C419 VTAIL.n298 VSUBS 0.02315f
C420 VTAIL.n299 VSUBS 0.01244f
C421 VTAIL.n300 VSUBS 0.01244f
C422 VTAIL.n301 VSUBS 0.013172f
C423 VTAIL.n302 VSUBS 0.029403f
C424 VTAIL.n303 VSUBS 0.029403f
C425 VTAIL.n304 VSUBS 0.029403f
C426 VTAIL.n305 VSUBS 0.012806f
C427 VTAIL.n306 VSUBS 0.01244f
C428 VTAIL.n307 VSUBS 0.02315f
C429 VTAIL.n308 VSUBS 0.02315f
C430 VTAIL.n309 VSUBS 0.01244f
C431 VTAIL.n310 VSUBS 0.013172f
C432 VTAIL.n311 VSUBS 0.029403f
C433 VTAIL.n312 VSUBS 0.029403f
C434 VTAIL.n313 VSUBS 0.013172f
C435 VTAIL.n314 VSUBS 0.01244f
C436 VTAIL.n315 VSUBS 0.02315f
C437 VTAIL.n316 VSUBS 0.02315f
C438 VTAIL.n317 VSUBS 0.01244f
C439 VTAIL.n318 VSUBS 0.013172f
C440 VTAIL.n319 VSUBS 0.029403f
C441 VTAIL.n320 VSUBS 0.029403f
C442 VTAIL.n321 VSUBS 0.013172f
C443 VTAIL.n322 VSUBS 0.01244f
C444 VTAIL.n323 VSUBS 0.02315f
C445 VTAIL.n324 VSUBS 0.02315f
C446 VTAIL.n325 VSUBS 0.01244f
C447 VTAIL.n326 VSUBS 0.013172f
C448 VTAIL.n327 VSUBS 0.029403f
C449 VTAIL.n328 VSUBS 0.07152f
C450 VTAIL.n329 VSUBS 0.013172f
C451 VTAIL.n330 VSUBS 0.01244f
C452 VTAIL.n331 VSUBS 0.051612f
C453 VTAIL.n332 VSUBS 0.035923f
C454 VTAIL.n333 VSUBS 1.91894f
C455 VTAIL.n334 VSUBS 0.025536f
C456 VTAIL.n335 VSUBS 0.02315f
C457 VTAIL.n336 VSUBS 0.01244f
C458 VTAIL.n337 VSUBS 0.029403f
C459 VTAIL.n338 VSUBS 0.013172f
C460 VTAIL.n339 VSUBS 0.02315f
C461 VTAIL.n340 VSUBS 0.01244f
C462 VTAIL.n341 VSUBS 0.029403f
C463 VTAIL.n342 VSUBS 0.013172f
C464 VTAIL.n343 VSUBS 0.02315f
C465 VTAIL.n344 VSUBS 0.01244f
C466 VTAIL.n345 VSUBS 0.029403f
C467 VTAIL.n346 VSUBS 0.012806f
C468 VTAIL.n347 VSUBS 0.02315f
C469 VTAIL.n348 VSUBS 0.012806f
C470 VTAIL.n349 VSUBS 0.01244f
C471 VTAIL.n350 VSUBS 0.029403f
C472 VTAIL.n351 VSUBS 0.029403f
C473 VTAIL.n352 VSUBS 0.013172f
C474 VTAIL.n353 VSUBS 0.02315f
C475 VTAIL.n354 VSUBS 0.01244f
C476 VTAIL.n355 VSUBS 0.029403f
C477 VTAIL.n356 VSUBS 0.013172f
C478 VTAIL.n357 VSUBS 0.02315f
C479 VTAIL.n358 VSUBS 0.01244f
C480 VTAIL.n359 VSUBS 0.029403f
C481 VTAIL.n360 VSUBS 0.013172f
C482 VTAIL.n361 VSUBS 0.02315f
C483 VTAIL.n362 VSUBS 0.01244f
C484 VTAIL.n363 VSUBS 0.029403f
C485 VTAIL.n364 VSUBS 0.013172f
C486 VTAIL.n365 VSUBS 0.02315f
C487 VTAIL.n366 VSUBS 0.01244f
C488 VTAIL.n367 VSUBS 0.029403f
C489 VTAIL.n368 VSUBS 0.013172f
C490 VTAIL.n369 VSUBS 1.9637f
C491 VTAIL.n370 VSUBS 0.01244f
C492 VTAIL.t2 VSUBS 0.063212f
C493 VTAIL.n371 VSUBS 0.194733f
C494 VTAIL.n372 VSUBS 0.018705f
C495 VTAIL.n373 VSUBS 0.022052f
C496 VTAIL.n374 VSUBS 0.029403f
C497 VTAIL.n375 VSUBS 0.013172f
C498 VTAIL.n376 VSUBS 0.01244f
C499 VTAIL.n377 VSUBS 0.02315f
C500 VTAIL.n378 VSUBS 0.02315f
C501 VTAIL.n379 VSUBS 0.01244f
C502 VTAIL.n380 VSUBS 0.013172f
C503 VTAIL.n381 VSUBS 0.029403f
C504 VTAIL.n382 VSUBS 0.029403f
C505 VTAIL.n383 VSUBS 0.013172f
C506 VTAIL.n384 VSUBS 0.01244f
C507 VTAIL.n385 VSUBS 0.02315f
C508 VTAIL.n386 VSUBS 0.02315f
C509 VTAIL.n387 VSUBS 0.01244f
C510 VTAIL.n388 VSUBS 0.013172f
C511 VTAIL.n389 VSUBS 0.029403f
C512 VTAIL.n390 VSUBS 0.029403f
C513 VTAIL.n391 VSUBS 0.013172f
C514 VTAIL.n392 VSUBS 0.01244f
C515 VTAIL.n393 VSUBS 0.02315f
C516 VTAIL.n394 VSUBS 0.02315f
C517 VTAIL.n395 VSUBS 0.01244f
C518 VTAIL.n396 VSUBS 0.013172f
C519 VTAIL.n397 VSUBS 0.029403f
C520 VTAIL.n398 VSUBS 0.029403f
C521 VTAIL.n399 VSUBS 0.013172f
C522 VTAIL.n400 VSUBS 0.01244f
C523 VTAIL.n401 VSUBS 0.02315f
C524 VTAIL.n402 VSUBS 0.02315f
C525 VTAIL.n403 VSUBS 0.01244f
C526 VTAIL.n404 VSUBS 0.013172f
C527 VTAIL.n405 VSUBS 0.029403f
C528 VTAIL.n406 VSUBS 0.029403f
C529 VTAIL.n407 VSUBS 0.013172f
C530 VTAIL.n408 VSUBS 0.01244f
C531 VTAIL.n409 VSUBS 0.02315f
C532 VTAIL.n410 VSUBS 0.02315f
C533 VTAIL.n411 VSUBS 0.01244f
C534 VTAIL.n412 VSUBS 0.013172f
C535 VTAIL.n413 VSUBS 0.029403f
C536 VTAIL.n414 VSUBS 0.029403f
C537 VTAIL.n415 VSUBS 0.013172f
C538 VTAIL.n416 VSUBS 0.01244f
C539 VTAIL.n417 VSUBS 0.02315f
C540 VTAIL.n418 VSUBS 0.02315f
C541 VTAIL.n419 VSUBS 0.01244f
C542 VTAIL.n420 VSUBS 0.013172f
C543 VTAIL.n421 VSUBS 0.029403f
C544 VTAIL.n422 VSUBS 0.029403f
C545 VTAIL.n423 VSUBS 0.013172f
C546 VTAIL.n424 VSUBS 0.01244f
C547 VTAIL.n425 VSUBS 0.02315f
C548 VTAIL.n426 VSUBS 0.02315f
C549 VTAIL.n427 VSUBS 0.01244f
C550 VTAIL.n428 VSUBS 0.013172f
C551 VTAIL.n429 VSUBS 0.029403f
C552 VTAIL.n430 VSUBS 0.029403f
C553 VTAIL.n431 VSUBS 0.013172f
C554 VTAIL.n432 VSUBS 0.01244f
C555 VTAIL.n433 VSUBS 0.02315f
C556 VTAIL.n434 VSUBS 0.02315f
C557 VTAIL.n435 VSUBS 0.01244f
C558 VTAIL.n436 VSUBS 0.013172f
C559 VTAIL.n437 VSUBS 0.029403f
C560 VTAIL.n438 VSUBS 0.07152f
C561 VTAIL.n439 VSUBS 0.013172f
C562 VTAIL.n440 VSUBS 0.01244f
C563 VTAIL.n441 VSUBS 0.051612f
C564 VTAIL.n442 VSUBS 0.035923f
C565 VTAIL.n443 VSUBS 1.91894f
C566 VTAIL.t5 VSUBS 0.358924f
C567 VTAIL.t4 VSUBS 0.358924f
C568 VTAIL.n444 VSUBS 2.85185f
C569 VTAIL.n445 VSUBS 0.914901f
C570 VTAIL.n446 VSUBS 0.025536f
C571 VTAIL.n447 VSUBS 0.02315f
C572 VTAIL.n448 VSUBS 0.01244f
C573 VTAIL.n449 VSUBS 0.029403f
C574 VTAIL.n450 VSUBS 0.013172f
C575 VTAIL.n451 VSUBS 0.02315f
C576 VTAIL.n452 VSUBS 0.01244f
C577 VTAIL.n453 VSUBS 0.029403f
C578 VTAIL.n454 VSUBS 0.013172f
C579 VTAIL.n455 VSUBS 0.02315f
C580 VTAIL.n456 VSUBS 0.01244f
C581 VTAIL.n457 VSUBS 0.029403f
C582 VTAIL.n458 VSUBS 0.012806f
C583 VTAIL.n459 VSUBS 0.02315f
C584 VTAIL.n460 VSUBS 0.012806f
C585 VTAIL.n461 VSUBS 0.01244f
C586 VTAIL.n462 VSUBS 0.029403f
C587 VTAIL.n463 VSUBS 0.029403f
C588 VTAIL.n464 VSUBS 0.013172f
C589 VTAIL.n465 VSUBS 0.02315f
C590 VTAIL.n466 VSUBS 0.01244f
C591 VTAIL.n467 VSUBS 0.029403f
C592 VTAIL.n468 VSUBS 0.013172f
C593 VTAIL.n469 VSUBS 0.02315f
C594 VTAIL.n470 VSUBS 0.01244f
C595 VTAIL.n471 VSUBS 0.029403f
C596 VTAIL.n472 VSUBS 0.013172f
C597 VTAIL.n473 VSUBS 0.02315f
C598 VTAIL.n474 VSUBS 0.01244f
C599 VTAIL.n475 VSUBS 0.029403f
C600 VTAIL.n476 VSUBS 0.013172f
C601 VTAIL.n477 VSUBS 0.02315f
C602 VTAIL.n478 VSUBS 0.01244f
C603 VTAIL.n479 VSUBS 0.029403f
C604 VTAIL.n480 VSUBS 0.013172f
C605 VTAIL.n481 VSUBS 1.9637f
C606 VTAIL.n482 VSUBS 0.01244f
C607 VTAIL.t6 VSUBS 0.063212f
C608 VTAIL.n483 VSUBS 0.194733f
C609 VTAIL.n484 VSUBS 0.018705f
C610 VTAIL.n485 VSUBS 0.022052f
C611 VTAIL.n486 VSUBS 0.029403f
C612 VTAIL.n487 VSUBS 0.013172f
C613 VTAIL.n488 VSUBS 0.01244f
C614 VTAIL.n489 VSUBS 0.02315f
C615 VTAIL.n490 VSUBS 0.02315f
C616 VTAIL.n491 VSUBS 0.01244f
C617 VTAIL.n492 VSUBS 0.013172f
C618 VTAIL.n493 VSUBS 0.029403f
C619 VTAIL.n494 VSUBS 0.029403f
C620 VTAIL.n495 VSUBS 0.013172f
C621 VTAIL.n496 VSUBS 0.01244f
C622 VTAIL.n497 VSUBS 0.02315f
C623 VTAIL.n498 VSUBS 0.02315f
C624 VTAIL.n499 VSUBS 0.01244f
C625 VTAIL.n500 VSUBS 0.013172f
C626 VTAIL.n501 VSUBS 0.029403f
C627 VTAIL.n502 VSUBS 0.029403f
C628 VTAIL.n503 VSUBS 0.013172f
C629 VTAIL.n504 VSUBS 0.01244f
C630 VTAIL.n505 VSUBS 0.02315f
C631 VTAIL.n506 VSUBS 0.02315f
C632 VTAIL.n507 VSUBS 0.01244f
C633 VTAIL.n508 VSUBS 0.013172f
C634 VTAIL.n509 VSUBS 0.029403f
C635 VTAIL.n510 VSUBS 0.029403f
C636 VTAIL.n511 VSUBS 0.013172f
C637 VTAIL.n512 VSUBS 0.01244f
C638 VTAIL.n513 VSUBS 0.02315f
C639 VTAIL.n514 VSUBS 0.02315f
C640 VTAIL.n515 VSUBS 0.01244f
C641 VTAIL.n516 VSUBS 0.013172f
C642 VTAIL.n517 VSUBS 0.029403f
C643 VTAIL.n518 VSUBS 0.029403f
C644 VTAIL.n519 VSUBS 0.013172f
C645 VTAIL.n520 VSUBS 0.01244f
C646 VTAIL.n521 VSUBS 0.02315f
C647 VTAIL.n522 VSUBS 0.02315f
C648 VTAIL.n523 VSUBS 0.01244f
C649 VTAIL.n524 VSUBS 0.013172f
C650 VTAIL.n525 VSUBS 0.029403f
C651 VTAIL.n526 VSUBS 0.029403f
C652 VTAIL.n527 VSUBS 0.013172f
C653 VTAIL.n528 VSUBS 0.01244f
C654 VTAIL.n529 VSUBS 0.02315f
C655 VTAIL.n530 VSUBS 0.02315f
C656 VTAIL.n531 VSUBS 0.01244f
C657 VTAIL.n532 VSUBS 0.013172f
C658 VTAIL.n533 VSUBS 0.029403f
C659 VTAIL.n534 VSUBS 0.029403f
C660 VTAIL.n535 VSUBS 0.013172f
C661 VTAIL.n536 VSUBS 0.01244f
C662 VTAIL.n537 VSUBS 0.02315f
C663 VTAIL.n538 VSUBS 0.02315f
C664 VTAIL.n539 VSUBS 0.01244f
C665 VTAIL.n540 VSUBS 0.013172f
C666 VTAIL.n541 VSUBS 0.029403f
C667 VTAIL.n542 VSUBS 0.029403f
C668 VTAIL.n543 VSUBS 0.013172f
C669 VTAIL.n544 VSUBS 0.01244f
C670 VTAIL.n545 VSUBS 0.02315f
C671 VTAIL.n546 VSUBS 0.02315f
C672 VTAIL.n547 VSUBS 0.01244f
C673 VTAIL.n548 VSUBS 0.013172f
C674 VTAIL.n549 VSUBS 0.029403f
C675 VTAIL.n550 VSUBS 0.07152f
C676 VTAIL.n551 VSUBS 0.013172f
C677 VTAIL.n552 VSUBS 0.01244f
C678 VTAIL.n553 VSUBS 0.051612f
C679 VTAIL.n554 VSUBS 0.035923f
C680 VTAIL.n555 VSUBS 0.215798f
C681 VTAIL.n556 VSUBS 0.025536f
C682 VTAIL.n557 VSUBS 0.02315f
C683 VTAIL.n558 VSUBS 0.01244f
C684 VTAIL.n559 VSUBS 0.029403f
C685 VTAIL.n560 VSUBS 0.013172f
C686 VTAIL.n561 VSUBS 0.02315f
C687 VTAIL.n562 VSUBS 0.01244f
C688 VTAIL.n563 VSUBS 0.029403f
C689 VTAIL.n564 VSUBS 0.013172f
C690 VTAIL.n565 VSUBS 0.02315f
C691 VTAIL.n566 VSUBS 0.01244f
C692 VTAIL.n567 VSUBS 0.029403f
C693 VTAIL.n568 VSUBS 0.012806f
C694 VTAIL.n569 VSUBS 0.02315f
C695 VTAIL.n570 VSUBS 0.012806f
C696 VTAIL.n571 VSUBS 0.01244f
C697 VTAIL.n572 VSUBS 0.029403f
C698 VTAIL.n573 VSUBS 0.029403f
C699 VTAIL.n574 VSUBS 0.013172f
C700 VTAIL.n575 VSUBS 0.02315f
C701 VTAIL.n576 VSUBS 0.01244f
C702 VTAIL.n577 VSUBS 0.029403f
C703 VTAIL.n578 VSUBS 0.013172f
C704 VTAIL.n579 VSUBS 0.02315f
C705 VTAIL.n580 VSUBS 0.01244f
C706 VTAIL.n581 VSUBS 0.029403f
C707 VTAIL.n582 VSUBS 0.013172f
C708 VTAIL.n583 VSUBS 0.02315f
C709 VTAIL.n584 VSUBS 0.01244f
C710 VTAIL.n585 VSUBS 0.029403f
C711 VTAIL.n586 VSUBS 0.013172f
C712 VTAIL.n587 VSUBS 0.02315f
C713 VTAIL.n588 VSUBS 0.01244f
C714 VTAIL.n589 VSUBS 0.029403f
C715 VTAIL.n590 VSUBS 0.013172f
C716 VTAIL.n591 VSUBS 1.9637f
C717 VTAIL.n592 VSUBS 0.01244f
C718 VTAIL.t8 VSUBS 0.063212f
C719 VTAIL.n593 VSUBS 0.194733f
C720 VTAIL.n594 VSUBS 0.018705f
C721 VTAIL.n595 VSUBS 0.022052f
C722 VTAIL.n596 VSUBS 0.029403f
C723 VTAIL.n597 VSUBS 0.013172f
C724 VTAIL.n598 VSUBS 0.01244f
C725 VTAIL.n599 VSUBS 0.02315f
C726 VTAIL.n600 VSUBS 0.02315f
C727 VTAIL.n601 VSUBS 0.01244f
C728 VTAIL.n602 VSUBS 0.013172f
C729 VTAIL.n603 VSUBS 0.029403f
C730 VTAIL.n604 VSUBS 0.029403f
C731 VTAIL.n605 VSUBS 0.013172f
C732 VTAIL.n606 VSUBS 0.01244f
C733 VTAIL.n607 VSUBS 0.02315f
C734 VTAIL.n608 VSUBS 0.02315f
C735 VTAIL.n609 VSUBS 0.01244f
C736 VTAIL.n610 VSUBS 0.013172f
C737 VTAIL.n611 VSUBS 0.029403f
C738 VTAIL.n612 VSUBS 0.029403f
C739 VTAIL.n613 VSUBS 0.013172f
C740 VTAIL.n614 VSUBS 0.01244f
C741 VTAIL.n615 VSUBS 0.02315f
C742 VTAIL.n616 VSUBS 0.02315f
C743 VTAIL.n617 VSUBS 0.01244f
C744 VTAIL.n618 VSUBS 0.013172f
C745 VTAIL.n619 VSUBS 0.029403f
C746 VTAIL.n620 VSUBS 0.029403f
C747 VTAIL.n621 VSUBS 0.013172f
C748 VTAIL.n622 VSUBS 0.01244f
C749 VTAIL.n623 VSUBS 0.02315f
C750 VTAIL.n624 VSUBS 0.02315f
C751 VTAIL.n625 VSUBS 0.01244f
C752 VTAIL.n626 VSUBS 0.013172f
C753 VTAIL.n627 VSUBS 0.029403f
C754 VTAIL.n628 VSUBS 0.029403f
C755 VTAIL.n629 VSUBS 0.013172f
C756 VTAIL.n630 VSUBS 0.01244f
C757 VTAIL.n631 VSUBS 0.02315f
C758 VTAIL.n632 VSUBS 0.02315f
C759 VTAIL.n633 VSUBS 0.01244f
C760 VTAIL.n634 VSUBS 0.013172f
C761 VTAIL.n635 VSUBS 0.029403f
C762 VTAIL.n636 VSUBS 0.029403f
C763 VTAIL.n637 VSUBS 0.013172f
C764 VTAIL.n638 VSUBS 0.01244f
C765 VTAIL.n639 VSUBS 0.02315f
C766 VTAIL.n640 VSUBS 0.02315f
C767 VTAIL.n641 VSUBS 0.01244f
C768 VTAIL.n642 VSUBS 0.013172f
C769 VTAIL.n643 VSUBS 0.029403f
C770 VTAIL.n644 VSUBS 0.029403f
C771 VTAIL.n645 VSUBS 0.013172f
C772 VTAIL.n646 VSUBS 0.01244f
C773 VTAIL.n647 VSUBS 0.02315f
C774 VTAIL.n648 VSUBS 0.02315f
C775 VTAIL.n649 VSUBS 0.01244f
C776 VTAIL.n650 VSUBS 0.013172f
C777 VTAIL.n651 VSUBS 0.029403f
C778 VTAIL.n652 VSUBS 0.029403f
C779 VTAIL.n653 VSUBS 0.013172f
C780 VTAIL.n654 VSUBS 0.01244f
C781 VTAIL.n655 VSUBS 0.02315f
C782 VTAIL.n656 VSUBS 0.02315f
C783 VTAIL.n657 VSUBS 0.01244f
C784 VTAIL.n658 VSUBS 0.013172f
C785 VTAIL.n659 VSUBS 0.029403f
C786 VTAIL.n660 VSUBS 0.07152f
C787 VTAIL.n661 VSUBS 0.013172f
C788 VTAIL.n662 VSUBS 0.01244f
C789 VTAIL.n663 VSUBS 0.051612f
C790 VTAIL.n664 VSUBS 0.035923f
C791 VTAIL.n665 VSUBS 0.215798f
C792 VTAIL.t14 VSUBS 0.358924f
C793 VTAIL.t10 VSUBS 0.358924f
C794 VTAIL.n666 VSUBS 2.85185f
C795 VTAIL.n667 VSUBS 0.914901f
C796 VTAIL.n668 VSUBS 0.025536f
C797 VTAIL.n669 VSUBS 0.02315f
C798 VTAIL.n670 VSUBS 0.01244f
C799 VTAIL.n671 VSUBS 0.029403f
C800 VTAIL.n672 VSUBS 0.013172f
C801 VTAIL.n673 VSUBS 0.02315f
C802 VTAIL.n674 VSUBS 0.01244f
C803 VTAIL.n675 VSUBS 0.029403f
C804 VTAIL.n676 VSUBS 0.013172f
C805 VTAIL.n677 VSUBS 0.02315f
C806 VTAIL.n678 VSUBS 0.01244f
C807 VTAIL.n679 VSUBS 0.029403f
C808 VTAIL.n680 VSUBS 0.012806f
C809 VTAIL.n681 VSUBS 0.02315f
C810 VTAIL.n682 VSUBS 0.012806f
C811 VTAIL.n683 VSUBS 0.01244f
C812 VTAIL.n684 VSUBS 0.029403f
C813 VTAIL.n685 VSUBS 0.029403f
C814 VTAIL.n686 VSUBS 0.013172f
C815 VTAIL.n687 VSUBS 0.02315f
C816 VTAIL.n688 VSUBS 0.01244f
C817 VTAIL.n689 VSUBS 0.029403f
C818 VTAIL.n690 VSUBS 0.013172f
C819 VTAIL.n691 VSUBS 0.02315f
C820 VTAIL.n692 VSUBS 0.01244f
C821 VTAIL.n693 VSUBS 0.029403f
C822 VTAIL.n694 VSUBS 0.013172f
C823 VTAIL.n695 VSUBS 0.02315f
C824 VTAIL.n696 VSUBS 0.01244f
C825 VTAIL.n697 VSUBS 0.029403f
C826 VTAIL.n698 VSUBS 0.013172f
C827 VTAIL.n699 VSUBS 0.02315f
C828 VTAIL.n700 VSUBS 0.01244f
C829 VTAIL.n701 VSUBS 0.029403f
C830 VTAIL.n702 VSUBS 0.013172f
C831 VTAIL.n703 VSUBS 1.9637f
C832 VTAIL.n704 VSUBS 0.01244f
C833 VTAIL.t9 VSUBS 0.063212f
C834 VTAIL.n705 VSUBS 0.194733f
C835 VTAIL.n706 VSUBS 0.018705f
C836 VTAIL.n707 VSUBS 0.022052f
C837 VTAIL.n708 VSUBS 0.029403f
C838 VTAIL.n709 VSUBS 0.013172f
C839 VTAIL.n710 VSUBS 0.01244f
C840 VTAIL.n711 VSUBS 0.02315f
C841 VTAIL.n712 VSUBS 0.02315f
C842 VTAIL.n713 VSUBS 0.01244f
C843 VTAIL.n714 VSUBS 0.013172f
C844 VTAIL.n715 VSUBS 0.029403f
C845 VTAIL.n716 VSUBS 0.029403f
C846 VTAIL.n717 VSUBS 0.013172f
C847 VTAIL.n718 VSUBS 0.01244f
C848 VTAIL.n719 VSUBS 0.02315f
C849 VTAIL.n720 VSUBS 0.02315f
C850 VTAIL.n721 VSUBS 0.01244f
C851 VTAIL.n722 VSUBS 0.013172f
C852 VTAIL.n723 VSUBS 0.029403f
C853 VTAIL.n724 VSUBS 0.029403f
C854 VTAIL.n725 VSUBS 0.013172f
C855 VTAIL.n726 VSUBS 0.01244f
C856 VTAIL.n727 VSUBS 0.02315f
C857 VTAIL.n728 VSUBS 0.02315f
C858 VTAIL.n729 VSUBS 0.01244f
C859 VTAIL.n730 VSUBS 0.013172f
C860 VTAIL.n731 VSUBS 0.029403f
C861 VTAIL.n732 VSUBS 0.029403f
C862 VTAIL.n733 VSUBS 0.013172f
C863 VTAIL.n734 VSUBS 0.01244f
C864 VTAIL.n735 VSUBS 0.02315f
C865 VTAIL.n736 VSUBS 0.02315f
C866 VTAIL.n737 VSUBS 0.01244f
C867 VTAIL.n738 VSUBS 0.013172f
C868 VTAIL.n739 VSUBS 0.029403f
C869 VTAIL.n740 VSUBS 0.029403f
C870 VTAIL.n741 VSUBS 0.013172f
C871 VTAIL.n742 VSUBS 0.01244f
C872 VTAIL.n743 VSUBS 0.02315f
C873 VTAIL.n744 VSUBS 0.02315f
C874 VTAIL.n745 VSUBS 0.01244f
C875 VTAIL.n746 VSUBS 0.013172f
C876 VTAIL.n747 VSUBS 0.029403f
C877 VTAIL.n748 VSUBS 0.029403f
C878 VTAIL.n749 VSUBS 0.013172f
C879 VTAIL.n750 VSUBS 0.01244f
C880 VTAIL.n751 VSUBS 0.02315f
C881 VTAIL.n752 VSUBS 0.02315f
C882 VTAIL.n753 VSUBS 0.01244f
C883 VTAIL.n754 VSUBS 0.013172f
C884 VTAIL.n755 VSUBS 0.029403f
C885 VTAIL.n756 VSUBS 0.029403f
C886 VTAIL.n757 VSUBS 0.013172f
C887 VTAIL.n758 VSUBS 0.01244f
C888 VTAIL.n759 VSUBS 0.02315f
C889 VTAIL.n760 VSUBS 0.02315f
C890 VTAIL.n761 VSUBS 0.01244f
C891 VTAIL.n762 VSUBS 0.013172f
C892 VTAIL.n763 VSUBS 0.029403f
C893 VTAIL.n764 VSUBS 0.029403f
C894 VTAIL.n765 VSUBS 0.013172f
C895 VTAIL.n766 VSUBS 0.01244f
C896 VTAIL.n767 VSUBS 0.02315f
C897 VTAIL.n768 VSUBS 0.02315f
C898 VTAIL.n769 VSUBS 0.01244f
C899 VTAIL.n770 VSUBS 0.013172f
C900 VTAIL.n771 VSUBS 0.029403f
C901 VTAIL.n772 VSUBS 0.07152f
C902 VTAIL.n773 VSUBS 0.013172f
C903 VTAIL.n774 VSUBS 0.01244f
C904 VTAIL.n775 VSUBS 0.051612f
C905 VTAIL.n776 VSUBS 0.035923f
C906 VTAIL.n777 VSUBS 1.91894f
C907 VTAIL.n778 VSUBS 0.025536f
C908 VTAIL.n779 VSUBS 0.02315f
C909 VTAIL.n780 VSUBS 0.01244f
C910 VTAIL.n781 VSUBS 0.029403f
C911 VTAIL.n782 VSUBS 0.013172f
C912 VTAIL.n783 VSUBS 0.02315f
C913 VTAIL.n784 VSUBS 0.01244f
C914 VTAIL.n785 VSUBS 0.029403f
C915 VTAIL.n786 VSUBS 0.013172f
C916 VTAIL.n787 VSUBS 0.02315f
C917 VTAIL.n788 VSUBS 0.01244f
C918 VTAIL.n789 VSUBS 0.029403f
C919 VTAIL.n790 VSUBS 0.012806f
C920 VTAIL.n791 VSUBS 0.02315f
C921 VTAIL.n792 VSUBS 0.013172f
C922 VTAIL.n793 VSUBS 0.029403f
C923 VTAIL.n794 VSUBS 0.013172f
C924 VTAIL.n795 VSUBS 0.02315f
C925 VTAIL.n796 VSUBS 0.01244f
C926 VTAIL.n797 VSUBS 0.029403f
C927 VTAIL.n798 VSUBS 0.013172f
C928 VTAIL.n799 VSUBS 0.02315f
C929 VTAIL.n800 VSUBS 0.01244f
C930 VTAIL.n801 VSUBS 0.029403f
C931 VTAIL.n802 VSUBS 0.013172f
C932 VTAIL.n803 VSUBS 0.02315f
C933 VTAIL.n804 VSUBS 0.01244f
C934 VTAIL.n805 VSUBS 0.029403f
C935 VTAIL.n806 VSUBS 0.013172f
C936 VTAIL.n807 VSUBS 0.02315f
C937 VTAIL.n808 VSUBS 0.01244f
C938 VTAIL.n809 VSUBS 0.029403f
C939 VTAIL.n810 VSUBS 0.013172f
C940 VTAIL.n811 VSUBS 1.9637f
C941 VTAIL.n812 VSUBS 0.01244f
C942 VTAIL.t0 VSUBS 0.063212f
C943 VTAIL.n813 VSUBS 0.194733f
C944 VTAIL.n814 VSUBS 0.018705f
C945 VTAIL.n815 VSUBS 0.022052f
C946 VTAIL.n816 VSUBS 0.029403f
C947 VTAIL.n817 VSUBS 0.013172f
C948 VTAIL.n818 VSUBS 0.01244f
C949 VTAIL.n819 VSUBS 0.02315f
C950 VTAIL.n820 VSUBS 0.02315f
C951 VTAIL.n821 VSUBS 0.01244f
C952 VTAIL.n822 VSUBS 0.013172f
C953 VTAIL.n823 VSUBS 0.029403f
C954 VTAIL.n824 VSUBS 0.029403f
C955 VTAIL.n825 VSUBS 0.013172f
C956 VTAIL.n826 VSUBS 0.01244f
C957 VTAIL.n827 VSUBS 0.02315f
C958 VTAIL.n828 VSUBS 0.02315f
C959 VTAIL.n829 VSUBS 0.01244f
C960 VTAIL.n830 VSUBS 0.013172f
C961 VTAIL.n831 VSUBS 0.029403f
C962 VTAIL.n832 VSUBS 0.029403f
C963 VTAIL.n833 VSUBS 0.013172f
C964 VTAIL.n834 VSUBS 0.01244f
C965 VTAIL.n835 VSUBS 0.02315f
C966 VTAIL.n836 VSUBS 0.02315f
C967 VTAIL.n837 VSUBS 0.01244f
C968 VTAIL.n838 VSUBS 0.013172f
C969 VTAIL.n839 VSUBS 0.029403f
C970 VTAIL.n840 VSUBS 0.029403f
C971 VTAIL.n841 VSUBS 0.013172f
C972 VTAIL.n842 VSUBS 0.01244f
C973 VTAIL.n843 VSUBS 0.02315f
C974 VTAIL.n844 VSUBS 0.02315f
C975 VTAIL.n845 VSUBS 0.01244f
C976 VTAIL.n846 VSUBS 0.013172f
C977 VTAIL.n847 VSUBS 0.029403f
C978 VTAIL.n848 VSUBS 0.029403f
C979 VTAIL.n849 VSUBS 0.013172f
C980 VTAIL.n850 VSUBS 0.01244f
C981 VTAIL.n851 VSUBS 0.02315f
C982 VTAIL.n852 VSUBS 0.02315f
C983 VTAIL.n853 VSUBS 0.01244f
C984 VTAIL.n854 VSUBS 0.01244f
C985 VTAIL.n855 VSUBS 0.013172f
C986 VTAIL.n856 VSUBS 0.029403f
C987 VTAIL.n857 VSUBS 0.029403f
C988 VTAIL.n858 VSUBS 0.029403f
C989 VTAIL.n859 VSUBS 0.012806f
C990 VTAIL.n860 VSUBS 0.01244f
C991 VTAIL.n861 VSUBS 0.02315f
C992 VTAIL.n862 VSUBS 0.02315f
C993 VTAIL.n863 VSUBS 0.01244f
C994 VTAIL.n864 VSUBS 0.013172f
C995 VTAIL.n865 VSUBS 0.029403f
C996 VTAIL.n866 VSUBS 0.029403f
C997 VTAIL.n867 VSUBS 0.013172f
C998 VTAIL.n868 VSUBS 0.01244f
C999 VTAIL.n869 VSUBS 0.02315f
C1000 VTAIL.n870 VSUBS 0.02315f
C1001 VTAIL.n871 VSUBS 0.01244f
C1002 VTAIL.n872 VSUBS 0.013172f
C1003 VTAIL.n873 VSUBS 0.029403f
C1004 VTAIL.n874 VSUBS 0.029403f
C1005 VTAIL.n875 VSUBS 0.013172f
C1006 VTAIL.n876 VSUBS 0.01244f
C1007 VTAIL.n877 VSUBS 0.02315f
C1008 VTAIL.n878 VSUBS 0.02315f
C1009 VTAIL.n879 VSUBS 0.01244f
C1010 VTAIL.n880 VSUBS 0.013172f
C1011 VTAIL.n881 VSUBS 0.029403f
C1012 VTAIL.n882 VSUBS 0.07152f
C1013 VTAIL.n883 VSUBS 0.013172f
C1014 VTAIL.n884 VSUBS 0.01244f
C1015 VTAIL.n885 VSUBS 0.051612f
C1016 VTAIL.n886 VSUBS 0.035923f
C1017 VTAIL.n887 VSUBS 1.91459f
C1018 VP.n0 VSUBS 0.038244f
C1019 VP.t7 VSUBS 3.4339f
C1020 VP.n1 VSUBS 0.023579f
C1021 VP.n2 VSUBS 0.02901f
C1022 VP.t3 VSUBS 3.4339f
C1023 VP.n3 VSUBS 0.057353f
C1024 VP.n4 VSUBS 0.02901f
C1025 VP.t2 VSUBS 3.4339f
C1026 VP.n5 VSUBS 1.19097f
C1027 VP.n6 VSUBS 0.02901f
C1028 VP.n7 VSUBS 0.056707f
C1029 VP.n8 VSUBS 0.038244f
C1030 VP.t0 VSUBS 3.4339f
C1031 VP.n9 VSUBS 0.023579f
C1032 VP.n10 VSUBS 0.02901f
C1033 VP.t1 VSUBS 3.4339f
C1034 VP.n11 VSUBS 0.057353f
C1035 VP.n12 VSUBS 0.02901f
C1036 VP.t6 VSUBS 3.4339f
C1037 VP.n13 VSUBS 1.26564f
C1038 VP.t5 VSUBS 3.60998f
C1039 VP.n14 VSUBS 1.25638f
C1040 VP.n15 VSUBS 0.246616f
C1041 VP.n16 VSUBS 0.041048f
C1042 VP.n17 VSUBS 0.057353f
C1043 VP.n18 VSUBS 0.02343f
C1044 VP.n19 VSUBS 0.02901f
C1045 VP.n20 VSUBS 0.02901f
C1046 VP.n21 VSUBS 0.02901f
C1047 VP.n22 VSUBS 0.041048f
C1048 VP.n23 VSUBS 1.19097f
C1049 VP.n24 VSUBS 0.039986f
C1050 VP.n25 VSUBS 0.057851f
C1051 VP.n26 VSUBS 0.02901f
C1052 VP.n27 VSUBS 0.02901f
C1053 VP.n28 VSUBS 0.02901f
C1054 VP.n29 VSUBS 0.056707f
C1055 VP.n30 VSUBS 0.042111f
C1056 VP.n31 VSUBS 1.27728f
C1057 VP.n32 VSUBS 1.83109f
C1058 VP.n33 VSUBS 1.8502f
C1059 VP.t4 VSUBS 3.4339f
C1060 VP.n34 VSUBS 1.27728f
C1061 VP.n35 VSUBS 0.042111f
C1062 VP.n36 VSUBS 0.038244f
C1063 VP.n37 VSUBS 0.02901f
C1064 VP.n38 VSUBS 0.02901f
C1065 VP.n39 VSUBS 0.023579f
C1066 VP.n40 VSUBS 0.057851f
C1067 VP.n41 VSUBS 0.039986f
C1068 VP.n42 VSUBS 0.02901f
C1069 VP.n43 VSUBS 0.02901f
C1070 VP.n44 VSUBS 0.041048f
C1071 VP.n45 VSUBS 0.057353f
C1072 VP.n46 VSUBS 0.02343f
C1073 VP.n47 VSUBS 0.02901f
C1074 VP.n48 VSUBS 0.02901f
C1075 VP.n49 VSUBS 0.02901f
C1076 VP.n50 VSUBS 0.041048f
C1077 VP.n51 VSUBS 1.19097f
C1078 VP.n52 VSUBS 0.039986f
C1079 VP.n53 VSUBS 0.057851f
C1080 VP.n54 VSUBS 0.02901f
C1081 VP.n55 VSUBS 0.02901f
C1082 VP.n56 VSUBS 0.02901f
C1083 VP.n57 VSUBS 0.056707f
C1084 VP.n58 VSUBS 0.042111f
C1085 VP.n59 VSUBS 1.27728f
C1086 VP.n60 VSUBS 0.041075f
C1087 B.n0 VSUBS 0.003923f
C1088 B.n1 VSUBS 0.003923f
C1089 B.n2 VSUBS 0.006204f
C1090 B.n3 VSUBS 0.006204f
C1091 B.n4 VSUBS 0.006204f
C1092 B.n5 VSUBS 0.006204f
C1093 B.n6 VSUBS 0.006204f
C1094 B.n7 VSUBS 0.006204f
C1095 B.n8 VSUBS 0.006204f
C1096 B.n9 VSUBS 0.006204f
C1097 B.n10 VSUBS 0.006204f
C1098 B.n11 VSUBS 0.006204f
C1099 B.n12 VSUBS 0.006204f
C1100 B.n13 VSUBS 0.006204f
C1101 B.n14 VSUBS 0.006204f
C1102 B.n15 VSUBS 0.006204f
C1103 B.n16 VSUBS 0.006204f
C1104 B.n17 VSUBS 0.006204f
C1105 B.n18 VSUBS 0.006204f
C1106 B.n19 VSUBS 0.006204f
C1107 B.n20 VSUBS 0.006204f
C1108 B.n21 VSUBS 0.006204f
C1109 B.n22 VSUBS 0.006204f
C1110 B.n23 VSUBS 0.006204f
C1111 B.n24 VSUBS 0.013845f
C1112 B.n25 VSUBS 0.006204f
C1113 B.n26 VSUBS 0.006204f
C1114 B.n27 VSUBS 0.006204f
C1115 B.n28 VSUBS 0.006204f
C1116 B.n29 VSUBS 0.006204f
C1117 B.n30 VSUBS 0.006204f
C1118 B.n31 VSUBS 0.006204f
C1119 B.n32 VSUBS 0.006204f
C1120 B.n33 VSUBS 0.006204f
C1121 B.n34 VSUBS 0.006204f
C1122 B.n35 VSUBS 0.006204f
C1123 B.n36 VSUBS 0.006204f
C1124 B.n37 VSUBS 0.006204f
C1125 B.n38 VSUBS 0.006204f
C1126 B.n39 VSUBS 0.006204f
C1127 B.n40 VSUBS 0.006204f
C1128 B.n41 VSUBS 0.006204f
C1129 B.n42 VSUBS 0.006204f
C1130 B.n43 VSUBS 0.006204f
C1131 B.n44 VSUBS 0.006204f
C1132 B.n45 VSUBS 0.006204f
C1133 B.n46 VSUBS 0.006204f
C1134 B.n47 VSUBS 0.006204f
C1135 B.n48 VSUBS 0.006204f
C1136 B.n49 VSUBS 0.006204f
C1137 B.n50 VSUBS 0.006204f
C1138 B.n51 VSUBS 0.006204f
C1139 B.n52 VSUBS 0.006204f
C1140 B.n53 VSUBS 0.006204f
C1141 B.n54 VSUBS 0.006204f
C1142 B.n55 VSUBS 0.006204f
C1143 B.n56 VSUBS 0.005839f
C1144 B.n57 VSUBS 0.006204f
C1145 B.t11 VSUBS 0.346189f
C1146 B.t10 VSUBS 0.372096f
C1147 B.t9 VSUBS 1.65743f
C1148 B.n58 VSUBS 0.550047f
C1149 B.n59 VSUBS 0.306678f
C1150 B.n60 VSUBS 0.014373f
C1151 B.n61 VSUBS 0.006204f
C1152 B.n62 VSUBS 0.006204f
C1153 B.n63 VSUBS 0.006204f
C1154 B.n64 VSUBS 0.006204f
C1155 B.t2 VSUBS 0.346192f
C1156 B.t1 VSUBS 0.372099f
C1157 B.t0 VSUBS 1.65743f
C1158 B.n65 VSUBS 0.550044f
C1159 B.n66 VSUBS 0.306674f
C1160 B.n67 VSUBS 0.006204f
C1161 B.n68 VSUBS 0.006204f
C1162 B.n69 VSUBS 0.006204f
C1163 B.n70 VSUBS 0.006204f
C1164 B.n71 VSUBS 0.006204f
C1165 B.n72 VSUBS 0.006204f
C1166 B.n73 VSUBS 0.006204f
C1167 B.n74 VSUBS 0.006204f
C1168 B.n75 VSUBS 0.006204f
C1169 B.n76 VSUBS 0.006204f
C1170 B.n77 VSUBS 0.006204f
C1171 B.n78 VSUBS 0.006204f
C1172 B.n79 VSUBS 0.006204f
C1173 B.n80 VSUBS 0.006204f
C1174 B.n81 VSUBS 0.006204f
C1175 B.n82 VSUBS 0.006204f
C1176 B.n83 VSUBS 0.006204f
C1177 B.n84 VSUBS 0.006204f
C1178 B.n85 VSUBS 0.006204f
C1179 B.n86 VSUBS 0.006204f
C1180 B.n87 VSUBS 0.006204f
C1181 B.n88 VSUBS 0.006204f
C1182 B.n89 VSUBS 0.006204f
C1183 B.n90 VSUBS 0.006204f
C1184 B.n91 VSUBS 0.006204f
C1185 B.n92 VSUBS 0.006204f
C1186 B.n93 VSUBS 0.006204f
C1187 B.n94 VSUBS 0.006204f
C1188 B.n95 VSUBS 0.006204f
C1189 B.n96 VSUBS 0.006204f
C1190 B.n97 VSUBS 0.006204f
C1191 B.n98 VSUBS 0.014984f
C1192 B.n99 VSUBS 0.006204f
C1193 B.n100 VSUBS 0.006204f
C1194 B.n101 VSUBS 0.006204f
C1195 B.n102 VSUBS 0.006204f
C1196 B.n103 VSUBS 0.006204f
C1197 B.n104 VSUBS 0.006204f
C1198 B.n105 VSUBS 0.006204f
C1199 B.n106 VSUBS 0.006204f
C1200 B.n107 VSUBS 0.006204f
C1201 B.n108 VSUBS 0.006204f
C1202 B.n109 VSUBS 0.006204f
C1203 B.n110 VSUBS 0.006204f
C1204 B.n111 VSUBS 0.006204f
C1205 B.n112 VSUBS 0.006204f
C1206 B.n113 VSUBS 0.006204f
C1207 B.n114 VSUBS 0.006204f
C1208 B.n115 VSUBS 0.006204f
C1209 B.n116 VSUBS 0.006204f
C1210 B.n117 VSUBS 0.006204f
C1211 B.n118 VSUBS 0.006204f
C1212 B.n119 VSUBS 0.006204f
C1213 B.n120 VSUBS 0.006204f
C1214 B.n121 VSUBS 0.006204f
C1215 B.n122 VSUBS 0.006204f
C1216 B.n123 VSUBS 0.006204f
C1217 B.n124 VSUBS 0.006204f
C1218 B.n125 VSUBS 0.006204f
C1219 B.n126 VSUBS 0.006204f
C1220 B.n127 VSUBS 0.006204f
C1221 B.n128 VSUBS 0.006204f
C1222 B.n129 VSUBS 0.006204f
C1223 B.n130 VSUBS 0.006204f
C1224 B.n131 VSUBS 0.006204f
C1225 B.n132 VSUBS 0.006204f
C1226 B.n133 VSUBS 0.006204f
C1227 B.n134 VSUBS 0.006204f
C1228 B.n135 VSUBS 0.006204f
C1229 B.n136 VSUBS 0.006204f
C1230 B.n137 VSUBS 0.006204f
C1231 B.n138 VSUBS 0.006204f
C1232 B.n139 VSUBS 0.006204f
C1233 B.n140 VSUBS 0.006204f
C1234 B.n141 VSUBS 0.006204f
C1235 B.n142 VSUBS 0.006204f
C1236 B.n143 VSUBS 0.006204f
C1237 B.n144 VSUBS 0.014984f
C1238 B.n145 VSUBS 0.006204f
C1239 B.n146 VSUBS 0.006204f
C1240 B.n147 VSUBS 0.006204f
C1241 B.n148 VSUBS 0.006204f
C1242 B.n149 VSUBS 0.006204f
C1243 B.n150 VSUBS 0.006204f
C1244 B.n151 VSUBS 0.006204f
C1245 B.n152 VSUBS 0.006204f
C1246 B.n153 VSUBS 0.006204f
C1247 B.n154 VSUBS 0.006204f
C1248 B.n155 VSUBS 0.006204f
C1249 B.n156 VSUBS 0.006204f
C1250 B.n157 VSUBS 0.006204f
C1251 B.n158 VSUBS 0.006204f
C1252 B.n159 VSUBS 0.006204f
C1253 B.n160 VSUBS 0.006204f
C1254 B.n161 VSUBS 0.006204f
C1255 B.n162 VSUBS 0.006204f
C1256 B.n163 VSUBS 0.006204f
C1257 B.n164 VSUBS 0.006204f
C1258 B.n165 VSUBS 0.006204f
C1259 B.n166 VSUBS 0.006204f
C1260 B.n167 VSUBS 0.006204f
C1261 B.n168 VSUBS 0.006204f
C1262 B.n169 VSUBS 0.006204f
C1263 B.n170 VSUBS 0.006204f
C1264 B.n171 VSUBS 0.006204f
C1265 B.n172 VSUBS 0.006204f
C1266 B.n173 VSUBS 0.006204f
C1267 B.n174 VSUBS 0.006204f
C1268 B.n175 VSUBS 0.006204f
C1269 B.n176 VSUBS 0.006204f
C1270 B.t4 VSUBS 0.346192f
C1271 B.t5 VSUBS 0.372099f
C1272 B.t3 VSUBS 1.65743f
C1273 B.n177 VSUBS 0.550044f
C1274 B.n178 VSUBS 0.306674f
C1275 B.n179 VSUBS 0.006204f
C1276 B.n180 VSUBS 0.006204f
C1277 B.n181 VSUBS 0.006204f
C1278 B.n182 VSUBS 0.006204f
C1279 B.t7 VSUBS 0.346189f
C1280 B.t8 VSUBS 0.372096f
C1281 B.t6 VSUBS 1.65743f
C1282 B.n183 VSUBS 0.550047f
C1283 B.n184 VSUBS 0.306678f
C1284 B.n185 VSUBS 0.014373f
C1285 B.n186 VSUBS 0.006204f
C1286 B.n187 VSUBS 0.006204f
C1287 B.n188 VSUBS 0.006204f
C1288 B.n189 VSUBS 0.006204f
C1289 B.n190 VSUBS 0.006204f
C1290 B.n191 VSUBS 0.006204f
C1291 B.n192 VSUBS 0.006204f
C1292 B.n193 VSUBS 0.006204f
C1293 B.n194 VSUBS 0.006204f
C1294 B.n195 VSUBS 0.006204f
C1295 B.n196 VSUBS 0.006204f
C1296 B.n197 VSUBS 0.006204f
C1297 B.n198 VSUBS 0.006204f
C1298 B.n199 VSUBS 0.006204f
C1299 B.n200 VSUBS 0.006204f
C1300 B.n201 VSUBS 0.006204f
C1301 B.n202 VSUBS 0.006204f
C1302 B.n203 VSUBS 0.006204f
C1303 B.n204 VSUBS 0.006204f
C1304 B.n205 VSUBS 0.006204f
C1305 B.n206 VSUBS 0.006204f
C1306 B.n207 VSUBS 0.006204f
C1307 B.n208 VSUBS 0.006204f
C1308 B.n209 VSUBS 0.006204f
C1309 B.n210 VSUBS 0.006204f
C1310 B.n211 VSUBS 0.006204f
C1311 B.n212 VSUBS 0.006204f
C1312 B.n213 VSUBS 0.006204f
C1313 B.n214 VSUBS 0.006204f
C1314 B.n215 VSUBS 0.006204f
C1315 B.n216 VSUBS 0.006204f
C1316 B.n217 VSUBS 0.014984f
C1317 B.n218 VSUBS 0.006204f
C1318 B.n219 VSUBS 0.006204f
C1319 B.n220 VSUBS 0.006204f
C1320 B.n221 VSUBS 0.006204f
C1321 B.n222 VSUBS 0.006204f
C1322 B.n223 VSUBS 0.006204f
C1323 B.n224 VSUBS 0.006204f
C1324 B.n225 VSUBS 0.006204f
C1325 B.n226 VSUBS 0.006204f
C1326 B.n227 VSUBS 0.006204f
C1327 B.n228 VSUBS 0.006204f
C1328 B.n229 VSUBS 0.006204f
C1329 B.n230 VSUBS 0.006204f
C1330 B.n231 VSUBS 0.006204f
C1331 B.n232 VSUBS 0.006204f
C1332 B.n233 VSUBS 0.006204f
C1333 B.n234 VSUBS 0.006204f
C1334 B.n235 VSUBS 0.006204f
C1335 B.n236 VSUBS 0.006204f
C1336 B.n237 VSUBS 0.006204f
C1337 B.n238 VSUBS 0.006204f
C1338 B.n239 VSUBS 0.006204f
C1339 B.n240 VSUBS 0.006204f
C1340 B.n241 VSUBS 0.006204f
C1341 B.n242 VSUBS 0.006204f
C1342 B.n243 VSUBS 0.006204f
C1343 B.n244 VSUBS 0.006204f
C1344 B.n245 VSUBS 0.006204f
C1345 B.n246 VSUBS 0.006204f
C1346 B.n247 VSUBS 0.006204f
C1347 B.n248 VSUBS 0.006204f
C1348 B.n249 VSUBS 0.006204f
C1349 B.n250 VSUBS 0.006204f
C1350 B.n251 VSUBS 0.006204f
C1351 B.n252 VSUBS 0.006204f
C1352 B.n253 VSUBS 0.006204f
C1353 B.n254 VSUBS 0.006204f
C1354 B.n255 VSUBS 0.006204f
C1355 B.n256 VSUBS 0.006204f
C1356 B.n257 VSUBS 0.006204f
C1357 B.n258 VSUBS 0.006204f
C1358 B.n259 VSUBS 0.006204f
C1359 B.n260 VSUBS 0.006204f
C1360 B.n261 VSUBS 0.006204f
C1361 B.n262 VSUBS 0.006204f
C1362 B.n263 VSUBS 0.006204f
C1363 B.n264 VSUBS 0.006204f
C1364 B.n265 VSUBS 0.006204f
C1365 B.n266 VSUBS 0.006204f
C1366 B.n267 VSUBS 0.006204f
C1367 B.n268 VSUBS 0.006204f
C1368 B.n269 VSUBS 0.006204f
C1369 B.n270 VSUBS 0.006204f
C1370 B.n271 VSUBS 0.006204f
C1371 B.n272 VSUBS 0.006204f
C1372 B.n273 VSUBS 0.006204f
C1373 B.n274 VSUBS 0.006204f
C1374 B.n275 VSUBS 0.006204f
C1375 B.n276 VSUBS 0.006204f
C1376 B.n277 VSUBS 0.006204f
C1377 B.n278 VSUBS 0.006204f
C1378 B.n279 VSUBS 0.006204f
C1379 B.n280 VSUBS 0.006204f
C1380 B.n281 VSUBS 0.006204f
C1381 B.n282 VSUBS 0.006204f
C1382 B.n283 VSUBS 0.006204f
C1383 B.n284 VSUBS 0.006204f
C1384 B.n285 VSUBS 0.006204f
C1385 B.n286 VSUBS 0.006204f
C1386 B.n287 VSUBS 0.006204f
C1387 B.n288 VSUBS 0.006204f
C1388 B.n289 VSUBS 0.006204f
C1389 B.n290 VSUBS 0.006204f
C1390 B.n291 VSUBS 0.006204f
C1391 B.n292 VSUBS 0.006204f
C1392 B.n293 VSUBS 0.006204f
C1393 B.n294 VSUBS 0.006204f
C1394 B.n295 VSUBS 0.006204f
C1395 B.n296 VSUBS 0.006204f
C1396 B.n297 VSUBS 0.006204f
C1397 B.n298 VSUBS 0.006204f
C1398 B.n299 VSUBS 0.006204f
C1399 B.n300 VSUBS 0.006204f
C1400 B.n301 VSUBS 0.006204f
C1401 B.n302 VSUBS 0.006204f
C1402 B.n303 VSUBS 0.006204f
C1403 B.n304 VSUBS 0.013845f
C1404 B.n305 VSUBS 0.013845f
C1405 B.n306 VSUBS 0.014984f
C1406 B.n307 VSUBS 0.006204f
C1407 B.n308 VSUBS 0.006204f
C1408 B.n309 VSUBS 0.006204f
C1409 B.n310 VSUBS 0.006204f
C1410 B.n311 VSUBS 0.006204f
C1411 B.n312 VSUBS 0.006204f
C1412 B.n313 VSUBS 0.006204f
C1413 B.n314 VSUBS 0.006204f
C1414 B.n315 VSUBS 0.006204f
C1415 B.n316 VSUBS 0.006204f
C1416 B.n317 VSUBS 0.006204f
C1417 B.n318 VSUBS 0.006204f
C1418 B.n319 VSUBS 0.006204f
C1419 B.n320 VSUBS 0.006204f
C1420 B.n321 VSUBS 0.006204f
C1421 B.n322 VSUBS 0.006204f
C1422 B.n323 VSUBS 0.006204f
C1423 B.n324 VSUBS 0.006204f
C1424 B.n325 VSUBS 0.006204f
C1425 B.n326 VSUBS 0.006204f
C1426 B.n327 VSUBS 0.006204f
C1427 B.n328 VSUBS 0.006204f
C1428 B.n329 VSUBS 0.006204f
C1429 B.n330 VSUBS 0.006204f
C1430 B.n331 VSUBS 0.006204f
C1431 B.n332 VSUBS 0.006204f
C1432 B.n333 VSUBS 0.006204f
C1433 B.n334 VSUBS 0.006204f
C1434 B.n335 VSUBS 0.006204f
C1435 B.n336 VSUBS 0.006204f
C1436 B.n337 VSUBS 0.006204f
C1437 B.n338 VSUBS 0.006204f
C1438 B.n339 VSUBS 0.006204f
C1439 B.n340 VSUBS 0.006204f
C1440 B.n341 VSUBS 0.006204f
C1441 B.n342 VSUBS 0.006204f
C1442 B.n343 VSUBS 0.006204f
C1443 B.n344 VSUBS 0.006204f
C1444 B.n345 VSUBS 0.006204f
C1445 B.n346 VSUBS 0.006204f
C1446 B.n347 VSUBS 0.006204f
C1447 B.n348 VSUBS 0.006204f
C1448 B.n349 VSUBS 0.006204f
C1449 B.n350 VSUBS 0.006204f
C1450 B.n351 VSUBS 0.006204f
C1451 B.n352 VSUBS 0.006204f
C1452 B.n353 VSUBS 0.006204f
C1453 B.n354 VSUBS 0.006204f
C1454 B.n355 VSUBS 0.006204f
C1455 B.n356 VSUBS 0.006204f
C1456 B.n357 VSUBS 0.006204f
C1457 B.n358 VSUBS 0.006204f
C1458 B.n359 VSUBS 0.006204f
C1459 B.n360 VSUBS 0.006204f
C1460 B.n361 VSUBS 0.006204f
C1461 B.n362 VSUBS 0.006204f
C1462 B.n363 VSUBS 0.006204f
C1463 B.n364 VSUBS 0.006204f
C1464 B.n365 VSUBS 0.006204f
C1465 B.n366 VSUBS 0.006204f
C1466 B.n367 VSUBS 0.006204f
C1467 B.n368 VSUBS 0.006204f
C1468 B.n369 VSUBS 0.006204f
C1469 B.n370 VSUBS 0.006204f
C1470 B.n371 VSUBS 0.006204f
C1471 B.n372 VSUBS 0.006204f
C1472 B.n373 VSUBS 0.006204f
C1473 B.n374 VSUBS 0.006204f
C1474 B.n375 VSUBS 0.006204f
C1475 B.n376 VSUBS 0.006204f
C1476 B.n377 VSUBS 0.006204f
C1477 B.n378 VSUBS 0.006204f
C1478 B.n379 VSUBS 0.006204f
C1479 B.n380 VSUBS 0.006204f
C1480 B.n381 VSUBS 0.006204f
C1481 B.n382 VSUBS 0.006204f
C1482 B.n383 VSUBS 0.006204f
C1483 B.n384 VSUBS 0.006204f
C1484 B.n385 VSUBS 0.006204f
C1485 B.n386 VSUBS 0.006204f
C1486 B.n387 VSUBS 0.006204f
C1487 B.n388 VSUBS 0.006204f
C1488 B.n389 VSUBS 0.006204f
C1489 B.n390 VSUBS 0.006204f
C1490 B.n391 VSUBS 0.006204f
C1491 B.n392 VSUBS 0.006204f
C1492 B.n393 VSUBS 0.006204f
C1493 B.n394 VSUBS 0.006204f
C1494 B.n395 VSUBS 0.006204f
C1495 B.n396 VSUBS 0.006204f
C1496 B.n397 VSUBS 0.006204f
C1497 B.n398 VSUBS 0.006204f
C1498 B.n399 VSUBS 0.006204f
C1499 B.n400 VSUBS 0.005839f
C1500 B.n401 VSUBS 0.006204f
C1501 B.n402 VSUBS 0.006204f
C1502 B.n403 VSUBS 0.003467f
C1503 B.n404 VSUBS 0.006204f
C1504 B.n405 VSUBS 0.006204f
C1505 B.n406 VSUBS 0.006204f
C1506 B.n407 VSUBS 0.006204f
C1507 B.n408 VSUBS 0.006204f
C1508 B.n409 VSUBS 0.006204f
C1509 B.n410 VSUBS 0.006204f
C1510 B.n411 VSUBS 0.006204f
C1511 B.n412 VSUBS 0.006204f
C1512 B.n413 VSUBS 0.006204f
C1513 B.n414 VSUBS 0.006204f
C1514 B.n415 VSUBS 0.006204f
C1515 B.n416 VSUBS 0.003467f
C1516 B.n417 VSUBS 0.014373f
C1517 B.n418 VSUBS 0.005839f
C1518 B.n419 VSUBS 0.006204f
C1519 B.n420 VSUBS 0.006204f
C1520 B.n421 VSUBS 0.006204f
C1521 B.n422 VSUBS 0.006204f
C1522 B.n423 VSUBS 0.006204f
C1523 B.n424 VSUBS 0.006204f
C1524 B.n425 VSUBS 0.006204f
C1525 B.n426 VSUBS 0.006204f
C1526 B.n427 VSUBS 0.006204f
C1527 B.n428 VSUBS 0.006204f
C1528 B.n429 VSUBS 0.006204f
C1529 B.n430 VSUBS 0.006204f
C1530 B.n431 VSUBS 0.006204f
C1531 B.n432 VSUBS 0.006204f
C1532 B.n433 VSUBS 0.006204f
C1533 B.n434 VSUBS 0.006204f
C1534 B.n435 VSUBS 0.006204f
C1535 B.n436 VSUBS 0.006204f
C1536 B.n437 VSUBS 0.006204f
C1537 B.n438 VSUBS 0.006204f
C1538 B.n439 VSUBS 0.006204f
C1539 B.n440 VSUBS 0.006204f
C1540 B.n441 VSUBS 0.006204f
C1541 B.n442 VSUBS 0.006204f
C1542 B.n443 VSUBS 0.006204f
C1543 B.n444 VSUBS 0.006204f
C1544 B.n445 VSUBS 0.006204f
C1545 B.n446 VSUBS 0.006204f
C1546 B.n447 VSUBS 0.006204f
C1547 B.n448 VSUBS 0.006204f
C1548 B.n449 VSUBS 0.006204f
C1549 B.n450 VSUBS 0.006204f
C1550 B.n451 VSUBS 0.006204f
C1551 B.n452 VSUBS 0.006204f
C1552 B.n453 VSUBS 0.006204f
C1553 B.n454 VSUBS 0.006204f
C1554 B.n455 VSUBS 0.006204f
C1555 B.n456 VSUBS 0.006204f
C1556 B.n457 VSUBS 0.006204f
C1557 B.n458 VSUBS 0.006204f
C1558 B.n459 VSUBS 0.006204f
C1559 B.n460 VSUBS 0.006204f
C1560 B.n461 VSUBS 0.006204f
C1561 B.n462 VSUBS 0.006204f
C1562 B.n463 VSUBS 0.006204f
C1563 B.n464 VSUBS 0.006204f
C1564 B.n465 VSUBS 0.006204f
C1565 B.n466 VSUBS 0.006204f
C1566 B.n467 VSUBS 0.006204f
C1567 B.n468 VSUBS 0.006204f
C1568 B.n469 VSUBS 0.006204f
C1569 B.n470 VSUBS 0.006204f
C1570 B.n471 VSUBS 0.006204f
C1571 B.n472 VSUBS 0.006204f
C1572 B.n473 VSUBS 0.006204f
C1573 B.n474 VSUBS 0.006204f
C1574 B.n475 VSUBS 0.006204f
C1575 B.n476 VSUBS 0.006204f
C1576 B.n477 VSUBS 0.006204f
C1577 B.n478 VSUBS 0.006204f
C1578 B.n479 VSUBS 0.006204f
C1579 B.n480 VSUBS 0.006204f
C1580 B.n481 VSUBS 0.006204f
C1581 B.n482 VSUBS 0.006204f
C1582 B.n483 VSUBS 0.006204f
C1583 B.n484 VSUBS 0.006204f
C1584 B.n485 VSUBS 0.006204f
C1585 B.n486 VSUBS 0.006204f
C1586 B.n487 VSUBS 0.006204f
C1587 B.n488 VSUBS 0.006204f
C1588 B.n489 VSUBS 0.006204f
C1589 B.n490 VSUBS 0.006204f
C1590 B.n491 VSUBS 0.006204f
C1591 B.n492 VSUBS 0.006204f
C1592 B.n493 VSUBS 0.006204f
C1593 B.n494 VSUBS 0.006204f
C1594 B.n495 VSUBS 0.006204f
C1595 B.n496 VSUBS 0.006204f
C1596 B.n497 VSUBS 0.006204f
C1597 B.n498 VSUBS 0.006204f
C1598 B.n499 VSUBS 0.006204f
C1599 B.n500 VSUBS 0.006204f
C1600 B.n501 VSUBS 0.006204f
C1601 B.n502 VSUBS 0.006204f
C1602 B.n503 VSUBS 0.006204f
C1603 B.n504 VSUBS 0.006204f
C1604 B.n505 VSUBS 0.006204f
C1605 B.n506 VSUBS 0.006204f
C1606 B.n507 VSUBS 0.006204f
C1607 B.n508 VSUBS 0.006204f
C1608 B.n509 VSUBS 0.006204f
C1609 B.n510 VSUBS 0.006204f
C1610 B.n511 VSUBS 0.006204f
C1611 B.n512 VSUBS 0.006204f
C1612 B.n513 VSUBS 0.014984f
C1613 B.n514 VSUBS 0.013845f
C1614 B.n515 VSUBS 0.013845f
C1615 B.n516 VSUBS 0.006204f
C1616 B.n517 VSUBS 0.006204f
C1617 B.n518 VSUBS 0.006204f
C1618 B.n519 VSUBS 0.006204f
C1619 B.n520 VSUBS 0.006204f
C1620 B.n521 VSUBS 0.006204f
C1621 B.n522 VSUBS 0.006204f
C1622 B.n523 VSUBS 0.006204f
C1623 B.n524 VSUBS 0.006204f
C1624 B.n525 VSUBS 0.006204f
C1625 B.n526 VSUBS 0.006204f
C1626 B.n527 VSUBS 0.006204f
C1627 B.n528 VSUBS 0.006204f
C1628 B.n529 VSUBS 0.006204f
C1629 B.n530 VSUBS 0.006204f
C1630 B.n531 VSUBS 0.006204f
C1631 B.n532 VSUBS 0.006204f
C1632 B.n533 VSUBS 0.006204f
C1633 B.n534 VSUBS 0.006204f
C1634 B.n535 VSUBS 0.006204f
C1635 B.n536 VSUBS 0.006204f
C1636 B.n537 VSUBS 0.006204f
C1637 B.n538 VSUBS 0.006204f
C1638 B.n539 VSUBS 0.006204f
C1639 B.n540 VSUBS 0.006204f
C1640 B.n541 VSUBS 0.006204f
C1641 B.n542 VSUBS 0.006204f
C1642 B.n543 VSUBS 0.006204f
C1643 B.n544 VSUBS 0.006204f
C1644 B.n545 VSUBS 0.006204f
C1645 B.n546 VSUBS 0.006204f
C1646 B.n547 VSUBS 0.006204f
C1647 B.n548 VSUBS 0.006204f
C1648 B.n549 VSUBS 0.006204f
C1649 B.n550 VSUBS 0.006204f
C1650 B.n551 VSUBS 0.006204f
C1651 B.n552 VSUBS 0.006204f
C1652 B.n553 VSUBS 0.006204f
C1653 B.n554 VSUBS 0.006204f
C1654 B.n555 VSUBS 0.006204f
C1655 B.n556 VSUBS 0.006204f
C1656 B.n557 VSUBS 0.006204f
C1657 B.n558 VSUBS 0.006204f
C1658 B.n559 VSUBS 0.006204f
C1659 B.n560 VSUBS 0.006204f
C1660 B.n561 VSUBS 0.006204f
C1661 B.n562 VSUBS 0.006204f
C1662 B.n563 VSUBS 0.006204f
C1663 B.n564 VSUBS 0.006204f
C1664 B.n565 VSUBS 0.006204f
C1665 B.n566 VSUBS 0.006204f
C1666 B.n567 VSUBS 0.006204f
C1667 B.n568 VSUBS 0.006204f
C1668 B.n569 VSUBS 0.006204f
C1669 B.n570 VSUBS 0.006204f
C1670 B.n571 VSUBS 0.006204f
C1671 B.n572 VSUBS 0.006204f
C1672 B.n573 VSUBS 0.006204f
C1673 B.n574 VSUBS 0.006204f
C1674 B.n575 VSUBS 0.006204f
C1675 B.n576 VSUBS 0.006204f
C1676 B.n577 VSUBS 0.006204f
C1677 B.n578 VSUBS 0.006204f
C1678 B.n579 VSUBS 0.006204f
C1679 B.n580 VSUBS 0.006204f
C1680 B.n581 VSUBS 0.006204f
C1681 B.n582 VSUBS 0.006204f
C1682 B.n583 VSUBS 0.006204f
C1683 B.n584 VSUBS 0.006204f
C1684 B.n585 VSUBS 0.006204f
C1685 B.n586 VSUBS 0.006204f
C1686 B.n587 VSUBS 0.006204f
C1687 B.n588 VSUBS 0.006204f
C1688 B.n589 VSUBS 0.006204f
C1689 B.n590 VSUBS 0.006204f
C1690 B.n591 VSUBS 0.006204f
C1691 B.n592 VSUBS 0.006204f
C1692 B.n593 VSUBS 0.006204f
C1693 B.n594 VSUBS 0.006204f
C1694 B.n595 VSUBS 0.006204f
C1695 B.n596 VSUBS 0.006204f
C1696 B.n597 VSUBS 0.006204f
C1697 B.n598 VSUBS 0.006204f
C1698 B.n599 VSUBS 0.006204f
C1699 B.n600 VSUBS 0.006204f
C1700 B.n601 VSUBS 0.006204f
C1701 B.n602 VSUBS 0.006204f
C1702 B.n603 VSUBS 0.006204f
C1703 B.n604 VSUBS 0.006204f
C1704 B.n605 VSUBS 0.006204f
C1705 B.n606 VSUBS 0.006204f
C1706 B.n607 VSUBS 0.006204f
C1707 B.n608 VSUBS 0.006204f
C1708 B.n609 VSUBS 0.006204f
C1709 B.n610 VSUBS 0.006204f
C1710 B.n611 VSUBS 0.006204f
C1711 B.n612 VSUBS 0.006204f
C1712 B.n613 VSUBS 0.006204f
C1713 B.n614 VSUBS 0.006204f
C1714 B.n615 VSUBS 0.006204f
C1715 B.n616 VSUBS 0.006204f
C1716 B.n617 VSUBS 0.006204f
C1717 B.n618 VSUBS 0.006204f
C1718 B.n619 VSUBS 0.006204f
C1719 B.n620 VSUBS 0.006204f
C1720 B.n621 VSUBS 0.006204f
C1721 B.n622 VSUBS 0.006204f
C1722 B.n623 VSUBS 0.006204f
C1723 B.n624 VSUBS 0.006204f
C1724 B.n625 VSUBS 0.006204f
C1725 B.n626 VSUBS 0.006204f
C1726 B.n627 VSUBS 0.006204f
C1727 B.n628 VSUBS 0.006204f
C1728 B.n629 VSUBS 0.006204f
C1729 B.n630 VSUBS 0.006204f
C1730 B.n631 VSUBS 0.006204f
C1731 B.n632 VSUBS 0.006204f
C1732 B.n633 VSUBS 0.006204f
C1733 B.n634 VSUBS 0.006204f
C1734 B.n635 VSUBS 0.006204f
C1735 B.n636 VSUBS 0.006204f
C1736 B.n637 VSUBS 0.006204f
C1737 B.n638 VSUBS 0.006204f
C1738 B.n639 VSUBS 0.006204f
C1739 B.n640 VSUBS 0.006204f
C1740 B.n641 VSUBS 0.006204f
C1741 B.n642 VSUBS 0.006204f
C1742 B.n643 VSUBS 0.006204f
C1743 B.n644 VSUBS 0.006204f
C1744 B.n645 VSUBS 0.006204f
C1745 B.n646 VSUBS 0.006204f
C1746 B.n647 VSUBS 0.006204f
C1747 B.n648 VSUBS 0.006204f
C1748 B.n649 VSUBS 0.013845f
C1749 B.n650 VSUBS 0.014586f
C1750 B.n651 VSUBS 0.014243f
C1751 B.n652 VSUBS 0.006204f
C1752 B.n653 VSUBS 0.006204f
C1753 B.n654 VSUBS 0.006204f
C1754 B.n655 VSUBS 0.006204f
C1755 B.n656 VSUBS 0.006204f
C1756 B.n657 VSUBS 0.006204f
C1757 B.n658 VSUBS 0.006204f
C1758 B.n659 VSUBS 0.006204f
C1759 B.n660 VSUBS 0.006204f
C1760 B.n661 VSUBS 0.006204f
C1761 B.n662 VSUBS 0.006204f
C1762 B.n663 VSUBS 0.006204f
C1763 B.n664 VSUBS 0.006204f
C1764 B.n665 VSUBS 0.006204f
C1765 B.n666 VSUBS 0.006204f
C1766 B.n667 VSUBS 0.006204f
C1767 B.n668 VSUBS 0.006204f
C1768 B.n669 VSUBS 0.006204f
C1769 B.n670 VSUBS 0.006204f
C1770 B.n671 VSUBS 0.006204f
C1771 B.n672 VSUBS 0.006204f
C1772 B.n673 VSUBS 0.006204f
C1773 B.n674 VSUBS 0.006204f
C1774 B.n675 VSUBS 0.006204f
C1775 B.n676 VSUBS 0.006204f
C1776 B.n677 VSUBS 0.006204f
C1777 B.n678 VSUBS 0.006204f
C1778 B.n679 VSUBS 0.006204f
C1779 B.n680 VSUBS 0.006204f
C1780 B.n681 VSUBS 0.006204f
C1781 B.n682 VSUBS 0.006204f
C1782 B.n683 VSUBS 0.006204f
C1783 B.n684 VSUBS 0.006204f
C1784 B.n685 VSUBS 0.006204f
C1785 B.n686 VSUBS 0.006204f
C1786 B.n687 VSUBS 0.006204f
C1787 B.n688 VSUBS 0.006204f
C1788 B.n689 VSUBS 0.006204f
C1789 B.n690 VSUBS 0.006204f
C1790 B.n691 VSUBS 0.006204f
C1791 B.n692 VSUBS 0.006204f
C1792 B.n693 VSUBS 0.006204f
C1793 B.n694 VSUBS 0.006204f
C1794 B.n695 VSUBS 0.006204f
C1795 B.n696 VSUBS 0.006204f
C1796 B.n697 VSUBS 0.006204f
C1797 B.n698 VSUBS 0.006204f
C1798 B.n699 VSUBS 0.006204f
C1799 B.n700 VSUBS 0.006204f
C1800 B.n701 VSUBS 0.006204f
C1801 B.n702 VSUBS 0.006204f
C1802 B.n703 VSUBS 0.006204f
C1803 B.n704 VSUBS 0.006204f
C1804 B.n705 VSUBS 0.006204f
C1805 B.n706 VSUBS 0.006204f
C1806 B.n707 VSUBS 0.006204f
C1807 B.n708 VSUBS 0.006204f
C1808 B.n709 VSUBS 0.006204f
C1809 B.n710 VSUBS 0.006204f
C1810 B.n711 VSUBS 0.006204f
C1811 B.n712 VSUBS 0.006204f
C1812 B.n713 VSUBS 0.006204f
C1813 B.n714 VSUBS 0.006204f
C1814 B.n715 VSUBS 0.006204f
C1815 B.n716 VSUBS 0.006204f
C1816 B.n717 VSUBS 0.006204f
C1817 B.n718 VSUBS 0.006204f
C1818 B.n719 VSUBS 0.006204f
C1819 B.n720 VSUBS 0.006204f
C1820 B.n721 VSUBS 0.006204f
C1821 B.n722 VSUBS 0.006204f
C1822 B.n723 VSUBS 0.006204f
C1823 B.n724 VSUBS 0.006204f
C1824 B.n725 VSUBS 0.006204f
C1825 B.n726 VSUBS 0.006204f
C1826 B.n727 VSUBS 0.006204f
C1827 B.n728 VSUBS 0.006204f
C1828 B.n729 VSUBS 0.006204f
C1829 B.n730 VSUBS 0.006204f
C1830 B.n731 VSUBS 0.006204f
C1831 B.n732 VSUBS 0.006204f
C1832 B.n733 VSUBS 0.006204f
C1833 B.n734 VSUBS 0.006204f
C1834 B.n735 VSUBS 0.006204f
C1835 B.n736 VSUBS 0.006204f
C1836 B.n737 VSUBS 0.006204f
C1837 B.n738 VSUBS 0.006204f
C1838 B.n739 VSUBS 0.006204f
C1839 B.n740 VSUBS 0.006204f
C1840 B.n741 VSUBS 0.006204f
C1841 B.n742 VSUBS 0.006204f
C1842 B.n743 VSUBS 0.006204f
C1843 B.n744 VSUBS 0.006204f
C1844 B.n745 VSUBS 0.006204f
C1845 B.n746 VSUBS 0.005839f
C1846 B.n747 VSUBS 0.014373f
C1847 B.n748 VSUBS 0.003467f
C1848 B.n749 VSUBS 0.006204f
C1849 B.n750 VSUBS 0.006204f
C1850 B.n751 VSUBS 0.006204f
C1851 B.n752 VSUBS 0.006204f
C1852 B.n753 VSUBS 0.006204f
C1853 B.n754 VSUBS 0.006204f
C1854 B.n755 VSUBS 0.006204f
C1855 B.n756 VSUBS 0.006204f
C1856 B.n757 VSUBS 0.006204f
C1857 B.n758 VSUBS 0.006204f
C1858 B.n759 VSUBS 0.006204f
C1859 B.n760 VSUBS 0.006204f
C1860 B.n761 VSUBS 0.003467f
C1861 B.n762 VSUBS 0.006204f
C1862 B.n763 VSUBS 0.006204f
C1863 B.n764 VSUBS 0.006204f
C1864 B.n765 VSUBS 0.006204f
C1865 B.n766 VSUBS 0.006204f
C1866 B.n767 VSUBS 0.006204f
C1867 B.n768 VSUBS 0.006204f
C1868 B.n769 VSUBS 0.006204f
C1869 B.n770 VSUBS 0.006204f
C1870 B.n771 VSUBS 0.006204f
C1871 B.n772 VSUBS 0.006204f
C1872 B.n773 VSUBS 0.006204f
C1873 B.n774 VSUBS 0.006204f
C1874 B.n775 VSUBS 0.006204f
C1875 B.n776 VSUBS 0.006204f
C1876 B.n777 VSUBS 0.006204f
C1877 B.n778 VSUBS 0.006204f
C1878 B.n779 VSUBS 0.006204f
C1879 B.n780 VSUBS 0.006204f
C1880 B.n781 VSUBS 0.006204f
C1881 B.n782 VSUBS 0.006204f
C1882 B.n783 VSUBS 0.006204f
C1883 B.n784 VSUBS 0.006204f
C1884 B.n785 VSUBS 0.006204f
C1885 B.n786 VSUBS 0.006204f
C1886 B.n787 VSUBS 0.006204f
C1887 B.n788 VSUBS 0.006204f
C1888 B.n789 VSUBS 0.006204f
C1889 B.n790 VSUBS 0.006204f
C1890 B.n791 VSUBS 0.006204f
C1891 B.n792 VSUBS 0.006204f
C1892 B.n793 VSUBS 0.006204f
C1893 B.n794 VSUBS 0.006204f
C1894 B.n795 VSUBS 0.006204f
C1895 B.n796 VSUBS 0.006204f
C1896 B.n797 VSUBS 0.006204f
C1897 B.n798 VSUBS 0.006204f
C1898 B.n799 VSUBS 0.006204f
C1899 B.n800 VSUBS 0.006204f
C1900 B.n801 VSUBS 0.006204f
C1901 B.n802 VSUBS 0.006204f
C1902 B.n803 VSUBS 0.006204f
C1903 B.n804 VSUBS 0.006204f
C1904 B.n805 VSUBS 0.006204f
C1905 B.n806 VSUBS 0.006204f
C1906 B.n807 VSUBS 0.006204f
C1907 B.n808 VSUBS 0.006204f
C1908 B.n809 VSUBS 0.006204f
C1909 B.n810 VSUBS 0.006204f
C1910 B.n811 VSUBS 0.006204f
C1911 B.n812 VSUBS 0.006204f
C1912 B.n813 VSUBS 0.006204f
C1913 B.n814 VSUBS 0.006204f
C1914 B.n815 VSUBS 0.006204f
C1915 B.n816 VSUBS 0.006204f
C1916 B.n817 VSUBS 0.006204f
C1917 B.n818 VSUBS 0.006204f
C1918 B.n819 VSUBS 0.006204f
C1919 B.n820 VSUBS 0.006204f
C1920 B.n821 VSUBS 0.006204f
C1921 B.n822 VSUBS 0.006204f
C1922 B.n823 VSUBS 0.006204f
C1923 B.n824 VSUBS 0.006204f
C1924 B.n825 VSUBS 0.006204f
C1925 B.n826 VSUBS 0.006204f
C1926 B.n827 VSUBS 0.006204f
C1927 B.n828 VSUBS 0.006204f
C1928 B.n829 VSUBS 0.006204f
C1929 B.n830 VSUBS 0.006204f
C1930 B.n831 VSUBS 0.006204f
C1931 B.n832 VSUBS 0.006204f
C1932 B.n833 VSUBS 0.006204f
C1933 B.n834 VSUBS 0.006204f
C1934 B.n835 VSUBS 0.006204f
C1935 B.n836 VSUBS 0.006204f
C1936 B.n837 VSUBS 0.006204f
C1937 B.n838 VSUBS 0.006204f
C1938 B.n839 VSUBS 0.006204f
C1939 B.n840 VSUBS 0.006204f
C1940 B.n841 VSUBS 0.006204f
C1941 B.n842 VSUBS 0.006204f
C1942 B.n843 VSUBS 0.006204f
C1943 B.n844 VSUBS 0.006204f
C1944 B.n845 VSUBS 0.006204f
C1945 B.n846 VSUBS 0.006204f
C1946 B.n847 VSUBS 0.006204f
C1947 B.n848 VSUBS 0.006204f
C1948 B.n849 VSUBS 0.006204f
C1949 B.n850 VSUBS 0.006204f
C1950 B.n851 VSUBS 0.006204f
C1951 B.n852 VSUBS 0.006204f
C1952 B.n853 VSUBS 0.006204f
C1953 B.n854 VSUBS 0.006204f
C1954 B.n855 VSUBS 0.006204f
C1955 B.n856 VSUBS 0.006204f
C1956 B.n857 VSUBS 0.014984f
C1957 B.n858 VSUBS 0.014984f
C1958 B.n859 VSUBS 0.013845f
C1959 B.n860 VSUBS 0.006204f
C1960 B.n861 VSUBS 0.006204f
C1961 B.n862 VSUBS 0.006204f
C1962 B.n863 VSUBS 0.006204f
C1963 B.n864 VSUBS 0.006204f
C1964 B.n865 VSUBS 0.006204f
C1965 B.n866 VSUBS 0.006204f
C1966 B.n867 VSUBS 0.006204f
C1967 B.n868 VSUBS 0.006204f
C1968 B.n869 VSUBS 0.006204f
C1969 B.n870 VSUBS 0.006204f
C1970 B.n871 VSUBS 0.006204f
C1971 B.n872 VSUBS 0.006204f
C1972 B.n873 VSUBS 0.006204f
C1973 B.n874 VSUBS 0.006204f
C1974 B.n875 VSUBS 0.006204f
C1975 B.n876 VSUBS 0.006204f
C1976 B.n877 VSUBS 0.006204f
C1977 B.n878 VSUBS 0.006204f
C1978 B.n879 VSUBS 0.006204f
C1979 B.n880 VSUBS 0.006204f
C1980 B.n881 VSUBS 0.006204f
C1981 B.n882 VSUBS 0.006204f
C1982 B.n883 VSUBS 0.006204f
C1983 B.n884 VSUBS 0.006204f
C1984 B.n885 VSUBS 0.006204f
C1985 B.n886 VSUBS 0.006204f
C1986 B.n887 VSUBS 0.006204f
C1987 B.n888 VSUBS 0.006204f
C1988 B.n889 VSUBS 0.006204f
C1989 B.n890 VSUBS 0.006204f
C1990 B.n891 VSUBS 0.006204f
C1991 B.n892 VSUBS 0.006204f
C1992 B.n893 VSUBS 0.006204f
C1993 B.n894 VSUBS 0.006204f
C1994 B.n895 VSUBS 0.006204f
C1995 B.n896 VSUBS 0.006204f
C1996 B.n897 VSUBS 0.006204f
C1997 B.n898 VSUBS 0.006204f
C1998 B.n899 VSUBS 0.006204f
C1999 B.n900 VSUBS 0.006204f
C2000 B.n901 VSUBS 0.006204f
C2001 B.n902 VSUBS 0.006204f
C2002 B.n903 VSUBS 0.006204f
C2003 B.n904 VSUBS 0.006204f
C2004 B.n905 VSUBS 0.006204f
C2005 B.n906 VSUBS 0.006204f
C2006 B.n907 VSUBS 0.006204f
C2007 B.n908 VSUBS 0.006204f
C2008 B.n909 VSUBS 0.006204f
C2009 B.n910 VSUBS 0.006204f
C2010 B.n911 VSUBS 0.006204f
C2011 B.n912 VSUBS 0.006204f
C2012 B.n913 VSUBS 0.006204f
C2013 B.n914 VSUBS 0.006204f
C2014 B.n915 VSUBS 0.006204f
C2015 B.n916 VSUBS 0.006204f
C2016 B.n917 VSUBS 0.006204f
C2017 B.n918 VSUBS 0.006204f
C2018 B.n919 VSUBS 0.006204f
C2019 B.n920 VSUBS 0.006204f
C2020 B.n921 VSUBS 0.006204f
C2021 B.n922 VSUBS 0.006204f
C2022 B.n923 VSUBS 0.006204f
C2023 B.n924 VSUBS 0.006204f
C2024 B.n925 VSUBS 0.006204f
C2025 B.n926 VSUBS 0.006204f
C2026 B.n927 VSUBS 0.014048f
.ends

