* NGSPICE file created from diff_pair_sample_0701.ext - technology: sky130A

.subckt diff_pair_sample_0701 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=0 ps=0 w=3.77 l=1.93
X1 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=0 ps=0 w=3.77 l=1.93
X2 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=0 ps=0 w=3.77 l=1.93
X3 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=0 ps=0 w=3.77 l=1.93
X4 VDD2.t1 VN.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=1.4703 ps=8.32 w=3.77 l=1.93
X5 VDD2.t0 VN.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=1.4703 ps=8.32 w=3.77 l=1.93
X6 VDD1.t1 VP.t0 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=1.4703 ps=8.32 w=3.77 l=1.93
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.4703 pd=8.32 as=1.4703 ps=8.32 w=3.77 l=1.93
R0 B.n404 B.n403 585
R1 B.n155 B.n64 585
R2 B.n154 B.n153 585
R3 B.n152 B.n151 585
R4 B.n150 B.n149 585
R5 B.n148 B.n147 585
R6 B.n146 B.n145 585
R7 B.n144 B.n143 585
R8 B.n142 B.n141 585
R9 B.n140 B.n139 585
R10 B.n138 B.n137 585
R11 B.n136 B.n135 585
R12 B.n134 B.n133 585
R13 B.n132 B.n131 585
R14 B.n130 B.n129 585
R15 B.n128 B.n127 585
R16 B.n126 B.n125 585
R17 B.n123 B.n122 585
R18 B.n121 B.n120 585
R19 B.n119 B.n118 585
R20 B.n117 B.n116 585
R21 B.n115 B.n114 585
R22 B.n113 B.n112 585
R23 B.n111 B.n110 585
R24 B.n109 B.n108 585
R25 B.n107 B.n106 585
R26 B.n105 B.n104 585
R27 B.n102 B.n101 585
R28 B.n100 B.n99 585
R29 B.n98 B.n97 585
R30 B.n96 B.n95 585
R31 B.n94 B.n93 585
R32 B.n92 B.n91 585
R33 B.n90 B.n89 585
R34 B.n88 B.n87 585
R35 B.n86 B.n85 585
R36 B.n84 B.n83 585
R37 B.n82 B.n81 585
R38 B.n80 B.n79 585
R39 B.n78 B.n77 585
R40 B.n76 B.n75 585
R41 B.n74 B.n73 585
R42 B.n72 B.n71 585
R43 B.n70 B.n69 585
R44 B.n402 B.n42 585
R45 B.n407 B.n42 585
R46 B.n401 B.n41 585
R47 B.n408 B.n41 585
R48 B.n400 B.n399 585
R49 B.n399 B.n37 585
R50 B.n398 B.n36 585
R51 B.n414 B.n36 585
R52 B.n397 B.n35 585
R53 B.n415 B.n35 585
R54 B.n396 B.n34 585
R55 B.n416 B.n34 585
R56 B.n395 B.n394 585
R57 B.n394 B.n33 585
R58 B.n393 B.n29 585
R59 B.n422 B.n29 585
R60 B.n392 B.n28 585
R61 B.n423 B.n28 585
R62 B.n391 B.n27 585
R63 B.n424 B.n27 585
R64 B.n390 B.n389 585
R65 B.n389 B.n23 585
R66 B.n388 B.n22 585
R67 B.n430 B.n22 585
R68 B.n387 B.n21 585
R69 B.n431 B.n21 585
R70 B.n386 B.n20 585
R71 B.n432 B.n20 585
R72 B.n385 B.n384 585
R73 B.n384 B.n16 585
R74 B.n383 B.n15 585
R75 B.n438 B.n15 585
R76 B.n382 B.n14 585
R77 B.n439 B.n14 585
R78 B.n381 B.n13 585
R79 B.n440 B.n13 585
R80 B.n380 B.n379 585
R81 B.n379 B.n12 585
R82 B.n378 B.n377 585
R83 B.n378 B.n8 585
R84 B.n376 B.n7 585
R85 B.n447 B.n7 585
R86 B.n375 B.n6 585
R87 B.n448 B.n6 585
R88 B.n374 B.n5 585
R89 B.n449 B.n5 585
R90 B.n373 B.n372 585
R91 B.n372 B.n4 585
R92 B.n371 B.n156 585
R93 B.n371 B.n370 585
R94 B.n361 B.n157 585
R95 B.n158 B.n157 585
R96 B.n363 B.n362 585
R97 B.n364 B.n363 585
R98 B.n360 B.n162 585
R99 B.n166 B.n162 585
R100 B.n359 B.n358 585
R101 B.n358 B.n357 585
R102 B.n164 B.n163 585
R103 B.n165 B.n164 585
R104 B.n350 B.n349 585
R105 B.n351 B.n350 585
R106 B.n348 B.n171 585
R107 B.n171 B.n170 585
R108 B.n347 B.n346 585
R109 B.n346 B.n345 585
R110 B.n173 B.n172 585
R111 B.n174 B.n173 585
R112 B.n338 B.n337 585
R113 B.n339 B.n338 585
R114 B.n336 B.n179 585
R115 B.n179 B.n178 585
R116 B.n335 B.n334 585
R117 B.n334 B.n333 585
R118 B.n181 B.n180 585
R119 B.n326 B.n181 585
R120 B.n325 B.n324 585
R121 B.n327 B.n325 585
R122 B.n323 B.n186 585
R123 B.n186 B.n185 585
R124 B.n322 B.n321 585
R125 B.n321 B.n320 585
R126 B.n188 B.n187 585
R127 B.n189 B.n188 585
R128 B.n313 B.n312 585
R129 B.n314 B.n313 585
R130 B.n311 B.n194 585
R131 B.n194 B.n193 585
R132 B.n306 B.n305 585
R133 B.n304 B.n218 585
R134 B.n303 B.n217 585
R135 B.n308 B.n217 585
R136 B.n302 B.n301 585
R137 B.n300 B.n299 585
R138 B.n298 B.n297 585
R139 B.n296 B.n295 585
R140 B.n294 B.n293 585
R141 B.n292 B.n291 585
R142 B.n290 B.n289 585
R143 B.n288 B.n287 585
R144 B.n286 B.n285 585
R145 B.n284 B.n283 585
R146 B.n282 B.n281 585
R147 B.n280 B.n279 585
R148 B.n278 B.n277 585
R149 B.n276 B.n275 585
R150 B.n274 B.n273 585
R151 B.n272 B.n271 585
R152 B.n270 B.n269 585
R153 B.n268 B.n267 585
R154 B.n266 B.n265 585
R155 B.n264 B.n263 585
R156 B.n262 B.n261 585
R157 B.n260 B.n259 585
R158 B.n258 B.n257 585
R159 B.n256 B.n255 585
R160 B.n254 B.n253 585
R161 B.n252 B.n251 585
R162 B.n250 B.n249 585
R163 B.n248 B.n247 585
R164 B.n246 B.n245 585
R165 B.n244 B.n243 585
R166 B.n242 B.n241 585
R167 B.n240 B.n239 585
R168 B.n238 B.n237 585
R169 B.n236 B.n235 585
R170 B.n234 B.n233 585
R171 B.n232 B.n231 585
R172 B.n230 B.n229 585
R173 B.n228 B.n227 585
R174 B.n226 B.n225 585
R175 B.n196 B.n195 585
R176 B.n310 B.n309 585
R177 B.n309 B.n308 585
R178 B.n192 B.n191 585
R179 B.n193 B.n192 585
R180 B.n316 B.n315 585
R181 B.n315 B.n314 585
R182 B.n317 B.n190 585
R183 B.n190 B.n189 585
R184 B.n319 B.n318 585
R185 B.n320 B.n319 585
R186 B.n184 B.n183 585
R187 B.n185 B.n184 585
R188 B.n329 B.n328 585
R189 B.n328 B.n327 585
R190 B.n330 B.n182 585
R191 B.n326 B.n182 585
R192 B.n332 B.n331 585
R193 B.n333 B.n332 585
R194 B.n177 B.n176 585
R195 B.n178 B.n177 585
R196 B.n341 B.n340 585
R197 B.n340 B.n339 585
R198 B.n342 B.n175 585
R199 B.n175 B.n174 585
R200 B.n344 B.n343 585
R201 B.n345 B.n344 585
R202 B.n169 B.n168 585
R203 B.n170 B.n169 585
R204 B.n353 B.n352 585
R205 B.n352 B.n351 585
R206 B.n354 B.n167 585
R207 B.n167 B.n165 585
R208 B.n356 B.n355 585
R209 B.n357 B.n356 585
R210 B.n161 B.n160 585
R211 B.n166 B.n161 585
R212 B.n366 B.n365 585
R213 B.n365 B.n364 585
R214 B.n367 B.n159 585
R215 B.n159 B.n158 585
R216 B.n369 B.n368 585
R217 B.n370 B.n369 585
R218 B.n3 B.n0 585
R219 B.n4 B.n3 585
R220 B.n446 B.n1 585
R221 B.n447 B.n446 585
R222 B.n445 B.n444 585
R223 B.n445 B.n8 585
R224 B.n443 B.n9 585
R225 B.n12 B.n9 585
R226 B.n442 B.n441 585
R227 B.n441 B.n440 585
R228 B.n11 B.n10 585
R229 B.n439 B.n11 585
R230 B.n437 B.n436 585
R231 B.n438 B.n437 585
R232 B.n435 B.n17 585
R233 B.n17 B.n16 585
R234 B.n434 B.n433 585
R235 B.n433 B.n432 585
R236 B.n19 B.n18 585
R237 B.n431 B.n19 585
R238 B.n429 B.n428 585
R239 B.n430 B.n429 585
R240 B.n427 B.n24 585
R241 B.n24 B.n23 585
R242 B.n426 B.n425 585
R243 B.n425 B.n424 585
R244 B.n26 B.n25 585
R245 B.n423 B.n26 585
R246 B.n421 B.n420 585
R247 B.n422 B.n421 585
R248 B.n419 B.n30 585
R249 B.n33 B.n30 585
R250 B.n418 B.n417 585
R251 B.n417 B.n416 585
R252 B.n32 B.n31 585
R253 B.n415 B.n32 585
R254 B.n413 B.n412 585
R255 B.n414 B.n413 585
R256 B.n411 B.n38 585
R257 B.n38 B.n37 585
R258 B.n410 B.n409 585
R259 B.n409 B.n408 585
R260 B.n40 B.n39 585
R261 B.n407 B.n40 585
R262 B.n450 B.n449 585
R263 B.n448 B.n2 585
R264 B.n69 B.n40 516.524
R265 B.n404 B.n42 516.524
R266 B.n309 B.n194 516.524
R267 B.n306 B.n192 516.524
R268 B.n406 B.n405 256.663
R269 B.n406 B.n63 256.663
R270 B.n406 B.n62 256.663
R271 B.n406 B.n61 256.663
R272 B.n406 B.n60 256.663
R273 B.n406 B.n59 256.663
R274 B.n406 B.n58 256.663
R275 B.n406 B.n57 256.663
R276 B.n406 B.n56 256.663
R277 B.n406 B.n55 256.663
R278 B.n406 B.n54 256.663
R279 B.n406 B.n53 256.663
R280 B.n406 B.n52 256.663
R281 B.n406 B.n51 256.663
R282 B.n406 B.n50 256.663
R283 B.n406 B.n49 256.663
R284 B.n406 B.n48 256.663
R285 B.n406 B.n47 256.663
R286 B.n406 B.n46 256.663
R287 B.n406 B.n45 256.663
R288 B.n406 B.n44 256.663
R289 B.n406 B.n43 256.663
R290 B.n308 B.n307 256.663
R291 B.n308 B.n197 256.663
R292 B.n308 B.n198 256.663
R293 B.n308 B.n199 256.663
R294 B.n308 B.n200 256.663
R295 B.n308 B.n201 256.663
R296 B.n308 B.n202 256.663
R297 B.n308 B.n203 256.663
R298 B.n308 B.n204 256.663
R299 B.n308 B.n205 256.663
R300 B.n308 B.n206 256.663
R301 B.n308 B.n207 256.663
R302 B.n308 B.n208 256.663
R303 B.n308 B.n209 256.663
R304 B.n308 B.n210 256.663
R305 B.n308 B.n211 256.663
R306 B.n308 B.n212 256.663
R307 B.n308 B.n213 256.663
R308 B.n308 B.n214 256.663
R309 B.n308 B.n215 256.663
R310 B.n308 B.n216 256.663
R311 B.n452 B.n451 256.663
R312 B.n67 B.t10 253.825
R313 B.n65 B.t2 253.825
R314 B.n222 B.t13 253.825
R315 B.n219 B.t6 253.825
R316 B.n65 B.t4 184.63
R317 B.n222 B.t15 184.63
R318 B.n67 B.t11 184.63
R319 B.n219 B.t9 184.63
R320 B.n73 B.n72 163.367
R321 B.n77 B.n76 163.367
R322 B.n81 B.n80 163.367
R323 B.n85 B.n84 163.367
R324 B.n89 B.n88 163.367
R325 B.n93 B.n92 163.367
R326 B.n97 B.n96 163.367
R327 B.n101 B.n100 163.367
R328 B.n106 B.n105 163.367
R329 B.n110 B.n109 163.367
R330 B.n114 B.n113 163.367
R331 B.n118 B.n117 163.367
R332 B.n122 B.n121 163.367
R333 B.n127 B.n126 163.367
R334 B.n131 B.n130 163.367
R335 B.n135 B.n134 163.367
R336 B.n139 B.n138 163.367
R337 B.n143 B.n142 163.367
R338 B.n147 B.n146 163.367
R339 B.n151 B.n150 163.367
R340 B.n153 B.n64 163.367
R341 B.n313 B.n194 163.367
R342 B.n313 B.n188 163.367
R343 B.n321 B.n188 163.367
R344 B.n321 B.n186 163.367
R345 B.n325 B.n186 163.367
R346 B.n325 B.n181 163.367
R347 B.n334 B.n181 163.367
R348 B.n334 B.n179 163.367
R349 B.n338 B.n179 163.367
R350 B.n338 B.n173 163.367
R351 B.n346 B.n173 163.367
R352 B.n346 B.n171 163.367
R353 B.n350 B.n171 163.367
R354 B.n350 B.n164 163.367
R355 B.n358 B.n164 163.367
R356 B.n358 B.n162 163.367
R357 B.n363 B.n162 163.367
R358 B.n363 B.n157 163.367
R359 B.n371 B.n157 163.367
R360 B.n372 B.n371 163.367
R361 B.n372 B.n5 163.367
R362 B.n6 B.n5 163.367
R363 B.n7 B.n6 163.367
R364 B.n378 B.n7 163.367
R365 B.n379 B.n378 163.367
R366 B.n379 B.n13 163.367
R367 B.n14 B.n13 163.367
R368 B.n15 B.n14 163.367
R369 B.n384 B.n15 163.367
R370 B.n384 B.n20 163.367
R371 B.n21 B.n20 163.367
R372 B.n22 B.n21 163.367
R373 B.n389 B.n22 163.367
R374 B.n389 B.n27 163.367
R375 B.n28 B.n27 163.367
R376 B.n29 B.n28 163.367
R377 B.n394 B.n29 163.367
R378 B.n394 B.n34 163.367
R379 B.n35 B.n34 163.367
R380 B.n36 B.n35 163.367
R381 B.n399 B.n36 163.367
R382 B.n399 B.n41 163.367
R383 B.n42 B.n41 163.367
R384 B.n218 B.n217 163.367
R385 B.n301 B.n217 163.367
R386 B.n299 B.n298 163.367
R387 B.n295 B.n294 163.367
R388 B.n291 B.n290 163.367
R389 B.n287 B.n286 163.367
R390 B.n283 B.n282 163.367
R391 B.n279 B.n278 163.367
R392 B.n275 B.n274 163.367
R393 B.n271 B.n270 163.367
R394 B.n267 B.n266 163.367
R395 B.n263 B.n262 163.367
R396 B.n259 B.n258 163.367
R397 B.n255 B.n254 163.367
R398 B.n251 B.n250 163.367
R399 B.n247 B.n246 163.367
R400 B.n243 B.n242 163.367
R401 B.n239 B.n238 163.367
R402 B.n235 B.n234 163.367
R403 B.n231 B.n230 163.367
R404 B.n227 B.n226 163.367
R405 B.n309 B.n196 163.367
R406 B.n315 B.n192 163.367
R407 B.n315 B.n190 163.367
R408 B.n319 B.n190 163.367
R409 B.n319 B.n184 163.367
R410 B.n328 B.n184 163.367
R411 B.n328 B.n182 163.367
R412 B.n332 B.n182 163.367
R413 B.n332 B.n177 163.367
R414 B.n340 B.n177 163.367
R415 B.n340 B.n175 163.367
R416 B.n344 B.n175 163.367
R417 B.n344 B.n169 163.367
R418 B.n352 B.n169 163.367
R419 B.n352 B.n167 163.367
R420 B.n356 B.n167 163.367
R421 B.n356 B.n161 163.367
R422 B.n365 B.n161 163.367
R423 B.n365 B.n159 163.367
R424 B.n369 B.n159 163.367
R425 B.n369 B.n3 163.367
R426 B.n450 B.n3 163.367
R427 B.n446 B.n2 163.367
R428 B.n446 B.n445 163.367
R429 B.n445 B.n9 163.367
R430 B.n441 B.n9 163.367
R431 B.n441 B.n11 163.367
R432 B.n437 B.n11 163.367
R433 B.n437 B.n17 163.367
R434 B.n433 B.n17 163.367
R435 B.n433 B.n19 163.367
R436 B.n429 B.n19 163.367
R437 B.n429 B.n24 163.367
R438 B.n425 B.n24 163.367
R439 B.n425 B.n26 163.367
R440 B.n421 B.n26 163.367
R441 B.n421 B.n30 163.367
R442 B.n417 B.n30 163.367
R443 B.n417 B.n32 163.367
R444 B.n413 B.n32 163.367
R445 B.n413 B.n38 163.367
R446 B.n409 B.n38 163.367
R447 B.n409 B.n40 163.367
R448 B.n308 B.n193 142.29
R449 B.n407 B.n406 142.29
R450 B.n66 B.t5 140.799
R451 B.n223 B.t14 140.799
R452 B.n68 B.t12 140.799
R453 B.n220 B.t8 140.799
R454 B.n314 B.n193 82.6981
R455 B.n314 B.n189 82.6981
R456 B.n320 B.n189 82.6981
R457 B.n320 B.n185 82.6981
R458 B.n327 B.n185 82.6981
R459 B.n327 B.n326 82.6981
R460 B.n333 B.n178 82.6981
R461 B.n339 B.n178 82.6981
R462 B.n339 B.n174 82.6981
R463 B.n345 B.n174 82.6981
R464 B.n345 B.n170 82.6981
R465 B.n351 B.n170 82.6981
R466 B.n351 B.n165 82.6981
R467 B.n357 B.n165 82.6981
R468 B.n357 B.n166 82.6981
R469 B.n364 B.n158 82.6981
R470 B.n370 B.n158 82.6981
R471 B.n370 B.n4 82.6981
R472 B.n449 B.n4 82.6981
R473 B.n449 B.n448 82.6981
R474 B.n448 B.n447 82.6981
R475 B.n447 B.n8 82.6981
R476 B.n12 B.n8 82.6981
R477 B.n440 B.n12 82.6981
R478 B.n439 B.n438 82.6981
R479 B.n438 B.n16 82.6981
R480 B.n432 B.n16 82.6981
R481 B.n432 B.n431 82.6981
R482 B.n431 B.n430 82.6981
R483 B.n430 B.n23 82.6981
R484 B.n424 B.n23 82.6981
R485 B.n424 B.n423 82.6981
R486 B.n423 B.n422 82.6981
R487 B.n416 B.n33 82.6981
R488 B.n416 B.n415 82.6981
R489 B.n415 B.n414 82.6981
R490 B.n414 B.n37 82.6981
R491 B.n408 B.n37 82.6981
R492 B.n408 B.n407 82.6981
R493 B.n69 B.n43 71.676
R494 B.n73 B.n44 71.676
R495 B.n77 B.n45 71.676
R496 B.n81 B.n46 71.676
R497 B.n85 B.n47 71.676
R498 B.n89 B.n48 71.676
R499 B.n93 B.n49 71.676
R500 B.n97 B.n50 71.676
R501 B.n101 B.n51 71.676
R502 B.n106 B.n52 71.676
R503 B.n110 B.n53 71.676
R504 B.n114 B.n54 71.676
R505 B.n118 B.n55 71.676
R506 B.n122 B.n56 71.676
R507 B.n127 B.n57 71.676
R508 B.n131 B.n58 71.676
R509 B.n135 B.n59 71.676
R510 B.n139 B.n60 71.676
R511 B.n143 B.n61 71.676
R512 B.n147 B.n62 71.676
R513 B.n151 B.n63 71.676
R514 B.n405 B.n64 71.676
R515 B.n405 B.n404 71.676
R516 B.n153 B.n63 71.676
R517 B.n150 B.n62 71.676
R518 B.n146 B.n61 71.676
R519 B.n142 B.n60 71.676
R520 B.n138 B.n59 71.676
R521 B.n134 B.n58 71.676
R522 B.n130 B.n57 71.676
R523 B.n126 B.n56 71.676
R524 B.n121 B.n55 71.676
R525 B.n117 B.n54 71.676
R526 B.n113 B.n53 71.676
R527 B.n109 B.n52 71.676
R528 B.n105 B.n51 71.676
R529 B.n100 B.n50 71.676
R530 B.n96 B.n49 71.676
R531 B.n92 B.n48 71.676
R532 B.n88 B.n47 71.676
R533 B.n84 B.n46 71.676
R534 B.n80 B.n45 71.676
R535 B.n76 B.n44 71.676
R536 B.n72 B.n43 71.676
R537 B.n307 B.n306 71.676
R538 B.n301 B.n197 71.676
R539 B.n298 B.n198 71.676
R540 B.n294 B.n199 71.676
R541 B.n290 B.n200 71.676
R542 B.n286 B.n201 71.676
R543 B.n282 B.n202 71.676
R544 B.n278 B.n203 71.676
R545 B.n274 B.n204 71.676
R546 B.n270 B.n205 71.676
R547 B.n266 B.n206 71.676
R548 B.n262 B.n207 71.676
R549 B.n258 B.n208 71.676
R550 B.n254 B.n209 71.676
R551 B.n250 B.n210 71.676
R552 B.n246 B.n211 71.676
R553 B.n242 B.n212 71.676
R554 B.n238 B.n213 71.676
R555 B.n234 B.n214 71.676
R556 B.n230 B.n215 71.676
R557 B.n226 B.n216 71.676
R558 B.n307 B.n218 71.676
R559 B.n299 B.n197 71.676
R560 B.n295 B.n198 71.676
R561 B.n291 B.n199 71.676
R562 B.n287 B.n200 71.676
R563 B.n283 B.n201 71.676
R564 B.n279 B.n202 71.676
R565 B.n275 B.n203 71.676
R566 B.n271 B.n204 71.676
R567 B.n267 B.n205 71.676
R568 B.n263 B.n206 71.676
R569 B.n259 B.n207 71.676
R570 B.n255 B.n208 71.676
R571 B.n251 B.n209 71.676
R572 B.n247 B.n210 71.676
R573 B.n243 B.n211 71.676
R574 B.n239 B.n212 71.676
R575 B.n235 B.n213 71.676
R576 B.n231 B.n214 71.676
R577 B.n227 B.n215 71.676
R578 B.n216 B.n196 71.676
R579 B.n451 B.n450 71.676
R580 B.n451 B.n2 71.676
R581 B.n326 B.t7 59.5914
R582 B.n33 B.t3 59.5914
R583 B.n103 B.n68 59.5399
R584 B.n124 B.n66 59.5399
R585 B.n224 B.n223 59.5399
R586 B.n221 B.n220 59.5399
R587 B.n166 B.t0 47.43
R588 B.t1 B.n439 47.43
R589 B.n68 B.n67 43.8308
R590 B.n66 B.n65 43.8308
R591 B.n223 B.n222 43.8308
R592 B.n220 B.n219 43.8308
R593 B.n364 B.t0 35.2686
R594 B.n440 B.t1 35.2686
R595 B.n305 B.n191 33.5615
R596 B.n311 B.n310 33.5615
R597 B.n403 B.n402 33.5615
R598 B.n70 B.n39 33.5615
R599 B.n333 B.t7 23.1072
R600 B.n422 B.t3 23.1072
R601 B B.n452 18.0485
R602 B.n316 B.n191 10.6151
R603 B.n317 B.n316 10.6151
R604 B.n318 B.n317 10.6151
R605 B.n318 B.n183 10.6151
R606 B.n329 B.n183 10.6151
R607 B.n330 B.n329 10.6151
R608 B.n331 B.n330 10.6151
R609 B.n331 B.n176 10.6151
R610 B.n341 B.n176 10.6151
R611 B.n342 B.n341 10.6151
R612 B.n343 B.n342 10.6151
R613 B.n343 B.n168 10.6151
R614 B.n353 B.n168 10.6151
R615 B.n354 B.n353 10.6151
R616 B.n355 B.n354 10.6151
R617 B.n355 B.n160 10.6151
R618 B.n366 B.n160 10.6151
R619 B.n367 B.n366 10.6151
R620 B.n368 B.n367 10.6151
R621 B.n368 B.n0 10.6151
R622 B.n305 B.n304 10.6151
R623 B.n304 B.n303 10.6151
R624 B.n303 B.n302 10.6151
R625 B.n302 B.n300 10.6151
R626 B.n300 B.n297 10.6151
R627 B.n297 B.n296 10.6151
R628 B.n296 B.n293 10.6151
R629 B.n293 B.n292 10.6151
R630 B.n292 B.n289 10.6151
R631 B.n289 B.n288 10.6151
R632 B.n288 B.n285 10.6151
R633 B.n285 B.n284 10.6151
R634 B.n284 B.n281 10.6151
R635 B.n281 B.n280 10.6151
R636 B.n280 B.n277 10.6151
R637 B.n277 B.n276 10.6151
R638 B.n273 B.n272 10.6151
R639 B.n272 B.n269 10.6151
R640 B.n269 B.n268 10.6151
R641 B.n268 B.n265 10.6151
R642 B.n265 B.n264 10.6151
R643 B.n264 B.n261 10.6151
R644 B.n261 B.n260 10.6151
R645 B.n260 B.n257 10.6151
R646 B.n257 B.n256 10.6151
R647 B.n253 B.n252 10.6151
R648 B.n252 B.n249 10.6151
R649 B.n249 B.n248 10.6151
R650 B.n248 B.n245 10.6151
R651 B.n245 B.n244 10.6151
R652 B.n244 B.n241 10.6151
R653 B.n241 B.n240 10.6151
R654 B.n240 B.n237 10.6151
R655 B.n237 B.n236 10.6151
R656 B.n236 B.n233 10.6151
R657 B.n233 B.n232 10.6151
R658 B.n232 B.n229 10.6151
R659 B.n229 B.n228 10.6151
R660 B.n228 B.n225 10.6151
R661 B.n225 B.n195 10.6151
R662 B.n310 B.n195 10.6151
R663 B.n312 B.n311 10.6151
R664 B.n312 B.n187 10.6151
R665 B.n322 B.n187 10.6151
R666 B.n323 B.n322 10.6151
R667 B.n324 B.n323 10.6151
R668 B.n324 B.n180 10.6151
R669 B.n335 B.n180 10.6151
R670 B.n336 B.n335 10.6151
R671 B.n337 B.n336 10.6151
R672 B.n337 B.n172 10.6151
R673 B.n347 B.n172 10.6151
R674 B.n348 B.n347 10.6151
R675 B.n349 B.n348 10.6151
R676 B.n349 B.n163 10.6151
R677 B.n359 B.n163 10.6151
R678 B.n360 B.n359 10.6151
R679 B.n362 B.n360 10.6151
R680 B.n362 B.n361 10.6151
R681 B.n361 B.n156 10.6151
R682 B.n373 B.n156 10.6151
R683 B.n374 B.n373 10.6151
R684 B.n375 B.n374 10.6151
R685 B.n376 B.n375 10.6151
R686 B.n377 B.n376 10.6151
R687 B.n380 B.n377 10.6151
R688 B.n381 B.n380 10.6151
R689 B.n382 B.n381 10.6151
R690 B.n383 B.n382 10.6151
R691 B.n385 B.n383 10.6151
R692 B.n386 B.n385 10.6151
R693 B.n387 B.n386 10.6151
R694 B.n388 B.n387 10.6151
R695 B.n390 B.n388 10.6151
R696 B.n391 B.n390 10.6151
R697 B.n392 B.n391 10.6151
R698 B.n393 B.n392 10.6151
R699 B.n395 B.n393 10.6151
R700 B.n396 B.n395 10.6151
R701 B.n397 B.n396 10.6151
R702 B.n398 B.n397 10.6151
R703 B.n400 B.n398 10.6151
R704 B.n401 B.n400 10.6151
R705 B.n402 B.n401 10.6151
R706 B.n444 B.n1 10.6151
R707 B.n444 B.n443 10.6151
R708 B.n443 B.n442 10.6151
R709 B.n442 B.n10 10.6151
R710 B.n436 B.n10 10.6151
R711 B.n436 B.n435 10.6151
R712 B.n435 B.n434 10.6151
R713 B.n434 B.n18 10.6151
R714 B.n428 B.n18 10.6151
R715 B.n428 B.n427 10.6151
R716 B.n427 B.n426 10.6151
R717 B.n426 B.n25 10.6151
R718 B.n420 B.n25 10.6151
R719 B.n420 B.n419 10.6151
R720 B.n419 B.n418 10.6151
R721 B.n418 B.n31 10.6151
R722 B.n412 B.n31 10.6151
R723 B.n412 B.n411 10.6151
R724 B.n411 B.n410 10.6151
R725 B.n410 B.n39 10.6151
R726 B.n71 B.n70 10.6151
R727 B.n74 B.n71 10.6151
R728 B.n75 B.n74 10.6151
R729 B.n78 B.n75 10.6151
R730 B.n79 B.n78 10.6151
R731 B.n82 B.n79 10.6151
R732 B.n83 B.n82 10.6151
R733 B.n86 B.n83 10.6151
R734 B.n87 B.n86 10.6151
R735 B.n90 B.n87 10.6151
R736 B.n91 B.n90 10.6151
R737 B.n94 B.n91 10.6151
R738 B.n95 B.n94 10.6151
R739 B.n98 B.n95 10.6151
R740 B.n99 B.n98 10.6151
R741 B.n102 B.n99 10.6151
R742 B.n107 B.n104 10.6151
R743 B.n108 B.n107 10.6151
R744 B.n111 B.n108 10.6151
R745 B.n112 B.n111 10.6151
R746 B.n115 B.n112 10.6151
R747 B.n116 B.n115 10.6151
R748 B.n119 B.n116 10.6151
R749 B.n120 B.n119 10.6151
R750 B.n123 B.n120 10.6151
R751 B.n128 B.n125 10.6151
R752 B.n129 B.n128 10.6151
R753 B.n132 B.n129 10.6151
R754 B.n133 B.n132 10.6151
R755 B.n136 B.n133 10.6151
R756 B.n137 B.n136 10.6151
R757 B.n140 B.n137 10.6151
R758 B.n141 B.n140 10.6151
R759 B.n144 B.n141 10.6151
R760 B.n145 B.n144 10.6151
R761 B.n148 B.n145 10.6151
R762 B.n149 B.n148 10.6151
R763 B.n152 B.n149 10.6151
R764 B.n154 B.n152 10.6151
R765 B.n155 B.n154 10.6151
R766 B.n403 B.n155 10.6151
R767 B.n276 B.n221 9.36635
R768 B.n253 B.n224 9.36635
R769 B.n103 B.n102 9.36635
R770 B.n125 B.n124 9.36635
R771 B.n452 B.n0 8.11757
R772 B.n452 B.n1 8.11757
R773 B.n273 B.n221 1.24928
R774 B.n256 B.n224 1.24928
R775 B.n104 B.n103 1.24928
R776 B.n124 B.n123 1.24928
R777 VN VN.t1 142.774
R778 VN VN.t0 106.178
R779 VTAIL.n74 VTAIL.n60 289.615
R780 VTAIL.n14 VTAIL.n0 289.615
R781 VTAIL.n54 VTAIL.n40 289.615
R782 VTAIL.n34 VTAIL.n20 289.615
R783 VTAIL.n67 VTAIL.n66 185
R784 VTAIL.n64 VTAIL.n63 185
R785 VTAIL.n73 VTAIL.n72 185
R786 VTAIL.n75 VTAIL.n74 185
R787 VTAIL.n7 VTAIL.n6 185
R788 VTAIL.n4 VTAIL.n3 185
R789 VTAIL.n13 VTAIL.n12 185
R790 VTAIL.n15 VTAIL.n14 185
R791 VTAIL.n55 VTAIL.n54 185
R792 VTAIL.n53 VTAIL.n52 185
R793 VTAIL.n44 VTAIL.n43 185
R794 VTAIL.n47 VTAIL.n46 185
R795 VTAIL.n35 VTAIL.n34 185
R796 VTAIL.n33 VTAIL.n32 185
R797 VTAIL.n24 VTAIL.n23 185
R798 VTAIL.n27 VTAIL.n26 185
R799 VTAIL.t2 VTAIL.n65 147.888
R800 VTAIL.t1 VTAIL.n5 147.888
R801 VTAIL.t0 VTAIL.n45 147.888
R802 VTAIL.t3 VTAIL.n25 147.888
R803 VTAIL.n66 VTAIL.n63 104.615
R804 VTAIL.n73 VTAIL.n63 104.615
R805 VTAIL.n74 VTAIL.n73 104.615
R806 VTAIL.n6 VTAIL.n3 104.615
R807 VTAIL.n13 VTAIL.n3 104.615
R808 VTAIL.n14 VTAIL.n13 104.615
R809 VTAIL.n54 VTAIL.n53 104.615
R810 VTAIL.n53 VTAIL.n43 104.615
R811 VTAIL.n46 VTAIL.n43 104.615
R812 VTAIL.n34 VTAIL.n33 104.615
R813 VTAIL.n33 VTAIL.n23 104.615
R814 VTAIL.n26 VTAIL.n23 104.615
R815 VTAIL.n66 VTAIL.t2 52.3082
R816 VTAIL.n6 VTAIL.t1 52.3082
R817 VTAIL.n46 VTAIL.t0 52.3082
R818 VTAIL.n26 VTAIL.t3 52.3082
R819 VTAIL.n79 VTAIL.n78 30.8278
R820 VTAIL.n19 VTAIL.n18 30.8278
R821 VTAIL.n59 VTAIL.n58 30.8278
R822 VTAIL.n39 VTAIL.n38 30.8278
R823 VTAIL.n39 VTAIL.n19 19.5134
R824 VTAIL.n79 VTAIL.n59 17.5652
R825 VTAIL.n67 VTAIL.n65 15.6496
R826 VTAIL.n7 VTAIL.n5 15.6496
R827 VTAIL.n47 VTAIL.n45 15.6496
R828 VTAIL.n27 VTAIL.n25 15.6496
R829 VTAIL.n68 VTAIL.n64 12.8005
R830 VTAIL.n8 VTAIL.n4 12.8005
R831 VTAIL.n48 VTAIL.n44 12.8005
R832 VTAIL.n28 VTAIL.n24 12.8005
R833 VTAIL.n72 VTAIL.n71 12.0247
R834 VTAIL.n12 VTAIL.n11 12.0247
R835 VTAIL.n52 VTAIL.n51 12.0247
R836 VTAIL.n32 VTAIL.n31 12.0247
R837 VTAIL.n75 VTAIL.n62 11.249
R838 VTAIL.n15 VTAIL.n2 11.249
R839 VTAIL.n55 VTAIL.n42 11.249
R840 VTAIL.n35 VTAIL.n22 11.249
R841 VTAIL.n76 VTAIL.n60 10.4732
R842 VTAIL.n16 VTAIL.n0 10.4732
R843 VTAIL.n56 VTAIL.n40 10.4732
R844 VTAIL.n36 VTAIL.n20 10.4732
R845 VTAIL.n78 VTAIL.n77 9.45567
R846 VTAIL.n18 VTAIL.n17 9.45567
R847 VTAIL.n58 VTAIL.n57 9.45567
R848 VTAIL.n38 VTAIL.n37 9.45567
R849 VTAIL.n77 VTAIL.n76 9.3005
R850 VTAIL.n62 VTAIL.n61 9.3005
R851 VTAIL.n71 VTAIL.n70 9.3005
R852 VTAIL.n69 VTAIL.n68 9.3005
R853 VTAIL.n17 VTAIL.n16 9.3005
R854 VTAIL.n2 VTAIL.n1 9.3005
R855 VTAIL.n11 VTAIL.n10 9.3005
R856 VTAIL.n9 VTAIL.n8 9.3005
R857 VTAIL.n57 VTAIL.n56 9.3005
R858 VTAIL.n42 VTAIL.n41 9.3005
R859 VTAIL.n51 VTAIL.n50 9.3005
R860 VTAIL.n49 VTAIL.n48 9.3005
R861 VTAIL.n37 VTAIL.n36 9.3005
R862 VTAIL.n22 VTAIL.n21 9.3005
R863 VTAIL.n31 VTAIL.n30 9.3005
R864 VTAIL.n29 VTAIL.n28 9.3005
R865 VTAIL.n69 VTAIL.n65 4.40546
R866 VTAIL.n9 VTAIL.n5 4.40546
R867 VTAIL.n49 VTAIL.n45 4.40546
R868 VTAIL.n29 VTAIL.n25 4.40546
R869 VTAIL.n78 VTAIL.n60 3.49141
R870 VTAIL.n18 VTAIL.n0 3.49141
R871 VTAIL.n58 VTAIL.n40 3.49141
R872 VTAIL.n38 VTAIL.n20 3.49141
R873 VTAIL.n76 VTAIL.n75 2.71565
R874 VTAIL.n16 VTAIL.n15 2.71565
R875 VTAIL.n56 VTAIL.n55 2.71565
R876 VTAIL.n36 VTAIL.n35 2.71565
R877 VTAIL.n72 VTAIL.n62 1.93989
R878 VTAIL.n12 VTAIL.n2 1.93989
R879 VTAIL.n52 VTAIL.n42 1.93989
R880 VTAIL.n32 VTAIL.n22 1.93989
R881 VTAIL.n59 VTAIL.n39 1.44447
R882 VTAIL.n71 VTAIL.n64 1.16414
R883 VTAIL.n11 VTAIL.n4 1.16414
R884 VTAIL.n51 VTAIL.n44 1.16414
R885 VTAIL.n31 VTAIL.n24 1.16414
R886 VTAIL VTAIL.n19 1.01559
R887 VTAIL VTAIL.n79 0.429379
R888 VTAIL.n68 VTAIL.n67 0.388379
R889 VTAIL.n8 VTAIL.n7 0.388379
R890 VTAIL.n48 VTAIL.n47 0.388379
R891 VTAIL.n28 VTAIL.n27 0.388379
R892 VTAIL.n70 VTAIL.n69 0.155672
R893 VTAIL.n70 VTAIL.n61 0.155672
R894 VTAIL.n77 VTAIL.n61 0.155672
R895 VTAIL.n10 VTAIL.n9 0.155672
R896 VTAIL.n10 VTAIL.n1 0.155672
R897 VTAIL.n17 VTAIL.n1 0.155672
R898 VTAIL.n57 VTAIL.n41 0.155672
R899 VTAIL.n50 VTAIL.n41 0.155672
R900 VTAIL.n50 VTAIL.n49 0.155672
R901 VTAIL.n37 VTAIL.n21 0.155672
R902 VTAIL.n30 VTAIL.n21 0.155672
R903 VTAIL.n30 VTAIL.n29 0.155672
R904 VDD2.n33 VDD2.n19 289.615
R905 VDD2.n14 VDD2.n0 289.615
R906 VDD2.n34 VDD2.n33 185
R907 VDD2.n32 VDD2.n31 185
R908 VDD2.n23 VDD2.n22 185
R909 VDD2.n26 VDD2.n25 185
R910 VDD2.n7 VDD2.n6 185
R911 VDD2.n4 VDD2.n3 185
R912 VDD2.n13 VDD2.n12 185
R913 VDD2.n15 VDD2.n14 185
R914 VDD2.t0 VDD2.n24 147.888
R915 VDD2.t1 VDD2.n5 147.888
R916 VDD2.n33 VDD2.n32 104.615
R917 VDD2.n32 VDD2.n22 104.615
R918 VDD2.n25 VDD2.n22 104.615
R919 VDD2.n6 VDD2.n3 104.615
R920 VDD2.n13 VDD2.n3 104.615
R921 VDD2.n14 VDD2.n13 104.615
R922 VDD2.n38 VDD2.n18 78.3126
R923 VDD2.n25 VDD2.t0 52.3082
R924 VDD2.n6 VDD2.t1 52.3082
R925 VDD2.n38 VDD2.n37 47.5066
R926 VDD2.n26 VDD2.n24 15.6496
R927 VDD2.n7 VDD2.n5 15.6496
R928 VDD2.n27 VDD2.n23 12.8005
R929 VDD2.n8 VDD2.n4 12.8005
R930 VDD2.n31 VDD2.n30 12.0247
R931 VDD2.n12 VDD2.n11 12.0247
R932 VDD2.n34 VDD2.n21 11.249
R933 VDD2.n15 VDD2.n2 11.249
R934 VDD2.n35 VDD2.n19 10.4732
R935 VDD2.n16 VDD2.n0 10.4732
R936 VDD2.n37 VDD2.n36 9.45567
R937 VDD2.n18 VDD2.n17 9.45567
R938 VDD2.n36 VDD2.n35 9.3005
R939 VDD2.n21 VDD2.n20 9.3005
R940 VDD2.n30 VDD2.n29 9.3005
R941 VDD2.n28 VDD2.n27 9.3005
R942 VDD2.n17 VDD2.n16 9.3005
R943 VDD2.n2 VDD2.n1 9.3005
R944 VDD2.n11 VDD2.n10 9.3005
R945 VDD2.n9 VDD2.n8 9.3005
R946 VDD2.n28 VDD2.n24 4.40546
R947 VDD2.n9 VDD2.n5 4.40546
R948 VDD2.n37 VDD2.n19 3.49141
R949 VDD2.n18 VDD2.n0 3.49141
R950 VDD2.n35 VDD2.n34 2.71565
R951 VDD2.n16 VDD2.n15 2.71565
R952 VDD2.n31 VDD2.n21 1.93989
R953 VDD2.n12 VDD2.n2 1.93989
R954 VDD2.n30 VDD2.n23 1.16414
R955 VDD2.n11 VDD2.n4 1.16414
R956 VDD2 VDD2.n38 0.545759
R957 VDD2.n27 VDD2.n26 0.388379
R958 VDD2.n8 VDD2.n7 0.388379
R959 VDD2.n36 VDD2.n20 0.155672
R960 VDD2.n29 VDD2.n20 0.155672
R961 VDD2.n29 VDD2.n28 0.155672
R962 VDD2.n10 VDD2.n9 0.155672
R963 VDD2.n10 VDD2.n1 0.155672
R964 VDD2.n17 VDD2.n1 0.155672
R965 VP.n0 VP.t0 142.582
R966 VP.n0 VP.t1 105.938
R967 VP VP.n0 0.241678
R968 VDD1.n14 VDD1.n0 289.615
R969 VDD1.n33 VDD1.n19 289.615
R970 VDD1.n15 VDD1.n14 185
R971 VDD1.n13 VDD1.n12 185
R972 VDD1.n4 VDD1.n3 185
R973 VDD1.n7 VDD1.n6 185
R974 VDD1.n26 VDD1.n25 185
R975 VDD1.n23 VDD1.n22 185
R976 VDD1.n32 VDD1.n31 185
R977 VDD1.n34 VDD1.n33 185
R978 VDD1.t1 VDD1.n5 147.888
R979 VDD1.t0 VDD1.n24 147.888
R980 VDD1.n14 VDD1.n13 104.615
R981 VDD1.n13 VDD1.n3 104.615
R982 VDD1.n6 VDD1.n3 104.615
R983 VDD1.n25 VDD1.n22 104.615
R984 VDD1.n32 VDD1.n22 104.615
R985 VDD1.n33 VDD1.n32 104.615
R986 VDD1 VDD1.n37 79.3245
R987 VDD1.n6 VDD1.t1 52.3082
R988 VDD1.n25 VDD1.t0 52.3082
R989 VDD1 VDD1.n18 48.0518
R990 VDD1.n7 VDD1.n5 15.6496
R991 VDD1.n26 VDD1.n24 15.6496
R992 VDD1.n8 VDD1.n4 12.8005
R993 VDD1.n27 VDD1.n23 12.8005
R994 VDD1.n12 VDD1.n11 12.0247
R995 VDD1.n31 VDD1.n30 12.0247
R996 VDD1.n15 VDD1.n2 11.249
R997 VDD1.n34 VDD1.n21 11.249
R998 VDD1.n16 VDD1.n0 10.4732
R999 VDD1.n35 VDD1.n19 10.4732
R1000 VDD1.n18 VDD1.n17 9.45567
R1001 VDD1.n37 VDD1.n36 9.45567
R1002 VDD1.n17 VDD1.n16 9.3005
R1003 VDD1.n2 VDD1.n1 9.3005
R1004 VDD1.n11 VDD1.n10 9.3005
R1005 VDD1.n9 VDD1.n8 9.3005
R1006 VDD1.n36 VDD1.n35 9.3005
R1007 VDD1.n21 VDD1.n20 9.3005
R1008 VDD1.n30 VDD1.n29 9.3005
R1009 VDD1.n28 VDD1.n27 9.3005
R1010 VDD1.n9 VDD1.n5 4.40546
R1011 VDD1.n28 VDD1.n24 4.40546
R1012 VDD1.n18 VDD1.n0 3.49141
R1013 VDD1.n37 VDD1.n19 3.49141
R1014 VDD1.n16 VDD1.n15 2.71565
R1015 VDD1.n35 VDD1.n34 2.71565
R1016 VDD1.n12 VDD1.n2 1.93989
R1017 VDD1.n31 VDD1.n21 1.93989
R1018 VDD1.n11 VDD1.n4 1.16414
R1019 VDD1.n30 VDD1.n23 1.16414
R1020 VDD1.n8 VDD1.n7 0.388379
R1021 VDD1.n27 VDD1.n26 0.388379
R1022 VDD1.n17 VDD1.n1 0.155672
R1023 VDD1.n10 VDD1.n1 0.155672
R1024 VDD1.n10 VDD1.n9 0.155672
R1025 VDD1.n29 VDD1.n28 0.155672
R1026 VDD1.n29 VDD1.n20 0.155672
R1027 VDD1.n36 VDD1.n20 0.155672
C0 VN VDD1 0.152201f
C1 VTAIL VDD2 2.76119f
C2 VN VP 3.62183f
C3 VDD1 VDD2 0.593965f
C4 VTAIL VDD1 2.71345f
C5 VP VDD2 0.308945f
C6 VTAIL VP 1.0889f
C7 VDD1 VP 1.15616f
C8 VN VDD2 1.00098f
C9 VTAIL VN 1.07471f
C10 VDD2 B 2.68177f
C11 VDD1 B 4.11163f
C12 VTAIL B 3.540459f
C13 VN B 6.87798f
C14 VP B 4.85492f
C15 VDD1.n0 B 0.019141f
C16 VDD1.n1 B 0.014984f
C17 VDD1.n2 B 0.008052f
C18 VDD1.n3 B 0.019032f
C19 VDD1.n4 B 0.008526f
C20 VDD1.n5 B 0.056376f
C21 VDD1.t1 B 0.03131f
C22 VDD1.n6 B 0.014274f
C23 VDD1.n7 B 0.011201f
C24 VDD1.n8 B 0.008052f
C25 VDD1.n9 B 0.202397f
C26 VDD1.n10 B 0.014984f
C27 VDD1.n11 B 0.008052f
C28 VDD1.n12 B 0.008526f
C29 VDD1.n13 B 0.019032f
C30 VDD1.n14 B 0.037804f
C31 VDD1.n15 B 0.008526f
C32 VDD1.n16 B 0.008052f
C33 VDD1.n17 B 0.033202f
C34 VDD1.n18 B 0.031734f
C35 VDD1.n19 B 0.019141f
C36 VDD1.n20 B 0.014984f
C37 VDD1.n21 B 0.008052f
C38 VDD1.n22 B 0.019032f
C39 VDD1.n23 B 0.008526f
C40 VDD1.n24 B 0.056376f
C41 VDD1.t0 B 0.03131f
C42 VDD1.n25 B 0.014274f
C43 VDD1.n26 B 0.011201f
C44 VDD1.n27 B 0.008052f
C45 VDD1.n28 B 0.202397f
C46 VDD1.n29 B 0.014984f
C47 VDD1.n30 B 0.008052f
C48 VDD1.n31 B 0.008526f
C49 VDD1.n32 B 0.019032f
C50 VDD1.n33 B 0.037804f
C51 VDD1.n34 B 0.008526f
C52 VDD1.n35 B 0.008052f
C53 VDD1.n36 B 0.033202f
C54 VDD1.n37 B 0.281626f
C55 VP.t0 B 0.975967f
C56 VP.t1 B 0.69546f
C57 VP.n0 B 1.88498f
C58 VDD2.n0 B 0.020265f
C59 VDD2.n1 B 0.015864f
C60 VDD2.n2 B 0.008525f
C61 VDD2.n3 B 0.02015f
C62 VDD2.n4 B 0.009026f
C63 VDD2.n5 B 0.059687f
C64 VDD2.t1 B 0.03315f
C65 VDD2.n6 B 0.015112f
C66 VDD2.n7 B 0.011859f
C67 VDD2.n8 B 0.008525f
C68 VDD2.n9 B 0.214286f
C69 VDD2.n10 B 0.015864f
C70 VDD2.n11 B 0.008525f
C71 VDD2.n12 B 0.009026f
C72 VDD2.n13 B 0.02015f
C73 VDD2.n14 B 0.040024f
C74 VDD2.n15 B 0.009026f
C75 VDD2.n16 B 0.008525f
C76 VDD2.n17 B 0.035153f
C77 VDD2.n18 B 0.274893f
C78 VDD2.n19 B 0.020265f
C79 VDD2.n20 B 0.015864f
C80 VDD2.n21 B 0.008525f
C81 VDD2.n22 B 0.02015f
C82 VDD2.n23 B 0.009026f
C83 VDD2.n24 B 0.059687f
C84 VDD2.t0 B 0.03315f
C85 VDD2.n25 B 0.015112f
C86 VDD2.n26 B 0.011859f
C87 VDD2.n27 B 0.008525f
C88 VDD2.n28 B 0.214286f
C89 VDD2.n29 B 0.015864f
C90 VDD2.n30 B 0.008525f
C91 VDD2.n31 B 0.009026f
C92 VDD2.n32 B 0.02015f
C93 VDD2.n33 B 0.040024f
C94 VDD2.n34 B 0.009026f
C95 VDD2.n35 B 0.008525f
C96 VDD2.n36 B 0.035153f
C97 VDD2.n37 B 0.032945f
C98 VDD2.n38 B 1.28857f
C99 VTAIL.n0 B 0.023177f
C100 VTAIL.n1 B 0.018144f
C101 VTAIL.n2 B 0.00975f
C102 VTAIL.n3 B 0.023045f
C103 VTAIL.n4 B 0.010323f
C104 VTAIL.n5 B 0.068264f
C105 VTAIL.t1 B 0.037913f
C106 VTAIL.n6 B 0.017284f
C107 VTAIL.n7 B 0.013563f
C108 VTAIL.n8 B 0.00975f
C109 VTAIL.n9 B 0.245076f
C110 VTAIL.n10 B 0.018144f
C111 VTAIL.n11 B 0.00975f
C112 VTAIL.n12 B 0.010323f
C113 VTAIL.n13 B 0.023045f
C114 VTAIL.n14 B 0.045775f
C115 VTAIL.n15 B 0.010323f
C116 VTAIL.n16 B 0.00975f
C117 VTAIL.n17 B 0.040204f
C118 VTAIL.n18 B 0.025136f
C119 VTAIL.n19 B 0.738141f
C120 VTAIL.n20 B 0.023177f
C121 VTAIL.n21 B 0.018144f
C122 VTAIL.n22 B 0.00975f
C123 VTAIL.n23 B 0.023045f
C124 VTAIL.n24 B 0.010323f
C125 VTAIL.n25 B 0.068264f
C126 VTAIL.t3 B 0.037913f
C127 VTAIL.n26 B 0.017284f
C128 VTAIL.n27 B 0.013563f
C129 VTAIL.n28 B 0.00975f
C130 VTAIL.n29 B 0.245076f
C131 VTAIL.n30 B 0.018144f
C132 VTAIL.n31 B 0.00975f
C133 VTAIL.n32 B 0.010323f
C134 VTAIL.n33 B 0.023045f
C135 VTAIL.n34 B 0.045775f
C136 VTAIL.n35 B 0.010323f
C137 VTAIL.n36 B 0.00975f
C138 VTAIL.n37 B 0.040204f
C139 VTAIL.n38 B 0.025136f
C140 VTAIL.n39 B 0.763215f
C141 VTAIL.n40 B 0.023177f
C142 VTAIL.n41 B 0.018144f
C143 VTAIL.n42 B 0.00975f
C144 VTAIL.n43 B 0.023045f
C145 VTAIL.n44 B 0.010323f
C146 VTAIL.n45 B 0.068264f
C147 VTAIL.t0 B 0.037913f
C148 VTAIL.n46 B 0.017284f
C149 VTAIL.n47 B 0.013563f
C150 VTAIL.n48 B 0.00975f
C151 VTAIL.n49 B 0.245076f
C152 VTAIL.n50 B 0.018144f
C153 VTAIL.n51 B 0.00975f
C154 VTAIL.n52 B 0.010323f
C155 VTAIL.n53 B 0.023045f
C156 VTAIL.n54 B 0.045775f
C157 VTAIL.n55 B 0.010323f
C158 VTAIL.n56 B 0.00975f
C159 VTAIL.n57 B 0.040204f
C160 VTAIL.n58 B 0.025136f
C161 VTAIL.n59 B 0.649311f
C162 VTAIL.n60 B 0.023177f
C163 VTAIL.n61 B 0.018144f
C164 VTAIL.n62 B 0.00975f
C165 VTAIL.n63 B 0.023045f
C166 VTAIL.n64 B 0.010323f
C167 VTAIL.n65 B 0.068264f
C168 VTAIL.t2 B 0.037913f
C169 VTAIL.n66 B 0.017284f
C170 VTAIL.n67 B 0.013563f
C171 VTAIL.n68 B 0.00975f
C172 VTAIL.n69 B 0.245076f
C173 VTAIL.n70 B 0.018144f
C174 VTAIL.n71 B 0.00975f
C175 VTAIL.n72 B 0.010323f
C176 VTAIL.n73 B 0.023045f
C177 VTAIL.n74 B 0.045775f
C178 VTAIL.n75 B 0.010323f
C179 VTAIL.n76 B 0.00975f
C180 VTAIL.n77 B 0.040204f
C181 VTAIL.n78 B 0.025136f
C182 VTAIL.n79 B 0.589966f
C183 VN.t0 B 0.688773f
C184 VN.t1 B 0.970259f
.ends

