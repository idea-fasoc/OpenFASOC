// Decoder output to apply to DCO
//

module decode_dco(
    input prop_gain,
    output dc_swval,
    input dco_inval
);


endmodule : decode_dco
