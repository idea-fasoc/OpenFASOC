* NGSPICE file created from diff_pair_sample_1770.ext - technology: sky130A

.subckt diff_pair_sample_1770 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.95
X1 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=7.1565 ps=37.48 w=18.35 l=1.95
X2 VDD1.t1 VP.t0 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=7.1565 ps=37.48 w=18.35 l=1.95
X3 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=7.1565 ps=37.48 w=18.35 l=1.95
X4 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.95
X5 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.95
X6 VDD1.t0 VP.t1 VTAIL.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=7.1565 ps=37.48 w=18.35 l=1.95
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=7.1565 pd=37.48 as=0 ps=0 w=18.35 l=1.95
R0 B.n834 B.n833 585
R1 B.n370 B.n107 585
R2 B.n369 B.n368 585
R3 B.n367 B.n366 585
R4 B.n365 B.n364 585
R5 B.n363 B.n362 585
R6 B.n361 B.n360 585
R7 B.n359 B.n358 585
R8 B.n357 B.n356 585
R9 B.n355 B.n354 585
R10 B.n353 B.n352 585
R11 B.n351 B.n350 585
R12 B.n349 B.n348 585
R13 B.n347 B.n346 585
R14 B.n345 B.n344 585
R15 B.n343 B.n342 585
R16 B.n341 B.n340 585
R17 B.n339 B.n338 585
R18 B.n337 B.n336 585
R19 B.n335 B.n334 585
R20 B.n333 B.n332 585
R21 B.n331 B.n330 585
R22 B.n329 B.n328 585
R23 B.n327 B.n326 585
R24 B.n325 B.n324 585
R25 B.n323 B.n322 585
R26 B.n321 B.n320 585
R27 B.n319 B.n318 585
R28 B.n317 B.n316 585
R29 B.n315 B.n314 585
R30 B.n313 B.n312 585
R31 B.n311 B.n310 585
R32 B.n309 B.n308 585
R33 B.n307 B.n306 585
R34 B.n305 B.n304 585
R35 B.n303 B.n302 585
R36 B.n301 B.n300 585
R37 B.n299 B.n298 585
R38 B.n297 B.n296 585
R39 B.n295 B.n294 585
R40 B.n293 B.n292 585
R41 B.n291 B.n290 585
R42 B.n289 B.n288 585
R43 B.n287 B.n286 585
R44 B.n285 B.n284 585
R45 B.n283 B.n282 585
R46 B.n281 B.n280 585
R47 B.n279 B.n278 585
R48 B.n277 B.n276 585
R49 B.n275 B.n274 585
R50 B.n273 B.n272 585
R51 B.n271 B.n270 585
R52 B.n269 B.n268 585
R53 B.n267 B.n266 585
R54 B.n265 B.n264 585
R55 B.n263 B.n262 585
R56 B.n261 B.n260 585
R57 B.n259 B.n258 585
R58 B.n257 B.n256 585
R59 B.n255 B.n254 585
R60 B.n253 B.n252 585
R61 B.n251 B.n250 585
R62 B.n249 B.n248 585
R63 B.n247 B.n246 585
R64 B.n245 B.n244 585
R65 B.n243 B.n242 585
R66 B.n241 B.n240 585
R67 B.n239 B.n238 585
R68 B.n237 B.n236 585
R69 B.n235 B.n234 585
R70 B.n233 B.n232 585
R71 B.n231 B.n230 585
R72 B.n229 B.n228 585
R73 B.n227 B.n226 585
R74 B.n225 B.n224 585
R75 B.n223 B.n222 585
R76 B.n221 B.n220 585
R77 B.n219 B.n218 585
R78 B.n217 B.n216 585
R79 B.n215 B.n214 585
R80 B.n213 B.n212 585
R81 B.n211 B.n210 585
R82 B.n209 B.n208 585
R83 B.n207 B.n206 585
R84 B.n205 B.n204 585
R85 B.n203 B.n202 585
R86 B.n201 B.n200 585
R87 B.n199 B.n198 585
R88 B.n197 B.n196 585
R89 B.n195 B.n194 585
R90 B.n193 B.n192 585
R91 B.n191 B.n190 585
R92 B.n189 B.n188 585
R93 B.n187 B.n186 585
R94 B.n185 B.n184 585
R95 B.n183 B.n182 585
R96 B.n181 B.n180 585
R97 B.n179 B.n178 585
R98 B.n177 B.n176 585
R99 B.n175 B.n174 585
R100 B.n173 B.n172 585
R101 B.n171 B.n170 585
R102 B.n169 B.n168 585
R103 B.n167 B.n166 585
R104 B.n165 B.n164 585
R105 B.n163 B.n162 585
R106 B.n161 B.n160 585
R107 B.n159 B.n158 585
R108 B.n157 B.n156 585
R109 B.n155 B.n154 585
R110 B.n153 B.n152 585
R111 B.n151 B.n150 585
R112 B.n149 B.n148 585
R113 B.n147 B.n146 585
R114 B.n145 B.n144 585
R115 B.n143 B.n142 585
R116 B.n141 B.n140 585
R117 B.n139 B.n138 585
R118 B.n137 B.n136 585
R119 B.n135 B.n134 585
R120 B.n133 B.n132 585
R121 B.n131 B.n130 585
R122 B.n129 B.n128 585
R123 B.n127 B.n126 585
R124 B.n125 B.n124 585
R125 B.n123 B.n122 585
R126 B.n121 B.n120 585
R127 B.n119 B.n118 585
R128 B.n117 B.n116 585
R129 B.n115 B.n114 585
R130 B.n832 B.n42 585
R131 B.n837 B.n42 585
R132 B.n831 B.n41 585
R133 B.n838 B.n41 585
R134 B.n830 B.n829 585
R135 B.n829 B.n37 585
R136 B.n828 B.n36 585
R137 B.n844 B.n36 585
R138 B.n827 B.n35 585
R139 B.n845 B.n35 585
R140 B.n826 B.n34 585
R141 B.n846 B.n34 585
R142 B.n825 B.n824 585
R143 B.n824 B.n33 585
R144 B.n823 B.n29 585
R145 B.n852 B.n29 585
R146 B.n822 B.n28 585
R147 B.n853 B.n28 585
R148 B.n821 B.n27 585
R149 B.n854 B.n27 585
R150 B.n820 B.n819 585
R151 B.n819 B.n23 585
R152 B.n818 B.n22 585
R153 B.n860 B.n22 585
R154 B.n817 B.n21 585
R155 B.n861 B.n21 585
R156 B.n816 B.n20 585
R157 B.n862 B.n20 585
R158 B.n815 B.n814 585
R159 B.n814 B.n16 585
R160 B.n813 B.n15 585
R161 B.n868 B.n15 585
R162 B.n812 B.n14 585
R163 B.n869 B.n14 585
R164 B.n811 B.n13 585
R165 B.n870 B.n13 585
R166 B.n810 B.n809 585
R167 B.n809 B.n12 585
R168 B.n808 B.n807 585
R169 B.n808 B.n8 585
R170 B.n806 B.n7 585
R171 B.n877 B.n7 585
R172 B.n805 B.n6 585
R173 B.n878 B.n6 585
R174 B.n804 B.n5 585
R175 B.n879 B.n5 585
R176 B.n803 B.n802 585
R177 B.n802 B.n4 585
R178 B.n801 B.n371 585
R179 B.n801 B.n800 585
R180 B.n791 B.n372 585
R181 B.n373 B.n372 585
R182 B.n793 B.n792 585
R183 B.n794 B.n793 585
R184 B.n790 B.n377 585
R185 B.n381 B.n377 585
R186 B.n789 B.n788 585
R187 B.n788 B.n787 585
R188 B.n379 B.n378 585
R189 B.n380 B.n379 585
R190 B.n780 B.n779 585
R191 B.n781 B.n780 585
R192 B.n778 B.n386 585
R193 B.n386 B.n385 585
R194 B.n777 B.n776 585
R195 B.n776 B.n775 585
R196 B.n388 B.n387 585
R197 B.n389 B.n388 585
R198 B.n768 B.n767 585
R199 B.n769 B.n768 585
R200 B.n766 B.n394 585
R201 B.n394 B.n393 585
R202 B.n765 B.n764 585
R203 B.n764 B.n763 585
R204 B.n396 B.n395 585
R205 B.n756 B.n396 585
R206 B.n755 B.n754 585
R207 B.n757 B.n755 585
R208 B.n753 B.n401 585
R209 B.n401 B.n400 585
R210 B.n752 B.n751 585
R211 B.n751 B.n750 585
R212 B.n403 B.n402 585
R213 B.n404 B.n403 585
R214 B.n743 B.n742 585
R215 B.n744 B.n743 585
R216 B.n741 B.n409 585
R217 B.n409 B.n408 585
R218 B.n736 B.n735 585
R219 B.n734 B.n476 585
R220 B.n733 B.n475 585
R221 B.n738 B.n475 585
R222 B.n732 B.n731 585
R223 B.n730 B.n729 585
R224 B.n728 B.n727 585
R225 B.n726 B.n725 585
R226 B.n724 B.n723 585
R227 B.n722 B.n721 585
R228 B.n720 B.n719 585
R229 B.n718 B.n717 585
R230 B.n716 B.n715 585
R231 B.n714 B.n713 585
R232 B.n712 B.n711 585
R233 B.n710 B.n709 585
R234 B.n708 B.n707 585
R235 B.n706 B.n705 585
R236 B.n704 B.n703 585
R237 B.n702 B.n701 585
R238 B.n700 B.n699 585
R239 B.n698 B.n697 585
R240 B.n696 B.n695 585
R241 B.n694 B.n693 585
R242 B.n692 B.n691 585
R243 B.n690 B.n689 585
R244 B.n688 B.n687 585
R245 B.n686 B.n685 585
R246 B.n684 B.n683 585
R247 B.n682 B.n681 585
R248 B.n680 B.n679 585
R249 B.n678 B.n677 585
R250 B.n676 B.n675 585
R251 B.n674 B.n673 585
R252 B.n672 B.n671 585
R253 B.n670 B.n669 585
R254 B.n668 B.n667 585
R255 B.n666 B.n665 585
R256 B.n664 B.n663 585
R257 B.n662 B.n661 585
R258 B.n660 B.n659 585
R259 B.n658 B.n657 585
R260 B.n656 B.n655 585
R261 B.n654 B.n653 585
R262 B.n652 B.n651 585
R263 B.n650 B.n649 585
R264 B.n648 B.n647 585
R265 B.n646 B.n645 585
R266 B.n644 B.n643 585
R267 B.n642 B.n641 585
R268 B.n640 B.n639 585
R269 B.n638 B.n637 585
R270 B.n636 B.n635 585
R271 B.n634 B.n633 585
R272 B.n632 B.n631 585
R273 B.n630 B.n629 585
R274 B.n628 B.n627 585
R275 B.n626 B.n625 585
R276 B.n624 B.n623 585
R277 B.n622 B.n621 585
R278 B.n620 B.n619 585
R279 B.n617 B.n616 585
R280 B.n615 B.n614 585
R281 B.n613 B.n612 585
R282 B.n611 B.n610 585
R283 B.n609 B.n608 585
R284 B.n607 B.n606 585
R285 B.n605 B.n604 585
R286 B.n603 B.n602 585
R287 B.n601 B.n600 585
R288 B.n599 B.n598 585
R289 B.n596 B.n595 585
R290 B.n594 B.n593 585
R291 B.n592 B.n591 585
R292 B.n590 B.n589 585
R293 B.n588 B.n587 585
R294 B.n586 B.n585 585
R295 B.n584 B.n583 585
R296 B.n582 B.n581 585
R297 B.n580 B.n579 585
R298 B.n578 B.n577 585
R299 B.n576 B.n575 585
R300 B.n574 B.n573 585
R301 B.n572 B.n571 585
R302 B.n570 B.n569 585
R303 B.n568 B.n567 585
R304 B.n566 B.n565 585
R305 B.n564 B.n563 585
R306 B.n562 B.n561 585
R307 B.n560 B.n559 585
R308 B.n558 B.n557 585
R309 B.n556 B.n555 585
R310 B.n554 B.n553 585
R311 B.n552 B.n551 585
R312 B.n550 B.n549 585
R313 B.n548 B.n547 585
R314 B.n546 B.n545 585
R315 B.n544 B.n543 585
R316 B.n542 B.n541 585
R317 B.n540 B.n539 585
R318 B.n538 B.n537 585
R319 B.n536 B.n535 585
R320 B.n534 B.n533 585
R321 B.n532 B.n531 585
R322 B.n530 B.n529 585
R323 B.n528 B.n527 585
R324 B.n526 B.n525 585
R325 B.n524 B.n523 585
R326 B.n522 B.n521 585
R327 B.n520 B.n519 585
R328 B.n518 B.n517 585
R329 B.n516 B.n515 585
R330 B.n514 B.n513 585
R331 B.n512 B.n511 585
R332 B.n510 B.n509 585
R333 B.n508 B.n507 585
R334 B.n506 B.n505 585
R335 B.n504 B.n503 585
R336 B.n502 B.n501 585
R337 B.n500 B.n499 585
R338 B.n498 B.n497 585
R339 B.n496 B.n495 585
R340 B.n494 B.n493 585
R341 B.n492 B.n491 585
R342 B.n490 B.n489 585
R343 B.n488 B.n487 585
R344 B.n486 B.n485 585
R345 B.n484 B.n483 585
R346 B.n482 B.n481 585
R347 B.n411 B.n410 585
R348 B.n740 B.n739 585
R349 B.n739 B.n738 585
R350 B.n407 B.n406 585
R351 B.n408 B.n407 585
R352 B.n746 B.n745 585
R353 B.n745 B.n744 585
R354 B.n747 B.n405 585
R355 B.n405 B.n404 585
R356 B.n749 B.n748 585
R357 B.n750 B.n749 585
R358 B.n399 B.n398 585
R359 B.n400 B.n399 585
R360 B.n759 B.n758 585
R361 B.n758 B.n757 585
R362 B.n760 B.n397 585
R363 B.n756 B.n397 585
R364 B.n762 B.n761 585
R365 B.n763 B.n762 585
R366 B.n392 B.n391 585
R367 B.n393 B.n392 585
R368 B.n771 B.n770 585
R369 B.n770 B.n769 585
R370 B.n772 B.n390 585
R371 B.n390 B.n389 585
R372 B.n774 B.n773 585
R373 B.n775 B.n774 585
R374 B.n384 B.n383 585
R375 B.n385 B.n384 585
R376 B.n783 B.n782 585
R377 B.n782 B.n781 585
R378 B.n784 B.n382 585
R379 B.n382 B.n380 585
R380 B.n786 B.n785 585
R381 B.n787 B.n786 585
R382 B.n376 B.n375 585
R383 B.n381 B.n376 585
R384 B.n796 B.n795 585
R385 B.n795 B.n794 585
R386 B.n797 B.n374 585
R387 B.n374 B.n373 585
R388 B.n799 B.n798 585
R389 B.n800 B.n799 585
R390 B.n3 B.n0 585
R391 B.n4 B.n3 585
R392 B.n876 B.n1 585
R393 B.n877 B.n876 585
R394 B.n875 B.n874 585
R395 B.n875 B.n8 585
R396 B.n873 B.n9 585
R397 B.n12 B.n9 585
R398 B.n872 B.n871 585
R399 B.n871 B.n870 585
R400 B.n11 B.n10 585
R401 B.n869 B.n11 585
R402 B.n867 B.n866 585
R403 B.n868 B.n867 585
R404 B.n865 B.n17 585
R405 B.n17 B.n16 585
R406 B.n864 B.n863 585
R407 B.n863 B.n862 585
R408 B.n19 B.n18 585
R409 B.n861 B.n19 585
R410 B.n859 B.n858 585
R411 B.n860 B.n859 585
R412 B.n857 B.n24 585
R413 B.n24 B.n23 585
R414 B.n856 B.n855 585
R415 B.n855 B.n854 585
R416 B.n26 B.n25 585
R417 B.n853 B.n26 585
R418 B.n851 B.n850 585
R419 B.n852 B.n851 585
R420 B.n849 B.n30 585
R421 B.n33 B.n30 585
R422 B.n848 B.n847 585
R423 B.n847 B.n846 585
R424 B.n32 B.n31 585
R425 B.n845 B.n32 585
R426 B.n843 B.n842 585
R427 B.n844 B.n843 585
R428 B.n841 B.n38 585
R429 B.n38 B.n37 585
R430 B.n840 B.n839 585
R431 B.n839 B.n838 585
R432 B.n40 B.n39 585
R433 B.n837 B.n40 585
R434 B.n880 B.n879 585
R435 B.n878 B.n2 585
R436 B.n114 B.n40 516.524
R437 B.n834 B.n42 516.524
R438 B.n739 B.n409 516.524
R439 B.n736 B.n407 516.524
R440 B.n108 B.t4 436.099
R441 B.n479 B.t12 436.099
R442 B.n111 B.t7 436.099
R443 B.n477 B.t15 436.099
R444 B.n111 B.t6 433.586
R445 B.n108 B.t2 433.586
R446 B.n479 B.t9 433.586
R447 B.n477 B.t13 433.586
R448 B.n109 B.t5 391.88
R449 B.n480 B.t11 391.88
R450 B.n112 B.t8 391.88
R451 B.n478 B.t14 391.88
R452 B.n836 B.n835 256.663
R453 B.n836 B.n106 256.663
R454 B.n836 B.n105 256.663
R455 B.n836 B.n104 256.663
R456 B.n836 B.n103 256.663
R457 B.n836 B.n102 256.663
R458 B.n836 B.n101 256.663
R459 B.n836 B.n100 256.663
R460 B.n836 B.n99 256.663
R461 B.n836 B.n98 256.663
R462 B.n836 B.n97 256.663
R463 B.n836 B.n96 256.663
R464 B.n836 B.n95 256.663
R465 B.n836 B.n94 256.663
R466 B.n836 B.n93 256.663
R467 B.n836 B.n92 256.663
R468 B.n836 B.n91 256.663
R469 B.n836 B.n90 256.663
R470 B.n836 B.n89 256.663
R471 B.n836 B.n88 256.663
R472 B.n836 B.n87 256.663
R473 B.n836 B.n86 256.663
R474 B.n836 B.n85 256.663
R475 B.n836 B.n84 256.663
R476 B.n836 B.n83 256.663
R477 B.n836 B.n82 256.663
R478 B.n836 B.n81 256.663
R479 B.n836 B.n80 256.663
R480 B.n836 B.n79 256.663
R481 B.n836 B.n78 256.663
R482 B.n836 B.n77 256.663
R483 B.n836 B.n76 256.663
R484 B.n836 B.n75 256.663
R485 B.n836 B.n74 256.663
R486 B.n836 B.n73 256.663
R487 B.n836 B.n72 256.663
R488 B.n836 B.n71 256.663
R489 B.n836 B.n70 256.663
R490 B.n836 B.n69 256.663
R491 B.n836 B.n68 256.663
R492 B.n836 B.n67 256.663
R493 B.n836 B.n66 256.663
R494 B.n836 B.n65 256.663
R495 B.n836 B.n64 256.663
R496 B.n836 B.n63 256.663
R497 B.n836 B.n62 256.663
R498 B.n836 B.n61 256.663
R499 B.n836 B.n60 256.663
R500 B.n836 B.n59 256.663
R501 B.n836 B.n58 256.663
R502 B.n836 B.n57 256.663
R503 B.n836 B.n56 256.663
R504 B.n836 B.n55 256.663
R505 B.n836 B.n54 256.663
R506 B.n836 B.n53 256.663
R507 B.n836 B.n52 256.663
R508 B.n836 B.n51 256.663
R509 B.n836 B.n50 256.663
R510 B.n836 B.n49 256.663
R511 B.n836 B.n48 256.663
R512 B.n836 B.n47 256.663
R513 B.n836 B.n46 256.663
R514 B.n836 B.n45 256.663
R515 B.n836 B.n44 256.663
R516 B.n836 B.n43 256.663
R517 B.n738 B.n737 256.663
R518 B.n738 B.n412 256.663
R519 B.n738 B.n413 256.663
R520 B.n738 B.n414 256.663
R521 B.n738 B.n415 256.663
R522 B.n738 B.n416 256.663
R523 B.n738 B.n417 256.663
R524 B.n738 B.n418 256.663
R525 B.n738 B.n419 256.663
R526 B.n738 B.n420 256.663
R527 B.n738 B.n421 256.663
R528 B.n738 B.n422 256.663
R529 B.n738 B.n423 256.663
R530 B.n738 B.n424 256.663
R531 B.n738 B.n425 256.663
R532 B.n738 B.n426 256.663
R533 B.n738 B.n427 256.663
R534 B.n738 B.n428 256.663
R535 B.n738 B.n429 256.663
R536 B.n738 B.n430 256.663
R537 B.n738 B.n431 256.663
R538 B.n738 B.n432 256.663
R539 B.n738 B.n433 256.663
R540 B.n738 B.n434 256.663
R541 B.n738 B.n435 256.663
R542 B.n738 B.n436 256.663
R543 B.n738 B.n437 256.663
R544 B.n738 B.n438 256.663
R545 B.n738 B.n439 256.663
R546 B.n738 B.n440 256.663
R547 B.n738 B.n441 256.663
R548 B.n738 B.n442 256.663
R549 B.n738 B.n443 256.663
R550 B.n738 B.n444 256.663
R551 B.n738 B.n445 256.663
R552 B.n738 B.n446 256.663
R553 B.n738 B.n447 256.663
R554 B.n738 B.n448 256.663
R555 B.n738 B.n449 256.663
R556 B.n738 B.n450 256.663
R557 B.n738 B.n451 256.663
R558 B.n738 B.n452 256.663
R559 B.n738 B.n453 256.663
R560 B.n738 B.n454 256.663
R561 B.n738 B.n455 256.663
R562 B.n738 B.n456 256.663
R563 B.n738 B.n457 256.663
R564 B.n738 B.n458 256.663
R565 B.n738 B.n459 256.663
R566 B.n738 B.n460 256.663
R567 B.n738 B.n461 256.663
R568 B.n738 B.n462 256.663
R569 B.n738 B.n463 256.663
R570 B.n738 B.n464 256.663
R571 B.n738 B.n465 256.663
R572 B.n738 B.n466 256.663
R573 B.n738 B.n467 256.663
R574 B.n738 B.n468 256.663
R575 B.n738 B.n469 256.663
R576 B.n738 B.n470 256.663
R577 B.n738 B.n471 256.663
R578 B.n738 B.n472 256.663
R579 B.n738 B.n473 256.663
R580 B.n738 B.n474 256.663
R581 B.n882 B.n881 256.663
R582 B.n118 B.n117 163.367
R583 B.n122 B.n121 163.367
R584 B.n126 B.n125 163.367
R585 B.n130 B.n129 163.367
R586 B.n134 B.n133 163.367
R587 B.n138 B.n137 163.367
R588 B.n142 B.n141 163.367
R589 B.n146 B.n145 163.367
R590 B.n150 B.n149 163.367
R591 B.n154 B.n153 163.367
R592 B.n158 B.n157 163.367
R593 B.n162 B.n161 163.367
R594 B.n166 B.n165 163.367
R595 B.n170 B.n169 163.367
R596 B.n174 B.n173 163.367
R597 B.n178 B.n177 163.367
R598 B.n182 B.n181 163.367
R599 B.n186 B.n185 163.367
R600 B.n190 B.n189 163.367
R601 B.n194 B.n193 163.367
R602 B.n198 B.n197 163.367
R603 B.n202 B.n201 163.367
R604 B.n206 B.n205 163.367
R605 B.n210 B.n209 163.367
R606 B.n214 B.n213 163.367
R607 B.n218 B.n217 163.367
R608 B.n222 B.n221 163.367
R609 B.n226 B.n225 163.367
R610 B.n230 B.n229 163.367
R611 B.n234 B.n233 163.367
R612 B.n238 B.n237 163.367
R613 B.n242 B.n241 163.367
R614 B.n246 B.n245 163.367
R615 B.n250 B.n249 163.367
R616 B.n254 B.n253 163.367
R617 B.n258 B.n257 163.367
R618 B.n262 B.n261 163.367
R619 B.n266 B.n265 163.367
R620 B.n270 B.n269 163.367
R621 B.n274 B.n273 163.367
R622 B.n278 B.n277 163.367
R623 B.n282 B.n281 163.367
R624 B.n286 B.n285 163.367
R625 B.n290 B.n289 163.367
R626 B.n294 B.n293 163.367
R627 B.n298 B.n297 163.367
R628 B.n302 B.n301 163.367
R629 B.n306 B.n305 163.367
R630 B.n310 B.n309 163.367
R631 B.n314 B.n313 163.367
R632 B.n318 B.n317 163.367
R633 B.n322 B.n321 163.367
R634 B.n326 B.n325 163.367
R635 B.n330 B.n329 163.367
R636 B.n334 B.n333 163.367
R637 B.n338 B.n337 163.367
R638 B.n342 B.n341 163.367
R639 B.n346 B.n345 163.367
R640 B.n350 B.n349 163.367
R641 B.n354 B.n353 163.367
R642 B.n358 B.n357 163.367
R643 B.n362 B.n361 163.367
R644 B.n366 B.n365 163.367
R645 B.n368 B.n107 163.367
R646 B.n743 B.n409 163.367
R647 B.n743 B.n403 163.367
R648 B.n751 B.n403 163.367
R649 B.n751 B.n401 163.367
R650 B.n755 B.n401 163.367
R651 B.n755 B.n396 163.367
R652 B.n764 B.n396 163.367
R653 B.n764 B.n394 163.367
R654 B.n768 B.n394 163.367
R655 B.n768 B.n388 163.367
R656 B.n776 B.n388 163.367
R657 B.n776 B.n386 163.367
R658 B.n780 B.n386 163.367
R659 B.n780 B.n379 163.367
R660 B.n788 B.n379 163.367
R661 B.n788 B.n377 163.367
R662 B.n793 B.n377 163.367
R663 B.n793 B.n372 163.367
R664 B.n801 B.n372 163.367
R665 B.n802 B.n801 163.367
R666 B.n802 B.n5 163.367
R667 B.n6 B.n5 163.367
R668 B.n7 B.n6 163.367
R669 B.n808 B.n7 163.367
R670 B.n809 B.n808 163.367
R671 B.n809 B.n13 163.367
R672 B.n14 B.n13 163.367
R673 B.n15 B.n14 163.367
R674 B.n814 B.n15 163.367
R675 B.n814 B.n20 163.367
R676 B.n21 B.n20 163.367
R677 B.n22 B.n21 163.367
R678 B.n819 B.n22 163.367
R679 B.n819 B.n27 163.367
R680 B.n28 B.n27 163.367
R681 B.n29 B.n28 163.367
R682 B.n824 B.n29 163.367
R683 B.n824 B.n34 163.367
R684 B.n35 B.n34 163.367
R685 B.n36 B.n35 163.367
R686 B.n829 B.n36 163.367
R687 B.n829 B.n41 163.367
R688 B.n42 B.n41 163.367
R689 B.n476 B.n475 163.367
R690 B.n731 B.n475 163.367
R691 B.n729 B.n728 163.367
R692 B.n725 B.n724 163.367
R693 B.n721 B.n720 163.367
R694 B.n717 B.n716 163.367
R695 B.n713 B.n712 163.367
R696 B.n709 B.n708 163.367
R697 B.n705 B.n704 163.367
R698 B.n701 B.n700 163.367
R699 B.n697 B.n696 163.367
R700 B.n693 B.n692 163.367
R701 B.n689 B.n688 163.367
R702 B.n685 B.n684 163.367
R703 B.n681 B.n680 163.367
R704 B.n677 B.n676 163.367
R705 B.n673 B.n672 163.367
R706 B.n669 B.n668 163.367
R707 B.n665 B.n664 163.367
R708 B.n661 B.n660 163.367
R709 B.n657 B.n656 163.367
R710 B.n653 B.n652 163.367
R711 B.n649 B.n648 163.367
R712 B.n645 B.n644 163.367
R713 B.n641 B.n640 163.367
R714 B.n637 B.n636 163.367
R715 B.n633 B.n632 163.367
R716 B.n629 B.n628 163.367
R717 B.n625 B.n624 163.367
R718 B.n621 B.n620 163.367
R719 B.n616 B.n615 163.367
R720 B.n612 B.n611 163.367
R721 B.n608 B.n607 163.367
R722 B.n604 B.n603 163.367
R723 B.n600 B.n599 163.367
R724 B.n595 B.n594 163.367
R725 B.n591 B.n590 163.367
R726 B.n587 B.n586 163.367
R727 B.n583 B.n582 163.367
R728 B.n579 B.n578 163.367
R729 B.n575 B.n574 163.367
R730 B.n571 B.n570 163.367
R731 B.n567 B.n566 163.367
R732 B.n563 B.n562 163.367
R733 B.n559 B.n558 163.367
R734 B.n555 B.n554 163.367
R735 B.n551 B.n550 163.367
R736 B.n547 B.n546 163.367
R737 B.n543 B.n542 163.367
R738 B.n539 B.n538 163.367
R739 B.n535 B.n534 163.367
R740 B.n531 B.n530 163.367
R741 B.n527 B.n526 163.367
R742 B.n523 B.n522 163.367
R743 B.n519 B.n518 163.367
R744 B.n515 B.n514 163.367
R745 B.n511 B.n510 163.367
R746 B.n507 B.n506 163.367
R747 B.n503 B.n502 163.367
R748 B.n499 B.n498 163.367
R749 B.n495 B.n494 163.367
R750 B.n491 B.n490 163.367
R751 B.n487 B.n486 163.367
R752 B.n483 B.n482 163.367
R753 B.n739 B.n411 163.367
R754 B.n745 B.n407 163.367
R755 B.n745 B.n405 163.367
R756 B.n749 B.n405 163.367
R757 B.n749 B.n399 163.367
R758 B.n758 B.n399 163.367
R759 B.n758 B.n397 163.367
R760 B.n762 B.n397 163.367
R761 B.n762 B.n392 163.367
R762 B.n770 B.n392 163.367
R763 B.n770 B.n390 163.367
R764 B.n774 B.n390 163.367
R765 B.n774 B.n384 163.367
R766 B.n782 B.n384 163.367
R767 B.n782 B.n382 163.367
R768 B.n786 B.n382 163.367
R769 B.n786 B.n376 163.367
R770 B.n795 B.n376 163.367
R771 B.n795 B.n374 163.367
R772 B.n799 B.n374 163.367
R773 B.n799 B.n3 163.367
R774 B.n880 B.n3 163.367
R775 B.n876 B.n2 163.367
R776 B.n876 B.n875 163.367
R777 B.n875 B.n9 163.367
R778 B.n871 B.n9 163.367
R779 B.n871 B.n11 163.367
R780 B.n867 B.n11 163.367
R781 B.n867 B.n17 163.367
R782 B.n863 B.n17 163.367
R783 B.n863 B.n19 163.367
R784 B.n859 B.n19 163.367
R785 B.n859 B.n24 163.367
R786 B.n855 B.n24 163.367
R787 B.n855 B.n26 163.367
R788 B.n851 B.n26 163.367
R789 B.n851 B.n30 163.367
R790 B.n847 B.n30 163.367
R791 B.n847 B.n32 163.367
R792 B.n843 B.n32 163.367
R793 B.n843 B.n38 163.367
R794 B.n839 B.n38 163.367
R795 B.n839 B.n40 163.367
R796 B.n114 B.n43 71.676
R797 B.n118 B.n44 71.676
R798 B.n122 B.n45 71.676
R799 B.n126 B.n46 71.676
R800 B.n130 B.n47 71.676
R801 B.n134 B.n48 71.676
R802 B.n138 B.n49 71.676
R803 B.n142 B.n50 71.676
R804 B.n146 B.n51 71.676
R805 B.n150 B.n52 71.676
R806 B.n154 B.n53 71.676
R807 B.n158 B.n54 71.676
R808 B.n162 B.n55 71.676
R809 B.n166 B.n56 71.676
R810 B.n170 B.n57 71.676
R811 B.n174 B.n58 71.676
R812 B.n178 B.n59 71.676
R813 B.n182 B.n60 71.676
R814 B.n186 B.n61 71.676
R815 B.n190 B.n62 71.676
R816 B.n194 B.n63 71.676
R817 B.n198 B.n64 71.676
R818 B.n202 B.n65 71.676
R819 B.n206 B.n66 71.676
R820 B.n210 B.n67 71.676
R821 B.n214 B.n68 71.676
R822 B.n218 B.n69 71.676
R823 B.n222 B.n70 71.676
R824 B.n226 B.n71 71.676
R825 B.n230 B.n72 71.676
R826 B.n234 B.n73 71.676
R827 B.n238 B.n74 71.676
R828 B.n242 B.n75 71.676
R829 B.n246 B.n76 71.676
R830 B.n250 B.n77 71.676
R831 B.n254 B.n78 71.676
R832 B.n258 B.n79 71.676
R833 B.n262 B.n80 71.676
R834 B.n266 B.n81 71.676
R835 B.n270 B.n82 71.676
R836 B.n274 B.n83 71.676
R837 B.n278 B.n84 71.676
R838 B.n282 B.n85 71.676
R839 B.n286 B.n86 71.676
R840 B.n290 B.n87 71.676
R841 B.n294 B.n88 71.676
R842 B.n298 B.n89 71.676
R843 B.n302 B.n90 71.676
R844 B.n306 B.n91 71.676
R845 B.n310 B.n92 71.676
R846 B.n314 B.n93 71.676
R847 B.n318 B.n94 71.676
R848 B.n322 B.n95 71.676
R849 B.n326 B.n96 71.676
R850 B.n330 B.n97 71.676
R851 B.n334 B.n98 71.676
R852 B.n338 B.n99 71.676
R853 B.n342 B.n100 71.676
R854 B.n346 B.n101 71.676
R855 B.n350 B.n102 71.676
R856 B.n354 B.n103 71.676
R857 B.n358 B.n104 71.676
R858 B.n362 B.n105 71.676
R859 B.n366 B.n106 71.676
R860 B.n835 B.n107 71.676
R861 B.n835 B.n834 71.676
R862 B.n368 B.n106 71.676
R863 B.n365 B.n105 71.676
R864 B.n361 B.n104 71.676
R865 B.n357 B.n103 71.676
R866 B.n353 B.n102 71.676
R867 B.n349 B.n101 71.676
R868 B.n345 B.n100 71.676
R869 B.n341 B.n99 71.676
R870 B.n337 B.n98 71.676
R871 B.n333 B.n97 71.676
R872 B.n329 B.n96 71.676
R873 B.n325 B.n95 71.676
R874 B.n321 B.n94 71.676
R875 B.n317 B.n93 71.676
R876 B.n313 B.n92 71.676
R877 B.n309 B.n91 71.676
R878 B.n305 B.n90 71.676
R879 B.n301 B.n89 71.676
R880 B.n297 B.n88 71.676
R881 B.n293 B.n87 71.676
R882 B.n289 B.n86 71.676
R883 B.n285 B.n85 71.676
R884 B.n281 B.n84 71.676
R885 B.n277 B.n83 71.676
R886 B.n273 B.n82 71.676
R887 B.n269 B.n81 71.676
R888 B.n265 B.n80 71.676
R889 B.n261 B.n79 71.676
R890 B.n257 B.n78 71.676
R891 B.n253 B.n77 71.676
R892 B.n249 B.n76 71.676
R893 B.n245 B.n75 71.676
R894 B.n241 B.n74 71.676
R895 B.n237 B.n73 71.676
R896 B.n233 B.n72 71.676
R897 B.n229 B.n71 71.676
R898 B.n225 B.n70 71.676
R899 B.n221 B.n69 71.676
R900 B.n217 B.n68 71.676
R901 B.n213 B.n67 71.676
R902 B.n209 B.n66 71.676
R903 B.n205 B.n65 71.676
R904 B.n201 B.n64 71.676
R905 B.n197 B.n63 71.676
R906 B.n193 B.n62 71.676
R907 B.n189 B.n61 71.676
R908 B.n185 B.n60 71.676
R909 B.n181 B.n59 71.676
R910 B.n177 B.n58 71.676
R911 B.n173 B.n57 71.676
R912 B.n169 B.n56 71.676
R913 B.n165 B.n55 71.676
R914 B.n161 B.n54 71.676
R915 B.n157 B.n53 71.676
R916 B.n153 B.n52 71.676
R917 B.n149 B.n51 71.676
R918 B.n145 B.n50 71.676
R919 B.n141 B.n49 71.676
R920 B.n137 B.n48 71.676
R921 B.n133 B.n47 71.676
R922 B.n129 B.n46 71.676
R923 B.n125 B.n45 71.676
R924 B.n121 B.n44 71.676
R925 B.n117 B.n43 71.676
R926 B.n737 B.n736 71.676
R927 B.n731 B.n412 71.676
R928 B.n728 B.n413 71.676
R929 B.n724 B.n414 71.676
R930 B.n720 B.n415 71.676
R931 B.n716 B.n416 71.676
R932 B.n712 B.n417 71.676
R933 B.n708 B.n418 71.676
R934 B.n704 B.n419 71.676
R935 B.n700 B.n420 71.676
R936 B.n696 B.n421 71.676
R937 B.n692 B.n422 71.676
R938 B.n688 B.n423 71.676
R939 B.n684 B.n424 71.676
R940 B.n680 B.n425 71.676
R941 B.n676 B.n426 71.676
R942 B.n672 B.n427 71.676
R943 B.n668 B.n428 71.676
R944 B.n664 B.n429 71.676
R945 B.n660 B.n430 71.676
R946 B.n656 B.n431 71.676
R947 B.n652 B.n432 71.676
R948 B.n648 B.n433 71.676
R949 B.n644 B.n434 71.676
R950 B.n640 B.n435 71.676
R951 B.n636 B.n436 71.676
R952 B.n632 B.n437 71.676
R953 B.n628 B.n438 71.676
R954 B.n624 B.n439 71.676
R955 B.n620 B.n440 71.676
R956 B.n615 B.n441 71.676
R957 B.n611 B.n442 71.676
R958 B.n607 B.n443 71.676
R959 B.n603 B.n444 71.676
R960 B.n599 B.n445 71.676
R961 B.n594 B.n446 71.676
R962 B.n590 B.n447 71.676
R963 B.n586 B.n448 71.676
R964 B.n582 B.n449 71.676
R965 B.n578 B.n450 71.676
R966 B.n574 B.n451 71.676
R967 B.n570 B.n452 71.676
R968 B.n566 B.n453 71.676
R969 B.n562 B.n454 71.676
R970 B.n558 B.n455 71.676
R971 B.n554 B.n456 71.676
R972 B.n550 B.n457 71.676
R973 B.n546 B.n458 71.676
R974 B.n542 B.n459 71.676
R975 B.n538 B.n460 71.676
R976 B.n534 B.n461 71.676
R977 B.n530 B.n462 71.676
R978 B.n526 B.n463 71.676
R979 B.n522 B.n464 71.676
R980 B.n518 B.n465 71.676
R981 B.n514 B.n466 71.676
R982 B.n510 B.n467 71.676
R983 B.n506 B.n468 71.676
R984 B.n502 B.n469 71.676
R985 B.n498 B.n470 71.676
R986 B.n494 B.n471 71.676
R987 B.n490 B.n472 71.676
R988 B.n486 B.n473 71.676
R989 B.n482 B.n474 71.676
R990 B.n737 B.n476 71.676
R991 B.n729 B.n412 71.676
R992 B.n725 B.n413 71.676
R993 B.n721 B.n414 71.676
R994 B.n717 B.n415 71.676
R995 B.n713 B.n416 71.676
R996 B.n709 B.n417 71.676
R997 B.n705 B.n418 71.676
R998 B.n701 B.n419 71.676
R999 B.n697 B.n420 71.676
R1000 B.n693 B.n421 71.676
R1001 B.n689 B.n422 71.676
R1002 B.n685 B.n423 71.676
R1003 B.n681 B.n424 71.676
R1004 B.n677 B.n425 71.676
R1005 B.n673 B.n426 71.676
R1006 B.n669 B.n427 71.676
R1007 B.n665 B.n428 71.676
R1008 B.n661 B.n429 71.676
R1009 B.n657 B.n430 71.676
R1010 B.n653 B.n431 71.676
R1011 B.n649 B.n432 71.676
R1012 B.n645 B.n433 71.676
R1013 B.n641 B.n434 71.676
R1014 B.n637 B.n435 71.676
R1015 B.n633 B.n436 71.676
R1016 B.n629 B.n437 71.676
R1017 B.n625 B.n438 71.676
R1018 B.n621 B.n439 71.676
R1019 B.n616 B.n440 71.676
R1020 B.n612 B.n441 71.676
R1021 B.n608 B.n442 71.676
R1022 B.n604 B.n443 71.676
R1023 B.n600 B.n444 71.676
R1024 B.n595 B.n445 71.676
R1025 B.n591 B.n446 71.676
R1026 B.n587 B.n447 71.676
R1027 B.n583 B.n448 71.676
R1028 B.n579 B.n449 71.676
R1029 B.n575 B.n450 71.676
R1030 B.n571 B.n451 71.676
R1031 B.n567 B.n452 71.676
R1032 B.n563 B.n453 71.676
R1033 B.n559 B.n454 71.676
R1034 B.n555 B.n455 71.676
R1035 B.n551 B.n456 71.676
R1036 B.n547 B.n457 71.676
R1037 B.n543 B.n458 71.676
R1038 B.n539 B.n459 71.676
R1039 B.n535 B.n460 71.676
R1040 B.n531 B.n461 71.676
R1041 B.n527 B.n462 71.676
R1042 B.n523 B.n463 71.676
R1043 B.n519 B.n464 71.676
R1044 B.n515 B.n465 71.676
R1045 B.n511 B.n466 71.676
R1046 B.n507 B.n467 71.676
R1047 B.n503 B.n468 71.676
R1048 B.n499 B.n469 71.676
R1049 B.n495 B.n470 71.676
R1050 B.n491 B.n471 71.676
R1051 B.n487 B.n472 71.676
R1052 B.n483 B.n473 71.676
R1053 B.n474 B.n411 71.676
R1054 B.n881 B.n880 71.676
R1055 B.n881 B.n2 71.676
R1056 B.n113 B.n112 59.5399
R1057 B.n110 B.n109 59.5399
R1058 B.n597 B.n480 59.5399
R1059 B.n618 B.n478 59.5399
R1060 B.n738 B.n408 58.2016
R1061 B.n837 B.n836 58.2016
R1062 B.n112 B.n111 44.2187
R1063 B.n109 B.n108 44.2187
R1064 B.n480 B.n479 44.2187
R1065 B.n478 B.n477 44.2187
R1066 B.n735 B.n406 33.5615
R1067 B.n741 B.n740 33.5615
R1068 B.n833 B.n832 33.5615
R1069 B.n115 B.n39 33.5615
R1070 B.n744 B.n408 31.6619
R1071 B.n744 B.n404 31.6619
R1072 B.n750 B.n404 31.6619
R1073 B.n750 B.n400 31.6619
R1074 B.n757 B.n400 31.6619
R1075 B.n757 B.n756 31.6619
R1076 B.n763 B.n393 31.6619
R1077 B.n769 B.n393 31.6619
R1078 B.n769 B.n389 31.6619
R1079 B.n775 B.n389 31.6619
R1080 B.n775 B.n385 31.6619
R1081 B.n781 B.n385 31.6619
R1082 B.n781 B.n380 31.6619
R1083 B.n787 B.n380 31.6619
R1084 B.n787 B.n381 31.6619
R1085 B.n794 B.n373 31.6619
R1086 B.n800 B.n373 31.6619
R1087 B.n800 B.n4 31.6619
R1088 B.n879 B.n4 31.6619
R1089 B.n879 B.n878 31.6619
R1090 B.n878 B.n877 31.6619
R1091 B.n877 B.n8 31.6619
R1092 B.n12 B.n8 31.6619
R1093 B.n870 B.n12 31.6619
R1094 B.n869 B.n868 31.6619
R1095 B.n868 B.n16 31.6619
R1096 B.n862 B.n16 31.6619
R1097 B.n862 B.n861 31.6619
R1098 B.n861 B.n860 31.6619
R1099 B.n860 B.n23 31.6619
R1100 B.n854 B.n23 31.6619
R1101 B.n854 B.n853 31.6619
R1102 B.n853 B.n852 31.6619
R1103 B.n846 B.n33 31.6619
R1104 B.n846 B.n845 31.6619
R1105 B.n845 B.n844 31.6619
R1106 B.n844 B.n37 31.6619
R1107 B.n838 B.n37 31.6619
R1108 B.n838 B.n837 31.6619
R1109 B.n756 B.t10 20.0217
R1110 B.n33 B.t3 20.0217
R1111 B B.n882 18.0485
R1112 B.n381 B.t1 17.228
R1113 B.t0 B.n869 17.228
R1114 B.n794 B.t1 14.4344
R1115 B.n870 B.t0 14.4344
R1116 B.n763 B.t10 11.6407
R1117 B.n852 B.t3 11.6407
R1118 B.n746 B.n406 10.6151
R1119 B.n747 B.n746 10.6151
R1120 B.n748 B.n747 10.6151
R1121 B.n748 B.n398 10.6151
R1122 B.n759 B.n398 10.6151
R1123 B.n760 B.n759 10.6151
R1124 B.n761 B.n760 10.6151
R1125 B.n761 B.n391 10.6151
R1126 B.n771 B.n391 10.6151
R1127 B.n772 B.n771 10.6151
R1128 B.n773 B.n772 10.6151
R1129 B.n773 B.n383 10.6151
R1130 B.n783 B.n383 10.6151
R1131 B.n784 B.n783 10.6151
R1132 B.n785 B.n784 10.6151
R1133 B.n785 B.n375 10.6151
R1134 B.n796 B.n375 10.6151
R1135 B.n797 B.n796 10.6151
R1136 B.n798 B.n797 10.6151
R1137 B.n798 B.n0 10.6151
R1138 B.n735 B.n734 10.6151
R1139 B.n734 B.n733 10.6151
R1140 B.n733 B.n732 10.6151
R1141 B.n732 B.n730 10.6151
R1142 B.n730 B.n727 10.6151
R1143 B.n727 B.n726 10.6151
R1144 B.n726 B.n723 10.6151
R1145 B.n723 B.n722 10.6151
R1146 B.n722 B.n719 10.6151
R1147 B.n719 B.n718 10.6151
R1148 B.n718 B.n715 10.6151
R1149 B.n715 B.n714 10.6151
R1150 B.n714 B.n711 10.6151
R1151 B.n711 B.n710 10.6151
R1152 B.n710 B.n707 10.6151
R1153 B.n707 B.n706 10.6151
R1154 B.n706 B.n703 10.6151
R1155 B.n703 B.n702 10.6151
R1156 B.n702 B.n699 10.6151
R1157 B.n699 B.n698 10.6151
R1158 B.n698 B.n695 10.6151
R1159 B.n695 B.n694 10.6151
R1160 B.n694 B.n691 10.6151
R1161 B.n691 B.n690 10.6151
R1162 B.n690 B.n687 10.6151
R1163 B.n687 B.n686 10.6151
R1164 B.n686 B.n683 10.6151
R1165 B.n683 B.n682 10.6151
R1166 B.n682 B.n679 10.6151
R1167 B.n679 B.n678 10.6151
R1168 B.n678 B.n675 10.6151
R1169 B.n675 B.n674 10.6151
R1170 B.n674 B.n671 10.6151
R1171 B.n671 B.n670 10.6151
R1172 B.n670 B.n667 10.6151
R1173 B.n667 B.n666 10.6151
R1174 B.n666 B.n663 10.6151
R1175 B.n663 B.n662 10.6151
R1176 B.n662 B.n659 10.6151
R1177 B.n659 B.n658 10.6151
R1178 B.n658 B.n655 10.6151
R1179 B.n655 B.n654 10.6151
R1180 B.n654 B.n651 10.6151
R1181 B.n651 B.n650 10.6151
R1182 B.n650 B.n647 10.6151
R1183 B.n647 B.n646 10.6151
R1184 B.n646 B.n643 10.6151
R1185 B.n643 B.n642 10.6151
R1186 B.n642 B.n639 10.6151
R1187 B.n639 B.n638 10.6151
R1188 B.n638 B.n635 10.6151
R1189 B.n635 B.n634 10.6151
R1190 B.n634 B.n631 10.6151
R1191 B.n631 B.n630 10.6151
R1192 B.n630 B.n627 10.6151
R1193 B.n627 B.n626 10.6151
R1194 B.n626 B.n623 10.6151
R1195 B.n623 B.n622 10.6151
R1196 B.n622 B.n619 10.6151
R1197 B.n617 B.n614 10.6151
R1198 B.n614 B.n613 10.6151
R1199 B.n613 B.n610 10.6151
R1200 B.n610 B.n609 10.6151
R1201 B.n609 B.n606 10.6151
R1202 B.n606 B.n605 10.6151
R1203 B.n605 B.n602 10.6151
R1204 B.n602 B.n601 10.6151
R1205 B.n601 B.n598 10.6151
R1206 B.n596 B.n593 10.6151
R1207 B.n593 B.n592 10.6151
R1208 B.n592 B.n589 10.6151
R1209 B.n589 B.n588 10.6151
R1210 B.n588 B.n585 10.6151
R1211 B.n585 B.n584 10.6151
R1212 B.n584 B.n581 10.6151
R1213 B.n581 B.n580 10.6151
R1214 B.n580 B.n577 10.6151
R1215 B.n577 B.n576 10.6151
R1216 B.n576 B.n573 10.6151
R1217 B.n573 B.n572 10.6151
R1218 B.n572 B.n569 10.6151
R1219 B.n569 B.n568 10.6151
R1220 B.n568 B.n565 10.6151
R1221 B.n565 B.n564 10.6151
R1222 B.n564 B.n561 10.6151
R1223 B.n561 B.n560 10.6151
R1224 B.n560 B.n557 10.6151
R1225 B.n557 B.n556 10.6151
R1226 B.n556 B.n553 10.6151
R1227 B.n553 B.n552 10.6151
R1228 B.n552 B.n549 10.6151
R1229 B.n549 B.n548 10.6151
R1230 B.n548 B.n545 10.6151
R1231 B.n545 B.n544 10.6151
R1232 B.n544 B.n541 10.6151
R1233 B.n541 B.n540 10.6151
R1234 B.n540 B.n537 10.6151
R1235 B.n537 B.n536 10.6151
R1236 B.n536 B.n533 10.6151
R1237 B.n533 B.n532 10.6151
R1238 B.n532 B.n529 10.6151
R1239 B.n529 B.n528 10.6151
R1240 B.n528 B.n525 10.6151
R1241 B.n525 B.n524 10.6151
R1242 B.n524 B.n521 10.6151
R1243 B.n521 B.n520 10.6151
R1244 B.n520 B.n517 10.6151
R1245 B.n517 B.n516 10.6151
R1246 B.n516 B.n513 10.6151
R1247 B.n513 B.n512 10.6151
R1248 B.n512 B.n509 10.6151
R1249 B.n509 B.n508 10.6151
R1250 B.n508 B.n505 10.6151
R1251 B.n505 B.n504 10.6151
R1252 B.n504 B.n501 10.6151
R1253 B.n501 B.n500 10.6151
R1254 B.n500 B.n497 10.6151
R1255 B.n497 B.n496 10.6151
R1256 B.n496 B.n493 10.6151
R1257 B.n493 B.n492 10.6151
R1258 B.n492 B.n489 10.6151
R1259 B.n489 B.n488 10.6151
R1260 B.n488 B.n485 10.6151
R1261 B.n485 B.n484 10.6151
R1262 B.n484 B.n481 10.6151
R1263 B.n481 B.n410 10.6151
R1264 B.n740 B.n410 10.6151
R1265 B.n742 B.n741 10.6151
R1266 B.n742 B.n402 10.6151
R1267 B.n752 B.n402 10.6151
R1268 B.n753 B.n752 10.6151
R1269 B.n754 B.n753 10.6151
R1270 B.n754 B.n395 10.6151
R1271 B.n765 B.n395 10.6151
R1272 B.n766 B.n765 10.6151
R1273 B.n767 B.n766 10.6151
R1274 B.n767 B.n387 10.6151
R1275 B.n777 B.n387 10.6151
R1276 B.n778 B.n777 10.6151
R1277 B.n779 B.n778 10.6151
R1278 B.n779 B.n378 10.6151
R1279 B.n789 B.n378 10.6151
R1280 B.n790 B.n789 10.6151
R1281 B.n792 B.n790 10.6151
R1282 B.n792 B.n791 10.6151
R1283 B.n791 B.n371 10.6151
R1284 B.n803 B.n371 10.6151
R1285 B.n804 B.n803 10.6151
R1286 B.n805 B.n804 10.6151
R1287 B.n806 B.n805 10.6151
R1288 B.n807 B.n806 10.6151
R1289 B.n810 B.n807 10.6151
R1290 B.n811 B.n810 10.6151
R1291 B.n812 B.n811 10.6151
R1292 B.n813 B.n812 10.6151
R1293 B.n815 B.n813 10.6151
R1294 B.n816 B.n815 10.6151
R1295 B.n817 B.n816 10.6151
R1296 B.n818 B.n817 10.6151
R1297 B.n820 B.n818 10.6151
R1298 B.n821 B.n820 10.6151
R1299 B.n822 B.n821 10.6151
R1300 B.n823 B.n822 10.6151
R1301 B.n825 B.n823 10.6151
R1302 B.n826 B.n825 10.6151
R1303 B.n827 B.n826 10.6151
R1304 B.n828 B.n827 10.6151
R1305 B.n830 B.n828 10.6151
R1306 B.n831 B.n830 10.6151
R1307 B.n832 B.n831 10.6151
R1308 B.n874 B.n1 10.6151
R1309 B.n874 B.n873 10.6151
R1310 B.n873 B.n872 10.6151
R1311 B.n872 B.n10 10.6151
R1312 B.n866 B.n10 10.6151
R1313 B.n866 B.n865 10.6151
R1314 B.n865 B.n864 10.6151
R1315 B.n864 B.n18 10.6151
R1316 B.n858 B.n18 10.6151
R1317 B.n858 B.n857 10.6151
R1318 B.n857 B.n856 10.6151
R1319 B.n856 B.n25 10.6151
R1320 B.n850 B.n25 10.6151
R1321 B.n850 B.n849 10.6151
R1322 B.n849 B.n848 10.6151
R1323 B.n848 B.n31 10.6151
R1324 B.n842 B.n31 10.6151
R1325 B.n842 B.n841 10.6151
R1326 B.n841 B.n840 10.6151
R1327 B.n840 B.n39 10.6151
R1328 B.n116 B.n115 10.6151
R1329 B.n119 B.n116 10.6151
R1330 B.n120 B.n119 10.6151
R1331 B.n123 B.n120 10.6151
R1332 B.n124 B.n123 10.6151
R1333 B.n127 B.n124 10.6151
R1334 B.n128 B.n127 10.6151
R1335 B.n131 B.n128 10.6151
R1336 B.n132 B.n131 10.6151
R1337 B.n135 B.n132 10.6151
R1338 B.n136 B.n135 10.6151
R1339 B.n139 B.n136 10.6151
R1340 B.n140 B.n139 10.6151
R1341 B.n143 B.n140 10.6151
R1342 B.n144 B.n143 10.6151
R1343 B.n147 B.n144 10.6151
R1344 B.n148 B.n147 10.6151
R1345 B.n151 B.n148 10.6151
R1346 B.n152 B.n151 10.6151
R1347 B.n155 B.n152 10.6151
R1348 B.n156 B.n155 10.6151
R1349 B.n159 B.n156 10.6151
R1350 B.n160 B.n159 10.6151
R1351 B.n163 B.n160 10.6151
R1352 B.n164 B.n163 10.6151
R1353 B.n167 B.n164 10.6151
R1354 B.n168 B.n167 10.6151
R1355 B.n171 B.n168 10.6151
R1356 B.n172 B.n171 10.6151
R1357 B.n175 B.n172 10.6151
R1358 B.n176 B.n175 10.6151
R1359 B.n179 B.n176 10.6151
R1360 B.n180 B.n179 10.6151
R1361 B.n183 B.n180 10.6151
R1362 B.n184 B.n183 10.6151
R1363 B.n187 B.n184 10.6151
R1364 B.n188 B.n187 10.6151
R1365 B.n191 B.n188 10.6151
R1366 B.n192 B.n191 10.6151
R1367 B.n195 B.n192 10.6151
R1368 B.n196 B.n195 10.6151
R1369 B.n199 B.n196 10.6151
R1370 B.n200 B.n199 10.6151
R1371 B.n203 B.n200 10.6151
R1372 B.n204 B.n203 10.6151
R1373 B.n207 B.n204 10.6151
R1374 B.n208 B.n207 10.6151
R1375 B.n211 B.n208 10.6151
R1376 B.n212 B.n211 10.6151
R1377 B.n215 B.n212 10.6151
R1378 B.n216 B.n215 10.6151
R1379 B.n219 B.n216 10.6151
R1380 B.n220 B.n219 10.6151
R1381 B.n223 B.n220 10.6151
R1382 B.n224 B.n223 10.6151
R1383 B.n227 B.n224 10.6151
R1384 B.n228 B.n227 10.6151
R1385 B.n231 B.n228 10.6151
R1386 B.n232 B.n231 10.6151
R1387 B.n236 B.n235 10.6151
R1388 B.n239 B.n236 10.6151
R1389 B.n240 B.n239 10.6151
R1390 B.n243 B.n240 10.6151
R1391 B.n244 B.n243 10.6151
R1392 B.n247 B.n244 10.6151
R1393 B.n248 B.n247 10.6151
R1394 B.n251 B.n248 10.6151
R1395 B.n252 B.n251 10.6151
R1396 B.n256 B.n255 10.6151
R1397 B.n259 B.n256 10.6151
R1398 B.n260 B.n259 10.6151
R1399 B.n263 B.n260 10.6151
R1400 B.n264 B.n263 10.6151
R1401 B.n267 B.n264 10.6151
R1402 B.n268 B.n267 10.6151
R1403 B.n271 B.n268 10.6151
R1404 B.n272 B.n271 10.6151
R1405 B.n275 B.n272 10.6151
R1406 B.n276 B.n275 10.6151
R1407 B.n279 B.n276 10.6151
R1408 B.n280 B.n279 10.6151
R1409 B.n283 B.n280 10.6151
R1410 B.n284 B.n283 10.6151
R1411 B.n287 B.n284 10.6151
R1412 B.n288 B.n287 10.6151
R1413 B.n291 B.n288 10.6151
R1414 B.n292 B.n291 10.6151
R1415 B.n295 B.n292 10.6151
R1416 B.n296 B.n295 10.6151
R1417 B.n299 B.n296 10.6151
R1418 B.n300 B.n299 10.6151
R1419 B.n303 B.n300 10.6151
R1420 B.n304 B.n303 10.6151
R1421 B.n307 B.n304 10.6151
R1422 B.n308 B.n307 10.6151
R1423 B.n311 B.n308 10.6151
R1424 B.n312 B.n311 10.6151
R1425 B.n315 B.n312 10.6151
R1426 B.n316 B.n315 10.6151
R1427 B.n319 B.n316 10.6151
R1428 B.n320 B.n319 10.6151
R1429 B.n323 B.n320 10.6151
R1430 B.n324 B.n323 10.6151
R1431 B.n327 B.n324 10.6151
R1432 B.n328 B.n327 10.6151
R1433 B.n331 B.n328 10.6151
R1434 B.n332 B.n331 10.6151
R1435 B.n335 B.n332 10.6151
R1436 B.n336 B.n335 10.6151
R1437 B.n339 B.n336 10.6151
R1438 B.n340 B.n339 10.6151
R1439 B.n343 B.n340 10.6151
R1440 B.n344 B.n343 10.6151
R1441 B.n347 B.n344 10.6151
R1442 B.n348 B.n347 10.6151
R1443 B.n351 B.n348 10.6151
R1444 B.n352 B.n351 10.6151
R1445 B.n355 B.n352 10.6151
R1446 B.n356 B.n355 10.6151
R1447 B.n359 B.n356 10.6151
R1448 B.n360 B.n359 10.6151
R1449 B.n363 B.n360 10.6151
R1450 B.n364 B.n363 10.6151
R1451 B.n367 B.n364 10.6151
R1452 B.n369 B.n367 10.6151
R1453 B.n370 B.n369 10.6151
R1454 B.n833 B.n370 10.6151
R1455 B.n619 B.n618 9.36635
R1456 B.n597 B.n596 9.36635
R1457 B.n232 B.n113 9.36635
R1458 B.n255 B.n110 9.36635
R1459 B.n882 B.n0 8.11757
R1460 B.n882 B.n1 8.11757
R1461 B.n618 B.n617 1.24928
R1462 B.n598 B.n597 1.24928
R1463 B.n235 B.n113 1.24928
R1464 B.n252 B.n110 1.24928
R1465 VN VN.t1 333.582
R1466 VN VN.t0 285.889
R1467 VTAIL.n402 VTAIL.n306 289.615
R1468 VTAIL.n96 VTAIL.n0 289.615
R1469 VTAIL.n300 VTAIL.n204 289.615
R1470 VTAIL.n198 VTAIL.n102 289.615
R1471 VTAIL.n338 VTAIL.n337 185
R1472 VTAIL.n343 VTAIL.n342 185
R1473 VTAIL.n345 VTAIL.n344 185
R1474 VTAIL.n334 VTAIL.n333 185
R1475 VTAIL.n351 VTAIL.n350 185
R1476 VTAIL.n353 VTAIL.n352 185
R1477 VTAIL.n330 VTAIL.n329 185
R1478 VTAIL.n359 VTAIL.n358 185
R1479 VTAIL.n361 VTAIL.n360 185
R1480 VTAIL.n326 VTAIL.n325 185
R1481 VTAIL.n367 VTAIL.n366 185
R1482 VTAIL.n369 VTAIL.n368 185
R1483 VTAIL.n322 VTAIL.n321 185
R1484 VTAIL.n375 VTAIL.n374 185
R1485 VTAIL.n377 VTAIL.n376 185
R1486 VTAIL.n318 VTAIL.n317 185
R1487 VTAIL.n384 VTAIL.n383 185
R1488 VTAIL.n385 VTAIL.n316 185
R1489 VTAIL.n387 VTAIL.n386 185
R1490 VTAIL.n314 VTAIL.n313 185
R1491 VTAIL.n393 VTAIL.n392 185
R1492 VTAIL.n395 VTAIL.n394 185
R1493 VTAIL.n310 VTAIL.n309 185
R1494 VTAIL.n401 VTAIL.n400 185
R1495 VTAIL.n403 VTAIL.n402 185
R1496 VTAIL.n32 VTAIL.n31 185
R1497 VTAIL.n37 VTAIL.n36 185
R1498 VTAIL.n39 VTAIL.n38 185
R1499 VTAIL.n28 VTAIL.n27 185
R1500 VTAIL.n45 VTAIL.n44 185
R1501 VTAIL.n47 VTAIL.n46 185
R1502 VTAIL.n24 VTAIL.n23 185
R1503 VTAIL.n53 VTAIL.n52 185
R1504 VTAIL.n55 VTAIL.n54 185
R1505 VTAIL.n20 VTAIL.n19 185
R1506 VTAIL.n61 VTAIL.n60 185
R1507 VTAIL.n63 VTAIL.n62 185
R1508 VTAIL.n16 VTAIL.n15 185
R1509 VTAIL.n69 VTAIL.n68 185
R1510 VTAIL.n71 VTAIL.n70 185
R1511 VTAIL.n12 VTAIL.n11 185
R1512 VTAIL.n78 VTAIL.n77 185
R1513 VTAIL.n79 VTAIL.n10 185
R1514 VTAIL.n81 VTAIL.n80 185
R1515 VTAIL.n8 VTAIL.n7 185
R1516 VTAIL.n87 VTAIL.n86 185
R1517 VTAIL.n89 VTAIL.n88 185
R1518 VTAIL.n4 VTAIL.n3 185
R1519 VTAIL.n95 VTAIL.n94 185
R1520 VTAIL.n97 VTAIL.n96 185
R1521 VTAIL.n301 VTAIL.n300 185
R1522 VTAIL.n299 VTAIL.n298 185
R1523 VTAIL.n208 VTAIL.n207 185
R1524 VTAIL.n293 VTAIL.n292 185
R1525 VTAIL.n291 VTAIL.n290 185
R1526 VTAIL.n212 VTAIL.n211 185
R1527 VTAIL.n285 VTAIL.n284 185
R1528 VTAIL.n283 VTAIL.n214 185
R1529 VTAIL.n282 VTAIL.n281 185
R1530 VTAIL.n217 VTAIL.n215 185
R1531 VTAIL.n276 VTAIL.n275 185
R1532 VTAIL.n274 VTAIL.n273 185
R1533 VTAIL.n221 VTAIL.n220 185
R1534 VTAIL.n268 VTAIL.n267 185
R1535 VTAIL.n266 VTAIL.n265 185
R1536 VTAIL.n225 VTAIL.n224 185
R1537 VTAIL.n260 VTAIL.n259 185
R1538 VTAIL.n258 VTAIL.n257 185
R1539 VTAIL.n229 VTAIL.n228 185
R1540 VTAIL.n252 VTAIL.n251 185
R1541 VTAIL.n250 VTAIL.n249 185
R1542 VTAIL.n233 VTAIL.n232 185
R1543 VTAIL.n244 VTAIL.n243 185
R1544 VTAIL.n242 VTAIL.n241 185
R1545 VTAIL.n237 VTAIL.n236 185
R1546 VTAIL.n199 VTAIL.n198 185
R1547 VTAIL.n197 VTAIL.n196 185
R1548 VTAIL.n106 VTAIL.n105 185
R1549 VTAIL.n191 VTAIL.n190 185
R1550 VTAIL.n189 VTAIL.n188 185
R1551 VTAIL.n110 VTAIL.n109 185
R1552 VTAIL.n183 VTAIL.n182 185
R1553 VTAIL.n181 VTAIL.n112 185
R1554 VTAIL.n180 VTAIL.n179 185
R1555 VTAIL.n115 VTAIL.n113 185
R1556 VTAIL.n174 VTAIL.n173 185
R1557 VTAIL.n172 VTAIL.n171 185
R1558 VTAIL.n119 VTAIL.n118 185
R1559 VTAIL.n166 VTAIL.n165 185
R1560 VTAIL.n164 VTAIL.n163 185
R1561 VTAIL.n123 VTAIL.n122 185
R1562 VTAIL.n158 VTAIL.n157 185
R1563 VTAIL.n156 VTAIL.n155 185
R1564 VTAIL.n127 VTAIL.n126 185
R1565 VTAIL.n150 VTAIL.n149 185
R1566 VTAIL.n148 VTAIL.n147 185
R1567 VTAIL.n131 VTAIL.n130 185
R1568 VTAIL.n142 VTAIL.n141 185
R1569 VTAIL.n140 VTAIL.n139 185
R1570 VTAIL.n135 VTAIL.n134 185
R1571 VTAIL.n339 VTAIL.t3 147.659
R1572 VTAIL.n33 VTAIL.t0 147.659
R1573 VTAIL.n238 VTAIL.t1 147.659
R1574 VTAIL.n136 VTAIL.t2 147.659
R1575 VTAIL.n343 VTAIL.n337 104.615
R1576 VTAIL.n344 VTAIL.n343 104.615
R1577 VTAIL.n344 VTAIL.n333 104.615
R1578 VTAIL.n351 VTAIL.n333 104.615
R1579 VTAIL.n352 VTAIL.n351 104.615
R1580 VTAIL.n352 VTAIL.n329 104.615
R1581 VTAIL.n359 VTAIL.n329 104.615
R1582 VTAIL.n360 VTAIL.n359 104.615
R1583 VTAIL.n360 VTAIL.n325 104.615
R1584 VTAIL.n367 VTAIL.n325 104.615
R1585 VTAIL.n368 VTAIL.n367 104.615
R1586 VTAIL.n368 VTAIL.n321 104.615
R1587 VTAIL.n375 VTAIL.n321 104.615
R1588 VTAIL.n376 VTAIL.n375 104.615
R1589 VTAIL.n376 VTAIL.n317 104.615
R1590 VTAIL.n384 VTAIL.n317 104.615
R1591 VTAIL.n385 VTAIL.n384 104.615
R1592 VTAIL.n386 VTAIL.n385 104.615
R1593 VTAIL.n386 VTAIL.n313 104.615
R1594 VTAIL.n393 VTAIL.n313 104.615
R1595 VTAIL.n394 VTAIL.n393 104.615
R1596 VTAIL.n394 VTAIL.n309 104.615
R1597 VTAIL.n401 VTAIL.n309 104.615
R1598 VTAIL.n402 VTAIL.n401 104.615
R1599 VTAIL.n37 VTAIL.n31 104.615
R1600 VTAIL.n38 VTAIL.n37 104.615
R1601 VTAIL.n38 VTAIL.n27 104.615
R1602 VTAIL.n45 VTAIL.n27 104.615
R1603 VTAIL.n46 VTAIL.n45 104.615
R1604 VTAIL.n46 VTAIL.n23 104.615
R1605 VTAIL.n53 VTAIL.n23 104.615
R1606 VTAIL.n54 VTAIL.n53 104.615
R1607 VTAIL.n54 VTAIL.n19 104.615
R1608 VTAIL.n61 VTAIL.n19 104.615
R1609 VTAIL.n62 VTAIL.n61 104.615
R1610 VTAIL.n62 VTAIL.n15 104.615
R1611 VTAIL.n69 VTAIL.n15 104.615
R1612 VTAIL.n70 VTAIL.n69 104.615
R1613 VTAIL.n70 VTAIL.n11 104.615
R1614 VTAIL.n78 VTAIL.n11 104.615
R1615 VTAIL.n79 VTAIL.n78 104.615
R1616 VTAIL.n80 VTAIL.n79 104.615
R1617 VTAIL.n80 VTAIL.n7 104.615
R1618 VTAIL.n87 VTAIL.n7 104.615
R1619 VTAIL.n88 VTAIL.n87 104.615
R1620 VTAIL.n88 VTAIL.n3 104.615
R1621 VTAIL.n95 VTAIL.n3 104.615
R1622 VTAIL.n96 VTAIL.n95 104.615
R1623 VTAIL.n300 VTAIL.n299 104.615
R1624 VTAIL.n299 VTAIL.n207 104.615
R1625 VTAIL.n292 VTAIL.n207 104.615
R1626 VTAIL.n292 VTAIL.n291 104.615
R1627 VTAIL.n291 VTAIL.n211 104.615
R1628 VTAIL.n284 VTAIL.n211 104.615
R1629 VTAIL.n284 VTAIL.n283 104.615
R1630 VTAIL.n283 VTAIL.n282 104.615
R1631 VTAIL.n282 VTAIL.n215 104.615
R1632 VTAIL.n275 VTAIL.n215 104.615
R1633 VTAIL.n275 VTAIL.n274 104.615
R1634 VTAIL.n274 VTAIL.n220 104.615
R1635 VTAIL.n267 VTAIL.n220 104.615
R1636 VTAIL.n267 VTAIL.n266 104.615
R1637 VTAIL.n266 VTAIL.n224 104.615
R1638 VTAIL.n259 VTAIL.n224 104.615
R1639 VTAIL.n259 VTAIL.n258 104.615
R1640 VTAIL.n258 VTAIL.n228 104.615
R1641 VTAIL.n251 VTAIL.n228 104.615
R1642 VTAIL.n251 VTAIL.n250 104.615
R1643 VTAIL.n250 VTAIL.n232 104.615
R1644 VTAIL.n243 VTAIL.n232 104.615
R1645 VTAIL.n243 VTAIL.n242 104.615
R1646 VTAIL.n242 VTAIL.n236 104.615
R1647 VTAIL.n198 VTAIL.n197 104.615
R1648 VTAIL.n197 VTAIL.n105 104.615
R1649 VTAIL.n190 VTAIL.n105 104.615
R1650 VTAIL.n190 VTAIL.n189 104.615
R1651 VTAIL.n189 VTAIL.n109 104.615
R1652 VTAIL.n182 VTAIL.n109 104.615
R1653 VTAIL.n182 VTAIL.n181 104.615
R1654 VTAIL.n181 VTAIL.n180 104.615
R1655 VTAIL.n180 VTAIL.n113 104.615
R1656 VTAIL.n173 VTAIL.n113 104.615
R1657 VTAIL.n173 VTAIL.n172 104.615
R1658 VTAIL.n172 VTAIL.n118 104.615
R1659 VTAIL.n165 VTAIL.n118 104.615
R1660 VTAIL.n165 VTAIL.n164 104.615
R1661 VTAIL.n164 VTAIL.n122 104.615
R1662 VTAIL.n157 VTAIL.n122 104.615
R1663 VTAIL.n157 VTAIL.n156 104.615
R1664 VTAIL.n156 VTAIL.n126 104.615
R1665 VTAIL.n149 VTAIL.n126 104.615
R1666 VTAIL.n149 VTAIL.n148 104.615
R1667 VTAIL.n148 VTAIL.n130 104.615
R1668 VTAIL.n141 VTAIL.n130 104.615
R1669 VTAIL.n141 VTAIL.n140 104.615
R1670 VTAIL.n140 VTAIL.n134 104.615
R1671 VTAIL.t3 VTAIL.n337 52.3082
R1672 VTAIL.t0 VTAIL.n31 52.3082
R1673 VTAIL.t1 VTAIL.n236 52.3082
R1674 VTAIL.t2 VTAIL.n134 52.3082
R1675 VTAIL.n407 VTAIL.n406 34.3187
R1676 VTAIL.n101 VTAIL.n100 34.3187
R1677 VTAIL.n305 VTAIL.n304 34.3187
R1678 VTAIL.n203 VTAIL.n202 34.3187
R1679 VTAIL.n203 VTAIL.n101 32.1169
R1680 VTAIL.n407 VTAIL.n305 30.1514
R1681 VTAIL.n339 VTAIL.n338 15.6677
R1682 VTAIL.n33 VTAIL.n32 15.6677
R1683 VTAIL.n238 VTAIL.n237 15.6677
R1684 VTAIL.n136 VTAIL.n135 15.6677
R1685 VTAIL.n387 VTAIL.n316 13.1884
R1686 VTAIL.n81 VTAIL.n10 13.1884
R1687 VTAIL.n285 VTAIL.n214 13.1884
R1688 VTAIL.n183 VTAIL.n112 13.1884
R1689 VTAIL.n342 VTAIL.n341 12.8005
R1690 VTAIL.n383 VTAIL.n382 12.8005
R1691 VTAIL.n388 VTAIL.n314 12.8005
R1692 VTAIL.n36 VTAIL.n35 12.8005
R1693 VTAIL.n77 VTAIL.n76 12.8005
R1694 VTAIL.n82 VTAIL.n8 12.8005
R1695 VTAIL.n286 VTAIL.n212 12.8005
R1696 VTAIL.n281 VTAIL.n216 12.8005
R1697 VTAIL.n241 VTAIL.n240 12.8005
R1698 VTAIL.n184 VTAIL.n110 12.8005
R1699 VTAIL.n179 VTAIL.n114 12.8005
R1700 VTAIL.n139 VTAIL.n138 12.8005
R1701 VTAIL.n345 VTAIL.n336 12.0247
R1702 VTAIL.n381 VTAIL.n318 12.0247
R1703 VTAIL.n392 VTAIL.n391 12.0247
R1704 VTAIL.n39 VTAIL.n30 12.0247
R1705 VTAIL.n75 VTAIL.n12 12.0247
R1706 VTAIL.n86 VTAIL.n85 12.0247
R1707 VTAIL.n290 VTAIL.n289 12.0247
R1708 VTAIL.n280 VTAIL.n217 12.0247
R1709 VTAIL.n244 VTAIL.n235 12.0247
R1710 VTAIL.n188 VTAIL.n187 12.0247
R1711 VTAIL.n178 VTAIL.n115 12.0247
R1712 VTAIL.n142 VTAIL.n133 12.0247
R1713 VTAIL.n346 VTAIL.n334 11.249
R1714 VTAIL.n378 VTAIL.n377 11.249
R1715 VTAIL.n395 VTAIL.n312 11.249
R1716 VTAIL.n40 VTAIL.n28 11.249
R1717 VTAIL.n72 VTAIL.n71 11.249
R1718 VTAIL.n89 VTAIL.n6 11.249
R1719 VTAIL.n293 VTAIL.n210 11.249
R1720 VTAIL.n277 VTAIL.n276 11.249
R1721 VTAIL.n245 VTAIL.n233 11.249
R1722 VTAIL.n191 VTAIL.n108 11.249
R1723 VTAIL.n175 VTAIL.n174 11.249
R1724 VTAIL.n143 VTAIL.n131 11.249
R1725 VTAIL.n350 VTAIL.n349 10.4732
R1726 VTAIL.n374 VTAIL.n320 10.4732
R1727 VTAIL.n396 VTAIL.n310 10.4732
R1728 VTAIL.n44 VTAIL.n43 10.4732
R1729 VTAIL.n68 VTAIL.n14 10.4732
R1730 VTAIL.n90 VTAIL.n4 10.4732
R1731 VTAIL.n294 VTAIL.n208 10.4732
R1732 VTAIL.n273 VTAIL.n219 10.4732
R1733 VTAIL.n249 VTAIL.n248 10.4732
R1734 VTAIL.n192 VTAIL.n106 10.4732
R1735 VTAIL.n171 VTAIL.n117 10.4732
R1736 VTAIL.n147 VTAIL.n146 10.4732
R1737 VTAIL.n353 VTAIL.n332 9.69747
R1738 VTAIL.n373 VTAIL.n322 9.69747
R1739 VTAIL.n400 VTAIL.n399 9.69747
R1740 VTAIL.n47 VTAIL.n26 9.69747
R1741 VTAIL.n67 VTAIL.n16 9.69747
R1742 VTAIL.n94 VTAIL.n93 9.69747
R1743 VTAIL.n298 VTAIL.n297 9.69747
R1744 VTAIL.n272 VTAIL.n221 9.69747
R1745 VTAIL.n252 VTAIL.n231 9.69747
R1746 VTAIL.n196 VTAIL.n195 9.69747
R1747 VTAIL.n170 VTAIL.n119 9.69747
R1748 VTAIL.n150 VTAIL.n129 9.69747
R1749 VTAIL.n406 VTAIL.n405 9.45567
R1750 VTAIL.n100 VTAIL.n99 9.45567
R1751 VTAIL.n304 VTAIL.n303 9.45567
R1752 VTAIL.n202 VTAIL.n201 9.45567
R1753 VTAIL.n405 VTAIL.n404 9.3005
R1754 VTAIL.n308 VTAIL.n307 9.3005
R1755 VTAIL.n399 VTAIL.n398 9.3005
R1756 VTAIL.n397 VTAIL.n396 9.3005
R1757 VTAIL.n312 VTAIL.n311 9.3005
R1758 VTAIL.n391 VTAIL.n390 9.3005
R1759 VTAIL.n389 VTAIL.n388 9.3005
R1760 VTAIL.n328 VTAIL.n327 9.3005
R1761 VTAIL.n357 VTAIL.n356 9.3005
R1762 VTAIL.n355 VTAIL.n354 9.3005
R1763 VTAIL.n332 VTAIL.n331 9.3005
R1764 VTAIL.n349 VTAIL.n348 9.3005
R1765 VTAIL.n347 VTAIL.n346 9.3005
R1766 VTAIL.n336 VTAIL.n335 9.3005
R1767 VTAIL.n341 VTAIL.n340 9.3005
R1768 VTAIL.n363 VTAIL.n362 9.3005
R1769 VTAIL.n365 VTAIL.n364 9.3005
R1770 VTAIL.n324 VTAIL.n323 9.3005
R1771 VTAIL.n371 VTAIL.n370 9.3005
R1772 VTAIL.n373 VTAIL.n372 9.3005
R1773 VTAIL.n320 VTAIL.n319 9.3005
R1774 VTAIL.n379 VTAIL.n378 9.3005
R1775 VTAIL.n381 VTAIL.n380 9.3005
R1776 VTAIL.n382 VTAIL.n315 9.3005
R1777 VTAIL.n99 VTAIL.n98 9.3005
R1778 VTAIL.n2 VTAIL.n1 9.3005
R1779 VTAIL.n93 VTAIL.n92 9.3005
R1780 VTAIL.n91 VTAIL.n90 9.3005
R1781 VTAIL.n6 VTAIL.n5 9.3005
R1782 VTAIL.n85 VTAIL.n84 9.3005
R1783 VTAIL.n83 VTAIL.n82 9.3005
R1784 VTAIL.n22 VTAIL.n21 9.3005
R1785 VTAIL.n51 VTAIL.n50 9.3005
R1786 VTAIL.n49 VTAIL.n48 9.3005
R1787 VTAIL.n26 VTAIL.n25 9.3005
R1788 VTAIL.n43 VTAIL.n42 9.3005
R1789 VTAIL.n41 VTAIL.n40 9.3005
R1790 VTAIL.n30 VTAIL.n29 9.3005
R1791 VTAIL.n35 VTAIL.n34 9.3005
R1792 VTAIL.n57 VTAIL.n56 9.3005
R1793 VTAIL.n59 VTAIL.n58 9.3005
R1794 VTAIL.n18 VTAIL.n17 9.3005
R1795 VTAIL.n65 VTAIL.n64 9.3005
R1796 VTAIL.n67 VTAIL.n66 9.3005
R1797 VTAIL.n14 VTAIL.n13 9.3005
R1798 VTAIL.n73 VTAIL.n72 9.3005
R1799 VTAIL.n75 VTAIL.n74 9.3005
R1800 VTAIL.n76 VTAIL.n9 9.3005
R1801 VTAIL.n264 VTAIL.n263 9.3005
R1802 VTAIL.n223 VTAIL.n222 9.3005
R1803 VTAIL.n270 VTAIL.n269 9.3005
R1804 VTAIL.n272 VTAIL.n271 9.3005
R1805 VTAIL.n219 VTAIL.n218 9.3005
R1806 VTAIL.n278 VTAIL.n277 9.3005
R1807 VTAIL.n280 VTAIL.n279 9.3005
R1808 VTAIL.n216 VTAIL.n213 9.3005
R1809 VTAIL.n303 VTAIL.n302 9.3005
R1810 VTAIL.n206 VTAIL.n205 9.3005
R1811 VTAIL.n297 VTAIL.n296 9.3005
R1812 VTAIL.n295 VTAIL.n294 9.3005
R1813 VTAIL.n210 VTAIL.n209 9.3005
R1814 VTAIL.n289 VTAIL.n288 9.3005
R1815 VTAIL.n287 VTAIL.n286 9.3005
R1816 VTAIL.n262 VTAIL.n261 9.3005
R1817 VTAIL.n227 VTAIL.n226 9.3005
R1818 VTAIL.n256 VTAIL.n255 9.3005
R1819 VTAIL.n254 VTAIL.n253 9.3005
R1820 VTAIL.n231 VTAIL.n230 9.3005
R1821 VTAIL.n248 VTAIL.n247 9.3005
R1822 VTAIL.n246 VTAIL.n245 9.3005
R1823 VTAIL.n235 VTAIL.n234 9.3005
R1824 VTAIL.n240 VTAIL.n239 9.3005
R1825 VTAIL.n162 VTAIL.n161 9.3005
R1826 VTAIL.n121 VTAIL.n120 9.3005
R1827 VTAIL.n168 VTAIL.n167 9.3005
R1828 VTAIL.n170 VTAIL.n169 9.3005
R1829 VTAIL.n117 VTAIL.n116 9.3005
R1830 VTAIL.n176 VTAIL.n175 9.3005
R1831 VTAIL.n178 VTAIL.n177 9.3005
R1832 VTAIL.n114 VTAIL.n111 9.3005
R1833 VTAIL.n201 VTAIL.n200 9.3005
R1834 VTAIL.n104 VTAIL.n103 9.3005
R1835 VTAIL.n195 VTAIL.n194 9.3005
R1836 VTAIL.n193 VTAIL.n192 9.3005
R1837 VTAIL.n108 VTAIL.n107 9.3005
R1838 VTAIL.n187 VTAIL.n186 9.3005
R1839 VTAIL.n185 VTAIL.n184 9.3005
R1840 VTAIL.n160 VTAIL.n159 9.3005
R1841 VTAIL.n125 VTAIL.n124 9.3005
R1842 VTAIL.n154 VTAIL.n153 9.3005
R1843 VTAIL.n152 VTAIL.n151 9.3005
R1844 VTAIL.n129 VTAIL.n128 9.3005
R1845 VTAIL.n146 VTAIL.n145 9.3005
R1846 VTAIL.n144 VTAIL.n143 9.3005
R1847 VTAIL.n133 VTAIL.n132 9.3005
R1848 VTAIL.n138 VTAIL.n137 9.3005
R1849 VTAIL.n354 VTAIL.n330 8.92171
R1850 VTAIL.n370 VTAIL.n369 8.92171
R1851 VTAIL.n403 VTAIL.n308 8.92171
R1852 VTAIL.n48 VTAIL.n24 8.92171
R1853 VTAIL.n64 VTAIL.n63 8.92171
R1854 VTAIL.n97 VTAIL.n2 8.92171
R1855 VTAIL.n301 VTAIL.n206 8.92171
R1856 VTAIL.n269 VTAIL.n268 8.92171
R1857 VTAIL.n253 VTAIL.n229 8.92171
R1858 VTAIL.n199 VTAIL.n104 8.92171
R1859 VTAIL.n167 VTAIL.n166 8.92171
R1860 VTAIL.n151 VTAIL.n127 8.92171
R1861 VTAIL.n358 VTAIL.n357 8.14595
R1862 VTAIL.n366 VTAIL.n324 8.14595
R1863 VTAIL.n404 VTAIL.n306 8.14595
R1864 VTAIL.n52 VTAIL.n51 8.14595
R1865 VTAIL.n60 VTAIL.n18 8.14595
R1866 VTAIL.n98 VTAIL.n0 8.14595
R1867 VTAIL.n302 VTAIL.n204 8.14595
R1868 VTAIL.n265 VTAIL.n223 8.14595
R1869 VTAIL.n257 VTAIL.n256 8.14595
R1870 VTAIL.n200 VTAIL.n102 8.14595
R1871 VTAIL.n163 VTAIL.n121 8.14595
R1872 VTAIL.n155 VTAIL.n154 8.14595
R1873 VTAIL.n361 VTAIL.n328 7.3702
R1874 VTAIL.n365 VTAIL.n326 7.3702
R1875 VTAIL.n55 VTAIL.n22 7.3702
R1876 VTAIL.n59 VTAIL.n20 7.3702
R1877 VTAIL.n264 VTAIL.n225 7.3702
R1878 VTAIL.n260 VTAIL.n227 7.3702
R1879 VTAIL.n162 VTAIL.n123 7.3702
R1880 VTAIL.n158 VTAIL.n125 7.3702
R1881 VTAIL.n362 VTAIL.n361 6.59444
R1882 VTAIL.n362 VTAIL.n326 6.59444
R1883 VTAIL.n56 VTAIL.n55 6.59444
R1884 VTAIL.n56 VTAIL.n20 6.59444
R1885 VTAIL.n261 VTAIL.n225 6.59444
R1886 VTAIL.n261 VTAIL.n260 6.59444
R1887 VTAIL.n159 VTAIL.n123 6.59444
R1888 VTAIL.n159 VTAIL.n158 6.59444
R1889 VTAIL.n358 VTAIL.n328 5.81868
R1890 VTAIL.n366 VTAIL.n365 5.81868
R1891 VTAIL.n406 VTAIL.n306 5.81868
R1892 VTAIL.n52 VTAIL.n22 5.81868
R1893 VTAIL.n60 VTAIL.n59 5.81868
R1894 VTAIL.n100 VTAIL.n0 5.81868
R1895 VTAIL.n304 VTAIL.n204 5.81868
R1896 VTAIL.n265 VTAIL.n264 5.81868
R1897 VTAIL.n257 VTAIL.n227 5.81868
R1898 VTAIL.n202 VTAIL.n102 5.81868
R1899 VTAIL.n163 VTAIL.n162 5.81868
R1900 VTAIL.n155 VTAIL.n125 5.81868
R1901 VTAIL.n357 VTAIL.n330 5.04292
R1902 VTAIL.n369 VTAIL.n324 5.04292
R1903 VTAIL.n404 VTAIL.n403 5.04292
R1904 VTAIL.n51 VTAIL.n24 5.04292
R1905 VTAIL.n63 VTAIL.n18 5.04292
R1906 VTAIL.n98 VTAIL.n97 5.04292
R1907 VTAIL.n302 VTAIL.n301 5.04292
R1908 VTAIL.n268 VTAIL.n223 5.04292
R1909 VTAIL.n256 VTAIL.n229 5.04292
R1910 VTAIL.n200 VTAIL.n199 5.04292
R1911 VTAIL.n166 VTAIL.n121 5.04292
R1912 VTAIL.n154 VTAIL.n127 5.04292
R1913 VTAIL.n340 VTAIL.n339 4.38563
R1914 VTAIL.n34 VTAIL.n33 4.38563
R1915 VTAIL.n239 VTAIL.n238 4.38563
R1916 VTAIL.n137 VTAIL.n136 4.38563
R1917 VTAIL.n354 VTAIL.n353 4.26717
R1918 VTAIL.n370 VTAIL.n322 4.26717
R1919 VTAIL.n400 VTAIL.n308 4.26717
R1920 VTAIL.n48 VTAIL.n47 4.26717
R1921 VTAIL.n64 VTAIL.n16 4.26717
R1922 VTAIL.n94 VTAIL.n2 4.26717
R1923 VTAIL.n298 VTAIL.n206 4.26717
R1924 VTAIL.n269 VTAIL.n221 4.26717
R1925 VTAIL.n253 VTAIL.n252 4.26717
R1926 VTAIL.n196 VTAIL.n104 4.26717
R1927 VTAIL.n167 VTAIL.n119 4.26717
R1928 VTAIL.n151 VTAIL.n150 4.26717
R1929 VTAIL.n350 VTAIL.n332 3.49141
R1930 VTAIL.n374 VTAIL.n373 3.49141
R1931 VTAIL.n399 VTAIL.n310 3.49141
R1932 VTAIL.n44 VTAIL.n26 3.49141
R1933 VTAIL.n68 VTAIL.n67 3.49141
R1934 VTAIL.n93 VTAIL.n4 3.49141
R1935 VTAIL.n297 VTAIL.n208 3.49141
R1936 VTAIL.n273 VTAIL.n272 3.49141
R1937 VTAIL.n249 VTAIL.n231 3.49141
R1938 VTAIL.n195 VTAIL.n106 3.49141
R1939 VTAIL.n171 VTAIL.n170 3.49141
R1940 VTAIL.n147 VTAIL.n129 3.49141
R1941 VTAIL.n349 VTAIL.n334 2.71565
R1942 VTAIL.n377 VTAIL.n320 2.71565
R1943 VTAIL.n396 VTAIL.n395 2.71565
R1944 VTAIL.n43 VTAIL.n28 2.71565
R1945 VTAIL.n71 VTAIL.n14 2.71565
R1946 VTAIL.n90 VTAIL.n89 2.71565
R1947 VTAIL.n294 VTAIL.n293 2.71565
R1948 VTAIL.n276 VTAIL.n219 2.71565
R1949 VTAIL.n248 VTAIL.n233 2.71565
R1950 VTAIL.n192 VTAIL.n191 2.71565
R1951 VTAIL.n174 VTAIL.n117 2.71565
R1952 VTAIL.n146 VTAIL.n131 2.71565
R1953 VTAIL.n346 VTAIL.n345 1.93989
R1954 VTAIL.n378 VTAIL.n318 1.93989
R1955 VTAIL.n392 VTAIL.n312 1.93989
R1956 VTAIL.n40 VTAIL.n39 1.93989
R1957 VTAIL.n72 VTAIL.n12 1.93989
R1958 VTAIL.n86 VTAIL.n6 1.93989
R1959 VTAIL.n290 VTAIL.n210 1.93989
R1960 VTAIL.n277 VTAIL.n217 1.93989
R1961 VTAIL.n245 VTAIL.n244 1.93989
R1962 VTAIL.n188 VTAIL.n108 1.93989
R1963 VTAIL.n175 VTAIL.n115 1.93989
R1964 VTAIL.n143 VTAIL.n142 1.93989
R1965 VTAIL.n305 VTAIL.n203 1.45309
R1966 VTAIL.n342 VTAIL.n336 1.16414
R1967 VTAIL.n383 VTAIL.n381 1.16414
R1968 VTAIL.n391 VTAIL.n314 1.16414
R1969 VTAIL.n36 VTAIL.n30 1.16414
R1970 VTAIL.n77 VTAIL.n75 1.16414
R1971 VTAIL.n85 VTAIL.n8 1.16414
R1972 VTAIL.n289 VTAIL.n212 1.16414
R1973 VTAIL.n281 VTAIL.n280 1.16414
R1974 VTAIL.n241 VTAIL.n235 1.16414
R1975 VTAIL.n187 VTAIL.n110 1.16414
R1976 VTAIL.n179 VTAIL.n178 1.16414
R1977 VTAIL.n139 VTAIL.n133 1.16414
R1978 VTAIL VTAIL.n101 1.0199
R1979 VTAIL VTAIL.n407 0.43369
R1980 VTAIL.n341 VTAIL.n338 0.388379
R1981 VTAIL.n382 VTAIL.n316 0.388379
R1982 VTAIL.n388 VTAIL.n387 0.388379
R1983 VTAIL.n35 VTAIL.n32 0.388379
R1984 VTAIL.n76 VTAIL.n10 0.388379
R1985 VTAIL.n82 VTAIL.n81 0.388379
R1986 VTAIL.n286 VTAIL.n285 0.388379
R1987 VTAIL.n216 VTAIL.n214 0.388379
R1988 VTAIL.n240 VTAIL.n237 0.388379
R1989 VTAIL.n184 VTAIL.n183 0.388379
R1990 VTAIL.n114 VTAIL.n112 0.388379
R1991 VTAIL.n138 VTAIL.n135 0.388379
R1992 VTAIL.n340 VTAIL.n335 0.155672
R1993 VTAIL.n347 VTAIL.n335 0.155672
R1994 VTAIL.n348 VTAIL.n347 0.155672
R1995 VTAIL.n348 VTAIL.n331 0.155672
R1996 VTAIL.n355 VTAIL.n331 0.155672
R1997 VTAIL.n356 VTAIL.n355 0.155672
R1998 VTAIL.n356 VTAIL.n327 0.155672
R1999 VTAIL.n363 VTAIL.n327 0.155672
R2000 VTAIL.n364 VTAIL.n363 0.155672
R2001 VTAIL.n364 VTAIL.n323 0.155672
R2002 VTAIL.n371 VTAIL.n323 0.155672
R2003 VTAIL.n372 VTAIL.n371 0.155672
R2004 VTAIL.n372 VTAIL.n319 0.155672
R2005 VTAIL.n379 VTAIL.n319 0.155672
R2006 VTAIL.n380 VTAIL.n379 0.155672
R2007 VTAIL.n380 VTAIL.n315 0.155672
R2008 VTAIL.n389 VTAIL.n315 0.155672
R2009 VTAIL.n390 VTAIL.n389 0.155672
R2010 VTAIL.n390 VTAIL.n311 0.155672
R2011 VTAIL.n397 VTAIL.n311 0.155672
R2012 VTAIL.n398 VTAIL.n397 0.155672
R2013 VTAIL.n398 VTAIL.n307 0.155672
R2014 VTAIL.n405 VTAIL.n307 0.155672
R2015 VTAIL.n34 VTAIL.n29 0.155672
R2016 VTAIL.n41 VTAIL.n29 0.155672
R2017 VTAIL.n42 VTAIL.n41 0.155672
R2018 VTAIL.n42 VTAIL.n25 0.155672
R2019 VTAIL.n49 VTAIL.n25 0.155672
R2020 VTAIL.n50 VTAIL.n49 0.155672
R2021 VTAIL.n50 VTAIL.n21 0.155672
R2022 VTAIL.n57 VTAIL.n21 0.155672
R2023 VTAIL.n58 VTAIL.n57 0.155672
R2024 VTAIL.n58 VTAIL.n17 0.155672
R2025 VTAIL.n65 VTAIL.n17 0.155672
R2026 VTAIL.n66 VTAIL.n65 0.155672
R2027 VTAIL.n66 VTAIL.n13 0.155672
R2028 VTAIL.n73 VTAIL.n13 0.155672
R2029 VTAIL.n74 VTAIL.n73 0.155672
R2030 VTAIL.n74 VTAIL.n9 0.155672
R2031 VTAIL.n83 VTAIL.n9 0.155672
R2032 VTAIL.n84 VTAIL.n83 0.155672
R2033 VTAIL.n84 VTAIL.n5 0.155672
R2034 VTAIL.n91 VTAIL.n5 0.155672
R2035 VTAIL.n92 VTAIL.n91 0.155672
R2036 VTAIL.n92 VTAIL.n1 0.155672
R2037 VTAIL.n99 VTAIL.n1 0.155672
R2038 VTAIL.n303 VTAIL.n205 0.155672
R2039 VTAIL.n296 VTAIL.n205 0.155672
R2040 VTAIL.n296 VTAIL.n295 0.155672
R2041 VTAIL.n295 VTAIL.n209 0.155672
R2042 VTAIL.n288 VTAIL.n209 0.155672
R2043 VTAIL.n288 VTAIL.n287 0.155672
R2044 VTAIL.n287 VTAIL.n213 0.155672
R2045 VTAIL.n279 VTAIL.n213 0.155672
R2046 VTAIL.n279 VTAIL.n278 0.155672
R2047 VTAIL.n278 VTAIL.n218 0.155672
R2048 VTAIL.n271 VTAIL.n218 0.155672
R2049 VTAIL.n271 VTAIL.n270 0.155672
R2050 VTAIL.n270 VTAIL.n222 0.155672
R2051 VTAIL.n263 VTAIL.n222 0.155672
R2052 VTAIL.n263 VTAIL.n262 0.155672
R2053 VTAIL.n262 VTAIL.n226 0.155672
R2054 VTAIL.n255 VTAIL.n226 0.155672
R2055 VTAIL.n255 VTAIL.n254 0.155672
R2056 VTAIL.n254 VTAIL.n230 0.155672
R2057 VTAIL.n247 VTAIL.n230 0.155672
R2058 VTAIL.n247 VTAIL.n246 0.155672
R2059 VTAIL.n246 VTAIL.n234 0.155672
R2060 VTAIL.n239 VTAIL.n234 0.155672
R2061 VTAIL.n201 VTAIL.n103 0.155672
R2062 VTAIL.n194 VTAIL.n103 0.155672
R2063 VTAIL.n194 VTAIL.n193 0.155672
R2064 VTAIL.n193 VTAIL.n107 0.155672
R2065 VTAIL.n186 VTAIL.n107 0.155672
R2066 VTAIL.n186 VTAIL.n185 0.155672
R2067 VTAIL.n185 VTAIL.n111 0.155672
R2068 VTAIL.n177 VTAIL.n111 0.155672
R2069 VTAIL.n177 VTAIL.n176 0.155672
R2070 VTAIL.n176 VTAIL.n116 0.155672
R2071 VTAIL.n169 VTAIL.n116 0.155672
R2072 VTAIL.n169 VTAIL.n168 0.155672
R2073 VTAIL.n168 VTAIL.n120 0.155672
R2074 VTAIL.n161 VTAIL.n120 0.155672
R2075 VTAIL.n161 VTAIL.n160 0.155672
R2076 VTAIL.n160 VTAIL.n124 0.155672
R2077 VTAIL.n153 VTAIL.n124 0.155672
R2078 VTAIL.n153 VTAIL.n152 0.155672
R2079 VTAIL.n152 VTAIL.n128 0.155672
R2080 VTAIL.n145 VTAIL.n128 0.155672
R2081 VTAIL.n145 VTAIL.n144 0.155672
R2082 VTAIL.n144 VTAIL.n132 0.155672
R2083 VTAIL.n137 VTAIL.n132 0.155672
R2084 VDD2.n197 VDD2.n101 289.615
R2085 VDD2.n96 VDD2.n0 289.615
R2086 VDD2.n198 VDD2.n197 185
R2087 VDD2.n196 VDD2.n195 185
R2088 VDD2.n105 VDD2.n104 185
R2089 VDD2.n190 VDD2.n189 185
R2090 VDD2.n188 VDD2.n187 185
R2091 VDD2.n109 VDD2.n108 185
R2092 VDD2.n182 VDD2.n181 185
R2093 VDD2.n180 VDD2.n111 185
R2094 VDD2.n179 VDD2.n178 185
R2095 VDD2.n114 VDD2.n112 185
R2096 VDD2.n173 VDD2.n172 185
R2097 VDD2.n171 VDD2.n170 185
R2098 VDD2.n118 VDD2.n117 185
R2099 VDD2.n165 VDD2.n164 185
R2100 VDD2.n163 VDD2.n162 185
R2101 VDD2.n122 VDD2.n121 185
R2102 VDD2.n157 VDD2.n156 185
R2103 VDD2.n155 VDD2.n154 185
R2104 VDD2.n126 VDD2.n125 185
R2105 VDD2.n149 VDD2.n148 185
R2106 VDD2.n147 VDD2.n146 185
R2107 VDD2.n130 VDD2.n129 185
R2108 VDD2.n141 VDD2.n140 185
R2109 VDD2.n139 VDD2.n138 185
R2110 VDD2.n134 VDD2.n133 185
R2111 VDD2.n32 VDD2.n31 185
R2112 VDD2.n37 VDD2.n36 185
R2113 VDD2.n39 VDD2.n38 185
R2114 VDD2.n28 VDD2.n27 185
R2115 VDD2.n45 VDD2.n44 185
R2116 VDD2.n47 VDD2.n46 185
R2117 VDD2.n24 VDD2.n23 185
R2118 VDD2.n53 VDD2.n52 185
R2119 VDD2.n55 VDD2.n54 185
R2120 VDD2.n20 VDD2.n19 185
R2121 VDD2.n61 VDD2.n60 185
R2122 VDD2.n63 VDD2.n62 185
R2123 VDD2.n16 VDD2.n15 185
R2124 VDD2.n69 VDD2.n68 185
R2125 VDD2.n71 VDD2.n70 185
R2126 VDD2.n12 VDD2.n11 185
R2127 VDD2.n78 VDD2.n77 185
R2128 VDD2.n79 VDD2.n10 185
R2129 VDD2.n81 VDD2.n80 185
R2130 VDD2.n8 VDD2.n7 185
R2131 VDD2.n87 VDD2.n86 185
R2132 VDD2.n89 VDD2.n88 185
R2133 VDD2.n4 VDD2.n3 185
R2134 VDD2.n95 VDD2.n94 185
R2135 VDD2.n97 VDD2.n96 185
R2136 VDD2.n135 VDD2.t0 147.659
R2137 VDD2.n33 VDD2.t1 147.659
R2138 VDD2.n197 VDD2.n196 104.615
R2139 VDD2.n196 VDD2.n104 104.615
R2140 VDD2.n189 VDD2.n104 104.615
R2141 VDD2.n189 VDD2.n188 104.615
R2142 VDD2.n188 VDD2.n108 104.615
R2143 VDD2.n181 VDD2.n108 104.615
R2144 VDD2.n181 VDD2.n180 104.615
R2145 VDD2.n180 VDD2.n179 104.615
R2146 VDD2.n179 VDD2.n112 104.615
R2147 VDD2.n172 VDD2.n112 104.615
R2148 VDD2.n172 VDD2.n171 104.615
R2149 VDD2.n171 VDD2.n117 104.615
R2150 VDD2.n164 VDD2.n117 104.615
R2151 VDD2.n164 VDD2.n163 104.615
R2152 VDD2.n163 VDD2.n121 104.615
R2153 VDD2.n156 VDD2.n121 104.615
R2154 VDD2.n156 VDD2.n155 104.615
R2155 VDD2.n155 VDD2.n125 104.615
R2156 VDD2.n148 VDD2.n125 104.615
R2157 VDD2.n148 VDD2.n147 104.615
R2158 VDD2.n147 VDD2.n129 104.615
R2159 VDD2.n140 VDD2.n129 104.615
R2160 VDD2.n140 VDD2.n139 104.615
R2161 VDD2.n139 VDD2.n133 104.615
R2162 VDD2.n37 VDD2.n31 104.615
R2163 VDD2.n38 VDD2.n37 104.615
R2164 VDD2.n38 VDD2.n27 104.615
R2165 VDD2.n45 VDD2.n27 104.615
R2166 VDD2.n46 VDD2.n45 104.615
R2167 VDD2.n46 VDD2.n23 104.615
R2168 VDD2.n53 VDD2.n23 104.615
R2169 VDD2.n54 VDD2.n53 104.615
R2170 VDD2.n54 VDD2.n19 104.615
R2171 VDD2.n61 VDD2.n19 104.615
R2172 VDD2.n62 VDD2.n61 104.615
R2173 VDD2.n62 VDD2.n15 104.615
R2174 VDD2.n69 VDD2.n15 104.615
R2175 VDD2.n70 VDD2.n69 104.615
R2176 VDD2.n70 VDD2.n11 104.615
R2177 VDD2.n78 VDD2.n11 104.615
R2178 VDD2.n79 VDD2.n78 104.615
R2179 VDD2.n80 VDD2.n79 104.615
R2180 VDD2.n80 VDD2.n7 104.615
R2181 VDD2.n87 VDD2.n7 104.615
R2182 VDD2.n88 VDD2.n87 104.615
R2183 VDD2.n88 VDD2.n3 104.615
R2184 VDD2.n95 VDD2.n3 104.615
R2185 VDD2.n96 VDD2.n95 104.615
R2186 VDD2.n202 VDD2.n100 94.4069
R2187 VDD2.t0 VDD2.n133 52.3082
R2188 VDD2.t1 VDD2.n31 52.3082
R2189 VDD2.n202 VDD2.n201 50.9975
R2190 VDD2.n135 VDD2.n134 15.6677
R2191 VDD2.n33 VDD2.n32 15.6677
R2192 VDD2.n182 VDD2.n111 13.1884
R2193 VDD2.n81 VDD2.n10 13.1884
R2194 VDD2.n183 VDD2.n109 12.8005
R2195 VDD2.n178 VDD2.n113 12.8005
R2196 VDD2.n138 VDD2.n137 12.8005
R2197 VDD2.n36 VDD2.n35 12.8005
R2198 VDD2.n77 VDD2.n76 12.8005
R2199 VDD2.n82 VDD2.n8 12.8005
R2200 VDD2.n187 VDD2.n186 12.0247
R2201 VDD2.n177 VDD2.n114 12.0247
R2202 VDD2.n141 VDD2.n132 12.0247
R2203 VDD2.n39 VDD2.n30 12.0247
R2204 VDD2.n75 VDD2.n12 12.0247
R2205 VDD2.n86 VDD2.n85 12.0247
R2206 VDD2.n190 VDD2.n107 11.249
R2207 VDD2.n174 VDD2.n173 11.249
R2208 VDD2.n142 VDD2.n130 11.249
R2209 VDD2.n40 VDD2.n28 11.249
R2210 VDD2.n72 VDD2.n71 11.249
R2211 VDD2.n89 VDD2.n6 11.249
R2212 VDD2.n191 VDD2.n105 10.4732
R2213 VDD2.n170 VDD2.n116 10.4732
R2214 VDD2.n146 VDD2.n145 10.4732
R2215 VDD2.n44 VDD2.n43 10.4732
R2216 VDD2.n68 VDD2.n14 10.4732
R2217 VDD2.n90 VDD2.n4 10.4732
R2218 VDD2.n195 VDD2.n194 9.69747
R2219 VDD2.n169 VDD2.n118 9.69747
R2220 VDD2.n149 VDD2.n128 9.69747
R2221 VDD2.n47 VDD2.n26 9.69747
R2222 VDD2.n67 VDD2.n16 9.69747
R2223 VDD2.n94 VDD2.n93 9.69747
R2224 VDD2.n201 VDD2.n200 9.45567
R2225 VDD2.n100 VDD2.n99 9.45567
R2226 VDD2.n161 VDD2.n160 9.3005
R2227 VDD2.n120 VDD2.n119 9.3005
R2228 VDD2.n167 VDD2.n166 9.3005
R2229 VDD2.n169 VDD2.n168 9.3005
R2230 VDD2.n116 VDD2.n115 9.3005
R2231 VDD2.n175 VDD2.n174 9.3005
R2232 VDD2.n177 VDD2.n176 9.3005
R2233 VDD2.n113 VDD2.n110 9.3005
R2234 VDD2.n200 VDD2.n199 9.3005
R2235 VDD2.n103 VDD2.n102 9.3005
R2236 VDD2.n194 VDD2.n193 9.3005
R2237 VDD2.n192 VDD2.n191 9.3005
R2238 VDD2.n107 VDD2.n106 9.3005
R2239 VDD2.n186 VDD2.n185 9.3005
R2240 VDD2.n184 VDD2.n183 9.3005
R2241 VDD2.n159 VDD2.n158 9.3005
R2242 VDD2.n124 VDD2.n123 9.3005
R2243 VDD2.n153 VDD2.n152 9.3005
R2244 VDD2.n151 VDD2.n150 9.3005
R2245 VDD2.n128 VDD2.n127 9.3005
R2246 VDD2.n145 VDD2.n144 9.3005
R2247 VDD2.n143 VDD2.n142 9.3005
R2248 VDD2.n132 VDD2.n131 9.3005
R2249 VDD2.n137 VDD2.n136 9.3005
R2250 VDD2.n99 VDD2.n98 9.3005
R2251 VDD2.n2 VDD2.n1 9.3005
R2252 VDD2.n93 VDD2.n92 9.3005
R2253 VDD2.n91 VDD2.n90 9.3005
R2254 VDD2.n6 VDD2.n5 9.3005
R2255 VDD2.n85 VDD2.n84 9.3005
R2256 VDD2.n83 VDD2.n82 9.3005
R2257 VDD2.n22 VDD2.n21 9.3005
R2258 VDD2.n51 VDD2.n50 9.3005
R2259 VDD2.n49 VDD2.n48 9.3005
R2260 VDD2.n26 VDD2.n25 9.3005
R2261 VDD2.n43 VDD2.n42 9.3005
R2262 VDD2.n41 VDD2.n40 9.3005
R2263 VDD2.n30 VDD2.n29 9.3005
R2264 VDD2.n35 VDD2.n34 9.3005
R2265 VDD2.n57 VDD2.n56 9.3005
R2266 VDD2.n59 VDD2.n58 9.3005
R2267 VDD2.n18 VDD2.n17 9.3005
R2268 VDD2.n65 VDD2.n64 9.3005
R2269 VDD2.n67 VDD2.n66 9.3005
R2270 VDD2.n14 VDD2.n13 9.3005
R2271 VDD2.n73 VDD2.n72 9.3005
R2272 VDD2.n75 VDD2.n74 9.3005
R2273 VDD2.n76 VDD2.n9 9.3005
R2274 VDD2.n198 VDD2.n103 8.92171
R2275 VDD2.n166 VDD2.n165 8.92171
R2276 VDD2.n150 VDD2.n126 8.92171
R2277 VDD2.n48 VDD2.n24 8.92171
R2278 VDD2.n64 VDD2.n63 8.92171
R2279 VDD2.n97 VDD2.n2 8.92171
R2280 VDD2.n199 VDD2.n101 8.14595
R2281 VDD2.n162 VDD2.n120 8.14595
R2282 VDD2.n154 VDD2.n153 8.14595
R2283 VDD2.n52 VDD2.n51 8.14595
R2284 VDD2.n60 VDD2.n18 8.14595
R2285 VDD2.n98 VDD2.n0 8.14595
R2286 VDD2.n161 VDD2.n122 7.3702
R2287 VDD2.n157 VDD2.n124 7.3702
R2288 VDD2.n55 VDD2.n22 7.3702
R2289 VDD2.n59 VDD2.n20 7.3702
R2290 VDD2.n158 VDD2.n122 6.59444
R2291 VDD2.n158 VDD2.n157 6.59444
R2292 VDD2.n56 VDD2.n55 6.59444
R2293 VDD2.n56 VDD2.n20 6.59444
R2294 VDD2.n201 VDD2.n101 5.81868
R2295 VDD2.n162 VDD2.n161 5.81868
R2296 VDD2.n154 VDD2.n124 5.81868
R2297 VDD2.n52 VDD2.n22 5.81868
R2298 VDD2.n60 VDD2.n59 5.81868
R2299 VDD2.n100 VDD2.n0 5.81868
R2300 VDD2.n199 VDD2.n198 5.04292
R2301 VDD2.n165 VDD2.n120 5.04292
R2302 VDD2.n153 VDD2.n126 5.04292
R2303 VDD2.n51 VDD2.n24 5.04292
R2304 VDD2.n63 VDD2.n18 5.04292
R2305 VDD2.n98 VDD2.n97 5.04292
R2306 VDD2.n136 VDD2.n135 4.38563
R2307 VDD2.n34 VDD2.n33 4.38563
R2308 VDD2.n195 VDD2.n103 4.26717
R2309 VDD2.n166 VDD2.n118 4.26717
R2310 VDD2.n150 VDD2.n149 4.26717
R2311 VDD2.n48 VDD2.n47 4.26717
R2312 VDD2.n64 VDD2.n16 4.26717
R2313 VDD2.n94 VDD2.n2 4.26717
R2314 VDD2.n194 VDD2.n105 3.49141
R2315 VDD2.n170 VDD2.n169 3.49141
R2316 VDD2.n146 VDD2.n128 3.49141
R2317 VDD2.n44 VDD2.n26 3.49141
R2318 VDD2.n68 VDD2.n67 3.49141
R2319 VDD2.n93 VDD2.n4 3.49141
R2320 VDD2.n191 VDD2.n190 2.71565
R2321 VDD2.n173 VDD2.n116 2.71565
R2322 VDD2.n145 VDD2.n130 2.71565
R2323 VDD2.n43 VDD2.n28 2.71565
R2324 VDD2.n71 VDD2.n14 2.71565
R2325 VDD2.n90 VDD2.n89 2.71565
R2326 VDD2.n187 VDD2.n107 1.93989
R2327 VDD2.n174 VDD2.n114 1.93989
R2328 VDD2.n142 VDD2.n141 1.93989
R2329 VDD2.n40 VDD2.n39 1.93989
R2330 VDD2.n72 VDD2.n12 1.93989
R2331 VDD2.n86 VDD2.n6 1.93989
R2332 VDD2.n186 VDD2.n109 1.16414
R2333 VDD2.n178 VDD2.n177 1.16414
R2334 VDD2.n138 VDD2.n132 1.16414
R2335 VDD2.n36 VDD2.n30 1.16414
R2336 VDD2.n77 VDD2.n75 1.16414
R2337 VDD2.n85 VDD2.n8 1.16414
R2338 VDD2 VDD2.n202 0.550069
R2339 VDD2.n183 VDD2.n182 0.388379
R2340 VDD2.n113 VDD2.n111 0.388379
R2341 VDD2.n137 VDD2.n134 0.388379
R2342 VDD2.n35 VDD2.n32 0.388379
R2343 VDD2.n76 VDD2.n10 0.388379
R2344 VDD2.n82 VDD2.n81 0.388379
R2345 VDD2.n200 VDD2.n102 0.155672
R2346 VDD2.n193 VDD2.n102 0.155672
R2347 VDD2.n193 VDD2.n192 0.155672
R2348 VDD2.n192 VDD2.n106 0.155672
R2349 VDD2.n185 VDD2.n106 0.155672
R2350 VDD2.n185 VDD2.n184 0.155672
R2351 VDD2.n184 VDD2.n110 0.155672
R2352 VDD2.n176 VDD2.n110 0.155672
R2353 VDD2.n176 VDD2.n175 0.155672
R2354 VDD2.n175 VDD2.n115 0.155672
R2355 VDD2.n168 VDD2.n115 0.155672
R2356 VDD2.n168 VDD2.n167 0.155672
R2357 VDD2.n167 VDD2.n119 0.155672
R2358 VDD2.n160 VDD2.n119 0.155672
R2359 VDD2.n160 VDD2.n159 0.155672
R2360 VDD2.n159 VDD2.n123 0.155672
R2361 VDD2.n152 VDD2.n123 0.155672
R2362 VDD2.n152 VDD2.n151 0.155672
R2363 VDD2.n151 VDD2.n127 0.155672
R2364 VDD2.n144 VDD2.n127 0.155672
R2365 VDD2.n144 VDD2.n143 0.155672
R2366 VDD2.n143 VDD2.n131 0.155672
R2367 VDD2.n136 VDD2.n131 0.155672
R2368 VDD2.n34 VDD2.n29 0.155672
R2369 VDD2.n41 VDD2.n29 0.155672
R2370 VDD2.n42 VDD2.n41 0.155672
R2371 VDD2.n42 VDD2.n25 0.155672
R2372 VDD2.n49 VDD2.n25 0.155672
R2373 VDD2.n50 VDD2.n49 0.155672
R2374 VDD2.n50 VDD2.n21 0.155672
R2375 VDD2.n57 VDD2.n21 0.155672
R2376 VDD2.n58 VDD2.n57 0.155672
R2377 VDD2.n58 VDD2.n17 0.155672
R2378 VDD2.n65 VDD2.n17 0.155672
R2379 VDD2.n66 VDD2.n65 0.155672
R2380 VDD2.n66 VDD2.n13 0.155672
R2381 VDD2.n73 VDD2.n13 0.155672
R2382 VDD2.n74 VDD2.n73 0.155672
R2383 VDD2.n74 VDD2.n9 0.155672
R2384 VDD2.n83 VDD2.n9 0.155672
R2385 VDD2.n84 VDD2.n83 0.155672
R2386 VDD2.n84 VDD2.n5 0.155672
R2387 VDD2.n91 VDD2.n5 0.155672
R2388 VDD2.n92 VDD2.n91 0.155672
R2389 VDD2.n92 VDD2.n1 0.155672
R2390 VDD2.n99 VDD2.n1 0.155672
R2391 VP.n0 VP.t0 333.392
R2392 VP.n0 VP.t1 285.649
R2393 VP VP.n0 0.241678
R2394 VDD1.n96 VDD1.n0 289.615
R2395 VDD1.n197 VDD1.n101 289.615
R2396 VDD1.n97 VDD1.n96 185
R2397 VDD1.n95 VDD1.n94 185
R2398 VDD1.n4 VDD1.n3 185
R2399 VDD1.n89 VDD1.n88 185
R2400 VDD1.n87 VDD1.n86 185
R2401 VDD1.n8 VDD1.n7 185
R2402 VDD1.n81 VDD1.n80 185
R2403 VDD1.n79 VDD1.n10 185
R2404 VDD1.n78 VDD1.n77 185
R2405 VDD1.n13 VDD1.n11 185
R2406 VDD1.n72 VDD1.n71 185
R2407 VDD1.n70 VDD1.n69 185
R2408 VDD1.n17 VDD1.n16 185
R2409 VDD1.n64 VDD1.n63 185
R2410 VDD1.n62 VDD1.n61 185
R2411 VDD1.n21 VDD1.n20 185
R2412 VDD1.n56 VDD1.n55 185
R2413 VDD1.n54 VDD1.n53 185
R2414 VDD1.n25 VDD1.n24 185
R2415 VDD1.n48 VDD1.n47 185
R2416 VDD1.n46 VDD1.n45 185
R2417 VDD1.n29 VDD1.n28 185
R2418 VDD1.n40 VDD1.n39 185
R2419 VDD1.n38 VDD1.n37 185
R2420 VDD1.n33 VDD1.n32 185
R2421 VDD1.n133 VDD1.n132 185
R2422 VDD1.n138 VDD1.n137 185
R2423 VDD1.n140 VDD1.n139 185
R2424 VDD1.n129 VDD1.n128 185
R2425 VDD1.n146 VDD1.n145 185
R2426 VDD1.n148 VDD1.n147 185
R2427 VDD1.n125 VDD1.n124 185
R2428 VDD1.n154 VDD1.n153 185
R2429 VDD1.n156 VDD1.n155 185
R2430 VDD1.n121 VDD1.n120 185
R2431 VDD1.n162 VDD1.n161 185
R2432 VDD1.n164 VDD1.n163 185
R2433 VDD1.n117 VDD1.n116 185
R2434 VDD1.n170 VDD1.n169 185
R2435 VDD1.n172 VDD1.n171 185
R2436 VDD1.n113 VDD1.n112 185
R2437 VDD1.n179 VDD1.n178 185
R2438 VDD1.n180 VDD1.n111 185
R2439 VDD1.n182 VDD1.n181 185
R2440 VDD1.n109 VDD1.n108 185
R2441 VDD1.n188 VDD1.n187 185
R2442 VDD1.n190 VDD1.n189 185
R2443 VDD1.n105 VDD1.n104 185
R2444 VDD1.n196 VDD1.n195 185
R2445 VDD1.n198 VDD1.n197 185
R2446 VDD1.n34 VDD1.t1 147.659
R2447 VDD1.n134 VDD1.t0 147.659
R2448 VDD1.n96 VDD1.n95 104.615
R2449 VDD1.n95 VDD1.n3 104.615
R2450 VDD1.n88 VDD1.n3 104.615
R2451 VDD1.n88 VDD1.n87 104.615
R2452 VDD1.n87 VDD1.n7 104.615
R2453 VDD1.n80 VDD1.n7 104.615
R2454 VDD1.n80 VDD1.n79 104.615
R2455 VDD1.n79 VDD1.n78 104.615
R2456 VDD1.n78 VDD1.n11 104.615
R2457 VDD1.n71 VDD1.n11 104.615
R2458 VDD1.n71 VDD1.n70 104.615
R2459 VDD1.n70 VDD1.n16 104.615
R2460 VDD1.n63 VDD1.n16 104.615
R2461 VDD1.n63 VDD1.n62 104.615
R2462 VDD1.n62 VDD1.n20 104.615
R2463 VDD1.n55 VDD1.n20 104.615
R2464 VDD1.n55 VDD1.n54 104.615
R2465 VDD1.n54 VDD1.n24 104.615
R2466 VDD1.n47 VDD1.n24 104.615
R2467 VDD1.n47 VDD1.n46 104.615
R2468 VDD1.n46 VDD1.n28 104.615
R2469 VDD1.n39 VDD1.n28 104.615
R2470 VDD1.n39 VDD1.n38 104.615
R2471 VDD1.n38 VDD1.n32 104.615
R2472 VDD1.n138 VDD1.n132 104.615
R2473 VDD1.n139 VDD1.n138 104.615
R2474 VDD1.n139 VDD1.n128 104.615
R2475 VDD1.n146 VDD1.n128 104.615
R2476 VDD1.n147 VDD1.n146 104.615
R2477 VDD1.n147 VDD1.n124 104.615
R2478 VDD1.n154 VDD1.n124 104.615
R2479 VDD1.n155 VDD1.n154 104.615
R2480 VDD1.n155 VDD1.n120 104.615
R2481 VDD1.n162 VDD1.n120 104.615
R2482 VDD1.n163 VDD1.n162 104.615
R2483 VDD1.n163 VDD1.n116 104.615
R2484 VDD1.n170 VDD1.n116 104.615
R2485 VDD1.n171 VDD1.n170 104.615
R2486 VDD1.n171 VDD1.n112 104.615
R2487 VDD1.n179 VDD1.n112 104.615
R2488 VDD1.n180 VDD1.n179 104.615
R2489 VDD1.n181 VDD1.n180 104.615
R2490 VDD1.n181 VDD1.n108 104.615
R2491 VDD1.n188 VDD1.n108 104.615
R2492 VDD1.n189 VDD1.n188 104.615
R2493 VDD1.n189 VDD1.n104 104.615
R2494 VDD1.n196 VDD1.n104 104.615
R2495 VDD1.n197 VDD1.n196 104.615
R2496 VDD1 VDD1.n201 95.4231
R2497 VDD1.t1 VDD1.n32 52.3082
R2498 VDD1.t0 VDD1.n132 52.3082
R2499 VDD1 VDD1.n100 51.547
R2500 VDD1.n34 VDD1.n33 15.6677
R2501 VDD1.n134 VDD1.n133 15.6677
R2502 VDD1.n81 VDD1.n10 13.1884
R2503 VDD1.n182 VDD1.n111 13.1884
R2504 VDD1.n82 VDD1.n8 12.8005
R2505 VDD1.n77 VDD1.n12 12.8005
R2506 VDD1.n37 VDD1.n36 12.8005
R2507 VDD1.n137 VDD1.n136 12.8005
R2508 VDD1.n178 VDD1.n177 12.8005
R2509 VDD1.n183 VDD1.n109 12.8005
R2510 VDD1.n86 VDD1.n85 12.0247
R2511 VDD1.n76 VDD1.n13 12.0247
R2512 VDD1.n40 VDD1.n31 12.0247
R2513 VDD1.n140 VDD1.n131 12.0247
R2514 VDD1.n176 VDD1.n113 12.0247
R2515 VDD1.n187 VDD1.n186 12.0247
R2516 VDD1.n89 VDD1.n6 11.249
R2517 VDD1.n73 VDD1.n72 11.249
R2518 VDD1.n41 VDD1.n29 11.249
R2519 VDD1.n141 VDD1.n129 11.249
R2520 VDD1.n173 VDD1.n172 11.249
R2521 VDD1.n190 VDD1.n107 11.249
R2522 VDD1.n90 VDD1.n4 10.4732
R2523 VDD1.n69 VDD1.n15 10.4732
R2524 VDD1.n45 VDD1.n44 10.4732
R2525 VDD1.n145 VDD1.n144 10.4732
R2526 VDD1.n169 VDD1.n115 10.4732
R2527 VDD1.n191 VDD1.n105 10.4732
R2528 VDD1.n94 VDD1.n93 9.69747
R2529 VDD1.n68 VDD1.n17 9.69747
R2530 VDD1.n48 VDD1.n27 9.69747
R2531 VDD1.n148 VDD1.n127 9.69747
R2532 VDD1.n168 VDD1.n117 9.69747
R2533 VDD1.n195 VDD1.n194 9.69747
R2534 VDD1.n100 VDD1.n99 9.45567
R2535 VDD1.n201 VDD1.n200 9.45567
R2536 VDD1.n60 VDD1.n59 9.3005
R2537 VDD1.n19 VDD1.n18 9.3005
R2538 VDD1.n66 VDD1.n65 9.3005
R2539 VDD1.n68 VDD1.n67 9.3005
R2540 VDD1.n15 VDD1.n14 9.3005
R2541 VDD1.n74 VDD1.n73 9.3005
R2542 VDD1.n76 VDD1.n75 9.3005
R2543 VDD1.n12 VDD1.n9 9.3005
R2544 VDD1.n99 VDD1.n98 9.3005
R2545 VDD1.n2 VDD1.n1 9.3005
R2546 VDD1.n93 VDD1.n92 9.3005
R2547 VDD1.n91 VDD1.n90 9.3005
R2548 VDD1.n6 VDD1.n5 9.3005
R2549 VDD1.n85 VDD1.n84 9.3005
R2550 VDD1.n83 VDD1.n82 9.3005
R2551 VDD1.n58 VDD1.n57 9.3005
R2552 VDD1.n23 VDD1.n22 9.3005
R2553 VDD1.n52 VDD1.n51 9.3005
R2554 VDD1.n50 VDD1.n49 9.3005
R2555 VDD1.n27 VDD1.n26 9.3005
R2556 VDD1.n44 VDD1.n43 9.3005
R2557 VDD1.n42 VDD1.n41 9.3005
R2558 VDD1.n31 VDD1.n30 9.3005
R2559 VDD1.n36 VDD1.n35 9.3005
R2560 VDD1.n200 VDD1.n199 9.3005
R2561 VDD1.n103 VDD1.n102 9.3005
R2562 VDD1.n194 VDD1.n193 9.3005
R2563 VDD1.n192 VDD1.n191 9.3005
R2564 VDD1.n107 VDD1.n106 9.3005
R2565 VDD1.n186 VDD1.n185 9.3005
R2566 VDD1.n184 VDD1.n183 9.3005
R2567 VDD1.n123 VDD1.n122 9.3005
R2568 VDD1.n152 VDD1.n151 9.3005
R2569 VDD1.n150 VDD1.n149 9.3005
R2570 VDD1.n127 VDD1.n126 9.3005
R2571 VDD1.n144 VDD1.n143 9.3005
R2572 VDD1.n142 VDD1.n141 9.3005
R2573 VDD1.n131 VDD1.n130 9.3005
R2574 VDD1.n136 VDD1.n135 9.3005
R2575 VDD1.n158 VDD1.n157 9.3005
R2576 VDD1.n160 VDD1.n159 9.3005
R2577 VDD1.n119 VDD1.n118 9.3005
R2578 VDD1.n166 VDD1.n165 9.3005
R2579 VDD1.n168 VDD1.n167 9.3005
R2580 VDD1.n115 VDD1.n114 9.3005
R2581 VDD1.n174 VDD1.n173 9.3005
R2582 VDD1.n176 VDD1.n175 9.3005
R2583 VDD1.n177 VDD1.n110 9.3005
R2584 VDD1.n97 VDD1.n2 8.92171
R2585 VDD1.n65 VDD1.n64 8.92171
R2586 VDD1.n49 VDD1.n25 8.92171
R2587 VDD1.n149 VDD1.n125 8.92171
R2588 VDD1.n165 VDD1.n164 8.92171
R2589 VDD1.n198 VDD1.n103 8.92171
R2590 VDD1.n98 VDD1.n0 8.14595
R2591 VDD1.n61 VDD1.n19 8.14595
R2592 VDD1.n53 VDD1.n52 8.14595
R2593 VDD1.n153 VDD1.n152 8.14595
R2594 VDD1.n161 VDD1.n119 8.14595
R2595 VDD1.n199 VDD1.n101 8.14595
R2596 VDD1.n60 VDD1.n21 7.3702
R2597 VDD1.n56 VDD1.n23 7.3702
R2598 VDD1.n156 VDD1.n123 7.3702
R2599 VDD1.n160 VDD1.n121 7.3702
R2600 VDD1.n57 VDD1.n21 6.59444
R2601 VDD1.n57 VDD1.n56 6.59444
R2602 VDD1.n157 VDD1.n156 6.59444
R2603 VDD1.n157 VDD1.n121 6.59444
R2604 VDD1.n100 VDD1.n0 5.81868
R2605 VDD1.n61 VDD1.n60 5.81868
R2606 VDD1.n53 VDD1.n23 5.81868
R2607 VDD1.n153 VDD1.n123 5.81868
R2608 VDD1.n161 VDD1.n160 5.81868
R2609 VDD1.n201 VDD1.n101 5.81868
R2610 VDD1.n98 VDD1.n97 5.04292
R2611 VDD1.n64 VDD1.n19 5.04292
R2612 VDD1.n52 VDD1.n25 5.04292
R2613 VDD1.n152 VDD1.n125 5.04292
R2614 VDD1.n164 VDD1.n119 5.04292
R2615 VDD1.n199 VDD1.n198 5.04292
R2616 VDD1.n35 VDD1.n34 4.38563
R2617 VDD1.n135 VDD1.n134 4.38563
R2618 VDD1.n94 VDD1.n2 4.26717
R2619 VDD1.n65 VDD1.n17 4.26717
R2620 VDD1.n49 VDD1.n48 4.26717
R2621 VDD1.n149 VDD1.n148 4.26717
R2622 VDD1.n165 VDD1.n117 4.26717
R2623 VDD1.n195 VDD1.n103 4.26717
R2624 VDD1.n93 VDD1.n4 3.49141
R2625 VDD1.n69 VDD1.n68 3.49141
R2626 VDD1.n45 VDD1.n27 3.49141
R2627 VDD1.n145 VDD1.n127 3.49141
R2628 VDD1.n169 VDD1.n168 3.49141
R2629 VDD1.n194 VDD1.n105 3.49141
R2630 VDD1.n90 VDD1.n89 2.71565
R2631 VDD1.n72 VDD1.n15 2.71565
R2632 VDD1.n44 VDD1.n29 2.71565
R2633 VDD1.n144 VDD1.n129 2.71565
R2634 VDD1.n172 VDD1.n115 2.71565
R2635 VDD1.n191 VDD1.n190 2.71565
R2636 VDD1.n86 VDD1.n6 1.93989
R2637 VDD1.n73 VDD1.n13 1.93989
R2638 VDD1.n41 VDD1.n40 1.93989
R2639 VDD1.n141 VDD1.n140 1.93989
R2640 VDD1.n173 VDD1.n113 1.93989
R2641 VDD1.n187 VDD1.n107 1.93989
R2642 VDD1.n85 VDD1.n8 1.16414
R2643 VDD1.n77 VDD1.n76 1.16414
R2644 VDD1.n37 VDD1.n31 1.16414
R2645 VDD1.n137 VDD1.n131 1.16414
R2646 VDD1.n178 VDD1.n176 1.16414
R2647 VDD1.n186 VDD1.n109 1.16414
R2648 VDD1.n82 VDD1.n81 0.388379
R2649 VDD1.n12 VDD1.n10 0.388379
R2650 VDD1.n36 VDD1.n33 0.388379
R2651 VDD1.n136 VDD1.n133 0.388379
R2652 VDD1.n177 VDD1.n111 0.388379
R2653 VDD1.n183 VDD1.n182 0.388379
R2654 VDD1.n99 VDD1.n1 0.155672
R2655 VDD1.n92 VDD1.n1 0.155672
R2656 VDD1.n92 VDD1.n91 0.155672
R2657 VDD1.n91 VDD1.n5 0.155672
R2658 VDD1.n84 VDD1.n5 0.155672
R2659 VDD1.n84 VDD1.n83 0.155672
R2660 VDD1.n83 VDD1.n9 0.155672
R2661 VDD1.n75 VDD1.n9 0.155672
R2662 VDD1.n75 VDD1.n74 0.155672
R2663 VDD1.n74 VDD1.n14 0.155672
R2664 VDD1.n67 VDD1.n14 0.155672
R2665 VDD1.n67 VDD1.n66 0.155672
R2666 VDD1.n66 VDD1.n18 0.155672
R2667 VDD1.n59 VDD1.n18 0.155672
R2668 VDD1.n59 VDD1.n58 0.155672
R2669 VDD1.n58 VDD1.n22 0.155672
R2670 VDD1.n51 VDD1.n22 0.155672
R2671 VDD1.n51 VDD1.n50 0.155672
R2672 VDD1.n50 VDD1.n26 0.155672
R2673 VDD1.n43 VDD1.n26 0.155672
R2674 VDD1.n43 VDD1.n42 0.155672
R2675 VDD1.n42 VDD1.n30 0.155672
R2676 VDD1.n35 VDD1.n30 0.155672
R2677 VDD1.n135 VDD1.n130 0.155672
R2678 VDD1.n142 VDD1.n130 0.155672
R2679 VDD1.n143 VDD1.n142 0.155672
R2680 VDD1.n143 VDD1.n126 0.155672
R2681 VDD1.n150 VDD1.n126 0.155672
R2682 VDD1.n151 VDD1.n150 0.155672
R2683 VDD1.n151 VDD1.n122 0.155672
R2684 VDD1.n158 VDD1.n122 0.155672
R2685 VDD1.n159 VDD1.n158 0.155672
R2686 VDD1.n159 VDD1.n118 0.155672
R2687 VDD1.n166 VDD1.n118 0.155672
R2688 VDD1.n167 VDD1.n166 0.155672
R2689 VDD1.n167 VDD1.n114 0.155672
R2690 VDD1.n174 VDD1.n114 0.155672
R2691 VDD1.n175 VDD1.n174 0.155672
R2692 VDD1.n175 VDD1.n110 0.155672
R2693 VDD1.n184 VDD1.n110 0.155672
R2694 VDD1.n185 VDD1.n184 0.155672
R2695 VDD1.n185 VDD1.n106 0.155672
R2696 VDD1.n192 VDD1.n106 0.155672
R2697 VDD1.n193 VDD1.n192 0.155672
R2698 VDD1.n193 VDD1.n102 0.155672
R2699 VDD1.n200 VDD1.n102 0.155672
C0 VDD2 VN 3.91482f
C1 VDD2 VTAIL 6.83703f
C2 VN VTAIL 3.25044f
C3 VDD1 VP 4.06912f
C4 VDD2 VP 0.306432f
C5 VP VN 6.32517f
C6 VDD1 VDD2 0.598491f
C7 VP VTAIL 3.26492f
C8 VDD1 VN 0.147824f
C9 VDD1 VTAIL 6.79354f
C10 VDD2 B 5.343853f
C11 VDD1 B 8.45047f
C12 VTAIL B 9.565072f
C13 VN B 11.657411f
C14 VP B 6.014319f
C15 VDD1.n0 B 0.029675f
C16 VDD1.n1 B 0.020054f
C17 VDD1.n2 B 0.010776f
C18 VDD1.n3 B 0.02547f
C19 VDD1.n4 B 0.01141f
C20 VDD1.n5 B 0.020054f
C21 VDD1.n6 B 0.010776f
C22 VDD1.n7 B 0.02547f
C23 VDD1.n8 B 0.01141f
C24 VDD1.n9 B 0.020054f
C25 VDD1.n10 B 0.011093f
C26 VDD1.n11 B 0.02547f
C27 VDD1.n12 B 0.010776f
C28 VDD1.n13 B 0.01141f
C29 VDD1.n14 B 0.020054f
C30 VDD1.n15 B 0.010776f
C31 VDD1.n16 B 0.02547f
C32 VDD1.n17 B 0.01141f
C33 VDD1.n18 B 0.020054f
C34 VDD1.n19 B 0.010776f
C35 VDD1.n20 B 0.02547f
C36 VDD1.n21 B 0.01141f
C37 VDD1.n22 B 0.020054f
C38 VDD1.n23 B 0.010776f
C39 VDD1.n24 B 0.02547f
C40 VDD1.n25 B 0.01141f
C41 VDD1.n26 B 0.020054f
C42 VDD1.n27 B 0.010776f
C43 VDD1.n28 B 0.02547f
C44 VDD1.n29 B 0.01141f
C45 VDD1.n30 B 0.020054f
C46 VDD1.n31 B 0.010776f
C47 VDD1.n32 B 0.019103f
C48 VDD1.n33 B 0.015046f
C49 VDD1.t1 B 0.042228f
C50 VDD1.n34 B 0.147637f
C51 VDD1.n35 B 1.6126f
C52 VDD1.n36 B 0.010776f
C53 VDD1.n37 B 0.01141f
C54 VDD1.n38 B 0.02547f
C55 VDD1.n39 B 0.02547f
C56 VDD1.n40 B 0.01141f
C57 VDD1.n41 B 0.010776f
C58 VDD1.n42 B 0.020054f
C59 VDD1.n43 B 0.020054f
C60 VDD1.n44 B 0.010776f
C61 VDD1.n45 B 0.01141f
C62 VDD1.n46 B 0.02547f
C63 VDD1.n47 B 0.02547f
C64 VDD1.n48 B 0.01141f
C65 VDD1.n49 B 0.010776f
C66 VDD1.n50 B 0.020054f
C67 VDD1.n51 B 0.020054f
C68 VDD1.n52 B 0.010776f
C69 VDD1.n53 B 0.01141f
C70 VDD1.n54 B 0.02547f
C71 VDD1.n55 B 0.02547f
C72 VDD1.n56 B 0.01141f
C73 VDD1.n57 B 0.010776f
C74 VDD1.n58 B 0.020054f
C75 VDD1.n59 B 0.020054f
C76 VDD1.n60 B 0.010776f
C77 VDD1.n61 B 0.01141f
C78 VDD1.n62 B 0.02547f
C79 VDD1.n63 B 0.02547f
C80 VDD1.n64 B 0.01141f
C81 VDD1.n65 B 0.010776f
C82 VDD1.n66 B 0.020054f
C83 VDD1.n67 B 0.020054f
C84 VDD1.n68 B 0.010776f
C85 VDD1.n69 B 0.01141f
C86 VDD1.n70 B 0.02547f
C87 VDD1.n71 B 0.02547f
C88 VDD1.n72 B 0.01141f
C89 VDD1.n73 B 0.010776f
C90 VDD1.n74 B 0.020054f
C91 VDD1.n75 B 0.020054f
C92 VDD1.n76 B 0.010776f
C93 VDD1.n77 B 0.01141f
C94 VDD1.n78 B 0.02547f
C95 VDD1.n79 B 0.02547f
C96 VDD1.n80 B 0.02547f
C97 VDD1.n81 B 0.011093f
C98 VDD1.n82 B 0.010776f
C99 VDD1.n83 B 0.020054f
C100 VDD1.n84 B 0.020054f
C101 VDD1.n85 B 0.010776f
C102 VDD1.n86 B 0.01141f
C103 VDD1.n87 B 0.02547f
C104 VDD1.n88 B 0.02547f
C105 VDD1.n89 B 0.01141f
C106 VDD1.n90 B 0.010776f
C107 VDD1.n91 B 0.020054f
C108 VDD1.n92 B 0.020054f
C109 VDD1.n93 B 0.010776f
C110 VDD1.n94 B 0.01141f
C111 VDD1.n95 B 0.02547f
C112 VDD1.n96 B 0.057771f
C113 VDD1.n97 B 0.01141f
C114 VDD1.n98 B 0.010776f
C115 VDD1.n99 B 0.049366f
C116 VDD1.n100 B 0.047319f
C117 VDD1.n101 B 0.029675f
C118 VDD1.n102 B 0.020054f
C119 VDD1.n103 B 0.010776f
C120 VDD1.n104 B 0.02547f
C121 VDD1.n105 B 0.01141f
C122 VDD1.n106 B 0.020054f
C123 VDD1.n107 B 0.010776f
C124 VDD1.n108 B 0.02547f
C125 VDD1.n109 B 0.01141f
C126 VDD1.n110 B 0.020054f
C127 VDD1.n111 B 0.011093f
C128 VDD1.n112 B 0.02547f
C129 VDD1.n113 B 0.01141f
C130 VDD1.n114 B 0.020054f
C131 VDD1.n115 B 0.010776f
C132 VDD1.n116 B 0.02547f
C133 VDD1.n117 B 0.01141f
C134 VDD1.n118 B 0.020054f
C135 VDD1.n119 B 0.010776f
C136 VDD1.n120 B 0.02547f
C137 VDD1.n121 B 0.01141f
C138 VDD1.n122 B 0.020054f
C139 VDD1.n123 B 0.010776f
C140 VDD1.n124 B 0.02547f
C141 VDD1.n125 B 0.01141f
C142 VDD1.n126 B 0.020054f
C143 VDD1.n127 B 0.010776f
C144 VDD1.n128 B 0.02547f
C145 VDD1.n129 B 0.01141f
C146 VDD1.n130 B 0.020054f
C147 VDD1.n131 B 0.010776f
C148 VDD1.n132 B 0.019103f
C149 VDD1.n133 B 0.015046f
C150 VDD1.t0 B 0.042228f
C151 VDD1.n134 B 0.147637f
C152 VDD1.n135 B 1.6126f
C153 VDD1.n136 B 0.010776f
C154 VDD1.n137 B 0.01141f
C155 VDD1.n138 B 0.02547f
C156 VDD1.n139 B 0.02547f
C157 VDD1.n140 B 0.01141f
C158 VDD1.n141 B 0.010776f
C159 VDD1.n142 B 0.020054f
C160 VDD1.n143 B 0.020054f
C161 VDD1.n144 B 0.010776f
C162 VDD1.n145 B 0.01141f
C163 VDD1.n146 B 0.02547f
C164 VDD1.n147 B 0.02547f
C165 VDD1.n148 B 0.01141f
C166 VDD1.n149 B 0.010776f
C167 VDD1.n150 B 0.020054f
C168 VDD1.n151 B 0.020054f
C169 VDD1.n152 B 0.010776f
C170 VDD1.n153 B 0.01141f
C171 VDD1.n154 B 0.02547f
C172 VDD1.n155 B 0.02547f
C173 VDD1.n156 B 0.01141f
C174 VDD1.n157 B 0.010776f
C175 VDD1.n158 B 0.020054f
C176 VDD1.n159 B 0.020054f
C177 VDD1.n160 B 0.010776f
C178 VDD1.n161 B 0.01141f
C179 VDD1.n162 B 0.02547f
C180 VDD1.n163 B 0.02547f
C181 VDD1.n164 B 0.01141f
C182 VDD1.n165 B 0.010776f
C183 VDD1.n166 B 0.020054f
C184 VDD1.n167 B 0.020054f
C185 VDD1.n168 B 0.010776f
C186 VDD1.n169 B 0.01141f
C187 VDD1.n170 B 0.02547f
C188 VDD1.n171 B 0.02547f
C189 VDD1.n172 B 0.01141f
C190 VDD1.n173 B 0.010776f
C191 VDD1.n174 B 0.020054f
C192 VDD1.n175 B 0.020054f
C193 VDD1.n176 B 0.010776f
C194 VDD1.n177 B 0.010776f
C195 VDD1.n178 B 0.01141f
C196 VDD1.n179 B 0.02547f
C197 VDD1.n180 B 0.02547f
C198 VDD1.n181 B 0.02547f
C199 VDD1.n182 B 0.011093f
C200 VDD1.n183 B 0.010776f
C201 VDD1.n184 B 0.020054f
C202 VDD1.n185 B 0.020054f
C203 VDD1.n186 B 0.010776f
C204 VDD1.n187 B 0.01141f
C205 VDD1.n188 B 0.02547f
C206 VDD1.n189 B 0.02547f
C207 VDD1.n190 B 0.01141f
C208 VDD1.n191 B 0.010776f
C209 VDD1.n192 B 0.020054f
C210 VDD1.n193 B 0.020054f
C211 VDD1.n194 B 0.010776f
C212 VDD1.n195 B 0.01141f
C213 VDD1.n196 B 0.02547f
C214 VDD1.n197 B 0.057771f
C215 VDD1.n198 B 0.01141f
C216 VDD1.n199 B 0.010776f
C217 VDD1.n200 B 0.049366f
C218 VDD1.n201 B 0.767798f
C219 VP.t0 B 4.24305f
C220 VP.t1 B 3.80957f
C221 VP.n0 B 5.5887f
C222 VDD2.n0 B 0.02933f
C223 VDD2.n1 B 0.01982f
C224 VDD2.n2 B 0.010651f
C225 VDD2.n3 B 0.025174f
C226 VDD2.n4 B 0.011277f
C227 VDD2.n5 B 0.01982f
C228 VDD2.n6 B 0.010651f
C229 VDD2.n7 B 0.025174f
C230 VDD2.n8 B 0.011277f
C231 VDD2.n9 B 0.01982f
C232 VDD2.n10 B 0.010964f
C233 VDD2.n11 B 0.025174f
C234 VDD2.n12 B 0.011277f
C235 VDD2.n13 B 0.01982f
C236 VDD2.n14 B 0.010651f
C237 VDD2.n15 B 0.025174f
C238 VDD2.n16 B 0.011277f
C239 VDD2.n17 B 0.01982f
C240 VDD2.n18 B 0.010651f
C241 VDD2.n19 B 0.025174f
C242 VDD2.n20 B 0.011277f
C243 VDD2.n21 B 0.01982f
C244 VDD2.n22 B 0.010651f
C245 VDD2.n23 B 0.025174f
C246 VDD2.n24 B 0.011277f
C247 VDD2.n25 B 0.01982f
C248 VDD2.n26 B 0.010651f
C249 VDD2.n27 B 0.025174f
C250 VDD2.n28 B 0.011277f
C251 VDD2.n29 B 0.01982f
C252 VDD2.n30 B 0.010651f
C253 VDD2.n31 B 0.018881f
C254 VDD2.n32 B 0.014871f
C255 VDD2.t1 B 0.041737f
C256 VDD2.n33 B 0.14592f
C257 VDD2.n34 B 1.59384f
C258 VDD2.n35 B 0.010651f
C259 VDD2.n36 B 0.011277f
C260 VDD2.n37 B 0.025174f
C261 VDD2.n38 B 0.025174f
C262 VDD2.n39 B 0.011277f
C263 VDD2.n40 B 0.010651f
C264 VDD2.n41 B 0.01982f
C265 VDD2.n42 B 0.01982f
C266 VDD2.n43 B 0.010651f
C267 VDD2.n44 B 0.011277f
C268 VDD2.n45 B 0.025174f
C269 VDD2.n46 B 0.025174f
C270 VDD2.n47 B 0.011277f
C271 VDD2.n48 B 0.010651f
C272 VDD2.n49 B 0.01982f
C273 VDD2.n50 B 0.01982f
C274 VDD2.n51 B 0.010651f
C275 VDD2.n52 B 0.011277f
C276 VDD2.n53 B 0.025174f
C277 VDD2.n54 B 0.025174f
C278 VDD2.n55 B 0.011277f
C279 VDD2.n56 B 0.010651f
C280 VDD2.n57 B 0.01982f
C281 VDD2.n58 B 0.01982f
C282 VDD2.n59 B 0.010651f
C283 VDD2.n60 B 0.011277f
C284 VDD2.n61 B 0.025174f
C285 VDD2.n62 B 0.025174f
C286 VDD2.n63 B 0.011277f
C287 VDD2.n64 B 0.010651f
C288 VDD2.n65 B 0.01982f
C289 VDD2.n66 B 0.01982f
C290 VDD2.n67 B 0.010651f
C291 VDD2.n68 B 0.011277f
C292 VDD2.n69 B 0.025174f
C293 VDD2.n70 B 0.025174f
C294 VDD2.n71 B 0.011277f
C295 VDD2.n72 B 0.010651f
C296 VDD2.n73 B 0.01982f
C297 VDD2.n74 B 0.01982f
C298 VDD2.n75 B 0.010651f
C299 VDD2.n76 B 0.010651f
C300 VDD2.n77 B 0.011277f
C301 VDD2.n78 B 0.025174f
C302 VDD2.n79 B 0.025174f
C303 VDD2.n80 B 0.025174f
C304 VDD2.n81 B 0.010964f
C305 VDD2.n82 B 0.010651f
C306 VDD2.n83 B 0.01982f
C307 VDD2.n84 B 0.01982f
C308 VDD2.n85 B 0.010651f
C309 VDD2.n86 B 0.011277f
C310 VDD2.n87 B 0.025174f
C311 VDD2.n88 B 0.025174f
C312 VDD2.n89 B 0.011277f
C313 VDD2.n90 B 0.010651f
C314 VDD2.n91 B 0.01982f
C315 VDD2.n92 B 0.01982f
C316 VDD2.n93 B 0.010651f
C317 VDD2.n94 B 0.011277f
C318 VDD2.n95 B 0.025174f
C319 VDD2.n96 B 0.057099f
C320 VDD2.n97 B 0.011277f
C321 VDD2.n98 B 0.010651f
C322 VDD2.n99 B 0.048792f
C323 VDD2.n100 B 0.721593f
C324 VDD2.n101 B 0.02933f
C325 VDD2.n102 B 0.01982f
C326 VDD2.n103 B 0.010651f
C327 VDD2.n104 B 0.025174f
C328 VDD2.n105 B 0.011277f
C329 VDD2.n106 B 0.01982f
C330 VDD2.n107 B 0.010651f
C331 VDD2.n108 B 0.025174f
C332 VDD2.n109 B 0.011277f
C333 VDD2.n110 B 0.01982f
C334 VDD2.n111 B 0.010964f
C335 VDD2.n112 B 0.025174f
C336 VDD2.n113 B 0.010651f
C337 VDD2.n114 B 0.011277f
C338 VDD2.n115 B 0.01982f
C339 VDD2.n116 B 0.010651f
C340 VDD2.n117 B 0.025174f
C341 VDD2.n118 B 0.011277f
C342 VDD2.n119 B 0.01982f
C343 VDD2.n120 B 0.010651f
C344 VDD2.n121 B 0.025174f
C345 VDD2.n122 B 0.011277f
C346 VDD2.n123 B 0.01982f
C347 VDD2.n124 B 0.010651f
C348 VDD2.n125 B 0.025174f
C349 VDD2.n126 B 0.011277f
C350 VDD2.n127 B 0.01982f
C351 VDD2.n128 B 0.010651f
C352 VDD2.n129 B 0.025174f
C353 VDD2.n130 B 0.011277f
C354 VDD2.n131 B 0.01982f
C355 VDD2.n132 B 0.010651f
C356 VDD2.n133 B 0.018881f
C357 VDD2.n134 B 0.014871f
C358 VDD2.t0 B 0.041737f
C359 VDD2.n135 B 0.14592f
C360 VDD2.n136 B 1.59384f
C361 VDD2.n137 B 0.010651f
C362 VDD2.n138 B 0.011277f
C363 VDD2.n139 B 0.025174f
C364 VDD2.n140 B 0.025174f
C365 VDD2.n141 B 0.011277f
C366 VDD2.n142 B 0.010651f
C367 VDD2.n143 B 0.01982f
C368 VDD2.n144 B 0.01982f
C369 VDD2.n145 B 0.010651f
C370 VDD2.n146 B 0.011277f
C371 VDD2.n147 B 0.025174f
C372 VDD2.n148 B 0.025174f
C373 VDD2.n149 B 0.011277f
C374 VDD2.n150 B 0.010651f
C375 VDD2.n151 B 0.01982f
C376 VDD2.n152 B 0.01982f
C377 VDD2.n153 B 0.010651f
C378 VDD2.n154 B 0.011277f
C379 VDD2.n155 B 0.025174f
C380 VDD2.n156 B 0.025174f
C381 VDD2.n157 B 0.011277f
C382 VDD2.n158 B 0.010651f
C383 VDD2.n159 B 0.01982f
C384 VDD2.n160 B 0.01982f
C385 VDD2.n161 B 0.010651f
C386 VDD2.n162 B 0.011277f
C387 VDD2.n163 B 0.025174f
C388 VDD2.n164 B 0.025174f
C389 VDD2.n165 B 0.011277f
C390 VDD2.n166 B 0.010651f
C391 VDD2.n167 B 0.01982f
C392 VDD2.n168 B 0.01982f
C393 VDD2.n169 B 0.010651f
C394 VDD2.n170 B 0.011277f
C395 VDD2.n171 B 0.025174f
C396 VDD2.n172 B 0.025174f
C397 VDD2.n173 B 0.011277f
C398 VDD2.n174 B 0.010651f
C399 VDD2.n175 B 0.01982f
C400 VDD2.n176 B 0.01982f
C401 VDD2.n177 B 0.010651f
C402 VDD2.n178 B 0.011277f
C403 VDD2.n179 B 0.025174f
C404 VDD2.n180 B 0.025174f
C405 VDD2.n181 B 0.025174f
C406 VDD2.n182 B 0.010964f
C407 VDD2.n183 B 0.010651f
C408 VDD2.n184 B 0.01982f
C409 VDD2.n185 B 0.01982f
C410 VDD2.n186 B 0.010651f
C411 VDD2.n187 B 0.011277f
C412 VDD2.n188 B 0.025174f
C413 VDD2.n189 B 0.025174f
C414 VDD2.n190 B 0.011277f
C415 VDD2.n191 B 0.010651f
C416 VDD2.n192 B 0.01982f
C417 VDD2.n193 B 0.01982f
C418 VDD2.n194 B 0.010651f
C419 VDD2.n195 B 0.011277f
C420 VDD2.n196 B 0.025174f
C421 VDD2.n197 B 0.057099f
C422 VDD2.n198 B 0.011277f
C423 VDD2.n199 B 0.010651f
C424 VDD2.n200 B 0.048792f
C425 VDD2.n201 B 0.045969f
C426 VDD2.n202 B 2.8517f
C427 VTAIL.n0 B 0.029028f
C428 VTAIL.n1 B 0.019616f
C429 VTAIL.n2 B 0.010541f
C430 VTAIL.n3 B 0.024914f
C431 VTAIL.n4 B 0.011161f
C432 VTAIL.n5 B 0.019616f
C433 VTAIL.n6 B 0.010541f
C434 VTAIL.n7 B 0.024914f
C435 VTAIL.n8 B 0.011161f
C436 VTAIL.n9 B 0.019616f
C437 VTAIL.n10 B 0.010851f
C438 VTAIL.n11 B 0.024914f
C439 VTAIL.n12 B 0.011161f
C440 VTAIL.n13 B 0.019616f
C441 VTAIL.n14 B 0.010541f
C442 VTAIL.n15 B 0.024914f
C443 VTAIL.n16 B 0.011161f
C444 VTAIL.n17 B 0.019616f
C445 VTAIL.n18 B 0.010541f
C446 VTAIL.n19 B 0.024914f
C447 VTAIL.n20 B 0.011161f
C448 VTAIL.n21 B 0.019616f
C449 VTAIL.n22 B 0.010541f
C450 VTAIL.n23 B 0.024914f
C451 VTAIL.n24 B 0.011161f
C452 VTAIL.n25 B 0.019616f
C453 VTAIL.n26 B 0.010541f
C454 VTAIL.n27 B 0.024914f
C455 VTAIL.n28 B 0.011161f
C456 VTAIL.n29 B 0.019616f
C457 VTAIL.n30 B 0.010541f
C458 VTAIL.n31 B 0.018686f
C459 VTAIL.n32 B 0.014718f
C460 VTAIL.t0 B 0.041306f
C461 VTAIL.n33 B 0.144414f
C462 VTAIL.n34 B 1.57739f
C463 VTAIL.n35 B 0.010541f
C464 VTAIL.n36 B 0.011161f
C465 VTAIL.n37 B 0.024914f
C466 VTAIL.n38 B 0.024914f
C467 VTAIL.n39 B 0.011161f
C468 VTAIL.n40 B 0.010541f
C469 VTAIL.n41 B 0.019616f
C470 VTAIL.n42 B 0.019616f
C471 VTAIL.n43 B 0.010541f
C472 VTAIL.n44 B 0.011161f
C473 VTAIL.n45 B 0.024914f
C474 VTAIL.n46 B 0.024914f
C475 VTAIL.n47 B 0.011161f
C476 VTAIL.n48 B 0.010541f
C477 VTAIL.n49 B 0.019616f
C478 VTAIL.n50 B 0.019616f
C479 VTAIL.n51 B 0.010541f
C480 VTAIL.n52 B 0.011161f
C481 VTAIL.n53 B 0.024914f
C482 VTAIL.n54 B 0.024914f
C483 VTAIL.n55 B 0.011161f
C484 VTAIL.n56 B 0.010541f
C485 VTAIL.n57 B 0.019616f
C486 VTAIL.n58 B 0.019616f
C487 VTAIL.n59 B 0.010541f
C488 VTAIL.n60 B 0.011161f
C489 VTAIL.n61 B 0.024914f
C490 VTAIL.n62 B 0.024914f
C491 VTAIL.n63 B 0.011161f
C492 VTAIL.n64 B 0.010541f
C493 VTAIL.n65 B 0.019616f
C494 VTAIL.n66 B 0.019616f
C495 VTAIL.n67 B 0.010541f
C496 VTAIL.n68 B 0.011161f
C497 VTAIL.n69 B 0.024914f
C498 VTAIL.n70 B 0.024914f
C499 VTAIL.n71 B 0.011161f
C500 VTAIL.n72 B 0.010541f
C501 VTAIL.n73 B 0.019616f
C502 VTAIL.n74 B 0.019616f
C503 VTAIL.n75 B 0.010541f
C504 VTAIL.n76 B 0.010541f
C505 VTAIL.n77 B 0.011161f
C506 VTAIL.n78 B 0.024914f
C507 VTAIL.n79 B 0.024914f
C508 VTAIL.n80 B 0.024914f
C509 VTAIL.n81 B 0.010851f
C510 VTAIL.n82 B 0.010541f
C511 VTAIL.n83 B 0.019616f
C512 VTAIL.n84 B 0.019616f
C513 VTAIL.n85 B 0.010541f
C514 VTAIL.n86 B 0.011161f
C515 VTAIL.n87 B 0.024914f
C516 VTAIL.n88 B 0.024914f
C517 VTAIL.n89 B 0.011161f
C518 VTAIL.n90 B 0.010541f
C519 VTAIL.n91 B 0.019616f
C520 VTAIL.n92 B 0.019616f
C521 VTAIL.n93 B 0.010541f
C522 VTAIL.n94 B 0.011161f
C523 VTAIL.n95 B 0.024914f
C524 VTAIL.n96 B 0.05651f
C525 VTAIL.n97 B 0.011161f
C526 VTAIL.n98 B 0.010541f
C527 VTAIL.n99 B 0.048289f
C528 VTAIL.n100 B 0.031972f
C529 VTAIL.n101 B 1.59763f
C530 VTAIL.n102 B 0.029028f
C531 VTAIL.n103 B 0.019616f
C532 VTAIL.n104 B 0.010541f
C533 VTAIL.n105 B 0.024914f
C534 VTAIL.n106 B 0.011161f
C535 VTAIL.n107 B 0.019616f
C536 VTAIL.n108 B 0.010541f
C537 VTAIL.n109 B 0.024914f
C538 VTAIL.n110 B 0.011161f
C539 VTAIL.n111 B 0.019616f
C540 VTAIL.n112 B 0.010851f
C541 VTAIL.n113 B 0.024914f
C542 VTAIL.n114 B 0.010541f
C543 VTAIL.n115 B 0.011161f
C544 VTAIL.n116 B 0.019616f
C545 VTAIL.n117 B 0.010541f
C546 VTAIL.n118 B 0.024914f
C547 VTAIL.n119 B 0.011161f
C548 VTAIL.n120 B 0.019616f
C549 VTAIL.n121 B 0.010541f
C550 VTAIL.n122 B 0.024914f
C551 VTAIL.n123 B 0.011161f
C552 VTAIL.n124 B 0.019616f
C553 VTAIL.n125 B 0.010541f
C554 VTAIL.n126 B 0.024914f
C555 VTAIL.n127 B 0.011161f
C556 VTAIL.n128 B 0.019616f
C557 VTAIL.n129 B 0.010541f
C558 VTAIL.n130 B 0.024914f
C559 VTAIL.n131 B 0.011161f
C560 VTAIL.n132 B 0.019616f
C561 VTAIL.n133 B 0.010541f
C562 VTAIL.n134 B 0.018686f
C563 VTAIL.n135 B 0.014718f
C564 VTAIL.t2 B 0.041306f
C565 VTAIL.n136 B 0.144414f
C566 VTAIL.n137 B 1.57739f
C567 VTAIL.n138 B 0.010541f
C568 VTAIL.n139 B 0.011161f
C569 VTAIL.n140 B 0.024914f
C570 VTAIL.n141 B 0.024914f
C571 VTAIL.n142 B 0.011161f
C572 VTAIL.n143 B 0.010541f
C573 VTAIL.n144 B 0.019616f
C574 VTAIL.n145 B 0.019616f
C575 VTAIL.n146 B 0.010541f
C576 VTAIL.n147 B 0.011161f
C577 VTAIL.n148 B 0.024914f
C578 VTAIL.n149 B 0.024914f
C579 VTAIL.n150 B 0.011161f
C580 VTAIL.n151 B 0.010541f
C581 VTAIL.n152 B 0.019616f
C582 VTAIL.n153 B 0.019616f
C583 VTAIL.n154 B 0.010541f
C584 VTAIL.n155 B 0.011161f
C585 VTAIL.n156 B 0.024914f
C586 VTAIL.n157 B 0.024914f
C587 VTAIL.n158 B 0.011161f
C588 VTAIL.n159 B 0.010541f
C589 VTAIL.n160 B 0.019616f
C590 VTAIL.n161 B 0.019616f
C591 VTAIL.n162 B 0.010541f
C592 VTAIL.n163 B 0.011161f
C593 VTAIL.n164 B 0.024914f
C594 VTAIL.n165 B 0.024914f
C595 VTAIL.n166 B 0.011161f
C596 VTAIL.n167 B 0.010541f
C597 VTAIL.n168 B 0.019616f
C598 VTAIL.n169 B 0.019616f
C599 VTAIL.n170 B 0.010541f
C600 VTAIL.n171 B 0.011161f
C601 VTAIL.n172 B 0.024914f
C602 VTAIL.n173 B 0.024914f
C603 VTAIL.n174 B 0.011161f
C604 VTAIL.n175 B 0.010541f
C605 VTAIL.n176 B 0.019616f
C606 VTAIL.n177 B 0.019616f
C607 VTAIL.n178 B 0.010541f
C608 VTAIL.n179 B 0.011161f
C609 VTAIL.n180 B 0.024914f
C610 VTAIL.n181 B 0.024914f
C611 VTAIL.n182 B 0.024914f
C612 VTAIL.n183 B 0.010851f
C613 VTAIL.n184 B 0.010541f
C614 VTAIL.n185 B 0.019616f
C615 VTAIL.n186 B 0.019616f
C616 VTAIL.n187 B 0.010541f
C617 VTAIL.n188 B 0.011161f
C618 VTAIL.n189 B 0.024914f
C619 VTAIL.n190 B 0.024914f
C620 VTAIL.n191 B 0.011161f
C621 VTAIL.n192 B 0.010541f
C622 VTAIL.n193 B 0.019616f
C623 VTAIL.n194 B 0.019616f
C624 VTAIL.n195 B 0.010541f
C625 VTAIL.n196 B 0.011161f
C626 VTAIL.n197 B 0.024914f
C627 VTAIL.n198 B 0.05651f
C628 VTAIL.n199 B 0.011161f
C629 VTAIL.n200 B 0.010541f
C630 VTAIL.n201 B 0.048289f
C631 VTAIL.n202 B 0.031972f
C632 VTAIL.n203 B 1.62502f
C633 VTAIL.n204 B 0.029028f
C634 VTAIL.n205 B 0.019616f
C635 VTAIL.n206 B 0.010541f
C636 VTAIL.n207 B 0.024914f
C637 VTAIL.n208 B 0.011161f
C638 VTAIL.n209 B 0.019616f
C639 VTAIL.n210 B 0.010541f
C640 VTAIL.n211 B 0.024914f
C641 VTAIL.n212 B 0.011161f
C642 VTAIL.n213 B 0.019616f
C643 VTAIL.n214 B 0.010851f
C644 VTAIL.n215 B 0.024914f
C645 VTAIL.n216 B 0.010541f
C646 VTAIL.n217 B 0.011161f
C647 VTAIL.n218 B 0.019616f
C648 VTAIL.n219 B 0.010541f
C649 VTAIL.n220 B 0.024914f
C650 VTAIL.n221 B 0.011161f
C651 VTAIL.n222 B 0.019616f
C652 VTAIL.n223 B 0.010541f
C653 VTAIL.n224 B 0.024914f
C654 VTAIL.n225 B 0.011161f
C655 VTAIL.n226 B 0.019616f
C656 VTAIL.n227 B 0.010541f
C657 VTAIL.n228 B 0.024914f
C658 VTAIL.n229 B 0.011161f
C659 VTAIL.n230 B 0.019616f
C660 VTAIL.n231 B 0.010541f
C661 VTAIL.n232 B 0.024914f
C662 VTAIL.n233 B 0.011161f
C663 VTAIL.n234 B 0.019616f
C664 VTAIL.n235 B 0.010541f
C665 VTAIL.n236 B 0.018686f
C666 VTAIL.n237 B 0.014718f
C667 VTAIL.t1 B 0.041306f
C668 VTAIL.n238 B 0.144414f
C669 VTAIL.n239 B 1.57739f
C670 VTAIL.n240 B 0.010541f
C671 VTAIL.n241 B 0.011161f
C672 VTAIL.n242 B 0.024914f
C673 VTAIL.n243 B 0.024914f
C674 VTAIL.n244 B 0.011161f
C675 VTAIL.n245 B 0.010541f
C676 VTAIL.n246 B 0.019616f
C677 VTAIL.n247 B 0.019616f
C678 VTAIL.n248 B 0.010541f
C679 VTAIL.n249 B 0.011161f
C680 VTAIL.n250 B 0.024914f
C681 VTAIL.n251 B 0.024914f
C682 VTAIL.n252 B 0.011161f
C683 VTAIL.n253 B 0.010541f
C684 VTAIL.n254 B 0.019616f
C685 VTAIL.n255 B 0.019616f
C686 VTAIL.n256 B 0.010541f
C687 VTAIL.n257 B 0.011161f
C688 VTAIL.n258 B 0.024914f
C689 VTAIL.n259 B 0.024914f
C690 VTAIL.n260 B 0.011161f
C691 VTAIL.n261 B 0.010541f
C692 VTAIL.n262 B 0.019616f
C693 VTAIL.n263 B 0.019616f
C694 VTAIL.n264 B 0.010541f
C695 VTAIL.n265 B 0.011161f
C696 VTAIL.n266 B 0.024914f
C697 VTAIL.n267 B 0.024914f
C698 VTAIL.n268 B 0.011161f
C699 VTAIL.n269 B 0.010541f
C700 VTAIL.n270 B 0.019616f
C701 VTAIL.n271 B 0.019616f
C702 VTAIL.n272 B 0.010541f
C703 VTAIL.n273 B 0.011161f
C704 VTAIL.n274 B 0.024914f
C705 VTAIL.n275 B 0.024914f
C706 VTAIL.n276 B 0.011161f
C707 VTAIL.n277 B 0.010541f
C708 VTAIL.n278 B 0.019616f
C709 VTAIL.n279 B 0.019616f
C710 VTAIL.n280 B 0.010541f
C711 VTAIL.n281 B 0.011161f
C712 VTAIL.n282 B 0.024914f
C713 VTAIL.n283 B 0.024914f
C714 VTAIL.n284 B 0.024914f
C715 VTAIL.n285 B 0.010851f
C716 VTAIL.n286 B 0.010541f
C717 VTAIL.n287 B 0.019616f
C718 VTAIL.n288 B 0.019616f
C719 VTAIL.n289 B 0.010541f
C720 VTAIL.n290 B 0.011161f
C721 VTAIL.n291 B 0.024914f
C722 VTAIL.n292 B 0.024914f
C723 VTAIL.n293 B 0.011161f
C724 VTAIL.n294 B 0.010541f
C725 VTAIL.n295 B 0.019616f
C726 VTAIL.n296 B 0.019616f
C727 VTAIL.n297 B 0.010541f
C728 VTAIL.n298 B 0.011161f
C729 VTAIL.n299 B 0.024914f
C730 VTAIL.n300 B 0.05651f
C731 VTAIL.n301 B 0.011161f
C732 VTAIL.n302 B 0.010541f
C733 VTAIL.n303 B 0.048289f
C734 VTAIL.n304 B 0.031972f
C735 VTAIL.n305 B 1.50078f
C736 VTAIL.n306 B 0.029028f
C737 VTAIL.n307 B 0.019616f
C738 VTAIL.n308 B 0.010541f
C739 VTAIL.n309 B 0.024914f
C740 VTAIL.n310 B 0.011161f
C741 VTAIL.n311 B 0.019616f
C742 VTAIL.n312 B 0.010541f
C743 VTAIL.n313 B 0.024914f
C744 VTAIL.n314 B 0.011161f
C745 VTAIL.n315 B 0.019616f
C746 VTAIL.n316 B 0.010851f
C747 VTAIL.n317 B 0.024914f
C748 VTAIL.n318 B 0.011161f
C749 VTAIL.n319 B 0.019616f
C750 VTAIL.n320 B 0.010541f
C751 VTAIL.n321 B 0.024914f
C752 VTAIL.n322 B 0.011161f
C753 VTAIL.n323 B 0.019616f
C754 VTAIL.n324 B 0.010541f
C755 VTAIL.n325 B 0.024914f
C756 VTAIL.n326 B 0.011161f
C757 VTAIL.n327 B 0.019616f
C758 VTAIL.n328 B 0.010541f
C759 VTAIL.n329 B 0.024914f
C760 VTAIL.n330 B 0.011161f
C761 VTAIL.n331 B 0.019616f
C762 VTAIL.n332 B 0.010541f
C763 VTAIL.n333 B 0.024914f
C764 VTAIL.n334 B 0.011161f
C765 VTAIL.n335 B 0.019616f
C766 VTAIL.n336 B 0.010541f
C767 VTAIL.n337 B 0.018686f
C768 VTAIL.n338 B 0.014718f
C769 VTAIL.t3 B 0.041306f
C770 VTAIL.n339 B 0.144414f
C771 VTAIL.n340 B 1.57739f
C772 VTAIL.n341 B 0.010541f
C773 VTAIL.n342 B 0.011161f
C774 VTAIL.n343 B 0.024914f
C775 VTAIL.n344 B 0.024914f
C776 VTAIL.n345 B 0.011161f
C777 VTAIL.n346 B 0.010541f
C778 VTAIL.n347 B 0.019616f
C779 VTAIL.n348 B 0.019616f
C780 VTAIL.n349 B 0.010541f
C781 VTAIL.n350 B 0.011161f
C782 VTAIL.n351 B 0.024914f
C783 VTAIL.n352 B 0.024914f
C784 VTAIL.n353 B 0.011161f
C785 VTAIL.n354 B 0.010541f
C786 VTAIL.n355 B 0.019616f
C787 VTAIL.n356 B 0.019616f
C788 VTAIL.n357 B 0.010541f
C789 VTAIL.n358 B 0.011161f
C790 VTAIL.n359 B 0.024914f
C791 VTAIL.n360 B 0.024914f
C792 VTAIL.n361 B 0.011161f
C793 VTAIL.n362 B 0.010541f
C794 VTAIL.n363 B 0.019616f
C795 VTAIL.n364 B 0.019616f
C796 VTAIL.n365 B 0.010541f
C797 VTAIL.n366 B 0.011161f
C798 VTAIL.n367 B 0.024914f
C799 VTAIL.n368 B 0.024914f
C800 VTAIL.n369 B 0.011161f
C801 VTAIL.n370 B 0.010541f
C802 VTAIL.n371 B 0.019616f
C803 VTAIL.n372 B 0.019616f
C804 VTAIL.n373 B 0.010541f
C805 VTAIL.n374 B 0.011161f
C806 VTAIL.n375 B 0.024914f
C807 VTAIL.n376 B 0.024914f
C808 VTAIL.n377 B 0.011161f
C809 VTAIL.n378 B 0.010541f
C810 VTAIL.n379 B 0.019616f
C811 VTAIL.n380 B 0.019616f
C812 VTAIL.n381 B 0.010541f
C813 VTAIL.n382 B 0.010541f
C814 VTAIL.n383 B 0.011161f
C815 VTAIL.n384 B 0.024914f
C816 VTAIL.n385 B 0.024914f
C817 VTAIL.n386 B 0.024914f
C818 VTAIL.n387 B 0.010851f
C819 VTAIL.n388 B 0.010541f
C820 VTAIL.n389 B 0.019616f
C821 VTAIL.n390 B 0.019616f
C822 VTAIL.n391 B 0.010541f
C823 VTAIL.n392 B 0.011161f
C824 VTAIL.n393 B 0.024914f
C825 VTAIL.n394 B 0.024914f
C826 VTAIL.n395 B 0.011161f
C827 VTAIL.n396 B 0.010541f
C828 VTAIL.n397 B 0.019616f
C829 VTAIL.n398 B 0.019616f
C830 VTAIL.n399 B 0.010541f
C831 VTAIL.n400 B 0.011161f
C832 VTAIL.n401 B 0.024914f
C833 VTAIL.n402 B 0.05651f
C834 VTAIL.n403 B 0.011161f
C835 VTAIL.n404 B 0.010541f
C836 VTAIL.n405 B 0.048289f
C837 VTAIL.n406 B 0.031972f
C838 VTAIL.n407 B 1.43635f
C839 VN.t0 B 3.74127f
C840 VN.t1 B 4.16954f
.ends

