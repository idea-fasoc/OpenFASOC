* NGSPICE file created from diff_pair_sample_1220.ext - technology: sky130A

.subckt diff_pair_sample_1220 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VN.t0 VDD2.t0 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=2.7654 ps=17.09 w=16.76 l=0.86
X1 B.t11 B.t9 B.t10 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=0 ps=0 w=16.76 l=0.86
X2 B.t8 B.t6 B.t7 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=0 ps=0 w=16.76 l=0.86
X3 VTAIL.t3 VP.t0 VDD1.t3 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=2.7654 ps=17.09 w=16.76 l=0.86
X4 VDD2.t1 VN.t1 VTAIL.t6 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=2.7654 pd=17.09 as=6.5364 ps=34.3 w=16.76 l=0.86
X5 VTAIL.t5 VN.t2 VDD2.t3 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=2.7654 ps=17.09 w=16.76 l=0.86
X6 B.t5 B.t3 B.t4 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=0 ps=0 w=16.76 l=0.86
X7 VDD2.t2 VN.t3 VTAIL.t4 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=2.7654 pd=17.09 as=6.5364 ps=34.3 w=16.76 l=0.86
X8 B.t2 B.t0 B.t1 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=0 ps=0 w=16.76 l=0.86
X9 VDD1.t2 VP.t1 VTAIL.t1 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=2.7654 pd=17.09 as=6.5364 ps=34.3 w=16.76 l=0.86
X10 VTAIL.t0 VP.t2 VDD1.t1 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=6.5364 pd=34.3 as=2.7654 ps=17.09 w=16.76 l=0.86
X11 VDD1.t0 VP.t3 VTAIL.t2 w_n1684_n4320# sky130_fd_pr__pfet_01v8 ad=2.7654 pd=17.09 as=6.5364 ps=34.3 w=16.76 l=0.86
R0 VN.n0 VN.t0 536.904
R1 VN.n1 VN.t1 536.904
R2 VN.n0 VN.t3 536.856
R3 VN.n1 VN.t2 536.856
R4 VN VN.n1 89.664
R5 VN VN.n0 44.7132
R6 VDD2.n2 VDD2.n0 109.856
R7 VDD2.n2 VDD2.n1 68.6161
R8 VDD2.n1 VDD2.t3 1.93994
R9 VDD2.n1 VDD2.t1 1.93994
R10 VDD2.n0 VDD2.t0 1.93994
R11 VDD2.n0 VDD2.t2 1.93994
R12 VDD2 VDD2.n2 0.0586897
R13 VTAIL.n746 VTAIL.n658 756.745
R14 VTAIL.n88 VTAIL.n0 756.745
R15 VTAIL.n182 VTAIL.n94 756.745
R16 VTAIL.n276 VTAIL.n188 756.745
R17 VTAIL.n652 VTAIL.n564 756.745
R18 VTAIL.n558 VTAIL.n470 756.745
R19 VTAIL.n464 VTAIL.n376 756.745
R20 VTAIL.n370 VTAIL.n282 756.745
R21 VTAIL.n689 VTAIL.n688 585
R22 VTAIL.n686 VTAIL.n685 585
R23 VTAIL.n695 VTAIL.n694 585
R24 VTAIL.n697 VTAIL.n696 585
R25 VTAIL.n682 VTAIL.n681 585
R26 VTAIL.n703 VTAIL.n702 585
R27 VTAIL.n705 VTAIL.n704 585
R28 VTAIL.n678 VTAIL.n677 585
R29 VTAIL.n711 VTAIL.n710 585
R30 VTAIL.n713 VTAIL.n712 585
R31 VTAIL.n674 VTAIL.n673 585
R32 VTAIL.n719 VTAIL.n718 585
R33 VTAIL.n721 VTAIL.n720 585
R34 VTAIL.n670 VTAIL.n669 585
R35 VTAIL.n727 VTAIL.n726 585
R36 VTAIL.n730 VTAIL.n729 585
R37 VTAIL.n728 VTAIL.n666 585
R38 VTAIL.n735 VTAIL.n665 585
R39 VTAIL.n737 VTAIL.n736 585
R40 VTAIL.n739 VTAIL.n738 585
R41 VTAIL.n662 VTAIL.n661 585
R42 VTAIL.n745 VTAIL.n744 585
R43 VTAIL.n747 VTAIL.n746 585
R44 VTAIL.n31 VTAIL.n30 585
R45 VTAIL.n28 VTAIL.n27 585
R46 VTAIL.n37 VTAIL.n36 585
R47 VTAIL.n39 VTAIL.n38 585
R48 VTAIL.n24 VTAIL.n23 585
R49 VTAIL.n45 VTAIL.n44 585
R50 VTAIL.n47 VTAIL.n46 585
R51 VTAIL.n20 VTAIL.n19 585
R52 VTAIL.n53 VTAIL.n52 585
R53 VTAIL.n55 VTAIL.n54 585
R54 VTAIL.n16 VTAIL.n15 585
R55 VTAIL.n61 VTAIL.n60 585
R56 VTAIL.n63 VTAIL.n62 585
R57 VTAIL.n12 VTAIL.n11 585
R58 VTAIL.n69 VTAIL.n68 585
R59 VTAIL.n72 VTAIL.n71 585
R60 VTAIL.n70 VTAIL.n8 585
R61 VTAIL.n77 VTAIL.n7 585
R62 VTAIL.n79 VTAIL.n78 585
R63 VTAIL.n81 VTAIL.n80 585
R64 VTAIL.n4 VTAIL.n3 585
R65 VTAIL.n87 VTAIL.n86 585
R66 VTAIL.n89 VTAIL.n88 585
R67 VTAIL.n125 VTAIL.n124 585
R68 VTAIL.n122 VTAIL.n121 585
R69 VTAIL.n131 VTAIL.n130 585
R70 VTAIL.n133 VTAIL.n132 585
R71 VTAIL.n118 VTAIL.n117 585
R72 VTAIL.n139 VTAIL.n138 585
R73 VTAIL.n141 VTAIL.n140 585
R74 VTAIL.n114 VTAIL.n113 585
R75 VTAIL.n147 VTAIL.n146 585
R76 VTAIL.n149 VTAIL.n148 585
R77 VTAIL.n110 VTAIL.n109 585
R78 VTAIL.n155 VTAIL.n154 585
R79 VTAIL.n157 VTAIL.n156 585
R80 VTAIL.n106 VTAIL.n105 585
R81 VTAIL.n163 VTAIL.n162 585
R82 VTAIL.n166 VTAIL.n165 585
R83 VTAIL.n164 VTAIL.n102 585
R84 VTAIL.n171 VTAIL.n101 585
R85 VTAIL.n173 VTAIL.n172 585
R86 VTAIL.n175 VTAIL.n174 585
R87 VTAIL.n98 VTAIL.n97 585
R88 VTAIL.n181 VTAIL.n180 585
R89 VTAIL.n183 VTAIL.n182 585
R90 VTAIL.n219 VTAIL.n218 585
R91 VTAIL.n216 VTAIL.n215 585
R92 VTAIL.n225 VTAIL.n224 585
R93 VTAIL.n227 VTAIL.n226 585
R94 VTAIL.n212 VTAIL.n211 585
R95 VTAIL.n233 VTAIL.n232 585
R96 VTAIL.n235 VTAIL.n234 585
R97 VTAIL.n208 VTAIL.n207 585
R98 VTAIL.n241 VTAIL.n240 585
R99 VTAIL.n243 VTAIL.n242 585
R100 VTAIL.n204 VTAIL.n203 585
R101 VTAIL.n249 VTAIL.n248 585
R102 VTAIL.n251 VTAIL.n250 585
R103 VTAIL.n200 VTAIL.n199 585
R104 VTAIL.n257 VTAIL.n256 585
R105 VTAIL.n260 VTAIL.n259 585
R106 VTAIL.n258 VTAIL.n196 585
R107 VTAIL.n265 VTAIL.n195 585
R108 VTAIL.n267 VTAIL.n266 585
R109 VTAIL.n269 VTAIL.n268 585
R110 VTAIL.n192 VTAIL.n191 585
R111 VTAIL.n275 VTAIL.n274 585
R112 VTAIL.n277 VTAIL.n276 585
R113 VTAIL.n653 VTAIL.n652 585
R114 VTAIL.n651 VTAIL.n650 585
R115 VTAIL.n568 VTAIL.n567 585
R116 VTAIL.n645 VTAIL.n644 585
R117 VTAIL.n643 VTAIL.n642 585
R118 VTAIL.n641 VTAIL.n571 585
R119 VTAIL.n575 VTAIL.n572 585
R120 VTAIL.n636 VTAIL.n635 585
R121 VTAIL.n634 VTAIL.n633 585
R122 VTAIL.n577 VTAIL.n576 585
R123 VTAIL.n628 VTAIL.n627 585
R124 VTAIL.n626 VTAIL.n625 585
R125 VTAIL.n581 VTAIL.n580 585
R126 VTAIL.n620 VTAIL.n619 585
R127 VTAIL.n618 VTAIL.n617 585
R128 VTAIL.n585 VTAIL.n584 585
R129 VTAIL.n612 VTAIL.n611 585
R130 VTAIL.n610 VTAIL.n609 585
R131 VTAIL.n589 VTAIL.n588 585
R132 VTAIL.n604 VTAIL.n603 585
R133 VTAIL.n602 VTAIL.n601 585
R134 VTAIL.n593 VTAIL.n592 585
R135 VTAIL.n596 VTAIL.n595 585
R136 VTAIL.n559 VTAIL.n558 585
R137 VTAIL.n557 VTAIL.n556 585
R138 VTAIL.n474 VTAIL.n473 585
R139 VTAIL.n551 VTAIL.n550 585
R140 VTAIL.n549 VTAIL.n548 585
R141 VTAIL.n547 VTAIL.n477 585
R142 VTAIL.n481 VTAIL.n478 585
R143 VTAIL.n542 VTAIL.n541 585
R144 VTAIL.n540 VTAIL.n539 585
R145 VTAIL.n483 VTAIL.n482 585
R146 VTAIL.n534 VTAIL.n533 585
R147 VTAIL.n532 VTAIL.n531 585
R148 VTAIL.n487 VTAIL.n486 585
R149 VTAIL.n526 VTAIL.n525 585
R150 VTAIL.n524 VTAIL.n523 585
R151 VTAIL.n491 VTAIL.n490 585
R152 VTAIL.n518 VTAIL.n517 585
R153 VTAIL.n516 VTAIL.n515 585
R154 VTAIL.n495 VTAIL.n494 585
R155 VTAIL.n510 VTAIL.n509 585
R156 VTAIL.n508 VTAIL.n507 585
R157 VTAIL.n499 VTAIL.n498 585
R158 VTAIL.n502 VTAIL.n501 585
R159 VTAIL.n465 VTAIL.n464 585
R160 VTAIL.n463 VTAIL.n462 585
R161 VTAIL.n380 VTAIL.n379 585
R162 VTAIL.n457 VTAIL.n456 585
R163 VTAIL.n455 VTAIL.n454 585
R164 VTAIL.n453 VTAIL.n383 585
R165 VTAIL.n387 VTAIL.n384 585
R166 VTAIL.n448 VTAIL.n447 585
R167 VTAIL.n446 VTAIL.n445 585
R168 VTAIL.n389 VTAIL.n388 585
R169 VTAIL.n440 VTAIL.n439 585
R170 VTAIL.n438 VTAIL.n437 585
R171 VTAIL.n393 VTAIL.n392 585
R172 VTAIL.n432 VTAIL.n431 585
R173 VTAIL.n430 VTAIL.n429 585
R174 VTAIL.n397 VTAIL.n396 585
R175 VTAIL.n424 VTAIL.n423 585
R176 VTAIL.n422 VTAIL.n421 585
R177 VTAIL.n401 VTAIL.n400 585
R178 VTAIL.n416 VTAIL.n415 585
R179 VTAIL.n414 VTAIL.n413 585
R180 VTAIL.n405 VTAIL.n404 585
R181 VTAIL.n408 VTAIL.n407 585
R182 VTAIL.n371 VTAIL.n370 585
R183 VTAIL.n369 VTAIL.n368 585
R184 VTAIL.n286 VTAIL.n285 585
R185 VTAIL.n363 VTAIL.n362 585
R186 VTAIL.n361 VTAIL.n360 585
R187 VTAIL.n359 VTAIL.n289 585
R188 VTAIL.n293 VTAIL.n290 585
R189 VTAIL.n354 VTAIL.n353 585
R190 VTAIL.n352 VTAIL.n351 585
R191 VTAIL.n295 VTAIL.n294 585
R192 VTAIL.n346 VTAIL.n345 585
R193 VTAIL.n344 VTAIL.n343 585
R194 VTAIL.n299 VTAIL.n298 585
R195 VTAIL.n338 VTAIL.n337 585
R196 VTAIL.n336 VTAIL.n335 585
R197 VTAIL.n303 VTAIL.n302 585
R198 VTAIL.n330 VTAIL.n329 585
R199 VTAIL.n328 VTAIL.n327 585
R200 VTAIL.n307 VTAIL.n306 585
R201 VTAIL.n322 VTAIL.n321 585
R202 VTAIL.n320 VTAIL.n319 585
R203 VTAIL.n311 VTAIL.n310 585
R204 VTAIL.n314 VTAIL.n313 585
R205 VTAIL.t1 VTAIL.n594 327.466
R206 VTAIL.t0 VTAIL.n500 327.466
R207 VTAIL.t6 VTAIL.n406 327.466
R208 VTAIL.t5 VTAIL.n312 327.466
R209 VTAIL.t4 VTAIL.n687 327.466
R210 VTAIL.t7 VTAIL.n29 327.466
R211 VTAIL.t2 VTAIL.n123 327.466
R212 VTAIL.t3 VTAIL.n217 327.466
R213 VTAIL.n688 VTAIL.n685 171.744
R214 VTAIL.n695 VTAIL.n685 171.744
R215 VTAIL.n696 VTAIL.n695 171.744
R216 VTAIL.n696 VTAIL.n681 171.744
R217 VTAIL.n703 VTAIL.n681 171.744
R218 VTAIL.n704 VTAIL.n703 171.744
R219 VTAIL.n704 VTAIL.n677 171.744
R220 VTAIL.n711 VTAIL.n677 171.744
R221 VTAIL.n712 VTAIL.n711 171.744
R222 VTAIL.n712 VTAIL.n673 171.744
R223 VTAIL.n719 VTAIL.n673 171.744
R224 VTAIL.n720 VTAIL.n719 171.744
R225 VTAIL.n720 VTAIL.n669 171.744
R226 VTAIL.n727 VTAIL.n669 171.744
R227 VTAIL.n729 VTAIL.n727 171.744
R228 VTAIL.n729 VTAIL.n728 171.744
R229 VTAIL.n728 VTAIL.n665 171.744
R230 VTAIL.n737 VTAIL.n665 171.744
R231 VTAIL.n738 VTAIL.n737 171.744
R232 VTAIL.n738 VTAIL.n661 171.744
R233 VTAIL.n745 VTAIL.n661 171.744
R234 VTAIL.n746 VTAIL.n745 171.744
R235 VTAIL.n30 VTAIL.n27 171.744
R236 VTAIL.n37 VTAIL.n27 171.744
R237 VTAIL.n38 VTAIL.n37 171.744
R238 VTAIL.n38 VTAIL.n23 171.744
R239 VTAIL.n45 VTAIL.n23 171.744
R240 VTAIL.n46 VTAIL.n45 171.744
R241 VTAIL.n46 VTAIL.n19 171.744
R242 VTAIL.n53 VTAIL.n19 171.744
R243 VTAIL.n54 VTAIL.n53 171.744
R244 VTAIL.n54 VTAIL.n15 171.744
R245 VTAIL.n61 VTAIL.n15 171.744
R246 VTAIL.n62 VTAIL.n61 171.744
R247 VTAIL.n62 VTAIL.n11 171.744
R248 VTAIL.n69 VTAIL.n11 171.744
R249 VTAIL.n71 VTAIL.n69 171.744
R250 VTAIL.n71 VTAIL.n70 171.744
R251 VTAIL.n70 VTAIL.n7 171.744
R252 VTAIL.n79 VTAIL.n7 171.744
R253 VTAIL.n80 VTAIL.n79 171.744
R254 VTAIL.n80 VTAIL.n3 171.744
R255 VTAIL.n87 VTAIL.n3 171.744
R256 VTAIL.n88 VTAIL.n87 171.744
R257 VTAIL.n124 VTAIL.n121 171.744
R258 VTAIL.n131 VTAIL.n121 171.744
R259 VTAIL.n132 VTAIL.n131 171.744
R260 VTAIL.n132 VTAIL.n117 171.744
R261 VTAIL.n139 VTAIL.n117 171.744
R262 VTAIL.n140 VTAIL.n139 171.744
R263 VTAIL.n140 VTAIL.n113 171.744
R264 VTAIL.n147 VTAIL.n113 171.744
R265 VTAIL.n148 VTAIL.n147 171.744
R266 VTAIL.n148 VTAIL.n109 171.744
R267 VTAIL.n155 VTAIL.n109 171.744
R268 VTAIL.n156 VTAIL.n155 171.744
R269 VTAIL.n156 VTAIL.n105 171.744
R270 VTAIL.n163 VTAIL.n105 171.744
R271 VTAIL.n165 VTAIL.n163 171.744
R272 VTAIL.n165 VTAIL.n164 171.744
R273 VTAIL.n164 VTAIL.n101 171.744
R274 VTAIL.n173 VTAIL.n101 171.744
R275 VTAIL.n174 VTAIL.n173 171.744
R276 VTAIL.n174 VTAIL.n97 171.744
R277 VTAIL.n181 VTAIL.n97 171.744
R278 VTAIL.n182 VTAIL.n181 171.744
R279 VTAIL.n218 VTAIL.n215 171.744
R280 VTAIL.n225 VTAIL.n215 171.744
R281 VTAIL.n226 VTAIL.n225 171.744
R282 VTAIL.n226 VTAIL.n211 171.744
R283 VTAIL.n233 VTAIL.n211 171.744
R284 VTAIL.n234 VTAIL.n233 171.744
R285 VTAIL.n234 VTAIL.n207 171.744
R286 VTAIL.n241 VTAIL.n207 171.744
R287 VTAIL.n242 VTAIL.n241 171.744
R288 VTAIL.n242 VTAIL.n203 171.744
R289 VTAIL.n249 VTAIL.n203 171.744
R290 VTAIL.n250 VTAIL.n249 171.744
R291 VTAIL.n250 VTAIL.n199 171.744
R292 VTAIL.n257 VTAIL.n199 171.744
R293 VTAIL.n259 VTAIL.n257 171.744
R294 VTAIL.n259 VTAIL.n258 171.744
R295 VTAIL.n258 VTAIL.n195 171.744
R296 VTAIL.n267 VTAIL.n195 171.744
R297 VTAIL.n268 VTAIL.n267 171.744
R298 VTAIL.n268 VTAIL.n191 171.744
R299 VTAIL.n275 VTAIL.n191 171.744
R300 VTAIL.n276 VTAIL.n275 171.744
R301 VTAIL.n652 VTAIL.n651 171.744
R302 VTAIL.n651 VTAIL.n567 171.744
R303 VTAIL.n644 VTAIL.n567 171.744
R304 VTAIL.n644 VTAIL.n643 171.744
R305 VTAIL.n643 VTAIL.n571 171.744
R306 VTAIL.n575 VTAIL.n571 171.744
R307 VTAIL.n635 VTAIL.n575 171.744
R308 VTAIL.n635 VTAIL.n634 171.744
R309 VTAIL.n634 VTAIL.n576 171.744
R310 VTAIL.n627 VTAIL.n576 171.744
R311 VTAIL.n627 VTAIL.n626 171.744
R312 VTAIL.n626 VTAIL.n580 171.744
R313 VTAIL.n619 VTAIL.n580 171.744
R314 VTAIL.n619 VTAIL.n618 171.744
R315 VTAIL.n618 VTAIL.n584 171.744
R316 VTAIL.n611 VTAIL.n584 171.744
R317 VTAIL.n611 VTAIL.n610 171.744
R318 VTAIL.n610 VTAIL.n588 171.744
R319 VTAIL.n603 VTAIL.n588 171.744
R320 VTAIL.n603 VTAIL.n602 171.744
R321 VTAIL.n602 VTAIL.n592 171.744
R322 VTAIL.n595 VTAIL.n592 171.744
R323 VTAIL.n558 VTAIL.n557 171.744
R324 VTAIL.n557 VTAIL.n473 171.744
R325 VTAIL.n550 VTAIL.n473 171.744
R326 VTAIL.n550 VTAIL.n549 171.744
R327 VTAIL.n549 VTAIL.n477 171.744
R328 VTAIL.n481 VTAIL.n477 171.744
R329 VTAIL.n541 VTAIL.n481 171.744
R330 VTAIL.n541 VTAIL.n540 171.744
R331 VTAIL.n540 VTAIL.n482 171.744
R332 VTAIL.n533 VTAIL.n482 171.744
R333 VTAIL.n533 VTAIL.n532 171.744
R334 VTAIL.n532 VTAIL.n486 171.744
R335 VTAIL.n525 VTAIL.n486 171.744
R336 VTAIL.n525 VTAIL.n524 171.744
R337 VTAIL.n524 VTAIL.n490 171.744
R338 VTAIL.n517 VTAIL.n490 171.744
R339 VTAIL.n517 VTAIL.n516 171.744
R340 VTAIL.n516 VTAIL.n494 171.744
R341 VTAIL.n509 VTAIL.n494 171.744
R342 VTAIL.n509 VTAIL.n508 171.744
R343 VTAIL.n508 VTAIL.n498 171.744
R344 VTAIL.n501 VTAIL.n498 171.744
R345 VTAIL.n464 VTAIL.n463 171.744
R346 VTAIL.n463 VTAIL.n379 171.744
R347 VTAIL.n456 VTAIL.n379 171.744
R348 VTAIL.n456 VTAIL.n455 171.744
R349 VTAIL.n455 VTAIL.n383 171.744
R350 VTAIL.n387 VTAIL.n383 171.744
R351 VTAIL.n447 VTAIL.n387 171.744
R352 VTAIL.n447 VTAIL.n446 171.744
R353 VTAIL.n446 VTAIL.n388 171.744
R354 VTAIL.n439 VTAIL.n388 171.744
R355 VTAIL.n439 VTAIL.n438 171.744
R356 VTAIL.n438 VTAIL.n392 171.744
R357 VTAIL.n431 VTAIL.n392 171.744
R358 VTAIL.n431 VTAIL.n430 171.744
R359 VTAIL.n430 VTAIL.n396 171.744
R360 VTAIL.n423 VTAIL.n396 171.744
R361 VTAIL.n423 VTAIL.n422 171.744
R362 VTAIL.n422 VTAIL.n400 171.744
R363 VTAIL.n415 VTAIL.n400 171.744
R364 VTAIL.n415 VTAIL.n414 171.744
R365 VTAIL.n414 VTAIL.n404 171.744
R366 VTAIL.n407 VTAIL.n404 171.744
R367 VTAIL.n370 VTAIL.n369 171.744
R368 VTAIL.n369 VTAIL.n285 171.744
R369 VTAIL.n362 VTAIL.n285 171.744
R370 VTAIL.n362 VTAIL.n361 171.744
R371 VTAIL.n361 VTAIL.n289 171.744
R372 VTAIL.n293 VTAIL.n289 171.744
R373 VTAIL.n353 VTAIL.n293 171.744
R374 VTAIL.n353 VTAIL.n352 171.744
R375 VTAIL.n352 VTAIL.n294 171.744
R376 VTAIL.n345 VTAIL.n294 171.744
R377 VTAIL.n345 VTAIL.n344 171.744
R378 VTAIL.n344 VTAIL.n298 171.744
R379 VTAIL.n337 VTAIL.n298 171.744
R380 VTAIL.n337 VTAIL.n336 171.744
R381 VTAIL.n336 VTAIL.n302 171.744
R382 VTAIL.n329 VTAIL.n302 171.744
R383 VTAIL.n329 VTAIL.n328 171.744
R384 VTAIL.n328 VTAIL.n306 171.744
R385 VTAIL.n321 VTAIL.n306 171.744
R386 VTAIL.n321 VTAIL.n320 171.744
R387 VTAIL.n320 VTAIL.n310 171.744
R388 VTAIL.n313 VTAIL.n310 171.744
R389 VTAIL.n688 VTAIL.t4 85.8723
R390 VTAIL.n30 VTAIL.t7 85.8723
R391 VTAIL.n124 VTAIL.t2 85.8723
R392 VTAIL.n218 VTAIL.t3 85.8723
R393 VTAIL.n595 VTAIL.t1 85.8723
R394 VTAIL.n501 VTAIL.t0 85.8723
R395 VTAIL.n407 VTAIL.t6 85.8723
R396 VTAIL.n313 VTAIL.t5 85.8723
R397 VTAIL.n751 VTAIL.n750 31.4096
R398 VTAIL.n93 VTAIL.n92 31.4096
R399 VTAIL.n187 VTAIL.n186 31.4096
R400 VTAIL.n281 VTAIL.n280 31.4096
R401 VTAIL.n657 VTAIL.n656 31.4096
R402 VTAIL.n563 VTAIL.n562 31.4096
R403 VTAIL.n469 VTAIL.n468 31.4096
R404 VTAIL.n375 VTAIL.n374 31.4096
R405 VTAIL.n751 VTAIL.n657 27.841
R406 VTAIL.n375 VTAIL.n281 27.841
R407 VTAIL.n689 VTAIL.n687 16.3895
R408 VTAIL.n31 VTAIL.n29 16.3895
R409 VTAIL.n125 VTAIL.n123 16.3895
R410 VTAIL.n219 VTAIL.n217 16.3895
R411 VTAIL.n596 VTAIL.n594 16.3895
R412 VTAIL.n502 VTAIL.n500 16.3895
R413 VTAIL.n408 VTAIL.n406 16.3895
R414 VTAIL.n314 VTAIL.n312 16.3895
R415 VTAIL.n736 VTAIL.n735 13.1884
R416 VTAIL.n78 VTAIL.n77 13.1884
R417 VTAIL.n172 VTAIL.n171 13.1884
R418 VTAIL.n266 VTAIL.n265 13.1884
R419 VTAIL.n642 VTAIL.n641 13.1884
R420 VTAIL.n548 VTAIL.n547 13.1884
R421 VTAIL.n454 VTAIL.n453 13.1884
R422 VTAIL.n360 VTAIL.n359 13.1884
R423 VTAIL.n690 VTAIL.n686 12.8005
R424 VTAIL.n734 VTAIL.n666 12.8005
R425 VTAIL.n739 VTAIL.n664 12.8005
R426 VTAIL.n32 VTAIL.n28 12.8005
R427 VTAIL.n76 VTAIL.n8 12.8005
R428 VTAIL.n81 VTAIL.n6 12.8005
R429 VTAIL.n126 VTAIL.n122 12.8005
R430 VTAIL.n170 VTAIL.n102 12.8005
R431 VTAIL.n175 VTAIL.n100 12.8005
R432 VTAIL.n220 VTAIL.n216 12.8005
R433 VTAIL.n264 VTAIL.n196 12.8005
R434 VTAIL.n269 VTAIL.n194 12.8005
R435 VTAIL.n645 VTAIL.n570 12.8005
R436 VTAIL.n640 VTAIL.n572 12.8005
R437 VTAIL.n597 VTAIL.n593 12.8005
R438 VTAIL.n551 VTAIL.n476 12.8005
R439 VTAIL.n546 VTAIL.n478 12.8005
R440 VTAIL.n503 VTAIL.n499 12.8005
R441 VTAIL.n457 VTAIL.n382 12.8005
R442 VTAIL.n452 VTAIL.n384 12.8005
R443 VTAIL.n409 VTAIL.n405 12.8005
R444 VTAIL.n363 VTAIL.n288 12.8005
R445 VTAIL.n358 VTAIL.n290 12.8005
R446 VTAIL.n315 VTAIL.n311 12.8005
R447 VTAIL.n694 VTAIL.n693 12.0247
R448 VTAIL.n731 VTAIL.n730 12.0247
R449 VTAIL.n740 VTAIL.n662 12.0247
R450 VTAIL.n36 VTAIL.n35 12.0247
R451 VTAIL.n73 VTAIL.n72 12.0247
R452 VTAIL.n82 VTAIL.n4 12.0247
R453 VTAIL.n130 VTAIL.n129 12.0247
R454 VTAIL.n167 VTAIL.n166 12.0247
R455 VTAIL.n176 VTAIL.n98 12.0247
R456 VTAIL.n224 VTAIL.n223 12.0247
R457 VTAIL.n261 VTAIL.n260 12.0247
R458 VTAIL.n270 VTAIL.n192 12.0247
R459 VTAIL.n646 VTAIL.n568 12.0247
R460 VTAIL.n637 VTAIL.n636 12.0247
R461 VTAIL.n601 VTAIL.n600 12.0247
R462 VTAIL.n552 VTAIL.n474 12.0247
R463 VTAIL.n543 VTAIL.n542 12.0247
R464 VTAIL.n507 VTAIL.n506 12.0247
R465 VTAIL.n458 VTAIL.n380 12.0247
R466 VTAIL.n449 VTAIL.n448 12.0247
R467 VTAIL.n413 VTAIL.n412 12.0247
R468 VTAIL.n364 VTAIL.n286 12.0247
R469 VTAIL.n355 VTAIL.n354 12.0247
R470 VTAIL.n319 VTAIL.n318 12.0247
R471 VTAIL.n697 VTAIL.n684 11.249
R472 VTAIL.n726 VTAIL.n668 11.249
R473 VTAIL.n744 VTAIL.n743 11.249
R474 VTAIL.n39 VTAIL.n26 11.249
R475 VTAIL.n68 VTAIL.n10 11.249
R476 VTAIL.n86 VTAIL.n85 11.249
R477 VTAIL.n133 VTAIL.n120 11.249
R478 VTAIL.n162 VTAIL.n104 11.249
R479 VTAIL.n180 VTAIL.n179 11.249
R480 VTAIL.n227 VTAIL.n214 11.249
R481 VTAIL.n256 VTAIL.n198 11.249
R482 VTAIL.n274 VTAIL.n273 11.249
R483 VTAIL.n650 VTAIL.n649 11.249
R484 VTAIL.n633 VTAIL.n574 11.249
R485 VTAIL.n604 VTAIL.n591 11.249
R486 VTAIL.n556 VTAIL.n555 11.249
R487 VTAIL.n539 VTAIL.n480 11.249
R488 VTAIL.n510 VTAIL.n497 11.249
R489 VTAIL.n462 VTAIL.n461 11.249
R490 VTAIL.n445 VTAIL.n386 11.249
R491 VTAIL.n416 VTAIL.n403 11.249
R492 VTAIL.n368 VTAIL.n367 11.249
R493 VTAIL.n351 VTAIL.n292 11.249
R494 VTAIL.n322 VTAIL.n309 11.249
R495 VTAIL.n698 VTAIL.n682 10.4732
R496 VTAIL.n725 VTAIL.n670 10.4732
R497 VTAIL.n747 VTAIL.n660 10.4732
R498 VTAIL.n40 VTAIL.n24 10.4732
R499 VTAIL.n67 VTAIL.n12 10.4732
R500 VTAIL.n89 VTAIL.n2 10.4732
R501 VTAIL.n134 VTAIL.n118 10.4732
R502 VTAIL.n161 VTAIL.n106 10.4732
R503 VTAIL.n183 VTAIL.n96 10.4732
R504 VTAIL.n228 VTAIL.n212 10.4732
R505 VTAIL.n255 VTAIL.n200 10.4732
R506 VTAIL.n277 VTAIL.n190 10.4732
R507 VTAIL.n653 VTAIL.n566 10.4732
R508 VTAIL.n632 VTAIL.n577 10.4732
R509 VTAIL.n605 VTAIL.n589 10.4732
R510 VTAIL.n559 VTAIL.n472 10.4732
R511 VTAIL.n538 VTAIL.n483 10.4732
R512 VTAIL.n511 VTAIL.n495 10.4732
R513 VTAIL.n465 VTAIL.n378 10.4732
R514 VTAIL.n444 VTAIL.n389 10.4732
R515 VTAIL.n417 VTAIL.n401 10.4732
R516 VTAIL.n371 VTAIL.n284 10.4732
R517 VTAIL.n350 VTAIL.n295 10.4732
R518 VTAIL.n323 VTAIL.n307 10.4732
R519 VTAIL.n702 VTAIL.n701 9.69747
R520 VTAIL.n722 VTAIL.n721 9.69747
R521 VTAIL.n748 VTAIL.n658 9.69747
R522 VTAIL.n44 VTAIL.n43 9.69747
R523 VTAIL.n64 VTAIL.n63 9.69747
R524 VTAIL.n90 VTAIL.n0 9.69747
R525 VTAIL.n138 VTAIL.n137 9.69747
R526 VTAIL.n158 VTAIL.n157 9.69747
R527 VTAIL.n184 VTAIL.n94 9.69747
R528 VTAIL.n232 VTAIL.n231 9.69747
R529 VTAIL.n252 VTAIL.n251 9.69747
R530 VTAIL.n278 VTAIL.n188 9.69747
R531 VTAIL.n654 VTAIL.n564 9.69747
R532 VTAIL.n629 VTAIL.n628 9.69747
R533 VTAIL.n609 VTAIL.n608 9.69747
R534 VTAIL.n560 VTAIL.n470 9.69747
R535 VTAIL.n535 VTAIL.n534 9.69747
R536 VTAIL.n515 VTAIL.n514 9.69747
R537 VTAIL.n466 VTAIL.n376 9.69747
R538 VTAIL.n441 VTAIL.n440 9.69747
R539 VTAIL.n421 VTAIL.n420 9.69747
R540 VTAIL.n372 VTAIL.n282 9.69747
R541 VTAIL.n347 VTAIL.n346 9.69747
R542 VTAIL.n327 VTAIL.n326 9.69747
R543 VTAIL.n750 VTAIL.n749 9.45567
R544 VTAIL.n92 VTAIL.n91 9.45567
R545 VTAIL.n186 VTAIL.n185 9.45567
R546 VTAIL.n280 VTAIL.n279 9.45567
R547 VTAIL.n656 VTAIL.n655 9.45567
R548 VTAIL.n562 VTAIL.n561 9.45567
R549 VTAIL.n468 VTAIL.n467 9.45567
R550 VTAIL.n374 VTAIL.n373 9.45567
R551 VTAIL.n749 VTAIL.n748 9.3005
R552 VTAIL.n660 VTAIL.n659 9.3005
R553 VTAIL.n743 VTAIL.n742 9.3005
R554 VTAIL.n741 VTAIL.n740 9.3005
R555 VTAIL.n664 VTAIL.n663 9.3005
R556 VTAIL.n709 VTAIL.n708 9.3005
R557 VTAIL.n707 VTAIL.n706 9.3005
R558 VTAIL.n680 VTAIL.n679 9.3005
R559 VTAIL.n701 VTAIL.n700 9.3005
R560 VTAIL.n699 VTAIL.n698 9.3005
R561 VTAIL.n684 VTAIL.n683 9.3005
R562 VTAIL.n693 VTAIL.n692 9.3005
R563 VTAIL.n691 VTAIL.n690 9.3005
R564 VTAIL.n676 VTAIL.n675 9.3005
R565 VTAIL.n715 VTAIL.n714 9.3005
R566 VTAIL.n717 VTAIL.n716 9.3005
R567 VTAIL.n672 VTAIL.n671 9.3005
R568 VTAIL.n723 VTAIL.n722 9.3005
R569 VTAIL.n725 VTAIL.n724 9.3005
R570 VTAIL.n668 VTAIL.n667 9.3005
R571 VTAIL.n732 VTAIL.n731 9.3005
R572 VTAIL.n734 VTAIL.n733 9.3005
R573 VTAIL.n91 VTAIL.n90 9.3005
R574 VTAIL.n2 VTAIL.n1 9.3005
R575 VTAIL.n85 VTAIL.n84 9.3005
R576 VTAIL.n83 VTAIL.n82 9.3005
R577 VTAIL.n6 VTAIL.n5 9.3005
R578 VTAIL.n51 VTAIL.n50 9.3005
R579 VTAIL.n49 VTAIL.n48 9.3005
R580 VTAIL.n22 VTAIL.n21 9.3005
R581 VTAIL.n43 VTAIL.n42 9.3005
R582 VTAIL.n41 VTAIL.n40 9.3005
R583 VTAIL.n26 VTAIL.n25 9.3005
R584 VTAIL.n35 VTAIL.n34 9.3005
R585 VTAIL.n33 VTAIL.n32 9.3005
R586 VTAIL.n18 VTAIL.n17 9.3005
R587 VTAIL.n57 VTAIL.n56 9.3005
R588 VTAIL.n59 VTAIL.n58 9.3005
R589 VTAIL.n14 VTAIL.n13 9.3005
R590 VTAIL.n65 VTAIL.n64 9.3005
R591 VTAIL.n67 VTAIL.n66 9.3005
R592 VTAIL.n10 VTAIL.n9 9.3005
R593 VTAIL.n74 VTAIL.n73 9.3005
R594 VTAIL.n76 VTAIL.n75 9.3005
R595 VTAIL.n185 VTAIL.n184 9.3005
R596 VTAIL.n96 VTAIL.n95 9.3005
R597 VTAIL.n179 VTAIL.n178 9.3005
R598 VTAIL.n177 VTAIL.n176 9.3005
R599 VTAIL.n100 VTAIL.n99 9.3005
R600 VTAIL.n145 VTAIL.n144 9.3005
R601 VTAIL.n143 VTAIL.n142 9.3005
R602 VTAIL.n116 VTAIL.n115 9.3005
R603 VTAIL.n137 VTAIL.n136 9.3005
R604 VTAIL.n135 VTAIL.n134 9.3005
R605 VTAIL.n120 VTAIL.n119 9.3005
R606 VTAIL.n129 VTAIL.n128 9.3005
R607 VTAIL.n127 VTAIL.n126 9.3005
R608 VTAIL.n112 VTAIL.n111 9.3005
R609 VTAIL.n151 VTAIL.n150 9.3005
R610 VTAIL.n153 VTAIL.n152 9.3005
R611 VTAIL.n108 VTAIL.n107 9.3005
R612 VTAIL.n159 VTAIL.n158 9.3005
R613 VTAIL.n161 VTAIL.n160 9.3005
R614 VTAIL.n104 VTAIL.n103 9.3005
R615 VTAIL.n168 VTAIL.n167 9.3005
R616 VTAIL.n170 VTAIL.n169 9.3005
R617 VTAIL.n279 VTAIL.n278 9.3005
R618 VTAIL.n190 VTAIL.n189 9.3005
R619 VTAIL.n273 VTAIL.n272 9.3005
R620 VTAIL.n271 VTAIL.n270 9.3005
R621 VTAIL.n194 VTAIL.n193 9.3005
R622 VTAIL.n239 VTAIL.n238 9.3005
R623 VTAIL.n237 VTAIL.n236 9.3005
R624 VTAIL.n210 VTAIL.n209 9.3005
R625 VTAIL.n231 VTAIL.n230 9.3005
R626 VTAIL.n229 VTAIL.n228 9.3005
R627 VTAIL.n214 VTAIL.n213 9.3005
R628 VTAIL.n223 VTAIL.n222 9.3005
R629 VTAIL.n221 VTAIL.n220 9.3005
R630 VTAIL.n206 VTAIL.n205 9.3005
R631 VTAIL.n245 VTAIL.n244 9.3005
R632 VTAIL.n247 VTAIL.n246 9.3005
R633 VTAIL.n202 VTAIL.n201 9.3005
R634 VTAIL.n253 VTAIL.n252 9.3005
R635 VTAIL.n255 VTAIL.n254 9.3005
R636 VTAIL.n198 VTAIL.n197 9.3005
R637 VTAIL.n262 VTAIL.n261 9.3005
R638 VTAIL.n264 VTAIL.n263 9.3005
R639 VTAIL.n622 VTAIL.n621 9.3005
R640 VTAIL.n624 VTAIL.n623 9.3005
R641 VTAIL.n579 VTAIL.n578 9.3005
R642 VTAIL.n630 VTAIL.n629 9.3005
R643 VTAIL.n632 VTAIL.n631 9.3005
R644 VTAIL.n574 VTAIL.n573 9.3005
R645 VTAIL.n638 VTAIL.n637 9.3005
R646 VTAIL.n640 VTAIL.n639 9.3005
R647 VTAIL.n655 VTAIL.n654 9.3005
R648 VTAIL.n566 VTAIL.n565 9.3005
R649 VTAIL.n649 VTAIL.n648 9.3005
R650 VTAIL.n647 VTAIL.n646 9.3005
R651 VTAIL.n570 VTAIL.n569 9.3005
R652 VTAIL.n583 VTAIL.n582 9.3005
R653 VTAIL.n616 VTAIL.n615 9.3005
R654 VTAIL.n614 VTAIL.n613 9.3005
R655 VTAIL.n587 VTAIL.n586 9.3005
R656 VTAIL.n608 VTAIL.n607 9.3005
R657 VTAIL.n606 VTAIL.n605 9.3005
R658 VTAIL.n591 VTAIL.n590 9.3005
R659 VTAIL.n600 VTAIL.n599 9.3005
R660 VTAIL.n598 VTAIL.n597 9.3005
R661 VTAIL.n528 VTAIL.n527 9.3005
R662 VTAIL.n530 VTAIL.n529 9.3005
R663 VTAIL.n485 VTAIL.n484 9.3005
R664 VTAIL.n536 VTAIL.n535 9.3005
R665 VTAIL.n538 VTAIL.n537 9.3005
R666 VTAIL.n480 VTAIL.n479 9.3005
R667 VTAIL.n544 VTAIL.n543 9.3005
R668 VTAIL.n546 VTAIL.n545 9.3005
R669 VTAIL.n561 VTAIL.n560 9.3005
R670 VTAIL.n472 VTAIL.n471 9.3005
R671 VTAIL.n555 VTAIL.n554 9.3005
R672 VTAIL.n553 VTAIL.n552 9.3005
R673 VTAIL.n476 VTAIL.n475 9.3005
R674 VTAIL.n489 VTAIL.n488 9.3005
R675 VTAIL.n522 VTAIL.n521 9.3005
R676 VTAIL.n520 VTAIL.n519 9.3005
R677 VTAIL.n493 VTAIL.n492 9.3005
R678 VTAIL.n514 VTAIL.n513 9.3005
R679 VTAIL.n512 VTAIL.n511 9.3005
R680 VTAIL.n497 VTAIL.n496 9.3005
R681 VTAIL.n506 VTAIL.n505 9.3005
R682 VTAIL.n504 VTAIL.n503 9.3005
R683 VTAIL.n434 VTAIL.n433 9.3005
R684 VTAIL.n436 VTAIL.n435 9.3005
R685 VTAIL.n391 VTAIL.n390 9.3005
R686 VTAIL.n442 VTAIL.n441 9.3005
R687 VTAIL.n444 VTAIL.n443 9.3005
R688 VTAIL.n386 VTAIL.n385 9.3005
R689 VTAIL.n450 VTAIL.n449 9.3005
R690 VTAIL.n452 VTAIL.n451 9.3005
R691 VTAIL.n467 VTAIL.n466 9.3005
R692 VTAIL.n378 VTAIL.n377 9.3005
R693 VTAIL.n461 VTAIL.n460 9.3005
R694 VTAIL.n459 VTAIL.n458 9.3005
R695 VTAIL.n382 VTAIL.n381 9.3005
R696 VTAIL.n395 VTAIL.n394 9.3005
R697 VTAIL.n428 VTAIL.n427 9.3005
R698 VTAIL.n426 VTAIL.n425 9.3005
R699 VTAIL.n399 VTAIL.n398 9.3005
R700 VTAIL.n420 VTAIL.n419 9.3005
R701 VTAIL.n418 VTAIL.n417 9.3005
R702 VTAIL.n403 VTAIL.n402 9.3005
R703 VTAIL.n412 VTAIL.n411 9.3005
R704 VTAIL.n410 VTAIL.n409 9.3005
R705 VTAIL.n340 VTAIL.n339 9.3005
R706 VTAIL.n342 VTAIL.n341 9.3005
R707 VTAIL.n297 VTAIL.n296 9.3005
R708 VTAIL.n348 VTAIL.n347 9.3005
R709 VTAIL.n350 VTAIL.n349 9.3005
R710 VTAIL.n292 VTAIL.n291 9.3005
R711 VTAIL.n356 VTAIL.n355 9.3005
R712 VTAIL.n358 VTAIL.n357 9.3005
R713 VTAIL.n373 VTAIL.n372 9.3005
R714 VTAIL.n284 VTAIL.n283 9.3005
R715 VTAIL.n367 VTAIL.n366 9.3005
R716 VTAIL.n365 VTAIL.n364 9.3005
R717 VTAIL.n288 VTAIL.n287 9.3005
R718 VTAIL.n301 VTAIL.n300 9.3005
R719 VTAIL.n334 VTAIL.n333 9.3005
R720 VTAIL.n332 VTAIL.n331 9.3005
R721 VTAIL.n305 VTAIL.n304 9.3005
R722 VTAIL.n326 VTAIL.n325 9.3005
R723 VTAIL.n324 VTAIL.n323 9.3005
R724 VTAIL.n309 VTAIL.n308 9.3005
R725 VTAIL.n318 VTAIL.n317 9.3005
R726 VTAIL.n316 VTAIL.n315 9.3005
R727 VTAIL.n705 VTAIL.n680 8.92171
R728 VTAIL.n718 VTAIL.n672 8.92171
R729 VTAIL.n47 VTAIL.n22 8.92171
R730 VTAIL.n60 VTAIL.n14 8.92171
R731 VTAIL.n141 VTAIL.n116 8.92171
R732 VTAIL.n154 VTAIL.n108 8.92171
R733 VTAIL.n235 VTAIL.n210 8.92171
R734 VTAIL.n248 VTAIL.n202 8.92171
R735 VTAIL.n625 VTAIL.n579 8.92171
R736 VTAIL.n612 VTAIL.n587 8.92171
R737 VTAIL.n531 VTAIL.n485 8.92171
R738 VTAIL.n518 VTAIL.n493 8.92171
R739 VTAIL.n437 VTAIL.n391 8.92171
R740 VTAIL.n424 VTAIL.n399 8.92171
R741 VTAIL.n343 VTAIL.n297 8.92171
R742 VTAIL.n330 VTAIL.n305 8.92171
R743 VTAIL.n706 VTAIL.n678 8.14595
R744 VTAIL.n717 VTAIL.n674 8.14595
R745 VTAIL.n48 VTAIL.n20 8.14595
R746 VTAIL.n59 VTAIL.n16 8.14595
R747 VTAIL.n142 VTAIL.n114 8.14595
R748 VTAIL.n153 VTAIL.n110 8.14595
R749 VTAIL.n236 VTAIL.n208 8.14595
R750 VTAIL.n247 VTAIL.n204 8.14595
R751 VTAIL.n624 VTAIL.n581 8.14595
R752 VTAIL.n613 VTAIL.n585 8.14595
R753 VTAIL.n530 VTAIL.n487 8.14595
R754 VTAIL.n519 VTAIL.n491 8.14595
R755 VTAIL.n436 VTAIL.n393 8.14595
R756 VTAIL.n425 VTAIL.n397 8.14595
R757 VTAIL.n342 VTAIL.n299 8.14595
R758 VTAIL.n331 VTAIL.n303 8.14595
R759 VTAIL.n710 VTAIL.n709 7.3702
R760 VTAIL.n714 VTAIL.n713 7.3702
R761 VTAIL.n52 VTAIL.n51 7.3702
R762 VTAIL.n56 VTAIL.n55 7.3702
R763 VTAIL.n146 VTAIL.n145 7.3702
R764 VTAIL.n150 VTAIL.n149 7.3702
R765 VTAIL.n240 VTAIL.n239 7.3702
R766 VTAIL.n244 VTAIL.n243 7.3702
R767 VTAIL.n621 VTAIL.n620 7.3702
R768 VTAIL.n617 VTAIL.n616 7.3702
R769 VTAIL.n527 VTAIL.n526 7.3702
R770 VTAIL.n523 VTAIL.n522 7.3702
R771 VTAIL.n433 VTAIL.n432 7.3702
R772 VTAIL.n429 VTAIL.n428 7.3702
R773 VTAIL.n339 VTAIL.n338 7.3702
R774 VTAIL.n335 VTAIL.n334 7.3702
R775 VTAIL.n710 VTAIL.n676 6.59444
R776 VTAIL.n713 VTAIL.n676 6.59444
R777 VTAIL.n52 VTAIL.n18 6.59444
R778 VTAIL.n55 VTAIL.n18 6.59444
R779 VTAIL.n146 VTAIL.n112 6.59444
R780 VTAIL.n149 VTAIL.n112 6.59444
R781 VTAIL.n240 VTAIL.n206 6.59444
R782 VTAIL.n243 VTAIL.n206 6.59444
R783 VTAIL.n620 VTAIL.n583 6.59444
R784 VTAIL.n617 VTAIL.n583 6.59444
R785 VTAIL.n526 VTAIL.n489 6.59444
R786 VTAIL.n523 VTAIL.n489 6.59444
R787 VTAIL.n432 VTAIL.n395 6.59444
R788 VTAIL.n429 VTAIL.n395 6.59444
R789 VTAIL.n338 VTAIL.n301 6.59444
R790 VTAIL.n335 VTAIL.n301 6.59444
R791 VTAIL.n709 VTAIL.n678 5.81868
R792 VTAIL.n714 VTAIL.n674 5.81868
R793 VTAIL.n51 VTAIL.n20 5.81868
R794 VTAIL.n56 VTAIL.n16 5.81868
R795 VTAIL.n145 VTAIL.n114 5.81868
R796 VTAIL.n150 VTAIL.n110 5.81868
R797 VTAIL.n239 VTAIL.n208 5.81868
R798 VTAIL.n244 VTAIL.n204 5.81868
R799 VTAIL.n621 VTAIL.n581 5.81868
R800 VTAIL.n616 VTAIL.n585 5.81868
R801 VTAIL.n527 VTAIL.n487 5.81868
R802 VTAIL.n522 VTAIL.n491 5.81868
R803 VTAIL.n433 VTAIL.n393 5.81868
R804 VTAIL.n428 VTAIL.n397 5.81868
R805 VTAIL.n339 VTAIL.n299 5.81868
R806 VTAIL.n334 VTAIL.n303 5.81868
R807 VTAIL.n706 VTAIL.n705 5.04292
R808 VTAIL.n718 VTAIL.n717 5.04292
R809 VTAIL.n48 VTAIL.n47 5.04292
R810 VTAIL.n60 VTAIL.n59 5.04292
R811 VTAIL.n142 VTAIL.n141 5.04292
R812 VTAIL.n154 VTAIL.n153 5.04292
R813 VTAIL.n236 VTAIL.n235 5.04292
R814 VTAIL.n248 VTAIL.n247 5.04292
R815 VTAIL.n625 VTAIL.n624 5.04292
R816 VTAIL.n613 VTAIL.n612 5.04292
R817 VTAIL.n531 VTAIL.n530 5.04292
R818 VTAIL.n519 VTAIL.n518 5.04292
R819 VTAIL.n437 VTAIL.n436 5.04292
R820 VTAIL.n425 VTAIL.n424 5.04292
R821 VTAIL.n343 VTAIL.n342 5.04292
R822 VTAIL.n331 VTAIL.n330 5.04292
R823 VTAIL.n702 VTAIL.n680 4.26717
R824 VTAIL.n721 VTAIL.n672 4.26717
R825 VTAIL.n750 VTAIL.n658 4.26717
R826 VTAIL.n44 VTAIL.n22 4.26717
R827 VTAIL.n63 VTAIL.n14 4.26717
R828 VTAIL.n92 VTAIL.n0 4.26717
R829 VTAIL.n138 VTAIL.n116 4.26717
R830 VTAIL.n157 VTAIL.n108 4.26717
R831 VTAIL.n186 VTAIL.n94 4.26717
R832 VTAIL.n232 VTAIL.n210 4.26717
R833 VTAIL.n251 VTAIL.n202 4.26717
R834 VTAIL.n280 VTAIL.n188 4.26717
R835 VTAIL.n656 VTAIL.n564 4.26717
R836 VTAIL.n628 VTAIL.n579 4.26717
R837 VTAIL.n609 VTAIL.n587 4.26717
R838 VTAIL.n562 VTAIL.n470 4.26717
R839 VTAIL.n534 VTAIL.n485 4.26717
R840 VTAIL.n515 VTAIL.n493 4.26717
R841 VTAIL.n468 VTAIL.n376 4.26717
R842 VTAIL.n440 VTAIL.n391 4.26717
R843 VTAIL.n421 VTAIL.n399 4.26717
R844 VTAIL.n374 VTAIL.n282 4.26717
R845 VTAIL.n346 VTAIL.n297 4.26717
R846 VTAIL.n327 VTAIL.n305 4.26717
R847 VTAIL.n691 VTAIL.n687 3.70982
R848 VTAIL.n33 VTAIL.n29 3.70982
R849 VTAIL.n127 VTAIL.n123 3.70982
R850 VTAIL.n221 VTAIL.n217 3.70982
R851 VTAIL.n598 VTAIL.n594 3.70982
R852 VTAIL.n504 VTAIL.n500 3.70982
R853 VTAIL.n410 VTAIL.n406 3.70982
R854 VTAIL.n316 VTAIL.n312 3.70982
R855 VTAIL.n701 VTAIL.n682 3.49141
R856 VTAIL.n722 VTAIL.n670 3.49141
R857 VTAIL.n748 VTAIL.n747 3.49141
R858 VTAIL.n43 VTAIL.n24 3.49141
R859 VTAIL.n64 VTAIL.n12 3.49141
R860 VTAIL.n90 VTAIL.n89 3.49141
R861 VTAIL.n137 VTAIL.n118 3.49141
R862 VTAIL.n158 VTAIL.n106 3.49141
R863 VTAIL.n184 VTAIL.n183 3.49141
R864 VTAIL.n231 VTAIL.n212 3.49141
R865 VTAIL.n252 VTAIL.n200 3.49141
R866 VTAIL.n278 VTAIL.n277 3.49141
R867 VTAIL.n654 VTAIL.n653 3.49141
R868 VTAIL.n629 VTAIL.n577 3.49141
R869 VTAIL.n608 VTAIL.n589 3.49141
R870 VTAIL.n560 VTAIL.n559 3.49141
R871 VTAIL.n535 VTAIL.n483 3.49141
R872 VTAIL.n514 VTAIL.n495 3.49141
R873 VTAIL.n466 VTAIL.n465 3.49141
R874 VTAIL.n441 VTAIL.n389 3.49141
R875 VTAIL.n420 VTAIL.n401 3.49141
R876 VTAIL.n372 VTAIL.n371 3.49141
R877 VTAIL.n347 VTAIL.n295 3.49141
R878 VTAIL.n326 VTAIL.n307 3.49141
R879 VTAIL.n698 VTAIL.n697 2.71565
R880 VTAIL.n726 VTAIL.n725 2.71565
R881 VTAIL.n744 VTAIL.n660 2.71565
R882 VTAIL.n40 VTAIL.n39 2.71565
R883 VTAIL.n68 VTAIL.n67 2.71565
R884 VTAIL.n86 VTAIL.n2 2.71565
R885 VTAIL.n134 VTAIL.n133 2.71565
R886 VTAIL.n162 VTAIL.n161 2.71565
R887 VTAIL.n180 VTAIL.n96 2.71565
R888 VTAIL.n228 VTAIL.n227 2.71565
R889 VTAIL.n256 VTAIL.n255 2.71565
R890 VTAIL.n274 VTAIL.n190 2.71565
R891 VTAIL.n650 VTAIL.n566 2.71565
R892 VTAIL.n633 VTAIL.n632 2.71565
R893 VTAIL.n605 VTAIL.n604 2.71565
R894 VTAIL.n556 VTAIL.n472 2.71565
R895 VTAIL.n539 VTAIL.n538 2.71565
R896 VTAIL.n511 VTAIL.n510 2.71565
R897 VTAIL.n462 VTAIL.n378 2.71565
R898 VTAIL.n445 VTAIL.n444 2.71565
R899 VTAIL.n417 VTAIL.n416 2.71565
R900 VTAIL.n368 VTAIL.n284 2.71565
R901 VTAIL.n351 VTAIL.n350 2.71565
R902 VTAIL.n323 VTAIL.n322 2.71565
R903 VTAIL.n694 VTAIL.n684 1.93989
R904 VTAIL.n730 VTAIL.n668 1.93989
R905 VTAIL.n743 VTAIL.n662 1.93989
R906 VTAIL.n36 VTAIL.n26 1.93989
R907 VTAIL.n72 VTAIL.n10 1.93989
R908 VTAIL.n85 VTAIL.n4 1.93989
R909 VTAIL.n130 VTAIL.n120 1.93989
R910 VTAIL.n166 VTAIL.n104 1.93989
R911 VTAIL.n179 VTAIL.n98 1.93989
R912 VTAIL.n224 VTAIL.n214 1.93989
R913 VTAIL.n260 VTAIL.n198 1.93989
R914 VTAIL.n273 VTAIL.n192 1.93989
R915 VTAIL.n649 VTAIL.n568 1.93989
R916 VTAIL.n636 VTAIL.n574 1.93989
R917 VTAIL.n601 VTAIL.n591 1.93989
R918 VTAIL.n555 VTAIL.n474 1.93989
R919 VTAIL.n542 VTAIL.n480 1.93989
R920 VTAIL.n507 VTAIL.n497 1.93989
R921 VTAIL.n461 VTAIL.n380 1.93989
R922 VTAIL.n448 VTAIL.n386 1.93989
R923 VTAIL.n413 VTAIL.n403 1.93989
R924 VTAIL.n367 VTAIL.n286 1.93989
R925 VTAIL.n354 VTAIL.n292 1.93989
R926 VTAIL.n319 VTAIL.n309 1.93989
R927 VTAIL.n693 VTAIL.n686 1.16414
R928 VTAIL.n731 VTAIL.n666 1.16414
R929 VTAIL.n740 VTAIL.n739 1.16414
R930 VTAIL.n35 VTAIL.n28 1.16414
R931 VTAIL.n73 VTAIL.n8 1.16414
R932 VTAIL.n82 VTAIL.n81 1.16414
R933 VTAIL.n129 VTAIL.n122 1.16414
R934 VTAIL.n167 VTAIL.n102 1.16414
R935 VTAIL.n176 VTAIL.n175 1.16414
R936 VTAIL.n223 VTAIL.n216 1.16414
R937 VTAIL.n261 VTAIL.n196 1.16414
R938 VTAIL.n270 VTAIL.n269 1.16414
R939 VTAIL.n646 VTAIL.n645 1.16414
R940 VTAIL.n637 VTAIL.n572 1.16414
R941 VTAIL.n600 VTAIL.n593 1.16414
R942 VTAIL.n552 VTAIL.n551 1.16414
R943 VTAIL.n543 VTAIL.n478 1.16414
R944 VTAIL.n506 VTAIL.n499 1.16414
R945 VTAIL.n458 VTAIL.n457 1.16414
R946 VTAIL.n449 VTAIL.n384 1.16414
R947 VTAIL.n412 VTAIL.n405 1.16414
R948 VTAIL.n364 VTAIL.n363 1.16414
R949 VTAIL.n355 VTAIL.n290 1.16414
R950 VTAIL.n318 VTAIL.n311 1.16414
R951 VTAIL.n469 VTAIL.n375 1.02636
R952 VTAIL.n657 VTAIL.n563 1.02636
R953 VTAIL.n281 VTAIL.n187 1.02636
R954 VTAIL VTAIL.n93 0.571621
R955 VTAIL.n563 VTAIL.n469 0.470328
R956 VTAIL.n187 VTAIL.n93 0.470328
R957 VTAIL VTAIL.n751 0.455241
R958 VTAIL.n690 VTAIL.n689 0.388379
R959 VTAIL.n735 VTAIL.n734 0.388379
R960 VTAIL.n736 VTAIL.n664 0.388379
R961 VTAIL.n32 VTAIL.n31 0.388379
R962 VTAIL.n77 VTAIL.n76 0.388379
R963 VTAIL.n78 VTAIL.n6 0.388379
R964 VTAIL.n126 VTAIL.n125 0.388379
R965 VTAIL.n171 VTAIL.n170 0.388379
R966 VTAIL.n172 VTAIL.n100 0.388379
R967 VTAIL.n220 VTAIL.n219 0.388379
R968 VTAIL.n265 VTAIL.n264 0.388379
R969 VTAIL.n266 VTAIL.n194 0.388379
R970 VTAIL.n642 VTAIL.n570 0.388379
R971 VTAIL.n641 VTAIL.n640 0.388379
R972 VTAIL.n597 VTAIL.n596 0.388379
R973 VTAIL.n548 VTAIL.n476 0.388379
R974 VTAIL.n547 VTAIL.n546 0.388379
R975 VTAIL.n503 VTAIL.n502 0.388379
R976 VTAIL.n454 VTAIL.n382 0.388379
R977 VTAIL.n453 VTAIL.n452 0.388379
R978 VTAIL.n409 VTAIL.n408 0.388379
R979 VTAIL.n360 VTAIL.n288 0.388379
R980 VTAIL.n359 VTAIL.n358 0.388379
R981 VTAIL.n315 VTAIL.n314 0.388379
R982 VTAIL.n692 VTAIL.n691 0.155672
R983 VTAIL.n692 VTAIL.n683 0.155672
R984 VTAIL.n699 VTAIL.n683 0.155672
R985 VTAIL.n700 VTAIL.n699 0.155672
R986 VTAIL.n700 VTAIL.n679 0.155672
R987 VTAIL.n707 VTAIL.n679 0.155672
R988 VTAIL.n708 VTAIL.n707 0.155672
R989 VTAIL.n708 VTAIL.n675 0.155672
R990 VTAIL.n715 VTAIL.n675 0.155672
R991 VTAIL.n716 VTAIL.n715 0.155672
R992 VTAIL.n716 VTAIL.n671 0.155672
R993 VTAIL.n723 VTAIL.n671 0.155672
R994 VTAIL.n724 VTAIL.n723 0.155672
R995 VTAIL.n724 VTAIL.n667 0.155672
R996 VTAIL.n732 VTAIL.n667 0.155672
R997 VTAIL.n733 VTAIL.n732 0.155672
R998 VTAIL.n733 VTAIL.n663 0.155672
R999 VTAIL.n741 VTAIL.n663 0.155672
R1000 VTAIL.n742 VTAIL.n741 0.155672
R1001 VTAIL.n742 VTAIL.n659 0.155672
R1002 VTAIL.n749 VTAIL.n659 0.155672
R1003 VTAIL.n34 VTAIL.n33 0.155672
R1004 VTAIL.n34 VTAIL.n25 0.155672
R1005 VTAIL.n41 VTAIL.n25 0.155672
R1006 VTAIL.n42 VTAIL.n41 0.155672
R1007 VTAIL.n42 VTAIL.n21 0.155672
R1008 VTAIL.n49 VTAIL.n21 0.155672
R1009 VTAIL.n50 VTAIL.n49 0.155672
R1010 VTAIL.n50 VTAIL.n17 0.155672
R1011 VTAIL.n57 VTAIL.n17 0.155672
R1012 VTAIL.n58 VTAIL.n57 0.155672
R1013 VTAIL.n58 VTAIL.n13 0.155672
R1014 VTAIL.n65 VTAIL.n13 0.155672
R1015 VTAIL.n66 VTAIL.n65 0.155672
R1016 VTAIL.n66 VTAIL.n9 0.155672
R1017 VTAIL.n74 VTAIL.n9 0.155672
R1018 VTAIL.n75 VTAIL.n74 0.155672
R1019 VTAIL.n75 VTAIL.n5 0.155672
R1020 VTAIL.n83 VTAIL.n5 0.155672
R1021 VTAIL.n84 VTAIL.n83 0.155672
R1022 VTAIL.n84 VTAIL.n1 0.155672
R1023 VTAIL.n91 VTAIL.n1 0.155672
R1024 VTAIL.n128 VTAIL.n127 0.155672
R1025 VTAIL.n128 VTAIL.n119 0.155672
R1026 VTAIL.n135 VTAIL.n119 0.155672
R1027 VTAIL.n136 VTAIL.n135 0.155672
R1028 VTAIL.n136 VTAIL.n115 0.155672
R1029 VTAIL.n143 VTAIL.n115 0.155672
R1030 VTAIL.n144 VTAIL.n143 0.155672
R1031 VTAIL.n144 VTAIL.n111 0.155672
R1032 VTAIL.n151 VTAIL.n111 0.155672
R1033 VTAIL.n152 VTAIL.n151 0.155672
R1034 VTAIL.n152 VTAIL.n107 0.155672
R1035 VTAIL.n159 VTAIL.n107 0.155672
R1036 VTAIL.n160 VTAIL.n159 0.155672
R1037 VTAIL.n160 VTAIL.n103 0.155672
R1038 VTAIL.n168 VTAIL.n103 0.155672
R1039 VTAIL.n169 VTAIL.n168 0.155672
R1040 VTAIL.n169 VTAIL.n99 0.155672
R1041 VTAIL.n177 VTAIL.n99 0.155672
R1042 VTAIL.n178 VTAIL.n177 0.155672
R1043 VTAIL.n178 VTAIL.n95 0.155672
R1044 VTAIL.n185 VTAIL.n95 0.155672
R1045 VTAIL.n222 VTAIL.n221 0.155672
R1046 VTAIL.n222 VTAIL.n213 0.155672
R1047 VTAIL.n229 VTAIL.n213 0.155672
R1048 VTAIL.n230 VTAIL.n229 0.155672
R1049 VTAIL.n230 VTAIL.n209 0.155672
R1050 VTAIL.n237 VTAIL.n209 0.155672
R1051 VTAIL.n238 VTAIL.n237 0.155672
R1052 VTAIL.n238 VTAIL.n205 0.155672
R1053 VTAIL.n245 VTAIL.n205 0.155672
R1054 VTAIL.n246 VTAIL.n245 0.155672
R1055 VTAIL.n246 VTAIL.n201 0.155672
R1056 VTAIL.n253 VTAIL.n201 0.155672
R1057 VTAIL.n254 VTAIL.n253 0.155672
R1058 VTAIL.n254 VTAIL.n197 0.155672
R1059 VTAIL.n262 VTAIL.n197 0.155672
R1060 VTAIL.n263 VTAIL.n262 0.155672
R1061 VTAIL.n263 VTAIL.n193 0.155672
R1062 VTAIL.n271 VTAIL.n193 0.155672
R1063 VTAIL.n272 VTAIL.n271 0.155672
R1064 VTAIL.n272 VTAIL.n189 0.155672
R1065 VTAIL.n279 VTAIL.n189 0.155672
R1066 VTAIL.n655 VTAIL.n565 0.155672
R1067 VTAIL.n648 VTAIL.n565 0.155672
R1068 VTAIL.n648 VTAIL.n647 0.155672
R1069 VTAIL.n647 VTAIL.n569 0.155672
R1070 VTAIL.n639 VTAIL.n569 0.155672
R1071 VTAIL.n639 VTAIL.n638 0.155672
R1072 VTAIL.n638 VTAIL.n573 0.155672
R1073 VTAIL.n631 VTAIL.n573 0.155672
R1074 VTAIL.n631 VTAIL.n630 0.155672
R1075 VTAIL.n630 VTAIL.n578 0.155672
R1076 VTAIL.n623 VTAIL.n578 0.155672
R1077 VTAIL.n623 VTAIL.n622 0.155672
R1078 VTAIL.n622 VTAIL.n582 0.155672
R1079 VTAIL.n615 VTAIL.n582 0.155672
R1080 VTAIL.n615 VTAIL.n614 0.155672
R1081 VTAIL.n614 VTAIL.n586 0.155672
R1082 VTAIL.n607 VTAIL.n586 0.155672
R1083 VTAIL.n607 VTAIL.n606 0.155672
R1084 VTAIL.n606 VTAIL.n590 0.155672
R1085 VTAIL.n599 VTAIL.n590 0.155672
R1086 VTAIL.n599 VTAIL.n598 0.155672
R1087 VTAIL.n561 VTAIL.n471 0.155672
R1088 VTAIL.n554 VTAIL.n471 0.155672
R1089 VTAIL.n554 VTAIL.n553 0.155672
R1090 VTAIL.n553 VTAIL.n475 0.155672
R1091 VTAIL.n545 VTAIL.n475 0.155672
R1092 VTAIL.n545 VTAIL.n544 0.155672
R1093 VTAIL.n544 VTAIL.n479 0.155672
R1094 VTAIL.n537 VTAIL.n479 0.155672
R1095 VTAIL.n537 VTAIL.n536 0.155672
R1096 VTAIL.n536 VTAIL.n484 0.155672
R1097 VTAIL.n529 VTAIL.n484 0.155672
R1098 VTAIL.n529 VTAIL.n528 0.155672
R1099 VTAIL.n528 VTAIL.n488 0.155672
R1100 VTAIL.n521 VTAIL.n488 0.155672
R1101 VTAIL.n521 VTAIL.n520 0.155672
R1102 VTAIL.n520 VTAIL.n492 0.155672
R1103 VTAIL.n513 VTAIL.n492 0.155672
R1104 VTAIL.n513 VTAIL.n512 0.155672
R1105 VTAIL.n512 VTAIL.n496 0.155672
R1106 VTAIL.n505 VTAIL.n496 0.155672
R1107 VTAIL.n505 VTAIL.n504 0.155672
R1108 VTAIL.n467 VTAIL.n377 0.155672
R1109 VTAIL.n460 VTAIL.n377 0.155672
R1110 VTAIL.n460 VTAIL.n459 0.155672
R1111 VTAIL.n459 VTAIL.n381 0.155672
R1112 VTAIL.n451 VTAIL.n381 0.155672
R1113 VTAIL.n451 VTAIL.n450 0.155672
R1114 VTAIL.n450 VTAIL.n385 0.155672
R1115 VTAIL.n443 VTAIL.n385 0.155672
R1116 VTAIL.n443 VTAIL.n442 0.155672
R1117 VTAIL.n442 VTAIL.n390 0.155672
R1118 VTAIL.n435 VTAIL.n390 0.155672
R1119 VTAIL.n435 VTAIL.n434 0.155672
R1120 VTAIL.n434 VTAIL.n394 0.155672
R1121 VTAIL.n427 VTAIL.n394 0.155672
R1122 VTAIL.n427 VTAIL.n426 0.155672
R1123 VTAIL.n426 VTAIL.n398 0.155672
R1124 VTAIL.n419 VTAIL.n398 0.155672
R1125 VTAIL.n419 VTAIL.n418 0.155672
R1126 VTAIL.n418 VTAIL.n402 0.155672
R1127 VTAIL.n411 VTAIL.n402 0.155672
R1128 VTAIL.n411 VTAIL.n410 0.155672
R1129 VTAIL.n373 VTAIL.n283 0.155672
R1130 VTAIL.n366 VTAIL.n283 0.155672
R1131 VTAIL.n366 VTAIL.n365 0.155672
R1132 VTAIL.n365 VTAIL.n287 0.155672
R1133 VTAIL.n357 VTAIL.n287 0.155672
R1134 VTAIL.n357 VTAIL.n356 0.155672
R1135 VTAIL.n356 VTAIL.n291 0.155672
R1136 VTAIL.n349 VTAIL.n291 0.155672
R1137 VTAIL.n349 VTAIL.n348 0.155672
R1138 VTAIL.n348 VTAIL.n296 0.155672
R1139 VTAIL.n341 VTAIL.n296 0.155672
R1140 VTAIL.n341 VTAIL.n340 0.155672
R1141 VTAIL.n340 VTAIL.n300 0.155672
R1142 VTAIL.n333 VTAIL.n300 0.155672
R1143 VTAIL.n333 VTAIL.n332 0.155672
R1144 VTAIL.n332 VTAIL.n304 0.155672
R1145 VTAIL.n325 VTAIL.n304 0.155672
R1146 VTAIL.n325 VTAIL.n324 0.155672
R1147 VTAIL.n324 VTAIL.n308 0.155672
R1148 VTAIL.n317 VTAIL.n308 0.155672
R1149 VTAIL.n317 VTAIL.n316 0.155672
R1150 B.n128 B.t0 671.542
R1151 B.n288 B.t3 671.542
R1152 B.n46 B.t9 671.542
R1153 B.n40 B.t6 671.542
R1154 B.n376 B.n375 585
R1155 B.n374 B.n95 585
R1156 B.n373 B.n372 585
R1157 B.n371 B.n96 585
R1158 B.n370 B.n369 585
R1159 B.n368 B.n97 585
R1160 B.n367 B.n366 585
R1161 B.n365 B.n98 585
R1162 B.n364 B.n363 585
R1163 B.n362 B.n99 585
R1164 B.n361 B.n360 585
R1165 B.n359 B.n100 585
R1166 B.n358 B.n357 585
R1167 B.n356 B.n101 585
R1168 B.n355 B.n354 585
R1169 B.n353 B.n102 585
R1170 B.n352 B.n351 585
R1171 B.n350 B.n103 585
R1172 B.n349 B.n348 585
R1173 B.n347 B.n104 585
R1174 B.n346 B.n345 585
R1175 B.n344 B.n105 585
R1176 B.n343 B.n342 585
R1177 B.n341 B.n106 585
R1178 B.n340 B.n339 585
R1179 B.n338 B.n107 585
R1180 B.n337 B.n336 585
R1181 B.n335 B.n108 585
R1182 B.n334 B.n333 585
R1183 B.n332 B.n109 585
R1184 B.n331 B.n330 585
R1185 B.n329 B.n110 585
R1186 B.n328 B.n327 585
R1187 B.n326 B.n111 585
R1188 B.n325 B.n324 585
R1189 B.n323 B.n112 585
R1190 B.n322 B.n321 585
R1191 B.n320 B.n113 585
R1192 B.n319 B.n318 585
R1193 B.n317 B.n114 585
R1194 B.n316 B.n315 585
R1195 B.n314 B.n115 585
R1196 B.n313 B.n312 585
R1197 B.n311 B.n116 585
R1198 B.n310 B.n309 585
R1199 B.n308 B.n117 585
R1200 B.n307 B.n306 585
R1201 B.n305 B.n118 585
R1202 B.n304 B.n303 585
R1203 B.n302 B.n119 585
R1204 B.n301 B.n300 585
R1205 B.n299 B.n120 585
R1206 B.n298 B.n297 585
R1207 B.n296 B.n121 585
R1208 B.n295 B.n294 585
R1209 B.n293 B.n122 585
R1210 B.n292 B.n291 585
R1211 B.n287 B.n123 585
R1212 B.n286 B.n285 585
R1213 B.n284 B.n124 585
R1214 B.n283 B.n282 585
R1215 B.n281 B.n125 585
R1216 B.n280 B.n279 585
R1217 B.n278 B.n126 585
R1218 B.n277 B.n276 585
R1219 B.n274 B.n127 585
R1220 B.n273 B.n272 585
R1221 B.n271 B.n130 585
R1222 B.n270 B.n269 585
R1223 B.n268 B.n131 585
R1224 B.n267 B.n266 585
R1225 B.n265 B.n132 585
R1226 B.n264 B.n263 585
R1227 B.n262 B.n133 585
R1228 B.n261 B.n260 585
R1229 B.n259 B.n134 585
R1230 B.n258 B.n257 585
R1231 B.n256 B.n135 585
R1232 B.n255 B.n254 585
R1233 B.n253 B.n136 585
R1234 B.n252 B.n251 585
R1235 B.n250 B.n137 585
R1236 B.n249 B.n248 585
R1237 B.n247 B.n138 585
R1238 B.n246 B.n245 585
R1239 B.n244 B.n139 585
R1240 B.n243 B.n242 585
R1241 B.n241 B.n140 585
R1242 B.n240 B.n239 585
R1243 B.n238 B.n141 585
R1244 B.n237 B.n236 585
R1245 B.n235 B.n142 585
R1246 B.n234 B.n233 585
R1247 B.n232 B.n143 585
R1248 B.n231 B.n230 585
R1249 B.n229 B.n144 585
R1250 B.n228 B.n227 585
R1251 B.n226 B.n145 585
R1252 B.n225 B.n224 585
R1253 B.n223 B.n146 585
R1254 B.n222 B.n221 585
R1255 B.n220 B.n147 585
R1256 B.n219 B.n218 585
R1257 B.n217 B.n148 585
R1258 B.n216 B.n215 585
R1259 B.n214 B.n149 585
R1260 B.n213 B.n212 585
R1261 B.n211 B.n150 585
R1262 B.n210 B.n209 585
R1263 B.n208 B.n151 585
R1264 B.n207 B.n206 585
R1265 B.n205 B.n152 585
R1266 B.n204 B.n203 585
R1267 B.n202 B.n153 585
R1268 B.n201 B.n200 585
R1269 B.n199 B.n154 585
R1270 B.n198 B.n197 585
R1271 B.n196 B.n155 585
R1272 B.n195 B.n194 585
R1273 B.n193 B.n156 585
R1274 B.n192 B.n191 585
R1275 B.n377 B.n94 585
R1276 B.n379 B.n378 585
R1277 B.n380 B.n93 585
R1278 B.n382 B.n381 585
R1279 B.n383 B.n92 585
R1280 B.n385 B.n384 585
R1281 B.n386 B.n91 585
R1282 B.n388 B.n387 585
R1283 B.n389 B.n90 585
R1284 B.n391 B.n390 585
R1285 B.n392 B.n89 585
R1286 B.n394 B.n393 585
R1287 B.n395 B.n88 585
R1288 B.n397 B.n396 585
R1289 B.n398 B.n87 585
R1290 B.n400 B.n399 585
R1291 B.n401 B.n86 585
R1292 B.n403 B.n402 585
R1293 B.n404 B.n85 585
R1294 B.n406 B.n405 585
R1295 B.n407 B.n84 585
R1296 B.n409 B.n408 585
R1297 B.n410 B.n83 585
R1298 B.n412 B.n411 585
R1299 B.n413 B.n82 585
R1300 B.n415 B.n414 585
R1301 B.n416 B.n81 585
R1302 B.n418 B.n417 585
R1303 B.n419 B.n80 585
R1304 B.n421 B.n420 585
R1305 B.n422 B.n79 585
R1306 B.n424 B.n423 585
R1307 B.n425 B.n78 585
R1308 B.n427 B.n426 585
R1309 B.n428 B.n77 585
R1310 B.n430 B.n429 585
R1311 B.n431 B.n76 585
R1312 B.n433 B.n432 585
R1313 B.n616 B.n11 585
R1314 B.n615 B.n614 585
R1315 B.n613 B.n12 585
R1316 B.n612 B.n611 585
R1317 B.n610 B.n13 585
R1318 B.n609 B.n608 585
R1319 B.n607 B.n14 585
R1320 B.n606 B.n605 585
R1321 B.n604 B.n15 585
R1322 B.n603 B.n602 585
R1323 B.n601 B.n16 585
R1324 B.n600 B.n599 585
R1325 B.n598 B.n17 585
R1326 B.n597 B.n596 585
R1327 B.n595 B.n18 585
R1328 B.n594 B.n593 585
R1329 B.n592 B.n19 585
R1330 B.n591 B.n590 585
R1331 B.n589 B.n20 585
R1332 B.n588 B.n587 585
R1333 B.n586 B.n21 585
R1334 B.n585 B.n584 585
R1335 B.n583 B.n22 585
R1336 B.n582 B.n581 585
R1337 B.n580 B.n23 585
R1338 B.n579 B.n578 585
R1339 B.n577 B.n24 585
R1340 B.n576 B.n575 585
R1341 B.n574 B.n25 585
R1342 B.n573 B.n572 585
R1343 B.n571 B.n26 585
R1344 B.n570 B.n569 585
R1345 B.n568 B.n27 585
R1346 B.n567 B.n566 585
R1347 B.n565 B.n28 585
R1348 B.n564 B.n563 585
R1349 B.n562 B.n29 585
R1350 B.n561 B.n560 585
R1351 B.n559 B.n30 585
R1352 B.n558 B.n557 585
R1353 B.n556 B.n31 585
R1354 B.n555 B.n554 585
R1355 B.n553 B.n32 585
R1356 B.n552 B.n551 585
R1357 B.n550 B.n33 585
R1358 B.n549 B.n548 585
R1359 B.n547 B.n34 585
R1360 B.n546 B.n545 585
R1361 B.n544 B.n35 585
R1362 B.n543 B.n542 585
R1363 B.n541 B.n36 585
R1364 B.n540 B.n539 585
R1365 B.n538 B.n37 585
R1366 B.n537 B.n536 585
R1367 B.n535 B.n38 585
R1368 B.n534 B.n533 585
R1369 B.n531 B.n39 585
R1370 B.n530 B.n529 585
R1371 B.n528 B.n42 585
R1372 B.n527 B.n526 585
R1373 B.n525 B.n43 585
R1374 B.n524 B.n523 585
R1375 B.n522 B.n44 585
R1376 B.n521 B.n520 585
R1377 B.n519 B.n45 585
R1378 B.n517 B.n516 585
R1379 B.n515 B.n48 585
R1380 B.n514 B.n513 585
R1381 B.n512 B.n49 585
R1382 B.n511 B.n510 585
R1383 B.n509 B.n50 585
R1384 B.n508 B.n507 585
R1385 B.n506 B.n51 585
R1386 B.n505 B.n504 585
R1387 B.n503 B.n52 585
R1388 B.n502 B.n501 585
R1389 B.n500 B.n53 585
R1390 B.n499 B.n498 585
R1391 B.n497 B.n54 585
R1392 B.n496 B.n495 585
R1393 B.n494 B.n55 585
R1394 B.n493 B.n492 585
R1395 B.n491 B.n56 585
R1396 B.n490 B.n489 585
R1397 B.n488 B.n57 585
R1398 B.n487 B.n486 585
R1399 B.n485 B.n58 585
R1400 B.n484 B.n483 585
R1401 B.n482 B.n59 585
R1402 B.n481 B.n480 585
R1403 B.n479 B.n60 585
R1404 B.n478 B.n477 585
R1405 B.n476 B.n61 585
R1406 B.n475 B.n474 585
R1407 B.n473 B.n62 585
R1408 B.n472 B.n471 585
R1409 B.n470 B.n63 585
R1410 B.n469 B.n468 585
R1411 B.n467 B.n64 585
R1412 B.n466 B.n465 585
R1413 B.n464 B.n65 585
R1414 B.n463 B.n462 585
R1415 B.n461 B.n66 585
R1416 B.n460 B.n459 585
R1417 B.n458 B.n67 585
R1418 B.n457 B.n456 585
R1419 B.n455 B.n68 585
R1420 B.n454 B.n453 585
R1421 B.n452 B.n69 585
R1422 B.n451 B.n450 585
R1423 B.n449 B.n70 585
R1424 B.n448 B.n447 585
R1425 B.n446 B.n71 585
R1426 B.n445 B.n444 585
R1427 B.n443 B.n72 585
R1428 B.n442 B.n441 585
R1429 B.n440 B.n73 585
R1430 B.n439 B.n438 585
R1431 B.n437 B.n74 585
R1432 B.n436 B.n435 585
R1433 B.n434 B.n75 585
R1434 B.n618 B.n617 585
R1435 B.n619 B.n10 585
R1436 B.n621 B.n620 585
R1437 B.n622 B.n9 585
R1438 B.n624 B.n623 585
R1439 B.n625 B.n8 585
R1440 B.n627 B.n626 585
R1441 B.n628 B.n7 585
R1442 B.n630 B.n629 585
R1443 B.n631 B.n6 585
R1444 B.n633 B.n632 585
R1445 B.n634 B.n5 585
R1446 B.n636 B.n635 585
R1447 B.n637 B.n4 585
R1448 B.n639 B.n638 585
R1449 B.n640 B.n3 585
R1450 B.n642 B.n641 585
R1451 B.n643 B.n0 585
R1452 B.n2 B.n1 585
R1453 B.n166 B.n165 585
R1454 B.n168 B.n167 585
R1455 B.n169 B.n164 585
R1456 B.n171 B.n170 585
R1457 B.n172 B.n163 585
R1458 B.n174 B.n173 585
R1459 B.n175 B.n162 585
R1460 B.n177 B.n176 585
R1461 B.n178 B.n161 585
R1462 B.n180 B.n179 585
R1463 B.n181 B.n160 585
R1464 B.n183 B.n182 585
R1465 B.n184 B.n159 585
R1466 B.n186 B.n185 585
R1467 B.n187 B.n158 585
R1468 B.n189 B.n188 585
R1469 B.n190 B.n157 585
R1470 B.n192 B.n157 502.111
R1471 B.n377 B.n376 502.111
R1472 B.n432 B.n75 502.111
R1473 B.n618 B.n11 502.111
R1474 B.n288 B.t4 484.344
R1475 B.n46 B.t11 484.344
R1476 B.n128 B.t1 484.344
R1477 B.n40 B.t8 484.344
R1478 B.n289 B.t5 461.264
R1479 B.n47 B.t10 461.264
R1480 B.n129 B.t2 461.264
R1481 B.n41 B.t7 461.264
R1482 B.n645 B.n644 256.663
R1483 B.n644 B.n643 235.042
R1484 B.n644 B.n2 235.042
R1485 B.n193 B.n192 163.367
R1486 B.n194 B.n193 163.367
R1487 B.n194 B.n155 163.367
R1488 B.n198 B.n155 163.367
R1489 B.n199 B.n198 163.367
R1490 B.n200 B.n199 163.367
R1491 B.n200 B.n153 163.367
R1492 B.n204 B.n153 163.367
R1493 B.n205 B.n204 163.367
R1494 B.n206 B.n205 163.367
R1495 B.n206 B.n151 163.367
R1496 B.n210 B.n151 163.367
R1497 B.n211 B.n210 163.367
R1498 B.n212 B.n211 163.367
R1499 B.n212 B.n149 163.367
R1500 B.n216 B.n149 163.367
R1501 B.n217 B.n216 163.367
R1502 B.n218 B.n217 163.367
R1503 B.n218 B.n147 163.367
R1504 B.n222 B.n147 163.367
R1505 B.n223 B.n222 163.367
R1506 B.n224 B.n223 163.367
R1507 B.n224 B.n145 163.367
R1508 B.n228 B.n145 163.367
R1509 B.n229 B.n228 163.367
R1510 B.n230 B.n229 163.367
R1511 B.n230 B.n143 163.367
R1512 B.n234 B.n143 163.367
R1513 B.n235 B.n234 163.367
R1514 B.n236 B.n235 163.367
R1515 B.n236 B.n141 163.367
R1516 B.n240 B.n141 163.367
R1517 B.n241 B.n240 163.367
R1518 B.n242 B.n241 163.367
R1519 B.n242 B.n139 163.367
R1520 B.n246 B.n139 163.367
R1521 B.n247 B.n246 163.367
R1522 B.n248 B.n247 163.367
R1523 B.n248 B.n137 163.367
R1524 B.n252 B.n137 163.367
R1525 B.n253 B.n252 163.367
R1526 B.n254 B.n253 163.367
R1527 B.n254 B.n135 163.367
R1528 B.n258 B.n135 163.367
R1529 B.n259 B.n258 163.367
R1530 B.n260 B.n259 163.367
R1531 B.n260 B.n133 163.367
R1532 B.n264 B.n133 163.367
R1533 B.n265 B.n264 163.367
R1534 B.n266 B.n265 163.367
R1535 B.n266 B.n131 163.367
R1536 B.n270 B.n131 163.367
R1537 B.n271 B.n270 163.367
R1538 B.n272 B.n271 163.367
R1539 B.n272 B.n127 163.367
R1540 B.n277 B.n127 163.367
R1541 B.n278 B.n277 163.367
R1542 B.n279 B.n278 163.367
R1543 B.n279 B.n125 163.367
R1544 B.n283 B.n125 163.367
R1545 B.n284 B.n283 163.367
R1546 B.n285 B.n284 163.367
R1547 B.n285 B.n123 163.367
R1548 B.n292 B.n123 163.367
R1549 B.n293 B.n292 163.367
R1550 B.n294 B.n293 163.367
R1551 B.n294 B.n121 163.367
R1552 B.n298 B.n121 163.367
R1553 B.n299 B.n298 163.367
R1554 B.n300 B.n299 163.367
R1555 B.n300 B.n119 163.367
R1556 B.n304 B.n119 163.367
R1557 B.n305 B.n304 163.367
R1558 B.n306 B.n305 163.367
R1559 B.n306 B.n117 163.367
R1560 B.n310 B.n117 163.367
R1561 B.n311 B.n310 163.367
R1562 B.n312 B.n311 163.367
R1563 B.n312 B.n115 163.367
R1564 B.n316 B.n115 163.367
R1565 B.n317 B.n316 163.367
R1566 B.n318 B.n317 163.367
R1567 B.n318 B.n113 163.367
R1568 B.n322 B.n113 163.367
R1569 B.n323 B.n322 163.367
R1570 B.n324 B.n323 163.367
R1571 B.n324 B.n111 163.367
R1572 B.n328 B.n111 163.367
R1573 B.n329 B.n328 163.367
R1574 B.n330 B.n329 163.367
R1575 B.n330 B.n109 163.367
R1576 B.n334 B.n109 163.367
R1577 B.n335 B.n334 163.367
R1578 B.n336 B.n335 163.367
R1579 B.n336 B.n107 163.367
R1580 B.n340 B.n107 163.367
R1581 B.n341 B.n340 163.367
R1582 B.n342 B.n341 163.367
R1583 B.n342 B.n105 163.367
R1584 B.n346 B.n105 163.367
R1585 B.n347 B.n346 163.367
R1586 B.n348 B.n347 163.367
R1587 B.n348 B.n103 163.367
R1588 B.n352 B.n103 163.367
R1589 B.n353 B.n352 163.367
R1590 B.n354 B.n353 163.367
R1591 B.n354 B.n101 163.367
R1592 B.n358 B.n101 163.367
R1593 B.n359 B.n358 163.367
R1594 B.n360 B.n359 163.367
R1595 B.n360 B.n99 163.367
R1596 B.n364 B.n99 163.367
R1597 B.n365 B.n364 163.367
R1598 B.n366 B.n365 163.367
R1599 B.n366 B.n97 163.367
R1600 B.n370 B.n97 163.367
R1601 B.n371 B.n370 163.367
R1602 B.n372 B.n371 163.367
R1603 B.n372 B.n95 163.367
R1604 B.n376 B.n95 163.367
R1605 B.n432 B.n431 163.367
R1606 B.n431 B.n430 163.367
R1607 B.n430 B.n77 163.367
R1608 B.n426 B.n77 163.367
R1609 B.n426 B.n425 163.367
R1610 B.n425 B.n424 163.367
R1611 B.n424 B.n79 163.367
R1612 B.n420 B.n79 163.367
R1613 B.n420 B.n419 163.367
R1614 B.n419 B.n418 163.367
R1615 B.n418 B.n81 163.367
R1616 B.n414 B.n81 163.367
R1617 B.n414 B.n413 163.367
R1618 B.n413 B.n412 163.367
R1619 B.n412 B.n83 163.367
R1620 B.n408 B.n83 163.367
R1621 B.n408 B.n407 163.367
R1622 B.n407 B.n406 163.367
R1623 B.n406 B.n85 163.367
R1624 B.n402 B.n85 163.367
R1625 B.n402 B.n401 163.367
R1626 B.n401 B.n400 163.367
R1627 B.n400 B.n87 163.367
R1628 B.n396 B.n87 163.367
R1629 B.n396 B.n395 163.367
R1630 B.n395 B.n394 163.367
R1631 B.n394 B.n89 163.367
R1632 B.n390 B.n89 163.367
R1633 B.n390 B.n389 163.367
R1634 B.n389 B.n388 163.367
R1635 B.n388 B.n91 163.367
R1636 B.n384 B.n91 163.367
R1637 B.n384 B.n383 163.367
R1638 B.n383 B.n382 163.367
R1639 B.n382 B.n93 163.367
R1640 B.n378 B.n93 163.367
R1641 B.n378 B.n377 163.367
R1642 B.n614 B.n11 163.367
R1643 B.n614 B.n613 163.367
R1644 B.n613 B.n612 163.367
R1645 B.n612 B.n13 163.367
R1646 B.n608 B.n13 163.367
R1647 B.n608 B.n607 163.367
R1648 B.n607 B.n606 163.367
R1649 B.n606 B.n15 163.367
R1650 B.n602 B.n15 163.367
R1651 B.n602 B.n601 163.367
R1652 B.n601 B.n600 163.367
R1653 B.n600 B.n17 163.367
R1654 B.n596 B.n17 163.367
R1655 B.n596 B.n595 163.367
R1656 B.n595 B.n594 163.367
R1657 B.n594 B.n19 163.367
R1658 B.n590 B.n19 163.367
R1659 B.n590 B.n589 163.367
R1660 B.n589 B.n588 163.367
R1661 B.n588 B.n21 163.367
R1662 B.n584 B.n21 163.367
R1663 B.n584 B.n583 163.367
R1664 B.n583 B.n582 163.367
R1665 B.n582 B.n23 163.367
R1666 B.n578 B.n23 163.367
R1667 B.n578 B.n577 163.367
R1668 B.n577 B.n576 163.367
R1669 B.n576 B.n25 163.367
R1670 B.n572 B.n25 163.367
R1671 B.n572 B.n571 163.367
R1672 B.n571 B.n570 163.367
R1673 B.n570 B.n27 163.367
R1674 B.n566 B.n27 163.367
R1675 B.n566 B.n565 163.367
R1676 B.n565 B.n564 163.367
R1677 B.n564 B.n29 163.367
R1678 B.n560 B.n29 163.367
R1679 B.n560 B.n559 163.367
R1680 B.n559 B.n558 163.367
R1681 B.n558 B.n31 163.367
R1682 B.n554 B.n31 163.367
R1683 B.n554 B.n553 163.367
R1684 B.n553 B.n552 163.367
R1685 B.n552 B.n33 163.367
R1686 B.n548 B.n33 163.367
R1687 B.n548 B.n547 163.367
R1688 B.n547 B.n546 163.367
R1689 B.n546 B.n35 163.367
R1690 B.n542 B.n35 163.367
R1691 B.n542 B.n541 163.367
R1692 B.n541 B.n540 163.367
R1693 B.n540 B.n37 163.367
R1694 B.n536 B.n37 163.367
R1695 B.n536 B.n535 163.367
R1696 B.n535 B.n534 163.367
R1697 B.n534 B.n39 163.367
R1698 B.n529 B.n39 163.367
R1699 B.n529 B.n528 163.367
R1700 B.n528 B.n527 163.367
R1701 B.n527 B.n43 163.367
R1702 B.n523 B.n43 163.367
R1703 B.n523 B.n522 163.367
R1704 B.n522 B.n521 163.367
R1705 B.n521 B.n45 163.367
R1706 B.n516 B.n45 163.367
R1707 B.n516 B.n515 163.367
R1708 B.n515 B.n514 163.367
R1709 B.n514 B.n49 163.367
R1710 B.n510 B.n49 163.367
R1711 B.n510 B.n509 163.367
R1712 B.n509 B.n508 163.367
R1713 B.n508 B.n51 163.367
R1714 B.n504 B.n51 163.367
R1715 B.n504 B.n503 163.367
R1716 B.n503 B.n502 163.367
R1717 B.n502 B.n53 163.367
R1718 B.n498 B.n53 163.367
R1719 B.n498 B.n497 163.367
R1720 B.n497 B.n496 163.367
R1721 B.n496 B.n55 163.367
R1722 B.n492 B.n55 163.367
R1723 B.n492 B.n491 163.367
R1724 B.n491 B.n490 163.367
R1725 B.n490 B.n57 163.367
R1726 B.n486 B.n57 163.367
R1727 B.n486 B.n485 163.367
R1728 B.n485 B.n484 163.367
R1729 B.n484 B.n59 163.367
R1730 B.n480 B.n59 163.367
R1731 B.n480 B.n479 163.367
R1732 B.n479 B.n478 163.367
R1733 B.n478 B.n61 163.367
R1734 B.n474 B.n61 163.367
R1735 B.n474 B.n473 163.367
R1736 B.n473 B.n472 163.367
R1737 B.n472 B.n63 163.367
R1738 B.n468 B.n63 163.367
R1739 B.n468 B.n467 163.367
R1740 B.n467 B.n466 163.367
R1741 B.n466 B.n65 163.367
R1742 B.n462 B.n65 163.367
R1743 B.n462 B.n461 163.367
R1744 B.n461 B.n460 163.367
R1745 B.n460 B.n67 163.367
R1746 B.n456 B.n67 163.367
R1747 B.n456 B.n455 163.367
R1748 B.n455 B.n454 163.367
R1749 B.n454 B.n69 163.367
R1750 B.n450 B.n69 163.367
R1751 B.n450 B.n449 163.367
R1752 B.n449 B.n448 163.367
R1753 B.n448 B.n71 163.367
R1754 B.n444 B.n71 163.367
R1755 B.n444 B.n443 163.367
R1756 B.n443 B.n442 163.367
R1757 B.n442 B.n73 163.367
R1758 B.n438 B.n73 163.367
R1759 B.n438 B.n437 163.367
R1760 B.n437 B.n436 163.367
R1761 B.n436 B.n75 163.367
R1762 B.n619 B.n618 163.367
R1763 B.n620 B.n619 163.367
R1764 B.n620 B.n9 163.367
R1765 B.n624 B.n9 163.367
R1766 B.n625 B.n624 163.367
R1767 B.n626 B.n625 163.367
R1768 B.n626 B.n7 163.367
R1769 B.n630 B.n7 163.367
R1770 B.n631 B.n630 163.367
R1771 B.n632 B.n631 163.367
R1772 B.n632 B.n5 163.367
R1773 B.n636 B.n5 163.367
R1774 B.n637 B.n636 163.367
R1775 B.n638 B.n637 163.367
R1776 B.n638 B.n3 163.367
R1777 B.n642 B.n3 163.367
R1778 B.n643 B.n642 163.367
R1779 B.n165 B.n2 163.367
R1780 B.n168 B.n165 163.367
R1781 B.n169 B.n168 163.367
R1782 B.n170 B.n169 163.367
R1783 B.n170 B.n163 163.367
R1784 B.n174 B.n163 163.367
R1785 B.n175 B.n174 163.367
R1786 B.n176 B.n175 163.367
R1787 B.n176 B.n161 163.367
R1788 B.n180 B.n161 163.367
R1789 B.n181 B.n180 163.367
R1790 B.n182 B.n181 163.367
R1791 B.n182 B.n159 163.367
R1792 B.n186 B.n159 163.367
R1793 B.n187 B.n186 163.367
R1794 B.n188 B.n187 163.367
R1795 B.n188 B.n157 163.367
R1796 B.n275 B.n129 59.5399
R1797 B.n290 B.n289 59.5399
R1798 B.n518 B.n47 59.5399
R1799 B.n532 B.n41 59.5399
R1800 B.n617 B.n616 32.6249
R1801 B.n434 B.n433 32.6249
R1802 B.n375 B.n94 32.6249
R1803 B.n191 B.n190 32.6249
R1804 B.n129 B.n128 23.0793
R1805 B.n289 B.n288 23.0793
R1806 B.n47 B.n46 23.0793
R1807 B.n41 B.n40 23.0793
R1808 B B.n645 18.0485
R1809 B.n617 B.n10 10.6151
R1810 B.n621 B.n10 10.6151
R1811 B.n622 B.n621 10.6151
R1812 B.n623 B.n622 10.6151
R1813 B.n623 B.n8 10.6151
R1814 B.n627 B.n8 10.6151
R1815 B.n628 B.n627 10.6151
R1816 B.n629 B.n628 10.6151
R1817 B.n629 B.n6 10.6151
R1818 B.n633 B.n6 10.6151
R1819 B.n634 B.n633 10.6151
R1820 B.n635 B.n634 10.6151
R1821 B.n635 B.n4 10.6151
R1822 B.n639 B.n4 10.6151
R1823 B.n640 B.n639 10.6151
R1824 B.n641 B.n640 10.6151
R1825 B.n641 B.n0 10.6151
R1826 B.n616 B.n615 10.6151
R1827 B.n615 B.n12 10.6151
R1828 B.n611 B.n12 10.6151
R1829 B.n611 B.n610 10.6151
R1830 B.n610 B.n609 10.6151
R1831 B.n609 B.n14 10.6151
R1832 B.n605 B.n14 10.6151
R1833 B.n605 B.n604 10.6151
R1834 B.n604 B.n603 10.6151
R1835 B.n603 B.n16 10.6151
R1836 B.n599 B.n16 10.6151
R1837 B.n599 B.n598 10.6151
R1838 B.n598 B.n597 10.6151
R1839 B.n597 B.n18 10.6151
R1840 B.n593 B.n18 10.6151
R1841 B.n593 B.n592 10.6151
R1842 B.n592 B.n591 10.6151
R1843 B.n591 B.n20 10.6151
R1844 B.n587 B.n20 10.6151
R1845 B.n587 B.n586 10.6151
R1846 B.n586 B.n585 10.6151
R1847 B.n585 B.n22 10.6151
R1848 B.n581 B.n22 10.6151
R1849 B.n581 B.n580 10.6151
R1850 B.n580 B.n579 10.6151
R1851 B.n579 B.n24 10.6151
R1852 B.n575 B.n24 10.6151
R1853 B.n575 B.n574 10.6151
R1854 B.n574 B.n573 10.6151
R1855 B.n573 B.n26 10.6151
R1856 B.n569 B.n26 10.6151
R1857 B.n569 B.n568 10.6151
R1858 B.n568 B.n567 10.6151
R1859 B.n567 B.n28 10.6151
R1860 B.n563 B.n28 10.6151
R1861 B.n563 B.n562 10.6151
R1862 B.n562 B.n561 10.6151
R1863 B.n561 B.n30 10.6151
R1864 B.n557 B.n30 10.6151
R1865 B.n557 B.n556 10.6151
R1866 B.n556 B.n555 10.6151
R1867 B.n555 B.n32 10.6151
R1868 B.n551 B.n32 10.6151
R1869 B.n551 B.n550 10.6151
R1870 B.n550 B.n549 10.6151
R1871 B.n549 B.n34 10.6151
R1872 B.n545 B.n34 10.6151
R1873 B.n545 B.n544 10.6151
R1874 B.n544 B.n543 10.6151
R1875 B.n543 B.n36 10.6151
R1876 B.n539 B.n36 10.6151
R1877 B.n539 B.n538 10.6151
R1878 B.n538 B.n537 10.6151
R1879 B.n537 B.n38 10.6151
R1880 B.n533 B.n38 10.6151
R1881 B.n531 B.n530 10.6151
R1882 B.n530 B.n42 10.6151
R1883 B.n526 B.n42 10.6151
R1884 B.n526 B.n525 10.6151
R1885 B.n525 B.n524 10.6151
R1886 B.n524 B.n44 10.6151
R1887 B.n520 B.n44 10.6151
R1888 B.n520 B.n519 10.6151
R1889 B.n517 B.n48 10.6151
R1890 B.n513 B.n48 10.6151
R1891 B.n513 B.n512 10.6151
R1892 B.n512 B.n511 10.6151
R1893 B.n511 B.n50 10.6151
R1894 B.n507 B.n50 10.6151
R1895 B.n507 B.n506 10.6151
R1896 B.n506 B.n505 10.6151
R1897 B.n505 B.n52 10.6151
R1898 B.n501 B.n52 10.6151
R1899 B.n501 B.n500 10.6151
R1900 B.n500 B.n499 10.6151
R1901 B.n499 B.n54 10.6151
R1902 B.n495 B.n54 10.6151
R1903 B.n495 B.n494 10.6151
R1904 B.n494 B.n493 10.6151
R1905 B.n493 B.n56 10.6151
R1906 B.n489 B.n56 10.6151
R1907 B.n489 B.n488 10.6151
R1908 B.n488 B.n487 10.6151
R1909 B.n487 B.n58 10.6151
R1910 B.n483 B.n58 10.6151
R1911 B.n483 B.n482 10.6151
R1912 B.n482 B.n481 10.6151
R1913 B.n481 B.n60 10.6151
R1914 B.n477 B.n60 10.6151
R1915 B.n477 B.n476 10.6151
R1916 B.n476 B.n475 10.6151
R1917 B.n475 B.n62 10.6151
R1918 B.n471 B.n62 10.6151
R1919 B.n471 B.n470 10.6151
R1920 B.n470 B.n469 10.6151
R1921 B.n469 B.n64 10.6151
R1922 B.n465 B.n64 10.6151
R1923 B.n465 B.n464 10.6151
R1924 B.n464 B.n463 10.6151
R1925 B.n463 B.n66 10.6151
R1926 B.n459 B.n66 10.6151
R1927 B.n459 B.n458 10.6151
R1928 B.n458 B.n457 10.6151
R1929 B.n457 B.n68 10.6151
R1930 B.n453 B.n68 10.6151
R1931 B.n453 B.n452 10.6151
R1932 B.n452 B.n451 10.6151
R1933 B.n451 B.n70 10.6151
R1934 B.n447 B.n70 10.6151
R1935 B.n447 B.n446 10.6151
R1936 B.n446 B.n445 10.6151
R1937 B.n445 B.n72 10.6151
R1938 B.n441 B.n72 10.6151
R1939 B.n441 B.n440 10.6151
R1940 B.n440 B.n439 10.6151
R1941 B.n439 B.n74 10.6151
R1942 B.n435 B.n74 10.6151
R1943 B.n435 B.n434 10.6151
R1944 B.n433 B.n76 10.6151
R1945 B.n429 B.n76 10.6151
R1946 B.n429 B.n428 10.6151
R1947 B.n428 B.n427 10.6151
R1948 B.n427 B.n78 10.6151
R1949 B.n423 B.n78 10.6151
R1950 B.n423 B.n422 10.6151
R1951 B.n422 B.n421 10.6151
R1952 B.n421 B.n80 10.6151
R1953 B.n417 B.n80 10.6151
R1954 B.n417 B.n416 10.6151
R1955 B.n416 B.n415 10.6151
R1956 B.n415 B.n82 10.6151
R1957 B.n411 B.n82 10.6151
R1958 B.n411 B.n410 10.6151
R1959 B.n410 B.n409 10.6151
R1960 B.n409 B.n84 10.6151
R1961 B.n405 B.n84 10.6151
R1962 B.n405 B.n404 10.6151
R1963 B.n404 B.n403 10.6151
R1964 B.n403 B.n86 10.6151
R1965 B.n399 B.n86 10.6151
R1966 B.n399 B.n398 10.6151
R1967 B.n398 B.n397 10.6151
R1968 B.n397 B.n88 10.6151
R1969 B.n393 B.n88 10.6151
R1970 B.n393 B.n392 10.6151
R1971 B.n392 B.n391 10.6151
R1972 B.n391 B.n90 10.6151
R1973 B.n387 B.n90 10.6151
R1974 B.n387 B.n386 10.6151
R1975 B.n386 B.n385 10.6151
R1976 B.n385 B.n92 10.6151
R1977 B.n381 B.n92 10.6151
R1978 B.n381 B.n380 10.6151
R1979 B.n380 B.n379 10.6151
R1980 B.n379 B.n94 10.6151
R1981 B.n166 B.n1 10.6151
R1982 B.n167 B.n166 10.6151
R1983 B.n167 B.n164 10.6151
R1984 B.n171 B.n164 10.6151
R1985 B.n172 B.n171 10.6151
R1986 B.n173 B.n172 10.6151
R1987 B.n173 B.n162 10.6151
R1988 B.n177 B.n162 10.6151
R1989 B.n178 B.n177 10.6151
R1990 B.n179 B.n178 10.6151
R1991 B.n179 B.n160 10.6151
R1992 B.n183 B.n160 10.6151
R1993 B.n184 B.n183 10.6151
R1994 B.n185 B.n184 10.6151
R1995 B.n185 B.n158 10.6151
R1996 B.n189 B.n158 10.6151
R1997 B.n190 B.n189 10.6151
R1998 B.n191 B.n156 10.6151
R1999 B.n195 B.n156 10.6151
R2000 B.n196 B.n195 10.6151
R2001 B.n197 B.n196 10.6151
R2002 B.n197 B.n154 10.6151
R2003 B.n201 B.n154 10.6151
R2004 B.n202 B.n201 10.6151
R2005 B.n203 B.n202 10.6151
R2006 B.n203 B.n152 10.6151
R2007 B.n207 B.n152 10.6151
R2008 B.n208 B.n207 10.6151
R2009 B.n209 B.n208 10.6151
R2010 B.n209 B.n150 10.6151
R2011 B.n213 B.n150 10.6151
R2012 B.n214 B.n213 10.6151
R2013 B.n215 B.n214 10.6151
R2014 B.n215 B.n148 10.6151
R2015 B.n219 B.n148 10.6151
R2016 B.n220 B.n219 10.6151
R2017 B.n221 B.n220 10.6151
R2018 B.n221 B.n146 10.6151
R2019 B.n225 B.n146 10.6151
R2020 B.n226 B.n225 10.6151
R2021 B.n227 B.n226 10.6151
R2022 B.n227 B.n144 10.6151
R2023 B.n231 B.n144 10.6151
R2024 B.n232 B.n231 10.6151
R2025 B.n233 B.n232 10.6151
R2026 B.n233 B.n142 10.6151
R2027 B.n237 B.n142 10.6151
R2028 B.n238 B.n237 10.6151
R2029 B.n239 B.n238 10.6151
R2030 B.n239 B.n140 10.6151
R2031 B.n243 B.n140 10.6151
R2032 B.n244 B.n243 10.6151
R2033 B.n245 B.n244 10.6151
R2034 B.n245 B.n138 10.6151
R2035 B.n249 B.n138 10.6151
R2036 B.n250 B.n249 10.6151
R2037 B.n251 B.n250 10.6151
R2038 B.n251 B.n136 10.6151
R2039 B.n255 B.n136 10.6151
R2040 B.n256 B.n255 10.6151
R2041 B.n257 B.n256 10.6151
R2042 B.n257 B.n134 10.6151
R2043 B.n261 B.n134 10.6151
R2044 B.n262 B.n261 10.6151
R2045 B.n263 B.n262 10.6151
R2046 B.n263 B.n132 10.6151
R2047 B.n267 B.n132 10.6151
R2048 B.n268 B.n267 10.6151
R2049 B.n269 B.n268 10.6151
R2050 B.n269 B.n130 10.6151
R2051 B.n273 B.n130 10.6151
R2052 B.n274 B.n273 10.6151
R2053 B.n276 B.n126 10.6151
R2054 B.n280 B.n126 10.6151
R2055 B.n281 B.n280 10.6151
R2056 B.n282 B.n281 10.6151
R2057 B.n282 B.n124 10.6151
R2058 B.n286 B.n124 10.6151
R2059 B.n287 B.n286 10.6151
R2060 B.n291 B.n287 10.6151
R2061 B.n295 B.n122 10.6151
R2062 B.n296 B.n295 10.6151
R2063 B.n297 B.n296 10.6151
R2064 B.n297 B.n120 10.6151
R2065 B.n301 B.n120 10.6151
R2066 B.n302 B.n301 10.6151
R2067 B.n303 B.n302 10.6151
R2068 B.n303 B.n118 10.6151
R2069 B.n307 B.n118 10.6151
R2070 B.n308 B.n307 10.6151
R2071 B.n309 B.n308 10.6151
R2072 B.n309 B.n116 10.6151
R2073 B.n313 B.n116 10.6151
R2074 B.n314 B.n313 10.6151
R2075 B.n315 B.n314 10.6151
R2076 B.n315 B.n114 10.6151
R2077 B.n319 B.n114 10.6151
R2078 B.n320 B.n319 10.6151
R2079 B.n321 B.n320 10.6151
R2080 B.n321 B.n112 10.6151
R2081 B.n325 B.n112 10.6151
R2082 B.n326 B.n325 10.6151
R2083 B.n327 B.n326 10.6151
R2084 B.n327 B.n110 10.6151
R2085 B.n331 B.n110 10.6151
R2086 B.n332 B.n331 10.6151
R2087 B.n333 B.n332 10.6151
R2088 B.n333 B.n108 10.6151
R2089 B.n337 B.n108 10.6151
R2090 B.n338 B.n337 10.6151
R2091 B.n339 B.n338 10.6151
R2092 B.n339 B.n106 10.6151
R2093 B.n343 B.n106 10.6151
R2094 B.n344 B.n343 10.6151
R2095 B.n345 B.n344 10.6151
R2096 B.n345 B.n104 10.6151
R2097 B.n349 B.n104 10.6151
R2098 B.n350 B.n349 10.6151
R2099 B.n351 B.n350 10.6151
R2100 B.n351 B.n102 10.6151
R2101 B.n355 B.n102 10.6151
R2102 B.n356 B.n355 10.6151
R2103 B.n357 B.n356 10.6151
R2104 B.n357 B.n100 10.6151
R2105 B.n361 B.n100 10.6151
R2106 B.n362 B.n361 10.6151
R2107 B.n363 B.n362 10.6151
R2108 B.n363 B.n98 10.6151
R2109 B.n367 B.n98 10.6151
R2110 B.n368 B.n367 10.6151
R2111 B.n369 B.n368 10.6151
R2112 B.n369 B.n96 10.6151
R2113 B.n373 B.n96 10.6151
R2114 B.n374 B.n373 10.6151
R2115 B.n375 B.n374 10.6151
R2116 B.n645 B.n0 8.11757
R2117 B.n645 B.n1 8.11757
R2118 B.n532 B.n531 6.5566
R2119 B.n519 B.n518 6.5566
R2120 B.n276 B.n275 6.5566
R2121 B.n291 B.n290 6.5566
R2122 B.n533 B.n532 4.05904
R2123 B.n518 B.n517 4.05904
R2124 B.n275 B.n274 4.05904
R2125 B.n290 B.n122 4.05904
R2126 VP.n1 VP.t2 536.904
R2127 VP.n1 VP.t1 536.856
R2128 VP.n3 VP.t0 515.909
R2129 VP.n5 VP.t3 515.909
R2130 VP.n6 VP.n5 161.3
R2131 VP.n4 VP.n0 161.3
R2132 VP.n3 VP.n2 161.3
R2133 VP.n2 VP.n1 89.2833
R2134 VP.n4 VP.n3 24.1005
R2135 VP.n5 VP.n4 24.1005
R2136 VP.n2 VP.n0 0.189894
R2137 VP.n6 VP.n0 0.189894
R2138 VP VP.n6 0.0516364
R2139 VDD1 VDD1.n1 110.382
R2140 VDD1 VDD1.n0 68.6743
R2141 VDD1.n0 VDD1.t1 1.93994
R2142 VDD1.n0 VDD1.t2 1.93994
R2143 VDD1.n1 VDD1.t3 1.93994
R2144 VDD1.n1 VDD1.t0 1.93994
C0 B VDD2 1.10666f
C1 B VTAIL 5.25966f
C2 VP VN 5.81814f
C3 VDD2 VN 4.70939f
C4 VTAIL VN 4.15181f
C5 B VN 0.830993f
C6 VDD1 w_n1684_n4320# 1.22469f
C7 VP w_n1684_n4320# 2.82837f
C8 w_n1684_n4320# VDD2 1.24241f
C9 VTAIL w_n1684_n4320# 5.28209f
C10 VP VDD1 4.84525f
C11 VDD1 VDD2 0.603454f
C12 VTAIL VDD1 8.227599f
C13 VP VDD2 0.28306f
C14 B w_n1684_n4320# 8.43904f
C15 VP VTAIL 4.16592f
C16 VTAIL VDD2 8.27015f
C17 B VDD1 1.0828f
C18 w_n1684_n4320# VN 2.61629f
C19 VDD1 VN 0.146902f
C20 B VP 1.17484f
C21 VDD2 VSUBS 0.812724f
C22 VDD1 VSUBS 5.630316f
C23 VTAIL VSUBS 1.125299f
C24 VN VSUBS 6.11953f
C25 VP VSUBS 1.555025f
C26 B VSUBS 3.1596f
C27 w_n1684_n4320# VSUBS 89.0567f
C28 VDD1.t1 VSUBS 0.363932f
C29 VDD1.t2 VSUBS 0.363932f
C30 VDD1.n0 VSUBS 2.99258f
C31 VDD1.t3 VSUBS 0.363932f
C32 VDD1.t0 VSUBS 0.363932f
C33 VDD1.n1 VSUBS 3.85871f
C34 VP.n0 VSUBS 0.05457f
C35 VP.t1 VSUBS 2.26582f
C36 VP.t2 VSUBS 2.2659f
C37 VP.n1 VSUBS 2.93877f
C38 VP.n2 VSUBS 3.83821f
C39 VP.t0 VSUBS 2.23278f
C40 VP.n3 VSUBS 0.842862f
C41 VP.n4 VSUBS 0.012383f
C42 VP.t3 VSUBS 2.23278f
C43 VP.n5 VSUBS 0.842862f
C44 VP.n6 VSUBS 0.04229f
C45 B.n0 VSUBS 0.006714f
C46 B.n1 VSUBS 0.006714f
C47 B.n2 VSUBS 0.009929f
C48 B.n3 VSUBS 0.007609f
C49 B.n4 VSUBS 0.007609f
C50 B.n5 VSUBS 0.007609f
C51 B.n6 VSUBS 0.007609f
C52 B.n7 VSUBS 0.007609f
C53 B.n8 VSUBS 0.007609f
C54 B.n9 VSUBS 0.007609f
C55 B.n10 VSUBS 0.007609f
C56 B.n11 VSUBS 0.018373f
C57 B.n12 VSUBS 0.007609f
C58 B.n13 VSUBS 0.007609f
C59 B.n14 VSUBS 0.007609f
C60 B.n15 VSUBS 0.007609f
C61 B.n16 VSUBS 0.007609f
C62 B.n17 VSUBS 0.007609f
C63 B.n18 VSUBS 0.007609f
C64 B.n19 VSUBS 0.007609f
C65 B.n20 VSUBS 0.007609f
C66 B.n21 VSUBS 0.007609f
C67 B.n22 VSUBS 0.007609f
C68 B.n23 VSUBS 0.007609f
C69 B.n24 VSUBS 0.007609f
C70 B.n25 VSUBS 0.007609f
C71 B.n26 VSUBS 0.007609f
C72 B.n27 VSUBS 0.007609f
C73 B.n28 VSUBS 0.007609f
C74 B.n29 VSUBS 0.007609f
C75 B.n30 VSUBS 0.007609f
C76 B.n31 VSUBS 0.007609f
C77 B.n32 VSUBS 0.007609f
C78 B.n33 VSUBS 0.007609f
C79 B.n34 VSUBS 0.007609f
C80 B.n35 VSUBS 0.007609f
C81 B.n36 VSUBS 0.007609f
C82 B.n37 VSUBS 0.007609f
C83 B.n38 VSUBS 0.007609f
C84 B.n39 VSUBS 0.007609f
C85 B.t7 VSUBS 0.349085f
C86 B.t8 VSUBS 0.364447f
C87 B.t6 VSUBS 0.642276f
C88 B.n40 VSUBS 0.468163f
C89 B.n41 VSUBS 0.333261f
C90 B.n42 VSUBS 0.007609f
C91 B.n43 VSUBS 0.007609f
C92 B.n44 VSUBS 0.007609f
C93 B.n45 VSUBS 0.007609f
C94 B.t10 VSUBS 0.349088f
C95 B.t11 VSUBS 0.364451f
C96 B.t9 VSUBS 0.642276f
C97 B.n46 VSUBS 0.46816f
C98 B.n47 VSUBS 0.333257f
C99 B.n48 VSUBS 0.007609f
C100 B.n49 VSUBS 0.007609f
C101 B.n50 VSUBS 0.007609f
C102 B.n51 VSUBS 0.007609f
C103 B.n52 VSUBS 0.007609f
C104 B.n53 VSUBS 0.007609f
C105 B.n54 VSUBS 0.007609f
C106 B.n55 VSUBS 0.007609f
C107 B.n56 VSUBS 0.007609f
C108 B.n57 VSUBS 0.007609f
C109 B.n58 VSUBS 0.007609f
C110 B.n59 VSUBS 0.007609f
C111 B.n60 VSUBS 0.007609f
C112 B.n61 VSUBS 0.007609f
C113 B.n62 VSUBS 0.007609f
C114 B.n63 VSUBS 0.007609f
C115 B.n64 VSUBS 0.007609f
C116 B.n65 VSUBS 0.007609f
C117 B.n66 VSUBS 0.007609f
C118 B.n67 VSUBS 0.007609f
C119 B.n68 VSUBS 0.007609f
C120 B.n69 VSUBS 0.007609f
C121 B.n70 VSUBS 0.007609f
C122 B.n71 VSUBS 0.007609f
C123 B.n72 VSUBS 0.007609f
C124 B.n73 VSUBS 0.007609f
C125 B.n74 VSUBS 0.007609f
C126 B.n75 VSUBS 0.018373f
C127 B.n76 VSUBS 0.007609f
C128 B.n77 VSUBS 0.007609f
C129 B.n78 VSUBS 0.007609f
C130 B.n79 VSUBS 0.007609f
C131 B.n80 VSUBS 0.007609f
C132 B.n81 VSUBS 0.007609f
C133 B.n82 VSUBS 0.007609f
C134 B.n83 VSUBS 0.007609f
C135 B.n84 VSUBS 0.007609f
C136 B.n85 VSUBS 0.007609f
C137 B.n86 VSUBS 0.007609f
C138 B.n87 VSUBS 0.007609f
C139 B.n88 VSUBS 0.007609f
C140 B.n89 VSUBS 0.007609f
C141 B.n90 VSUBS 0.007609f
C142 B.n91 VSUBS 0.007609f
C143 B.n92 VSUBS 0.007609f
C144 B.n93 VSUBS 0.007609f
C145 B.n94 VSUBS 0.01811f
C146 B.n95 VSUBS 0.007609f
C147 B.n96 VSUBS 0.007609f
C148 B.n97 VSUBS 0.007609f
C149 B.n98 VSUBS 0.007609f
C150 B.n99 VSUBS 0.007609f
C151 B.n100 VSUBS 0.007609f
C152 B.n101 VSUBS 0.007609f
C153 B.n102 VSUBS 0.007609f
C154 B.n103 VSUBS 0.007609f
C155 B.n104 VSUBS 0.007609f
C156 B.n105 VSUBS 0.007609f
C157 B.n106 VSUBS 0.007609f
C158 B.n107 VSUBS 0.007609f
C159 B.n108 VSUBS 0.007609f
C160 B.n109 VSUBS 0.007609f
C161 B.n110 VSUBS 0.007609f
C162 B.n111 VSUBS 0.007609f
C163 B.n112 VSUBS 0.007609f
C164 B.n113 VSUBS 0.007609f
C165 B.n114 VSUBS 0.007609f
C166 B.n115 VSUBS 0.007609f
C167 B.n116 VSUBS 0.007609f
C168 B.n117 VSUBS 0.007609f
C169 B.n118 VSUBS 0.007609f
C170 B.n119 VSUBS 0.007609f
C171 B.n120 VSUBS 0.007609f
C172 B.n121 VSUBS 0.007609f
C173 B.n122 VSUBS 0.005259f
C174 B.n123 VSUBS 0.007609f
C175 B.n124 VSUBS 0.007609f
C176 B.n125 VSUBS 0.007609f
C177 B.n126 VSUBS 0.007609f
C178 B.n127 VSUBS 0.007609f
C179 B.t2 VSUBS 0.349085f
C180 B.t1 VSUBS 0.364447f
C181 B.t0 VSUBS 0.642276f
C182 B.n128 VSUBS 0.468163f
C183 B.n129 VSUBS 0.333261f
C184 B.n130 VSUBS 0.007609f
C185 B.n131 VSUBS 0.007609f
C186 B.n132 VSUBS 0.007609f
C187 B.n133 VSUBS 0.007609f
C188 B.n134 VSUBS 0.007609f
C189 B.n135 VSUBS 0.007609f
C190 B.n136 VSUBS 0.007609f
C191 B.n137 VSUBS 0.007609f
C192 B.n138 VSUBS 0.007609f
C193 B.n139 VSUBS 0.007609f
C194 B.n140 VSUBS 0.007609f
C195 B.n141 VSUBS 0.007609f
C196 B.n142 VSUBS 0.007609f
C197 B.n143 VSUBS 0.007609f
C198 B.n144 VSUBS 0.007609f
C199 B.n145 VSUBS 0.007609f
C200 B.n146 VSUBS 0.007609f
C201 B.n147 VSUBS 0.007609f
C202 B.n148 VSUBS 0.007609f
C203 B.n149 VSUBS 0.007609f
C204 B.n150 VSUBS 0.007609f
C205 B.n151 VSUBS 0.007609f
C206 B.n152 VSUBS 0.007609f
C207 B.n153 VSUBS 0.007609f
C208 B.n154 VSUBS 0.007609f
C209 B.n155 VSUBS 0.007609f
C210 B.n156 VSUBS 0.007609f
C211 B.n157 VSUBS 0.01721f
C212 B.n158 VSUBS 0.007609f
C213 B.n159 VSUBS 0.007609f
C214 B.n160 VSUBS 0.007609f
C215 B.n161 VSUBS 0.007609f
C216 B.n162 VSUBS 0.007609f
C217 B.n163 VSUBS 0.007609f
C218 B.n164 VSUBS 0.007609f
C219 B.n165 VSUBS 0.007609f
C220 B.n166 VSUBS 0.007609f
C221 B.n167 VSUBS 0.007609f
C222 B.n168 VSUBS 0.007609f
C223 B.n169 VSUBS 0.007609f
C224 B.n170 VSUBS 0.007609f
C225 B.n171 VSUBS 0.007609f
C226 B.n172 VSUBS 0.007609f
C227 B.n173 VSUBS 0.007609f
C228 B.n174 VSUBS 0.007609f
C229 B.n175 VSUBS 0.007609f
C230 B.n176 VSUBS 0.007609f
C231 B.n177 VSUBS 0.007609f
C232 B.n178 VSUBS 0.007609f
C233 B.n179 VSUBS 0.007609f
C234 B.n180 VSUBS 0.007609f
C235 B.n181 VSUBS 0.007609f
C236 B.n182 VSUBS 0.007609f
C237 B.n183 VSUBS 0.007609f
C238 B.n184 VSUBS 0.007609f
C239 B.n185 VSUBS 0.007609f
C240 B.n186 VSUBS 0.007609f
C241 B.n187 VSUBS 0.007609f
C242 B.n188 VSUBS 0.007609f
C243 B.n189 VSUBS 0.007609f
C244 B.n190 VSUBS 0.01721f
C245 B.n191 VSUBS 0.018373f
C246 B.n192 VSUBS 0.018373f
C247 B.n193 VSUBS 0.007609f
C248 B.n194 VSUBS 0.007609f
C249 B.n195 VSUBS 0.007609f
C250 B.n196 VSUBS 0.007609f
C251 B.n197 VSUBS 0.007609f
C252 B.n198 VSUBS 0.007609f
C253 B.n199 VSUBS 0.007609f
C254 B.n200 VSUBS 0.007609f
C255 B.n201 VSUBS 0.007609f
C256 B.n202 VSUBS 0.007609f
C257 B.n203 VSUBS 0.007609f
C258 B.n204 VSUBS 0.007609f
C259 B.n205 VSUBS 0.007609f
C260 B.n206 VSUBS 0.007609f
C261 B.n207 VSUBS 0.007609f
C262 B.n208 VSUBS 0.007609f
C263 B.n209 VSUBS 0.007609f
C264 B.n210 VSUBS 0.007609f
C265 B.n211 VSUBS 0.007609f
C266 B.n212 VSUBS 0.007609f
C267 B.n213 VSUBS 0.007609f
C268 B.n214 VSUBS 0.007609f
C269 B.n215 VSUBS 0.007609f
C270 B.n216 VSUBS 0.007609f
C271 B.n217 VSUBS 0.007609f
C272 B.n218 VSUBS 0.007609f
C273 B.n219 VSUBS 0.007609f
C274 B.n220 VSUBS 0.007609f
C275 B.n221 VSUBS 0.007609f
C276 B.n222 VSUBS 0.007609f
C277 B.n223 VSUBS 0.007609f
C278 B.n224 VSUBS 0.007609f
C279 B.n225 VSUBS 0.007609f
C280 B.n226 VSUBS 0.007609f
C281 B.n227 VSUBS 0.007609f
C282 B.n228 VSUBS 0.007609f
C283 B.n229 VSUBS 0.007609f
C284 B.n230 VSUBS 0.007609f
C285 B.n231 VSUBS 0.007609f
C286 B.n232 VSUBS 0.007609f
C287 B.n233 VSUBS 0.007609f
C288 B.n234 VSUBS 0.007609f
C289 B.n235 VSUBS 0.007609f
C290 B.n236 VSUBS 0.007609f
C291 B.n237 VSUBS 0.007609f
C292 B.n238 VSUBS 0.007609f
C293 B.n239 VSUBS 0.007609f
C294 B.n240 VSUBS 0.007609f
C295 B.n241 VSUBS 0.007609f
C296 B.n242 VSUBS 0.007609f
C297 B.n243 VSUBS 0.007609f
C298 B.n244 VSUBS 0.007609f
C299 B.n245 VSUBS 0.007609f
C300 B.n246 VSUBS 0.007609f
C301 B.n247 VSUBS 0.007609f
C302 B.n248 VSUBS 0.007609f
C303 B.n249 VSUBS 0.007609f
C304 B.n250 VSUBS 0.007609f
C305 B.n251 VSUBS 0.007609f
C306 B.n252 VSUBS 0.007609f
C307 B.n253 VSUBS 0.007609f
C308 B.n254 VSUBS 0.007609f
C309 B.n255 VSUBS 0.007609f
C310 B.n256 VSUBS 0.007609f
C311 B.n257 VSUBS 0.007609f
C312 B.n258 VSUBS 0.007609f
C313 B.n259 VSUBS 0.007609f
C314 B.n260 VSUBS 0.007609f
C315 B.n261 VSUBS 0.007609f
C316 B.n262 VSUBS 0.007609f
C317 B.n263 VSUBS 0.007609f
C318 B.n264 VSUBS 0.007609f
C319 B.n265 VSUBS 0.007609f
C320 B.n266 VSUBS 0.007609f
C321 B.n267 VSUBS 0.007609f
C322 B.n268 VSUBS 0.007609f
C323 B.n269 VSUBS 0.007609f
C324 B.n270 VSUBS 0.007609f
C325 B.n271 VSUBS 0.007609f
C326 B.n272 VSUBS 0.007609f
C327 B.n273 VSUBS 0.007609f
C328 B.n274 VSUBS 0.005259f
C329 B.n275 VSUBS 0.017629f
C330 B.n276 VSUBS 0.006154f
C331 B.n277 VSUBS 0.007609f
C332 B.n278 VSUBS 0.007609f
C333 B.n279 VSUBS 0.007609f
C334 B.n280 VSUBS 0.007609f
C335 B.n281 VSUBS 0.007609f
C336 B.n282 VSUBS 0.007609f
C337 B.n283 VSUBS 0.007609f
C338 B.n284 VSUBS 0.007609f
C339 B.n285 VSUBS 0.007609f
C340 B.n286 VSUBS 0.007609f
C341 B.n287 VSUBS 0.007609f
C342 B.t5 VSUBS 0.349088f
C343 B.t4 VSUBS 0.364451f
C344 B.t3 VSUBS 0.642276f
C345 B.n288 VSUBS 0.46816f
C346 B.n289 VSUBS 0.333257f
C347 B.n290 VSUBS 0.017629f
C348 B.n291 VSUBS 0.006154f
C349 B.n292 VSUBS 0.007609f
C350 B.n293 VSUBS 0.007609f
C351 B.n294 VSUBS 0.007609f
C352 B.n295 VSUBS 0.007609f
C353 B.n296 VSUBS 0.007609f
C354 B.n297 VSUBS 0.007609f
C355 B.n298 VSUBS 0.007609f
C356 B.n299 VSUBS 0.007609f
C357 B.n300 VSUBS 0.007609f
C358 B.n301 VSUBS 0.007609f
C359 B.n302 VSUBS 0.007609f
C360 B.n303 VSUBS 0.007609f
C361 B.n304 VSUBS 0.007609f
C362 B.n305 VSUBS 0.007609f
C363 B.n306 VSUBS 0.007609f
C364 B.n307 VSUBS 0.007609f
C365 B.n308 VSUBS 0.007609f
C366 B.n309 VSUBS 0.007609f
C367 B.n310 VSUBS 0.007609f
C368 B.n311 VSUBS 0.007609f
C369 B.n312 VSUBS 0.007609f
C370 B.n313 VSUBS 0.007609f
C371 B.n314 VSUBS 0.007609f
C372 B.n315 VSUBS 0.007609f
C373 B.n316 VSUBS 0.007609f
C374 B.n317 VSUBS 0.007609f
C375 B.n318 VSUBS 0.007609f
C376 B.n319 VSUBS 0.007609f
C377 B.n320 VSUBS 0.007609f
C378 B.n321 VSUBS 0.007609f
C379 B.n322 VSUBS 0.007609f
C380 B.n323 VSUBS 0.007609f
C381 B.n324 VSUBS 0.007609f
C382 B.n325 VSUBS 0.007609f
C383 B.n326 VSUBS 0.007609f
C384 B.n327 VSUBS 0.007609f
C385 B.n328 VSUBS 0.007609f
C386 B.n329 VSUBS 0.007609f
C387 B.n330 VSUBS 0.007609f
C388 B.n331 VSUBS 0.007609f
C389 B.n332 VSUBS 0.007609f
C390 B.n333 VSUBS 0.007609f
C391 B.n334 VSUBS 0.007609f
C392 B.n335 VSUBS 0.007609f
C393 B.n336 VSUBS 0.007609f
C394 B.n337 VSUBS 0.007609f
C395 B.n338 VSUBS 0.007609f
C396 B.n339 VSUBS 0.007609f
C397 B.n340 VSUBS 0.007609f
C398 B.n341 VSUBS 0.007609f
C399 B.n342 VSUBS 0.007609f
C400 B.n343 VSUBS 0.007609f
C401 B.n344 VSUBS 0.007609f
C402 B.n345 VSUBS 0.007609f
C403 B.n346 VSUBS 0.007609f
C404 B.n347 VSUBS 0.007609f
C405 B.n348 VSUBS 0.007609f
C406 B.n349 VSUBS 0.007609f
C407 B.n350 VSUBS 0.007609f
C408 B.n351 VSUBS 0.007609f
C409 B.n352 VSUBS 0.007609f
C410 B.n353 VSUBS 0.007609f
C411 B.n354 VSUBS 0.007609f
C412 B.n355 VSUBS 0.007609f
C413 B.n356 VSUBS 0.007609f
C414 B.n357 VSUBS 0.007609f
C415 B.n358 VSUBS 0.007609f
C416 B.n359 VSUBS 0.007609f
C417 B.n360 VSUBS 0.007609f
C418 B.n361 VSUBS 0.007609f
C419 B.n362 VSUBS 0.007609f
C420 B.n363 VSUBS 0.007609f
C421 B.n364 VSUBS 0.007609f
C422 B.n365 VSUBS 0.007609f
C423 B.n366 VSUBS 0.007609f
C424 B.n367 VSUBS 0.007609f
C425 B.n368 VSUBS 0.007609f
C426 B.n369 VSUBS 0.007609f
C427 B.n370 VSUBS 0.007609f
C428 B.n371 VSUBS 0.007609f
C429 B.n372 VSUBS 0.007609f
C430 B.n373 VSUBS 0.007609f
C431 B.n374 VSUBS 0.007609f
C432 B.n375 VSUBS 0.017473f
C433 B.n376 VSUBS 0.018373f
C434 B.n377 VSUBS 0.01721f
C435 B.n378 VSUBS 0.007609f
C436 B.n379 VSUBS 0.007609f
C437 B.n380 VSUBS 0.007609f
C438 B.n381 VSUBS 0.007609f
C439 B.n382 VSUBS 0.007609f
C440 B.n383 VSUBS 0.007609f
C441 B.n384 VSUBS 0.007609f
C442 B.n385 VSUBS 0.007609f
C443 B.n386 VSUBS 0.007609f
C444 B.n387 VSUBS 0.007609f
C445 B.n388 VSUBS 0.007609f
C446 B.n389 VSUBS 0.007609f
C447 B.n390 VSUBS 0.007609f
C448 B.n391 VSUBS 0.007609f
C449 B.n392 VSUBS 0.007609f
C450 B.n393 VSUBS 0.007609f
C451 B.n394 VSUBS 0.007609f
C452 B.n395 VSUBS 0.007609f
C453 B.n396 VSUBS 0.007609f
C454 B.n397 VSUBS 0.007609f
C455 B.n398 VSUBS 0.007609f
C456 B.n399 VSUBS 0.007609f
C457 B.n400 VSUBS 0.007609f
C458 B.n401 VSUBS 0.007609f
C459 B.n402 VSUBS 0.007609f
C460 B.n403 VSUBS 0.007609f
C461 B.n404 VSUBS 0.007609f
C462 B.n405 VSUBS 0.007609f
C463 B.n406 VSUBS 0.007609f
C464 B.n407 VSUBS 0.007609f
C465 B.n408 VSUBS 0.007609f
C466 B.n409 VSUBS 0.007609f
C467 B.n410 VSUBS 0.007609f
C468 B.n411 VSUBS 0.007609f
C469 B.n412 VSUBS 0.007609f
C470 B.n413 VSUBS 0.007609f
C471 B.n414 VSUBS 0.007609f
C472 B.n415 VSUBS 0.007609f
C473 B.n416 VSUBS 0.007609f
C474 B.n417 VSUBS 0.007609f
C475 B.n418 VSUBS 0.007609f
C476 B.n419 VSUBS 0.007609f
C477 B.n420 VSUBS 0.007609f
C478 B.n421 VSUBS 0.007609f
C479 B.n422 VSUBS 0.007609f
C480 B.n423 VSUBS 0.007609f
C481 B.n424 VSUBS 0.007609f
C482 B.n425 VSUBS 0.007609f
C483 B.n426 VSUBS 0.007609f
C484 B.n427 VSUBS 0.007609f
C485 B.n428 VSUBS 0.007609f
C486 B.n429 VSUBS 0.007609f
C487 B.n430 VSUBS 0.007609f
C488 B.n431 VSUBS 0.007609f
C489 B.n432 VSUBS 0.01721f
C490 B.n433 VSUBS 0.01721f
C491 B.n434 VSUBS 0.018373f
C492 B.n435 VSUBS 0.007609f
C493 B.n436 VSUBS 0.007609f
C494 B.n437 VSUBS 0.007609f
C495 B.n438 VSUBS 0.007609f
C496 B.n439 VSUBS 0.007609f
C497 B.n440 VSUBS 0.007609f
C498 B.n441 VSUBS 0.007609f
C499 B.n442 VSUBS 0.007609f
C500 B.n443 VSUBS 0.007609f
C501 B.n444 VSUBS 0.007609f
C502 B.n445 VSUBS 0.007609f
C503 B.n446 VSUBS 0.007609f
C504 B.n447 VSUBS 0.007609f
C505 B.n448 VSUBS 0.007609f
C506 B.n449 VSUBS 0.007609f
C507 B.n450 VSUBS 0.007609f
C508 B.n451 VSUBS 0.007609f
C509 B.n452 VSUBS 0.007609f
C510 B.n453 VSUBS 0.007609f
C511 B.n454 VSUBS 0.007609f
C512 B.n455 VSUBS 0.007609f
C513 B.n456 VSUBS 0.007609f
C514 B.n457 VSUBS 0.007609f
C515 B.n458 VSUBS 0.007609f
C516 B.n459 VSUBS 0.007609f
C517 B.n460 VSUBS 0.007609f
C518 B.n461 VSUBS 0.007609f
C519 B.n462 VSUBS 0.007609f
C520 B.n463 VSUBS 0.007609f
C521 B.n464 VSUBS 0.007609f
C522 B.n465 VSUBS 0.007609f
C523 B.n466 VSUBS 0.007609f
C524 B.n467 VSUBS 0.007609f
C525 B.n468 VSUBS 0.007609f
C526 B.n469 VSUBS 0.007609f
C527 B.n470 VSUBS 0.007609f
C528 B.n471 VSUBS 0.007609f
C529 B.n472 VSUBS 0.007609f
C530 B.n473 VSUBS 0.007609f
C531 B.n474 VSUBS 0.007609f
C532 B.n475 VSUBS 0.007609f
C533 B.n476 VSUBS 0.007609f
C534 B.n477 VSUBS 0.007609f
C535 B.n478 VSUBS 0.007609f
C536 B.n479 VSUBS 0.007609f
C537 B.n480 VSUBS 0.007609f
C538 B.n481 VSUBS 0.007609f
C539 B.n482 VSUBS 0.007609f
C540 B.n483 VSUBS 0.007609f
C541 B.n484 VSUBS 0.007609f
C542 B.n485 VSUBS 0.007609f
C543 B.n486 VSUBS 0.007609f
C544 B.n487 VSUBS 0.007609f
C545 B.n488 VSUBS 0.007609f
C546 B.n489 VSUBS 0.007609f
C547 B.n490 VSUBS 0.007609f
C548 B.n491 VSUBS 0.007609f
C549 B.n492 VSUBS 0.007609f
C550 B.n493 VSUBS 0.007609f
C551 B.n494 VSUBS 0.007609f
C552 B.n495 VSUBS 0.007609f
C553 B.n496 VSUBS 0.007609f
C554 B.n497 VSUBS 0.007609f
C555 B.n498 VSUBS 0.007609f
C556 B.n499 VSUBS 0.007609f
C557 B.n500 VSUBS 0.007609f
C558 B.n501 VSUBS 0.007609f
C559 B.n502 VSUBS 0.007609f
C560 B.n503 VSUBS 0.007609f
C561 B.n504 VSUBS 0.007609f
C562 B.n505 VSUBS 0.007609f
C563 B.n506 VSUBS 0.007609f
C564 B.n507 VSUBS 0.007609f
C565 B.n508 VSUBS 0.007609f
C566 B.n509 VSUBS 0.007609f
C567 B.n510 VSUBS 0.007609f
C568 B.n511 VSUBS 0.007609f
C569 B.n512 VSUBS 0.007609f
C570 B.n513 VSUBS 0.007609f
C571 B.n514 VSUBS 0.007609f
C572 B.n515 VSUBS 0.007609f
C573 B.n516 VSUBS 0.007609f
C574 B.n517 VSUBS 0.005259f
C575 B.n518 VSUBS 0.017629f
C576 B.n519 VSUBS 0.006154f
C577 B.n520 VSUBS 0.007609f
C578 B.n521 VSUBS 0.007609f
C579 B.n522 VSUBS 0.007609f
C580 B.n523 VSUBS 0.007609f
C581 B.n524 VSUBS 0.007609f
C582 B.n525 VSUBS 0.007609f
C583 B.n526 VSUBS 0.007609f
C584 B.n527 VSUBS 0.007609f
C585 B.n528 VSUBS 0.007609f
C586 B.n529 VSUBS 0.007609f
C587 B.n530 VSUBS 0.007609f
C588 B.n531 VSUBS 0.006154f
C589 B.n532 VSUBS 0.017629f
C590 B.n533 VSUBS 0.005259f
C591 B.n534 VSUBS 0.007609f
C592 B.n535 VSUBS 0.007609f
C593 B.n536 VSUBS 0.007609f
C594 B.n537 VSUBS 0.007609f
C595 B.n538 VSUBS 0.007609f
C596 B.n539 VSUBS 0.007609f
C597 B.n540 VSUBS 0.007609f
C598 B.n541 VSUBS 0.007609f
C599 B.n542 VSUBS 0.007609f
C600 B.n543 VSUBS 0.007609f
C601 B.n544 VSUBS 0.007609f
C602 B.n545 VSUBS 0.007609f
C603 B.n546 VSUBS 0.007609f
C604 B.n547 VSUBS 0.007609f
C605 B.n548 VSUBS 0.007609f
C606 B.n549 VSUBS 0.007609f
C607 B.n550 VSUBS 0.007609f
C608 B.n551 VSUBS 0.007609f
C609 B.n552 VSUBS 0.007609f
C610 B.n553 VSUBS 0.007609f
C611 B.n554 VSUBS 0.007609f
C612 B.n555 VSUBS 0.007609f
C613 B.n556 VSUBS 0.007609f
C614 B.n557 VSUBS 0.007609f
C615 B.n558 VSUBS 0.007609f
C616 B.n559 VSUBS 0.007609f
C617 B.n560 VSUBS 0.007609f
C618 B.n561 VSUBS 0.007609f
C619 B.n562 VSUBS 0.007609f
C620 B.n563 VSUBS 0.007609f
C621 B.n564 VSUBS 0.007609f
C622 B.n565 VSUBS 0.007609f
C623 B.n566 VSUBS 0.007609f
C624 B.n567 VSUBS 0.007609f
C625 B.n568 VSUBS 0.007609f
C626 B.n569 VSUBS 0.007609f
C627 B.n570 VSUBS 0.007609f
C628 B.n571 VSUBS 0.007609f
C629 B.n572 VSUBS 0.007609f
C630 B.n573 VSUBS 0.007609f
C631 B.n574 VSUBS 0.007609f
C632 B.n575 VSUBS 0.007609f
C633 B.n576 VSUBS 0.007609f
C634 B.n577 VSUBS 0.007609f
C635 B.n578 VSUBS 0.007609f
C636 B.n579 VSUBS 0.007609f
C637 B.n580 VSUBS 0.007609f
C638 B.n581 VSUBS 0.007609f
C639 B.n582 VSUBS 0.007609f
C640 B.n583 VSUBS 0.007609f
C641 B.n584 VSUBS 0.007609f
C642 B.n585 VSUBS 0.007609f
C643 B.n586 VSUBS 0.007609f
C644 B.n587 VSUBS 0.007609f
C645 B.n588 VSUBS 0.007609f
C646 B.n589 VSUBS 0.007609f
C647 B.n590 VSUBS 0.007609f
C648 B.n591 VSUBS 0.007609f
C649 B.n592 VSUBS 0.007609f
C650 B.n593 VSUBS 0.007609f
C651 B.n594 VSUBS 0.007609f
C652 B.n595 VSUBS 0.007609f
C653 B.n596 VSUBS 0.007609f
C654 B.n597 VSUBS 0.007609f
C655 B.n598 VSUBS 0.007609f
C656 B.n599 VSUBS 0.007609f
C657 B.n600 VSUBS 0.007609f
C658 B.n601 VSUBS 0.007609f
C659 B.n602 VSUBS 0.007609f
C660 B.n603 VSUBS 0.007609f
C661 B.n604 VSUBS 0.007609f
C662 B.n605 VSUBS 0.007609f
C663 B.n606 VSUBS 0.007609f
C664 B.n607 VSUBS 0.007609f
C665 B.n608 VSUBS 0.007609f
C666 B.n609 VSUBS 0.007609f
C667 B.n610 VSUBS 0.007609f
C668 B.n611 VSUBS 0.007609f
C669 B.n612 VSUBS 0.007609f
C670 B.n613 VSUBS 0.007609f
C671 B.n614 VSUBS 0.007609f
C672 B.n615 VSUBS 0.007609f
C673 B.n616 VSUBS 0.018373f
C674 B.n617 VSUBS 0.01721f
C675 B.n618 VSUBS 0.01721f
C676 B.n619 VSUBS 0.007609f
C677 B.n620 VSUBS 0.007609f
C678 B.n621 VSUBS 0.007609f
C679 B.n622 VSUBS 0.007609f
C680 B.n623 VSUBS 0.007609f
C681 B.n624 VSUBS 0.007609f
C682 B.n625 VSUBS 0.007609f
C683 B.n626 VSUBS 0.007609f
C684 B.n627 VSUBS 0.007609f
C685 B.n628 VSUBS 0.007609f
C686 B.n629 VSUBS 0.007609f
C687 B.n630 VSUBS 0.007609f
C688 B.n631 VSUBS 0.007609f
C689 B.n632 VSUBS 0.007609f
C690 B.n633 VSUBS 0.007609f
C691 B.n634 VSUBS 0.007609f
C692 B.n635 VSUBS 0.007609f
C693 B.n636 VSUBS 0.007609f
C694 B.n637 VSUBS 0.007609f
C695 B.n638 VSUBS 0.007609f
C696 B.n639 VSUBS 0.007609f
C697 B.n640 VSUBS 0.007609f
C698 B.n641 VSUBS 0.007609f
C699 B.n642 VSUBS 0.007609f
C700 B.n643 VSUBS 0.009929f
C701 B.n644 VSUBS 0.010577f
C702 B.n645 VSUBS 0.021033f
C703 VTAIL.n0 VSUBS 0.023261f
C704 VTAIL.n1 VSUBS 0.022286f
C705 VTAIL.n2 VSUBS 0.011976f
C706 VTAIL.n3 VSUBS 0.028306f
C707 VTAIL.n4 VSUBS 0.01268f
C708 VTAIL.n5 VSUBS 0.022286f
C709 VTAIL.n6 VSUBS 0.011976f
C710 VTAIL.n7 VSUBS 0.028306f
C711 VTAIL.n8 VSUBS 0.01268f
C712 VTAIL.n9 VSUBS 0.022286f
C713 VTAIL.n10 VSUBS 0.011976f
C714 VTAIL.n11 VSUBS 0.028306f
C715 VTAIL.n12 VSUBS 0.01268f
C716 VTAIL.n13 VSUBS 0.022286f
C717 VTAIL.n14 VSUBS 0.011976f
C718 VTAIL.n15 VSUBS 0.028306f
C719 VTAIL.n16 VSUBS 0.01268f
C720 VTAIL.n17 VSUBS 0.022286f
C721 VTAIL.n18 VSUBS 0.011976f
C722 VTAIL.n19 VSUBS 0.028306f
C723 VTAIL.n20 VSUBS 0.01268f
C724 VTAIL.n21 VSUBS 0.022286f
C725 VTAIL.n22 VSUBS 0.011976f
C726 VTAIL.n23 VSUBS 0.028306f
C727 VTAIL.n24 VSUBS 0.01268f
C728 VTAIL.n25 VSUBS 0.022286f
C729 VTAIL.n26 VSUBS 0.011976f
C730 VTAIL.n27 VSUBS 0.028306f
C731 VTAIL.n28 VSUBS 0.01268f
C732 VTAIL.n29 VSUBS 0.168669f
C733 VTAIL.t7 VSUBS 0.060696f
C734 VTAIL.n30 VSUBS 0.02123f
C735 VTAIL.n31 VSUBS 0.018007f
C736 VTAIL.n32 VSUBS 0.011976f
C737 VTAIL.n33 VSUBS 1.6011f
C738 VTAIL.n34 VSUBS 0.022286f
C739 VTAIL.n35 VSUBS 0.011976f
C740 VTAIL.n36 VSUBS 0.01268f
C741 VTAIL.n37 VSUBS 0.028306f
C742 VTAIL.n38 VSUBS 0.028306f
C743 VTAIL.n39 VSUBS 0.01268f
C744 VTAIL.n40 VSUBS 0.011976f
C745 VTAIL.n41 VSUBS 0.022286f
C746 VTAIL.n42 VSUBS 0.022286f
C747 VTAIL.n43 VSUBS 0.011976f
C748 VTAIL.n44 VSUBS 0.01268f
C749 VTAIL.n45 VSUBS 0.028306f
C750 VTAIL.n46 VSUBS 0.028306f
C751 VTAIL.n47 VSUBS 0.01268f
C752 VTAIL.n48 VSUBS 0.011976f
C753 VTAIL.n49 VSUBS 0.022286f
C754 VTAIL.n50 VSUBS 0.022286f
C755 VTAIL.n51 VSUBS 0.011976f
C756 VTAIL.n52 VSUBS 0.01268f
C757 VTAIL.n53 VSUBS 0.028306f
C758 VTAIL.n54 VSUBS 0.028306f
C759 VTAIL.n55 VSUBS 0.01268f
C760 VTAIL.n56 VSUBS 0.011976f
C761 VTAIL.n57 VSUBS 0.022286f
C762 VTAIL.n58 VSUBS 0.022286f
C763 VTAIL.n59 VSUBS 0.011976f
C764 VTAIL.n60 VSUBS 0.01268f
C765 VTAIL.n61 VSUBS 0.028306f
C766 VTAIL.n62 VSUBS 0.028306f
C767 VTAIL.n63 VSUBS 0.01268f
C768 VTAIL.n64 VSUBS 0.011976f
C769 VTAIL.n65 VSUBS 0.022286f
C770 VTAIL.n66 VSUBS 0.022286f
C771 VTAIL.n67 VSUBS 0.011976f
C772 VTAIL.n68 VSUBS 0.01268f
C773 VTAIL.n69 VSUBS 0.028306f
C774 VTAIL.n70 VSUBS 0.028306f
C775 VTAIL.n71 VSUBS 0.028306f
C776 VTAIL.n72 VSUBS 0.01268f
C777 VTAIL.n73 VSUBS 0.011976f
C778 VTAIL.n74 VSUBS 0.022286f
C779 VTAIL.n75 VSUBS 0.022286f
C780 VTAIL.n76 VSUBS 0.011976f
C781 VTAIL.n77 VSUBS 0.012328f
C782 VTAIL.n78 VSUBS 0.012328f
C783 VTAIL.n79 VSUBS 0.028306f
C784 VTAIL.n80 VSUBS 0.028306f
C785 VTAIL.n81 VSUBS 0.01268f
C786 VTAIL.n82 VSUBS 0.011976f
C787 VTAIL.n83 VSUBS 0.022286f
C788 VTAIL.n84 VSUBS 0.022286f
C789 VTAIL.n85 VSUBS 0.011976f
C790 VTAIL.n86 VSUBS 0.01268f
C791 VTAIL.n87 VSUBS 0.028306f
C792 VTAIL.n88 VSUBS 0.064348f
C793 VTAIL.n89 VSUBS 0.01268f
C794 VTAIL.n90 VSUBS 0.011976f
C795 VTAIL.n91 VSUBS 0.050296f
C796 VTAIL.n92 VSUBS 0.032137f
C797 VTAIL.n93 VSUBS 0.0931f
C798 VTAIL.n94 VSUBS 0.023261f
C799 VTAIL.n95 VSUBS 0.022286f
C800 VTAIL.n96 VSUBS 0.011976f
C801 VTAIL.n97 VSUBS 0.028306f
C802 VTAIL.n98 VSUBS 0.01268f
C803 VTAIL.n99 VSUBS 0.022286f
C804 VTAIL.n100 VSUBS 0.011976f
C805 VTAIL.n101 VSUBS 0.028306f
C806 VTAIL.n102 VSUBS 0.01268f
C807 VTAIL.n103 VSUBS 0.022286f
C808 VTAIL.n104 VSUBS 0.011976f
C809 VTAIL.n105 VSUBS 0.028306f
C810 VTAIL.n106 VSUBS 0.01268f
C811 VTAIL.n107 VSUBS 0.022286f
C812 VTAIL.n108 VSUBS 0.011976f
C813 VTAIL.n109 VSUBS 0.028306f
C814 VTAIL.n110 VSUBS 0.01268f
C815 VTAIL.n111 VSUBS 0.022286f
C816 VTAIL.n112 VSUBS 0.011976f
C817 VTAIL.n113 VSUBS 0.028306f
C818 VTAIL.n114 VSUBS 0.01268f
C819 VTAIL.n115 VSUBS 0.022286f
C820 VTAIL.n116 VSUBS 0.011976f
C821 VTAIL.n117 VSUBS 0.028306f
C822 VTAIL.n118 VSUBS 0.01268f
C823 VTAIL.n119 VSUBS 0.022286f
C824 VTAIL.n120 VSUBS 0.011976f
C825 VTAIL.n121 VSUBS 0.028306f
C826 VTAIL.n122 VSUBS 0.01268f
C827 VTAIL.n123 VSUBS 0.168669f
C828 VTAIL.t2 VSUBS 0.060696f
C829 VTAIL.n124 VSUBS 0.02123f
C830 VTAIL.n125 VSUBS 0.018007f
C831 VTAIL.n126 VSUBS 0.011976f
C832 VTAIL.n127 VSUBS 1.6011f
C833 VTAIL.n128 VSUBS 0.022286f
C834 VTAIL.n129 VSUBS 0.011976f
C835 VTAIL.n130 VSUBS 0.01268f
C836 VTAIL.n131 VSUBS 0.028306f
C837 VTAIL.n132 VSUBS 0.028306f
C838 VTAIL.n133 VSUBS 0.01268f
C839 VTAIL.n134 VSUBS 0.011976f
C840 VTAIL.n135 VSUBS 0.022286f
C841 VTAIL.n136 VSUBS 0.022286f
C842 VTAIL.n137 VSUBS 0.011976f
C843 VTAIL.n138 VSUBS 0.01268f
C844 VTAIL.n139 VSUBS 0.028306f
C845 VTAIL.n140 VSUBS 0.028306f
C846 VTAIL.n141 VSUBS 0.01268f
C847 VTAIL.n142 VSUBS 0.011976f
C848 VTAIL.n143 VSUBS 0.022286f
C849 VTAIL.n144 VSUBS 0.022286f
C850 VTAIL.n145 VSUBS 0.011976f
C851 VTAIL.n146 VSUBS 0.01268f
C852 VTAIL.n147 VSUBS 0.028306f
C853 VTAIL.n148 VSUBS 0.028306f
C854 VTAIL.n149 VSUBS 0.01268f
C855 VTAIL.n150 VSUBS 0.011976f
C856 VTAIL.n151 VSUBS 0.022286f
C857 VTAIL.n152 VSUBS 0.022286f
C858 VTAIL.n153 VSUBS 0.011976f
C859 VTAIL.n154 VSUBS 0.01268f
C860 VTAIL.n155 VSUBS 0.028306f
C861 VTAIL.n156 VSUBS 0.028306f
C862 VTAIL.n157 VSUBS 0.01268f
C863 VTAIL.n158 VSUBS 0.011976f
C864 VTAIL.n159 VSUBS 0.022286f
C865 VTAIL.n160 VSUBS 0.022286f
C866 VTAIL.n161 VSUBS 0.011976f
C867 VTAIL.n162 VSUBS 0.01268f
C868 VTAIL.n163 VSUBS 0.028306f
C869 VTAIL.n164 VSUBS 0.028306f
C870 VTAIL.n165 VSUBS 0.028306f
C871 VTAIL.n166 VSUBS 0.01268f
C872 VTAIL.n167 VSUBS 0.011976f
C873 VTAIL.n168 VSUBS 0.022286f
C874 VTAIL.n169 VSUBS 0.022286f
C875 VTAIL.n170 VSUBS 0.011976f
C876 VTAIL.n171 VSUBS 0.012328f
C877 VTAIL.n172 VSUBS 0.012328f
C878 VTAIL.n173 VSUBS 0.028306f
C879 VTAIL.n174 VSUBS 0.028306f
C880 VTAIL.n175 VSUBS 0.01268f
C881 VTAIL.n176 VSUBS 0.011976f
C882 VTAIL.n177 VSUBS 0.022286f
C883 VTAIL.n178 VSUBS 0.022286f
C884 VTAIL.n179 VSUBS 0.011976f
C885 VTAIL.n180 VSUBS 0.01268f
C886 VTAIL.n181 VSUBS 0.028306f
C887 VTAIL.n182 VSUBS 0.064348f
C888 VTAIL.n183 VSUBS 0.01268f
C889 VTAIL.n184 VSUBS 0.011976f
C890 VTAIL.n185 VSUBS 0.050296f
C891 VTAIL.n186 VSUBS 0.032137f
C892 VTAIL.n187 VSUBS 0.125756f
C893 VTAIL.n188 VSUBS 0.023261f
C894 VTAIL.n189 VSUBS 0.022286f
C895 VTAIL.n190 VSUBS 0.011976f
C896 VTAIL.n191 VSUBS 0.028306f
C897 VTAIL.n192 VSUBS 0.01268f
C898 VTAIL.n193 VSUBS 0.022286f
C899 VTAIL.n194 VSUBS 0.011976f
C900 VTAIL.n195 VSUBS 0.028306f
C901 VTAIL.n196 VSUBS 0.01268f
C902 VTAIL.n197 VSUBS 0.022286f
C903 VTAIL.n198 VSUBS 0.011976f
C904 VTAIL.n199 VSUBS 0.028306f
C905 VTAIL.n200 VSUBS 0.01268f
C906 VTAIL.n201 VSUBS 0.022286f
C907 VTAIL.n202 VSUBS 0.011976f
C908 VTAIL.n203 VSUBS 0.028306f
C909 VTAIL.n204 VSUBS 0.01268f
C910 VTAIL.n205 VSUBS 0.022286f
C911 VTAIL.n206 VSUBS 0.011976f
C912 VTAIL.n207 VSUBS 0.028306f
C913 VTAIL.n208 VSUBS 0.01268f
C914 VTAIL.n209 VSUBS 0.022286f
C915 VTAIL.n210 VSUBS 0.011976f
C916 VTAIL.n211 VSUBS 0.028306f
C917 VTAIL.n212 VSUBS 0.01268f
C918 VTAIL.n213 VSUBS 0.022286f
C919 VTAIL.n214 VSUBS 0.011976f
C920 VTAIL.n215 VSUBS 0.028306f
C921 VTAIL.n216 VSUBS 0.01268f
C922 VTAIL.n217 VSUBS 0.168669f
C923 VTAIL.t3 VSUBS 0.060696f
C924 VTAIL.n218 VSUBS 0.02123f
C925 VTAIL.n219 VSUBS 0.018007f
C926 VTAIL.n220 VSUBS 0.011976f
C927 VTAIL.n221 VSUBS 1.6011f
C928 VTAIL.n222 VSUBS 0.022286f
C929 VTAIL.n223 VSUBS 0.011976f
C930 VTAIL.n224 VSUBS 0.01268f
C931 VTAIL.n225 VSUBS 0.028306f
C932 VTAIL.n226 VSUBS 0.028306f
C933 VTAIL.n227 VSUBS 0.01268f
C934 VTAIL.n228 VSUBS 0.011976f
C935 VTAIL.n229 VSUBS 0.022286f
C936 VTAIL.n230 VSUBS 0.022286f
C937 VTAIL.n231 VSUBS 0.011976f
C938 VTAIL.n232 VSUBS 0.01268f
C939 VTAIL.n233 VSUBS 0.028306f
C940 VTAIL.n234 VSUBS 0.028306f
C941 VTAIL.n235 VSUBS 0.01268f
C942 VTAIL.n236 VSUBS 0.011976f
C943 VTAIL.n237 VSUBS 0.022286f
C944 VTAIL.n238 VSUBS 0.022286f
C945 VTAIL.n239 VSUBS 0.011976f
C946 VTAIL.n240 VSUBS 0.01268f
C947 VTAIL.n241 VSUBS 0.028306f
C948 VTAIL.n242 VSUBS 0.028306f
C949 VTAIL.n243 VSUBS 0.01268f
C950 VTAIL.n244 VSUBS 0.011976f
C951 VTAIL.n245 VSUBS 0.022286f
C952 VTAIL.n246 VSUBS 0.022286f
C953 VTAIL.n247 VSUBS 0.011976f
C954 VTAIL.n248 VSUBS 0.01268f
C955 VTAIL.n249 VSUBS 0.028306f
C956 VTAIL.n250 VSUBS 0.028306f
C957 VTAIL.n251 VSUBS 0.01268f
C958 VTAIL.n252 VSUBS 0.011976f
C959 VTAIL.n253 VSUBS 0.022286f
C960 VTAIL.n254 VSUBS 0.022286f
C961 VTAIL.n255 VSUBS 0.011976f
C962 VTAIL.n256 VSUBS 0.01268f
C963 VTAIL.n257 VSUBS 0.028306f
C964 VTAIL.n258 VSUBS 0.028306f
C965 VTAIL.n259 VSUBS 0.028306f
C966 VTAIL.n260 VSUBS 0.01268f
C967 VTAIL.n261 VSUBS 0.011976f
C968 VTAIL.n262 VSUBS 0.022286f
C969 VTAIL.n263 VSUBS 0.022286f
C970 VTAIL.n264 VSUBS 0.011976f
C971 VTAIL.n265 VSUBS 0.012328f
C972 VTAIL.n266 VSUBS 0.012328f
C973 VTAIL.n267 VSUBS 0.028306f
C974 VTAIL.n268 VSUBS 0.028306f
C975 VTAIL.n269 VSUBS 0.01268f
C976 VTAIL.n270 VSUBS 0.011976f
C977 VTAIL.n271 VSUBS 0.022286f
C978 VTAIL.n272 VSUBS 0.022286f
C979 VTAIL.n273 VSUBS 0.011976f
C980 VTAIL.n274 VSUBS 0.01268f
C981 VTAIL.n275 VSUBS 0.028306f
C982 VTAIL.n276 VSUBS 0.064348f
C983 VTAIL.n277 VSUBS 0.01268f
C984 VTAIL.n278 VSUBS 0.011976f
C985 VTAIL.n279 VSUBS 0.050296f
C986 VTAIL.n280 VSUBS 0.032137f
C987 VTAIL.n281 VSUBS 1.50598f
C988 VTAIL.n282 VSUBS 0.023261f
C989 VTAIL.n283 VSUBS 0.022286f
C990 VTAIL.n284 VSUBS 0.011976f
C991 VTAIL.n285 VSUBS 0.028306f
C992 VTAIL.n286 VSUBS 0.01268f
C993 VTAIL.n287 VSUBS 0.022286f
C994 VTAIL.n288 VSUBS 0.011976f
C995 VTAIL.n289 VSUBS 0.028306f
C996 VTAIL.n290 VSUBS 0.01268f
C997 VTAIL.n291 VSUBS 0.022286f
C998 VTAIL.n292 VSUBS 0.011976f
C999 VTAIL.n293 VSUBS 0.028306f
C1000 VTAIL.n294 VSUBS 0.028306f
C1001 VTAIL.n295 VSUBS 0.01268f
C1002 VTAIL.n296 VSUBS 0.022286f
C1003 VTAIL.n297 VSUBS 0.011976f
C1004 VTAIL.n298 VSUBS 0.028306f
C1005 VTAIL.n299 VSUBS 0.01268f
C1006 VTAIL.n300 VSUBS 0.022286f
C1007 VTAIL.n301 VSUBS 0.011976f
C1008 VTAIL.n302 VSUBS 0.028306f
C1009 VTAIL.n303 VSUBS 0.01268f
C1010 VTAIL.n304 VSUBS 0.022286f
C1011 VTAIL.n305 VSUBS 0.011976f
C1012 VTAIL.n306 VSUBS 0.028306f
C1013 VTAIL.n307 VSUBS 0.01268f
C1014 VTAIL.n308 VSUBS 0.022286f
C1015 VTAIL.n309 VSUBS 0.011976f
C1016 VTAIL.n310 VSUBS 0.028306f
C1017 VTAIL.n311 VSUBS 0.01268f
C1018 VTAIL.n312 VSUBS 0.168669f
C1019 VTAIL.t5 VSUBS 0.060696f
C1020 VTAIL.n313 VSUBS 0.02123f
C1021 VTAIL.n314 VSUBS 0.018007f
C1022 VTAIL.n315 VSUBS 0.011976f
C1023 VTAIL.n316 VSUBS 1.6011f
C1024 VTAIL.n317 VSUBS 0.022286f
C1025 VTAIL.n318 VSUBS 0.011976f
C1026 VTAIL.n319 VSUBS 0.01268f
C1027 VTAIL.n320 VSUBS 0.028306f
C1028 VTAIL.n321 VSUBS 0.028306f
C1029 VTAIL.n322 VSUBS 0.01268f
C1030 VTAIL.n323 VSUBS 0.011976f
C1031 VTAIL.n324 VSUBS 0.022286f
C1032 VTAIL.n325 VSUBS 0.022286f
C1033 VTAIL.n326 VSUBS 0.011976f
C1034 VTAIL.n327 VSUBS 0.01268f
C1035 VTAIL.n328 VSUBS 0.028306f
C1036 VTAIL.n329 VSUBS 0.028306f
C1037 VTAIL.n330 VSUBS 0.01268f
C1038 VTAIL.n331 VSUBS 0.011976f
C1039 VTAIL.n332 VSUBS 0.022286f
C1040 VTAIL.n333 VSUBS 0.022286f
C1041 VTAIL.n334 VSUBS 0.011976f
C1042 VTAIL.n335 VSUBS 0.01268f
C1043 VTAIL.n336 VSUBS 0.028306f
C1044 VTAIL.n337 VSUBS 0.028306f
C1045 VTAIL.n338 VSUBS 0.01268f
C1046 VTAIL.n339 VSUBS 0.011976f
C1047 VTAIL.n340 VSUBS 0.022286f
C1048 VTAIL.n341 VSUBS 0.022286f
C1049 VTAIL.n342 VSUBS 0.011976f
C1050 VTAIL.n343 VSUBS 0.01268f
C1051 VTAIL.n344 VSUBS 0.028306f
C1052 VTAIL.n345 VSUBS 0.028306f
C1053 VTAIL.n346 VSUBS 0.01268f
C1054 VTAIL.n347 VSUBS 0.011976f
C1055 VTAIL.n348 VSUBS 0.022286f
C1056 VTAIL.n349 VSUBS 0.022286f
C1057 VTAIL.n350 VSUBS 0.011976f
C1058 VTAIL.n351 VSUBS 0.01268f
C1059 VTAIL.n352 VSUBS 0.028306f
C1060 VTAIL.n353 VSUBS 0.028306f
C1061 VTAIL.n354 VSUBS 0.01268f
C1062 VTAIL.n355 VSUBS 0.011976f
C1063 VTAIL.n356 VSUBS 0.022286f
C1064 VTAIL.n357 VSUBS 0.022286f
C1065 VTAIL.n358 VSUBS 0.011976f
C1066 VTAIL.n359 VSUBS 0.012328f
C1067 VTAIL.n360 VSUBS 0.012328f
C1068 VTAIL.n361 VSUBS 0.028306f
C1069 VTAIL.n362 VSUBS 0.028306f
C1070 VTAIL.n363 VSUBS 0.01268f
C1071 VTAIL.n364 VSUBS 0.011976f
C1072 VTAIL.n365 VSUBS 0.022286f
C1073 VTAIL.n366 VSUBS 0.022286f
C1074 VTAIL.n367 VSUBS 0.011976f
C1075 VTAIL.n368 VSUBS 0.01268f
C1076 VTAIL.n369 VSUBS 0.028306f
C1077 VTAIL.n370 VSUBS 0.064348f
C1078 VTAIL.n371 VSUBS 0.01268f
C1079 VTAIL.n372 VSUBS 0.011976f
C1080 VTAIL.n373 VSUBS 0.050296f
C1081 VTAIL.n374 VSUBS 0.032137f
C1082 VTAIL.n375 VSUBS 1.50598f
C1083 VTAIL.n376 VSUBS 0.023261f
C1084 VTAIL.n377 VSUBS 0.022286f
C1085 VTAIL.n378 VSUBS 0.011976f
C1086 VTAIL.n379 VSUBS 0.028306f
C1087 VTAIL.n380 VSUBS 0.01268f
C1088 VTAIL.n381 VSUBS 0.022286f
C1089 VTAIL.n382 VSUBS 0.011976f
C1090 VTAIL.n383 VSUBS 0.028306f
C1091 VTAIL.n384 VSUBS 0.01268f
C1092 VTAIL.n385 VSUBS 0.022286f
C1093 VTAIL.n386 VSUBS 0.011976f
C1094 VTAIL.n387 VSUBS 0.028306f
C1095 VTAIL.n388 VSUBS 0.028306f
C1096 VTAIL.n389 VSUBS 0.01268f
C1097 VTAIL.n390 VSUBS 0.022286f
C1098 VTAIL.n391 VSUBS 0.011976f
C1099 VTAIL.n392 VSUBS 0.028306f
C1100 VTAIL.n393 VSUBS 0.01268f
C1101 VTAIL.n394 VSUBS 0.022286f
C1102 VTAIL.n395 VSUBS 0.011976f
C1103 VTAIL.n396 VSUBS 0.028306f
C1104 VTAIL.n397 VSUBS 0.01268f
C1105 VTAIL.n398 VSUBS 0.022286f
C1106 VTAIL.n399 VSUBS 0.011976f
C1107 VTAIL.n400 VSUBS 0.028306f
C1108 VTAIL.n401 VSUBS 0.01268f
C1109 VTAIL.n402 VSUBS 0.022286f
C1110 VTAIL.n403 VSUBS 0.011976f
C1111 VTAIL.n404 VSUBS 0.028306f
C1112 VTAIL.n405 VSUBS 0.01268f
C1113 VTAIL.n406 VSUBS 0.168669f
C1114 VTAIL.t6 VSUBS 0.060696f
C1115 VTAIL.n407 VSUBS 0.02123f
C1116 VTAIL.n408 VSUBS 0.018007f
C1117 VTAIL.n409 VSUBS 0.011976f
C1118 VTAIL.n410 VSUBS 1.6011f
C1119 VTAIL.n411 VSUBS 0.022286f
C1120 VTAIL.n412 VSUBS 0.011976f
C1121 VTAIL.n413 VSUBS 0.01268f
C1122 VTAIL.n414 VSUBS 0.028306f
C1123 VTAIL.n415 VSUBS 0.028306f
C1124 VTAIL.n416 VSUBS 0.01268f
C1125 VTAIL.n417 VSUBS 0.011976f
C1126 VTAIL.n418 VSUBS 0.022286f
C1127 VTAIL.n419 VSUBS 0.022286f
C1128 VTAIL.n420 VSUBS 0.011976f
C1129 VTAIL.n421 VSUBS 0.01268f
C1130 VTAIL.n422 VSUBS 0.028306f
C1131 VTAIL.n423 VSUBS 0.028306f
C1132 VTAIL.n424 VSUBS 0.01268f
C1133 VTAIL.n425 VSUBS 0.011976f
C1134 VTAIL.n426 VSUBS 0.022286f
C1135 VTAIL.n427 VSUBS 0.022286f
C1136 VTAIL.n428 VSUBS 0.011976f
C1137 VTAIL.n429 VSUBS 0.01268f
C1138 VTAIL.n430 VSUBS 0.028306f
C1139 VTAIL.n431 VSUBS 0.028306f
C1140 VTAIL.n432 VSUBS 0.01268f
C1141 VTAIL.n433 VSUBS 0.011976f
C1142 VTAIL.n434 VSUBS 0.022286f
C1143 VTAIL.n435 VSUBS 0.022286f
C1144 VTAIL.n436 VSUBS 0.011976f
C1145 VTAIL.n437 VSUBS 0.01268f
C1146 VTAIL.n438 VSUBS 0.028306f
C1147 VTAIL.n439 VSUBS 0.028306f
C1148 VTAIL.n440 VSUBS 0.01268f
C1149 VTAIL.n441 VSUBS 0.011976f
C1150 VTAIL.n442 VSUBS 0.022286f
C1151 VTAIL.n443 VSUBS 0.022286f
C1152 VTAIL.n444 VSUBS 0.011976f
C1153 VTAIL.n445 VSUBS 0.01268f
C1154 VTAIL.n446 VSUBS 0.028306f
C1155 VTAIL.n447 VSUBS 0.028306f
C1156 VTAIL.n448 VSUBS 0.01268f
C1157 VTAIL.n449 VSUBS 0.011976f
C1158 VTAIL.n450 VSUBS 0.022286f
C1159 VTAIL.n451 VSUBS 0.022286f
C1160 VTAIL.n452 VSUBS 0.011976f
C1161 VTAIL.n453 VSUBS 0.012328f
C1162 VTAIL.n454 VSUBS 0.012328f
C1163 VTAIL.n455 VSUBS 0.028306f
C1164 VTAIL.n456 VSUBS 0.028306f
C1165 VTAIL.n457 VSUBS 0.01268f
C1166 VTAIL.n458 VSUBS 0.011976f
C1167 VTAIL.n459 VSUBS 0.022286f
C1168 VTAIL.n460 VSUBS 0.022286f
C1169 VTAIL.n461 VSUBS 0.011976f
C1170 VTAIL.n462 VSUBS 0.01268f
C1171 VTAIL.n463 VSUBS 0.028306f
C1172 VTAIL.n464 VSUBS 0.064348f
C1173 VTAIL.n465 VSUBS 0.01268f
C1174 VTAIL.n466 VSUBS 0.011976f
C1175 VTAIL.n467 VSUBS 0.050296f
C1176 VTAIL.n468 VSUBS 0.032137f
C1177 VTAIL.n469 VSUBS 0.125756f
C1178 VTAIL.n470 VSUBS 0.023261f
C1179 VTAIL.n471 VSUBS 0.022286f
C1180 VTAIL.n472 VSUBS 0.011976f
C1181 VTAIL.n473 VSUBS 0.028306f
C1182 VTAIL.n474 VSUBS 0.01268f
C1183 VTAIL.n475 VSUBS 0.022286f
C1184 VTAIL.n476 VSUBS 0.011976f
C1185 VTAIL.n477 VSUBS 0.028306f
C1186 VTAIL.n478 VSUBS 0.01268f
C1187 VTAIL.n479 VSUBS 0.022286f
C1188 VTAIL.n480 VSUBS 0.011976f
C1189 VTAIL.n481 VSUBS 0.028306f
C1190 VTAIL.n482 VSUBS 0.028306f
C1191 VTAIL.n483 VSUBS 0.01268f
C1192 VTAIL.n484 VSUBS 0.022286f
C1193 VTAIL.n485 VSUBS 0.011976f
C1194 VTAIL.n486 VSUBS 0.028306f
C1195 VTAIL.n487 VSUBS 0.01268f
C1196 VTAIL.n488 VSUBS 0.022286f
C1197 VTAIL.n489 VSUBS 0.011976f
C1198 VTAIL.n490 VSUBS 0.028306f
C1199 VTAIL.n491 VSUBS 0.01268f
C1200 VTAIL.n492 VSUBS 0.022286f
C1201 VTAIL.n493 VSUBS 0.011976f
C1202 VTAIL.n494 VSUBS 0.028306f
C1203 VTAIL.n495 VSUBS 0.01268f
C1204 VTAIL.n496 VSUBS 0.022286f
C1205 VTAIL.n497 VSUBS 0.011976f
C1206 VTAIL.n498 VSUBS 0.028306f
C1207 VTAIL.n499 VSUBS 0.01268f
C1208 VTAIL.n500 VSUBS 0.168669f
C1209 VTAIL.t0 VSUBS 0.060696f
C1210 VTAIL.n501 VSUBS 0.02123f
C1211 VTAIL.n502 VSUBS 0.018007f
C1212 VTAIL.n503 VSUBS 0.011976f
C1213 VTAIL.n504 VSUBS 1.6011f
C1214 VTAIL.n505 VSUBS 0.022286f
C1215 VTAIL.n506 VSUBS 0.011976f
C1216 VTAIL.n507 VSUBS 0.01268f
C1217 VTAIL.n508 VSUBS 0.028306f
C1218 VTAIL.n509 VSUBS 0.028306f
C1219 VTAIL.n510 VSUBS 0.01268f
C1220 VTAIL.n511 VSUBS 0.011976f
C1221 VTAIL.n512 VSUBS 0.022286f
C1222 VTAIL.n513 VSUBS 0.022286f
C1223 VTAIL.n514 VSUBS 0.011976f
C1224 VTAIL.n515 VSUBS 0.01268f
C1225 VTAIL.n516 VSUBS 0.028306f
C1226 VTAIL.n517 VSUBS 0.028306f
C1227 VTAIL.n518 VSUBS 0.01268f
C1228 VTAIL.n519 VSUBS 0.011976f
C1229 VTAIL.n520 VSUBS 0.022286f
C1230 VTAIL.n521 VSUBS 0.022286f
C1231 VTAIL.n522 VSUBS 0.011976f
C1232 VTAIL.n523 VSUBS 0.01268f
C1233 VTAIL.n524 VSUBS 0.028306f
C1234 VTAIL.n525 VSUBS 0.028306f
C1235 VTAIL.n526 VSUBS 0.01268f
C1236 VTAIL.n527 VSUBS 0.011976f
C1237 VTAIL.n528 VSUBS 0.022286f
C1238 VTAIL.n529 VSUBS 0.022286f
C1239 VTAIL.n530 VSUBS 0.011976f
C1240 VTAIL.n531 VSUBS 0.01268f
C1241 VTAIL.n532 VSUBS 0.028306f
C1242 VTAIL.n533 VSUBS 0.028306f
C1243 VTAIL.n534 VSUBS 0.01268f
C1244 VTAIL.n535 VSUBS 0.011976f
C1245 VTAIL.n536 VSUBS 0.022286f
C1246 VTAIL.n537 VSUBS 0.022286f
C1247 VTAIL.n538 VSUBS 0.011976f
C1248 VTAIL.n539 VSUBS 0.01268f
C1249 VTAIL.n540 VSUBS 0.028306f
C1250 VTAIL.n541 VSUBS 0.028306f
C1251 VTAIL.n542 VSUBS 0.01268f
C1252 VTAIL.n543 VSUBS 0.011976f
C1253 VTAIL.n544 VSUBS 0.022286f
C1254 VTAIL.n545 VSUBS 0.022286f
C1255 VTAIL.n546 VSUBS 0.011976f
C1256 VTAIL.n547 VSUBS 0.012328f
C1257 VTAIL.n548 VSUBS 0.012328f
C1258 VTAIL.n549 VSUBS 0.028306f
C1259 VTAIL.n550 VSUBS 0.028306f
C1260 VTAIL.n551 VSUBS 0.01268f
C1261 VTAIL.n552 VSUBS 0.011976f
C1262 VTAIL.n553 VSUBS 0.022286f
C1263 VTAIL.n554 VSUBS 0.022286f
C1264 VTAIL.n555 VSUBS 0.011976f
C1265 VTAIL.n556 VSUBS 0.01268f
C1266 VTAIL.n557 VSUBS 0.028306f
C1267 VTAIL.n558 VSUBS 0.064348f
C1268 VTAIL.n559 VSUBS 0.01268f
C1269 VTAIL.n560 VSUBS 0.011976f
C1270 VTAIL.n561 VSUBS 0.050296f
C1271 VTAIL.n562 VSUBS 0.032137f
C1272 VTAIL.n563 VSUBS 0.125756f
C1273 VTAIL.n564 VSUBS 0.023261f
C1274 VTAIL.n565 VSUBS 0.022286f
C1275 VTAIL.n566 VSUBS 0.011976f
C1276 VTAIL.n567 VSUBS 0.028306f
C1277 VTAIL.n568 VSUBS 0.01268f
C1278 VTAIL.n569 VSUBS 0.022286f
C1279 VTAIL.n570 VSUBS 0.011976f
C1280 VTAIL.n571 VSUBS 0.028306f
C1281 VTAIL.n572 VSUBS 0.01268f
C1282 VTAIL.n573 VSUBS 0.022286f
C1283 VTAIL.n574 VSUBS 0.011976f
C1284 VTAIL.n575 VSUBS 0.028306f
C1285 VTAIL.n576 VSUBS 0.028306f
C1286 VTAIL.n577 VSUBS 0.01268f
C1287 VTAIL.n578 VSUBS 0.022286f
C1288 VTAIL.n579 VSUBS 0.011976f
C1289 VTAIL.n580 VSUBS 0.028306f
C1290 VTAIL.n581 VSUBS 0.01268f
C1291 VTAIL.n582 VSUBS 0.022286f
C1292 VTAIL.n583 VSUBS 0.011976f
C1293 VTAIL.n584 VSUBS 0.028306f
C1294 VTAIL.n585 VSUBS 0.01268f
C1295 VTAIL.n586 VSUBS 0.022286f
C1296 VTAIL.n587 VSUBS 0.011976f
C1297 VTAIL.n588 VSUBS 0.028306f
C1298 VTAIL.n589 VSUBS 0.01268f
C1299 VTAIL.n590 VSUBS 0.022286f
C1300 VTAIL.n591 VSUBS 0.011976f
C1301 VTAIL.n592 VSUBS 0.028306f
C1302 VTAIL.n593 VSUBS 0.01268f
C1303 VTAIL.n594 VSUBS 0.168669f
C1304 VTAIL.t1 VSUBS 0.060696f
C1305 VTAIL.n595 VSUBS 0.02123f
C1306 VTAIL.n596 VSUBS 0.018007f
C1307 VTAIL.n597 VSUBS 0.011976f
C1308 VTAIL.n598 VSUBS 1.6011f
C1309 VTAIL.n599 VSUBS 0.022286f
C1310 VTAIL.n600 VSUBS 0.011976f
C1311 VTAIL.n601 VSUBS 0.01268f
C1312 VTAIL.n602 VSUBS 0.028306f
C1313 VTAIL.n603 VSUBS 0.028306f
C1314 VTAIL.n604 VSUBS 0.01268f
C1315 VTAIL.n605 VSUBS 0.011976f
C1316 VTAIL.n606 VSUBS 0.022286f
C1317 VTAIL.n607 VSUBS 0.022286f
C1318 VTAIL.n608 VSUBS 0.011976f
C1319 VTAIL.n609 VSUBS 0.01268f
C1320 VTAIL.n610 VSUBS 0.028306f
C1321 VTAIL.n611 VSUBS 0.028306f
C1322 VTAIL.n612 VSUBS 0.01268f
C1323 VTAIL.n613 VSUBS 0.011976f
C1324 VTAIL.n614 VSUBS 0.022286f
C1325 VTAIL.n615 VSUBS 0.022286f
C1326 VTAIL.n616 VSUBS 0.011976f
C1327 VTAIL.n617 VSUBS 0.01268f
C1328 VTAIL.n618 VSUBS 0.028306f
C1329 VTAIL.n619 VSUBS 0.028306f
C1330 VTAIL.n620 VSUBS 0.01268f
C1331 VTAIL.n621 VSUBS 0.011976f
C1332 VTAIL.n622 VSUBS 0.022286f
C1333 VTAIL.n623 VSUBS 0.022286f
C1334 VTAIL.n624 VSUBS 0.011976f
C1335 VTAIL.n625 VSUBS 0.01268f
C1336 VTAIL.n626 VSUBS 0.028306f
C1337 VTAIL.n627 VSUBS 0.028306f
C1338 VTAIL.n628 VSUBS 0.01268f
C1339 VTAIL.n629 VSUBS 0.011976f
C1340 VTAIL.n630 VSUBS 0.022286f
C1341 VTAIL.n631 VSUBS 0.022286f
C1342 VTAIL.n632 VSUBS 0.011976f
C1343 VTAIL.n633 VSUBS 0.01268f
C1344 VTAIL.n634 VSUBS 0.028306f
C1345 VTAIL.n635 VSUBS 0.028306f
C1346 VTAIL.n636 VSUBS 0.01268f
C1347 VTAIL.n637 VSUBS 0.011976f
C1348 VTAIL.n638 VSUBS 0.022286f
C1349 VTAIL.n639 VSUBS 0.022286f
C1350 VTAIL.n640 VSUBS 0.011976f
C1351 VTAIL.n641 VSUBS 0.012328f
C1352 VTAIL.n642 VSUBS 0.012328f
C1353 VTAIL.n643 VSUBS 0.028306f
C1354 VTAIL.n644 VSUBS 0.028306f
C1355 VTAIL.n645 VSUBS 0.01268f
C1356 VTAIL.n646 VSUBS 0.011976f
C1357 VTAIL.n647 VSUBS 0.022286f
C1358 VTAIL.n648 VSUBS 0.022286f
C1359 VTAIL.n649 VSUBS 0.011976f
C1360 VTAIL.n650 VSUBS 0.01268f
C1361 VTAIL.n651 VSUBS 0.028306f
C1362 VTAIL.n652 VSUBS 0.064348f
C1363 VTAIL.n653 VSUBS 0.01268f
C1364 VTAIL.n654 VSUBS 0.011976f
C1365 VTAIL.n655 VSUBS 0.050296f
C1366 VTAIL.n656 VSUBS 0.032137f
C1367 VTAIL.n657 VSUBS 1.50598f
C1368 VTAIL.n658 VSUBS 0.023261f
C1369 VTAIL.n659 VSUBS 0.022286f
C1370 VTAIL.n660 VSUBS 0.011976f
C1371 VTAIL.n661 VSUBS 0.028306f
C1372 VTAIL.n662 VSUBS 0.01268f
C1373 VTAIL.n663 VSUBS 0.022286f
C1374 VTAIL.n664 VSUBS 0.011976f
C1375 VTAIL.n665 VSUBS 0.028306f
C1376 VTAIL.n666 VSUBS 0.01268f
C1377 VTAIL.n667 VSUBS 0.022286f
C1378 VTAIL.n668 VSUBS 0.011976f
C1379 VTAIL.n669 VSUBS 0.028306f
C1380 VTAIL.n670 VSUBS 0.01268f
C1381 VTAIL.n671 VSUBS 0.022286f
C1382 VTAIL.n672 VSUBS 0.011976f
C1383 VTAIL.n673 VSUBS 0.028306f
C1384 VTAIL.n674 VSUBS 0.01268f
C1385 VTAIL.n675 VSUBS 0.022286f
C1386 VTAIL.n676 VSUBS 0.011976f
C1387 VTAIL.n677 VSUBS 0.028306f
C1388 VTAIL.n678 VSUBS 0.01268f
C1389 VTAIL.n679 VSUBS 0.022286f
C1390 VTAIL.n680 VSUBS 0.011976f
C1391 VTAIL.n681 VSUBS 0.028306f
C1392 VTAIL.n682 VSUBS 0.01268f
C1393 VTAIL.n683 VSUBS 0.022286f
C1394 VTAIL.n684 VSUBS 0.011976f
C1395 VTAIL.n685 VSUBS 0.028306f
C1396 VTAIL.n686 VSUBS 0.01268f
C1397 VTAIL.n687 VSUBS 0.168669f
C1398 VTAIL.t4 VSUBS 0.060696f
C1399 VTAIL.n688 VSUBS 0.02123f
C1400 VTAIL.n689 VSUBS 0.018007f
C1401 VTAIL.n690 VSUBS 0.011976f
C1402 VTAIL.n691 VSUBS 1.6011f
C1403 VTAIL.n692 VSUBS 0.022286f
C1404 VTAIL.n693 VSUBS 0.011976f
C1405 VTAIL.n694 VSUBS 0.01268f
C1406 VTAIL.n695 VSUBS 0.028306f
C1407 VTAIL.n696 VSUBS 0.028306f
C1408 VTAIL.n697 VSUBS 0.01268f
C1409 VTAIL.n698 VSUBS 0.011976f
C1410 VTAIL.n699 VSUBS 0.022286f
C1411 VTAIL.n700 VSUBS 0.022286f
C1412 VTAIL.n701 VSUBS 0.011976f
C1413 VTAIL.n702 VSUBS 0.01268f
C1414 VTAIL.n703 VSUBS 0.028306f
C1415 VTAIL.n704 VSUBS 0.028306f
C1416 VTAIL.n705 VSUBS 0.01268f
C1417 VTAIL.n706 VSUBS 0.011976f
C1418 VTAIL.n707 VSUBS 0.022286f
C1419 VTAIL.n708 VSUBS 0.022286f
C1420 VTAIL.n709 VSUBS 0.011976f
C1421 VTAIL.n710 VSUBS 0.01268f
C1422 VTAIL.n711 VSUBS 0.028306f
C1423 VTAIL.n712 VSUBS 0.028306f
C1424 VTAIL.n713 VSUBS 0.01268f
C1425 VTAIL.n714 VSUBS 0.011976f
C1426 VTAIL.n715 VSUBS 0.022286f
C1427 VTAIL.n716 VSUBS 0.022286f
C1428 VTAIL.n717 VSUBS 0.011976f
C1429 VTAIL.n718 VSUBS 0.01268f
C1430 VTAIL.n719 VSUBS 0.028306f
C1431 VTAIL.n720 VSUBS 0.028306f
C1432 VTAIL.n721 VSUBS 0.01268f
C1433 VTAIL.n722 VSUBS 0.011976f
C1434 VTAIL.n723 VSUBS 0.022286f
C1435 VTAIL.n724 VSUBS 0.022286f
C1436 VTAIL.n725 VSUBS 0.011976f
C1437 VTAIL.n726 VSUBS 0.01268f
C1438 VTAIL.n727 VSUBS 0.028306f
C1439 VTAIL.n728 VSUBS 0.028306f
C1440 VTAIL.n729 VSUBS 0.028306f
C1441 VTAIL.n730 VSUBS 0.01268f
C1442 VTAIL.n731 VSUBS 0.011976f
C1443 VTAIL.n732 VSUBS 0.022286f
C1444 VTAIL.n733 VSUBS 0.022286f
C1445 VTAIL.n734 VSUBS 0.011976f
C1446 VTAIL.n735 VSUBS 0.012328f
C1447 VTAIL.n736 VSUBS 0.012328f
C1448 VTAIL.n737 VSUBS 0.028306f
C1449 VTAIL.n738 VSUBS 0.028306f
C1450 VTAIL.n739 VSUBS 0.01268f
C1451 VTAIL.n740 VSUBS 0.011976f
C1452 VTAIL.n741 VSUBS 0.022286f
C1453 VTAIL.n742 VSUBS 0.022286f
C1454 VTAIL.n743 VSUBS 0.011976f
C1455 VTAIL.n744 VSUBS 0.01268f
C1456 VTAIL.n745 VSUBS 0.028306f
C1457 VTAIL.n746 VSUBS 0.064348f
C1458 VTAIL.n747 VSUBS 0.01268f
C1459 VTAIL.n748 VSUBS 0.011976f
C1460 VTAIL.n749 VSUBS 0.050296f
C1461 VTAIL.n750 VSUBS 0.032137f
C1462 VTAIL.n751 VSUBS 1.46496f
C1463 VDD2.t0 VSUBS 0.366795f
C1464 VDD2.t2 VSUBS 0.366795f
C1465 VDD2.n0 VSUBS 3.86139f
C1466 VDD2.t3 VSUBS 0.366795f
C1467 VDD2.t1 VSUBS 0.366795f
C1468 VDD2.n1 VSUBS 3.01558f
C1469 VDD2.n2 VSUBS 4.55835f
C1470 VN.t0 VSUBS 2.21761f
C1471 VN.t3 VSUBS 2.21753f
C1472 VN.n0 VSUBS 1.59775f
C1473 VN.t1 VSUBS 2.21761f
C1474 VN.t2 VSUBS 2.21753f
C1475 VN.n1 VSUBS 2.89911f
.ends

