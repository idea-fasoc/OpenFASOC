* NGSPICE file created from diff_pair_sample_1586.ext - technology: sky130A

.subckt diff_pair_sample_1586 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=0 ps=0 w=15.41 l=1.86
X1 VDD1.t1 VP.t0 VTAIL.t3 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=6.0099 ps=31.6 w=15.41 l=1.86
X2 B.t8 B.t6 B.t7 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=0 ps=0 w=15.41 l=1.86
X3 B.t5 B.t3 B.t4 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=0 ps=0 w=15.41 l=1.86
X4 VDD2.t1 VN.t0 VTAIL.t1 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=6.0099 ps=31.6 w=15.41 l=1.86
X5 B.t2 B.t0 B.t1 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=0 ps=0 w=15.41 l=1.86
X6 VDD1.t0 VP.t1 VTAIL.t2 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=6.0099 ps=31.6 w=15.41 l=1.86
X7 VDD2.t0 VN.t1 VTAIL.t0 w_n1846_n4050# sky130_fd_pr__pfet_01v8 ad=6.0099 pd=31.6 as=6.0099 ps=31.6 w=15.41 l=1.86
R0 B.n433 B.n432 585
R1 B.n434 B.n73 585
R2 B.n436 B.n435 585
R3 B.n437 B.n72 585
R4 B.n439 B.n438 585
R5 B.n440 B.n71 585
R6 B.n442 B.n441 585
R7 B.n443 B.n70 585
R8 B.n445 B.n444 585
R9 B.n446 B.n69 585
R10 B.n448 B.n447 585
R11 B.n449 B.n68 585
R12 B.n451 B.n450 585
R13 B.n452 B.n67 585
R14 B.n454 B.n453 585
R15 B.n455 B.n66 585
R16 B.n457 B.n456 585
R17 B.n458 B.n65 585
R18 B.n460 B.n459 585
R19 B.n461 B.n64 585
R20 B.n463 B.n462 585
R21 B.n464 B.n63 585
R22 B.n466 B.n465 585
R23 B.n467 B.n62 585
R24 B.n469 B.n468 585
R25 B.n470 B.n61 585
R26 B.n472 B.n471 585
R27 B.n473 B.n60 585
R28 B.n475 B.n474 585
R29 B.n476 B.n59 585
R30 B.n478 B.n477 585
R31 B.n479 B.n58 585
R32 B.n481 B.n480 585
R33 B.n482 B.n57 585
R34 B.n484 B.n483 585
R35 B.n485 B.n56 585
R36 B.n487 B.n486 585
R37 B.n488 B.n55 585
R38 B.n490 B.n489 585
R39 B.n491 B.n54 585
R40 B.n493 B.n492 585
R41 B.n494 B.n53 585
R42 B.n496 B.n495 585
R43 B.n497 B.n52 585
R44 B.n499 B.n498 585
R45 B.n500 B.n51 585
R46 B.n502 B.n501 585
R47 B.n503 B.n50 585
R48 B.n505 B.n504 585
R49 B.n506 B.n49 585
R50 B.n508 B.n507 585
R51 B.n509 B.n46 585
R52 B.n512 B.n511 585
R53 B.n513 B.n45 585
R54 B.n515 B.n514 585
R55 B.n516 B.n44 585
R56 B.n518 B.n517 585
R57 B.n519 B.n43 585
R58 B.n521 B.n520 585
R59 B.n522 B.n39 585
R60 B.n524 B.n523 585
R61 B.n525 B.n38 585
R62 B.n527 B.n526 585
R63 B.n528 B.n37 585
R64 B.n530 B.n529 585
R65 B.n531 B.n36 585
R66 B.n533 B.n532 585
R67 B.n534 B.n35 585
R68 B.n536 B.n535 585
R69 B.n537 B.n34 585
R70 B.n539 B.n538 585
R71 B.n540 B.n33 585
R72 B.n542 B.n541 585
R73 B.n543 B.n32 585
R74 B.n545 B.n544 585
R75 B.n546 B.n31 585
R76 B.n548 B.n547 585
R77 B.n549 B.n30 585
R78 B.n551 B.n550 585
R79 B.n552 B.n29 585
R80 B.n554 B.n553 585
R81 B.n555 B.n28 585
R82 B.n557 B.n556 585
R83 B.n558 B.n27 585
R84 B.n560 B.n559 585
R85 B.n561 B.n26 585
R86 B.n563 B.n562 585
R87 B.n564 B.n25 585
R88 B.n566 B.n565 585
R89 B.n567 B.n24 585
R90 B.n569 B.n568 585
R91 B.n570 B.n23 585
R92 B.n572 B.n571 585
R93 B.n573 B.n22 585
R94 B.n575 B.n574 585
R95 B.n576 B.n21 585
R96 B.n578 B.n577 585
R97 B.n579 B.n20 585
R98 B.n581 B.n580 585
R99 B.n582 B.n19 585
R100 B.n584 B.n583 585
R101 B.n585 B.n18 585
R102 B.n587 B.n586 585
R103 B.n588 B.n17 585
R104 B.n590 B.n589 585
R105 B.n591 B.n16 585
R106 B.n593 B.n592 585
R107 B.n594 B.n15 585
R108 B.n596 B.n595 585
R109 B.n597 B.n14 585
R110 B.n599 B.n598 585
R111 B.n600 B.n13 585
R112 B.n602 B.n601 585
R113 B.n431 B.n74 585
R114 B.n430 B.n429 585
R115 B.n428 B.n75 585
R116 B.n427 B.n426 585
R117 B.n425 B.n76 585
R118 B.n424 B.n423 585
R119 B.n422 B.n77 585
R120 B.n421 B.n420 585
R121 B.n419 B.n78 585
R122 B.n418 B.n417 585
R123 B.n416 B.n79 585
R124 B.n415 B.n414 585
R125 B.n413 B.n80 585
R126 B.n412 B.n411 585
R127 B.n410 B.n81 585
R128 B.n409 B.n408 585
R129 B.n407 B.n82 585
R130 B.n406 B.n405 585
R131 B.n404 B.n83 585
R132 B.n403 B.n402 585
R133 B.n401 B.n84 585
R134 B.n400 B.n399 585
R135 B.n398 B.n85 585
R136 B.n397 B.n396 585
R137 B.n395 B.n86 585
R138 B.n394 B.n393 585
R139 B.n392 B.n87 585
R140 B.n391 B.n390 585
R141 B.n389 B.n88 585
R142 B.n388 B.n387 585
R143 B.n386 B.n89 585
R144 B.n385 B.n384 585
R145 B.n383 B.n90 585
R146 B.n382 B.n381 585
R147 B.n380 B.n91 585
R148 B.n379 B.n378 585
R149 B.n377 B.n92 585
R150 B.n376 B.n375 585
R151 B.n374 B.n93 585
R152 B.n373 B.n372 585
R153 B.n371 B.n94 585
R154 B.n370 B.n369 585
R155 B.n368 B.n95 585
R156 B.n195 B.n194 585
R157 B.n196 B.n153 585
R158 B.n198 B.n197 585
R159 B.n199 B.n152 585
R160 B.n201 B.n200 585
R161 B.n202 B.n151 585
R162 B.n204 B.n203 585
R163 B.n205 B.n150 585
R164 B.n207 B.n206 585
R165 B.n208 B.n149 585
R166 B.n210 B.n209 585
R167 B.n211 B.n148 585
R168 B.n213 B.n212 585
R169 B.n214 B.n147 585
R170 B.n216 B.n215 585
R171 B.n217 B.n146 585
R172 B.n219 B.n218 585
R173 B.n220 B.n145 585
R174 B.n222 B.n221 585
R175 B.n223 B.n144 585
R176 B.n225 B.n224 585
R177 B.n226 B.n143 585
R178 B.n228 B.n227 585
R179 B.n229 B.n142 585
R180 B.n231 B.n230 585
R181 B.n232 B.n141 585
R182 B.n234 B.n233 585
R183 B.n235 B.n140 585
R184 B.n237 B.n236 585
R185 B.n238 B.n139 585
R186 B.n240 B.n239 585
R187 B.n241 B.n138 585
R188 B.n243 B.n242 585
R189 B.n244 B.n137 585
R190 B.n246 B.n245 585
R191 B.n247 B.n136 585
R192 B.n249 B.n248 585
R193 B.n250 B.n135 585
R194 B.n252 B.n251 585
R195 B.n253 B.n134 585
R196 B.n255 B.n254 585
R197 B.n256 B.n133 585
R198 B.n258 B.n257 585
R199 B.n259 B.n132 585
R200 B.n261 B.n260 585
R201 B.n262 B.n131 585
R202 B.n264 B.n263 585
R203 B.n265 B.n130 585
R204 B.n267 B.n266 585
R205 B.n268 B.n129 585
R206 B.n270 B.n269 585
R207 B.n271 B.n126 585
R208 B.n274 B.n273 585
R209 B.n275 B.n125 585
R210 B.n277 B.n276 585
R211 B.n278 B.n124 585
R212 B.n280 B.n279 585
R213 B.n281 B.n123 585
R214 B.n283 B.n282 585
R215 B.n284 B.n122 585
R216 B.n289 B.n288 585
R217 B.n290 B.n121 585
R218 B.n292 B.n291 585
R219 B.n293 B.n120 585
R220 B.n295 B.n294 585
R221 B.n296 B.n119 585
R222 B.n298 B.n297 585
R223 B.n299 B.n118 585
R224 B.n301 B.n300 585
R225 B.n302 B.n117 585
R226 B.n304 B.n303 585
R227 B.n305 B.n116 585
R228 B.n307 B.n306 585
R229 B.n308 B.n115 585
R230 B.n310 B.n309 585
R231 B.n311 B.n114 585
R232 B.n313 B.n312 585
R233 B.n314 B.n113 585
R234 B.n316 B.n315 585
R235 B.n317 B.n112 585
R236 B.n319 B.n318 585
R237 B.n320 B.n111 585
R238 B.n322 B.n321 585
R239 B.n323 B.n110 585
R240 B.n325 B.n324 585
R241 B.n326 B.n109 585
R242 B.n328 B.n327 585
R243 B.n329 B.n108 585
R244 B.n331 B.n330 585
R245 B.n332 B.n107 585
R246 B.n334 B.n333 585
R247 B.n335 B.n106 585
R248 B.n337 B.n336 585
R249 B.n338 B.n105 585
R250 B.n340 B.n339 585
R251 B.n341 B.n104 585
R252 B.n343 B.n342 585
R253 B.n344 B.n103 585
R254 B.n346 B.n345 585
R255 B.n347 B.n102 585
R256 B.n349 B.n348 585
R257 B.n350 B.n101 585
R258 B.n352 B.n351 585
R259 B.n353 B.n100 585
R260 B.n355 B.n354 585
R261 B.n356 B.n99 585
R262 B.n358 B.n357 585
R263 B.n359 B.n98 585
R264 B.n361 B.n360 585
R265 B.n362 B.n97 585
R266 B.n364 B.n363 585
R267 B.n365 B.n96 585
R268 B.n367 B.n366 585
R269 B.n193 B.n154 585
R270 B.n192 B.n191 585
R271 B.n190 B.n155 585
R272 B.n189 B.n188 585
R273 B.n187 B.n156 585
R274 B.n186 B.n185 585
R275 B.n184 B.n157 585
R276 B.n183 B.n182 585
R277 B.n181 B.n158 585
R278 B.n180 B.n179 585
R279 B.n178 B.n159 585
R280 B.n177 B.n176 585
R281 B.n175 B.n160 585
R282 B.n174 B.n173 585
R283 B.n172 B.n161 585
R284 B.n171 B.n170 585
R285 B.n169 B.n162 585
R286 B.n168 B.n167 585
R287 B.n166 B.n163 585
R288 B.n165 B.n164 585
R289 B.n2 B.n0 585
R290 B.n633 B.n1 585
R291 B.n632 B.n631 585
R292 B.n630 B.n3 585
R293 B.n629 B.n628 585
R294 B.n627 B.n4 585
R295 B.n626 B.n625 585
R296 B.n624 B.n5 585
R297 B.n623 B.n622 585
R298 B.n621 B.n6 585
R299 B.n620 B.n619 585
R300 B.n618 B.n7 585
R301 B.n617 B.n616 585
R302 B.n615 B.n8 585
R303 B.n614 B.n613 585
R304 B.n612 B.n9 585
R305 B.n611 B.n610 585
R306 B.n609 B.n10 585
R307 B.n608 B.n607 585
R308 B.n606 B.n11 585
R309 B.n605 B.n604 585
R310 B.n603 B.n12 585
R311 B.n635 B.n634 585
R312 B.n195 B.n154 487.695
R313 B.n603 B.n602 487.695
R314 B.n368 B.n367 487.695
R315 B.n433 B.n74 487.695
R316 B.n285 B.t8 479.435
R317 B.n47 B.t4 479.435
R318 B.n127 B.t2 479.435
R319 B.n40 B.t10 479.435
R320 B.n286 B.t7 436.962
R321 B.n48 B.t5 436.962
R322 B.n128 B.t1 436.962
R323 B.n41 B.t11 436.962
R324 B.n285 B.t6 406.236
R325 B.n127 B.t0 406.236
R326 B.n40 B.t9 406.236
R327 B.n47 B.t3 406.236
R328 B.n191 B.n154 163.367
R329 B.n191 B.n190 163.367
R330 B.n190 B.n189 163.367
R331 B.n189 B.n156 163.367
R332 B.n185 B.n156 163.367
R333 B.n185 B.n184 163.367
R334 B.n184 B.n183 163.367
R335 B.n183 B.n158 163.367
R336 B.n179 B.n158 163.367
R337 B.n179 B.n178 163.367
R338 B.n178 B.n177 163.367
R339 B.n177 B.n160 163.367
R340 B.n173 B.n160 163.367
R341 B.n173 B.n172 163.367
R342 B.n172 B.n171 163.367
R343 B.n171 B.n162 163.367
R344 B.n167 B.n162 163.367
R345 B.n167 B.n166 163.367
R346 B.n166 B.n165 163.367
R347 B.n165 B.n2 163.367
R348 B.n634 B.n2 163.367
R349 B.n634 B.n633 163.367
R350 B.n633 B.n632 163.367
R351 B.n632 B.n3 163.367
R352 B.n628 B.n3 163.367
R353 B.n628 B.n627 163.367
R354 B.n627 B.n626 163.367
R355 B.n626 B.n5 163.367
R356 B.n622 B.n5 163.367
R357 B.n622 B.n621 163.367
R358 B.n621 B.n620 163.367
R359 B.n620 B.n7 163.367
R360 B.n616 B.n7 163.367
R361 B.n616 B.n615 163.367
R362 B.n615 B.n614 163.367
R363 B.n614 B.n9 163.367
R364 B.n610 B.n9 163.367
R365 B.n610 B.n609 163.367
R366 B.n609 B.n608 163.367
R367 B.n608 B.n11 163.367
R368 B.n604 B.n11 163.367
R369 B.n604 B.n603 163.367
R370 B.n196 B.n195 163.367
R371 B.n197 B.n196 163.367
R372 B.n197 B.n152 163.367
R373 B.n201 B.n152 163.367
R374 B.n202 B.n201 163.367
R375 B.n203 B.n202 163.367
R376 B.n203 B.n150 163.367
R377 B.n207 B.n150 163.367
R378 B.n208 B.n207 163.367
R379 B.n209 B.n208 163.367
R380 B.n209 B.n148 163.367
R381 B.n213 B.n148 163.367
R382 B.n214 B.n213 163.367
R383 B.n215 B.n214 163.367
R384 B.n215 B.n146 163.367
R385 B.n219 B.n146 163.367
R386 B.n220 B.n219 163.367
R387 B.n221 B.n220 163.367
R388 B.n221 B.n144 163.367
R389 B.n225 B.n144 163.367
R390 B.n226 B.n225 163.367
R391 B.n227 B.n226 163.367
R392 B.n227 B.n142 163.367
R393 B.n231 B.n142 163.367
R394 B.n232 B.n231 163.367
R395 B.n233 B.n232 163.367
R396 B.n233 B.n140 163.367
R397 B.n237 B.n140 163.367
R398 B.n238 B.n237 163.367
R399 B.n239 B.n238 163.367
R400 B.n239 B.n138 163.367
R401 B.n243 B.n138 163.367
R402 B.n244 B.n243 163.367
R403 B.n245 B.n244 163.367
R404 B.n245 B.n136 163.367
R405 B.n249 B.n136 163.367
R406 B.n250 B.n249 163.367
R407 B.n251 B.n250 163.367
R408 B.n251 B.n134 163.367
R409 B.n255 B.n134 163.367
R410 B.n256 B.n255 163.367
R411 B.n257 B.n256 163.367
R412 B.n257 B.n132 163.367
R413 B.n261 B.n132 163.367
R414 B.n262 B.n261 163.367
R415 B.n263 B.n262 163.367
R416 B.n263 B.n130 163.367
R417 B.n267 B.n130 163.367
R418 B.n268 B.n267 163.367
R419 B.n269 B.n268 163.367
R420 B.n269 B.n126 163.367
R421 B.n274 B.n126 163.367
R422 B.n275 B.n274 163.367
R423 B.n276 B.n275 163.367
R424 B.n276 B.n124 163.367
R425 B.n280 B.n124 163.367
R426 B.n281 B.n280 163.367
R427 B.n282 B.n281 163.367
R428 B.n282 B.n122 163.367
R429 B.n289 B.n122 163.367
R430 B.n290 B.n289 163.367
R431 B.n291 B.n290 163.367
R432 B.n291 B.n120 163.367
R433 B.n295 B.n120 163.367
R434 B.n296 B.n295 163.367
R435 B.n297 B.n296 163.367
R436 B.n297 B.n118 163.367
R437 B.n301 B.n118 163.367
R438 B.n302 B.n301 163.367
R439 B.n303 B.n302 163.367
R440 B.n303 B.n116 163.367
R441 B.n307 B.n116 163.367
R442 B.n308 B.n307 163.367
R443 B.n309 B.n308 163.367
R444 B.n309 B.n114 163.367
R445 B.n313 B.n114 163.367
R446 B.n314 B.n313 163.367
R447 B.n315 B.n314 163.367
R448 B.n315 B.n112 163.367
R449 B.n319 B.n112 163.367
R450 B.n320 B.n319 163.367
R451 B.n321 B.n320 163.367
R452 B.n321 B.n110 163.367
R453 B.n325 B.n110 163.367
R454 B.n326 B.n325 163.367
R455 B.n327 B.n326 163.367
R456 B.n327 B.n108 163.367
R457 B.n331 B.n108 163.367
R458 B.n332 B.n331 163.367
R459 B.n333 B.n332 163.367
R460 B.n333 B.n106 163.367
R461 B.n337 B.n106 163.367
R462 B.n338 B.n337 163.367
R463 B.n339 B.n338 163.367
R464 B.n339 B.n104 163.367
R465 B.n343 B.n104 163.367
R466 B.n344 B.n343 163.367
R467 B.n345 B.n344 163.367
R468 B.n345 B.n102 163.367
R469 B.n349 B.n102 163.367
R470 B.n350 B.n349 163.367
R471 B.n351 B.n350 163.367
R472 B.n351 B.n100 163.367
R473 B.n355 B.n100 163.367
R474 B.n356 B.n355 163.367
R475 B.n357 B.n356 163.367
R476 B.n357 B.n98 163.367
R477 B.n361 B.n98 163.367
R478 B.n362 B.n361 163.367
R479 B.n363 B.n362 163.367
R480 B.n363 B.n96 163.367
R481 B.n367 B.n96 163.367
R482 B.n369 B.n368 163.367
R483 B.n369 B.n94 163.367
R484 B.n373 B.n94 163.367
R485 B.n374 B.n373 163.367
R486 B.n375 B.n374 163.367
R487 B.n375 B.n92 163.367
R488 B.n379 B.n92 163.367
R489 B.n380 B.n379 163.367
R490 B.n381 B.n380 163.367
R491 B.n381 B.n90 163.367
R492 B.n385 B.n90 163.367
R493 B.n386 B.n385 163.367
R494 B.n387 B.n386 163.367
R495 B.n387 B.n88 163.367
R496 B.n391 B.n88 163.367
R497 B.n392 B.n391 163.367
R498 B.n393 B.n392 163.367
R499 B.n393 B.n86 163.367
R500 B.n397 B.n86 163.367
R501 B.n398 B.n397 163.367
R502 B.n399 B.n398 163.367
R503 B.n399 B.n84 163.367
R504 B.n403 B.n84 163.367
R505 B.n404 B.n403 163.367
R506 B.n405 B.n404 163.367
R507 B.n405 B.n82 163.367
R508 B.n409 B.n82 163.367
R509 B.n410 B.n409 163.367
R510 B.n411 B.n410 163.367
R511 B.n411 B.n80 163.367
R512 B.n415 B.n80 163.367
R513 B.n416 B.n415 163.367
R514 B.n417 B.n416 163.367
R515 B.n417 B.n78 163.367
R516 B.n421 B.n78 163.367
R517 B.n422 B.n421 163.367
R518 B.n423 B.n422 163.367
R519 B.n423 B.n76 163.367
R520 B.n427 B.n76 163.367
R521 B.n428 B.n427 163.367
R522 B.n429 B.n428 163.367
R523 B.n429 B.n74 163.367
R524 B.n602 B.n13 163.367
R525 B.n598 B.n13 163.367
R526 B.n598 B.n597 163.367
R527 B.n597 B.n596 163.367
R528 B.n596 B.n15 163.367
R529 B.n592 B.n15 163.367
R530 B.n592 B.n591 163.367
R531 B.n591 B.n590 163.367
R532 B.n590 B.n17 163.367
R533 B.n586 B.n17 163.367
R534 B.n586 B.n585 163.367
R535 B.n585 B.n584 163.367
R536 B.n584 B.n19 163.367
R537 B.n580 B.n19 163.367
R538 B.n580 B.n579 163.367
R539 B.n579 B.n578 163.367
R540 B.n578 B.n21 163.367
R541 B.n574 B.n21 163.367
R542 B.n574 B.n573 163.367
R543 B.n573 B.n572 163.367
R544 B.n572 B.n23 163.367
R545 B.n568 B.n23 163.367
R546 B.n568 B.n567 163.367
R547 B.n567 B.n566 163.367
R548 B.n566 B.n25 163.367
R549 B.n562 B.n25 163.367
R550 B.n562 B.n561 163.367
R551 B.n561 B.n560 163.367
R552 B.n560 B.n27 163.367
R553 B.n556 B.n27 163.367
R554 B.n556 B.n555 163.367
R555 B.n555 B.n554 163.367
R556 B.n554 B.n29 163.367
R557 B.n550 B.n29 163.367
R558 B.n550 B.n549 163.367
R559 B.n549 B.n548 163.367
R560 B.n548 B.n31 163.367
R561 B.n544 B.n31 163.367
R562 B.n544 B.n543 163.367
R563 B.n543 B.n542 163.367
R564 B.n542 B.n33 163.367
R565 B.n538 B.n33 163.367
R566 B.n538 B.n537 163.367
R567 B.n537 B.n536 163.367
R568 B.n536 B.n35 163.367
R569 B.n532 B.n35 163.367
R570 B.n532 B.n531 163.367
R571 B.n531 B.n530 163.367
R572 B.n530 B.n37 163.367
R573 B.n526 B.n37 163.367
R574 B.n526 B.n525 163.367
R575 B.n525 B.n524 163.367
R576 B.n524 B.n39 163.367
R577 B.n520 B.n39 163.367
R578 B.n520 B.n519 163.367
R579 B.n519 B.n518 163.367
R580 B.n518 B.n44 163.367
R581 B.n514 B.n44 163.367
R582 B.n514 B.n513 163.367
R583 B.n513 B.n512 163.367
R584 B.n512 B.n46 163.367
R585 B.n507 B.n46 163.367
R586 B.n507 B.n506 163.367
R587 B.n506 B.n505 163.367
R588 B.n505 B.n50 163.367
R589 B.n501 B.n50 163.367
R590 B.n501 B.n500 163.367
R591 B.n500 B.n499 163.367
R592 B.n499 B.n52 163.367
R593 B.n495 B.n52 163.367
R594 B.n495 B.n494 163.367
R595 B.n494 B.n493 163.367
R596 B.n493 B.n54 163.367
R597 B.n489 B.n54 163.367
R598 B.n489 B.n488 163.367
R599 B.n488 B.n487 163.367
R600 B.n487 B.n56 163.367
R601 B.n483 B.n56 163.367
R602 B.n483 B.n482 163.367
R603 B.n482 B.n481 163.367
R604 B.n481 B.n58 163.367
R605 B.n477 B.n58 163.367
R606 B.n477 B.n476 163.367
R607 B.n476 B.n475 163.367
R608 B.n475 B.n60 163.367
R609 B.n471 B.n60 163.367
R610 B.n471 B.n470 163.367
R611 B.n470 B.n469 163.367
R612 B.n469 B.n62 163.367
R613 B.n465 B.n62 163.367
R614 B.n465 B.n464 163.367
R615 B.n464 B.n463 163.367
R616 B.n463 B.n64 163.367
R617 B.n459 B.n64 163.367
R618 B.n459 B.n458 163.367
R619 B.n458 B.n457 163.367
R620 B.n457 B.n66 163.367
R621 B.n453 B.n66 163.367
R622 B.n453 B.n452 163.367
R623 B.n452 B.n451 163.367
R624 B.n451 B.n68 163.367
R625 B.n447 B.n68 163.367
R626 B.n447 B.n446 163.367
R627 B.n446 B.n445 163.367
R628 B.n445 B.n70 163.367
R629 B.n441 B.n70 163.367
R630 B.n441 B.n440 163.367
R631 B.n440 B.n439 163.367
R632 B.n439 B.n72 163.367
R633 B.n435 B.n72 163.367
R634 B.n435 B.n434 163.367
R635 B.n434 B.n433 163.367
R636 B.n287 B.n286 59.5399
R637 B.n272 B.n128 59.5399
R638 B.n42 B.n41 59.5399
R639 B.n510 B.n48 59.5399
R640 B.n286 B.n285 42.4732
R641 B.n128 B.n127 42.4732
R642 B.n41 B.n40 42.4732
R643 B.n48 B.n47 42.4732
R644 B.n601 B.n12 31.6883
R645 B.n432 B.n431 31.6883
R646 B.n366 B.n95 31.6883
R647 B.n194 B.n193 31.6883
R648 B B.n635 18.0485
R649 B.n601 B.n600 10.6151
R650 B.n600 B.n599 10.6151
R651 B.n599 B.n14 10.6151
R652 B.n595 B.n14 10.6151
R653 B.n595 B.n594 10.6151
R654 B.n594 B.n593 10.6151
R655 B.n593 B.n16 10.6151
R656 B.n589 B.n16 10.6151
R657 B.n589 B.n588 10.6151
R658 B.n588 B.n587 10.6151
R659 B.n587 B.n18 10.6151
R660 B.n583 B.n18 10.6151
R661 B.n583 B.n582 10.6151
R662 B.n582 B.n581 10.6151
R663 B.n581 B.n20 10.6151
R664 B.n577 B.n20 10.6151
R665 B.n577 B.n576 10.6151
R666 B.n576 B.n575 10.6151
R667 B.n575 B.n22 10.6151
R668 B.n571 B.n22 10.6151
R669 B.n571 B.n570 10.6151
R670 B.n570 B.n569 10.6151
R671 B.n569 B.n24 10.6151
R672 B.n565 B.n24 10.6151
R673 B.n565 B.n564 10.6151
R674 B.n564 B.n563 10.6151
R675 B.n563 B.n26 10.6151
R676 B.n559 B.n26 10.6151
R677 B.n559 B.n558 10.6151
R678 B.n558 B.n557 10.6151
R679 B.n557 B.n28 10.6151
R680 B.n553 B.n28 10.6151
R681 B.n553 B.n552 10.6151
R682 B.n552 B.n551 10.6151
R683 B.n551 B.n30 10.6151
R684 B.n547 B.n30 10.6151
R685 B.n547 B.n546 10.6151
R686 B.n546 B.n545 10.6151
R687 B.n545 B.n32 10.6151
R688 B.n541 B.n32 10.6151
R689 B.n541 B.n540 10.6151
R690 B.n540 B.n539 10.6151
R691 B.n539 B.n34 10.6151
R692 B.n535 B.n34 10.6151
R693 B.n535 B.n534 10.6151
R694 B.n534 B.n533 10.6151
R695 B.n533 B.n36 10.6151
R696 B.n529 B.n36 10.6151
R697 B.n529 B.n528 10.6151
R698 B.n528 B.n527 10.6151
R699 B.n527 B.n38 10.6151
R700 B.n523 B.n522 10.6151
R701 B.n522 B.n521 10.6151
R702 B.n521 B.n43 10.6151
R703 B.n517 B.n43 10.6151
R704 B.n517 B.n516 10.6151
R705 B.n516 B.n515 10.6151
R706 B.n515 B.n45 10.6151
R707 B.n511 B.n45 10.6151
R708 B.n509 B.n508 10.6151
R709 B.n508 B.n49 10.6151
R710 B.n504 B.n49 10.6151
R711 B.n504 B.n503 10.6151
R712 B.n503 B.n502 10.6151
R713 B.n502 B.n51 10.6151
R714 B.n498 B.n51 10.6151
R715 B.n498 B.n497 10.6151
R716 B.n497 B.n496 10.6151
R717 B.n496 B.n53 10.6151
R718 B.n492 B.n53 10.6151
R719 B.n492 B.n491 10.6151
R720 B.n491 B.n490 10.6151
R721 B.n490 B.n55 10.6151
R722 B.n486 B.n55 10.6151
R723 B.n486 B.n485 10.6151
R724 B.n485 B.n484 10.6151
R725 B.n484 B.n57 10.6151
R726 B.n480 B.n57 10.6151
R727 B.n480 B.n479 10.6151
R728 B.n479 B.n478 10.6151
R729 B.n478 B.n59 10.6151
R730 B.n474 B.n59 10.6151
R731 B.n474 B.n473 10.6151
R732 B.n473 B.n472 10.6151
R733 B.n472 B.n61 10.6151
R734 B.n468 B.n61 10.6151
R735 B.n468 B.n467 10.6151
R736 B.n467 B.n466 10.6151
R737 B.n466 B.n63 10.6151
R738 B.n462 B.n63 10.6151
R739 B.n462 B.n461 10.6151
R740 B.n461 B.n460 10.6151
R741 B.n460 B.n65 10.6151
R742 B.n456 B.n65 10.6151
R743 B.n456 B.n455 10.6151
R744 B.n455 B.n454 10.6151
R745 B.n454 B.n67 10.6151
R746 B.n450 B.n67 10.6151
R747 B.n450 B.n449 10.6151
R748 B.n449 B.n448 10.6151
R749 B.n448 B.n69 10.6151
R750 B.n444 B.n69 10.6151
R751 B.n444 B.n443 10.6151
R752 B.n443 B.n442 10.6151
R753 B.n442 B.n71 10.6151
R754 B.n438 B.n71 10.6151
R755 B.n438 B.n437 10.6151
R756 B.n437 B.n436 10.6151
R757 B.n436 B.n73 10.6151
R758 B.n432 B.n73 10.6151
R759 B.n370 B.n95 10.6151
R760 B.n371 B.n370 10.6151
R761 B.n372 B.n371 10.6151
R762 B.n372 B.n93 10.6151
R763 B.n376 B.n93 10.6151
R764 B.n377 B.n376 10.6151
R765 B.n378 B.n377 10.6151
R766 B.n378 B.n91 10.6151
R767 B.n382 B.n91 10.6151
R768 B.n383 B.n382 10.6151
R769 B.n384 B.n383 10.6151
R770 B.n384 B.n89 10.6151
R771 B.n388 B.n89 10.6151
R772 B.n389 B.n388 10.6151
R773 B.n390 B.n389 10.6151
R774 B.n390 B.n87 10.6151
R775 B.n394 B.n87 10.6151
R776 B.n395 B.n394 10.6151
R777 B.n396 B.n395 10.6151
R778 B.n396 B.n85 10.6151
R779 B.n400 B.n85 10.6151
R780 B.n401 B.n400 10.6151
R781 B.n402 B.n401 10.6151
R782 B.n402 B.n83 10.6151
R783 B.n406 B.n83 10.6151
R784 B.n407 B.n406 10.6151
R785 B.n408 B.n407 10.6151
R786 B.n408 B.n81 10.6151
R787 B.n412 B.n81 10.6151
R788 B.n413 B.n412 10.6151
R789 B.n414 B.n413 10.6151
R790 B.n414 B.n79 10.6151
R791 B.n418 B.n79 10.6151
R792 B.n419 B.n418 10.6151
R793 B.n420 B.n419 10.6151
R794 B.n420 B.n77 10.6151
R795 B.n424 B.n77 10.6151
R796 B.n425 B.n424 10.6151
R797 B.n426 B.n425 10.6151
R798 B.n426 B.n75 10.6151
R799 B.n430 B.n75 10.6151
R800 B.n431 B.n430 10.6151
R801 B.n194 B.n153 10.6151
R802 B.n198 B.n153 10.6151
R803 B.n199 B.n198 10.6151
R804 B.n200 B.n199 10.6151
R805 B.n200 B.n151 10.6151
R806 B.n204 B.n151 10.6151
R807 B.n205 B.n204 10.6151
R808 B.n206 B.n205 10.6151
R809 B.n206 B.n149 10.6151
R810 B.n210 B.n149 10.6151
R811 B.n211 B.n210 10.6151
R812 B.n212 B.n211 10.6151
R813 B.n212 B.n147 10.6151
R814 B.n216 B.n147 10.6151
R815 B.n217 B.n216 10.6151
R816 B.n218 B.n217 10.6151
R817 B.n218 B.n145 10.6151
R818 B.n222 B.n145 10.6151
R819 B.n223 B.n222 10.6151
R820 B.n224 B.n223 10.6151
R821 B.n224 B.n143 10.6151
R822 B.n228 B.n143 10.6151
R823 B.n229 B.n228 10.6151
R824 B.n230 B.n229 10.6151
R825 B.n230 B.n141 10.6151
R826 B.n234 B.n141 10.6151
R827 B.n235 B.n234 10.6151
R828 B.n236 B.n235 10.6151
R829 B.n236 B.n139 10.6151
R830 B.n240 B.n139 10.6151
R831 B.n241 B.n240 10.6151
R832 B.n242 B.n241 10.6151
R833 B.n242 B.n137 10.6151
R834 B.n246 B.n137 10.6151
R835 B.n247 B.n246 10.6151
R836 B.n248 B.n247 10.6151
R837 B.n248 B.n135 10.6151
R838 B.n252 B.n135 10.6151
R839 B.n253 B.n252 10.6151
R840 B.n254 B.n253 10.6151
R841 B.n254 B.n133 10.6151
R842 B.n258 B.n133 10.6151
R843 B.n259 B.n258 10.6151
R844 B.n260 B.n259 10.6151
R845 B.n260 B.n131 10.6151
R846 B.n264 B.n131 10.6151
R847 B.n265 B.n264 10.6151
R848 B.n266 B.n265 10.6151
R849 B.n266 B.n129 10.6151
R850 B.n270 B.n129 10.6151
R851 B.n271 B.n270 10.6151
R852 B.n273 B.n125 10.6151
R853 B.n277 B.n125 10.6151
R854 B.n278 B.n277 10.6151
R855 B.n279 B.n278 10.6151
R856 B.n279 B.n123 10.6151
R857 B.n283 B.n123 10.6151
R858 B.n284 B.n283 10.6151
R859 B.n288 B.n284 10.6151
R860 B.n292 B.n121 10.6151
R861 B.n293 B.n292 10.6151
R862 B.n294 B.n293 10.6151
R863 B.n294 B.n119 10.6151
R864 B.n298 B.n119 10.6151
R865 B.n299 B.n298 10.6151
R866 B.n300 B.n299 10.6151
R867 B.n300 B.n117 10.6151
R868 B.n304 B.n117 10.6151
R869 B.n305 B.n304 10.6151
R870 B.n306 B.n305 10.6151
R871 B.n306 B.n115 10.6151
R872 B.n310 B.n115 10.6151
R873 B.n311 B.n310 10.6151
R874 B.n312 B.n311 10.6151
R875 B.n312 B.n113 10.6151
R876 B.n316 B.n113 10.6151
R877 B.n317 B.n316 10.6151
R878 B.n318 B.n317 10.6151
R879 B.n318 B.n111 10.6151
R880 B.n322 B.n111 10.6151
R881 B.n323 B.n322 10.6151
R882 B.n324 B.n323 10.6151
R883 B.n324 B.n109 10.6151
R884 B.n328 B.n109 10.6151
R885 B.n329 B.n328 10.6151
R886 B.n330 B.n329 10.6151
R887 B.n330 B.n107 10.6151
R888 B.n334 B.n107 10.6151
R889 B.n335 B.n334 10.6151
R890 B.n336 B.n335 10.6151
R891 B.n336 B.n105 10.6151
R892 B.n340 B.n105 10.6151
R893 B.n341 B.n340 10.6151
R894 B.n342 B.n341 10.6151
R895 B.n342 B.n103 10.6151
R896 B.n346 B.n103 10.6151
R897 B.n347 B.n346 10.6151
R898 B.n348 B.n347 10.6151
R899 B.n348 B.n101 10.6151
R900 B.n352 B.n101 10.6151
R901 B.n353 B.n352 10.6151
R902 B.n354 B.n353 10.6151
R903 B.n354 B.n99 10.6151
R904 B.n358 B.n99 10.6151
R905 B.n359 B.n358 10.6151
R906 B.n360 B.n359 10.6151
R907 B.n360 B.n97 10.6151
R908 B.n364 B.n97 10.6151
R909 B.n365 B.n364 10.6151
R910 B.n366 B.n365 10.6151
R911 B.n193 B.n192 10.6151
R912 B.n192 B.n155 10.6151
R913 B.n188 B.n155 10.6151
R914 B.n188 B.n187 10.6151
R915 B.n187 B.n186 10.6151
R916 B.n186 B.n157 10.6151
R917 B.n182 B.n157 10.6151
R918 B.n182 B.n181 10.6151
R919 B.n181 B.n180 10.6151
R920 B.n180 B.n159 10.6151
R921 B.n176 B.n159 10.6151
R922 B.n176 B.n175 10.6151
R923 B.n175 B.n174 10.6151
R924 B.n174 B.n161 10.6151
R925 B.n170 B.n161 10.6151
R926 B.n170 B.n169 10.6151
R927 B.n169 B.n168 10.6151
R928 B.n168 B.n163 10.6151
R929 B.n164 B.n163 10.6151
R930 B.n164 B.n0 10.6151
R931 B.n631 B.n1 10.6151
R932 B.n631 B.n630 10.6151
R933 B.n630 B.n629 10.6151
R934 B.n629 B.n4 10.6151
R935 B.n625 B.n4 10.6151
R936 B.n625 B.n624 10.6151
R937 B.n624 B.n623 10.6151
R938 B.n623 B.n6 10.6151
R939 B.n619 B.n6 10.6151
R940 B.n619 B.n618 10.6151
R941 B.n618 B.n617 10.6151
R942 B.n617 B.n8 10.6151
R943 B.n613 B.n8 10.6151
R944 B.n613 B.n612 10.6151
R945 B.n612 B.n611 10.6151
R946 B.n611 B.n10 10.6151
R947 B.n607 B.n10 10.6151
R948 B.n607 B.n606 10.6151
R949 B.n606 B.n605 10.6151
R950 B.n605 B.n12 10.6151
R951 B.n523 B.n42 6.5566
R952 B.n511 B.n510 6.5566
R953 B.n273 B.n272 6.5566
R954 B.n288 B.n287 6.5566
R955 B.n42 B.n38 4.05904
R956 B.n510 B.n509 4.05904
R957 B.n272 B.n271 4.05904
R958 B.n287 B.n121 4.05904
R959 B.n635 B.n0 2.81026
R960 B.n635 B.n1 2.81026
R961 VP.n0 VP.t0 303.805
R962 VP.n0 VP.t1 258.529
R963 VP VP.n0 0.241678
R964 VTAIL.n338 VTAIL.n258 756.745
R965 VTAIL.n80 VTAIL.n0 756.745
R966 VTAIL.n252 VTAIL.n172 756.745
R967 VTAIL.n166 VTAIL.n86 756.745
R968 VTAIL.n287 VTAIL.n286 585
R969 VTAIL.n289 VTAIL.n288 585
R970 VTAIL.n282 VTAIL.n281 585
R971 VTAIL.n295 VTAIL.n294 585
R972 VTAIL.n297 VTAIL.n296 585
R973 VTAIL.n278 VTAIL.n277 585
R974 VTAIL.n303 VTAIL.n302 585
R975 VTAIL.n305 VTAIL.n304 585
R976 VTAIL.n274 VTAIL.n273 585
R977 VTAIL.n311 VTAIL.n310 585
R978 VTAIL.n313 VTAIL.n312 585
R979 VTAIL.n270 VTAIL.n269 585
R980 VTAIL.n319 VTAIL.n318 585
R981 VTAIL.n321 VTAIL.n320 585
R982 VTAIL.n266 VTAIL.n265 585
R983 VTAIL.n328 VTAIL.n327 585
R984 VTAIL.n329 VTAIL.n264 585
R985 VTAIL.n331 VTAIL.n330 585
R986 VTAIL.n262 VTAIL.n261 585
R987 VTAIL.n337 VTAIL.n336 585
R988 VTAIL.n339 VTAIL.n338 585
R989 VTAIL.n29 VTAIL.n28 585
R990 VTAIL.n31 VTAIL.n30 585
R991 VTAIL.n24 VTAIL.n23 585
R992 VTAIL.n37 VTAIL.n36 585
R993 VTAIL.n39 VTAIL.n38 585
R994 VTAIL.n20 VTAIL.n19 585
R995 VTAIL.n45 VTAIL.n44 585
R996 VTAIL.n47 VTAIL.n46 585
R997 VTAIL.n16 VTAIL.n15 585
R998 VTAIL.n53 VTAIL.n52 585
R999 VTAIL.n55 VTAIL.n54 585
R1000 VTAIL.n12 VTAIL.n11 585
R1001 VTAIL.n61 VTAIL.n60 585
R1002 VTAIL.n63 VTAIL.n62 585
R1003 VTAIL.n8 VTAIL.n7 585
R1004 VTAIL.n70 VTAIL.n69 585
R1005 VTAIL.n71 VTAIL.n6 585
R1006 VTAIL.n73 VTAIL.n72 585
R1007 VTAIL.n4 VTAIL.n3 585
R1008 VTAIL.n79 VTAIL.n78 585
R1009 VTAIL.n81 VTAIL.n80 585
R1010 VTAIL.n253 VTAIL.n252 585
R1011 VTAIL.n251 VTAIL.n250 585
R1012 VTAIL.n176 VTAIL.n175 585
R1013 VTAIL.n180 VTAIL.n178 585
R1014 VTAIL.n245 VTAIL.n244 585
R1015 VTAIL.n243 VTAIL.n242 585
R1016 VTAIL.n182 VTAIL.n181 585
R1017 VTAIL.n237 VTAIL.n236 585
R1018 VTAIL.n235 VTAIL.n234 585
R1019 VTAIL.n186 VTAIL.n185 585
R1020 VTAIL.n229 VTAIL.n228 585
R1021 VTAIL.n227 VTAIL.n226 585
R1022 VTAIL.n190 VTAIL.n189 585
R1023 VTAIL.n221 VTAIL.n220 585
R1024 VTAIL.n219 VTAIL.n218 585
R1025 VTAIL.n194 VTAIL.n193 585
R1026 VTAIL.n213 VTAIL.n212 585
R1027 VTAIL.n211 VTAIL.n210 585
R1028 VTAIL.n198 VTAIL.n197 585
R1029 VTAIL.n205 VTAIL.n204 585
R1030 VTAIL.n203 VTAIL.n202 585
R1031 VTAIL.n167 VTAIL.n166 585
R1032 VTAIL.n165 VTAIL.n164 585
R1033 VTAIL.n90 VTAIL.n89 585
R1034 VTAIL.n94 VTAIL.n92 585
R1035 VTAIL.n159 VTAIL.n158 585
R1036 VTAIL.n157 VTAIL.n156 585
R1037 VTAIL.n96 VTAIL.n95 585
R1038 VTAIL.n151 VTAIL.n150 585
R1039 VTAIL.n149 VTAIL.n148 585
R1040 VTAIL.n100 VTAIL.n99 585
R1041 VTAIL.n143 VTAIL.n142 585
R1042 VTAIL.n141 VTAIL.n140 585
R1043 VTAIL.n104 VTAIL.n103 585
R1044 VTAIL.n135 VTAIL.n134 585
R1045 VTAIL.n133 VTAIL.n132 585
R1046 VTAIL.n108 VTAIL.n107 585
R1047 VTAIL.n127 VTAIL.n126 585
R1048 VTAIL.n125 VTAIL.n124 585
R1049 VTAIL.n112 VTAIL.n111 585
R1050 VTAIL.n119 VTAIL.n118 585
R1051 VTAIL.n117 VTAIL.n116 585
R1052 VTAIL.n285 VTAIL.t0 327.466
R1053 VTAIL.n27 VTAIL.t2 327.466
R1054 VTAIL.n201 VTAIL.t3 327.466
R1055 VTAIL.n115 VTAIL.t1 327.466
R1056 VTAIL.n288 VTAIL.n287 171.744
R1057 VTAIL.n288 VTAIL.n281 171.744
R1058 VTAIL.n295 VTAIL.n281 171.744
R1059 VTAIL.n296 VTAIL.n295 171.744
R1060 VTAIL.n296 VTAIL.n277 171.744
R1061 VTAIL.n303 VTAIL.n277 171.744
R1062 VTAIL.n304 VTAIL.n303 171.744
R1063 VTAIL.n304 VTAIL.n273 171.744
R1064 VTAIL.n311 VTAIL.n273 171.744
R1065 VTAIL.n312 VTAIL.n311 171.744
R1066 VTAIL.n312 VTAIL.n269 171.744
R1067 VTAIL.n319 VTAIL.n269 171.744
R1068 VTAIL.n320 VTAIL.n319 171.744
R1069 VTAIL.n320 VTAIL.n265 171.744
R1070 VTAIL.n328 VTAIL.n265 171.744
R1071 VTAIL.n329 VTAIL.n328 171.744
R1072 VTAIL.n330 VTAIL.n329 171.744
R1073 VTAIL.n330 VTAIL.n261 171.744
R1074 VTAIL.n337 VTAIL.n261 171.744
R1075 VTAIL.n338 VTAIL.n337 171.744
R1076 VTAIL.n30 VTAIL.n29 171.744
R1077 VTAIL.n30 VTAIL.n23 171.744
R1078 VTAIL.n37 VTAIL.n23 171.744
R1079 VTAIL.n38 VTAIL.n37 171.744
R1080 VTAIL.n38 VTAIL.n19 171.744
R1081 VTAIL.n45 VTAIL.n19 171.744
R1082 VTAIL.n46 VTAIL.n45 171.744
R1083 VTAIL.n46 VTAIL.n15 171.744
R1084 VTAIL.n53 VTAIL.n15 171.744
R1085 VTAIL.n54 VTAIL.n53 171.744
R1086 VTAIL.n54 VTAIL.n11 171.744
R1087 VTAIL.n61 VTAIL.n11 171.744
R1088 VTAIL.n62 VTAIL.n61 171.744
R1089 VTAIL.n62 VTAIL.n7 171.744
R1090 VTAIL.n70 VTAIL.n7 171.744
R1091 VTAIL.n71 VTAIL.n70 171.744
R1092 VTAIL.n72 VTAIL.n71 171.744
R1093 VTAIL.n72 VTAIL.n3 171.744
R1094 VTAIL.n79 VTAIL.n3 171.744
R1095 VTAIL.n80 VTAIL.n79 171.744
R1096 VTAIL.n252 VTAIL.n251 171.744
R1097 VTAIL.n251 VTAIL.n175 171.744
R1098 VTAIL.n180 VTAIL.n175 171.744
R1099 VTAIL.n244 VTAIL.n180 171.744
R1100 VTAIL.n244 VTAIL.n243 171.744
R1101 VTAIL.n243 VTAIL.n181 171.744
R1102 VTAIL.n236 VTAIL.n181 171.744
R1103 VTAIL.n236 VTAIL.n235 171.744
R1104 VTAIL.n235 VTAIL.n185 171.744
R1105 VTAIL.n228 VTAIL.n185 171.744
R1106 VTAIL.n228 VTAIL.n227 171.744
R1107 VTAIL.n227 VTAIL.n189 171.744
R1108 VTAIL.n220 VTAIL.n189 171.744
R1109 VTAIL.n220 VTAIL.n219 171.744
R1110 VTAIL.n219 VTAIL.n193 171.744
R1111 VTAIL.n212 VTAIL.n193 171.744
R1112 VTAIL.n212 VTAIL.n211 171.744
R1113 VTAIL.n211 VTAIL.n197 171.744
R1114 VTAIL.n204 VTAIL.n197 171.744
R1115 VTAIL.n204 VTAIL.n203 171.744
R1116 VTAIL.n166 VTAIL.n165 171.744
R1117 VTAIL.n165 VTAIL.n89 171.744
R1118 VTAIL.n94 VTAIL.n89 171.744
R1119 VTAIL.n158 VTAIL.n94 171.744
R1120 VTAIL.n158 VTAIL.n157 171.744
R1121 VTAIL.n157 VTAIL.n95 171.744
R1122 VTAIL.n150 VTAIL.n95 171.744
R1123 VTAIL.n150 VTAIL.n149 171.744
R1124 VTAIL.n149 VTAIL.n99 171.744
R1125 VTAIL.n142 VTAIL.n99 171.744
R1126 VTAIL.n142 VTAIL.n141 171.744
R1127 VTAIL.n141 VTAIL.n103 171.744
R1128 VTAIL.n134 VTAIL.n103 171.744
R1129 VTAIL.n134 VTAIL.n133 171.744
R1130 VTAIL.n133 VTAIL.n107 171.744
R1131 VTAIL.n126 VTAIL.n107 171.744
R1132 VTAIL.n126 VTAIL.n125 171.744
R1133 VTAIL.n125 VTAIL.n111 171.744
R1134 VTAIL.n118 VTAIL.n111 171.744
R1135 VTAIL.n118 VTAIL.n117 171.744
R1136 VTAIL.n287 VTAIL.t0 85.8723
R1137 VTAIL.n29 VTAIL.t2 85.8723
R1138 VTAIL.n203 VTAIL.t3 85.8723
R1139 VTAIL.n117 VTAIL.t1 85.8723
R1140 VTAIL.n343 VTAIL.n342 33.155
R1141 VTAIL.n85 VTAIL.n84 33.155
R1142 VTAIL.n257 VTAIL.n256 33.155
R1143 VTAIL.n171 VTAIL.n170 33.155
R1144 VTAIL.n171 VTAIL.n85 29.4272
R1145 VTAIL.n343 VTAIL.n257 27.5393
R1146 VTAIL.n286 VTAIL.n285 16.3895
R1147 VTAIL.n28 VTAIL.n27 16.3895
R1148 VTAIL.n202 VTAIL.n201 16.3895
R1149 VTAIL.n116 VTAIL.n115 16.3895
R1150 VTAIL.n331 VTAIL.n262 13.1884
R1151 VTAIL.n73 VTAIL.n4 13.1884
R1152 VTAIL.n178 VTAIL.n176 13.1884
R1153 VTAIL.n92 VTAIL.n90 13.1884
R1154 VTAIL.n289 VTAIL.n284 12.8005
R1155 VTAIL.n332 VTAIL.n264 12.8005
R1156 VTAIL.n336 VTAIL.n335 12.8005
R1157 VTAIL.n31 VTAIL.n26 12.8005
R1158 VTAIL.n74 VTAIL.n6 12.8005
R1159 VTAIL.n78 VTAIL.n77 12.8005
R1160 VTAIL.n250 VTAIL.n249 12.8005
R1161 VTAIL.n246 VTAIL.n245 12.8005
R1162 VTAIL.n205 VTAIL.n200 12.8005
R1163 VTAIL.n164 VTAIL.n163 12.8005
R1164 VTAIL.n160 VTAIL.n159 12.8005
R1165 VTAIL.n119 VTAIL.n114 12.8005
R1166 VTAIL.n290 VTAIL.n282 12.0247
R1167 VTAIL.n327 VTAIL.n326 12.0247
R1168 VTAIL.n339 VTAIL.n260 12.0247
R1169 VTAIL.n32 VTAIL.n24 12.0247
R1170 VTAIL.n69 VTAIL.n68 12.0247
R1171 VTAIL.n81 VTAIL.n2 12.0247
R1172 VTAIL.n253 VTAIL.n174 12.0247
R1173 VTAIL.n242 VTAIL.n179 12.0247
R1174 VTAIL.n206 VTAIL.n198 12.0247
R1175 VTAIL.n167 VTAIL.n88 12.0247
R1176 VTAIL.n156 VTAIL.n93 12.0247
R1177 VTAIL.n120 VTAIL.n112 12.0247
R1178 VTAIL.n294 VTAIL.n293 11.249
R1179 VTAIL.n325 VTAIL.n266 11.249
R1180 VTAIL.n340 VTAIL.n258 11.249
R1181 VTAIL.n36 VTAIL.n35 11.249
R1182 VTAIL.n67 VTAIL.n8 11.249
R1183 VTAIL.n82 VTAIL.n0 11.249
R1184 VTAIL.n254 VTAIL.n172 11.249
R1185 VTAIL.n241 VTAIL.n182 11.249
R1186 VTAIL.n210 VTAIL.n209 11.249
R1187 VTAIL.n168 VTAIL.n86 11.249
R1188 VTAIL.n155 VTAIL.n96 11.249
R1189 VTAIL.n124 VTAIL.n123 11.249
R1190 VTAIL.n297 VTAIL.n280 10.4732
R1191 VTAIL.n322 VTAIL.n321 10.4732
R1192 VTAIL.n39 VTAIL.n22 10.4732
R1193 VTAIL.n64 VTAIL.n63 10.4732
R1194 VTAIL.n238 VTAIL.n237 10.4732
R1195 VTAIL.n213 VTAIL.n196 10.4732
R1196 VTAIL.n152 VTAIL.n151 10.4732
R1197 VTAIL.n127 VTAIL.n110 10.4732
R1198 VTAIL.n298 VTAIL.n278 9.69747
R1199 VTAIL.n318 VTAIL.n268 9.69747
R1200 VTAIL.n40 VTAIL.n20 9.69747
R1201 VTAIL.n60 VTAIL.n10 9.69747
R1202 VTAIL.n234 VTAIL.n184 9.69747
R1203 VTAIL.n214 VTAIL.n194 9.69747
R1204 VTAIL.n148 VTAIL.n98 9.69747
R1205 VTAIL.n128 VTAIL.n108 9.69747
R1206 VTAIL.n342 VTAIL.n341 9.45567
R1207 VTAIL.n84 VTAIL.n83 9.45567
R1208 VTAIL.n256 VTAIL.n255 9.45567
R1209 VTAIL.n170 VTAIL.n169 9.45567
R1210 VTAIL.n341 VTAIL.n340 9.3005
R1211 VTAIL.n260 VTAIL.n259 9.3005
R1212 VTAIL.n335 VTAIL.n334 9.3005
R1213 VTAIL.n307 VTAIL.n306 9.3005
R1214 VTAIL.n276 VTAIL.n275 9.3005
R1215 VTAIL.n301 VTAIL.n300 9.3005
R1216 VTAIL.n299 VTAIL.n298 9.3005
R1217 VTAIL.n280 VTAIL.n279 9.3005
R1218 VTAIL.n293 VTAIL.n292 9.3005
R1219 VTAIL.n291 VTAIL.n290 9.3005
R1220 VTAIL.n284 VTAIL.n283 9.3005
R1221 VTAIL.n309 VTAIL.n308 9.3005
R1222 VTAIL.n272 VTAIL.n271 9.3005
R1223 VTAIL.n315 VTAIL.n314 9.3005
R1224 VTAIL.n317 VTAIL.n316 9.3005
R1225 VTAIL.n268 VTAIL.n267 9.3005
R1226 VTAIL.n323 VTAIL.n322 9.3005
R1227 VTAIL.n325 VTAIL.n324 9.3005
R1228 VTAIL.n326 VTAIL.n263 9.3005
R1229 VTAIL.n333 VTAIL.n332 9.3005
R1230 VTAIL.n83 VTAIL.n82 9.3005
R1231 VTAIL.n2 VTAIL.n1 9.3005
R1232 VTAIL.n77 VTAIL.n76 9.3005
R1233 VTAIL.n49 VTAIL.n48 9.3005
R1234 VTAIL.n18 VTAIL.n17 9.3005
R1235 VTAIL.n43 VTAIL.n42 9.3005
R1236 VTAIL.n41 VTAIL.n40 9.3005
R1237 VTAIL.n22 VTAIL.n21 9.3005
R1238 VTAIL.n35 VTAIL.n34 9.3005
R1239 VTAIL.n33 VTAIL.n32 9.3005
R1240 VTAIL.n26 VTAIL.n25 9.3005
R1241 VTAIL.n51 VTAIL.n50 9.3005
R1242 VTAIL.n14 VTAIL.n13 9.3005
R1243 VTAIL.n57 VTAIL.n56 9.3005
R1244 VTAIL.n59 VTAIL.n58 9.3005
R1245 VTAIL.n10 VTAIL.n9 9.3005
R1246 VTAIL.n65 VTAIL.n64 9.3005
R1247 VTAIL.n67 VTAIL.n66 9.3005
R1248 VTAIL.n68 VTAIL.n5 9.3005
R1249 VTAIL.n75 VTAIL.n74 9.3005
R1250 VTAIL.n188 VTAIL.n187 9.3005
R1251 VTAIL.n231 VTAIL.n230 9.3005
R1252 VTAIL.n233 VTAIL.n232 9.3005
R1253 VTAIL.n184 VTAIL.n183 9.3005
R1254 VTAIL.n239 VTAIL.n238 9.3005
R1255 VTAIL.n241 VTAIL.n240 9.3005
R1256 VTAIL.n179 VTAIL.n177 9.3005
R1257 VTAIL.n247 VTAIL.n246 9.3005
R1258 VTAIL.n255 VTAIL.n254 9.3005
R1259 VTAIL.n174 VTAIL.n173 9.3005
R1260 VTAIL.n249 VTAIL.n248 9.3005
R1261 VTAIL.n225 VTAIL.n224 9.3005
R1262 VTAIL.n223 VTAIL.n222 9.3005
R1263 VTAIL.n192 VTAIL.n191 9.3005
R1264 VTAIL.n217 VTAIL.n216 9.3005
R1265 VTAIL.n215 VTAIL.n214 9.3005
R1266 VTAIL.n196 VTAIL.n195 9.3005
R1267 VTAIL.n209 VTAIL.n208 9.3005
R1268 VTAIL.n207 VTAIL.n206 9.3005
R1269 VTAIL.n200 VTAIL.n199 9.3005
R1270 VTAIL.n102 VTAIL.n101 9.3005
R1271 VTAIL.n145 VTAIL.n144 9.3005
R1272 VTAIL.n147 VTAIL.n146 9.3005
R1273 VTAIL.n98 VTAIL.n97 9.3005
R1274 VTAIL.n153 VTAIL.n152 9.3005
R1275 VTAIL.n155 VTAIL.n154 9.3005
R1276 VTAIL.n93 VTAIL.n91 9.3005
R1277 VTAIL.n161 VTAIL.n160 9.3005
R1278 VTAIL.n169 VTAIL.n168 9.3005
R1279 VTAIL.n88 VTAIL.n87 9.3005
R1280 VTAIL.n163 VTAIL.n162 9.3005
R1281 VTAIL.n139 VTAIL.n138 9.3005
R1282 VTAIL.n137 VTAIL.n136 9.3005
R1283 VTAIL.n106 VTAIL.n105 9.3005
R1284 VTAIL.n131 VTAIL.n130 9.3005
R1285 VTAIL.n129 VTAIL.n128 9.3005
R1286 VTAIL.n110 VTAIL.n109 9.3005
R1287 VTAIL.n123 VTAIL.n122 9.3005
R1288 VTAIL.n121 VTAIL.n120 9.3005
R1289 VTAIL.n114 VTAIL.n113 9.3005
R1290 VTAIL.n302 VTAIL.n301 8.92171
R1291 VTAIL.n317 VTAIL.n270 8.92171
R1292 VTAIL.n44 VTAIL.n43 8.92171
R1293 VTAIL.n59 VTAIL.n12 8.92171
R1294 VTAIL.n233 VTAIL.n186 8.92171
R1295 VTAIL.n218 VTAIL.n217 8.92171
R1296 VTAIL.n147 VTAIL.n100 8.92171
R1297 VTAIL.n132 VTAIL.n131 8.92171
R1298 VTAIL.n305 VTAIL.n276 8.14595
R1299 VTAIL.n314 VTAIL.n313 8.14595
R1300 VTAIL.n47 VTAIL.n18 8.14595
R1301 VTAIL.n56 VTAIL.n55 8.14595
R1302 VTAIL.n230 VTAIL.n229 8.14595
R1303 VTAIL.n221 VTAIL.n192 8.14595
R1304 VTAIL.n144 VTAIL.n143 8.14595
R1305 VTAIL.n135 VTAIL.n106 8.14595
R1306 VTAIL.n306 VTAIL.n274 7.3702
R1307 VTAIL.n310 VTAIL.n272 7.3702
R1308 VTAIL.n48 VTAIL.n16 7.3702
R1309 VTAIL.n52 VTAIL.n14 7.3702
R1310 VTAIL.n226 VTAIL.n188 7.3702
R1311 VTAIL.n222 VTAIL.n190 7.3702
R1312 VTAIL.n140 VTAIL.n102 7.3702
R1313 VTAIL.n136 VTAIL.n104 7.3702
R1314 VTAIL.n309 VTAIL.n274 6.59444
R1315 VTAIL.n310 VTAIL.n309 6.59444
R1316 VTAIL.n51 VTAIL.n16 6.59444
R1317 VTAIL.n52 VTAIL.n51 6.59444
R1318 VTAIL.n226 VTAIL.n225 6.59444
R1319 VTAIL.n225 VTAIL.n190 6.59444
R1320 VTAIL.n140 VTAIL.n139 6.59444
R1321 VTAIL.n139 VTAIL.n104 6.59444
R1322 VTAIL.n306 VTAIL.n305 5.81868
R1323 VTAIL.n313 VTAIL.n272 5.81868
R1324 VTAIL.n48 VTAIL.n47 5.81868
R1325 VTAIL.n55 VTAIL.n14 5.81868
R1326 VTAIL.n229 VTAIL.n188 5.81868
R1327 VTAIL.n222 VTAIL.n221 5.81868
R1328 VTAIL.n143 VTAIL.n102 5.81868
R1329 VTAIL.n136 VTAIL.n135 5.81868
R1330 VTAIL.n302 VTAIL.n276 5.04292
R1331 VTAIL.n314 VTAIL.n270 5.04292
R1332 VTAIL.n44 VTAIL.n18 5.04292
R1333 VTAIL.n56 VTAIL.n12 5.04292
R1334 VTAIL.n230 VTAIL.n186 5.04292
R1335 VTAIL.n218 VTAIL.n192 5.04292
R1336 VTAIL.n144 VTAIL.n100 5.04292
R1337 VTAIL.n132 VTAIL.n106 5.04292
R1338 VTAIL.n301 VTAIL.n278 4.26717
R1339 VTAIL.n318 VTAIL.n317 4.26717
R1340 VTAIL.n43 VTAIL.n20 4.26717
R1341 VTAIL.n60 VTAIL.n59 4.26717
R1342 VTAIL.n234 VTAIL.n233 4.26717
R1343 VTAIL.n217 VTAIL.n194 4.26717
R1344 VTAIL.n148 VTAIL.n147 4.26717
R1345 VTAIL.n131 VTAIL.n108 4.26717
R1346 VTAIL.n285 VTAIL.n283 3.70982
R1347 VTAIL.n27 VTAIL.n25 3.70982
R1348 VTAIL.n201 VTAIL.n199 3.70982
R1349 VTAIL.n115 VTAIL.n113 3.70982
R1350 VTAIL.n298 VTAIL.n297 3.49141
R1351 VTAIL.n321 VTAIL.n268 3.49141
R1352 VTAIL.n40 VTAIL.n39 3.49141
R1353 VTAIL.n63 VTAIL.n10 3.49141
R1354 VTAIL.n237 VTAIL.n184 3.49141
R1355 VTAIL.n214 VTAIL.n213 3.49141
R1356 VTAIL.n151 VTAIL.n98 3.49141
R1357 VTAIL.n128 VTAIL.n127 3.49141
R1358 VTAIL.n294 VTAIL.n280 2.71565
R1359 VTAIL.n322 VTAIL.n266 2.71565
R1360 VTAIL.n342 VTAIL.n258 2.71565
R1361 VTAIL.n36 VTAIL.n22 2.71565
R1362 VTAIL.n64 VTAIL.n8 2.71565
R1363 VTAIL.n84 VTAIL.n0 2.71565
R1364 VTAIL.n256 VTAIL.n172 2.71565
R1365 VTAIL.n238 VTAIL.n182 2.71565
R1366 VTAIL.n210 VTAIL.n196 2.71565
R1367 VTAIL.n170 VTAIL.n86 2.71565
R1368 VTAIL.n152 VTAIL.n96 2.71565
R1369 VTAIL.n124 VTAIL.n110 2.71565
R1370 VTAIL.n293 VTAIL.n282 1.93989
R1371 VTAIL.n327 VTAIL.n325 1.93989
R1372 VTAIL.n340 VTAIL.n339 1.93989
R1373 VTAIL.n35 VTAIL.n24 1.93989
R1374 VTAIL.n69 VTAIL.n67 1.93989
R1375 VTAIL.n82 VTAIL.n81 1.93989
R1376 VTAIL.n254 VTAIL.n253 1.93989
R1377 VTAIL.n242 VTAIL.n241 1.93989
R1378 VTAIL.n209 VTAIL.n198 1.93989
R1379 VTAIL.n168 VTAIL.n167 1.93989
R1380 VTAIL.n156 VTAIL.n155 1.93989
R1381 VTAIL.n123 VTAIL.n112 1.93989
R1382 VTAIL.n257 VTAIL.n171 1.41429
R1383 VTAIL.n290 VTAIL.n289 1.16414
R1384 VTAIL.n326 VTAIL.n264 1.16414
R1385 VTAIL.n336 VTAIL.n260 1.16414
R1386 VTAIL.n32 VTAIL.n31 1.16414
R1387 VTAIL.n68 VTAIL.n6 1.16414
R1388 VTAIL.n78 VTAIL.n2 1.16414
R1389 VTAIL.n250 VTAIL.n174 1.16414
R1390 VTAIL.n245 VTAIL.n179 1.16414
R1391 VTAIL.n206 VTAIL.n205 1.16414
R1392 VTAIL.n164 VTAIL.n88 1.16414
R1393 VTAIL.n159 VTAIL.n93 1.16414
R1394 VTAIL.n120 VTAIL.n119 1.16414
R1395 VTAIL VTAIL.n85 1.0005
R1396 VTAIL VTAIL.n343 0.414293
R1397 VTAIL.n286 VTAIL.n284 0.388379
R1398 VTAIL.n332 VTAIL.n331 0.388379
R1399 VTAIL.n335 VTAIL.n262 0.388379
R1400 VTAIL.n28 VTAIL.n26 0.388379
R1401 VTAIL.n74 VTAIL.n73 0.388379
R1402 VTAIL.n77 VTAIL.n4 0.388379
R1403 VTAIL.n249 VTAIL.n176 0.388379
R1404 VTAIL.n246 VTAIL.n178 0.388379
R1405 VTAIL.n202 VTAIL.n200 0.388379
R1406 VTAIL.n163 VTAIL.n90 0.388379
R1407 VTAIL.n160 VTAIL.n92 0.388379
R1408 VTAIL.n116 VTAIL.n114 0.388379
R1409 VTAIL.n291 VTAIL.n283 0.155672
R1410 VTAIL.n292 VTAIL.n291 0.155672
R1411 VTAIL.n292 VTAIL.n279 0.155672
R1412 VTAIL.n299 VTAIL.n279 0.155672
R1413 VTAIL.n300 VTAIL.n299 0.155672
R1414 VTAIL.n300 VTAIL.n275 0.155672
R1415 VTAIL.n307 VTAIL.n275 0.155672
R1416 VTAIL.n308 VTAIL.n307 0.155672
R1417 VTAIL.n308 VTAIL.n271 0.155672
R1418 VTAIL.n315 VTAIL.n271 0.155672
R1419 VTAIL.n316 VTAIL.n315 0.155672
R1420 VTAIL.n316 VTAIL.n267 0.155672
R1421 VTAIL.n323 VTAIL.n267 0.155672
R1422 VTAIL.n324 VTAIL.n323 0.155672
R1423 VTAIL.n324 VTAIL.n263 0.155672
R1424 VTAIL.n333 VTAIL.n263 0.155672
R1425 VTAIL.n334 VTAIL.n333 0.155672
R1426 VTAIL.n334 VTAIL.n259 0.155672
R1427 VTAIL.n341 VTAIL.n259 0.155672
R1428 VTAIL.n33 VTAIL.n25 0.155672
R1429 VTAIL.n34 VTAIL.n33 0.155672
R1430 VTAIL.n34 VTAIL.n21 0.155672
R1431 VTAIL.n41 VTAIL.n21 0.155672
R1432 VTAIL.n42 VTAIL.n41 0.155672
R1433 VTAIL.n42 VTAIL.n17 0.155672
R1434 VTAIL.n49 VTAIL.n17 0.155672
R1435 VTAIL.n50 VTAIL.n49 0.155672
R1436 VTAIL.n50 VTAIL.n13 0.155672
R1437 VTAIL.n57 VTAIL.n13 0.155672
R1438 VTAIL.n58 VTAIL.n57 0.155672
R1439 VTAIL.n58 VTAIL.n9 0.155672
R1440 VTAIL.n65 VTAIL.n9 0.155672
R1441 VTAIL.n66 VTAIL.n65 0.155672
R1442 VTAIL.n66 VTAIL.n5 0.155672
R1443 VTAIL.n75 VTAIL.n5 0.155672
R1444 VTAIL.n76 VTAIL.n75 0.155672
R1445 VTAIL.n76 VTAIL.n1 0.155672
R1446 VTAIL.n83 VTAIL.n1 0.155672
R1447 VTAIL.n255 VTAIL.n173 0.155672
R1448 VTAIL.n248 VTAIL.n173 0.155672
R1449 VTAIL.n248 VTAIL.n247 0.155672
R1450 VTAIL.n247 VTAIL.n177 0.155672
R1451 VTAIL.n240 VTAIL.n177 0.155672
R1452 VTAIL.n240 VTAIL.n239 0.155672
R1453 VTAIL.n239 VTAIL.n183 0.155672
R1454 VTAIL.n232 VTAIL.n183 0.155672
R1455 VTAIL.n232 VTAIL.n231 0.155672
R1456 VTAIL.n231 VTAIL.n187 0.155672
R1457 VTAIL.n224 VTAIL.n187 0.155672
R1458 VTAIL.n224 VTAIL.n223 0.155672
R1459 VTAIL.n223 VTAIL.n191 0.155672
R1460 VTAIL.n216 VTAIL.n191 0.155672
R1461 VTAIL.n216 VTAIL.n215 0.155672
R1462 VTAIL.n215 VTAIL.n195 0.155672
R1463 VTAIL.n208 VTAIL.n195 0.155672
R1464 VTAIL.n208 VTAIL.n207 0.155672
R1465 VTAIL.n207 VTAIL.n199 0.155672
R1466 VTAIL.n169 VTAIL.n87 0.155672
R1467 VTAIL.n162 VTAIL.n87 0.155672
R1468 VTAIL.n162 VTAIL.n161 0.155672
R1469 VTAIL.n161 VTAIL.n91 0.155672
R1470 VTAIL.n154 VTAIL.n91 0.155672
R1471 VTAIL.n154 VTAIL.n153 0.155672
R1472 VTAIL.n153 VTAIL.n97 0.155672
R1473 VTAIL.n146 VTAIL.n97 0.155672
R1474 VTAIL.n146 VTAIL.n145 0.155672
R1475 VTAIL.n145 VTAIL.n101 0.155672
R1476 VTAIL.n138 VTAIL.n101 0.155672
R1477 VTAIL.n138 VTAIL.n137 0.155672
R1478 VTAIL.n137 VTAIL.n105 0.155672
R1479 VTAIL.n130 VTAIL.n105 0.155672
R1480 VTAIL.n130 VTAIL.n129 0.155672
R1481 VTAIL.n129 VTAIL.n109 0.155672
R1482 VTAIL.n122 VTAIL.n109 0.155672
R1483 VTAIL.n122 VTAIL.n121 0.155672
R1484 VTAIL.n121 VTAIL.n113 0.155672
R1485 VDD1.n80 VDD1.n0 756.745
R1486 VDD1.n165 VDD1.n85 756.745
R1487 VDD1.n81 VDD1.n80 585
R1488 VDD1.n79 VDD1.n78 585
R1489 VDD1.n4 VDD1.n3 585
R1490 VDD1.n8 VDD1.n6 585
R1491 VDD1.n73 VDD1.n72 585
R1492 VDD1.n71 VDD1.n70 585
R1493 VDD1.n10 VDD1.n9 585
R1494 VDD1.n65 VDD1.n64 585
R1495 VDD1.n63 VDD1.n62 585
R1496 VDD1.n14 VDD1.n13 585
R1497 VDD1.n57 VDD1.n56 585
R1498 VDD1.n55 VDD1.n54 585
R1499 VDD1.n18 VDD1.n17 585
R1500 VDD1.n49 VDD1.n48 585
R1501 VDD1.n47 VDD1.n46 585
R1502 VDD1.n22 VDD1.n21 585
R1503 VDD1.n41 VDD1.n40 585
R1504 VDD1.n39 VDD1.n38 585
R1505 VDD1.n26 VDD1.n25 585
R1506 VDD1.n33 VDD1.n32 585
R1507 VDD1.n31 VDD1.n30 585
R1508 VDD1.n114 VDD1.n113 585
R1509 VDD1.n116 VDD1.n115 585
R1510 VDD1.n109 VDD1.n108 585
R1511 VDD1.n122 VDD1.n121 585
R1512 VDD1.n124 VDD1.n123 585
R1513 VDD1.n105 VDD1.n104 585
R1514 VDD1.n130 VDD1.n129 585
R1515 VDD1.n132 VDD1.n131 585
R1516 VDD1.n101 VDD1.n100 585
R1517 VDD1.n138 VDD1.n137 585
R1518 VDD1.n140 VDD1.n139 585
R1519 VDD1.n97 VDD1.n96 585
R1520 VDD1.n146 VDD1.n145 585
R1521 VDD1.n148 VDD1.n147 585
R1522 VDD1.n93 VDD1.n92 585
R1523 VDD1.n155 VDD1.n154 585
R1524 VDD1.n156 VDD1.n91 585
R1525 VDD1.n158 VDD1.n157 585
R1526 VDD1.n89 VDD1.n88 585
R1527 VDD1.n164 VDD1.n163 585
R1528 VDD1.n166 VDD1.n165 585
R1529 VDD1.n29 VDD1.t1 327.466
R1530 VDD1.n112 VDD1.t0 327.466
R1531 VDD1.n80 VDD1.n79 171.744
R1532 VDD1.n79 VDD1.n3 171.744
R1533 VDD1.n8 VDD1.n3 171.744
R1534 VDD1.n72 VDD1.n8 171.744
R1535 VDD1.n72 VDD1.n71 171.744
R1536 VDD1.n71 VDD1.n9 171.744
R1537 VDD1.n64 VDD1.n9 171.744
R1538 VDD1.n64 VDD1.n63 171.744
R1539 VDD1.n63 VDD1.n13 171.744
R1540 VDD1.n56 VDD1.n13 171.744
R1541 VDD1.n56 VDD1.n55 171.744
R1542 VDD1.n55 VDD1.n17 171.744
R1543 VDD1.n48 VDD1.n17 171.744
R1544 VDD1.n48 VDD1.n47 171.744
R1545 VDD1.n47 VDD1.n21 171.744
R1546 VDD1.n40 VDD1.n21 171.744
R1547 VDD1.n40 VDD1.n39 171.744
R1548 VDD1.n39 VDD1.n25 171.744
R1549 VDD1.n32 VDD1.n25 171.744
R1550 VDD1.n32 VDD1.n31 171.744
R1551 VDD1.n115 VDD1.n114 171.744
R1552 VDD1.n115 VDD1.n108 171.744
R1553 VDD1.n122 VDD1.n108 171.744
R1554 VDD1.n123 VDD1.n122 171.744
R1555 VDD1.n123 VDD1.n104 171.744
R1556 VDD1.n130 VDD1.n104 171.744
R1557 VDD1.n131 VDD1.n130 171.744
R1558 VDD1.n131 VDD1.n100 171.744
R1559 VDD1.n138 VDD1.n100 171.744
R1560 VDD1.n139 VDD1.n138 171.744
R1561 VDD1.n139 VDD1.n96 171.744
R1562 VDD1.n146 VDD1.n96 171.744
R1563 VDD1.n147 VDD1.n146 171.744
R1564 VDD1.n147 VDD1.n92 171.744
R1565 VDD1.n155 VDD1.n92 171.744
R1566 VDD1.n156 VDD1.n155 171.744
R1567 VDD1.n157 VDD1.n156 171.744
R1568 VDD1.n157 VDD1.n88 171.744
R1569 VDD1.n164 VDD1.n88 171.744
R1570 VDD1.n165 VDD1.n164 171.744
R1571 VDD1 VDD1.n169 91.5504
R1572 VDD1.n31 VDD1.t1 85.8723
R1573 VDD1.n114 VDD1.t0 85.8723
R1574 VDD1 VDD1.n84 50.364
R1575 VDD1.n30 VDD1.n29 16.3895
R1576 VDD1.n113 VDD1.n112 16.3895
R1577 VDD1.n6 VDD1.n4 13.1884
R1578 VDD1.n158 VDD1.n89 13.1884
R1579 VDD1.n78 VDD1.n77 12.8005
R1580 VDD1.n74 VDD1.n73 12.8005
R1581 VDD1.n33 VDD1.n28 12.8005
R1582 VDD1.n116 VDD1.n111 12.8005
R1583 VDD1.n159 VDD1.n91 12.8005
R1584 VDD1.n163 VDD1.n162 12.8005
R1585 VDD1.n81 VDD1.n2 12.0247
R1586 VDD1.n70 VDD1.n7 12.0247
R1587 VDD1.n34 VDD1.n26 12.0247
R1588 VDD1.n117 VDD1.n109 12.0247
R1589 VDD1.n154 VDD1.n153 12.0247
R1590 VDD1.n166 VDD1.n87 12.0247
R1591 VDD1.n82 VDD1.n0 11.249
R1592 VDD1.n69 VDD1.n10 11.249
R1593 VDD1.n38 VDD1.n37 11.249
R1594 VDD1.n121 VDD1.n120 11.249
R1595 VDD1.n152 VDD1.n93 11.249
R1596 VDD1.n167 VDD1.n85 11.249
R1597 VDD1.n66 VDD1.n65 10.4732
R1598 VDD1.n41 VDD1.n24 10.4732
R1599 VDD1.n124 VDD1.n107 10.4732
R1600 VDD1.n149 VDD1.n148 10.4732
R1601 VDD1.n62 VDD1.n12 9.69747
R1602 VDD1.n42 VDD1.n22 9.69747
R1603 VDD1.n125 VDD1.n105 9.69747
R1604 VDD1.n145 VDD1.n95 9.69747
R1605 VDD1.n84 VDD1.n83 9.45567
R1606 VDD1.n169 VDD1.n168 9.45567
R1607 VDD1.n16 VDD1.n15 9.3005
R1608 VDD1.n59 VDD1.n58 9.3005
R1609 VDD1.n61 VDD1.n60 9.3005
R1610 VDD1.n12 VDD1.n11 9.3005
R1611 VDD1.n67 VDD1.n66 9.3005
R1612 VDD1.n69 VDD1.n68 9.3005
R1613 VDD1.n7 VDD1.n5 9.3005
R1614 VDD1.n75 VDD1.n74 9.3005
R1615 VDD1.n83 VDD1.n82 9.3005
R1616 VDD1.n2 VDD1.n1 9.3005
R1617 VDD1.n77 VDD1.n76 9.3005
R1618 VDD1.n53 VDD1.n52 9.3005
R1619 VDD1.n51 VDD1.n50 9.3005
R1620 VDD1.n20 VDD1.n19 9.3005
R1621 VDD1.n45 VDD1.n44 9.3005
R1622 VDD1.n43 VDD1.n42 9.3005
R1623 VDD1.n24 VDD1.n23 9.3005
R1624 VDD1.n37 VDD1.n36 9.3005
R1625 VDD1.n35 VDD1.n34 9.3005
R1626 VDD1.n28 VDD1.n27 9.3005
R1627 VDD1.n168 VDD1.n167 9.3005
R1628 VDD1.n87 VDD1.n86 9.3005
R1629 VDD1.n162 VDD1.n161 9.3005
R1630 VDD1.n134 VDD1.n133 9.3005
R1631 VDD1.n103 VDD1.n102 9.3005
R1632 VDD1.n128 VDD1.n127 9.3005
R1633 VDD1.n126 VDD1.n125 9.3005
R1634 VDD1.n107 VDD1.n106 9.3005
R1635 VDD1.n120 VDD1.n119 9.3005
R1636 VDD1.n118 VDD1.n117 9.3005
R1637 VDD1.n111 VDD1.n110 9.3005
R1638 VDD1.n136 VDD1.n135 9.3005
R1639 VDD1.n99 VDD1.n98 9.3005
R1640 VDD1.n142 VDD1.n141 9.3005
R1641 VDD1.n144 VDD1.n143 9.3005
R1642 VDD1.n95 VDD1.n94 9.3005
R1643 VDD1.n150 VDD1.n149 9.3005
R1644 VDD1.n152 VDD1.n151 9.3005
R1645 VDD1.n153 VDD1.n90 9.3005
R1646 VDD1.n160 VDD1.n159 9.3005
R1647 VDD1.n61 VDD1.n14 8.92171
R1648 VDD1.n46 VDD1.n45 8.92171
R1649 VDD1.n129 VDD1.n128 8.92171
R1650 VDD1.n144 VDD1.n97 8.92171
R1651 VDD1.n58 VDD1.n57 8.14595
R1652 VDD1.n49 VDD1.n20 8.14595
R1653 VDD1.n132 VDD1.n103 8.14595
R1654 VDD1.n141 VDD1.n140 8.14595
R1655 VDD1.n54 VDD1.n16 7.3702
R1656 VDD1.n50 VDD1.n18 7.3702
R1657 VDD1.n133 VDD1.n101 7.3702
R1658 VDD1.n137 VDD1.n99 7.3702
R1659 VDD1.n54 VDD1.n53 6.59444
R1660 VDD1.n53 VDD1.n18 6.59444
R1661 VDD1.n136 VDD1.n101 6.59444
R1662 VDD1.n137 VDD1.n136 6.59444
R1663 VDD1.n57 VDD1.n16 5.81868
R1664 VDD1.n50 VDD1.n49 5.81868
R1665 VDD1.n133 VDD1.n132 5.81868
R1666 VDD1.n140 VDD1.n99 5.81868
R1667 VDD1.n58 VDD1.n14 5.04292
R1668 VDD1.n46 VDD1.n20 5.04292
R1669 VDD1.n129 VDD1.n103 5.04292
R1670 VDD1.n141 VDD1.n97 5.04292
R1671 VDD1.n62 VDD1.n61 4.26717
R1672 VDD1.n45 VDD1.n22 4.26717
R1673 VDD1.n128 VDD1.n105 4.26717
R1674 VDD1.n145 VDD1.n144 4.26717
R1675 VDD1.n29 VDD1.n27 3.70982
R1676 VDD1.n112 VDD1.n110 3.70982
R1677 VDD1.n65 VDD1.n12 3.49141
R1678 VDD1.n42 VDD1.n41 3.49141
R1679 VDD1.n125 VDD1.n124 3.49141
R1680 VDD1.n148 VDD1.n95 3.49141
R1681 VDD1.n84 VDD1.n0 2.71565
R1682 VDD1.n66 VDD1.n10 2.71565
R1683 VDD1.n38 VDD1.n24 2.71565
R1684 VDD1.n121 VDD1.n107 2.71565
R1685 VDD1.n149 VDD1.n93 2.71565
R1686 VDD1.n169 VDD1.n85 2.71565
R1687 VDD1.n82 VDD1.n81 1.93989
R1688 VDD1.n70 VDD1.n69 1.93989
R1689 VDD1.n37 VDD1.n26 1.93989
R1690 VDD1.n120 VDD1.n109 1.93989
R1691 VDD1.n154 VDD1.n152 1.93989
R1692 VDD1.n167 VDD1.n166 1.93989
R1693 VDD1.n78 VDD1.n2 1.16414
R1694 VDD1.n73 VDD1.n7 1.16414
R1695 VDD1.n34 VDD1.n33 1.16414
R1696 VDD1.n117 VDD1.n116 1.16414
R1697 VDD1.n153 VDD1.n91 1.16414
R1698 VDD1.n163 VDD1.n87 1.16414
R1699 VDD1.n77 VDD1.n4 0.388379
R1700 VDD1.n74 VDD1.n6 0.388379
R1701 VDD1.n30 VDD1.n28 0.388379
R1702 VDD1.n113 VDD1.n111 0.388379
R1703 VDD1.n159 VDD1.n158 0.388379
R1704 VDD1.n162 VDD1.n89 0.388379
R1705 VDD1.n83 VDD1.n1 0.155672
R1706 VDD1.n76 VDD1.n1 0.155672
R1707 VDD1.n76 VDD1.n75 0.155672
R1708 VDD1.n75 VDD1.n5 0.155672
R1709 VDD1.n68 VDD1.n5 0.155672
R1710 VDD1.n68 VDD1.n67 0.155672
R1711 VDD1.n67 VDD1.n11 0.155672
R1712 VDD1.n60 VDD1.n11 0.155672
R1713 VDD1.n60 VDD1.n59 0.155672
R1714 VDD1.n59 VDD1.n15 0.155672
R1715 VDD1.n52 VDD1.n15 0.155672
R1716 VDD1.n52 VDD1.n51 0.155672
R1717 VDD1.n51 VDD1.n19 0.155672
R1718 VDD1.n44 VDD1.n19 0.155672
R1719 VDD1.n44 VDD1.n43 0.155672
R1720 VDD1.n43 VDD1.n23 0.155672
R1721 VDD1.n36 VDD1.n23 0.155672
R1722 VDD1.n36 VDD1.n35 0.155672
R1723 VDD1.n35 VDD1.n27 0.155672
R1724 VDD1.n118 VDD1.n110 0.155672
R1725 VDD1.n119 VDD1.n118 0.155672
R1726 VDD1.n119 VDD1.n106 0.155672
R1727 VDD1.n126 VDD1.n106 0.155672
R1728 VDD1.n127 VDD1.n126 0.155672
R1729 VDD1.n127 VDD1.n102 0.155672
R1730 VDD1.n134 VDD1.n102 0.155672
R1731 VDD1.n135 VDD1.n134 0.155672
R1732 VDD1.n135 VDD1.n98 0.155672
R1733 VDD1.n142 VDD1.n98 0.155672
R1734 VDD1.n143 VDD1.n142 0.155672
R1735 VDD1.n143 VDD1.n94 0.155672
R1736 VDD1.n150 VDD1.n94 0.155672
R1737 VDD1.n151 VDD1.n150 0.155672
R1738 VDD1.n151 VDD1.n90 0.155672
R1739 VDD1.n160 VDD1.n90 0.155672
R1740 VDD1.n161 VDD1.n160 0.155672
R1741 VDD1.n161 VDD1.n86 0.155672
R1742 VDD1.n168 VDD1.n86 0.155672
R1743 VN VN.t0 303.997
R1744 VN VN.t1 258.769
R1745 VDD2.n165 VDD2.n85 756.745
R1746 VDD2.n80 VDD2.n0 756.745
R1747 VDD2.n166 VDD2.n165 585
R1748 VDD2.n164 VDD2.n163 585
R1749 VDD2.n89 VDD2.n88 585
R1750 VDD2.n93 VDD2.n91 585
R1751 VDD2.n158 VDD2.n157 585
R1752 VDD2.n156 VDD2.n155 585
R1753 VDD2.n95 VDD2.n94 585
R1754 VDD2.n150 VDD2.n149 585
R1755 VDD2.n148 VDD2.n147 585
R1756 VDD2.n99 VDD2.n98 585
R1757 VDD2.n142 VDD2.n141 585
R1758 VDD2.n140 VDD2.n139 585
R1759 VDD2.n103 VDD2.n102 585
R1760 VDD2.n134 VDD2.n133 585
R1761 VDD2.n132 VDD2.n131 585
R1762 VDD2.n107 VDD2.n106 585
R1763 VDD2.n126 VDD2.n125 585
R1764 VDD2.n124 VDD2.n123 585
R1765 VDD2.n111 VDD2.n110 585
R1766 VDD2.n118 VDD2.n117 585
R1767 VDD2.n116 VDD2.n115 585
R1768 VDD2.n29 VDD2.n28 585
R1769 VDD2.n31 VDD2.n30 585
R1770 VDD2.n24 VDD2.n23 585
R1771 VDD2.n37 VDD2.n36 585
R1772 VDD2.n39 VDD2.n38 585
R1773 VDD2.n20 VDD2.n19 585
R1774 VDD2.n45 VDD2.n44 585
R1775 VDD2.n47 VDD2.n46 585
R1776 VDD2.n16 VDD2.n15 585
R1777 VDD2.n53 VDD2.n52 585
R1778 VDD2.n55 VDD2.n54 585
R1779 VDD2.n12 VDD2.n11 585
R1780 VDD2.n61 VDD2.n60 585
R1781 VDD2.n63 VDD2.n62 585
R1782 VDD2.n8 VDD2.n7 585
R1783 VDD2.n70 VDD2.n69 585
R1784 VDD2.n71 VDD2.n6 585
R1785 VDD2.n73 VDD2.n72 585
R1786 VDD2.n4 VDD2.n3 585
R1787 VDD2.n79 VDD2.n78 585
R1788 VDD2.n81 VDD2.n80 585
R1789 VDD2.n114 VDD2.t1 327.466
R1790 VDD2.n27 VDD2.t0 327.466
R1791 VDD2.n165 VDD2.n164 171.744
R1792 VDD2.n164 VDD2.n88 171.744
R1793 VDD2.n93 VDD2.n88 171.744
R1794 VDD2.n157 VDD2.n93 171.744
R1795 VDD2.n157 VDD2.n156 171.744
R1796 VDD2.n156 VDD2.n94 171.744
R1797 VDD2.n149 VDD2.n94 171.744
R1798 VDD2.n149 VDD2.n148 171.744
R1799 VDD2.n148 VDD2.n98 171.744
R1800 VDD2.n141 VDD2.n98 171.744
R1801 VDD2.n141 VDD2.n140 171.744
R1802 VDD2.n140 VDD2.n102 171.744
R1803 VDD2.n133 VDD2.n102 171.744
R1804 VDD2.n133 VDD2.n132 171.744
R1805 VDD2.n132 VDD2.n106 171.744
R1806 VDD2.n125 VDD2.n106 171.744
R1807 VDD2.n125 VDD2.n124 171.744
R1808 VDD2.n124 VDD2.n110 171.744
R1809 VDD2.n117 VDD2.n110 171.744
R1810 VDD2.n117 VDD2.n116 171.744
R1811 VDD2.n30 VDD2.n29 171.744
R1812 VDD2.n30 VDD2.n23 171.744
R1813 VDD2.n37 VDD2.n23 171.744
R1814 VDD2.n38 VDD2.n37 171.744
R1815 VDD2.n38 VDD2.n19 171.744
R1816 VDD2.n45 VDD2.n19 171.744
R1817 VDD2.n46 VDD2.n45 171.744
R1818 VDD2.n46 VDD2.n15 171.744
R1819 VDD2.n53 VDD2.n15 171.744
R1820 VDD2.n54 VDD2.n53 171.744
R1821 VDD2.n54 VDD2.n11 171.744
R1822 VDD2.n61 VDD2.n11 171.744
R1823 VDD2.n62 VDD2.n61 171.744
R1824 VDD2.n62 VDD2.n7 171.744
R1825 VDD2.n70 VDD2.n7 171.744
R1826 VDD2.n71 VDD2.n70 171.744
R1827 VDD2.n72 VDD2.n71 171.744
R1828 VDD2.n72 VDD2.n3 171.744
R1829 VDD2.n79 VDD2.n3 171.744
R1830 VDD2.n80 VDD2.n79 171.744
R1831 VDD2.n170 VDD2.n84 90.5536
R1832 VDD2.n116 VDD2.t1 85.8723
R1833 VDD2.n29 VDD2.t0 85.8723
R1834 VDD2.n170 VDD2.n169 49.8338
R1835 VDD2.n115 VDD2.n114 16.3895
R1836 VDD2.n28 VDD2.n27 16.3895
R1837 VDD2.n91 VDD2.n89 13.1884
R1838 VDD2.n73 VDD2.n4 13.1884
R1839 VDD2.n163 VDD2.n162 12.8005
R1840 VDD2.n159 VDD2.n158 12.8005
R1841 VDD2.n118 VDD2.n113 12.8005
R1842 VDD2.n31 VDD2.n26 12.8005
R1843 VDD2.n74 VDD2.n6 12.8005
R1844 VDD2.n78 VDD2.n77 12.8005
R1845 VDD2.n166 VDD2.n87 12.0247
R1846 VDD2.n155 VDD2.n92 12.0247
R1847 VDD2.n119 VDD2.n111 12.0247
R1848 VDD2.n32 VDD2.n24 12.0247
R1849 VDD2.n69 VDD2.n68 12.0247
R1850 VDD2.n81 VDD2.n2 12.0247
R1851 VDD2.n167 VDD2.n85 11.249
R1852 VDD2.n154 VDD2.n95 11.249
R1853 VDD2.n123 VDD2.n122 11.249
R1854 VDD2.n36 VDD2.n35 11.249
R1855 VDD2.n67 VDD2.n8 11.249
R1856 VDD2.n82 VDD2.n0 11.249
R1857 VDD2.n151 VDD2.n150 10.4732
R1858 VDD2.n126 VDD2.n109 10.4732
R1859 VDD2.n39 VDD2.n22 10.4732
R1860 VDD2.n64 VDD2.n63 10.4732
R1861 VDD2.n147 VDD2.n97 9.69747
R1862 VDD2.n127 VDD2.n107 9.69747
R1863 VDD2.n40 VDD2.n20 9.69747
R1864 VDD2.n60 VDD2.n10 9.69747
R1865 VDD2.n169 VDD2.n168 9.45567
R1866 VDD2.n84 VDD2.n83 9.45567
R1867 VDD2.n101 VDD2.n100 9.3005
R1868 VDD2.n144 VDD2.n143 9.3005
R1869 VDD2.n146 VDD2.n145 9.3005
R1870 VDD2.n97 VDD2.n96 9.3005
R1871 VDD2.n152 VDD2.n151 9.3005
R1872 VDD2.n154 VDD2.n153 9.3005
R1873 VDD2.n92 VDD2.n90 9.3005
R1874 VDD2.n160 VDD2.n159 9.3005
R1875 VDD2.n168 VDD2.n167 9.3005
R1876 VDD2.n87 VDD2.n86 9.3005
R1877 VDD2.n162 VDD2.n161 9.3005
R1878 VDD2.n138 VDD2.n137 9.3005
R1879 VDD2.n136 VDD2.n135 9.3005
R1880 VDD2.n105 VDD2.n104 9.3005
R1881 VDD2.n130 VDD2.n129 9.3005
R1882 VDD2.n128 VDD2.n127 9.3005
R1883 VDD2.n109 VDD2.n108 9.3005
R1884 VDD2.n122 VDD2.n121 9.3005
R1885 VDD2.n120 VDD2.n119 9.3005
R1886 VDD2.n113 VDD2.n112 9.3005
R1887 VDD2.n83 VDD2.n82 9.3005
R1888 VDD2.n2 VDD2.n1 9.3005
R1889 VDD2.n77 VDD2.n76 9.3005
R1890 VDD2.n49 VDD2.n48 9.3005
R1891 VDD2.n18 VDD2.n17 9.3005
R1892 VDD2.n43 VDD2.n42 9.3005
R1893 VDD2.n41 VDD2.n40 9.3005
R1894 VDD2.n22 VDD2.n21 9.3005
R1895 VDD2.n35 VDD2.n34 9.3005
R1896 VDD2.n33 VDD2.n32 9.3005
R1897 VDD2.n26 VDD2.n25 9.3005
R1898 VDD2.n51 VDD2.n50 9.3005
R1899 VDD2.n14 VDD2.n13 9.3005
R1900 VDD2.n57 VDD2.n56 9.3005
R1901 VDD2.n59 VDD2.n58 9.3005
R1902 VDD2.n10 VDD2.n9 9.3005
R1903 VDD2.n65 VDD2.n64 9.3005
R1904 VDD2.n67 VDD2.n66 9.3005
R1905 VDD2.n68 VDD2.n5 9.3005
R1906 VDD2.n75 VDD2.n74 9.3005
R1907 VDD2.n146 VDD2.n99 8.92171
R1908 VDD2.n131 VDD2.n130 8.92171
R1909 VDD2.n44 VDD2.n43 8.92171
R1910 VDD2.n59 VDD2.n12 8.92171
R1911 VDD2.n143 VDD2.n142 8.14595
R1912 VDD2.n134 VDD2.n105 8.14595
R1913 VDD2.n47 VDD2.n18 8.14595
R1914 VDD2.n56 VDD2.n55 8.14595
R1915 VDD2.n139 VDD2.n101 7.3702
R1916 VDD2.n135 VDD2.n103 7.3702
R1917 VDD2.n48 VDD2.n16 7.3702
R1918 VDD2.n52 VDD2.n14 7.3702
R1919 VDD2.n139 VDD2.n138 6.59444
R1920 VDD2.n138 VDD2.n103 6.59444
R1921 VDD2.n51 VDD2.n16 6.59444
R1922 VDD2.n52 VDD2.n51 6.59444
R1923 VDD2.n142 VDD2.n101 5.81868
R1924 VDD2.n135 VDD2.n134 5.81868
R1925 VDD2.n48 VDD2.n47 5.81868
R1926 VDD2.n55 VDD2.n14 5.81868
R1927 VDD2.n143 VDD2.n99 5.04292
R1928 VDD2.n131 VDD2.n105 5.04292
R1929 VDD2.n44 VDD2.n18 5.04292
R1930 VDD2.n56 VDD2.n12 5.04292
R1931 VDD2.n147 VDD2.n146 4.26717
R1932 VDD2.n130 VDD2.n107 4.26717
R1933 VDD2.n43 VDD2.n20 4.26717
R1934 VDD2.n60 VDD2.n59 4.26717
R1935 VDD2.n114 VDD2.n112 3.70982
R1936 VDD2.n27 VDD2.n25 3.70982
R1937 VDD2.n150 VDD2.n97 3.49141
R1938 VDD2.n127 VDD2.n126 3.49141
R1939 VDD2.n40 VDD2.n39 3.49141
R1940 VDD2.n63 VDD2.n10 3.49141
R1941 VDD2.n169 VDD2.n85 2.71565
R1942 VDD2.n151 VDD2.n95 2.71565
R1943 VDD2.n123 VDD2.n109 2.71565
R1944 VDD2.n36 VDD2.n22 2.71565
R1945 VDD2.n64 VDD2.n8 2.71565
R1946 VDD2.n84 VDD2.n0 2.71565
R1947 VDD2.n167 VDD2.n166 1.93989
R1948 VDD2.n155 VDD2.n154 1.93989
R1949 VDD2.n122 VDD2.n111 1.93989
R1950 VDD2.n35 VDD2.n24 1.93989
R1951 VDD2.n69 VDD2.n67 1.93989
R1952 VDD2.n82 VDD2.n81 1.93989
R1953 VDD2.n163 VDD2.n87 1.16414
R1954 VDD2.n158 VDD2.n92 1.16414
R1955 VDD2.n119 VDD2.n118 1.16414
R1956 VDD2.n32 VDD2.n31 1.16414
R1957 VDD2.n68 VDD2.n6 1.16414
R1958 VDD2.n78 VDD2.n2 1.16414
R1959 VDD2 VDD2.n170 0.530672
R1960 VDD2.n162 VDD2.n89 0.388379
R1961 VDD2.n159 VDD2.n91 0.388379
R1962 VDD2.n115 VDD2.n113 0.388379
R1963 VDD2.n28 VDD2.n26 0.388379
R1964 VDD2.n74 VDD2.n73 0.388379
R1965 VDD2.n77 VDD2.n4 0.388379
R1966 VDD2.n168 VDD2.n86 0.155672
R1967 VDD2.n161 VDD2.n86 0.155672
R1968 VDD2.n161 VDD2.n160 0.155672
R1969 VDD2.n160 VDD2.n90 0.155672
R1970 VDD2.n153 VDD2.n90 0.155672
R1971 VDD2.n153 VDD2.n152 0.155672
R1972 VDD2.n152 VDD2.n96 0.155672
R1973 VDD2.n145 VDD2.n96 0.155672
R1974 VDD2.n145 VDD2.n144 0.155672
R1975 VDD2.n144 VDD2.n100 0.155672
R1976 VDD2.n137 VDD2.n100 0.155672
R1977 VDD2.n137 VDD2.n136 0.155672
R1978 VDD2.n136 VDD2.n104 0.155672
R1979 VDD2.n129 VDD2.n104 0.155672
R1980 VDD2.n129 VDD2.n128 0.155672
R1981 VDD2.n128 VDD2.n108 0.155672
R1982 VDD2.n121 VDD2.n108 0.155672
R1983 VDD2.n121 VDD2.n120 0.155672
R1984 VDD2.n120 VDD2.n112 0.155672
R1985 VDD2.n33 VDD2.n25 0.155672
R1986 VDD2.n34 VDD2.n33 0.155672
R1987 VDD2.n34 VDD2.n21 0.155672
R1988 VDD2.n41 VDD2.n21 0.155672
R1989 VDD2.n42 VDD2.n41 0.155672
R1990 VDD2.n42 VDD2.n17 0.155672
R1991 VDD2.n49 VDD2.n17 0.155672
R1992 VDD2.n50 VDD2.n49 0.155672
R1993 VDD2.n50 VDD2.n13 0.155672
R1994 VDD2.n57 VDD2.n13 0.155672
R1995 VDD2.n58 VDD2.n57 0.155672
R1996 VDD2.n58 VDD2.n9 0.155672
R1997 VDD2.n65 VDD2.n9 0.155672
R1998 VDD2.n66 VDD2.n65 0.155672
R1999 VDD2.n66 VDD2.n5 0.155672
R2000 VDD2.n75 VDD2.n5 0.155672
R2001 VDD2.n76 VDD2.n75 0.155672
R2002 VDD2.n76 VDD2.n1 0.155672
R2003 VDD2.n83 VDD2.n1 0.155672
C0 VDD1 VTAIL 5.98375f
C1 VN VP 5.73993f
C2 VDD2 VN 3.29501f
C3 w_n1846_n4050# VP 2.78385f
C4 VDD2 w_n1846_n4050# 1.95634f
C5 B VP 1.34587f
C6 VTAIL VN 2.75722f
C7 VDD2 B 1.88969f
C8 VTAIL w_n1846_n4050# 3.28062f
C9 VDD1 VN 0.147783f
C10 B VTAIL 4.0532f
C11 VDD2 VP 0.302388f
C12 VDD1 w_n1846_n4050# 1.93936f
C13 VTAIL VP 2.77166f
C14 B VDD1 1.86615f
C15 VDD2 VTAIL 6.02733f
C16 w_n1846_n4050# VN 2.55031f
C17 VDD1 VP 3.44585f
C18 VDD2 VDD1 0.587653f
C19 B VN 0.964869f
C20 B w_n1846_n4050# 8.96564f
C21 VDD2 VSUBS 0.93791f
C22 VDD1 VSUBS 3.81813f
C23 VTAIL VSUBS 1.04907f
C24 VN VSUBS 8.47543f
C25 VP VSUBS 1.59288f
C26 B VSUBS 3.632232f
C27 w_n1846_n4050# VSUBS 91.6428f
C28 VDD2.n0 VSUBS 0.020937f
C29 VDD2.n1 VSUBS 0.019978f
C30 VDD2.n2 VSUBS 0.010735f
C31 VDD2.n3 VSUBS 0.025375f
C32 VDD2.n4 VSUBS 0.011051f
C33 VDD2.n5 VSUBS 0.019978f
C34 VDD2.n6 VSUBS 0.011367f
C35 VDD2.n7 VSUBS 0.025375f
C36 VDD2.n8 VSUBS 0.011367f
C37 VDD2.n9 VSUBS 0.019978f
C38 VDD2.n10 VSUBS 0.010735f
C39 VDD2.n11 VSUBS 0.025375f
C40 VDD2.n12 VSUBS 0.011367f
C41 VDD2.n13 VSUBS 0.019978f
C42 VDD2.n14 VSUBS 0.010735f
C43 VDD2.n15 VSUBS 0.025375f
C44 VDD2.n16 VSUBS 0.011367f
C45 VDD2.n17 VSUBS 0.019978f
C46 VDD2.n18 VSUBS 0.010735f
C47 VDD2.n19 VSUBS 0.025375f
C48 VDD2.n20 VSUBS 0.011367f
C49 VDD2.n21 VSUBS 0.019978f
C50 VDD2.n22 VSUBS 0.010735f
C51 VDD2.n23 VSUBS 0.025375f
C52 VDD2.n24 VSUBS 0.011367f
C53 VDD2.n25 VSUBS 1.31284f
C54 VDD2.n26 VSUBS 0.010735f
C55 VDD2.t0 VSUBS 0.054342f
C56 VDD2.n27 VSUBS 0.143245f
C57 VDD2.n28 VSUBS 0.016142f
C58 VDD2.n29 VSUBS 0.019031f
C59 VDD2.n30 VSUBS 0.025375f
C60 VDD2.n31 VSUBS 0.011367f
C61 VDD2.n32 VSUBS 0.010735f
C62 VDD2.n33 VSUBS 0.019978f
C63 VDD2.n34 VSUBS 0.019978f
C64 VDD2.n35 VSUBS 0.010735f
C65 VDD2.n36 VSUBS 0.011367f
C66 VDD2.n37 VSUBS 0.025375f
C67 VDD2.n38 VSUBS 0.025375f
C68 VDD2.n39 VSUBS 0.011367f
C69 VDD2.n40 VSUBS 0.010735f
C70 VDD2.n41 VSUBS 0.019978f
C71 VDD2.n42 VSUBS 0.019978f
C72 VDD2.n43 VSUBS 0.010735f
C73 VDD2.n44 VSUBS 0.011367f
C74 VDD2.n45 VSUBS 0.025375f
C75 VDD2.n46 VSUBS 0.025375f
C76 VDD2.n47 VSUBS 0.011367f
C77 VDD2.n48 VSUBS 0.010735f
C78 VDD2.n49 VSUBS 0.019978f
C79 VDD2.n50 VSUBS 0.019978f
C80 VDD2.n51 VSUBS 0.010735f
C81 VDD2.n52 VSUBS 0.011367f
C82 VDD2.n53 VSUBS 0.025375f
C83 VDD2.n54 VSUBS 0.025375f
C84 VDD2.n55 VSUBS 0.011367f
C85 VDD2.n56 VSUBS 0.010735f
C86 VDD2.n57 VSUBS 0.019978f
C87 VDD2.n58 VSUBS 0.019978f
C88 VDD2.n59 VSUBS 0.010735f
C89 VDD2.n60 VSUBS 0.011367f
C90 VDD2.n61 VSUBS 0.025375f
C91 VDD2.n62 VSUBS 0.025375f
C92 VDD2.n63 VSUBS 0.011367f
C93 VDD2.n64 VSUBS 0.010735f
C94 VDD2.n65 VSUBS 0.019978f
C95 VDD2.n66 VSUBS 0.019978f
C96 VDD2.n67 VSUBS 0.010735f
C97 VDD2.n68 VSUBS 0.010735f
C98 VDD2.n69 VSUBS 0.011367f
C99 VDD2.n70 VSUBS 0.025375f
C100 VDD2.n71 VSUBS 0.025375f
C101 VDD2.n72 VSUBS 0.025375f
C102 VDD2.n73 VSUBS 0.011051f
C103 VDD2.n74 VSUBS 0.010735f
C104 VDD2.n75 VSUBS 0.019978f
C105 VDD2.n76 VSUBS 0.019978f
C106 VDD2.n77 VSUBS 0.010735f
C107 VDD2.n78 VSUBS 0.011367f
C108 VDD2.n79 VSUBS 0.025375f
C109 VDD2.n80 VSUBS 0.057972f
C110 VDD2.n81 VSUBS 0.011367f
C111 VDD2.n82 VSUBS 0.010735f
C112 VDD2.n83 VSUBS 0.047543f
C113 VDD2.n84 VSUBS 0.638776f
C114 VDD2.n85 VSUBS 0.020937f
C115 VDD2.n86 VSUBS 0.019978f
C116 VDD2.n87 VSUBS 0.010735f
C117 VDD2.n88 VSUBS 0.025375f
C118 VDD2.n89 VSUBS 0.011051f
C119 VDD2.n90 VSUBS 0.019978f
C120 VDD2.n91 VSUBS 0.011051f
C121 VDD2.n92 VSUBS 0.010735f
C122 VDD2.n93 VSUBS 0.025375f
C123 VDD2.n94 VSUBS 0.025375f
C124 VDD2.n95 VSUBS 0.011367f
C125 VDD2.n96 VSUBS 0.019978f
C126 VDD2.n97 VSUBS 0.010735f
C127 VDD2.n98 VSUBS 0.025375f
C128 VDD2.n99 VSUBS 0.011367f
C129 VDD2.n100 VSUBS 0.019978f
C130 VDD2.n101 VSUBS 0.010735f
C131 VDD2.n102 VSUBS 0.025375f
C132 VDD2.n103 VSUBS 0.011367f
C133 VDD2.n104 VSUBS 0.019978f
C134 VDD2.n105 VSUBS 0.010735f
C135 VDD2.n106 VSUBS 0.025375f
C136 VDD2.n107 VSUBS 0.011367f
C137 VDD2.n108 VSUBS 0.019978f
C138 VDD2.n109 VSUBS 0.010735f
C139 VDD2.n110 VSUBS 0.025375f
C140 VDD2.n111 VSUBS 0.011367f
C141 VDD2.n112 VSUBS 1.31284f
C142 VDD2.n113 VSUBS 0.010735f
C143 VDD2.t1 VSUBS 0.054342f
C144 VDD2.n114 VSUBS 0.143245f
C145 VDD2.n115 VSUBS 0.016142f
C146 VDD2.n116 VSUBS 0.019031f
C147 VDD2.n117 VSUBS 0.025375f
C148 VDD2.n118 VSUBS 0.011367f
C149 VDD2.n119 VSUBS 0.010735f
C150 VDD2.n120 VSUBS 0.019978f
C151 VDD2.n121 VSUBS 0.019978f
C152 VDD2.n122 VSUBS 0.010735f
C153 VDD2.n123 VSUBS 0.011367f
C154 VDD2.n124 VSUBS 0.025375f
C155 VDD2.n125 VSUBS 0.025375f
C156 VDD2.n126 VSUBS 0.011367f
C157 VDD2.n127 VSUBS 0.010735f
C158 VDD2.n128 VSUBS 0.019978f
C159 VDD2.n129 VSUBS 0.019978f
C160 VDD2.n130 VSUBS 0.010735f
C161 VDD2.n131 VSUBS 0.011367f
C162 VDD2.n132 VSUBS 0.025375f
C163 VDD2.n133 VSUBS 0.025375f
C164 VDD2.n134 VSUBS 0.011367f
C165 VDD2.n135 VSUBS 0.010735f
C166 VDD2.n136 VSUBS 0.019978f
C167 VDD2.n137 VSUBS 0.019978f
C168 VDD2.n138 VSUBS 0.010735f
C169 VDD2.n139 VSUBS 0.011367f
C170 VDD2.n140 VSUBS 0.025375f
C171 VDD2.n141 VSUBS 0.025375f
C172 VDD2.n142 VSUBS 0.011367f
C173 VDD2.n143 VSUBS 0.010735f
C174 VDD2.n144 VSUBS 0.019978f
C175 VDD2.n145 VSUBS 0.019978f
C176 VDD2.n146 VSUBS 0.010735f
C177 VDD2.n147 VSUBS 0.011367f
C178 VDD2.n148 VSUBS 0.025375f
C179 VDD2.n149 VSUBS 0.025375f
C180 VDD2.n150 VSUBS 0.011367f
C181 VDD2.n151 VSUBS 0.010735f
C182 VDD2.n152 VSUBS 0.019978f
C183 VDD2.n153 VSUBS 0.019978f
C184 VDD2.n154 VSUBS 0.010735f
C185 VDD2.n155 VSUBS 0.011367f
C186 VDD2.n156 VSUBS 0.025375f
C187 VDD2.n157 VSUBS 0.025375f
C188 VDD2.n158 VSUBS 0.011367f
C189 VDD2.n159 VSUBS 0.010735f
C190 VDD2.n160 VSUBS 0.019978f
C191 VDD2.n161 VSUBS 0.019978f
C192 VDD2.n162 VSUBS 0.010735f
C193 VDD2.n163 VSUBS 0.011367f
C194 VDD2.n164 VSUBS 0.025375f
C195 VDD2.n165 VSUBS 0.057972f
C196 VDD2.n166 VSUBS 0.011367f
C197 VDD2.n167 VSUBS 0.010735f
C198 VDD2.n168 VSUBS 0.047543f
C199 VDD2.n169 VSUBS 0.042825f
C200 VDD2.n170 VSUBS 2.61256f
C201 VN.t1 VSUBS 3.83701f
C202 VN.t0 VSUBS 4.3347f
C203 VDD1.n0 VSUBS 0.020995f
C204 VDD1.n1 VSUBS 0.020034f
C205 VDD1.n2 VSUBS 0.010766f
C206 VDD1.n3 VSUBS 0.025446f
C207 VDD1.n4 VSUBS 0.011082f
C208 VDD1.n5 VSUBS 0.020034f
C209 VDD1.n6 VSUBS 0.011082f
C210 VDD1.n7 VSUBS 0.010766f
C211 VDD1.n8 VSUBS 0.025446f
C212 VDD1.n9 VSUBS 0.025446f
C213 VDD1.n10 VSUBS 0.011399f
C214 VDD1.n11 VSUBS 0.020034f
C215 VDD1.n12 VSUBS 0.010766f
C216 VDD1.n13 VSUBS 0.025446f
C217 VDD1.n14 VSUBS 0.011399f
C218 VDD1.n15 VSUBS 0.020034f
C219 VDD1.n16 VSUBS 0.010766f
C220 VDD1.n17 VSUBS 0.025446f
C221 VDD1.n18 VSUBS 0.011399f
C222 VDD1.n19 VSUBS 0.020034f
C223 VDD1.n20 VSUBS 0.010766f
C224 VDD1.n21 VSUBS 0.025446f
C225 VDD1.n22 VSUBS 0.011399f
C226 VDD1.n23 VSUBS 0.020034f
C227 VDD1.n24 VSUBS 0.010766f
C228 VDD1.n25 VSUBS 0.025446f
C229 VDD1.n26 VSUBS 0.011399f
C230 VDD1.n27 VSUBS 1.31651f
C231 VDD1.n28 VSUBS 0.010766f
C232 VDD1.t1 VSUBS 0.054494f
C233 VDD1.n29 VSUBS 0.143646f
C234 VDD1.n30 VSUBS 0.016187f
C235 VDD1.n31 VSUBS 0.019084f
C236 VDD1.n32 VSUBS 0.025446f
C237 VDD1.n33 VSUBS 0.011399f
C238 VDD1.n34 VSUBS 0.010766f
C239 VDD1.n35 VSUBS 0.020034f
C240 VDD1.n36 VSUBS 0.020034f
C241 VDD1.n37 VSUBS 0.010766f
C242 VDD1.n38 VSUBS 0.011399f
C243 VDD1.n39 VSUBS 0.025446f
C244 VDD1.n40 VSUBS 0.025446f
C245 VDD1.n41 VSUBS 0.011399f
C246 VDD1.n42 VSUBS 0.010766f
C247 VDD1.n43 VSUBS 0.020034f
C248 VDD1.n44 VSUBS 0.020034f
C249 VDD1.n45 VSUBS 0.010766f
C250 VDD1.n46 VSUBS 0.011399f
C251 VDD1.n47 VSUBS 0.025446f
C252 VDD1.n48 VSUBS 0.025446f
C253 VDD1.n49 VSUBS 0.011399f
C254 VDD1.n50 VSUBS 0.010766f
C255 VDD1.n51 VSUBS 0.020034f
C256 VDD1.n52 VSUBS 0.020034f
C257 VDD1.n53 VSUBS 0.010766f
C258 VDD1.n54 VSUBS 0.011399f
C259 VDD1.n55 VSUBS 0.025446f
C260 VDD1.n56 VSUBS 0.025446f
C261 VDD1.n57 VSUBS 0.011399f
C262 VDD1.n58 VSUBS 0.010766f
C263 VDD1.n59 VSUBS 0.020034f
C264 VDD1.n60 VSUBS 0.020034f
C265 VDD1.n61 VSUBS 0.010766f
C266 VDD1.n62 VSUBS 0.011399f
C267 VDD1.n63 VSUBS 0.025446f
C268 VDD1.n64 VSUBS 0.025446f
C269 VDD1.n65 VSUBS 0.011399f
C270 VDD1.n66 VSUBS 0.010766f
C271 VDD1.n67 VSUBS 0.020034f
C272 VDD1.n68 VSUBS 0.020034f
C273 VDD1.n69 VSUBS 0.010766f
C274 VDD1.n70 VSUBS 0.011399f
C275 VDD1.n71 VSUBS 0.025446f
C276 VDD1.n72 VSUBS 0.025446f
C277 VDD1.n73 VSUBS 0.011399f
C278 VDD1.n74 VSUBS 0.010766f
C279 VDD1.n75 VSUBS 0.020034f
C280 VDD1.n76 VSUBS 0.020034f
C281 VDD1.n77 VSUBS 0.010766f
C282 VDD1.n78 VSUBS 0.011399f
C283 VDD1.n79 VSUBS 0.025446f
C284 VDD1.n80 VSUBS 0.058134f
C285 VDD1.n81 VSUBS 0.011399f
C286 VDD1.n82 VSUBS 0.010766f
C287 VDD1.n83 VSUBS 0.047676f
C288 VDD1.n84 VSUBS 0.04372f
C289 VDD1.n85 VSUBS 0.020995f
C290 VDD1.n86 VSUBS 0.020034f
C291 VDD1.n87 VSUBS 0.010766f
C292 VDD1.n88 VSUBS 0.025446f
C293 VDD1.n89 VSUBS 0.011082f
C294 VDD1.n90 VSUBS 0.020034f
C295 VDD1.n91 VSUBS 0.011399f
C296 VDD1.n92 VSUBS 0.025446f
C297 VDD1.n93 VSUBS 0.011399f
C298 VDD1.n94 VSUBS 0.020034f
C299 VDD1.n95 VSUBS 0.010766f
C300 VDD1.n96 VSUBS 0.025446f
C301 VDD1.n97 VSUBS 0.011399f
C302 VDD1.n98 VSUBS 0.020034f
C303 VDD1.n99 VSUBS 0.010766f
C304 VDD1.n100 VSUBS 0.025446f
C305 VDD1.n101 VSUBS 0.011399f
C306 VDD1.n102 VSUBS 0.020034f
C307 VDD1.n103 VSUBS 0.010766f
C308 VDD1.n104 VSUBS 0.025446f
C309 VDD1.n105 VSUBS 0.011399f
C310 VDD1.n106 VSUBS 0.020034f
C311 VDD1.n107 VSUBS 0.010766f
C312 VDD1.n108 VSUBS 0.025446f
C313 VDD1.n109 VSUBS 0.011399f
C314 VDD1.n110 VSUBS 1.31651f
C315 VDD1.n111 VSUBS 0.010766f
C316 VDD1.t0 VSUBS 0.054494f
C317 VDD1.n112 VSUBS 0.143646f
C318 VDD1.n113 VSUBS 0.016187f
C319 VDD1.n114 VSUBS 0.019084f
C320 VDD1.n115 VSUBS 0.025446f
C321 VDD1.n116 VSUBS 0.011399f
C322 VDD1.n117 VSUBS 0.010766f
C323 VDD1.n118 VSUBS 0.020034f
C324 VDD1.n119 VSUBS 0.020034f
C325 VDD1.n120 VSUBS 0.010766f
C326 VDD1.n121 VSUBS 0.011399f
C327 VDD1.n122 VSUBS 0.025446f
C328 VDD1.n123 VSUBS 0.025446f
C329 VDD1.n124 VSUBS 0.011399f
C330 VDD1.n125 VSUBS 0.010766f
C331 VDD1.n126 VSUBS 0.020034f
C332 VDD1.n127 VSUBS 0.020034f
C333 VDD1.n128 VSUBS 0.010766f
C334 VDD1.n129 VSUBS 0.011399f
C335 VDD1.n130 VSUBS 0.025446f
C336 VDD1.n131 VSUBS 0.025446f
C337 VDD1.n132 VSUBS 0.011399f
C338 VDD1.n133 VSUBS 0.010766f
C339 VDD1.n134 VSUBS 0.020034f
C340 VDD1.n135 VSUBS 0.020034f
C341 VDD1.n136 VSUBS 0.010766f
C342 VDD1.n137 VSUBS 0.011399f
C343 VDD1.n138 VSUBS 0.025446f
C344 VDD1.n139 VSUBS 0.025446f
C345 VDD1.n140 VSUBS 0.011399f
C346 VDD1.n141 VSUBS 0.010766f
C347 VDD1.n142 VSUBS 0.020034f
C348 VDD1.n143 VSUBS 0.020034f
C349 VDD1.n144 VSUBS 0.010766f
C350 VDD1.n145 VSUBS 0.011399f
C351 VDD1.n146 VSUBS 0.025446f
C352 VDD1.n147 VSUBS 0.025446f
C353 VDD1.n148 VSUBS 0.011399f
C354 VDD1.n149 VSUBS 0.010766f
C355 VDD1.n150 VSUBS 0.020034f
C356 VDD1.n151 VSUBS 0.020034f
C357 VDD1.n152 VSUBS 0.010766f
C358 VDD1.n153 VSUBS 0.010766f
C359 VDD1.n154 VSUBS 0.011399f
C360 VDD1.n155 VSUBS 0.025446f
C361 VDD1.n156 VSUBS 0.025446f
C362 VDD1.n157 VSUBS 0.025446f
C363 VDD1.n158 VSUBS 0.011082f
C364 VDD1.n159 VSUBS 0.010766f
C365 VDD1.n160 VSUBS 0.020034f
C366 VDD1.n161 VSUBS 0.020034f
C367 VDD1.n162 VSUBS 0.010766f
C368 VDD1.n163 VSUBS 0.011399f
C369 VDD1.n164 VSUBS 0.025446f
C370 VDD1.n165 VSUBS 0.058134f
C371 VDD1.n166 VSUBS 0.011399f
C372 VDD1.n167 VSUBS 0.010766f
C373 VDD1.n168 VSUBS 0.047676f
C374 VDD1.n169 VSUBS 0.67641f
C375 VTAIL.n0 VSUBS 0.029726f
C376 VTAIL.n1 VSUBS 0.028366f
C377 VTAIL.n2 VSUBS 0.015243f
C378 VTAIL.n3 VSUBS 0.036028f
C379 VTAIL.n4 VSUBS 0.015691f
C380 VTAIL.n5 VSUBS 0.028366f
C381 VTAIL.n6 VSUBS 0.016139f
C382 VTAIL.n7 VSUBS 0.036028f
C383 VTAIL.n8 VSUBS 0.016139f
C384 VTAIL.n9 VSUBS 0.028366f
C385 VTAIL.n10 VSUBS 0.015243f
C386 VTAIL.n11 VSUBS 0.036028f
C387 VTAIL.n12 VSUBS 0.016139f
C388 VTAIL.n13 VSUBS 0.028366f
C389 VTAIL.n14 VSUBS 0.015243f
C390 VTAIL.n15 VSUBS 0.036028f
C391 VTAIL.n16 VSUBS 0.016139f
C392 VTAIL.n17 VSUBS 0.028366f
C393 VTAIL.n18 VSUBS 0.015243f
C394 VTAIL.n19 VSUBS 0.036028f
C395 VTAIL.n20 VSUBS 0.016139f
C396 VTAIL.n21 VSUBS 0.028366f
C397 VTAIL.n22 VSUBS 0.015243f
C398 VTAIL.n23 VSUBS 0.036028f
C399 VTAIL.n24 VSUBS 0.016139f
C400 VTAIL.n25 VSUBS 1.864f
C401 VTAIL.n26 VSUBS 0.015243f
C402 VTAIL.t2 VSUBS 0.077157f
C403 VTAIL.n27 VSUBS 0.203384f
C404 VTAIL.n28 VSUBS 0.022919f
C405 VTAIL.n29 VSUBS 0.027021f
C406 VTAIL.n30 VSUBS 0.036028f
C407 VTAIL.n31 VSUBS 0.016139f
C408 VTAIL.n32 VSUBS 0.015243f
C409 VTAIL.n33 VSUBS 0.028366f
C410 VTAIL.n34 VSUBS 0.028366f
C411 VTAIL.n35 VSUBS 0.015243f
C412 VTAIL.n36 VSUBS 0.016139f
C413 VTAIL.n37 VSUBS 0.036028f
C414 VTAIL.n38 VSUBS 0.036028f
C415 VTAIL.n39 VSUBS 0.016139f
C416 VTAIL.n40 VSUBS 0.015243f
C417 VTAIL.n41 VSUBS 0.028366f
C418 VTAIL.n42 VSUBS 0.028366f
C419 VTAIL.n43 VSUBS 0.015243f
C420 VTAIL.n44 VSUBS 0.016139f
C421 VTAIL.n45 VSUBS 0.036028f
C422 VTAIL.n46 VSUBS 0.036028f
C423 VTAIL.n47 VSUBS 0.016139f
C424 VTAIL.n48 VSUBS 0.015243f
C425 VTAIL.n49 VSUBS 0.028366f
C426 VTAIL.n50 VSUBS 0.028366f
C427 VTAIL.n51 VSUBS 0.015243f
C428 VTAIL.n52 VSUBS 0.016139f
C429 VTAIL.n53 VSUBS 0.036028f
C430 VTAIL.n54 VSUBS 0.036028f
C431 VTAIL.n55 VSUBS 0.016139f
C432 VTAIL.n56 VSUBS 0.015243f
C433 VTAIL.n57 VSUBS 0.028366f
C434 VTAIL.n58 VSUBS 0.028366f
C435 VTAIL.n59 VSUBS 0.015243f
C436 VTAIL.n60 VSUBS 0.016139f
C437 VTAIL.n61 VSUBS 0.036028f
C438 VTAIL.n62 VSUBS 0.036028f
C439 VTAIL.n63 VSUBS 0.016139f
C440 VTAIL.n64 VSUBS 0.015243f
C441 VTAIL.n65 VSUBS 0.028366f
C442 VTAIL.n66 VSUBS 0.028366f
C443 VTAIL.n67 VSUBS 0.015243f
C444 VTAIL.n68 VSUBS 0.015243f
C445 VTAIL.n69 VSUBS 0.016139f
C446 VTAIL.n70 VSUBS 0.036028f
C447 VTAIL.n71 VSUBS 0.036028f
C448 VTAIL.n72 VSUBS 0.036028f
C449 VTAIL.n73 VSUBS 0.015691f
C450 VTAIL.n74 VSUBS 0.015243f
C451 VTAIL.n75 VSUBS 0.028366f
C452 VTAIL.n76 VSUBS 0.028366f
C453 VTAIL.n77 VSUBS 0.015243f
C454 VTAIL.n78 VSUBS 0.016139f
C455 VTAIL.n79 VSUBS 0.036028f
C456 VTAIL.n80 VSUBS 0.08231f
C457 VTAIL.n81 VSUBS 0.016139f
C458 VTAIL.n82 VSUBS 0.015243f
C459 VTAIL.n83 VSUBS 0.067503f
C460 VTAIL.n84 VSUBS 0.041234f
C461 VTAIL.n85 VSUBS 2.06136f
C462 VTAIL.n86 VSUBS 0.029726f
C463 VTAIL.n87 VSUBS 0.028366f
C464 VTAIL.n88 VSUBS 0.015243f
C465 VTAIL.n89 VSUBS 0.036028f
C466 VTAIL.n90 VSUBS 0.015691f
C467 VTAIL.n91 VSUBS 0.028366f
C468 VTAIL.n92 VSUBS 0.015691f
C469 VTAIL.n93 VSUBS 0.015243f
C470 VTAIL.n94 VSUBS 0.036028f
C471 VTAIL.n95 VSUBS 0.036028f
C472 VTAIL.n96 VSUBS 0.016139f
C473 VTAIL.n97 VSUBS 0.028366f
C474 VTAIL.n98 VSUBS 0.015243f
C475 VTAIL.n99 VSUBS 0.036028f
C476 VTAIL.n100 VSUBS 0.016139f
C477 VTAIL.n101 VSUBS 0.028366f
C478 VTAIL.n102 VSUBS 0.015243f
C479 VTAIL.n103 VSUBS 0.036028f
C480 VTAIL.n104 VSUBS 0.016139f
C481 VTAIL.n105 VSUBS 0.028366f
C482 VTAIL.n106 VSUBS 0.015243f
C483 VTAIL.n107 VSUBS 0.036028f
C484 VTAIL.n108 VSUBS 0.016139f
C485 VTAIL.n109 VSUBS 0.028366f
C486 VTAIL.n110 VSUBS 0.015243f
C487 VTAIL.n111 VSUBS 0.036028f
C488 VTAIL.n112 VSUBS 0.016139f
C489 VTAIL.n113 VSUBS 1.864f
C490 VTAIL.n114 VSUBS 0.015243f
C491 VTAIL.t1 VSUBS 0.077157f
C492 VTAIL.n115 VSUBS 0.203384f
C493 VTAIL.n116 VSUBS 0.022919f
C494 VTAIL.n117 VSUBS 0.027021f
C495 VTAIL.n118 VSUBS 0.036028f
C496 VTAIL.n119 VSUBS 0.016139f
C497 VTAIL.n120 VSUBS 0.015243f
C498 VTAIL.n121 VSUBS 0.028366f
C499 VTAIL.n122 VSUBS 0.028366f
C500 VTAIL.n123 VSUBS 0.015243f
C501 VTAIL.n124 VSUBS 0.016139f
C502 VTAIL.n125 VSUBS 0.036028f
C503 VTAIL.n126 VSUBS 0.036028f
C504 VTAIL.n127 VSUBS 0.016139f
C505 VTAIL.n128 VSUBS 0.015243f
C506 VTAIL.n129 VSUBS 0.028366f
C507 VTAIL.n130 VSUBS 0.028366f
C508 VTAIL.n131 VSUBS 0.015243f
C509 VTAIL.n132 VSUBS 0.016139f
C510 VTAIL.n133 VSUBS 0.036028f
C511 VTAIL.n134 VSUBS 0.036028f
C512 VTAIL.n135 VSUBS 0.016139f
C513 VTAIL.n136 VSUBS 0.015243f
C514 VTAIL.n137 VSUBS 0.028366f
C515 VTAIL.n138 VSUBS 0.028366f
C516 VTAIL.n139 VSUBS 0.015243f
C517 VTAIL.n140 VSUBS 0.016139f
C518 VTAIL.n141 VSUBS 0.036028f
C519 VTAIL.n142 VSUBS 0.036028f
C520 VTAIL.n143 VSUBS 0.016139f
C521 VTAIL.n144 VSUBS 0.015243f
C522 VTAIL.n145 VSUBS 0.028366f
C523 VTAIL.n146 VSUBS 0.028366f
C524 VTAIL.n147 VSUBS 0.015243f
C525 VTAIL.n148 VSUBS 0.016139f
C526 VTAIL.n149 VSUBS 0.036028f
C527 VTAIL.n150 VSUBS 0.036028f
C528 VTAIL.n151 VSUBS 0.016139f
C529 VTAIL.n152 VSUBS 0.015243f
C530 VTAIL.n153 VSUBS 0.028366f
C531 VTAIL.n154 VSUBS 0.028366f
C532 VTAIL.n155 VSUBS 0.015243f
C533 VTAIL.n156 VSUBS 0.016139f
C534 VTAIL.n157 VSUBS 0.036028f
C535 VTAIL.n158 VSUBS 0.036028f
C536 VTAIL.n159 VSUBS 0.016139f
C537 VTAIL.n160 VSUBS 0.015243f
C538 VTAIL.n161 VSUBS 0.028366f
C539 VTAIL.n162 VSUBS 0.028366f
C540 VTAIL.n163 VSUBS 0.015243f
C541 VTAIL.n164 VSUBS 0.016139f
C542 VTAIL.n165 VSUBS 0.036028f
C543 VTAIL.n166 VSUBS 0.08231f
C544 VTAIL.n167 VSUBS 0.016139f
C545 VTAIL.n168 VSUBS 0.015243f
C546 VTAIL.n169 VSUBS 0.067503f
C547 VTAIL.n170 VSUBS 0.041234f
C548 VTAIL.n171 VSUBS 2.09918f
C549 VTAIL.n172 VSUBS 0.029726f
C550 VTAIL.n173 VSUBS 0.028366f
C551 VTAIL.n174 VSUBS 0.015243f
C552 VTAIL.n175 VSUBS 0.036028f
C553 VTAIL.n176 VSUBS 0.015691f
C554 VTAIL.n177 VSUBS 0.028366f
C555 VTAIL.n178 VSUBS 0.015691f
C556 VTAIL.n179 VSUBS 0.015243f
C557 VTAIL.n180 VSUBS 0.036028f
C558 VTAIL.n181 VSUBS 0.036028f
C559 VTAIL.n182 VSUBS 0.016139f
C560 VTAIL.n183 VSUBS 0.028366f
C561 VTAIL.n184 VSUBS 0.015243f
C562 VTAIL.n185 VSUBS 0.036028f
C563 VTAIL.n186 VSUBS 0.016139f
C564 VTAIL.n187 VSUBS 0.028366f
C565 VTAIL.n188 VSUBS 0.015243f
C566 VTAIL.n189 VSUBS 0.036028f
C567 VTAIL.n190 VSUBS 0.016139f
C568 VTAIL.n191 VSUBS 0.028366f
C569 VTAIL.n192 VSUBS 0.015243f
C570 VTAIL.n193 VSUBS 0.036028f
C571 VTAIL.n194 VSUBS 0.016139f
C572 VTAIL.n195 VSUBS 0.028366f
C573 VTAIL.n196 VSUBS 0.015243f
C574 VTAIL.n197 VSUBS 0.036028f
C575 VTAIL.n198 VSUBS 0.016139f
C576 VTAIL.n199 VSUBS 1.864f
C577 VTAIL.n200 VSUBS 0.015243f
C578 VTAIL.t3 VSUBS 0.077157f
C579 VTAIL.n201 VSUBS 0.203384f
C580 VTAIL.n202 VSUBS 0.022919f
C581 VTAIL.n203 VSUBS 0.027021f
C582 VTAIL.n204 VSUBS 0.036028f
C583 VTAIL.n205 VSUBS 0.016139f
C584 VTAIL.n206 VSUBS 0.015243f
C585 VTAIL.n207 VSUBS 0.028366f
C586 VTAIL.n208 VSUBS 0.028366f
C587 VTAIL.n209 VSUBS 0.015243f
C588 VTAIL.n210 VSUBS 0.016139f
C589 VTAIL.n211 VSUBS 0.036028f
C590 VTAIL.n212 VSUBS 0.036028f
C591 VTAIL.n213 VSUBS 0.016139f
C592 VTAIL.n214 VSUBS 0.015243f
C593 VTAIL.n215 VSUBS 0.028366f
C594 VTAIL.n216 VSUBS 0.028366f
C595 VTAIL.n217 VSUBS 0.015243f
C596 VTAIL.n218 VSUBS 0.016139f
C597 VTAIL.n219 VSUBS 0.036028f
C598 VTAIL.n220 VSUBS 0.036028f
C599 VTAIL.n221 VSUBS 0.016139f
C600 VTAIL.n222 VSUBS 0.015243f
C601 VTAIL.n223 VSUBS 0.028366f
C602 VTAIL.n224 VSUBS 0.028366f
C603 VTAIL.n225 VSUBS 0.015243f
C604 VTAIL.n226 VSUBS 0.016139f
C605 VTAIL.n227 VSUBS 0.036028f
C606 VTAIL.n228 VSUBS 0.036028f
C607 VTAIL.n229 VSUBS 0.016139f
C608 VTAIL.n230 VSUBS 0.015243f
C609 VTAIL.n231 VSUBS 0.028366f
C610 VTAIL.n232 VSUBS 0.028366f
C611 VTAIL.n233 VSUBS 0.015243f
C612 VTAIL.n234 VSUBS 0.016139f
C613 VTAIL.n235 VSUBS 0.036028f
C614 VTAIL.n236 VSUBS 0.036028f
C615 VTAIL.n237 VSUBS 0.016139f
C616 VTAIL.n238 VSUBS 0.015243f
C617 VTAIL.n239 VSUBS 0.028366f
C618 VTAIL.n240 VSUBS 0.028366f
C619 VTAIL.n241 VSUBS 0.015243f
C620 VTAIL.n242 VSUBS 0.016139f
C621 VTAIL.n243 VSUBS 0.036028f
C622 VTAIL.n244 VSUBS 0.036028f
C623 VTAIL.n245 VSUBS 0.016139f
C624 VTAIL.n246 VSUBS 0.015243f
C625 VTAIL.n247 VSUBS 0.028366f
C626 VTAIL.n248 VSUBS 0.028366f
C627 VTAIL.n249 VSUBS 0.015243f
C628 VTAIL.n250 VSUBS 0.016139f
C629 VTAIL.n251 VSUBS 0.036028f
C630 VTAIL.n252 VSUBS 0.08231f
C631 VTAIL.n253 VSUBS 0.016139f
C632 VTAIL.n254 VSUBS 0.015243f
C633 VTAIL.n255 VSUBS 0.067503f
C634 VTAIL.n256 VSUBS 0.041234f
C635 VTAIL.n257 VSUBS 1.92662f
C636 VTAIL.n258 VSUBS 0.029726f
C637 VTAIL.n259 VSUBS 0.028366f
C638 VTAIL.n260 VSUBS 0.015243f
C639 VTAIL.n261 VSUBS 0.036028f
C640 VTAIL.n262 VSUBS 0.015691f
C641 VTAIL.n263 VSUBS 0.028366f
C642 VTAIL.n264 VSUBS 0.016139f
C643 VTAIL.n265 VSUBS 0.036028f
C644 VTAIL.n266 VSUBS 0.016139f
C645 VTAIL.n267 VSUBS 0.028366f
C646 VTAIL.n268 VSUBS 0.015243f
C647 VTAIL.n269 VSUBS 0.036028f
C648 VTAIL.n270 VSUBS 0.016139f
C649 VTAIL.n271 VSUBS 0.028366f
C650 VTAIL.n272 VSUBS 0.015243f
C651 VTAIL.n273 VSUBS 0.036028f
C652 VTAIL.n274 VSUBS 0.016139f
C653 VTAIL.n275 VSUBS 0.028366f
C654 VTAIL.n276 VSUBS 0.015243f
C655 VTAIL.n277 VSUBS 0.036028f
C656 VTAIL.n278 VSUBS 0.016139f
C657 VTAIL.n279 VSUBS 0.028366f
C658 VTAIL.n280 VSUBS 0.015243f
C659 VTAIL.n281 VSUBS 0.036028f
C660 VTAIL.n282 VSUBS 0.016139f
C661 VTAIL.n283 VSUBS 1.864f
C662 VTAIL.n284 VSUBS 0.015243f
C663 VTAIL.t0 VSUBS 0.077157f
C664 VTAIL.n285 VSUBS 0.203384f
C665 VTAIL.n286 VSUBS 0.022919f
C666 VTAIL.n287 VSUBS 0.027021f
C667 VTAIL.n288 VSUBS 0.036028f
C668 VTAIL.n289 VSUBS 0.016139f
C669 VTAIL.n290 VSUBS 0.015243f
C670 VTAIL.n291 VSUBS 0.028366f
C671 VTAIL.n292 VSUBS 0.028366f
C672 VTAIL.n293 VSUBS 0.015243f
C673 VTAIL.n294 VSUBS 0.016139f
C674 VTAIL.n295 VSUBS 0.036028f
C675 VTAIL.n296 VSUBS 0.036028f
C676 VTAIL.n297 VSUBS 0.016139f
C677 VTAIL.n298 VSUBS 0.015243f
C678 VTAIL.n299 VSUBS 0.028366f
C679 VTAIL.n300 VSUBS 0.028366f
C680 VTAIL.n301 VSUBS 0.015243f
C681 VTAIL.n302 VSUBS 0.016139f
C682 VTAIL.n303 VSUBS 0.036028f
C683 VTAIL.n304 VSUBS 0.036028f
C684 VTAIL.n305 VSUBS 0.016139f
C685 VTAIL.n306 VSUBS 0.015243f
C686 VTAIL.n307 VSUBS 0.028366f
C687 VTAIL.n308 VSUBS 0.028366f
C688 VTAIL.n309 VSUBS 0.015243f
C689 VTAIL.n310 VSUBS 0.016139f
C690 VTAIL.n311 VSUBS 0.036028f
C691 VTAIL.n312 VSUBS 0.036028f
C692 VTAIL.n313 VSUBS 0.016139f
C693 VTAIL.n314 VSUBS 0.015243f
C694 VTAIL.n315 VSUBS 0.028366f
C695 VTAIL.n316 VSUBS 0.028366f
C696 VTAIL.n317 VSUBS 0.015243f
C697 VTAIL.n318 VSUBS 0.016139f
C698 VTAIL.n319 VSUBS 0.036028f
C699 VTAIL.n320 VSUBS 0.036028f
C700 VTAIL.n321 VSUBS 0.016139f
C701 VTAIL.n322 VSUBS 0.015243f
C702 VTAIL.n323 VSUBS 0.028366f
C703 VTAIL.n324 VSUBS 0.028366f
C704 VTAIL.n325 VSUBS 0.015243f
C705 VTAIL.n326 VSUBS 0.015243f
C706 VTAIL.n327 VSUBS 0.016139f
C707 VTAIL.n328 VSUBS 0.036028f
C708 VTAIL.n329 VSUBS 0.036028f
C709 VTAIL.n330 VSUBS 0.036028f
C710 VTAIL.n331 VSUBS 0.015691f
C711 VTAIL.n332 VSUBS 0.015243f
C712 VTAIL.n333 VSUBS 0.028366f
C713 VTAIL.n334 VSUBS 0.028366f
C714 VTAIL.n335 VSUBS 0.015243f
C715 VTAIL.n336 VSUBS 0.016139f
C716 VTAIL.n337 VSUBS 0.036028f
C717 VTAIL.n338 VSUBS 0.08231f
C718 VTAIL.n339 VSUBS 0.016139f
C719 VTAIL.n340 VSUBS 0.015243f
C720 VTAIL.n341 VSUBS 0.067503f
C721 VTAIL.n342 VSUBS 0.041234f
C722 VTAIL.n343 VSUBS 1.83522f
C723 VP.t0 VSUBS 4.43943f
C724 VP.t1 VSUBS 3.93286f
C725 VP.n0 VSUBS 6.25597f
C726 B.n0 VSUBS 0.003852f
C727 B.n1 VSUBS 0.003852f
C728 B.n2 VSUBS 0.006092f
C729 B.n3 VSUBS 0.006092f
C730 B.n4 VSUBS 0.006092f
C731 B.n5 VSUBS 0.006092f
C732 B.n6 VSUBS 0.006092f
C733 B.n7 VSUBS 0.006092f
C734 B.n8 VSUBS 0.006092f
C735 B.n9 VSUBS 0.006092f
C736 B.n10 VSUBS 0.006092f
C737 B.n11 VSUBS 0.006092f
C738 B.n12 VSUBS 0.013587f
C739 B.n13 VSUBS 0.006092f
C740 B.n14 VSUBS 0.006092f
C741 B.n15 VSUBS 0.006092f
C742 B.n16 VSUBS 0.006092f
C743 B.n17 VSUBS 0.006092f
C744 B.n18 VSUBS 0.006092f
C745 B.n19 VSUBS 0.006092f
C746 B.n20 VSUBS 0.006092f
C747 B.n21 VSUBS 0.006092f
C748 B.n22 VSUBS 0.006092f
C749 B.n23 VSUBS 0.006092f
C750 B.n24 VSUBS 0.006092f
C751 B.n25 VSUBS 0.006092f
C752 B.n26 VSUBS 0.006092f
C753 B.n27 VSUBS 0.006092f
C754 B.n28 VSUBS 0.006092f
C755 B.n29 VSUBS 0.006092f
C756 B.n30 VSUBS 0.006092f
C757 B.n31 VSUBS 0.006092f
C758 B.n32 VSUBS 0.006092f
C759 B.n33 VSUBS 0.006092f
C760 B.n34 VSUBS 0.006092f
C761 B.n35 VSUBS 0.006092f
C762 B.n36 VSUBS 0.006092f
C763 B.n37 VSUBS 0.006092f
C764 B.n38 VSUBS 0.004211f
C765 B.n39 VSUBS 0.006092f
C766 B.t11 VSUBS 0.251639f
C767 B.t10 VSUBS 0.27353f
C768 B.t9 VSUBS 1.09029f
C769 B.n40 VSUBS 0.408069f
C770 B.n41 VSUBS 0.255802f
C771 B.n42 VSUBS 0.014114f
C772 B.n43 VSUBS 0.006092f
C773 B.n44 VSUBS 0.006092f
C774 B.n45 VSUBS 0.006092f
C775 B.n46 VSUBS 0.006092f
C776 B.t5 VSUBS 0.251642f
C777 B.t4 VSUBS 0.273533f
C778 B.t3 VSUBS 1.09029f
C779 B.n47 VSUBS 0.408066f
C780 B.n48 VSUBS 0.255799f
C781 B.n49 VSUBS 0.006092f
C782 B.n50 VSUBS 0.006092f
C783 B.n51 VSUBS 0.006092f
C784 B.n52 VSUBS 0.006092f
C785 B.n53 VSUBS 0.006092f
C786 B.n54 VSUBS 0.006092f
C787 B.n55 VSUBS 0.006092f
C788 B.n56 VSUBS 0.006092f
C789 B.n57 VSUBS 0.006092f
C790 B.n58 VSUBS 0.006092f
C791 B.n59 VSUBS 0.006092f
C792 B.n60 VSUBS 0.006092f
C793 B.n61 VSUBS 0.006092f
C794 B.n62 VSUBS 0.006092f
C795 B.n63 VSUBS 0.006092f
C796 B.n64 VSUBS 0.006092f
C797 B.n65 VSUBS 0.006092f
C798 B.n66 VSUBS 0.006092f
C799 B.n67 VSUBS 0.006092f
C800 B.n68 VSUBS 0.006092f
C801 B.n69 VSUBS 0.006092f
C802 B.n70 VSUBS 0.006092f
C803 B.n71 VSUBS 0.006092f
C804 B.n72 VSUBS 0.006092f
C805 B.n73 VSUBS 0.006092f
C806 B.n74 VSUBS 0.013587f
C807 B.n75 VSUBS 0.006092f
C808 B.n76 VSUBS 0.006092f
C809 B.n77 VSUBS 0.006092f
C810 B.n78 VSUBS 0.006092f
C811 B.n79 VSUBS 0.006092f
C812 B.n80 VSUBS 0.006092f
C813 B.n81 VSUBS 0.006092f
C814 B.n82 VSUBS 0.006092f
C815 B.n83 VSUBS 0.006092f
C816 B.n84 VSUBS 0.006092f
C817 B.n85 VSUBS 0.006092f
C818 B.n86 VSUBS 0.006092f
C819 B.n87 VSUBS 0.006092f
C820 B.n88 VSUBS 0.006092f
C821 B.n89 VSUBS 0.006092f
C822 B.n90 VSUBS 0.006092f
C823 B.n91 VSUBS 0.006092f
C824 B.n92 VSUBS 0.006092f
C825 B.n93 VSUBS 0.006092f
C826 B.n94 VSUBS 0.006092f
C827 B.n95 VSUBS 0.013587f
C828 B.n96 VSUBS 0.006092f
C829 B.n97 VSUBS 0.006092f
C830 B.n98 VSUBS 0.006092f
C831 B.n99 VSUBS 0.006092f
C832 B.n100 VSUBS 0.006092f
C833 B.n101 VSUBS 0.006092f
C834 B.n102 VSUBS 0.006092f
C835 B.n103 VSUBS 0.006092f
C836 B.n104 VSUBS 0.006092f
C837 B.n105 VSUBS 0.006092f
C838 B.n106 VSUBS 0.006092f
C839 B.n107 VSUBS 0.006092f
C840 B.n108 VSUBS 0.006092f
C841 B.n109 VSUBS 0.006092f
C842 B.n110 VSUBS 0.006092f
C843 B.n111 VSUBS 0.006092f
C844 B.n112 VSUBS 0.006092f
C845 B.n113 VSUBS 0.006092f
C846 B.n114 VSUBS 0.006092f
C847 B.n115 VSUBS 0.006092f
C848 B.n116 VSUBS 0.006092f
C849 B.n117 VSUBS 0.006092f
C850 B.n118 VSUBS 0.006092f
C851 B.n119 VSUBS 0.006092f
C852 B.n120 VSUBS 0.006092f
C853 B.n121 VSUBS 0.004211f
C854 B.n122 VSUBS 0.006092f
C855 B.n123 VSUBS 0.006092f
C856 B.n124 VSUBS 0.006092f
C857 B.n125 VSUBS 0.006092f
C858 B.n126 VSUBS 0.006092f
C859 B.t1 VSUBS 0.251639f
C860 B.t2 VSUBS 0.27353f
C861 B.t0 VSUBS 1.09029f
C862 B.n127 VSUBS 0.408069f
C863 B.n128 VSUBS 0.255802f
C864 B.n129 VSUBS 0.006092f
C865 B.n130 VSUBS 0.006092f
C866 B.n131 VSUBS 0.006092f
C867 B.n132 VSUBS 0.006092f
C868 B.n133 VSUBS 0.006092f
C869 B.n134 VSUBS 0.006092f
C870 B.n135 VSUBS 0.006092f
C871 B.n136 VSUBS 0.006092f
C872 B.n137 VSUBS 0.006092f
C873 B.n138 VSUBS 0.006092f
C874 B.n139 VSUBS 0.006092f
C875 B.n140 VSUBS 0.006092f
C876 B.n141 VSUBS 0.006092f
C877 B.n142 VSUBS 0.006092f
C878 B.n143 VSUBS 0.006092f
C879 B.n144 VSUBS 0.006092f
C880 B.n145 VSUBS 0.006092f
C881 B.n146 VSUBS 0.006092f
C882 B.n147 VSUBS 0.006092f
C883 B.n148 VSUBS 0.006092f
C884 B.n149 VSUBS 0.006092f
C885 B.n150 VSUBS 0.006092f
C886 B.n151 VSUBS 0.006092f
C887 B.n152 VSUBS 0.006092f
C888 B.n153 VSUBS 0.006092f
C889 B.n154 VSUBS 0.013587f
C890 B.n155 VSUBS 0.006092f
C891 B.n156 VSUBS 0.006092f
C892 B.n157 VSUBS 0.006092f
C893 B.n158 VSUBS 0.006092f
C894 B.n159 VSUBS 0.006092f
C895 B.n160 VSUBS 0.006092f
C896 B.n161 VSUBS 0.006092f
C897 B.n162 VSUBS 0.006092f
C898 B.n163 VSUBS 0.006092f
C899 B.n164 VSUBS 0.006092f
C900 B.n165 VSUBS 0.006092f
C901 B.n166 VSUBS 0.006092f
C902 B.n167 VSUBS 0.006092f
C903 B.n168 VSUBS 0.006092f
C904 B.n169 VSUBS 0.006092f
C905 B.n170 VSUBS 0.006092f
C906 B.n171 VSUBS 0.006092f
C907 B.n172 VSUBS 0.006092f
C908 B.n173 VSUBS 0.006092f
C909 B.n174 VSUBS 0.006092f
C910 B.n175 VSUBS 0.006092f
C911 B.n176 VSUBS 0.006092f
C912 B.n177 VSUBS 0.006092f
C913 B.n178 VSUBS 0.006092f
C914 B.n179 VSUBS 0.006092f
C915 B.n180 VSUBS 0.006092f
C916 B.n181 VSUBS 0.006092f
C917 B.n182 VSUBS 0.006092f
C918 B.n183 VSUBS 0.006092f
C919 B.n184 VSUBS 0.006092f
C920 B.n185 VSUBS 0.006092f
C921 B.n186 VSUBS 0.006092f
C922 B.n187 VSUBS 0.006092f
C923 B.n188 VSUBS 0.006092f
C924 B.n189 VSUBS 0.006092f
C925 B.n190 VSUBS 0.006092f
C926 B.n191 VSUBS 0.006092f
C927 B.n192 VSUBS 0.006092f
C928 B.n193 VSUBS 0.013587f
C929 B.n194 VSUBS 0.014365f
C930 B.n195 VSUBS 0.014365f
C931 B.n196 VSUBS 0.006092f
C932 B.n197 VSUBS 0.006092f
C933 B.n198 VSUBS 0.006092f
C934 B.n199 VSUBS 0.006092f
C935 B.n200 VSUBS 0.006092f
C936 B.n201 VSUBS 0.006092f
C937 B.n202 VSUBS 0.006092f
C938 B.n203 VSUBS 0.006092f
C939 B.n204 VSUBS 0.006092f
C940 B.n205 VSUBS 0.006092f
C941 B.n206 VSUBS 0.006092f
C942 B.n207 VSUBS 0.006092f
C943 B.n208 VSUBS 0.006092f
C944 B.n209 VSUBS 0.006092f
C945 B.n210 VSUBS 0.006092f
C946 B.n211 VSUBS 0.006092f
C947 B.n212 VSUBS 0.006092f
C948 B.n213 VSUBS 0.006092f
C949 B.n214 VSUBS 0.006092f
C950 B.n215 VSUBS 0.006092f
C951 B.n216 VSUBS 0.006092f
C952 B.n217 VSUBS 0.006092f
C953 B.n218 VSUBS 0.006092f
C954 B.n219 VSUBS 0.006092f
C955 B.n220 VSUBS 0.006092f
C956 B.n221 VSUBS 0.006092f
C957 B.n222 VSUBS 0.006092f
C958 B.n223 VSUBS 0.006092f
C959 B.n224 VSUBS 0.006092f
C960 B.n225 VSUBS 0.006092f
C961 B.n226 VSUBS 0.006092f
C962 B.n227 VSUBS 0.006092f
C963 B.n228 VSUBS 0.006092f
C964 B.n229 VSUBS 0.006092f
C965 B.n230 VSUBS 0.006092f
C966 B.n231 VSUBS 0.006092f
C967 B.n232 VSUBS 0.006092f
C968 B.n233 VSUBS 0.006092f
C969 B.n234 VSUBS 0.006092f
C970 B.n235 VSUBS 0.006092f
C971 B.n236 VSUBS 0.006092f
C972 B.n237 VSUBS 0.006092f
C973 B.n238 VSUBS 0.006092f
C974 B.n239 VSUBS 0.006092f
C975 B.n240 VSUBS 0.006092f
C976 B.n241 VSUBS 0.006092f
C977 B.n242 VSUBS 0.006092f
C978 B.n243 VSUBS 0.006092f
C979 B.n244 VSUBS 0.006092f
C980 B.n245 VSUBS 0.006092f
C981 B.n246 VSUBS 0.006092f
C982 B.n247 VSUBS 0.006092f
C983 B.n248 VSUBS 0.006092f
C984 B.n249 VSUBS 0.006092f
C985 B.n250 VSUBS 0.006092f
C986 B.n251 VSUBS 0.006092f
C987 B.n252 VSUBS 0.006092f
C988 B.n253 VSUBS 0.006092f
C989 B.n254 VSUBS 0.006092f
C990 B.n255 VSUBS 0.006092f
C991 B.n256 VSUBS 0.006092f
C992 B.n257 VSUBS 0.006092f
C993 B.n258 VSUBS 0.006092f
C994 B.n259 VSUBS 0.006092f
C995 B.n260 VSUBS 0.006092f
C996 B.n261 VSUBS 0.006092f
C997 B.n262 VSUBS 0.006092f
C998 B.n263 VSUBS 0.006092f
C999 B.n264 VSUBS 0.006092f
C1000 B.n265 VSUBS 0.006092f
C1001 B.n266 VSUBS 0.006092f
C1002 B.n267 VSUBS 0.006092f
C1003 B.n268 VSUBS 0.006092f
C1004 B.n269 VSUBS 0.006092f
C1005 B.n270 VSUBS 0.006092f
C1006 B.n271 VSUBS 0.004211f
C1007 B.n272 VSUBS 0.014114f
C1008 B.n273 VSUBS 0.004927f
C1009 B.n274 VSUBS 0.006092f
C1010 B.n275 VSUBS 0.006092f
C1011 B.n276 VSUBS 0.006092f
C1012 B.n277 VSUBS 0.006092f
C1013 B.n278 VSUBS 0.006092f
C1014 B.n279 VSUBS 0.006092f
C1015 B.n280 VSUBS 0.006092f
C1016 B.n281 VSUBS 0.006092f
C1017 B.n282 VSUBS 0.006092f
C1018 B.n283 VSUBS 0.006092f
C1019 B.n284 VSUBS 0.006092f
C1020 B.t7 VSUBS 0.251642f
C1021 B.t8 VSUBS 0.273533f
C1022 B.t6 VSUBS 1.09029f
C1023 B.n285 VSUBS 0.408066f
C1024 B.n286 VSUBS 0.255799f
C1025 B.n287 VSUBS 0.014114f
C1026 B.n288 VSUBS 0.004927f
C1027 B.n289 VSUBS 0.006092f
C1028 B.n290 VSUBS 0.006092f
C1029 B.n291 VSUBS 0.006092f
C1030 B.n292 VSUBS 0.006092f
C1031 B.n293 VSUBS 0.006092f
C1032 B.n294 VSUBS 0.006092f
C1033 B.n295 VSUBS 0.006092f
C1034 B.n296 VSUBS 0.006092f
C1035 B.n297 VSUBS 0.006092f
C1036 B.n298 VSUBS 0.006092f
C1037 B.n299 VSUBS 0.006092f
C1038 B.n300 VSUBS 0.006092f
C1039 B.n301 VSUBS 0.006092f
C1040 B.n302 VSUBS 0.006092f
C1041 B.n303 VSUBS 0.006092f
C1042 B.n304 VSUBS 0.006092f
C1043 B.n305 VSUBS 0.006092f
C1044 B.n306 VSUBS 0.006092f
C1045 B.n307 VSUBS 0.006092f
C1046 B.n308 VSUBS 0.006092f
C1047 B.n309 VSUBS 0.006092f
C1048 B.n310 VSUBS 0.006092f
C1049 B.n311 VSUBS 0.006092f
C1050 B.n312 VSUBS 0.006092f
C1051 B.n313 VSUBS 0.006092f
C1052 B.n314 VSUBS 0.006092f
C1053 B.n315 VSUBS 0.006092f
C1054 B.n316 VSUBS 0.006092f
C1055 B.n317 VSUBS 0.006092f
C1056 B.n318 VSUBS 0.006092f
C1057 B.n319 VSUBS 0.006092f
C1058 B.n320 VSUBS 0.006092f
C1059 B.n321 VSUBS 0.006092f
C1060 B.n322 VSUBS 0.006092f
C1061 B.n323 VSUBS 0.006092f
C1062 B.n324 VSUBS 0.006092f
C1063 B.n325 VSUBS 0.006092f
C1064 B.n326 VSUBS 0.006092f
C1065 B.n327 VSUBS 0.006092f
C1066 B.n328 VSUBS 0.006092f
C1067 B.n329 VSUBS 0.006092f
C1068 B.n330 VSUBS 0.006092f
C1069 B.n331 VSUBS 0.006092f
C1070 B.n332 VSUBS 0.006092f
C1071 B.n333 VSUBS 0.006092f
C1072 B.n334 VSUBS 0.006092f
C1073 B.n335 VSUBS 0.006092f
C1074 B.n336 VSUBS 0.006092f
C1075 B.n337 VSUBS 0.006092f
C1076 B.n338 VSUBS 0.006092f
C1077 B.n339 VSUBS 0.006092f
C1078 B.n340 VSUBS 0.006092f
C1079 B.n341 VSUBS 0.006092f
C1080 B.n342 VSUBS 0.006092f
C1081 B.n343 VSUBS 0.006092f
C1082 B.n344 VSUBS 0.006092f
C1083 B.n345 VSUBS 0.006092f
C1084 B.n346 VSUBS 0.006092f
C1085 B.n347 VSUBS 0.006092f
C1086 B.n348 VSUBS 0.006092f
C1087 B.n349 VSUBS 0.006092f
C1088 B.n350 VSUBS 0.006092f
C1089 B.n351 VSUBS 0.006092f
C1090 B.n352 VSUBS 0.006092f
C1091 B.n353 VSUBS 0.006092f
C1092 B.n354 VSUBS 0.006092f
C1093 B.n355 VSUBS 0.006092f
C1094 B.n356 VSUBS 0.006092f
C1095 B.n357 VSUBS 0.006092f
C1096 B.n358 VSUBS 0.006092f
C1097 B.n359 VSUBS 0.006092f
C1098 B.n360 VSUBS 0.006092f
C1099 B.n361 VSUBS 0.006092f
C1100 B.n362 VSUBS 0.006092f
C1101 B.n363 VSUBS 0.006092f
C1102 B.n364 VSUBS 0.006092f
C1103 B.n365 VSUBS 0.006092f
C1104 B.n366 VSUBS 0.014365f
C1105 B.n367 VSUBS 0.014365f
C1106 B.n368 VSUBS 0.013587f
C1107 B.n369 VSUBS 0.006092f
C1108 B.n370 VSUBS 0.006092f
C1109 B.n371 VSUBS 0.006092f
C1110 B.n372 VSUBS 0.006092f
C1111 B.n373 VSUBS 0.006092f
C1112 B.n374 VSUBS 0.006092f
C1113 B.n375 VSUBS 0.006092f
C1114 B.n376 VSUBS 0.006092f
C1115 B.n377 VSUBS 0.006092f
C1116 B.n378 VSUBS 0.006092f
C1117 B.n379 VSUBS 0.006092f
C1118 B.n380 VSUBS 0.006092f
C1119 B.n381 VSUBS 0.006092f
C1120 B.n382 VSUBS 0.006092f
C1121 B.n383 VSUBS 0.006092f
C1122 B.n384 VSUBS 0.006092f
C1123 B.n385 VSUBS 0.006092f
C1124 B.n386 VSUBS 0.006092f
C1125 B.n387 VSUBS 0.006092f
C1126 B.n388 VSUBS 0.006092f
C1127 B.n389 VSUBS 0.006092f
C1128 B.n390 VSUBS 0.006092f
C1129 B.n391 VSUBS 0.006092f
C1130 B.n392 VSUBS 0.006092f
C1131 B.n393 VSUBS 0.006092f
C1132 B.n394 VSUBS 0.006092f
C1133 B.n395 VSUBS 0.006092f
C1134 B.n396 VSUBS 0.006092f
C1135 B.n397 VSUBS 0.006092f
C1136 B.n398 VSUBS 0.006092f
C1137 B.n399 VSUBS 0.006092f
C1138 B.n400 VSUBS 0.006092f
C1139 B.n401 VSUBS 0.006092f
C1140 B.n402 VSUBS 0.006092f
C1141 B.n403 VSUBS 0.006092f
C1142 B.n404 VSUBS 0.006092f
C1143 B.n405 VSUBS 0.006092f
C1144 B.n406 VSUBS 0.006092f
C1145 B.n407 VSUBS 0.006092f
C1146 B.n408 VSUBS 0.006092f
C1147 B.n409 VSUBS 0.006092f
C1148 B.n410 VSUBS 0.006092f
C1149 B.n411 VSUBS 0.006092f
C1150 B.n412 VSUBS 0.006092f
C1151 B.n413 VSUBS 0.006092f
C1152 B.n414 VSUBS 0.006092f
C1153 B.n415 VSUBS 0.006092f
C1154 B.n416 VSUBS 0.006092f
C1155 B.n417 VSUBS 0.006092f
C1156 B.n418 VSUBS 0.006092f
C1157 B.n419 VSUBS 0.006092f
C1158 B.n420 VSUBS 0.006092f
C1159 B.n421 VSUBS 0.006092f
C1160 B.n422 VSUBS 0.006092f
C1161 B.n423 VSUBS 0.006092f
C1162 B.n424 VSUBS 0.006092f
C1163 B.n425 VSUBS 0.006092f
C1164 B.n426 VSUBS 0.006092f
C1165 B.n427 VSUBS 0.006092f
C1166 B.n428 VSUBS 0.006092f
C1167 B.n429 VSUBS 0.006092f
C1168 B.n430 VSUBS 0.006092f
C1169 B.n431 VSUBS 0.014328f
C1170 B.n432 VSUBS 0.013623f
C1171 B.n433 VSUBS 0.014365f
C1172 B.n434 VSUBS 0.006092f
C1173 B.n435 VSUBS 0.006092f
C1174 B.n436 VSUBS 0.006092f
C1175 B.n437 VSUBS 0.006092f
C1176 B.n438 VSUBS 0.006092f
C1177 B.n439 VSUBS 0.006092f
C1178 B.n440 VSUBS 0.006092f
C1179 B.n441 VSUBS 0.006092f
C1180 B.n442 VSUBS 0.006092f
C1181 B.n443 VSUBS 0.006092f
C1182 B.n444 VSUBS 0.006092f
C1183 B.n445 VSUBS 0.006092f
C1184 B.n446 VSUBS 0.006092f
C1185 B.n447 VSUBS 0.006092f
C1186 B.n448 VSUBS 0.006092f
C1187 B.n449 VSUBS 0.006092f
C1188 B.n450 VSUBS 0.006092f
C1189 B.n451 VSUBS 0.006092f
C1190 B.n452 VSUBS 0.006092f
C1191 B.n453 VSUBS 0.006092f
C1192 B.n454 VSUBS 0.006092f
C1193 B.n455 VSUBS 0.006092f
C1194 B.n456 VSUBS 0.006092f
C1195 B.n457 VSUBS 0.006092f
C1196 B.n458 VSUBS 0.006092f
C1197 B.n459 VSUBS 0.006092f
C1198 B.n460 VSUBS 0.006092f
C1199 B.n461 VSUBS 0.006092f
C1200 B.n462 VSUBS 0.006092f
C1201 B.n463 VSUBS 0.006092f
C1202 B.n464 VSUBS 0.006092f
C1203 B.n465 VSUBS 0.006092f
C1204 B.n466 VSUBS 0.006092f
C1205 B.n467 VSUBS 0.006092f
C1206 B.n468 VSUBS 0.006092f
C1207 B.n469 VSUBS 0.006092f
C1208 B.n470 VSUBS 0.006092f
C1209 B.n471 VSUBS 0.006092f
C1210 B.n472 VSUBS 0.006092f
C1211 B.n473 VSUBS 0.006092f
C1212 B.n474 VSUBS 0.006092f
C1213 B.n475 VSUBS 0.006092f
C1214 B.n476 VSUBS 0.006092f
C1215 B.n477 VSUBS 0.006092f
C1216 B.n478 VSUBS 0.006092f
C1217 B.n479 VSUBS 0.006092f
C1218 B.n480 VSUBS 0.006092f
C1219 B.n481 VSUBS 0.006092f
C1220 B.n482 VSUBS 0.006092f
C1221 B.n483 VSUBS 0.006092f
C1222 B.n484 VSUBS 0.006092f
C1223 B.n485 VSUBS 0.006092f
C1224 B.n486 VSUBS 0.006092f
C1225 B.n487 VSUBS 0.006092f
C1226 B.n488 VSUBS 0.006092f
C1227 B.n489 VSUBS 0.006092f
C1228 B.n490 VSUBS 0.006092f
C1229 B.n491 VSUBS 0.006092f
C1230 B.n492 VSUBS 0.006092f
C1231 B.n493 VSUBS 0.006092f
C1232 B.n494 VSUBS 0.006092f
C1233 B.n495 VSUBS 0.006092f
C1234 B.n496 VSUBS 0.006092f
C1235 B.n497 VSUBS 0.006092f
C1236 B.n498 VSUBS 0.006092f
C1237 B.n499 VSUBS 0.006092f
C1238 B.n500 VSUBS 0.006092f
C1239 B.n501 VSUBS 0.006092f
C1240 B.n502 VSUBS 0.006092f
C1241 B.n503 VSUBS 0.006092f
C1242 B.n504 VSUBS 0.006092f
C1243 B.n505 VSUBS 0.006092f
C1244 B.n506 VSUBS 0.006092f
C1245 B.n507 VSUBS 0.006092f
C1246 B.n508 VSUBS 0.006092f
C1247 B.n509 VSUBS 0.004211f
C1248 B.n510 VSUBS 0.014114f
C1249 B.n511 VSUBS 0.004927f
C1250 B.n512 VSUBS 0.006092f
C1251 B.n513 VSUBS 0.006092f
C1252 B.n514 VSUBS 0.006092f
C1253 B.n515 VSUBS 0.006092f
C1254 B.n516 VSUBS 0.006092f
C1255 B.n517 VSUBS 0.006092f
C1256 B.n518 VSUBS 0.006092f
C1257 B.n519 VSUBS 0.006092f
C1258 B.n520 VSUBS 0.006092f
C1259 B.n521 VSUBS 0.006092f
C1260 B.n522 VSUBS 0.006092f
C1261 B.n523 VSUBS 0.004927f
C1262 B.n524 VSUBS 0.006092f
C1263 B.n525 VSUBS 0.006092f
C1264 B.n526 VSUBS 0.006092f
C1265 B.n527 VSUBS 0.006092f
C1266 B.n528 VSUBS 0.006092f
C1267 B.n529 VSUBS 0.006092f
C1268 B.n530 VSUBS 0.006092f
C1269 B.n531 VSUBS 0.006092f
C1270 B.n532 VSUBS 0.006092f
C1271 B.n533 VSUBS 0.006092f
C1272 B.n534 VSUBS 0.006092f
C1273 B.n535 VSUBS 0.006092f
C1274 B.n536 VSUBS 0.006092f
C1275 B.n537 VSUBS 0.006092f
C1276 B.n538 VSUBS 0.006092f
C1277 B.n539 VSUBS 0.006092f
C1278 B.n540 VSUBS 0.006092f
C1279 B.n541 VSUBS 0.006092f
C1280 B.n542 VSUBS 0.006092f
C1281 B.n543 VSUBS 0.006092f
C1282 B.n544 VSUBS 0.006092f
C1283 B.n545 VSUBS 0.006092f
C1284 B.n546 VSUBS 0.006092f
C1285 B.n547 VSUBS 0.006092f
C1286 B.n548 VSUBS 0.006092f
C1287 B.n549 VSUBS 0.006092f
C1288 B.n550 VSUBS 0.006092f
C1289 B.n551 VSUBS 0.006092f
C1290 B.n552 VSUBS 0.006092f
C1291 B.n553 VSUBS 0.006092f
C1292 B.n554 VSUBS 0.006092f
C1293 B.n555 VSUBS 0.006092f
C1294 B.n556 VSUBS 0.006092f
C1295 B.n557 VSUBS 0.006092f
C1296 B.n558 VSUBS 0.006092f
C1297 B.n559 VSUBS 0.006092f
C1298 B.n560 VSUBS 0.006092f
C1299 B.n561 VSUBS 0.006092f
C1300 B.n562 VSUBS 0.006092f
C1301 B.n563 VSUBS 0.006092f
C1302 B.n564 VSUBS 0.006092f
C1303 B.n565 VSUBS 0.006092f
C1304 B.n566 VSUBS 0.006092f
C1305 B.n567 VSUBS 0.006092f
C1306 B.n568 VSUBS 0.006092f
C1307 B.n569 VSUBS 0.006092f
C1308 B.n570 VSUBS 0.006092f
C1309 B.n571 VSUBS 0.006092f
C1310 B.n572 VSUBS 0.006092f
C1311 B.n573 VSUBS 0.006092f
C1312 B.n574 VSUBS 0.006092f
C1313 B.n575 VSUBS 0.006092f
C1314 B.n576 VSUBS 0.006092f
C1315 B.n577 VSUBS 0.006092f
C1316 B.n578 VSUBS 0.006092f
C1317 B.n579 VSUBS 0.006092f
C1318 B.n580 VSUBS 0.006092f
C1319 B.n581 VSUBS 0.006092f
C1320 B.n582 VSUBS 0.006092f
C1321 B.n583 VSUBS 0.006092f
C1322 B.n584 VSUBS 0.006092f
C1323 B.n585 VSUBS 0.006092f
C1324 B.n586 VSUBS 0.006092f
C1325 B.n587 VSUBS 0.006092f
C1326 B.n588 VSUBS 0.006092f
C1327 B.n589 VSUBS 0.006092f
C1328 B.n590 VSUBS 0.006092f
C1329 B.n591 VSUBS 0.006092f
C1330 B.n592 VSUBS 0.006092f
C1331 B.n593 VSUBS 0.006092f
C1332 B.n594 VSUBS 0.006092f
C1333 B.n595 VSUBS 0.006092f
C1334 B.n596 VSUBS 0.006092f
C1335 B.n597 VSUBS 0.006092f
C1336 B.n598 VSUBS 0.006092f
C1337 B.n599 VSUBS 0.006092f
C1338 B.n600 VSUBS 0.006092f
C1339 B.n601 VSUBS 0.014365f
C1340 B.n602 VSUBS 0.014365f
C1341 B.n603 VSUBS 0.013587f
C1342 B.n604 VSUBS 0.006092f
C1343 B.n605 VSUBS 0.006092f
C1344 B.n606 VSUBS 0.006092f
C1345 B.n607 VSUBS 0.006092f
C1346 B.n608 VSUBS 0.006092f
C1347 B.n609 VSUBS 0.006092f
C1348 B.n610 VSUBS 0.006092f
C1349 B.n611 VSUBS 0.006092f
C1350 B.n612 VSUBS 0.006092f
C1351 B.n613 VSUBS 0.006092f
C1352 B.n614 VSUBS 0.006092f
C1353 B.n615 VSUBS 0.006092f
C1354 B.n616 VSUBS 0.006092f
C1355 B.n617 VSUBS 0.006092f
C1356 B.n618 VSUBS 0.006092f
C1357 B.n619 VSUBS 0.006092f
C1358 B.n620 VSUBS 0.006092f
C1359 B.n621 VSUBS 0.006092f
C1360 B.n622 VSUBS 0.006092f
C1361 B.n623 VSUBS 0.006092f
C1362 B.n624 VSUBS 0.006092f
C1363 B.n625 VSUBS 0.006092f
C1364 B.n626 VSUBS 0.006092f
C1365 B.n627 VSUBS 0.006092f
C1366 B.n628 VSUBS 0.006092f
C1367 B.n629 VSUBS 0.006092f
C1368 B.n630 VSUBS 0.006092f
C1369 B.n631 VSUBS 0.006092f
C1370 B.n632 VSUBS 0.006092f
C1371 B.n633 VSUBS 0.006092f
C1372 B.n634 VSUBS 0.006092f
C1373 B.n635 VSUBS 0.013794f
.ends

