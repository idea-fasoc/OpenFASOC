* NGSPICE file created from diff_pair_sample_1461.ext - technology: sky130A

.subckt diff_pair_sample_1461 VTAIL VN VP B VDD2 VDD1
X0 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.88
X1 VDD1.t7 VP.t0 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.88
X2 VTAIL.t5 VN.t0 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.88
X3 VTAIL.t14 VN.t1 VDD2.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X4 VTAIL.t15 VN.t2 VDD2.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X5 VDD2.t4 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X6 VTAIL.t6 VP.t1 VDD1.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X7 VDD2.t3 VN.t4 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.88
X8 VDD1.t5 VP.t2 VTAIL.t8 B.t0 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X9 VDD1.t4 VP.t3 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X10 VDD1.t3 VP.t4 VTAIL.t10 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.88
X11 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.88
X12 VDD2.t2 VN.t5 VTAIL.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=5.9436 ps=31.26 w=15.24 l=0.88
X13 VTAIL.t2 VN.t6 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.88
X14 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.88
X15 VTAIL.t11 VP.t5 VDD1.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.88
X16 VTAIL.t12 VP.t6 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=2.5146 ps=15.57 w=15.24 l=0.88
X17 VTAIL.t13 VP.t7 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X18 VDD2.t0 VN.t7 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.5146 pd=15.57 as=2.5146 ps=15.57 w=15.24 l=0.88
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.9436 pd=31.26 as=0 ps=0 w=15.24 l=0.88
R0 B.n193 B.t19 619.404
R1 B.n187 B.t12 619.404
R2 B.n78 B.t16 619.404
R3 B.n85 B.t8 619.404
R4 B.n559 B.n558 585
R5 B.n561 B.n111 585
R6 B.n564 B.n563 585
R7 B.n565 B.n110 585
R8 B.n567 B.n566 585
R9 B.n569 B.n109 585
R10 B.n572 B.n571 585
R11 B.n573 B.n108 585
R12 B.n575 B.n574 585
R13 B.n577 B.n107 585
R14 B.n580 B.n579 585
R15 B.n581 B.n106 585
R16 B.n583 B.n582 585
R17 B.n585 B.n105 585
R18 B.n588 B.n587 585
R19 B.n589 B.n104 585
R20 B.n591 B.n590 585
R21 B.n593 B.n103 585
R22 B.n596 B.n595 585
R23 B.n597 B.n102 585
R24 B.n599 B.n598 585
R25 B.n601 B.n101 585
R26 B.n604 B.n603 585
R27 B.n605 B.n100 585
R28 B.n607 B.n606 585
R29 B.n609 B.n99 585
R30 B.n612 B.n611 585
R31 B.n613 B.n98 585
R32 B.n615 B.n614 585
R33 B.n617 B.n97 585
R34 B.n620 B.n619 585
R35 B.n621 B.n96 585
R36 B.n623 B.n622 585
R37 B.n625 B.n95 585
R38 B.n628 B.n627 585
R39 B.n629 B.n94 585
R40 B.n631 B.n630 585
R41 B.n633 B.n93 585
R42 B.n636 B.n635 585
R43 B.n637 B.n92 585
R44 B.n639 B.n638 585
R45 B.n641 B.n91 585
R46 B.n644 B.n643 585
R47 B.n645 B.n90 585
R48 B.n647 B.n646 585
R49 B.n649 B.n89 585
R50 B.n652 B.n651 585
R51 B.n653 B.n88 585
R52 B.n655 B.n654 585
R53 B.n657 B.n87 585
R54 B.n660 B.n659 585
R55 B.n662 B.n84 585
R56 B.n664 B.n663 585
R57 B.n666 B.n83 585
R58 B.n669 B.n668 585
R59 B.n670 B.n82 585
R60 B.n672 B.n671 585
R61 B.n674 B.n81 585
R62 B.n677 B.n676 585
R63 B.n678 B.n77 585
R64 B.n680 B.n679 585
R65 B.n682 B.n76 585
R66 B.n685 B.n684 585
R67 B.n686 B.n75 585
R68 B.n688 B.n687 585
R69 B.n690 B.n74 585
R70 B.n693 B.n692 585
R71 B.n694 B.n73 585
R72 B.n696 B.n695 585
R73 B.n698 B.n72 585
R74 B.n701 B.n700 585
R75 B.n702 B.n71 585
R76 B.n704 B.n703 585
R77 B.n706 B.n70 585
R78 B.n709 B.n708 585
R79 B.n710 B.n69 585
R80 B.n712 B.n711 585
R81 B.n714 B.n68 585
R82 B.n717 B.n716 585
R83 B.n718 B.n67 585
R84 B.n720 B.n719 585
R85 B.n722 B.n66 585
R86 B.n725 B.n724 585
R87 B.n726 B.n65 585
R88 B.n728 B.n727 585
R89 B.n730 B.n64 585
R90 B.n733 B.n732 585
R91 B.n734 B.n63 585
R92 B.n736 B.n735 585
R93 B.n738 B.n62 585
R94 B.n741 B.n740 585
R95 B.n742 B.n61 585
R96 B.n744 B.n743 585
R97 B.n746 B.n60 585
R98 B.n749 B.n748 585
R99 B.n750 B.n59 585
R100 B.n752 B.n751 585
R101 B.n754 B.n58 585
R102 B.n757 B.n756 585
R103 B.n758 B.n57 585
R104 B.n760 B.n759 585
R105 B.n762 B.n56 585
R106 B.n765 B.n764 585
R107 B.n766 B.n55 585
R108 B.n768 B.n767 585
R109 B.n770 B.n54 585
R110 B.n773 B.n772 585
R111 B.n774 B.n53 585
R112 B.n776 B.n775 585
R113 B.n778 B.n52 585
R114 B.n781 B.n780 585
R115 B.n782 B.n51 585
R116 B.n557 B.n49 585
R117 B.n785 B.n49 585
R118 B.n556 B.n48 585
R119 B.n786 B.n48 585
R120 B.n555 B.n47 585
R121 B.n787 B.n47 585
R122 B.n554 B.n553 585
R123 B.n553 B.n43 585
R124 B.n552 B.n42 585
R125 B.n793 B.n42 585
R126 B.n551 B.n41 585
R127 B.n794 B.n41 585
R128 B.n550 B.n40 585
R129 B.n795 B.n40 585
R130 B.n549 B.n548 585
R131 B.n548 B.n36 585
R132 B.n547 B.n35 585
R133 B.n801 B.n35 585
R134 B.n546 B.n34 585
R135 B.n802 B.n34 585
R136 B.n545 B.n33 585
R137 B.n803 B.n33 585
R138 B.n544 B.n543 585
R139 B.n543 B.n32 585
R140 B.n542 B.n28 585
R141 B.n809 B.n28 585
R142 B.n541 B.n27 585
R143 B.n810 B.n27 585
R144 B.n540 B.n26 585
R145 B.n811 B.n26 585
R146 B.n539 B.n538 585
R147 B.n538 B.n25 585
R148 B.n537 B.n21 585
R149 B.n817 B.n21 585
R150 B.n536 B.n20 585
R151 B.n818 B.n20 585
R152 B.n535 B.n19 585
R153 B.n819 B.n19 585
R154 B.n534 B.n533 585
R155 B.n533 B.n18 585
R156 B.n532 B.n14 585
R157 B.n825 B.n14 585
R158 B.n531 B.n13 585
R159 B.n826 B.n13 585
R160 B.n530 B.n12 585
R161 B.n827 B.n12 585
R162 B.n529 B.n528 585
R163 B.n528 B.n8 585
R164 B.n527 B.n7 585
R165 B.n833 B.n7 585
R166 B.n526 B.n6 585
R167 B.n834 B.n6 585
R168 B.n525 B.n5 585
R169 B.n835 B.n5 585
R170 B.n524 B.n523 585
R171 B.n523 B.n4 585
R172 B.n522 B.n112 585
R173 B.n522 B.n521 585
R174 B.n512 B.n113 585
R175 B.n114 B.n113 585
R176 B.n514 B.n513 585
R177 B.n515 B.n514 585
R178 B.n511 B.n119 585
R179 B.n119 B.n118 585
R180 B.n510 B.n509 585
R181 B.n509 B.n508 585
R182 B.n121 B.n120 585
R183 B.n501 B.n121 585
R184 B.n500 B.n499 585
R185 B.n502 B.n500 585
R186 B.n498 B.n126 585
R187 B.n126 B.n125 585
R188 B.n497 B.n496 585
R189 B.n496 B.n495 585
R190 B.n128 B.n127 585
R191 B.n488 B.n128 585
R192 B.n487 B.n486 585
R193 B.n489 B.n487 585
R194 B.n485 B.n133 585
R195 B.n133 B.n132 585
R196 B.n484 B.n483 585
R197 B.n483 B.n482 585
R198 B.n135 B.n134 585
R199 B.n475 B.n135 585
R200 B.n474 B.n473 585
R201 B.n476 B.n474 585
R202 B.n472 B.n140 585
R203 B.n140 B.n139 585
R204 B.n471 B.n470 585
R205 B.n470 B.n469 585
R206 B.n142 B.n141 585
R207 B.n143 B.n142 585
R208 B.n462 B.n461 585
R209 B.n463 B.n462 585
R210 B.n460 B.n147 585
R211 B.n151 B.n147 585
R212 B.n459 B.n458 585
R213 B.n458 B.n457 585
R214 B.n149 B.n148 585
R215 B.n150 B.n149 585
R216 B.n450 B.n449 585
R217 B.n451 B.n450 585
R218 B.n448 B.n156 585
R219 B.n156 B.n155 585
R220 B.n447 B.n446 585
R221 B.n446 B.n445 585
R222 B.n442 B.n160 585
R223 B.n441 B.n440 585
R224 B.n438 B.n161 585
R225 B.n438 B.n159 585
R226 B.n437 B.n436 585
R227 B.n435 B.n434 585
R228 B.n433 B.n163 585
R229 B.n431 B.n430 585
R230 B.n429 B.n164 585
R231 B.n428 B.n427 585
R232 B.n425 B.n165 585
R233 B.n423 B.n422 585
R234 B.n421 B.n166 585
R235 B.n420 B.n419 585
R236 B.n417 B.n167 585
R237 B.n415 B.n414 585
R238 B.n413 B.n168 585
R239 B.n412 B.n411 585
R240 B.n409 B.n169 585
R241 B.n407 B.n406 585
R242 B.n405 B.n170 585
R243 B.n404 B.n403 585
R244 B.n401 B.n171 585
R245 B.n399 B.n398 585
R246 B.n397 B.n172 585
R247 B.n396 B.n395 585
R248 B.n393 B.n173 585
R249 B.n391 B.n390 585
R250 B.n389 B.n174 585
R251 B.n388 B.n387 585
R252 B.n385 B.n175 585
R253 B.n383 B.n382 585
R254 B.n381 B.n176 585
R255 B.n380 B.n379 585
R256 B.n377 B.n177 585
R257 B.n375 B.n374 585
R258 B.n373 B.n178 585
R259 B.n372 B.n371 585
R260 B.n369 B.n179 585
R261 B.n367 B.n366 585
R262 B.n365 B.n180 585
R263 B.n364 B.n363 585
R264 B.n361 B.n181 585
R265 B.n359 B.n358 585
R266 B.n357 B.n182 585
R267 B.n356 B.n355 585
R268 B.n353 B.n183 585
R269 B.n351 B.n350 585
R270 B.n349 B.n184 585
R271 B.n348 B.n347 585
R272 B.n345 B.n185 585
R273 B.n343 B.n342 585
R274 B.n340 B.n186 585
R275 B.n339 B.n338 585
R276 B.n336 B.n189 585
R277 B.n334 B.n333 585
R278 B.n332 B.n190 585
R279 B.n331 B.n330 585
R280 B.n328 B.n191 585
R281 B.n326 B.n325 585
R282 B.n324 B.n192 585
R283 B.n323 B.n322 585
R284 B.n320 B.n319 585
R285 B.n318 B.n317 585
R286 B.n316 B.n197 585
R287 B.n314 B.n313 585
R288 B.n312 B.n198 585
R289 B.n311 B.n310 585
R290 B.n308 B.n199 585
R291 B.n306 B.n305 585
R292 B.n304 B.n200 585
R293 B.n303 B.n302 585
R294 B.n300 B.n201 585
R295 B.n298 B.n297 585
R296 B.n296 B.n202 585
R297 B.n295 B.n294 585
R298 B.n292 B.n203 585
R299 B.n290 B.n289 585
R300 B.n288 B.n204 585
R301 B.n287 B.n286 585
R302 B.n284 B.n205 585
R303 B.n282 B.n281 585
R304 B.n280 B.n206 585
R305 B.n279 B.n278 585
R306 B.n276 B.n207 585
R307 B.n274 B.n273 585
R308 B.n272 B.n208 585
R309 B.n271 B.n270 585
R310 B.n268 B.n209 585
R311 B.n266 B.n265 585
R312 B.n264 B.n210 585
R313 B.n263 B.n262 585
R314 B.n260 B.n211 585
R315 B.n258 B.n257 585
R316 B.n256 B.n212 585
R317 B.n255 B.n254 585
R318 B.n252 B.n213 585
R319 B.n250 B.n249 585
R320 B.n248 B.n214 585
R321 B.n247 B.n246 585
R322 B.n244 B.n215 585
R323 B.n242 B.n241 585
R324 B.n240 B.n216 585
R325 B.n239 B.n238 585
R326 B.n236 B.n217 585
R327 B.n234 B.n233 585
R328 B.n232 B.n218 585
R329 B.n231 B.n230 585
R330 B.n228 B.n219 585
R331 B.n226 B.n225 585
R332 B.n224 B.n220 585
R333 B.n223 B.n222 585
R334 B.n158 B.n157 585
R335 B.n159 B.n158 585
R336 B.n444 B.n443 585
R337 B.n445 B.n444 585
R338 B.n154 B.n153 585
R339 B.n155 B.n154 585
R340 B.n453 B.n452 585
R341 B.n452 B.n451 585
R342 B.n454 B.n152 585
R343 B.n152 B.n150 585
R344 B.n456 B.n455 585
R345 B.n457 B.n456 585
R346 B.n146 B.n145 585
R347 B.n151 B.n146 585
R348 B.n465 B.n464 585
R349 B.n464 B.n463 585
R350 B.n466 B.n144 585
R351 B.n144 B.n143 585
R352 B.n468 B.n467 585
R353 B.n469 B.n468 585
R354 B.n138 B.n137 585
R355 B.n139 B.n138 585
R356 B.n478 B.n477 585
R357 B.n477 B.n476 585
R358 B.n479 B.n136 585
R359 B.n475 B.n136 585
R360 B.n481 B.n480 585
R361 B.n482 B.n481 585
R362 B.n131 B.n130 585
R363 B.n132 B.n131 585
R364 B.n491 B.n490 585
R365 B.n490 B.n489 585
R366 B.n492 B.n129 585
R367 B.n488 B.n129 585
R368 B.n494 B.n493 585
R369 B.n495 B.n494 585
R370 B.n124 B.n123 585
R371 B.n125 B.n124 585
R372 B.n504 B.n503 585
R373 B.n503 B.n502 585
R374 B.n505 B.n122 585
R375 B.n501 B.n122 585
R376 B.n507 B.n506 585
R377 B.n508 B.n507 585
R378 B.n117 B.n116 585
R379 B.n118 B.n117 585
R380 B.n517 B.n516 585
R381 B.n516 B.n515 585
R382 B.n518 B.n115 585
R383 B.n115 B.n114 585
R384 B.n520 B.n519 585
R385 B.n521 B.n520 585
R386 B.n2 B.n0 585
R387 B.n4 B.n2 585
R388 B.n3 B.n1 585
R389 B.n834 B.n3 585
R390 B.n832 B.n831 585
R391 B.n833 B.n832 585
R392 B.n830 B.n9 585
R393 B.n9 B.n8 585
R394 B.n829 B.n828 585
R395 B.n828 B.n827 585
R396 B.n11 B.n10 585
R397 B.n826 B.n11 585
R398 B.n824 B.n823 585
R399 B.n825 B.n824 585
R400 B.n822 B.n15 585
R401 B.n18 B.n15 585
R402 B.n821 B.n820 585
R403 B.n820 B.n819 585
R404 B.n17 B.n16 585
R405 B.n818 B.n17 585
R406 B.n816 B.n815 585
R407 B.n817 B.n816 585
R408 B.n814 B.n22 585
R409 B.n25 B.n22 585
R410 B.n813 B.n812 585
R411 B.n812 B.n811 585
R412 B.n24 B.n23 585
R413 B.n810 B.n24 585
R414 B.n808 B.n807 585
R415 B.n809 B.n808 585
R416 B.n806 B.n29 585
R417 B.n32 B.n29 585
R418 B.n805 B.n804 585
R419 B.n804 B.n803 585
R420 B.n31 B.n30 585
R421 B.n802 B.n31 585
R422 B.n800 B.n799 585
R423 B.n801 B.n800 585
R424 B.n798 B.n37 585
R425 B.n37 B.n36 585
R426 B.n797 B.n796 585
R427 B.n796 B.n795 585
R428 B.n39 B.n38 585
R429 B.n794 B.n39 585
R430 B.n792 B.n791 585
R431 B.n793 B.n792 585
R432 B.n790 B.n44 585
R433 B.n44 B.n43 585
R434 B.n789 B.n788 585
R435 B.n788 B.n787 585
R436 B.n46 B.n45 585
R437 B.n786 B.n46 585
R438 B.n784 B.n783 585
R439 B.n785 B.n784 585
R440 B.n837 B.n836 585
R441 B.n836 B.n835 585
R442 B.n444 B.n160 473.281
R443 B.n784 B.n51 473.281
R444 B.n446 B.n158 473.281
R445 B.n559 B.n49 473.281
R446 B.n560 B.n50 256.663
R447 B.n562 B.n50 256.663
R448 B.n568 B.n50 256.663
R449 B.n570 B.n50 256.663
R450 B.n576 B.n50 256.663
R451 B.n578 B.n50 256.663
R452 B.n584 B.n50 256.663
R453 B.n586 B.n50 256.663
R454 B.n592 B.n50 256.663
R455 B.n594 B.n50 256.663
R456 B.n600 B.n50 256.663
R457 B.n602 B.n50 256.663
R458 B.n608 B.n50 256.663
R459 B.n610 B.n50 256.663
R460 B.n616 B.n50 256.663
R461 B.n618 B.n50 256.663
R462 B.n624 B.n50 256.663
R463 B.n626 B.n50 256.663
R464 B.n632 B.n50 256.663
R465 B.n634 B.n50 256.663
R466 B.n640 B.n50 256.663
R467 B.n642 B.n50 256.663
R468 B.n648 B.n50 256.663
R469 B.n650 B.n50 256.663
R470 B.n656 B.n50 256.663
R471 B.n658 B.n50 256.663
R472 B.n665 B.n50 256.663
R473 B.n667 B.n50 256.663
R474 B.n673 B.n50 256.663
R475 B.n675 B.n50 256.663
R476 B.n681 B.n50 256.663
R477 B.n683 B.n50 256.663
R478 B.n689 B.n50 256.663
R479 B.n691 B.n50 256.663
R480 B.n697 B.n50 256.663
R481 B.n699 B.n50 256.663
R482 B.n705 B.n50 256.663
R483 B.n707 B.n50 256.663
R484 B.n713 B.n50 256.663
R485 B.n715 B.n50 256.663
R486 B.n721 B.n50 256.663
R487 B.n723 B.n50 256.663
R488 B.n729 B.n50 256.663
R489 B.n731 B.n50 256.663
R490 B.n737 B.n50 256.663
R491 B.n739 B.n50 256.663
R492 B.n745 B.n50 256.663
R493 B.n747 B.n50 256.663
R494 B.n753 B.n50 256.663
R495 B.n755 B.n50 256.663
R496 B.n761 B.n50 256.663
R497 B.n763 B.n50 256.663
R498 B.n769 B.n50 256.663
R499 B.n771 B.n50 256.663
R500 B.n777 B.n50 256.663
R501 B.n779 B.n50 256.663
R502 B.n439 B.n159 256.663
R503 B.n162 B.n159 256.663
R504 B.n432 B.n159 256.663
R505 B.n426 B.n159 256.663
R506 B.n424 B.n159 256.663
R507 B.n418 B.n159 256.663
R508 B.n416 B.n159 256.663
R509 B.n410 B.n159 256.663
R510 B.n408 B.n159 256.663
R511 B.n402 B.n159 256.663
R512 B.n400 B.n159 256.663
R513 B.n394 B.n159 256.663
R514 B.n392 B.n159 256.663
R515 B.n386 B.n159 256.663
R516 B.n384 B.n159 256.663
R517 B.n378 B.n159 256.663
R518 B.n376 B.n159 256.663
R519 B.n370 B.n159 256.663
R520 B.n368 B.n159 256.663
R521 B.n362 B.n159 256.663
R522 B.n360 B.n159 256.663
R523 B.n354 B.n159 256.663
R524 B.n352 B.n159 256.663
R525 B.n346 B.n159 256.663
R526 B.n344 B.n159 256.663
R527 B.n337 B.n159 256.663
R528 B.n335 B.n159 256.663
R529 B.n329 B.n159 256.663
R530 B.n327 B.n159 256.663
R531 B.n321 B.n159 256.663
R532 B.n196 B.n159 256.663
R533 B.n315 B.n159 256.663
R534 B.n309 B.n159 256.663
R535 B.n307 B.n159 256.663
R536 B.n301 B.n159 256.663
R537 B.n299 B.n159 256.663
R538 B.n293 B.n159 256.663
R539 B.n291 B.n159 256.663
R540 B.n285 B.n159 256.663
R541 B.n283 B.n159 256.663
R542 B.n277 B.n159 256.663
R543 B.n275 B.n159 256.663
R544 B.n269 B.n159 256.663
R545 B.n267 B.n159 256.663
R546 B.n261 B.n159 256.663
R547 B.n259 B.n159 256.663
R548 B.n253 B.n159 256.663
R549 B.n251 B.n159 256.663
R550 B.n245 B.n159 256.663
R551 B.n243 B.n159 256.663
R552 B.n237 B.n159 256.663
R553 B.n235 B.n159 256.663
R554 B.n229 B.n159 256.663
R555 B.n227 B.n159 256.663
R556 B.n221 B.n159 256.663
R557 B.n444 B.n154 163.367
R558 B.n452 B.n154 163.367
R559 B.n452 B.n152 163.367
R560 B.n456 B.n152 163.367
R561 B.n456 B.n146 163.367
R562 B.n464 B.n146 163.367
R563 B.n464 B.n144 163.367
R564 B.n468 B.n144 163.367
R565 B.n468 B.n138 163.367
R566 B.n477 B.n138 163.367
R567 B.n477 B.n136 163.367
R568 B.n481 B.n136 163.367
R569 B.n481 B.n131 163.367
R570 B.n490 B.n131 163.367
R571 B.n490 B.n129 163.367
R572 B.n494 B.n129 163.367
R573 B.n494 B.n124 163.367
R574 B.n503 B.n124 163.367
R575 B.n503 B.n122 163.367
R576 B.n507 B.n122 163.367
R577 B.n507 B.n117 163.367
R578 B.n516 B.n117 163.367
R579 B.n516 B.n115 163.367
R580 B.n520 B.n115 163.367
R581 B.n520 B.n2 163.367
R582 B.n836 B.n2 163.367
R583 B.n836 B.n3 163.367
R584 B.n832 B.n3 163.367
R585 B.n832 B.n9 163.367
R586 B.n828 B.n9 163.367
R587 B.n828 B.n11 163.367
R588 B.n824 B.n11 163.367
R589 B.n824 B.n15 163.367
R590 B.n820 B.n15 163.367
R591 B.n820 B.n17 163.367
R592 B.n816 B.n17 163.367
R593 B.n816 B.n22 163.367
R594 B.n812 B.n22 163.367
R595 B.n812 B.n24 163.367
R596 B.n808 B.n24 163.367
R597 B.n808 B.n29 163.367
R598 B.n804 B.n29 163.367
R599 B.n804 B.n31 163.367
R600 B.n800 B.n31 163.367
R601 B.n800 B.n37 163.367
R602 B.n796 B.n37 163.367
R603 B.n796 B.n39 163.367
R604 B.n792 B.n39 163.367
R605 B.n792 B.n44 163.367
R606 B.n788 B.n44 163.367
R607 B.n788 B.n46 163.367
R608 B.n784 B.n46 163.367
R609 B.n440 B.n438 163.367
R610 B.n438 B.n437 163.367
R611 B.n434 B.n433 163.367
R612 B.n431 B.n164 163.367
R613 B.n427 B.n425 163.367
R614 B.n423 B.n166 163.367
R615 B.n419 B.n417 163.367
R616 B.n415 B.n168 163.367
R617 B.n411 B.n409 163.367
R618 B.n407 B.n170 163.367
R619 B.n403 B.n401 163.367
R620 B.n399 B.n172 163.367
R621 B.n395 B.n393 163.367
R622 B.n391 B.n174 163.367
R623 B.n387 B.n385 163.367
R624 B.n383 B.n176 163.367
R625 B.n379 B.n377 163.367
R626 B.n375 B.n178 163.367
R627 B.n371 B.n369 163.367
R628 B.n367 B.n180 163.367
R629 B.n363 B.n361 163.367
R630 B.n359 B.n182 163.367
R631 B.n355 B.n353 163.367
R632 B.n351 B.n184 163.367
R633 B.n347 B.n345 163.367
R634 B.n343 B.n186 163.367
R635 B.n338 B.n336 163.367
R636 B.n334 B.n190 163.367
R637 B.n330 B.n328 163.367
R638 B.n326 B.n192 163.367
R639 B.n322 B.n320 163.367
R640 B.n317 B.n316 163.367
R641 B.n314 B.n198 163.367
R642 B.n310 B.n308 163.367
R643 B.n306 B.n200 163.367
R644 B.n302 B.n300 163.367
R645 B.n298 B.n202 163.367
R646 B.n294 B.n292 163.367
R647 B.n290 B.n204 163.367
R648 B.n286 B.n284 163.367
R649 B.n282 B.n206 163.367
R650 B.n278 B.n276 163.367
R651 B.n274 B.n208 163.367
R652 B.n270 B.n268 163.367
R653 B.n266 B.n210 163.367
R654 B.n262 B.n260 163.367
R655 B.n258 B.n212 163.367
R656 B.n254 B.n252 163.367
R657 B.n250 B.n214 163.367
R658 B.n246 B.n244 163.367
R659 B.n242 B.n216 163.367
R660 B.n238 B.n236 163.367
R661 B.n234 B.n218 163.367
R662 B.n230 B.n228 163.367
R663 B.n226 B.n220 163.367
R664 B.n222 B.n158 163.367
R665 B.n446 B.n156 163.367
R666 B.n450 B.n156 163.367
R667 B.n450 B.n149 163.367
R668 B.n458 B.n149 163.367
R669 B.n458 B.n147 163.367
R670 B.n462 B.n147 163.367
R671 B.n462 B.n142 163.367
R672 B.n470 B.n142 163.367
R673 B.n470 B.n140 163.367
R674 B.n474 B.n140 163.367
R675 B.n474 B.n135 163.367
R676 B.n483 B.n135 163.367
R677 B.n483 B.n133 163.367
R678 B.n487 B.n133 163.367
R679 B.n487 B.n128 163.367
R680 B.n496 B.n128 163.367
R681 B.n496 B.n126 163.367
R682 B.n500 B.n126 163.367
R683 B.n500 B.n121 163.367
R684 B.n509 B.n121 163.367
R685 B.n509 B.n119 163.367
R686 B.n514 B.n119 163.367
R687 B.n514 B.n113 163.367
R688 B.n522 B.n113 163.367
R689 B.n523 B.n522 163.367
R690 B.n523 B.n5 163.367
R691 B.n6 B.n5 163.367
R692 B.n7 B.n6 163.367
R693 B.n528 B.n7 163.367
R694 B.n528 B.n12 163.367
R695 B.n13 B.n12 163.367
R696 B.n14 B.n13 163.367
R697 B.n533 B.n14 163.367
R698 B.n533 B.n19 163.367
R699 B.n20 B.n19 163.367
R700 B.n21 B.n20 163.367
R701 B.n538 B.n21 163.367
R702 B.n538 B.n26 163.367
R703 B.n27 B.n26 163.367
R704 B.n28 B.n27 163.367
R705 B.n543 B.n28 163.367
R706 B.n543 B.n33 163.367
R707 B.n34 B.n33 163.367
R708 B.n35 B.n34 163.367
R709 B.n548 B.n35 163.367
R710 B.n548 B.n40 163.367
R711 B.n41 B.n40 163.367
R712 B.n42 B.n41 163.367
R713 B.n553 B.n42 163.367
R714 B.n553 B.n47 163.367
R715 B.n48 B.n47 163.367
R716 B.n49 B.n48 163.367
R717 B.n780 B.n778 163.367
R718 B.n776 B.n53 163.367
R719 B.n772 B.n770 163.367
R720 B.n768 B.n55 163.367
R721 B.n764 B.n762 163.367
R722 B.n760 B.n57 163.367
R723 B.n756 B.n754 163.367
R724 B.n752 B.n59 163.367
R725 B.n748 B.n746 163.367
R726 B.n744 B.n61 163.367
R727 B.n740 B.n738 163.367
R728 B.n736 B.n63 163.367
R729 B.n732 B.n730 163.367
R730 B.n728 B.n65 163.367
R731 B.n724 B.n722 163.367
R732 B.n720 B.n67 163.367
R733 B.n716 B.n714 163.367
R734 B.n712 B.n69 163.367
R735 B.n708 B.n706 163.367
R736 B.n704 B.n71 163.367
R737 B.n700 B.n698 163.367
R738 B.n696 B.n73 163.367
R739 B.n692 B.n690 163.367
R740 B.n688 B.n75 163.367
R741 B.n684 B.n682 163.367
R742 B.n680 B.n77 163.367
R743 B.n676 B.n674 163.367
R744 B.n672 B.n82 163.367
R745 B.n668 B.n666 163.367
R746 B.n664 B.n84 163.367
R747 B.n659 B.n657 163.367
R748 B.n655 B.n88 163.367
R749 B.n651 B.n649 163.367
R750 B.n647 B.n90 163.367
R751 B.n643 B.n641 163.367
R752 B.n639 B.n92 163.367
R753 B.n635 B.n633 163.367
R754 B.n631 B.n94 163.367
R755 B.n627 B.n625 163.367
R756 B.n623 B.n96 163.367
R757 B.n619 B.n617 163.367
R758 B.n615 B.n98 163.367
R759 B.n611 B.n609 163.367
R760 B.n607 B.n100 163.367
R761 B.n603 B.n601 163.367
R762 B.n599 B.n102 163.367
R763 B.n595 B.n593 163.367
R764 B.n591 B.n104 163.367
R765 B.n587 B.n585 163.367
R766 B.n583 B.n106 163.367
R767 B.n579 B.n577 163.367
R768 B.n575 B.n108 163.367
R769 B.n571 B.n569 163.367
R770 B.n567 B.n110 163.367
R771 B.n563 B.n561 163.367
R772 B.n193 B.t21 96.3406
R773 B.n85 B.t10 96.3406
R774 B.n187 B.t15 96.3208
R775 B.n78 B.t17 96.3208
R776 B.n194 B.t20 72.8739
R777 B.n86 B.t11 72.8739
R778 B.n188 B.t14 72.8542
R779 B.n79 B.t18 72.8542
R780 B.n439 B.n160 71.676
R781 B.n437 B.n162 71.676
R782 B.n433 B.n432 71.676
R783 B.n426 B.n164 71.676
R784 B.n425 B.n424 71.676
R785 B.n418 B.n166 71.676
R786 B.n417 B.n416 71.676
R787 B.n410 B.n168 71.676
R788 B.n409 B.n408 71.676
R789 B.n402 B.n170 71.676
R790 B.n401 B.n400 71.676
R791 B.n394 B.n172 71.676
R792 B.n393 B.n392 71.676
R793 B.n386 B.n174 71.676
R794 B.n385 B.n384 71.676
R795 B.n378 B.n176 71.676
R796 B.n377 B.n376 71.676
R797 B.n370 B.n178 71.676
R798 B.n369 B.n368 71.676
R799 B.n362 B.n180 71.676
R800 B.n361 B.n360 71.676
R801 B.n354 B.n182 71.676
R802 B.n353 B.n352 71.676
R803 B.n346 B.n184 71.676
R804 B.n345 B.n344 71.676
R805 B.n337 B.n186 71.676
R806 B.n336 B.n335 71.676
R807 B.n329 B.n190 71.676
R808 B.n328 B.n327 71.676
R809 B.n321 B.n192 71.676
R810 B.n320 B.n196 71.676
R811 B.n316 B.n315 71.676
R812 B.n309 B.n198 71.676
R813 B.n308 B.n307 71.676
R814 B.n301 B.n200 71.676
R815 B.n300 B.n299 71.676
R816 B.n293 B.n202 71.676
R817 B.n292 B.n291 71.676
R818 B.n285 B.n204 71.676
R819 B.n284 B.n283 71.676
R820 B.n277 B.n206 71.676
R821 B.n276 B.n275 71.676
R822 B.n269 B.n208 71.676
R823 B.n268 B.n267 71.676
R824 B.n261 B.n210 71.676
R825 B.n260 B.n259 71.676
R826 B.n253 B.n212 71.676
R827 B.n252 B.n251 71.676
R828 B.n245 B.n214 71.676
R829 B.n244 B.n243 71.676
R830 B.n237 B.n216 71.676
R831 B.n236 B.n235 71.676
R832 B.n229 B.n218 71.676
R833 B.n228 B.n227 71.676
R834 B.n221 B.n220 71.676
R835 B.n779 B.n51 71.676
R836 B.n778 B.n777 71.676
R837 B.n771 B.n53 71.676
R838 B.n770 B.n769 71.676
R839 B.n763 B.n55 71.676
R840 B.n762 B.n761 71.676
R841 B.n755 B.n57 71.676
R842 B.n754 B.n753 71.676
R843 B.n747 B.n59 71.676
R844 B.n746 B.n745 71.676
R845 B.n739 B.n61 71.676
R846 B.n738 B.n737 71.676
R847 B.n731 B.n63 71.676
R848 B.n730 B.n729 71.676
R849 B.n723 B.n65 71.676
R850 B.n722 B.n721 71.676
R851 B.n715 B.n67 71.676
R852 B.n714 B.n713 71.676
R853 B.n707 B.n69 71.676
R854 B.n706 B.n705 71.676
R855 B.n699 B.n71 71.676
R856 B.n698 B.n697 71.676
R857 B.n691 B.n73 71.676
R858 B.n690 B.n689 71.676
R859 B.n683 B.n75 71.676
R860 B.n682 B.n681 71.676
R861 B.n675 B.n77 71.676
R862 B.n674 B.n673 71.676
R863 B.n667 B.n82 71.676
R864 B.n666 B.n665 71.676
R865 B.n658 B.n84 71.676
R866 B.n657 B.n656 71.676
R867 B.n650 B.n88 71.676
R868 B.n649 B.n648 71.676
R869 B.n642 B.n90 71.676
R870 B.n641 B.n640 71.676
R871 B.n634 B.n92 71.676
R872 B.n633 B.n632 71.676
R873 B.n626 B.n94 71.676
R874 B.n625 B.n624 71.676
R875 B.n618 B.n96 71.676
R876 B.n617 B.n616 71.676
R877 B.n610 B.n98 71.676
R878 B.n609 B.n608 71.676
R879 B.n602 B.n100 71.676
R880 B.n601 B.n600 71.676
R881 B.n594 B.n102 71.676
R882 B.n593 B.n592 71.676
R883 B.n586 B.n104 71.676
R884 B.n585 B.n584 71.676
R885 B.n578 B.n106 71.676
R886 B.n577 B.n576 71.676
R887 B.n570 B.n108 71.676
R888 B.n569 B.n568 71.676
R889 B.n562 B.n110 71.676
R890 B.n561 B.n560 71.676
R891 B.n560 B.n559 71.676
R892 B.n563 B.n562 71.676
R893 B.n568 B.n567 71.676
R894 B.n571 B.n570 71.676
R895 B.n576 B.n575 71.676
R896 B.n579 B.n578 71.676
R897 B.n584 B.n583 71.676
R898 B.n587 B.n586 71.676
R899 B.n592 B.n591 71.676
R900 B.n595 B.n594 71.676
R901 B.n600 B.n599 71.676
R902 B.n603 B.n602 71.676
R903 B.n608 B.n607 71.676
R904 B.n611 B.n610 71.676
R905 B.n616 B.n615 71.676
R906 B.n619 B.n618 71.676
R907 B.n624 B.n623 71.676
R908 B.n627 B.n626 71.676
R909 B.n632 B.n631 71.676
R910 B.n635 B.n634 71.676
R911 B.n640 B.n639 71.676
R912 B.n643 B.n642 71.676
R913 B.n648 B.n647 71.676
R914 B.n651 B.n650 71.676
R915 B.n656 B.n655 71.676
R916 B.n659 B.n658 71.676
R917 B.n665 B.n664 71.676
R918 B.n668 B.n667 71.676
R919 B.n673 B.n672 71.676
R920 B.n676 B.n675 71.676
R921 B.n681 B.n680 71.676
R922 B.n684 B.n683 71.676
R923 B.n689 B.n688 71.676
R924 B.n692 B.n691 71.676
R925 B.n697 B.n696 71.676
R926 B.n700 B.n699 71.676
R927 B.n705 B.n704 71.676
R928 B.n708 B.n707 71.676
R929 B.n713 B.n712 71.676
R930 B.n716 B.n715 71.676
R931 B.n721 B.n720 71.676
R932 B.n724 B.n723 71.676
R933 B.n729 B.n728 71.676
R934 B.n732 B.n731 71.676
R935 B.n737 B.n736 71.676
R936 B.n740 B.n739 71.676
R937 B.n745 B.n744 71.676
R938 B.n748 B.n747 71.676
R939 B.n753 B.n752 71.676
R940 B.n756 B.n755 71.676
R941 B.n761 B.n760 71.676
R942 B.n764 B.n763 71.676
R943 B.n769 B.n768 71.676
R944 B.n772 B.n771 71.676
R945 B.n777 B.n776 71.676
R946 B.n780 B.n779 71.676
R947 B.n440 B.n439 71.676
R948 B.n434 B.n162 71.676
R949 B.n432 B.n431 71.676
R950 B.n427 B.n426 71.676
R951 B.n424 B.n423 71.676
R952 B.n419 B.n418 71.676
R953 B.n416 B.n415 71.676
R954 B.n411 B.n410 71.676
R955 B.n408 B.n407 71.676
R956 B.n403 B.n402 71.676
R957 B.n400 B.n399 71.676
R958 B.n395 B.n394 71.676
R959 B.n392 B.n391 71.676
R960 B.n387 B.n386 71.676
R961 B.n384 B.n383 71.676
R962 B.n379 B.n378 71.676
R963 B.n376 B.n375 71.676
R964 B.n371 B.n370 71.676
R965 B.n368 B.n367 71.676
R966 B.n363 B.n362 71.676
R967 B.n360 B.n359 71.676
R968 B.n355 B.n354 71.676
R969 B.n352 B.n351 71.676
R970 B.n347 B.n346 71.676
R971 B.n344 B.n343 71.676
R972 B.n338 B.n337 71.676
R973 B.n335 B.n334 71.676
R974 B.n330 B.n329 71.676
R975 B.n327 B.n326 71.676
R976 B.n322 B.n321 71.676
R977 B.n317 B.n196 71.676
R978 B.n315 B.n314 71.676
R979 B.n310 B.n309 71.676
R980 B.n307 B.n306 71.676
R981 B.n302 B.n301 71.676
R982 B.n299 B.n298 71.676
R983 B.n294 B.n293 71.676
R984 B.n291 B.n290 71.676
R985 B.n286 B.n285 71.676
R986 B.n283 B.n282 71.676
R987 B.n278 B.n277 71.676
R988 B.n275 B.n274 71.676
R989 B.n270 B.n269 71.676
R990 B.n267 B.n266 71.676
R991 B.n262 B.n261 71.676
R992 B.n259 B.n258 71.676
R993 B.n254 B.n253 71.676
R994 B.n251 B.n250 71.676
R995 B.n246 B.n245 71.676
R996 B.n243 B.n242 71.676
R997 B.n238 B.n237 71.676
R998 B.n235 B.n234 71.676
R999 B.n230 B.n229 71.676
R1000 B.n227 B.n226 71.676
R1001 B.n222 B.n221 71.676
R1002 B.n445 B.n159 62.7351
R1003 B.n785 B.n50 62.7351
R1004 B.n195 B.n194 59.5399
R1005 B.n341 B.n188 59.5399
R1006 B.n80 B.n79 59.5399
R1007 B.n661 B.n86 59.5399
R1008 B.n445 B.n155 36.4616
R1009 B.n451 B.n155 36.4616
R1010 B.n451 B.n150 36.4616
R1011 B.n457 B.n150 36.4616
R1012 B.n457 B.n151 36.4616
R1013 B.n463 B.n143 36.4616
R1014 B.n469 B.n143 36.4616
R1015 B.n469 B.n139 36.4616
R1016 B.n476 B.n139 36.4616
R1017 B.n476 B.n475 36.4616
R1018 B.n482 B.n132 36.4616
R1019 B.n489 B.n132 36.4616
R1020 B.n489 B.n488 36.4616
R1021 B.n495 B.n125 36.4616
R1022 B.n502 B.n125 36.4616
R1023 B.n502 B.n501 36.4616
R1024 B.n508 B.n118 36.4616
R1025 B.n515 B.n118 36.4616
R1026 B.n521 B.n114 36.4616
R1027 B.n521 B.n4 36.4616
R1028 B.n835 B.n4 36.4616
R1029 B.n835 B.n834 36.4616
R1030 B.n834 B.n833 36.4616
R1031 B.n833 B.n8 36.4616
R1032 B.n827 B.n826 36.4616
R1033 B.n826 B.n825 36.4616
R1034 B.n819 B.n18 36.4616
R1035 B.n819 B.n818 36.4616
R1036 B.n818 B.n817 36.4616
R1037 B.n811 B.n25 36.4616
R1038 B.n811 B.n810 36.4616
R1039 B.n810 B.n809 36.4616
R1040 B.n803 B.n32 36.4616
R1041 B.n803 B.n802 36.4616
R1042 B.n802 B.n801 36.4616
R1043 B.n801 B.n36 36.4616
R1044 B.n795 B.n36 36.4616
R1045 B.n794 B.n793 36.4616
R1046 B.n793 B.n43 36.4616
R1047 B.n787 B.n43 36.4616
R1048 B.n787 B.n786 36.4616
R1049 B.n786 B.n785 36.4616
R1050 B.n475 B.t6 34.3169
R1051 B.n508 B.t5 34.3169
R1052 B.n825 B.t1 34.3169
R1053 B.n32 B.t3 34.3169
R1054 B.n783 B.n782 30.7517
R1055 B.n558 B.n557 30.7517
R1056 B.n447 B.n157 30.7517
R1057 B.n443 B.n442 30.7517
R1058 B.n463 B.t13 30.0273
R1059 B.n795 B.t9 30.0273
R1060 B.n194 B.n193 23.4672
R1061 B.n188 B.n187 23.4672
R1062 B.n79 B.n78 23.4672
R1063 B.n86 B.n85 23.4672
R1064 B.n515 B.t7 22.5206
R1065 B.n827 B.t2 22.5206
R1066 B.n488 B.t0 18.2311
R1067 B.n495 B.t0 18.2311
R1068 B.n817 B.t4 18.2311
R1069 B.n25 B.t4 18.2311
R1070 B B.n837 18.0485
R1071 B.t7 B.n114 13.9415
R1072 B.t2 B.n8 13.9415
R1073 B.n782 B.n781 10.6151
R1074 B.n781 B.n52 10.6151
R1075 B.n775 B.n52 10.6151
R1076 B.n775 B.n774 10.6151
R1077 B.n774 B.n773 10.6151
R1078 B.n773 B.n54 10.6151
R1079 B.n767 B.n54 10.6151
R1080 B.n767 B.n766 10.6151
R1081 B.n766 B.n765 10.6151
R1082 B.n765 B.n56 10.6151
R1083 B.n759 B.n56 10.6151
R1084 B.n759 B.n758 10.6151
R1085 B.n758 B.n757 10.6151
R1086 B.n757 B.n58 10.6151
R1087 B.n751 B.n58 10.6151
R1088 B.n751 B.n750 10.6151
R1089 B.n750 B.n749 10.6151
R1090 B.n749 B.n60 10.6151
R1091 B.n743 B.n60 10.6151
R1092 B.n743 B.n742 10.6151
R1093 B.n742 B.n741 10.6151
R1094 B.n741 B.n62 10.6151
R1095 B.n735 B.n62 10.6151
R1096 B.n735 B.n734 10.6151
R1097 B.n734 B.n733 10.6151
R1098 B.n733 B.n64 10.6151
R1099 B.n727 B.n64 10.6151
R1100 B.n727 B.n726 10.6151
R1101 B.n726 B.n725 10.6151
R1102 B.n725 B.n66 10.6151
R1103 B.n719 B.n66 10.6151
R1104 B.n719 B.n718 10.6151
R1105 B.n718 B.n717 10.6151
R1106 B.n717 B.n68 10.6151
R1107 B.n711 B.n68 10.6151
R1108 B.n711 B.n710 10.6151
R1109 B.n710 B.n709 10.6151
R1110 B.n709 B.n70 10.6151
R1111 B.n703 B.n70 10.6151
R1112 B.n703 B.n702 10.6151
R1113 B.n702 B.n701 10.6151
R1114 B.n701 B.n72 10.6151
R1115 B.n695 B.n72 10.6151
R1116 B.n695 B.n694 10.6151
R1117 B.n694 B.n693 10.6151
R1118 B.n693 B.n74 10.6151
R1119 B.n687 B.n74 10.6151
R1120 B.n687 B.n686 10.6151
R1121 B.n686 B.n685 10.6151
R1122 B.n685 B.n76 10.6151
R1123 B.n679 B.n678 10.6151
R1124 B.n678 B.n677 10.6151
R1125 B.n677 B.n81 10.6151
R1126 B.n671 B.n81 10.6151
R1127 B.n671 B.n670 10.6151
R1128 B.n670 B.n669 10.6151
R1129 B.n669 B.n83 10.6151
R1130 B.n663 B.n83 10.6151
R1131 B.n663 B.n662 10.6151
R1132 B.n660 B.n87 10.6151
R1133 B.n654 B.n87 10.6151
R1134 B.n654 B.n653 10.6151
R1135 B.n653 B.n652 10.6151
R1136 B.n652 B.n89 10.6151
R1137 B.n646 B.n89 10.6151
R1138 B.n646 B.n645 10.6151
R1139 B.n645 B.n644 10.6151
R1140 B.n644 B.n91 10.6151
R1141 B.n638 B.n91 10.6151
R1142 B.n638 B.n637 10.6151
R1143 B.n637 B.n636 10.6151
R1144 B.n636 B.n93 10.6151
R1145 B.n630 B.n93 10.6151
R1146 B.n630 B.n629 10.6151
R1147 B.n629 B.n628 10.6151
R1148 B.n628 B.n95 10.6151
R1149 B.n622 B.n95 10.6151
R1150 B.n622 B.n621 10.6151
R1151 B.n621 B.n620 10.6151
R1152 B.n620 B.n97 10.6151
R1153 B.n614 B.n97 10.6151
R1154 B.n614 B.n613 10.6151
R1155 B.n613 B.n612 10.6151
R1156 B.n612 B.n99 10.6151
R1157 B.n606 B.n99 10.6151
R1158 B.n606 B.n605 10.6151
R1159 B.n605 B.n604 10.6151
R1160 B.n604 B.n101 10.6151
R1161 B.n598 B.n101 10.6151
R1162 B.n598 B.n597 10.6151
R1163 B.n597 B.n596 10.6151
R1164 B.n596 B.n103 10.6151
R1165 B.n590 B.n103 10.6151
R1166 B.n590 B.n589 10.6151
R1167 B.n589 B.n588 10.6151
R1168 B.n588 B.n105 10.6151
R1169 B.n582 B.n105 10.6151
R1170 B.n582 B.n581 10.6151
R1171 B.n581 B.n580 10.6151
R1172 B.n580 B.n107 10.6151
R1173 B.n574 B.n107 10.6151
R1174 B.n574 B.n573 10.6151
R1175 B.n573 B.n572 10.6151
R1176 B.n572 B.n109 10.6151
R1177 B.n566 B.n109 10.6151
R1178 B.n566 B.n565 10.6151
R1179 B.n565 B.n564 10.6151
R1180 B.n564 B.n111 10.6151
R1181 B.n558 B.n111 10.6151
R1182 B.n448 B.n447 10.6151
R1183 B.n449 B.n448 10.6151
R1184 B.n449 B.n148 10.6151
R1185 B.n459 B.n148 10.6151
R1186 B.n460 B.n459 10.6151
R1187 B.n461 B.n460 10.6151
R1188 B.n461 B.n141 10.6151
R1189 B.n471 B.n141 10.6151
R1190 B.n472 B.n471 10.6151
R1191 B.n473 B.n472 10.6151
R1192 B.n473 B.n134 10.6151
R1193 B.n484 B.n134 10.6151
R1194 B.n485 B.n484 10.6151
R1195 B.n486 B.n485 10.6151
R1196 B.n486 B.n127 10.6151
R1197 B.n497 B.n127 10.6151
R1198 B.n498 B.n497 10.6151
R1199 B.n499 B.n498 10.6151
R1200 B.n499 B.n120 10.6151
R1201 B.n510 B.n120 10.6151
R1202 B.n511 B.n510 10.6151
R1203 B.n513 B.n511 10.6151
R1204 B.n513 B.n512 10.6151
R1205 B.n512 B.n112 10.6151
R1206 B.n524 B.n112 10.6151
R1207 B.n525 B.n524 10.6151
R1208 B.n526 B.n525 10.6151
R1209 B.n527 B.n526 10.6151
R1210 B.n529 B.n527 10.6151
R1211 B.n530 B.n529 10.6151
R1212 B.n531 B.n530 10.6151
R1213 B.n532 B.n531 10.6151
R1214 B.n534 B.n532 10.6151
R1215 B.n535 B.n534 10.6151
R1216 B.n536 B.n535 10.6151
R1217 B.n537 B.n536 10.6151
R1218 B.n539 B.n537 10.6151
R1219 B.n540 B.n539 10.6151
R1220 B.n541 B.n540 10.6151
R1221 B.n542 B.n541 10.6151
R1222 B.n544 B.n542 10.6151
R1223 B.n545 B.n544 10.6151
R1224 B.n546 B.n545 10.6151
R1225 B.n547 B.n546 10.6151
R1226 B.n549 B.n547 10.6151
R1227 B.n550 B.n549 10.6151
R1228 B.n551 B.n550 10.6151
R1229 B.n552 B.n551 10.6151
R1230 B.n554 B.n552 10.6151
R1231 B.n555 B.n554 10.6151
R1232 B.n556 B.n555 10.6151
R1233 B.n557 B.n556 10.6151
R1234 B.n442 B.n441 10.6151
R1235 B.n441 B.n161 10.6151
R1236 B.n436 B.n161 10.6151
R1237 B.n436 B.n435 10.6151
R1238 B.n435 B.n163 10.6151
R1239 B.n430 B.n163 10.6151
R1240 B.n430 B.n429 10.6151
R1241 B.n429 B.n428 10.6151
R1242 B.n428 B.n165 10.6151
R1243 B.n422 B.n165 10.6151
R1244 B.n422 B.n421 10.6151
R1245 B.n421 B.n420 10.6151
R1246 B.n420 B.n167 10.6151
R1247 B.n414 B.n167 10.6151
R1248 B.n414 B.n413 10.6151
R1249 B.n413 B.n412 10.6151
R1250 B.n412 B.n169 10.6151
R1251 B.n406 B.n169 10.6151
R1252 B.n406 B.n405 10.6151
R1253 B.n405 B.n404 10.6151
R1254 B.n404 B.n171 10.6151
R1255 B.n398 B.n171 10.6151
R1256 B.n398 B.n397 10.6151
R1257 B.n397 B.n396 10.6151
R1258 B.n396 B.n173 10.6151
R1259 B.n390 B.n173 10.6151
R1260 B.n390 B.n389 10.6151
R1261 B.n389 B.n388 10.6151
R1262 B.n388 B.n175 10.6151
R1263 B.n382 B.n175 10.6151
R1264 B.n382 B.n381 10.6151
R1265 B.n381 B.n380 10.6151
R1266 B.n380 B.n177 10.6151
R1267 B.n374 B.n177 10.6151
R1268 B.n374 B.n373 10.6151
R1269 B.n373 B.n372 10.6151
R1270 B.n372 B.n179 10.6151
R1271 B.n366 B.n179 10.6151
R1272 B.n366 B.n365 10.6151
R1273 B.n365 B.n364 10.6151
R1274 B.n364 B.n181 10.6151
R1275 B.n358 B.n181 10.6151
R1276 B.n358 B.n357 10.6151
R1277 B.n357 B.n356 10.6151
R1278 B.n356 B.n183 10.6151
R1279 B.n350 B.n183 10.6151
R1280 B.n350 B.n349 10.6151
R1281 B.n349 B.n348 10.6151
R1282 B.n348 B.n185 10.6151
R1283 B.n342 B.n185 10.6151
R1284 B.n340 B.n339 10.6151
R1285 B.n339 B.n189 10.6151
R1286 B.n333 B.n189 10.6151
R1287 B.n333 B.n332 10.6151
R1288 B.n332 B.n331 10.6151
R1289 B.n331 B.n191 10.6151
R1290 B.n325 B.n191 10.6151
R1291 B.n325 B.n324 10.6151
R1292 B.n324 B.n323 10.6151
R1293 B.n319 B.n318 10.6151
R1294 B.n318 B.n197 10.6151
R1295 B.n313 B.n197 10.6151
R1296 B.n313 B.n312 10.6151
R1297 B.n312 B.n311 10.6151
R1298 B.n311 B.n199 10.6151
R1299 B.n305 B.n199 10.6151
R1300 B.n305 B.n304 10.6151
R1301 B.n304 B.n303 10.6151
R1302 B.n303 B.n201 10.6151
R1303 B.n297 B.n201 10.6151
R1304 B.n297 B.n296 10.6151
R1305 B.n296 B.n295 10.6151
R1306 B.n295 B.n203 10.6151
R1307 B.n289 B.n203 10.6151
R1308 B.n289 B.n288 10.6151
R1309 B.n288 B.n287 10.6151
R1310 B.n287 B.n205 10.6151
R1311 B.n281 B.n205 10.6151
R1312 B.n281 B.n280 10.6151
R1313 B.n280 B.n279 10.6151
R1314 B.n279 B.n207 10.6151
R1315 B.n273 B.n207 10.6151
R1316 B.n273 B.n272 10.6151
R1317 B.n272 B.n271 10.6151
R1318 B.n271 B.n209 10.6151
R1319 B.n265 B.n209 10.6151
R1320 B.n265 B.n264 10.6151
R1321 B.n264 B.n263 10.6151
R1322 B.n263 B.n211 10.6151
R1323 B.n257 B.n211 10.6151
R1324 B.n257 B.n256 10.6151
R1325 B.n256 B.n255 10.6151
R1326 B.n255 B.n213 10.6151
R1327 B.n249 B.n213 10.6151
R1328 B.n249 B.n248 10.6151
R1329 B.n248 B.n247 10.6151
R1330 B.n247 B.n215 10.6151
R1331 B.n241 B.n215 10.6151
R1332 B.n241 B.n240 10.6151
R1333 B.n240 B.n239 10.6151
R1334 B.n239 B.n217 10.6151
R1335 B.n233 B.n217 10.6151
R1336 B.n233 B.n232 10.6151
R1337 B.n232 B.n231 10.6151
R1338 B.n231 B.n219 10.6151
R1339 B.n225 B.n219 10.6151
R1340 B.n225 B.n224 10.6151
R1341 B.n224 B.n223 10.6151
R1342 B.n223 B.n157 10.6151
R1343 B.n443 B.n153 10.6151
R1344 B.n453 B.n153 10.6151
R1345 B.n454 B.n453 10.6151
R1346 B.n455 B.n454 10.6151
R1347 B.n455 B.n145 10.6151
R1348 B.n465 B.n145 10.6151
R1349 B.n466 B.n465 10.6151
R1350 B.n467 B.n466 10.6151
R1351 B.n467 B.n137 10.6151
R1352 B.n478 B.n137 10.6151
R1353 B.n479 B.n478 10.6151
R1354 B.n480 B.n479 10.6151
R1355 B.n480 B.n130 10.6151
R1356 B.n491 B.n130 10.6151
R1357 B.n492 B.n491 10.6151
R1358 B.n493 B.n492 10.6151
R1359 B.n493 B.n123 10.6151
R1360 B.n504 B.n123 10.6151
R1361 B.n505 B.n504 10.6151
R1362 B.n506 B.n505 10.6151
R1363 B.n506 B.n116 10.6151
R1364 B.n517 B.n116 10.6151
R1365 B.n518 B.n517 10.6151
R1366 B.n519 B.n518 10.6151
R1367 B.n519 B.n0 10.6151
R1368 B.n831 B.n1 10.6151
R1369 B.n831 B.n830 10.6151
R1370 B.n830 B.n829 10.6151
R1371 B.n829 B.n10 10.6151
R1372 B.n823 B.n10 10.6151
R1373 B.n823 B.n822 10.6151
R1374 B.n822 B.n821 10.6151
R1375 B.n821 B.n16 10.6151
R1376 B.n815 B.n16 10.6151
R1377 B.n815 B.n814 10.6151
R1378 B.n814 B.n813 10.6151
R1379 B.n813 B.n23 10.6151
R1380 B.n807 B.n23 10.6151
R1381 B.n807 B.n806 10.6151
R1382 B.n806 B.n805 10.6151
R1383 B.n805 B.n30 10.6151
R1384 B.n799 B.n30 10.6151
R1385 B.n799 B.n798 10.6151
R1386 B.n798 B.n797 10.6151
R1387 B.n797 B.n38 10.6151
R1388 B.n791 B.n38 10.6151
R1389 B.n791 B.n790 10.6151
R1390 B.n790 B.n789 10.6151
R1391 B.n789 B.n45 10.6151
R1392 B.n783 B.n45 10.6151
R1393 B.n80 B.n76 9.36635
R1394 B.n661 B.n660 9.36635
R1395 B.n342 B.n341 9.36635
R1396 B.n319 B.n195 9.36635
R1397 B.n151 B.t13 6.43482
R1398 B.t9 B.n794 6.43482
R1399 B.n837 B.n0 2.81026
R1400 B.n837 B.n1 2.81026
R1401 B.n482 B.t6 2.14527
R1402 B.n501 B.t5 2.14527
R1403 B.n18 B.t1 2.14527
R1404 B.n809 B.t3 2.14527
R1405 B.n679 B.n80 1.24928
R1406 B.n662 B.n661 1.24928
R1407 B.n341 B.n340 1.24928
R1408 B.n323 B.n195 1.24928
R1409 VP.n7 VP.t6 484.625
R1410 VP.n17 VP.t5 462.009
R1411 VP.n29 VP.t4 462.009
R1412 VP.n15 VP.t0 462.009
R1413 VP.n22 VP.t2 417.368
R1414 VP.n1 VP.t7 417.368
R1415 VP.n5 VP.t1 417.368
R1416 VP.n8 VP.t3 417.368
R1417 VP.n30 VP.n29 161.3
R1418 VP.n9 VP.n6 161.3
R1419 VP.n11 VP.n10 161.3
R1420 VP.n13 VP.n12 161.3
R1421 VP.n14 VP.n4 161.3
R1422 VP.n16 VP.n15 161.3
R1423 VP.n28 VP.n0 161.3
R1424 VP.n27 VP.n26 161.3
R1425 VP.n25 VP.n24 161.3
R1426 VP.n23 VP.n2 161.3
R1427 VP.n21 VP.n20 161.3
R1428 VP.n19 VP.n3 161.3
R1429 VP.n18 VP.n17 161.3
R1430 VP.n24 VP.n23 56.5617
R1431 VP.n10 VP.n9 56.5617
R1432 VP.n18 VP.n16 45.349
R1433 VP.n21 VP.n3 44.4521
R1434 VP.n28 VP.n27 44.4521
R1435 VP.n14 VP.n13 44.4521
R1436 VP.n7 VP.n6 42.6379
R1437 VP.n8 VP.n7 36.5632
R1438 VP.n17 VP.n3 18.2581
R1439 VP.n29 VP.n28 18.2581
R1440 VP.n15 VP.n14 18.2581
R1441 VP.n23 VP.n22 17.4607
R1442 VP.n24 VP.n1 17.4607
R1443 VP.n10 VP.n5 17.4607
R1444 VP.n9 VP.n8 17.4607
R1445 VP.n22 VP.n21 7.13213
R1446 VP.n27 VP.n1 7.13213
R1447 VP.n13 VP.n5 7.13213
R1448 VP.n11 VP.n6 0.189894
R1449 VP.n12 VP.n11 0.189894
R1450 VP.n12 VP.n4 0.189894
R1451 VP.n16 VP.n4 0.189894
R1452 VP.n19 VP.n18 0.189894
R1453 VP.n20 VP.n19 0.189894
R1454 VP.n20 VP.n2 0.189894
R1455 VP.n25 VP.n2 0.189894
R1456 VP.n26 VP.n25 0.189894
R1457 VP.n26 VP.n0 0.189894
R1458 VP.n30 VP.n0 0.189894
R1459 VP VP.n30 0.0516364
R1460 VTAIL.n14 VTAIL.t7 43.5677
R1461 VTAIL.n11 VTAIL.t12 43.5677
R1462 VTAIL.n10 VTAIL.t4 43.5677
R1463 VTAIL.n7 VTAIL.t5 43.5677
R1464 VTAIL.n15 VTAIL.t3 43.5675
R1465 VTAIL.n2 VTAIL.t2 43.5675
R1466 VTAIL.n3 VTAIL.t10 43.5675
R1467 VTAIL.n6 VTAIL.t11 43.5675
R1468 VTAIL.n13 VTAIL.n12 42.2685
R1469 VTAIL.n9 VTAIL.n8 42.2685
R1470 VTAIL.n1 VTAIL.n0 42.2683
R1471 VTAIL.n5 VTAIL.n4 42.2683
R1472 VTAIL.n15 VTAIL.n14 26.5479
R1473 VTAIL.n7 VTAIL.n6 26.5479
R1474 VTAIL.n0 VTAIL.t1 1.29971
R1475 VTAIL.n0 VTAIL.t14 1.29971
R1476 VTAIL.n4 VTAIL.t8 1.29971
R1477 VTAIL.n4 VTAIL.t13 1.29971
R1478 VTAIL.n12 VTAIL.t9 1.29971
R1479 VTAIL.n12 VTAIL.t6 1.29971
R1480 VTAIL.n8 VTAIL.t0 1.29971
R1481 VTAIL.n8 VTAIL.t15 1.29971
R1482 VTAIL.n9 VTAIL.n7 1.0436
R1483 VTAIL.n10 VTAIL.n9 1.0436
R1484 VTAIL.n13 VTAIL.n11 1.0436
R1485 VTAIL.n14 VTAIL.n13 1.0436
R1486 VTAIL.n6 VTAIL.n5 1.0436
R1487 VTAIL.n5 VTAIL.n3 1.0436
R1488 VTAIL.n2 VTAIL.n1 1.0436
R1489 VTAIL VTAIL.n15 0.985414
R1490 VTAIL.n11 VTAIL.n10 0.470328
R1491 VTAIL.n3 VTAIL.n2 0.470328
R1492 VTAIL VTAIL.n1 0.0586897
R1493 VDD1 VDD1.n0 59.527
R1494 VDD1.n3 VDD1.n2 59.4133
R1495 VDD1.n3 VDD1.n1 59.4133
R1496 VDD1.n5 VDD1.n4 58.9473
R1497 VDD1.n5 VDD1.n3 42.1302
R1498 VDD1.n4 VDD1.t6 1.29971
R1499 VDD1.n4 VDD1.t7 1.29971
R1500 VDD1.n0 VDD1.t1 1.29971
R1501 VDD1.n0 VDD1.t4 1.29971
R1502 VDD1.n2 VDD1.t0 1.29971
R1503 VDD1.n2 VDD1.t3 1.29971
R1504 VDD1.n1 VDD1.t2 1.29971
R1505 VDD1.n1 VDD1.t5 1.29971
R1506 VDD1 VDD1.n5 0.463862
R1507 VN.n3 VN.t6 484.625
R1508 VN.n16 VN.t5 484.625
R1509 VN.n11 VN.t4 462.009
R1510 VN.n24 VN.t0 462.009
R1511 VN.n4 VN.t7 417.368
R1512 VN.n1 VN.t1 417.368
R1513 VN.n17 VN.t2 417.368
R1514 VN.n14 VN.t3 417.368
R1515 VN.n12 VN.n11 161.3
R1516 VN.n25 VN.n24 161.3
R1517 VN.n23 VN.n13 161.3
R1518 VN.n22 VN.n21 161.3
R1519 VN.n20 VN.n19 161.3
R1520 VN.n18 VN.n15 161.3
R1521 VN.n10 VN.n0 161.3
R1522 VN.n9 VN.n8 161.3
R1523 VN.n7 VN.n6 161.3
R1524 VN.n5 VN.n2 161.3
R1525 VN.n6 VN.n5 56.5617
R1526 VN.n19 VN.n18 56.5617
R1527 VN VN.n25 45.7297
R1528 VN.n10 VN.n9 44.4521
R1529 VN.n23 VN.n22 44.4521
R1530 VN.n16 VN.n15 42.6379
R1531 VN.n3 VN.n2 42.6379
R1532 VN.n4 VN.n3 36.5632
R1533 VN.n17 VN.n16 36.5632
R1534 VN.n11 VN.n10 18.2581
R1535 VN.n24 VN.n23 18.2581
R1536 VN.n5 VN.n4 17.4607
R1537 VN.n6 VN.n1 17.4607
R1538 VN.n18 VN.n17 17.4607
R1539 VN.n19 VN.n14 17.4607
R1540 VN.n9 VN.n1 7.13213
R1541 VN.n22 VN.n14 7.13213
R1542 VN.n25 VN.n13 0.189894
R1543 VN.n21 VN.n13 0.189894
R1544 VN.n21 VN.n20 0.189894
R1545 VN.n20 VN.n15 0.189894
R1546 VN.n7 VN.n2 0.189894
R1547 VN.n8 VN.n7 0.189894
R1548 VN.n8 VN.n0 0.189894
R1549 VN.n12 VN.n0 0.189894
R1550 VN VN.n12 0.0516364
R1551 VDD2.n2 VDD2.n1 59.4133
R1552 VDD2.n2 VDD2.n0 59.4133
R1553 VDD2 VDD2.n5 59.4106
R1554 VDD2.n4 VDD2.n3 58.9473
R1555 VDD2.n4 VDD2.n2 41.5472
R1556 VDD2.n5 VDD2.t5 1.29971
R1557 VDD2.n5 VDD2.t2 1.29971
R1558 VDD2.n3 VDD2.t7 1.29971
R1559 VDD2.n3 VDD2.t4 1.29971
R1560 VDD2.n1 VDD2.t6 1.29971
R1561 VDD2.n1 VDD2.t3 1.29971
R1562 VDD2.n0 VDD2.t1 1.29971
R1563 VDD2.n0 VDD2.t0 1.29971
R1564 VDD2 VDD2.n4 0.580241
C0 VTAIL VDD2 12.1912f
C1 VDD1 VTAIL 12.1483f
C2 VTAIL VP 7.43562f
C3 VDD2 VN 7.72176f
C4 VDD1 VN 0.148541f
C5 VN VP 6.15328f
C6 VDD1 VDD2 0.912839f
C7 VDD2 VP 0.336567f
C8 VDD1 VP 7.90926f
C9 VTAIL VN 7.42151f
C10 VDD2 B 3.917942f
C11 VDD1 B 4.170049f
C12 VTAIL B 10.930953f
C13 VN B 9.55025f
C14 VP B 7.551198f
C15 VDD2.t1 B 0.318603f
C16 VDD2.t0 B 0.318603f
C17 VDD2.n0 B 2.87514f
C18 VDD2.t6 B 0.318603f
C19 VDD2.t3 B 0.318603f
C20 VDD2.n1 B 2.87514f
C21 VDD2.n2 B 2.63914f
C22 VDD2.t7 B 0.318603f
C23 VDD2.t4 B 0.318603f
C24 VDD2.n3 B 2.87226f
C25 VDD2.n4 B 2.76264f
C26 VDD2.t5 B 0.318603f
C27 VDD2.t2 B 0.318603f
C28 VDD2.n5 B 2.87511f
C29 VN.n0 B 0.039942f
C30 VN.t1 B 1.46838f
C31 VN.n1 B 0.536971f
C32 VN.n2 B 0.171452f
C33 VN.t7 B 1.46838f
C34 VN.t6 B 1.54939f
C35 VN.n3 B 0.578388f
C36 VN.n4 B 0.580387f
C37 VN.n5 B 0.047458f
C38 VN.n6 B 0.047458f
C39 VN.n7 B 0.039942f
C40 VN.n8 B 0.039942f
C41 VN.n9 B 0.051048f
C42 VN.n10 B 0.017753f
C43 VN.t4 B 1.5219f
C44 VN.n11 B 0.579612f
C45 VN.n12 B 0.030954f
C46 VN.n13 B 0.039942f
C47 VN.t3 B 1.46838f
C48 VN.n14 B 0.536971f
C49 VN.n15 B 0.171452f
C50 VN.t2 B 1.46838f
C51 VN.t5 B 1.54939f
C52 VN.n16 B 0.578388f
C53 VN.n17 B 0.580387f
C54 VN.n18 B 0.047458f
C55 VN.n19 B 0.047458f
C56 VN.n20 B 0.039942f
C57 VN.n21 B 0.039942f
C58 VN.n22 B 0.051048f
C59 VN.n23 B 0.017753f
C60 VN.t0 B 1.5219f
C61 VN.n24 B 0.579612f
C62 VN.n25 B 1.89375f
C63 VDD1.t1 B 0.318639f
C64 VDD1.t4 B 0.318639f
C65 VDD1.n0 B 2.87625f
C66 VDD1.t2 B 0.318639f
C67 VDD1.t5 B 0.318639f
C68 VDD1.n1 B 2.87547f
C69 VDD1.t0 B 0.318639f
C70 VDD1.t3 B 0.318639f
C71 VDD1.n2 B 2.87547f
C72 VDD1.n3 B 2.69556f
C73 VDD1.t6 B 0.318639f
C74 VDD1.t7 B 0.318639f
C75 VDD1.n4 B 2.87259f
C76 VDD1.n5 B 2.79464f
C77 VTAIL.t1 B 0.230219f
C78 VTAIL.t14 B 0.230219f
C79 VTAIL.n0 B 2.01228f
C80 VTAIL.n1 B 0.268784f
C81 VTAIL.t2 B 2.56828f
C82 VTAIL.n2 B 0.366011f
C83 VTAIL.t10 B 2.56828f
C84 VTAIL.n3 B 0.366011f
C85 VTAIL.t8 B 0.230219f
C86 VTAIL.t13 B 0.230219f
C87 VTAIL.n4 B 2.01228f
C88 VTAIL.n5 B 0.329452f
C89 VTAIL.t11 B 2.56828f
C90 VTAIL.n6 B 1.47025f
C91 VTAIL.t5 B 2.5683f
C92 VTAIL.n7 B 1.47024f
C93 VTAIL.t0 B 0.230219f
C94 VTAIL.t15 B 0.230219f
C95 VTAIL.n8 B 2.01229f
C96 VTAIL.n9 B 0.329446f
C97 VTAIL.t4 B 2.5683f
C98 VTAIL.n10 B 0.365996f
C99 VTAIL.t12 B 2.5683f
C100 VTAIL.n11 B 0.365996f
C101 VTAIL.t9 B 0.230219f
C102 VTAIL.t6 B 0.230219f
C103 VTAIL.n12 B 2.01229f
C104 VTAIL.n13 B 0.329446f
C105 VTAIL.t7 B 2.56829f
C106 VTAIL.n14 B 1.47024f
C107 VTAIL.t3 B 2.56828f
C108 VTAIL.n15 B 1.46667f
C109 VP.n0 B 0.040424f
C110 VP.t7 B 1.48608f
C111 VP.n1 B 0.543446f
C112 VP.n2 B 0.040424f
C113 VP.t2 B 1.48608f
C114 VP.n3 B 0.017968f
C115 VP.n4 B 0.040424f
C116 VP.t0 B 1.54025f
C117 VP.t1 B 1.48608f
C118 VP.n5 B 0.543446f
C119 VP.n6 B 0.173519f
C120 VP.t3 B 1.48608f
C121 VP.t6 B 1.56807f
C122 VP.n7 B 0.585362f
C123 VP.n8 B 0.587385f
C124 VP.n9 B 0.04803f
C125 VP.n10 B 0.04803f
C126 VP.n11 B 0.040424f
C127 VP.n12 B 0.040424f
C128 VP.n13 B 0.051664f
C129 VP.n14 B 0.017968f
C130 VP.n15 B 0.586601f
C131 VP.n16 B 1.89016f
C132 VP.t5 B 1.54025f
C133 VP.n17 B 0.586601f
C134 VP.n18 B 1.9223f
C135 VP.n19 B 0.040424f
C136 VP.n20 B 0.040424f
C137 VP.n21 B 0.051664f
C138 VP.n22 B 0.543446f
C139 VP.n23 B 0.04803f
C140 VP.n24 B 0.04803f
C141 VP.n25 B 0.040424f
C142 VP.n26 B 0.040424f
C143 VP.n27 B 0.051664f
C144 VP.n28 B 0.017968f
C145 VP.t4 B 1.54025f
C146 VP.n29 B 0.586601f
C147 VP.n30 B 0.031327f
.ends

