* NGSPICE file created from diff_pair_sample_0894.ext - technology: sky130A

.subckt diff_pair_sample_0894 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VP.t0 VDD1.t4 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=1.56915 ps=9.84 w=9.51 l=1.03
X1 VTAIL.t2 VN.t0 VDD2.t5 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=1.56915 ps=9.84 w=9.51 l=1.03
X2 B.t11 B.t9 B.t10 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=1.03
X3 VDD2.t4 VN.t1 VTAIL.t0 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=1.03
X4 VDD1.t3 VP.t1 VTAIL.t10 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=1.03
X5 VDD2.t3 VN.t2 VTAIL.t4 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=1.03
X6 VDD2.t2 VN.t3 VTAIL.t5 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=1.03
X7 B.t8 B.t6 B.t7 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=1.03
X8 B.t5 B.t3 B.t4 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=1.03
X9 VDD2.t1 VN.t4 VTAIL.t3 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=1.03
X10 VTAIL.t1 VN.t5 VDD2.t0 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=1.56915 ps=9.84 w=9.51 l=1.03
X11 VTAIL.t9 VP.t2 VDD1.t2 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=1.56915 ps=9.84 w=9.51 l=1.03
X12 VDD1.t5 VP.t3 VTAIL.t8 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=1.56915 ps=9.84 w=9.51 l=1.03
X13 B.t2 B.t0 B.t1 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=3.7089 pd=19.8 as=0 ps=0 w=9.51 l=1.03
X14 VDD1.t0 VP.t4 VTAIL.t7 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=1.03
X15 VDD1.t1 VP.t5 VTAIL.t6 w_n2058_n2870# sky130_fd_pr__pfet_01v8 ad=1.56915 pd=9.84 as=3.7089 ps=19.8 w=9.51 l=1.03
R0 VP.n3 VP.t3 283.488
R1 VP.n8 VP.t1 260.889
R2 VP.n14 VP.t4 260.889
R3 VP.n6 VP.t5 260.889
R4 VP.n12 VP.t2 222.517
R5 VP.n4 VP.t0 222.517
R6 VP.n5 VP.n2 161.3
R7 VP.n13 VP.n0 161.3
R8 VP.n12 VP.n11 161.3
R9 VP.n10 VP.n1 161.3
R10 VP.n7 VP.n6 80.6037
R11 VP.n15 VP.n14 80.6037
R12 VP.n9 VP.n8 80.6037
R13 VP.n8 VP.n1 48.9345
R14 VP.n14 VP.n13 48.9345
R15 VP.n6 VP.n5 48.9345
R16 VP.n9 VP.n7 40.7514
R17 VP.n4 VP.n3 32.2627
R18 VP.n3 VP.n2 28.3407
R19 VP.n12 VP.n1 24.4675
R20 VP.n13 VP.n12 24.4675
R21 VP.n5 VP.n4 24.4675
R22 VP.n7 VP.n2 0.285035
R23 VP.n10 VP.n9 0.285035
R24 VP.n15 VP.n0 0.285035
R25 VP.n11 VP.n10 0.189894
R26 VP.n11 VP.n0 0.189894
R27 VP VP.n15 0.146778
R28 VDD1.n46 VDD1.n0 756.745
R29 VDD1.n97 VDD1.n51 756.745
R30 VDD1.n47 VDD1.n46 585
R31 VDD1.n45 VDD1.n44 585
R32 VDD1.n4 VDD1.n3 585
R33 VDD1.n39 VDD1.n38 585
R34 VDD1.n37 VDD1.n36 585
R35 VDD1.n8 VDD1.n7 585
R36 VDD1.n31 VDD1.n30 585
R37 VDD1.n29 VDD1.n28 585
R38 VDD1.n12 VDD1.n11 585
R39 VDD1.n23 VDD1.n22 585
R40 VDD1.n21 VDD1.n20 585
R41 VDD1.n16 VDD1.n15 585
R42 VDD1.n67 VDD1.n66 585
R43 VDD1.n72 VDD1.n71 585
R44 VDD1.n74 VDD1.n73 585
R45 VDD1.n63 VDD1.n62 585
R46 VDD1.n80 VDD1.n79 585
R47 VDD1.n82 VDD1.n81 585
R48 VDD1.n59 VDD1.n58 585
R49 VDD1.n88 VDD1.n87 585
R50 VDD1.n90 VDD1.n89 585
R51 VDD1.n55 VDD1.n54 585
R52 VDD1.n96 VDD1.n95 585
R53 VDD1.n98 VDD1.n97 585
R54 VDD1.n17 VDD1.t5 327.467
R55 VDD1.n68 VDD1.t3 327.467
R56 VDD1.n46 VDD1.n45 171.744
R57 VDD1.n45 VDD1.n3 171.744
R58 VDD1.n38 VDD1.n3 171.744
R59 VDD1.n38 VDD1.n37 171.744
R60 VDD1.n37 VDD1.n7 171.744
R61 VDD1.n30 VDD1.n7 171.744
R62 VDD1.n30 VDD1.n29 171.744
R63 VDD1.n29 VDD1.n11 171.744
R64 VDD1.n22 VDD1.n11 171.744
R65 VDD1.n22 VDD1.n21 171.744
R66 VDD1.n21 VDD1.n15 171.744
R67 VDD1.n72 VDD1.n66 171.744
R68 VDD1.n73 VDD1.n72 171.744
R69 VDD1.n73 VDD1.n62 171.744
R70 VDD1.n80 VDD1.n62 171.744
R71 VDD1.n81 VDD1.n80 171.744
R72 VDD1.n81 VDD1.n58 171.744
R73 VDD1.n88 VDD1.n58 171.744
R74 VDD1.n89 VDD1.n88 171.744
R75 VDD1.n89 VDD1.n54 171.744
R76 VDD1.n96 VDD1.n54 171.744
R77 VDD1.n97 VDD1.n96 171.744
R78 VDD1.t5 VDD1.n15 85.8723
R79 VDD1.t3 VDD1.n66 85.8723
R80 VDD1.n103 VDD1.n102 77.4541
R81 VDD1.n105 VDD1.n104 77.2163
R82 VDD1 VDD1.n50 48.0562
R83 VDD1.n103 VDD1.n101 47.9427
R84 VDD1.n105 VDD1.n103 36.8931
R85 VDD1.n17 VDD1.n16 16.3895
R86 VDD1.n68 VDD1.n67 16.3895
R87 VDD1.n20 VDD1.n19 12.8005
R88 VDD1.n71 VDD1.n70 12.8005
R89 VDD1.n23 VDD1.n14 12.0247
R90 VDD1.n74 VDD1.n65 12.0247
R91 VDD1.n24 VDD1.n12 11.249
R92 VDD1.n75 VDD1.n63 11.249
R93 VDD1.n28 VDD1.n27 10.4732
R94 VDD1.n79 VDD1.n78 10.4732
R95 VDD1.n50 VDD1.n0 9.69747
R96 VDD1.n31 VDD1.n10 9.69747
R97 VDD1.n82 VDD1.n61 9.69747
R98 VDD1.n101 VDD1.n51 9.69747
R99 VDD1.n50 VDD1.n49 9.45567
R100 VDD1.n101 VDD1.n100 9.45567
R101 VDD1.n43 VDD1.n42 9.3005
R102 VDD1.n2 VDD1.n1 9.3005
R103 VDD1.n49 VDD1.n48 9.3005
R104 VDD1.n41 VDD1.n40 9.3005
R105 VDD1.n6 VDD1.n5 9.3005
R106 VDD1.n35 VDD1.n34 9.3005
R107 VDD1.n33 VDD1.n32 9.3005
R108 VDD1.n10 VDD1.n9 9.3005
R109 VDD1.n27 VDD1.n26 9.3005
R110 VDD1.n25 VDD1.n24 9.3005
R111 VDD1.n14 VDD1.n13 9.3005
R112 VDD1.n19 VDD1.n18 9.3005
R113 VDD1.n92 VDD1.n91 9.3005
R114 VDD1.n94 VDD1.n93 9.3005
R115 VDD1.n53 VDD1.n52 9.3005
R116 VDD1.n100 VDD1.n99 9.3005
R117 VDD1.n86 VDD1.n85 9.3005
R118 VDD1.n84 VDD1.n83 9.3005
R119 VDD1.n61 VDD1.n60 9.3005
R120 VDD1.n78 VDD1.n77 9.3005
R121 VDD1.n76 VDD1.n75 9.3005
R122 VDD1.n65 VDD1.n64 9.3005
R123 VDD1.n70 VDD1.n69 9.3005
R124 VDD1.n57 VDD1.n56 9.3005
R125 VDD1.n48 VDD1.n47 8.92171
R126 VDD1.n32 VDD1.n8 8.92171
R127 VDD1.n83 VDD1.n59 8.92171
R128 VDD1.n99 VDD1.n98 8.92171
R129 VDD1.n44 VDD1.n2 8.14595
R130 VDD1.n36 VDD1.n35 8.14595
R131 VDD1.n87 VDD1.n86 8.14595
R132 VDD1.n95 VDD1.n53 8.14595
R133 VDD1.n43 VDD1.n4 7.3702
R134 VDD1.n39 VDD1.n6 7.3702
R135 VDD1.n90 VDD1.n57 7.3702
R136 VDD1.n94 VDD1.n55 7.3702
R137 VDD1.n40 VDD1.n4 6.59444
R138 VDD1.n40 VDD1.n39 6.59444
R139 VDD1.n91 VDD1.n90 6.59444
R140 VDD1.n91 VDD1.n55 6.59444
R141 VDD1.n44 VDD1.n43 5.81868
R142 VDD1.n36 VDD1.n6 5.81868
R143 VDD1.n87 VDD1.n57 5.81868
R144 VDD1.n95 VDD1.n94 5.81868
R145 VDD1.n47 VDD1.n2 5.04292
R146 VDD1.n35 VDD1.n8 5.04292
R147 VDD1.n86 VDD1.n59 5.04292
R148 VDD1.n98 VDD1.n53 5.04292
R149 VDD1.n48 VDD1.n0 4.26717
R150 VDD1.n32 VDD1.n31 4.26717
R151 VDD1.n83 VDD1.n82 4.26717
R152 VDD1.n99 VDD1.n51 4.26717
R153 VDD1.n18 VDD1.n17 3.70984
R154 VDD1.n69 VDD1.n68 3.70984
R155 VDD1.n28 VDD1.n10 3.49141
R156 VDD1.n79 VDD1.n61 3.49141
R157 VDD1.n104 VDD1.t4 3.41848
R158 VDD1.n104 VDD1.t1 3.41848
R159 VDD1.n102 VDD1.t2 3.41848
R160 VDD1.n102 VDD1.t0 3.41848
R161 VDD1.n27 VDD1.n12 2.71565
R162 VDD1.n78 VDD1.n63 2.71565
R163 VDD1.n24 VDD1.n23 1.93989
R164 VDD1.n75 VDD1.n74 1.93989
R165 VDD1.n20 VDD1.n14 1.16414
R166 VDD1.n71 VDD1.n65 1.16414
R167 VDD1.n19 VDD1.n16 0.388379
R168 VDD1.n70 VDD1.n67 0.388379
R169 VDD1 VDD1.n105 0.235414
R170 VDD1.n49 VDD1.n1 0.155672
R171 VDD1.n42 VDD1.n1 0.155672
R172 VDD1.n42 VDD1.n41 0.155672
R173 VDD1.n41 VDD1.n5 0.155672
R174 VDD1.n34 VDD1.n5 0.155672
R175 VDD1.n34 VDD1.n33 0.155672
R176 VDD1.n33 VDD1.n9 0.155672
R177 VDD1.n26 VDD1.n9 0.155672
R178 VDD1.n26 VDD1.n25 0.155672
R179 VDD1.n25 VDD1.n13 0.155672
R180 VDD1.n18 VDD1.n13 0.155672
R181 VDD1.n69 VDD1.n64 0.155672
R182 VDD1.n76 VDD1.n64 0.155672
R183 VDD1.n77 VDD1.n76 0.155672
R184 VDD1.n77 VDD1.n60 0.155672
R185 VDD1.n84 VDD1.n60 0.155672
R186 VDD1.n85 VDD1.n84 0.155672
R187 VDD1.n85 VDD1.n56 0.155672
R188 VDD1.n92 VDD1.n56 0.155672
R189 VDD1.n93 VDD1.n92 0.155672
R190 VDD1.n93 VDD1.n52 0.155672
R191 VDD1.n100 VDD1.n52 0.155672
R192 VTAIL.n210 VTAIL.n164 756.745
R193 VTAIL.n48 VTAIL.n2 756.745
R194 VTAIL.n158 VTAIL.n112 756.745
R195 VTAIL.n104 VTAIL.n58 756.745
R196 VTAIL.n180 VTAIL.n179 585
R197 VTAIL.n185 VTAIL.n184 585
R198 VTAIL.n187 VTAIL.n186 585
R199 VTAIL.n176 VTAIL.n175 585
R200 VTAIL.n193 VTAIL.n192 585
R201 VTAIL.n195 VTAIL.n194 585
R202 VTAIL.n172 VTAIL.n171 585
R203 VTAIL.n201 VTAIL.n200 585
R204 VTAIL.n203 VTAIL.n202 585
R205 VTAIL.n168 VTAIL.n167 585
R206 VTAIL.n209 VTAIL.n208 585
R207 VTAIL.n211 VTAIL.n210 585
R208 VTAIL.n18 VTAIL.n17 585
R209 VTAIL.n23 VTAIL.n22 585
R210 VTAIL.n25 VTAIL.n24 585
R211 VTAIL.n14 VTAIL.n13 585
R212 VTAIL.n31 VTAIL.n30 585
R213 VTAIL.n33 VTAIL.n32 585
R214 VTAIL.n10 VTAIL.n9 585
R215 VTAIL.n39 VTAIL.n38 585
R216 VTAIL.n41 VTAIL.n40 585
R217 VTAIL.n6 VTAIL.n5 585
R218 VTAIL.n47 VTAIL.n46 585
R219 VTAIL.n49 VTAIL.n48 585
R220 VTAIL.n159 VTAIL.n158 585
R221 VTAIL.n157 VTAIL.n156 585
R222 VTAIL.n116 VTAIL.n115 585
R223 VTAIL.n151 VTAIL.n150 585
R224 VTAIL.n149 VTAIL.n148 585
R225 VTAIL.n120 VTAIL.n119 585
R226 VTAIL.n143 VTAIL.n142 585
R227 VTAIL.n141 VTAIL.n140 585
R228 VTAIL.n124 VTAIL.n123 585
R229 VTAIL.n135 VTAIL.n134 585
R230 VTAIL.n133 VTAIL.n132 585
R231 VTAIL.n128 VTAIL.n127 585
R232 VTAIL.n105 VTAIL.n104 585
R233 VTAIL.n103 VTAIL.n102 585
R234 VTAIL.n62 VTAIL.n61 585
R235 VTAIL.n97 VTAIL.n96 585
R236 VTAIL.n95 VTAIL.n94 585
R237 VTAIL.n66 VTAIL.n65 585
R238 VTAIL.n89 VTAIL.n88 585
R239 VTAIL.n87 VTAIL.n86 585
R240 VTAIL.n70 VTAIL.n69 585
R241 VTAIL.n81 VTAIL.n80 585
R242 VTAIL.n79 VTAIL.n78 585
R243 VTAIL.n74 VTAIL.n73 585
R244 VTAIL.n181 VTAIL.t4 327.467
R245 VTAIL.n19 VTAIL.t7 327.467
R246 VTAIL.n75 VTAIL.t5 327.467
R247 VTAIL.n129 VTAIL.t6 327.467
R248 VTAIL.n185 VTAIL.n179 171.744
R249 VTAIL.n186 VTAIL.n185 171.744
R250 VTAIL.n186 VTAIL.n175 171.744
R251 VTAIL.n193 VTAIL.n175 171.744
R252 VTAIL.n194 VTAIL.n193 171.744
R253 VTAIL.n194 VTAIL.n171 171.744
R254 VTAIL.n201 VTAIL.n171 171.744
R255 VTAIL.n202 VTAIL.n201 171.744
R256 VTAIL.n202 VTAIL.n167 171.744
R257 VTAIL.n209 VTAIL.n167 171.744
R258 VTAIL.n210 VTAIL.n209 171.744
R259 VTAIL.n23 VTAIL.n17 171.744
R260 VTAIL.n24 VTAIL.n23 171.744
R261 VTAIL.n24 VTAIL.n13 171.744
R262 VTAIL.n31 VTAIL.n13 171.744
R263 VTAIL.n32 VTAIL.n31 171.744
R264 VTAIL.n32 VTAIL.n9 171.744
R265 VTAIL.n39 VTAIL.n9 171.744
R266 VTAIL.n40 VTAIL.n39 171.744
R267 VTAIL.n40 VTAIL.n5 171.744
R268 VTAIL.n47 VTAIL.n5 171.744
R269 VTAIL.n48 VTAIL.n47 171.744
R270 VTAIL.n158 VTAIL.n157 171.744
R271 VTAIL.n157 VTAIL.n115 171.744
R272 VTAIL.n150 VTAIL.n115 171.744
R273 VTAIL.n150 VTAIL.n149 171.744
R274 VTAIL.n149 VTAIL.n119 171.744
R275 VTAIL.n142 VTAIL.n119 171.744
R276 VTAIL.n142 VTAIL.n141 171.744
R277 VTAIL.n141 VTAIL.n123 171.744
R278 VTAIL.n134 VTAIL.n123 171.744
R279 VTAIL.n134 VTAIL.n133 171.744
R280 VTAIL.n133 VTAIL.n127 171.744
R281 VTAIL.n104 VTAIL.n103 171.744
R282 VTAIL.n103 VTAIL.n61 171.744
R283 VTAIL.n96 VTAIL.n61 171.744
R284 VTAIL.n96 VTAIL.n95 171.744
R285 VTAIL.n95 VTAIL.n65 171.744
R286 VTAIL.n88 VTAIL.n65 171.744
R287 VTAIL.n88 VTAIL.n87 171.744
R288 VTAIL.n87 VTAIL.n69 171.744
R289 VTAIL.n80 VTAIL.n69 171.744
R290 VTAIL.n80 VTAIL.n79 171.744
R291 VTAIL.n79 VTAIL.n73 171.744
R292 VTAIL.t4 VTAIL.n179 85.8723
R293 VTAIL.t7 VTAIL.n17 85.8723
R294 VTAIL.t6 VTAIL.n127 85.8723
R295 VTAIL.t5 VTAIL.n73 85.8723
R296 VTAIL.n1 VTAIL.n0 60.5375
R297 VTAIL.n55 VTAIL.n54 60.5375
R298 VTAIL.n111 VTAIL.n110 60.5375
R299 VTAIL.n57 VTAIL.n56 60.5375
R300 VTAIL.n215 VTAIL.n214 30.4399
R301 VTAIL.n53 VTAIL.n52 30.4399
R302 VTAIL.n163 VTAIL.n162 30.4399
R303 VTAIL.n109 VTAIL.n108 30.4399
R304 VTAIL.n57 VTAIL.n55 22.91
R305 VTAIL.n215 VTAIL.n163 21.7376
R306 VTAIL.n181 VTAIL.n180 16.3895
R307 VTAIL.n19 VTAIL.n18 16.3895
R308 VTAIL.n129 VTAIL.n128 16.3895
R309 VTAIL.n75 VTAIL.n74 16.3895
R310 VTAIL.n184 VTAIL.n183 12.8005
R311 VTAIL.n22 VTAIL.n21 12.8005
R312 VTAIL.n132 VTAIL.n131 12.8005
R313 VTAIL.n78 VTAIL.n77 12.8005
R314 VTAIL.n187 VTAIL.n178 12.0247
R315 VTAIL.n25 VTAIL.n16 12.0247
R316 VTAIL.n135 VTAIL.n126 12.0247
R317 VTAIL.n81 VTAIL.n72 12.0247
R318 VTAIL.n188 VTAIL.n176 11.249
R319 VTAIL.n26 VTAIL.n14 11.249
R320 VTAIL.n136 VTAIL.n124 11.249
R321 VTAIL.n82 VTAIL.n70 11.249
R322 VTAIL.n192 VTAIL.n191 10.4732
R323 VTAIL.n30 VTAIL.n29 10.4732
R324 VTAIL.n140 VTAIL.n139 10.4732
R325 VTAIL.n86 VTAIL.n85 10.4732
R326 VTAIL.n195 VTAIL.n174 9.69747
R327 VTAIL.n214 VTAIL.n164 9.69747
R328 VTAIL.n33 VTAIL.n12 9.69747
R329 VTAIL.n52 VTAIL.n2 9.69747
R330 VTAIL.n162 VTAIL.n112 9.69747
R331 VTAIL.n143 VTAIL.n122 9.69747
R332 VTAIL.n108 VTAIL.n58 9.69747
R333 VTAIL.n89 VTAIL.n68 9.69747
R334 VTAIL.n214 VTAIL.n213 9.45567
R335 VTAIL.n52 VTAIL.n51 9.45567
R336 VTAIL.n162 VTAIL.n161 9.45567
R337 VTAIL.n108 VTAIL.n107 9.45567
R338 VTAIL.n205 VTAIL.n204 9.3005
R339 VTAIL.n207 VTAIL.n206 9.3005
R340 VTAIL.n166 VTAIL.n165 9.3005
R341 VTAIL.n213 VTAIL.n212 9.3005
R342 VTAIL.n199 VTAIL.n198 9.3005
R343 VTAIL.n197 VTAIL.n196 9.3005
R344 VTAIL.n174 VTAIL.n173 9.3005
R345 VTAIL.n191 VTAIL.n190 9.3005
R346 VTAIL.n189 VTAIL.n188 9.3005
R347 VTAIL.n178 VTAIL.n177 9.3005
R348 VTAIL.n183 VTAIL.n182 9.3005
R349 VTAIL.n170 VTAIL.n169 9.3005
R350 VTAIL.n43 VTAIL.n42 9.3005
R351 VTAIL.n45 VTAIL.n44 9.3005
R352 VTAIL.n4 VTAIL.n3 9.3005
R353 VTAIL.n51 VTAIL.n50 9.3005
R354 VTAIL.n37 VTAIL.n36 9.3005
R355 VTAIL.n35 VTAIL.n34 9.3005
R356 VTAIL.n12 VTAIL.n11 9.3005
R357 VTAIL.n29 VTAIL.n28 9.3005
R358 VTAIL.n27 VTAIL.n26 9.3005
R359 VTAIL.n16 VTAIL.n15 9.3005
R360 VTAIL.n21 VTAIL.n20 9.3005
R361 VTAIL.n8 VTAIL.n7 9.3005
R362 VTAIL.n114 VTAIL.n113 9.3005
R363 VTAIL.n155 VTAIL.n154 9.3005
R364 VTAIL.n153 VTAIL.n152 9.3005
R365 VTAIL.n118 VTAIL.n117 9.3005
R366 VTAIL.n147 VTAIL.n146 9.3005
R367 VTAIL.n145 VTAIL.n144 9.3005
R368 VTAIL.n122 VTAIL.n121 9.3005
R369 VTAIL.n139 VTAIL.n138 9.3005
R370 VTAIL.n137 VTAIL.n136 9.3005
R371 VTAIL.n126 VTAIL.n125 9.3005
R372 VTAIL.n131 VTAIL.n130 9.3005
R373 VTAIL.n161 VTAIL.n160 9.3005
R374 VTAIL.n101 VTAIL.n100 9.3005
R375 VTAIL.n60 VTAIL.n59 9.3005
R376 VTAIL.n107 VTAIL.n106 9.3005
R377 VTAIL.n99 VTAIL.n98 9.3005
R378 VTAIL.n64 VTAIL.n63 9.3005
R379 VTAIL.n93 VTAIL.n92 9.3005
R380 VTAIL.n91 VTAIL.n90 9.3005
R381 VTAIL.n68 VTAIL.n67 9.3005
R382 VTAIL.n85 VTAIL.n84 9.3005
R383 VTAIL.n83 VTAIL.n82 9.3005
R384 VTAIL.n72 VTAIL.n71 9.3005
R385 VTAIL.n77 VTAIL.n76 9.3005
R386 VTAIL.n196 VTAIL.n172 8.92171
R387 VTAIL.n212 VTAIL.n211 8.92171
R388 VTAIL.n34 VTAIL.n10 8.92171
R389 VTAIL.n50 VTAIL.n49 8.92171
R390 VTAIL.n160 VTAIL.n159 8.92171
R391 VTAIL.n144 VTAIL.n120 8.92171
R392 VTAIL.n106 VTAIL.n105 8.92171
R393 VTAIL.n90 VTAIL.n66 8.92171
R394 VTAIL.n200 VTAIL.n199 8.14595
R395 VTAIL.n208 VTAIL.n166 8.14595
R396 VTAIL.n38 VTAIL.n37 8.14595
R397 VTAIL.n46 VTAIL.n4 8.14595
R398 VTAIL.n156 VTAIL.n114 8.14595
R399 VTAIL.n148 VTAIL.n147 8.14595
R400 VTAIL.n102 VTAIL.n60 8.14595
R401 VTAIL.n94 VTAIL.n93 8.14595
R402 VTAIL.n203 VTAIL.n170 7.3702
R403 VTAIL.n207 VTAIL.n168 7.3702
R404 VTAIL.n41 VTAIL.n8 7.3702
R405 VTAIL.n45 VTAIL.n6 7.3702
R406 VTAIL.n155 VTAIL.n116 7.3702
R407 VTAIL.n151 VTAIL.n118 7.3702
R408 VTAIL.n101 VTAIL.n62 7.3702
R409 VTAIL.n97 VTAIL.n64 7.3702
R410 VTAIL.n204 VTAIL.n203 6.59444
R411 VTAIL.n204 VTAIL.n168 6.59444
R412 VTAIL.n42 VTAIL.n41 6.59444
R413 VTAIL.n42 VTAIL.n6 6.59444
R414 VTAIL.n152 VTAIL.n116 6.59444
R415 VTAIL.n152 VTAIL.n151 6.59444
R416 VTAIL.n98 VTAIL.n62 6.59444
R417 VTAIL.n98 VTAIL.n97 6.59444
R418 VTAIL.n200 VTAIL.n170 5.81868
R419 VTAIL.n208 VTAIL.n207 5.81868
R420 VTAIL.n38 VTAIL.n8 5.81868
R421 VTAIL.n46 VTAIL.n45 5.81868
R422 VTAIL.n156 VTAIL.n155 5.81868
R423 VTAIL.n148 VTAIL.n118 5.81868
R424 VTAIL.n102 VTAIL.n101 5.81868
R425 VTAIL.n94 VTAIL.n64 5.81868
R426 VTAIL.n199 VTAIL.n172 5.04292
R427 VTAIL.n211 VTAIL.n166 5.04292
R428 VTAIL.n37 VTAIL.n10 5.04292
R429 VTAIL.n49 VTAIL.n4 5.04292
R430 VTAIL.n159 VTAIL.n114 5.04292
R431 VTAIL.n147 VTAIL.n120 5.04292
R432 VTAIL.n105 VTAIL.n60 5.04292
R433 VTAIL.n93 VTAIL.n66 5.04292
R434 VTAIL.n196 VTAIL.n195 4.26717
R435 VTAIL.n212 VTAIL.n164 4.26717
R436 VTAIL.n34 VTAIL.n33 4.26717
R437 VTAIL.n50 VTAIL.n2 4.26717
R438 VTAIL.n160 VTAIL.n112 4.26717
R439 VTAIL.n144 VTAIL.n143 4.26717
R440 VTAIL.n106 VTAIL.n58 4.26717
R441 VTAIL.n90 VTAIL.n89 4.26717
R442 VTAIL.n182 VTAIL.n181 3.70984
R443 VTAIL.n20 VTAIL.n19 3.70984
R444 VTAIL.n76 VTAIL.n75 3.70984
R445 VTAIL.n130 VTAIL.n129 3.70984
R446 VTAIL.n192 VTAIL.n174 3.49141
R447 VTAIL.n30 VTAIL.n12 3.49141
R448 VTAIL.n140 VTAIL.n122 3.49141
R449 VTAIL.n86 VTAIL.n68 3.49141
R450 VTAIL.n0 VTAIL.t0 3.41848
R451 VTAIL.n0 VTAIL.t2 3.41848
R452 VTAIL.n54 VTAIL.t10 3.41848
R453 VTAIL.n54 VTAIL.t9 3.41848
R454 VTAIL.n110 VTAIL.t8 3.41848
R455 VTAIL.n110 VTAIL.t11 3.41848
R456 VTAIL.n56 VTAIL.t3 3.41848
R457 VTAIL.n56 VTAIL.t1 3.41848
R458 VTAIL.n191 VTAIL.n176 2.71565
R459 VTAIL.n29 VTAIL.n14 2.71565
R460 VTAIL.n139 VTAIL.n124 2.71565
R461 VTAIL.n85 VTAIL.n70 2.71565
R462 VTAIL.n188 VTAIL.n187 1.93989
R463 VTAIL.n26 VTAIL.n25 1.93989
R464 VTAIL.n136 VTAIL.n135 1.93989
R465 VTAIL.n82 VTAIL.n81 1.93989
R466 VTAIL.n109 VTAIL.n57 1.17291
R467 VTAIL.n163 VTAIL.n111 1.17291
R468 VTAIL.n55 VTAIL.n53 1.17291
R469 VTAIL.n184 VTAIL.n178 1.16414
R470 VTAIL.n22 VTAIL.n16 1.16414
R471 VTAIL.n132 VTAIL.n126 1.16414
R472 VTAIL.n78 VTAIL.n72 1.16414
R473 VTAIL.n111 VTAIL.n109 1.05653
R474 VTAIL.n53 VTAIL.n1 1.05653
R475 VTAIL VTAIL.n215 0.821621
R476 VTAIL.n183 VTAIL.n180 0.388379
R477 VTAIL.n21 VTAIL.n18 0.388379
R478 VTAIL.n131 VTAIL.n128 0.388379
R479 VTAIL.n77 VTAIL.n74 0.388379
R480 VTAIL VTAIL.n1 0.351793
R481 VTAIL.n182 VTAIL.n177 0.155672
R482 VTAIL.n189 VTAIL.n177 0.155672
R483 VTAIL.n190 VTAIL.n189 0.155672
R484 VTAIL.n190 VTAIL.n173 0.155672
R485 VTAIL.n197 VTAIL.n173 0.155672
R486 VTAIL.n198 VTAIL.n197 0.155672
R487 VTAIL.n198 VTAIL.n169 0.155672
R488 VTAIL.n205 VTAIL.n169 0.155672
R489 VTAIL.n206 VTAIL.n205 0.155672
R490 VTAIL.n206 VTAIL.n165 0.155672
R491 VTAIL.n213 VTAIL.n165 0.155672
R492 VTAIL.n20 VTAIL.n15 0.155672
R493 VTAIL.n27 VTAIL.n15 0.155672
R494 VTAIL.n28 VTAIL.n27 0.155672
R495 VTAIL.n28 VTAIL.n11 0.155672
R496 VTAIL.n35 VTAIL.n11 0.155672
R497 VTAIL.n36 VTAIL.n35 0.155672
R498 VTAIL.n36 VTAIL.n7 0.155672
R499 VTAIL.n43 VTAIL.n7 0.155672
R500 VTAIL.n44 VTAIL.n43 0.155672
R501 VTAIL.n44 VTAIL.n3 0.155672
R502 VTAIL.n51 VTAIL.n3 0.155672
R503 VTAIL.n161 VTAIL.n113 0.155672
R504 VTAIL.n154 VTAIL.n113 0.155672
R505 VTAIL.n154 VTAIL.n153 0.155672
R506 VTAIL.n153 VTAIL.n117 0.155672
R507 VTAIL.n146 VTAIL.n117 0.155672
R508 VTAIL.n146 VTAIL.n145 0.155672
R509 VTAIL.n145 VTAIL.n121 0.155672
R510 VTAIL.n138 VTAIL.n121 0.155672
R511 VTAIL.n138 VTAIL.n137 0.155672
R512 VTAIL.n137 VTAIL.n125 0.155672
R513 VTAIL.n130 VTAIL.n125 0.155672
R514 VTAIL.n107 VTAIL.n59 0.155672
R515 VTAIL.n100 VTAIL.n59 0.155672
R516 VTAIL.n100 VTAIL.n99 0.155672
R517 VTAIL.n99 VTAIL.n63 0.155672
R518 VTAIL.n92 VTAIL.n63 0.155672
R519 VTAIL.n92 VTAIL.n91 0.155672
R520 VTAIL.n91 VTAIL.n67 0.155672
R521 VTAIL.n84 VTAIL.n67 0.155672
R522 VTAIL.n84 VTAIL.n83 0.155672
R523 VTAIL.n83 VTAIL.n71 0.155672
R524 VTAIL.n76 VTAIL.n71 0.155672
R525 VN.n1 VN.t1 283.488
R526 VN.n7 VN.t3 283.488
R527 VN.n4 VN.t2 260.889
R528 VN.n10 VN.t4 260.889
R529 VN.n2 VN.t0 222.517
R530 VN.n8 VN.t5 222.517
R531 VN.n9 VN.n6 161.3
R532 VN.n3 VN.n0 161.3
R533 VN.n11 VN.n10 80.6037
R534 VN.n5 VN.n4 80.6037
R535 VN.n4 VN.n3 48.9345
R536 VN.n10 VN.n9 48.9345
R537 VN VN.n11 41.0369
R538 VN.n2 VN.n1 32.2627
R539 VN.n8 VN.n7 32.2627
R540 VN.n7 VN.n6 28.3407
R541 VN.n1 VN.n0 28.3407
R542 VN.n3 VN.n2 24.4675
R543 VN.n9 VN.n8 24.4675
R544 VN.n11 VN.n6 0.285035
R545 VN.n5 VN.n0 0.285035
R546 VN VN.n5 0.146778
R547 VDD2.n99 VDD2.n53 756.745
R548 VDD2.n46 VDD2.n0 756.745
R549 VDD2.n100 VDD2.n99 585
R550 VDD2.n98 VDD2.n97 585
R551 VDD2.n57 VDD2.n56 585
R552 VDD2.n92 VDD2.n91 585
R553 VDD2.n90 VDD2.n89 585
R554 VDD2.n61 VDD2.n60 585
R555 VDD2.n84 VDD2.n83 585
R556 VDD2.n82 VDD2.n81 585
R557 VDD2.n65 VDD2.n64 585
R558 VDD2.n76 VDD2.n75 585
R559 VDD2.n74 VDD2.n73 585
R560 VDD2.n69 VDD2.n68 585
R561 VDD2.n16 VDD2.n15 585
R562 VDD2.n21 VDD2.n20 585
R563 VDD2.n23 VDD2.n22 585
R564 VDD2.n12 VDD2.n11 585
R565 VDD2.n29 VDD2.n28 585
R566 VDD2.n31 VDD2.n30 585
R567 VDD2.n8 VDD2.n7 585
R568 VDD2.n37 VDD2.n36 585
R569 VDD2.n39 VDD2.n38 585
R570 VDD2.n4 VDD2.n3 585
R571 VDD2.n45 VDD2.n44 585
R572 VDD2.n47 VDD2.n46 585
R573 VDD2.n70 VDD2.t1 327.467
R574 VDD2.n17 VDD2.t4 327.467
R575 VDD2.n99 VDD2.n98 171.744
R576 VDD2.n98 VDD2.n56 171.744
R577 VDD2.n91 VDD2.n56 171.744
R578 VDD2.n91 VDD2.n90 171.744
R579 VDD2.n90 VDD2.n60 171.744
R580 VDD2.n83 VDD2.n60 171.744
R581 VDD2.n83 VDD2.n82 171.744
R582 VDD2.n82 VDD2.n64 171.744
R583 VDD2.n75 VDD2.n64 171.744
R584 VDD2.n75 VDD2.n74 171.744
R585 VDD2.n74 VDD2.n68 171.744
R586 VDD2.n21 VDD2.n15 171.744
R587 VDD2.n22 VDD2.n21 171.744
R588 VDD2.n22 VDD2.n11 171.744
R589 VDD2.n29 VDD2.n11 171.744
R590 VDD2.n30 VDD2.n29 171.744
R591 VDD2.n30 VDD2.n7 171.744
R592 VDD2.n37 VDD2.n7 171.744
R593 VDD2.n38 VDD2.n37 171.744
R594 VDD2.n38 VDD2.n3 171.744
R595 VDD2.n45 VDD2.n3 171.744
R596 VDD2.n46 VDD2.n45 171.744
R597 VDD2.t1 VDD2.n68 85.8723
R598 VDD2.t4 VDD2.n15 85.8723
R599 VDD2.n52 VDD2.n51 77.4541
R600 VDD2 VDD2.n105 77.4512
R601 VDD2.n52 VDD2.n50 47.9427
R602 VDD2.n104 VDD2.n103 47.1187
R603 VDD2.n104 VDD2.n52 35.7239
R604 VDD2.n70 VDD2.n69 16.3895
R605 VDD2.n17 VDD2.n16 16.3895
R606 VDD2.n73 VDD2.n72 12.8005
R607 VDD2.n20 VDD2.n19 12.8005
R608 VDD2.n76 VDD2.n67 12.0247
R609 VDD2.n23 VDD2.n14 12.0247
R610 VDD2.n77 VDD2.n65 11.249
R611 VDD2.n24 VDD2.n12 11.249
R612 VDD2.n81 VDD2.n80 10.4732
R613 VDD2.n28 VDD2.n27 10.4732
R614 VDD2.n103 VDD2.n53 9.69747
R615 VDD2.n84 VDD2.n63 9.69747
R616 VDD2.n31 VDD2.n10 9.69747
R617 VDD2.n50 VDD2.n0 9.69747
R618 VDD2.n103 VDD2.n102 9.45567
R619 VDD2.n50 VDD2.n49 9.45567
R620 VDD2.n96 VDD2.n95 9.3005
R621 VDD2.n55 VDD2.n54 9.3005
R622 VDD2.n102 VDD2.n101 9.3005
R623 VDD2.n94 VDD2.n93 9.3005
R624 VDD2.n59 VDD2.n58 9.3005
R625 VDD2.n88 VDD2.n87 9.3005
R626 VDD2.n86 VDD2.n85 9.3005
R627 VDD2.n63 VDD2.n62 9.3005
R628 VDD2.n80 VDD2.n79 9.3005
R629 VDD2.n78 VDD2.n77 9.3005
R630 VDD2.n67 VDD2.n66 9.3005
R631 VDD2.n72 VDD2.n71 9.3005
R632 VDD2.n41 VDD2.n40 9.3005
R633 VDD2.n43 VDD2.n42 9.3005
R634 VDD2.n2 VDD2.n1 9.3005
R635 VDD2.n49 VDD2.n48 9.3005
R636 VDD2.n35 VDD2.n34 9.3005
R637 VDD2.n33 VDD2.n32 9.3005
R638 VDD2.n10 VDD2.n9 9.3005
R639 VDD2.n27 VDD2.n26 9.3005
R640 VDD2.n25 VDD2.n24 9.3005
R641 VDD2.n14 VDD2.n13 9.3005
R642 VDD2.n19 VDD2.n18 9.3005
R643 VDD2.n6 VDD2.n5 9.3005
R644 VDD2.n101 VDD2.n100 8.92171
R645 VDD2.n85 VDD2.n61 8.92171
R646 VDD2.n32 VDD2.n8 8.92171
R647 VDD2.n48 VDD2.n47 8.92171
R648 VDD2.n97 VDD2.n55 8.14595
R649 VDD2.n89 VDD2.n88 8.14595
R650 VDD2.n36 VDD2.n35 8.14595
R651 VDD2.n44 VDD2.n2 8.14595
R652 VDD2.n96 VDD2.n57 7.3702
R653 VDD2.n92 VDD2.n59 7.3702
R654 VDD2.n39 VDD2.n6 7.3702
R655 VDD2.n43 VDD2.n4 7.3702
R656 VDD2.n93 VDD2.n57 6.59444
R657 VDD2.n93 VDD2.n92 6.59444
R658 VDD2.n40 VDD2.n39 6.59444
R659 VDD2.n40 VDD2.n4 6.59444
R660 VDD2.n97 VDD2.n96 5.81868
R661 VDD2.n89 VDD2.n59 5.81868
R662 VDD2.n36 VDD2.n6 5.81868
R663 VDD2.n44 VDD2.n43 5.81868
R664 VDD2.n100 VDD2.n55 5.04292
R665 VDD2.n88 VDD2.n61 5.04292
R666 VDD2.n35 VDD2.n8 5.04292
R667 VDD2.n47 VDD2.n2 5.04292
R668 VDD2.n101 VDD2.n53 4.26717
R669 VDD2.n85 VDD2.n84 4.26717
R670 VDD2.n32 VDD2.n31 4.26717
R671 VDD2.n48 VDD2.n0 4.26717
R672 VDD2.n71 VDD2.n70 3.70984
R673 VDD2.n18 VDD2.n17 3.70984
R674 VDD2.n81 VDD2.n63 3.49141
R675 VDD2.n28 VDD2.n10 3.49141
R676 VDD2.n105 VDD2.t0 3.41848
R677 VDD2.n105 VDD2.t2 3.41848
R678 VDD2.n51 VDD2.t5 3.41848
R679 VDD2.n51 VDD2.t3 3.41848
R680 VDD2.n80 VDD2.n65 2.71565
R681 VDD2.n27 VDD2.n12 2.71565
R682 VDD2.n77 VDD2.n76 1.93989
R683 VDD2.n24 VDD2.n23 1.93989
R684 VDD2.n73 VDD2.n67 1.16414
R685 VDD2.n20 VDD2.n14 1.16414
R686 VDD2 VDD2.n104 0.938
R687 VDD2.n72 VDD2.n69 0.388379
R688 VDD2.n19 VDD2.n16 0.388379
R689 VDD2.n102 VDD2.n54 0.155672
R690 VDD2.n95 VDD2.n54 0.155672
R691 VDD2.n95 VDD2.n94 0.155672
R692 VDD2.n94 VDD2.n58 0.155672
R693 VDD2.n87 VDD2.n58 0.155672
R694 VDD2.n87 VDD2.n86 0.155672
R695 VDD2.n86 VDD2.n62 0.155672
R696 VDD2.n79 VDD2.n62 0.155672
R697 VDD2.n79 VDD2.n78 0.155672
R698 VDD2.n78 VDD2.n66 0.155672
R699 VDD2.n71 VDD2.n66 0.155672
R700 VDD2.n18 VDD2.n13 0.155672
R701 VDD2.n25 VDD2.n13 0.155672
R702 VDD2.n26 VDD2.n25 0.155672
R703 VDD2.n26 VDD2.n9 0.155672
R704 VDD2.n33 VDD2.n9 0.155672
R705 VDD2.n34 VDD2.n33 0.155672
R706 VDD2.n34 VDD2.n5 0.155672
R707 VDD2.n41 VDD2.n5 0.155672
R708 VDD2.n42 VDD2.n41 0.155672
R709 VDD2.n42 VDD2.n1 0.155672
R710 VDD2.n49 VDD2.n1 0.155672
R711 B.n364 B.n57 585
R712 B.n366 B.n365 585
R713 B.n367 B.n56 585
R714 B.n369 B.n368 585
R715 B.n370 B.n55 585
R716 B.n372 B.n371 585
R717 B.n373 B.n54 585
R718 B.n375 B.n374 585
R719 B.n376 B.n53 585
R720 B.n378 B.n377 585
R721 B.n379 B.n52 585
R722 B.n381 B.n380 585
R723 B.n382 B.n51 585
R724 B.n384 B.n383 585
R725 B.n385 B.n50 585
R726 B.n387 B.n386 585
R727 B.n388 B.n49 585
R728 B.n390 B.n389 585
R729 B.n391 B.n48 585
R730 B.n393 B.n392 585
R731 B.n394 B.n47 585
R732 B.n396 B.n395 585
R733 B.n397 B.n46 585
R734 B.n399 B.n398 585
R735 B.n400 B.n45 585
R736 B.n402 B.n401 585
R737 B.n403 B.n44 585
R738 B.n405 B.n404 585
R739 B.n406 B.n43 585
R740 B.n408 B.n407 585
R741 B.n409 B.n42 585
R742 B.n411 B.n410 585
R743 B.n412 B.n41 585
R744 B.n414 B.n413 585
R745 B.n416 B.n415 585
R746 B.n417 B.n37 585
R747 B.n419 B.n418 585
R748 B.n420 B.n36 585
R749 B.n422 B.n421 585
R750 B.n423 B.n35 585
R751 B.n425 B.n424 585
R752 B.n426 B.n34 585
R753 B.n428 B.n427 585
R754 B.n429 B.n31 585
R755 B.n432 B.n431 585
R756 B.n433 B.n30 585
R757 B.n435 B.n434 585
R758 B.n436 B.n29 585
R759 B.n438 B.n437 585
R760 B.n439 B.n28 585
R761 B.n441 B.n440 585
R762 B.n442 B.n27 585
R763 B.n444 B.n443 585
R764 B.n445 B.n26 585
R765 B.n447 B.n446 585
R766 B.n448 B.n25 585
R767 B.n450 B.n449 585
R768 B.n451 B.n24 585
R769 B.n453 B.n452 585
R770 B.n454 B.n23 585
R771 B.n456 B.n455 585
R772 B.n457 B.n22 585
R773 B.n459 B.n458 585
R774 B.n460 B.n21 585
R775 B.n462 B.n461 585
R776 B.n463 B.n20 585
R777 B.n465 B.n464 585
R778 B.n466 B.n19 585
R779 B.n468 B.n467 585
R780 B.n469 B.n18 585
R781 B.n471 B.n470 585
R782 B.n472 B.n17 585
R783 B.n474 B.n473 585
R784 B.n475 B.n16 585
R785 B.n477 B.n476 585
R786 B.n478 B.n15 585
R787 B.n480 B.n479 585
R788 B.n481 B.n14 585
R789 B.n363 B.n362 585
R790 B.n361 B.n58 585
R791 B.n360 B.n359 585
R792 B.n358 B.n59 585
R793 B.n357 B.n356 585
R794 B.n355 B.n60 585
R795 B.n354 B.n353 585
R796 B.n352 B.n61 585
R797 B.n351 B.n350 585
R798 B.n349 B.n62 585
R799 B.n348 B.n347 585
R800 B.n346 B.n63 585
R801 B.n345 B.n344 585
R802 B.n343 B.n64 585
R803 B.n342 B.n341 585
R804 B.n340 B.n65 585
R805 B.n339 B.n338 585
R806 B.n337 B.n66 585
R807 B.n336 B.n335 585
R808 B.n334 B.n67 585
R809 B.n333 B.n332 585
R810 B.n331 B.n68 585
R811 B.n330 B.n329 585
R812 B.n328 B.n69 585
R813 B.n327 B.n326 585
R814 B.n325 B.n70 585
R815 B.n324 B.n323 585
R816 B.n322 B.n71 585
R817 B.n321 B.n320 585
R818 B.n319 B.n72 585
R819 B.n318 B.n317 585
R820 B.n316 B.n73 585
R821 B.n315 B.n314 585
R822 B.n313 B.n74 585
R823 B.n312 B.n311 585
R824 B.n310 B.n75 585
R825 B.n309 B.n308 585
R826 B.n307 B.n76 585
R827 B.n306 B.n305 585
R828 B.n304 B.n77 585
R829 B.n303 B.n302 585
R830 B.n301 B.n78 585
R831 B.n300 B.n299 585
R832 B.n298 B.n79 585
R833 B.n297 B.n296 585
R834 B.n295 B.n80 585
R835 B.n294 B.n293 585
R836 B.n292 B.n81 585
R837 B.n291 B.n290 585
R838 B.n172 B.n125 585
R839 B.n174 B.n173 585
R840 B.n175 B.n124 585
R841 B.n177 B.n176 585
R842 B.n178 B.n123 585
R843 B.n180 B.n179 585
R844 B.n181 B.n122 585
R845 B.n183 B.n182 585
R846 B.n184 B.n121 585
R847 B.n186 B.n185 585
R848 B.n187 B.n120 585
R849 B.n189 B.n188 585
R850 B.n190 B.n119 585
R851 B.n192 B.n191 585
R852 B.n193 B.n118 585
R853 B.n195 B.n194 585
R854 B.n196 B.n117 585
R855 B.n198 B.n197 585
R856 B.n199 B.n116 585
R857 B.n201 B.n200 585
R858 B.n202 B.n115 585
R859 B.n204 B.n203 585
R860 B.n205 B.n114 585
R861 B.n207 B.n206 585
R862 B.n208 B.n113 585
R863 B.n210 B.n209 585
R864 B.n211 B.n112 585
R865 B.n213 B.n212 585
R866 B.n214 B.n111 585
R867 B.n216 B.n215 585
R868 B.n217 B.n110 585
R869 B.n219 B.n218 585
R870 B.n220 B.n109 585
R871 B.n222 B.n221 585
R872 B.n224 B.n223 585
R873 B.n225 B.n105 585
R874 B.n227 B.n226 585
R875 B.n228 B.n104 585
R876 B.n230 B.n229 585
R877 B.n231 B.n103 585
R878 B.n233 B.n232 585
R879 B.n234 B.n102 585
R880 B.n236 B.n235 585
R881 B.n237 B.n99 585
R882 B.n240 B.n239 585
R883 B.n241 B.n98 585
R884 B.n243 B.n242 585
R885 B.n244 B.n97 585
R886 B.n246 B.n245 585
R887 B.n247 B.n96 585
R888 B.n249 B.n248 585
R889 B.n250 B.n95 585
R890 B.n252 B.n251 585
R891 B.n253 B.n94 585
R892 B.n255 B.n254 585
R893 B.n256 B.n93 585
R894 B.n258 B.n257 585
R895 B.n259 B.n92 585
R896 B.n261 B.n260 585
R897 B.n262 B.n91 585
R898 B.n264 B.n263 585
R899 B.n265 B.n90 585
R900 B.n267 B.n266 585
R901 B.n268 B.n89 585
R902 B.n270 B.n269 585
R903 B.n271 B.n88 585
R904 B.n273 B.n272 585
R905 B.n274 B.n87 585
R906 B.n276 B.n275 585
R907 B.n277 B.n86 585
R908 B.n279 B.n278 585
R909 B.n280 B.n85 585
R910 B.n282 B.n281 585
R911 B.n283 B.n84 585
R912 B.n285 B.n284 585
R913 B.n286 B.n83 585
R914 B.n288 B.n287 585
R915 B.n289 B.n82 585
R916 B.n171 B.n170 585
R917 B.n169 B.n126 585
R918 B.n168 B.n167 585
R919 B.n166 B.n127 585
R920 B.n165 B.n164 585
R921 B.n163 B.n128 585
R922 B.n162 B.n161 585
R923 B.n160 B.n129 585
R924 B.n159 B.n158 585
R925 B.n157 B.n130 585
R926 B.n156 B.n155 585
R927 B.n154 B.n131 585
R928 B.n153 B.n152 585
R929 B.n151 B.n132 585
R930 B.n150 B.n149 585
R931 B.n148 B.n133 585
R932 B.n147 B.n146 585
R933 B.n145 B.n134 585
R934 B.n144 B.n143 585
R935 B.n142 B.n135 585
R936 B.n141 B.n140 585
R937 B.n139 B.n136 585
R938 B.n138 B.n137 585
R939 B.n2 B.n0 585
R940 B.n517 B.n1 585
R941 B.n516 B.n515 585
R942 B.n514 B.n3 585
R943 B.n513 B.n512 585
R944 B.n511 B.n4 585
R945 B.n510 B.n509 585
R946 B.n508 B.n5 585
R947 B.n507 B.n506 585
R948 B.n505 B.n6 585
R949 B.n504 B.n503 585
R950 B.n502 B.n7 585
R951 B.n501 B.n500 585
R952 B.n499 B.n8 585
R953 B.n498 B.n497 585
R954 B.n496 B.n9 585
R955 B.n495 B.n494 585
R956 B.n493 B.n10 585
R957 B.n492 B.n491 585
R958 B.n490 B.n11 585
R959 B.n489 B.n488 585
R960 B.n487 B.n12 585
R961 B.n486 B.n485 585
R962 B.n484 B.n13 585
R963 B.n483 B.n482 585
R964 B.n519 B.n518 585
R965 B.n170 B.n125 530.939
R966 B.n482 B.n481 530.939
R967 B.n290 B.n289 530.939
R968 B.n362 B.n57 530.939
R969 B.n100 B.t0 425.642
R970 B.n106 B.t6 425.642
R971 B.n32 B.t3 425.642
R972 B.n38 B.t9 425.642
R973 B.n100 B.t2 357.402
R974 B.n38 B.t10 357.402
R975 B.n106 B.t8 357.402
R976 B.n32 B.t4 357.402
R977 B.n101 B.t1 331.027
R978 B.n39 B.t11 331.027
R979 B.n107 B.t7 331.026
R980 B.n33 B.t5 331.026
R981 B.n170 B.n169 163.367
R982 B.n169 B.n168 163.367
R983 B.n168 B.n127 163.367
R984 B.n164 B.n127 163.367
R985 B.n164 B.n163 163.367
R986 B.n163 B.n162 163.367
R987 B.n162 B.n129 163.367
R988 B.n158 B.n129 163.367
R989 B.n158 B.n157 163.367
R990 B.n157 B.n156 163.367
R991 B.n156 B.n131 163.367
R992 B.n152 B.n131 163.367
R993 B.n152 B.n151 163.367
R994 B.n151 B.n150 163.367
R995 B.n150 B.n133 163.367
R996 B.n146 B.n133 163.367
R997 B.n146 B.n145 163.367
R998 B.n145 B.n144 163.367
R999 B.n144 B.n135 163.367
R1000 B.n140 B.n135 163.367
R1001 B.n140 B.n139 163.367
R1002 B.n139 B.n138 163.367
R1003 B.n138 B.n2 163.367
R1004 B.n518 B.n2 163.367
R1005 B.n518 B.n517 163.367
R1006 B.n517 B.n516 163.367
R1007 B.n516 B.n3 163.367
R1008 B.n512 B.n3 163.367
R1009 B.n512 B.n511 163.367
R1010 B.n511 B.n510 163.367
R1011 B.n510 B.n5 163.367
R1012 B.n506 B.n5 163.367
R1013 B.n506 B.n505 163.367
R1014 B.n505 B.n504 163.367
R1015 B.n504 B.n7 163.367
R1016 B.n500 B.n7 163.367
R1017 B.n500 B.n499 163.367
R1018 B.n499 B.n498 163.367
R1019 B.n498 B.n9 163.367
R1020 B.n494 B.n9 163.367
R1021 B.n494 B.n493 163.367
R1022 B.n493 B.n492 163.367
R1023 B.n492 B.n11 163.367
R1024 B.n488 B.n11 163.367
R1025 B.n488 B.n487 163.367
R1026 B.n487 B.n486 163.367
R1027 B.n486 B.n13 163.367
R1028 B.n482 B.n13 163.367
R1029 B.n174 B.n125 163.367
R1030 B.n175 B.n174 163.367
R1031 B.n176 B.n175 163.367
R1032 B.n176 B.n123 163.367
R1033 B.n180 B.n123 163.367
R1034 B.n181 B.n180 163.367
R1035 B.n182 B.n181 163.367
R1036 B.n182 B.n121 163.367
R1037 B.n186 B.n121 163.367
R1038 B.n187 B.n186 163.367
R1039 B.n188 B.n187 163.367
R1040 B.n188 B.n119 163.367
R1041 B.n192 B.n119 163.367
R1042 B.n193 B.n192 163.367
R1043 B.n194 B.n193 163.367
R1044 B.n194 B.n117 163.367
R1045 B.n198 B.n117 163.367
R1046 B.n199 B.n198 163.367
R1047 B.n200 B.n199 163.367
R1048 B.n200 B.n115 163.367
R1049 B.n204 B.n115 163.367
R1050 B.n205 B.n204 163.367
R1051 B.n206 B.n205 163.367
R1052 B.n206 B.n113 163.367
R1053 B.n210 B.n113 163.367
R1054 B.n211 B.n210 163.367
R1055 B.n212 B.n211 163.367
R1056 B.n212 B.n111 163.367
R1057 B.n216 B.n111 163.367
R1058 B.n217 B.n216 163.367
R1059 B.n218 B.n217 163.367
R1060 B.n218 B.n109 163.367
R1061 B.n222 B.n109 163.367
R1062 B.n223 B.n222 163.367
R1063 B.n223 B.n105 163.367
R1064 B.n227 B.n105 163.367
R1065 B.n228 B.n227 163.367
R1066 B.n229 B.n228 163.367
R1067 B.n229 B.n103 163.367
R1068 B.n233 B.n103 163.367
R1069 B.n234 B.n233 163.367
R1070 B.n235 B.n234 163.367
R1071 B.n235 B.n99 163.367
R1072 B.n240 B.n99 163.367
R1073 B.n241 B.n240 163.367
R1074 B.n242 B.n241 163.367
R1075 B.n242 B.n97 163.367
R1076 B.n246 B.n97 163.367
R1077 B.n247 B.n246 163.367
R1078 B.n248 B.n247 163.367
R1079 B.n248 B.n95 163.367
R1080 B.n252 B.n95 163.367
R1081 B.n253 B.n252 163.367
R1082 B.n254 B.n253 163.367
R1083 B.n254 B.n93 163.367
R1084 B.n258 B.n93 163.367
R1085 B.n259 B.n258 163.367
R1086 B.n260 B.n259 163.367
R1087 B.n260 B.n91 163.367
R1088 B.n264 B.n91 163.367
R1089 B.n265 B.n264 163.367
R1090 B.n266 B.n265 163.367
R1091 B.n266 B.n89 163.367
R1092 B.n270 B.n89 163.367
R1093 B.n271 B.n270 163.367
R1094 B.n272 B.n271 163.367
R1095 B.n272 B.n87 163.367
R1096 B.n276 B.n87 163.367
R1097 B.n277 B.n276 163.367
R1098 B.n278 B.n277 163.367
R1099 B.n278 B.n85 163.367
R1100 B.n282 B.n85 163.367
R1101 B.n283 B.n282 163.367
R1102 B.n284 B.n283 163.367
R1103 B.n284 B.n83 163.367
R1104 B.n288 B.n83 163.367
R1105 B.n289 B.n288 163.367
R1106 B.n290 B.n81 163.367
R1107 B.n294 B.n81 163.367
R1108 B.n295 B.n294 163.367
R1109 B.n296 B.n295 163.367
R1110 B.n296 B.n79 163.367
R1111 B.n300 B.n79 163.367
R1112 B.n301 B.n300 163.367
R1113 B.n302 B.n301 163.367
R1114 B.n302 B.n77 163.367
R1115 B.n306 B.n77 163.367
R1116 B.n307 B.n306 163.367
R1117 B.n308 B.n307 163.367
R1118 B.n308 B.n75 163.367
R1119 B.n312 B.n75 163.367
R1120 B.n313 B.n312 163.367
R1121 B.n314 B.n313 163.367
R1122 B.n314 B.n73 163.367
R1123 B.n318 B.n73 163.367
R1124 B.n319 B.n318 163.367
R1125 B.n320 B.n319 163.367
R1126 B.n320 B.n71 163.367
R1127 B.n324 B.n71 163.367
R1128 B.n325 B.n324 163.367
R1129 B.n326 B.n325 163.367
R1130 B.n326 B.n69 163.367
R1131 B.n330 B.n69 163.367
R1132 B.n331 B.n330 163.367
R1133 B.n332 B.n331 163.367
R1134 B.n332 B.n67 163.367
R1135 B.n336 B.n67 163.367
R1136 B.n337 B.n336 163.367
R1137 B.n338 B.n337 163.367
R1138 B.n338 B.n65 163.367
R1139 B.n342 B.n65 163.367
R1140 B.n343 B.n342 163.367
R1141 B.n344 B.n343 163.367
R1142 B.n344 B.n63 163.367
R1143 B.n348 B.n63 163.367
R1144 B.n349 B.n348 163.367
R1145 B.n350 B.n349 163.367
R1146 B.n350 B.n61 163.367
R1147 B.n354 B.n61 163.367
R1148 B.n355 B.n354 163.367
R1149 B.n356 B.n355 163.367
R1150 B.n356 B.n59 163.367
R1151 B.n360 B.n59 163.367
R1152 B.n361 B.n360 163.367
R1153 B.n362 B.n361 163.367
R1154 B.n481 B.n480 163.367
R1155 B.n480 B.n15 163.367
R1156 B.n476 B.n15 163.367
R1157 B.n476 B.n475 163.367
R1158 B.n475 B.n474 163.367
R1159 B.n474 B.n17 163.367
R1160 B.n470 B.n17 163.367
R1161 B.n470 B.n469 163.367
R1162 B.n469 B.n468 163.367
R1163 B.n468 B.n19 163.367
R1164 B.n464 B.n19 163.367
R1165 B.n464 B.n463 163.367
R1166 B.n463 B.n462 163.367
R1167 B.n462 B.n21 163.367
R1168 B.n458 B.n21 163.367
R1169 B.n458 B.n457 163.367
R1170 B.n457 B.n456 163.367
R1171 B.n456 B.n23 163.367
R1172 B.n452 B.n23 163.367
R1173 B.n452 B.n451 163.367
R1174 B.n451 B.n450 163.367
R1175 B.n450 B.n25 163.367
R1176 B.n446 B.n25 163.367
R1177 B.n446 B.n445 163.367
R1178 B.n445 B.n444 163.367
R1179 B.n444 B.n27 163.367
R1180 B.n440 B.n27 163.367
R1181 B.n440 B.n439 163.367
R1182 B.n439 B.n438 163.367
R1183 B.n438 B.n29 163.367
R1184 B.n434 B.n29 163.367
R1185 B.n434 B.n433 163.367
R1186 B.n433 B.n432 163.367
R1187 B.n432 B.n31 163.367
R1188 B.n427 B.n31 163.367
R1189 B.n427 B.n426 163.367
R1190 B.n426 B.n425 163.367
R1191 B.n425 B.n35 163.367
R1192 B.n421 B.n35 163.367
R1193 B.n421 B.n420 163.367
R1194 B.n420 B.n419 163.367
R1195 B.n419 B.n37 163.367
R1196 B.n415 B.n37 163.367
R1197 B.n415 B.n414 163.367
R1198 B.n414 B.n41 163.367
R1199 B.n410 B.n41 163.367
R1200 B.n410 B.n409 163.367
R1201 B.n409 B.n408 163.367
R1202 B.n408 B.n43 163.367
R1203 B.n404 B.n43 163.367
R1204 B.n404 B.n403 163.367
R1205 B.n403 B.n402 163.367
R1206 B.n402 B.n45 163.367
R1207 B.n398 B.n45 163.367
R1208 B.n398 B.n397 163.367
R1209 B.n397 B.n396 163.367
R1210 B.n396 B.n47 163.367
R1211 B.n392 B.n47 163.367
R1212 B.n392 B.n391 163.367
R1213 B.n391 B.n390 163.367
R1214 B.n390 B.n49 163.367
R1215 B.n386 B.n49 163.367
R1216 B.n386 B.n385 163.367
R1217 B.n385 B.n384 163.367
R1218 B.n384 B.n51 163.367
R1219 B.n380 B.n51 163.367
R1220 B.n380 B.n379 163.367
R1221 B.n379 B.n378 163.367
R1222 B.n378 B.n53 163.367
R1223 B.n374 B.n53 163.367
R1224 B.n374 B.n373 163.367
R1225 B.n373 B.n372 163.367
R1226 B.n372 B.n55 163.367
R1227 B.n368 B.n55 163.367
R1228 B.n368 B.n367 163.367
R1229 B.n367 B.n366 163.367
R1230 B.n366 B.n57 163.367
R1231 B.n238 B.n101 59.5399
R1232 B.n108 B.n107 59.5399
R1233 B.n430 B.n33 59.5399
R1234 B.n40 B.n39 59.5399
R1235 B.n483 B.n14 34.4981
R1236 B.n364 B.n363 34.4981
R1237 B.n291 B.n82 34.4981
R1238 B.n172 B.n171 34.4981
R1239 B.n101 B.n100 26.3763
R1240 B.n107 B.n106 26.3763
R1241 B.n33 B.n32 26.3763
R1242 B.n39 B.n38 26.3763
R1243 B B.n519 18.0485
R1244 B.n479 B.n14 10.6151
R1245 B.n479 B.n478 10.6151
R1246 B.n478 B.n477 10.6151
R1247 B.n477 B.n16 10.6151
R1248 B.n473 B.n16 10.6151
R1249 B.n473 B.n472 10.6151
R1250 B.n472 B.n471 10.6151
R1251 B.n471 B.n18 10.6151
R1252 B.n467 B.n18 10.6151
R1253 B.n467 B.n466 10.6151
R1254 B.n466 B.n465 10.6151
R1255 B.n465 B.n20 10.6151
R1256 B.n461 B.n20 10.6151
R1257 B.n461 B.n460 10.6151
R1258 B.n460 B.n459 10.6151
R1259 B.n459 B.n22 10.6151
R1260 B.n455 B.n22 10.6151
R1261 B.n455 B.n454 10.6151
R1262 B.n454 B.n453 10.6151
R1263 B.n453 B.n24 10.6151
R1264 B.n449 B.n24 10.6151
R1265 B.n449 B.n448 10.6151
R1266 B.n448 B.n447 10.6151
R1267 B.n447 B.n26 10.6151
R1268 B.n443 B.n26 10.6151
R1269 B.n443 B.n442 10.6151
R1270 B.n442 B.n441 10.6151
R1271 B.n441 B.n28 10.6151
R1272 B.n437 B.n28 10.6151
R1273 B.n437 B.n436 10.6151
R1274 B.n436 B.n435 10.6151
R1275 B.n435 B.n30 10.6151
R1276 B.n431 B.n30 10.6151
R1277 B.n429 B.n428 10.6151
R1278 B.n428 B.n34 10.6151
R1279 B.n424 B.n34 10.6151
R1280 B.n424 B.n423 10.6151
R1281 B.n423 B.n422 10.6151
R1282 B.n422 B.n36 10.6151
R1283 B.n418 B.n36 10.6151
R1284 B.n418 B.n417 10.6151
R1285 B.n417 B.n416 10.6151
R1286 B.n413 B.n412 10.6151
R1287 B.n412 B.n411 10.6151
R1288 B.n411 B.n42 10.6151
R1289 B.n407 B.n42 10.6151
R1290 B.n407 B.n406 10.6151
R1291 B.n406 B.n405 10.6151
R1292 B.n405 B.n44 10.6151
R1293 B.n401 B.n44 10.6151
R1294 B.n401 B.n400 10.6151
R1295 B.n400 B.n399 10.6151
R1296 B.n399 B.n46 10.6151
R1297 B.n395 B.n46 10.6151
R1298 B.n395 B.n394 10.6151
R1299 B.n394 B.n393 10.6151
R1300 B.n393 B.n48 10.6151
R1301 B.n389 B.n48 10.6151
R1302 B.n389 B.n388 10.6151
R1303 B.n388 B.n387 10.6151
R1304 B.n387 B.n50 10.6151
R1305 B.n383 B.n50 10.6151
R1306 B.n383 B.n382 10.6151
R1307 B.n382 B.n381 10.6151
R1308 B.n381 B.n52 10.6151
R1309 B.n377 B.n52 10.6151
R1310 B.n377 B.n376 10.6151
R1311 B.n376 B.n375 10.6151
R1312 B.n375 B.n54 10.6151
R1313 B.n371 B.n54 10.6151
R1314 B.n371 B.n370 10.6151
R1315 B.n370 B.n369 10.6151
R1316 B.n369 B.n56 10.6151
R1317 B.n365 B.n56 10.6151
R1318 B.n365 B.n364 10.6151
R1319 B.n292 B.n291 10.6151
R1320 B.n293 B.n292 10.6151
R1321 B.n293 B.n80 10.6151
R1322 B.n297 B.n80 10.6151
R1323 B.n298 B.n297 10.6151
R1324 B.n299 B.n298 10.6151
R1325 B.n299 B.n78 10.6151
R1326 B.n303 B.n78 10.6151
R1327 B.n304 B.n303 10.6151
R1328 B.n305 B.n304 10.6151
R1329 B.n305 B.n76 10.6151
R1330 B.n309 B.n76 10.6151
R1331 B.n310 B.n309 10.6151
R1332 B.n311 B.n310 10.6151
R1333 B.n311 B.n74 10.6151
R1334 B.n315 B.n74 10.6151
R1335 B.n316 B.n315 10.6151
R1336 B.n317 B.n316 10.6151
R1337 B.n317 B.n72 10.6151
R1338 B.n321 B.n72 10.6151
R1339 B.n322 B.n321 10.6151
R1340 B.n323 B.n322 10.6151
R1341 B.n323 B.n70 10.6151
R1342 B.n327 B.n70 10.6151
R1343 B.n328 B.n327 10.6151
R1344 B.n329 B.n328 10.6151
R1345 B.n329 B.n68 10.6151
R1346 B.n333 B.n68 10.6151
R1347 B.n334 B.n333 10.6151
R1348 B.n335 B.n334 10.6151
R1349 B.n335 B.n66 10.6151
R1350 B.n339 B.n66 10.6151
R1351 B.n340 B.n339 10.6151
R1352 B.n341 B.n340 10.6151
R1353 B.n341 B.n64 10.6151
R1354 B.n345 B.n64 10.6151
R1355 B.n346 B.n345 10.6151
R1356 B.n347 B.n346 10.6151
R1357 B.n347 B.n62 10.6151
R1358 B.n351 B.n62 10.6151
R1359 B.n352 B.n351 10.6151
R1360 B.n353 B.n352 10.6151
R1361 B.n353 B.n60 10.6151
R1362 B.n357 B.n60 10.6151
R1363 B.n358 B.n357 10.6151
R1364 B.n359 B.n358 10.6151
R1365 B.n359 B.n58 10.6151
R1366 B.n363 B.n58 10.6151
R1367 B.n173 B.n172 10.6151
R1368 B.n173 B.n124 10.6151
R1369 B.n177 B.n124 10.6151
R1370 B.n178 B.n177 10.6151
R1371 B.n179 B.n178 10.6151
R1372 B.n179 B.n122 10.6151
R1373 B.n183 B.n122 10.6151
R1374 B.n184 B.n183 10.6151
R1375 B.n185 B.n184 10.6151
R1376 B.n185 B.n120 10.6151
R1377 B.n189 B.n120 10.6151
R1378 B.n190 B.n189 10.6151
R1379 B.n191 B.n190 10.6151
R1380 B.n191 B.n118 10.6151
R1381 B.n195 B.n118 10.6151
R1382 B.n196 B.n195 10.6151
R1383 B.n197 B.n196 10.6151
R1384 B.n197 B.n116 10.6151
R1385 B.n201 B.n116 10.6151
R1386 B.n202 B.n201 10.6151
R1387 B.n203 B.n202 10.6151
R1388 B.n203 B.n114 10.6151
R1389 B.n207 B.n114 10.6151
R1390 B.n208 B.n207 10.6151
R1391 B.n209 B.n208 10.6151
R1392 B.n209 B.n112 10.6151
R1393 B.n213 B.n112 10.6151
R1394 B.n214 B.n213 10.6151
R1395 B.n215 B.n214 10.6151
R1396 B.n215 B.n110 10.6151
R1397 B.n219 B.n110 10.6151
R1398 B.n220 B.n219 10.6151
R1399 B.n221 B.n220 10.6151
R1400 B.n225 B.n224 10.6151
R1401 B.n226 B.n225 10.6151
R1402 B.n226 B.n104 10.6151
R1403 B.n230 B.n104 10.6151
R1404 B.n231 B.n230 10.6151
R1405 B.n232 B.n231 10.6151
R1406 B.n232 B.n102 10.6151
R1407 B.n236 B.n102 10.6151
R1408 B.n237 B.n236 10.6151
R1409 B.n239 B.n98 10.6151
R1410 B.n243 B.n98 10.6151
R1411 B.n244 B.n243 10.6151
R1412 B.n245 B.n244 10.6151
R1413 B.n245 B.n96 10.6151
R1414 B.n249 B.n96 10.6151
R1415 B.n250 B.n249 10.6151
R1416 B.n251 B.n250 10.6151
R1417 B.n251 B.n94 10.6151
R1418 B.n255 B.n94 10.6151
R1419 B.n256 B.n255 10.6151
R1420 B.n257 B.n256 10.6151
R1421 B.n257 B.n92 10.6151
R1422 B.n261 B.n92 10.6151
R1423 B.n262 B.n261 10.6151
R1424 B.n263 B.n262 10.6151
R1425 B.n263 B.n90 10.6151
R1426 B.n267 B.n90 10.6151
R1427 B.n268 B.n267 10.6151
R1428 B.n269 B.n268 10.6151
R1429 B.n269 B.n88 10.6151
R1430 B.n273 B.n88 10.6151
R1431 B.n274 B.n273 10.6151
R1432 B.n275 B.n274 10.6151
R1433 B.n275 B.n86 10.6151
R1434 B.n279 B.n86 10.6151
R1435 B.n280 B.n279 10.6151
R1436 B.n281 B.n280 10.6151
R1437 B.n281 B.n84 10.6151
R1438 B.n285 B.n84 10.6151
R1439 B.n286 B.n285 10.6151
R1440 B.n287 B.n286 10.6151
R1441 B.n287 B.n82 10.6151
R1442 B.n171 B.n126 10.6151
R1443 B.n167 B.n126 10.6151
R1444 B.n167 B.n166 10.6151
R1445 B.n166 B.n165 10.6151
R1446 B.n165 B.n128 10.6151
R1447 B.n161 B.n128 10.6151
R1448 B.n161 B.n160 10.6151
R1449 B.n160 B.n159 10.6151
R1450 B.n159 B.n130 10.6151
R1451 B.n155 B.n130 10.6151
R1452 B.n155 B.n154 10.6151
R1453 B.n154 B.n153 10.6151
R1454 B.n153 B.n132 10.6151
R1455 B.n149 B.n132 10.6151
R1456 B.n149 B.n148 10.6151
R1457 B.n148 B.n147 10.6151
R1458 B.n147 B.n134 10.6151
R1459 B.n143 B.n134 10.6151
R1460 B.n143 B.n142 10.6151
R1461 B.n142 B.n141 10.6151
R1462 B.n141 B.n136 10.6151
R1463 B.n137 B.n136 10.6151
R1464 B.n137 B.n0 10.6151
R1465 B.n515 B.n1 10.6151
R1466 B.n515 B.n514 10.6151
R1467 B.n514 B.n513 10.6151
R1468 B.n513 B.n4 10.6151
R1469 B.n509 B.n4 10.6151
R1470 B.n509 B.n508 10.6151
R1471 B.n508 B.n507 10.6151
R1472 B.n507 B.n6 10.6151
R1473 B.n503 B.n6 10.6151
R1474 B.n503 B.n502 10.6151
R1475 B.n502 B.n501 10.6151
R1476 B.n501 B.n8 10.6151
R1477 B.n497 B.n8 10.6151
R1478 B.n497 B.n496 10.6151
R1479 B.n496 B.n495 10.6151
R1480 B.n495 B.n10 10.6151
R1481 B.n491 B.n10 10.6151
R1482 B.n491 B.n490 10.6151
R1483 B.n490 B.n489 10.6151
R1484 B.n489 B.n12 10.6151
R1485 B.n485 B.n12 10.6151
R1486 B.n485 B.n484 10.6151
R1487 B.n484 B.n483 10.6151
R1488 B.n431 B.n430 9.36635
R1489 B.n413 B.n40 9.36635
R1490 B.n221 B.n108 9.36635
R1491 B.n239 B.n238 9.36635
R1492 B.n519 B.n0 2.81026
R1493 B.n519 B.n1 2.81026
R1494 B.n430 B.n429 1.24928
R1495 B.n416 B.n40 1.24928
R1496 B.n224 B.n108 1.24928
R1497 B.n238 B.n237 1.24928
C0 w_n2058_n2870# VDD2 1.75422f
C1 VTAIL VDD1 7.359479f
C2 VTAIL VN 4.02924f
C3 VP VDD2 0.325196f
C4 B VDD1 1.47395f
C5 VN B 0.805472f
C6 w_n2058_n2870# VDD1 1.71961f
C7 w_n2058_n2870# VN 3.47503f
C8 VP VDD1 4.32379f
C9 VN VP 4.94197f
C10 VTAIL B 2.44758f
C11 w_n2058_n2870# VTAIL 2.54878f
C12 VDD1 VDD2 0.831379f
C13 VN VDD2 4.150609f
C14 VTAIL VP 4.04367f
C15 w_n2058_n2870# B 6.81035f
C16 VN VDD1 0.148654f
C17 VP B 1.2345f
C18 VTAIL VDD2 7.398069f
C19 w_n2058_n2870# VP 3.73672f
C20 B VDD2 1.51068f
C21 VDD2 VSUBS 1.273683f
C22 VDD1 VSUBS 1.151609f
C23 VTAIL VSUBS 0.775091f
C24 VN VSUBS 4.438099f
C25 VP VSUBS 1.649231f
C26 B VSUBS 2.876425f
C27 w_n2058_n2870# VSUBS 73.0261f
C28 B.n0 VSUBS 0.004679f
C29 B.n1 VSUBS 0.004679f
C30 B.n2 VSUBS 0.007399f
C31 B.n3 VSUBS 0.007399f
C32 B.n4 VSUBS 0.007399f
C33 B.n5 VSUBS 0.007399f
C34 B.n6 VSUBS 0.007399f
C35 B.n7 VSUBS 0.007399f
C36 B.n8 VSUBS 0.007399f
C37 B.n9 VSUBS 0.007399f
C38 B.n10 VSUBS 0.007399f
C39 B.n11 VSUBS 0.007399f
C40 B.n12 VSUBS 0.007399f
C41 B.n13 VSUBS 0.007399f
C42 B.n14 VSUBS 0.018366f
C43 B.n15 VSUBS 0.007399f
C44 B.n16 VSUBS 0.007399f
C45 B.n17 VSUBS 0.007399f
C46 B.n18 VSUBS 0.007399f
C47 B.n19 VSUBS 0.007399f
C48 B.n20 VSUBS 0.007399f
C49 B.n21 VSUBS 0.007399f
C50 B.n22 VSUBS 0.007399f
C51 B.n23 VSUBS 0.007399f
C52 B.n24 VSUBS 0.007399f
C53 B.n25 VSUBS 0.007399f
C54 B.n26 VSUBS 0.007399f
C55 B.n27 VSUBS 0.007399f
C56 B.n28 VSUBS 0.007399f
C57 B.n29 VSUBS 0.007399f
C58 B.n30 VSUBS 0.007399f
C59 B.n31 VSUBS 0.007399f
C60 B.t5 VSUBS 0.166488f
C61 B.t4 VSUBS 0.181996f
C62 B.t3 VSUBS 0.446776f
C63 B.n32 VSUBS 0.285438f
C64 B.n33 VSUBS 0.220702f
C65 B.n34 VSUBS 0.007399f
C66 B.n35 VSUBS 0.007399f
C67 B.n36 VSUBS 0.007399f
C68 B.n37 VSUBS 0.007399f
C69 B.t11 VSUBS 0.16649f
C70 B.t10 VSUBS 0.181999f
C71 B.t9 VSUBS 0.446776f
C72 B.n38 VSUBS 0.285435f
C73 B.n39 VSUBS 0.220699f
C74 B.n40 VSUBS 0.017142f
C75 B.n41 VSUBS 0.007399f
C76 B.n42 VSUBS 0.007399f
C77 B.n43 VSUBS 0.007399f
C78 B.n44 VSUBS 0.007399f
C79 B.n45 VSUBS 0.007399f
C80 B.n46 VSUBS 0.007399f
C81 B.n47 VSUBS 0.007399f
C82 B.n48 VSUBS 0.007399f
C83 B.n49 VSUBS 0.007399f
C84 B.n50 VSUBS 0.007399f
C85 B.n51 VSUBS 0.007399f
C86 B.n52 VSUBS 0.007399f
C87 B.n53 VSUBS 0.007399f
C88 B.n54 VSUBS 0.007399f
C89 B.n55 VSUBS 0.007399f
C90 B.n56 VSUBS 0.007399f
C91 B.n57 VSUBS 0.018366f
C92 B.n58 VSUBS 0.007399f
C93 B.n59 VSUBS 0.007399f
C94 B.n60 VSUBS 0.007399f
C95 B.n61 VSUBS 0.007399f
C96 B.n62 VSUBS 0.007399f
C97 B.n63 VSUBS 0.007399f
C98 B.n64 VSUBS 0.007399f
C99 B.n65 VSUBS 0.007399f
C100 B.n66 VSUBS 0.007399f
C101 B.n67 VSUBS 0.007399f
C102 B.n68 VSUBS 0.007399f
C103 B.n69 VSUBS 0.007399f
C104 B.n70 VSUBS 0.007399f
C105 B.n71 VSUBS 0.007399f
C106 B.n72 VSUBS 0.007399f
C107 B.n73 VSUBS 0.007399f
C108 B.n74 VSUBS 0.007399f
C109 B.n75 VSUBS 0.007399f
C110 B.n76 VSUBS 0.007399f
C111 B.n77 VSUBS 0.007399f
C112 B.n78 VSUBS 0.007399f
C113 B.n79 VSUBS 0.007399f
C114 B.n80 VSUBS 0.007399f
C115 B.n81 VSUBS 0.007399f
C116 B.n82 VSUBS 0.018366f
C117 B.n83 VSUBS 0.007399f
C118 B.n84 VSUBS 0.007399f
C119 B.n85 VSUBS 0.007399f
C120 B.n86 VSUBS 0.007399f
C121 B.n87 VSUBS 0.007399f
C122 B.n88 VSUBS 0.007399f
C123 B.n89 VSUBS 0.007399f
C124 B.n90 VSUBS 0.007399f
C125 B.n91 VSUBS 0.007399f
C126 B.n92 VSUBS 0.007399f
C127 B.n93 VSUBS 0.007399f
C128 B.n94 VSUBS 0.007399f
C129 B.n95 VSUBS 0.007399f
C130 B.n96 VSUBS 0.007399f
C131 B.n97 VSUBS 0.007399f
C132 B.n98 VSUBS 0.007399f
C133 B.n99 VSUBS 0.007399f
C134 B.t1 VSUBS 0.16649f
C135 B.t2 VSUBS 0.181999f
C136 B.t0 VSUBS 0.446776f
C137 B.n100 VSUBS 0.285435f
C138 B.n101 VSUBS 0.220699f
C139 B.n102 VSUBS 0.007399f
C140 B.n103 VSUBS 0.007399f
C141 B.n104 VSUBS 0.007399f
C142 B.n105 VSUBS 0.007399f
C143 B.t7 VSUBS 0.166488f
C144 B.t8 VSUBS 0.181996f
C145 B.t6 VSUBS 0.446776f
C146 B.n106 VSUBS 0.285438f
C147 B.n107 VSUBS 0.220702f
C148 B.n108 VSUBS 0.017142f
C149 B.n109 VSUBS 0.007399f
C150 B.n110 VSUBS 0.007399f
C151 B.n111 VSUBS 0.007399f
C152 B.n112 VSUBS 0.007399f
C153 B.n113 VSUBS 0.007399f
C154 B.n114 VSUBS 0.007399f
C155 B.n115 VSUBS 0.007399f
C156 B.n116 VSUBS 0.007399f
C157 B.n117 VSUBS 0.007399f
C158 B.n118 VSUBS 0.007399f
C159 B.n119 VSUBS 0.007399f
C160 B.n120 VSUBS 0.007399f
C161 B.n121 VSUBS 0.007399f
C162 B.n122 VSUBS 0.007399f
C163 B.n123 VSUBS 0.007399f
C164 B.n124 VSUBS 0.007399f
C165 B.n125 VSUBS 0.018366f
C166 B.n126 VSUBS 0.007399f
C167 B.n127 VSUBS 0.007399f
C168 B.n128 VSUBS 0.007399f
C169 B.n129 VSUBS 0.007399f
C170 B.n130 VSUBS 0.007399f
C171 B.n131 VSUBS 0.007399f
C172 B.n132 VSUBS 0.007399f
C173 B.n133 VSUBS 0.007399f
C174 B.n134 VSUBS 0.007399f
C175 B.n135 VSUBS 0.007399f
C176 B.n136 VSUBS 0.007399f
C177 B.n137 VSUBS 0.007399f
C178 B.n138 VSUBS 0.007399f
C179 B.n139 VSUBS 0.007399f
C180 B.n140 VSUBS 0.007399f
C181 B.n141 VSUBS 0.007399f
C182 B.n142 VSUBS 0.007399f
C183 B.n143 VSUBS 0.007399f
C184 B.n144 VSUBS 0.007399f
C185 B.n145 VSUBS 0.007399f
C186 B.n146 VSUBS 0.007399f
C187 B.n147 VSUBS 0.007399f
C188 B.n148 VSUBS 0.007399f
C189 B.n149 VSUBS 0.007399f
C190 B.n150 VSUBS 0.007399f
C191 B.n151 VSUBS 0.007399f
C192 B.n152 VSUBS 0.007399f
C193 B.n153 VSUBS 0.007399f
C194 B.n154 VSUBS 0.007399f
C195 B.n155 VSUBS 0.007399f
C196 B.n156 VSUBS 0.007399f
C197 B.n157 VSUBS 0.007399f
C198 B.n158 VSUBS 0.007399f
C199 B.n159 VSUBS 0.007399f
C200 B.n160 VSUBS 0.007399f
C201 B.n161 VSUBS 0.007399f
C202 B.n162 VSUBS 0.007399f
C203 B.n163 VSUBS 0.007399f
C204 B.n164 VSUBS 0.007399f
C205 B.n165 VSUBS 0.007399f
C206 B.n166 VSUBS 0.007399f
C207 B.n167 VSUBS 0.007399f
C208 B.n168 VSUBS 0.007399f
C209 B.n169 VSUBS 0.007399f
C210 B.n170 VSUBS 0.017539f
C211 B.n171 VSUBS 0.017539f
C212 B.n172 VSUBS 0.018366f
C213 B.n173 VSUBS 0.007399f
C214 B.n174 VSUBS 0.007399f
C215 B.n175 VSUBS 0.007399f
C216 B.n176 VSUBS 0.007399f
C217 B.n177 VSUBS 0.007399f
C218 B.n178 VSUBS 0.007399f
C219 B.n179 VSUBS 0.007399f
C220 B.n180 VSUBS 0.007399f
C221 B.n181 VSUBS 0.007399f
C222 B.n182 VSUBS 0.007399f
C223 B.n183 VSUBS 0.007399f
C224 B.n184 VSUBS 0.007399f
C225 B.n185 VSUBS 0.007399f
C226 B.n186 VSUBS 0.007399f
C227 B.n187 VSUBS 0.007399f
C228 B.n188 VSUBS 0.007399f
C229 B.n189 VSUBS 0.007399f
C230 B.n190 VSUBS 0.007399f
C231 B.n191 VSUBS 0.007399f
C232 B.n192 VSUBS 0.007399f
C233 B.n193 VSUBS 0.007399f
C234 B.n194 VSUBS 0.007399f
C235 B.n195 VSUBS 0.007399f
C236 B.n196 VSUBS 0.007399f
C237 B.n197 VSUBS 0.007399f
C238 B.n198 VSUBS 0.007399f
C239 B.n199 VSUBS 0.007399f
C240 B.n200 VSUBS 0.007399f
C241 B.n201 VSUBS 0.007399f
C242 B.n202 VSUBS 0.007399f
C243 B.n203 VSUBS 0.007399f
C244 B.n204 VSUBS 0.007399f
C245 B.n205 VSUBS 0.007399f
C246 B.n206 VSUBS 0.007399f
C247 B.n207 VSUBS 0.007399f
C248 B.n208 VSUBS 0.007399f
C249 B.n209 VSUBS 0.007399f
C250 B.n210 VSUBS 0.007399f
C251 B.n211 VSUBS 0.007399f
C252 B.n212 VSUBS 0.007399f
C253 B.n213 VSUBS 0.007399f
C254 B.n214 VSUBS 0.007399f
C255 B.n215 VSUBS 0.007399f
C256 B.n216 VSUBS 0.007399f
C257 B.n217 VSUBS 0.007399f
C258 B.n218 VSUBS 0.007399f
C259 B.n219 VSUBS 0.007399f
C260 B.n220 VSUBS 0.007399f
C261 B.n221 VSUBS 0.006963f
C262 B.n222 VSUBS 0.007399f
C263 B.n223 VSUBS 0.007399f
C264 B.n224 VSUBS 0.004135f
C265 B.n225 VSUBS 0.007399f
C266 B.n226 VSUBS 0.007399f
C267 B.n227 VSUBS 0.007399f
C268 B.n228 VSUBS 0.007399f
C269 B.n229 VSUBS 0.007399f
C270 B.n230 VSUBS 0.007399f
C271 B.n231 VSUBS 0.007399f
C272 B.n232 VSUBS 0.007399f
C273 B.n233 VSUBS 0.007399f
C274 B.n234 VSUBS 0.007399f
C275 B.n235 VSUBS 0.007399f
C276 B.n236 VSUBS 0.007399f
C277 B.n237 VSUBS 0.004135f
C278 B.n238 VSUBS 0.017142f
C279 B.n239 VSUBS 0.006963f
C280 B.n240 VSUBS 0.007399f
C281 B.n241 VSUBS 0.007399f
C282 B.n242 VSUBS 0.007399f
C283 B.n243 VSUBS 0.007399f
C284 B.n244 VSUBS 0.007399f
C285 B.n245 VSUBS 0.007399f
C286 B.n246 VSUBS 0.007399f
C287 B.n247 VSUBS 0.007399f
C288 B.n248 VSUBS 0.007399f
C289 B.n249 VSUBS 0.007399f
C290 B.n250 VSUBS 0.007399f
C291 B.n251 VSUBS 0.007399f
C292 B.n252 VSUBS 0.007399f
C293 B.n253 VSUBS 0.007399f
C294 B.n254 VSUBS 0.007399f
C295 B.n255 VSUBS 0.007399f
C296 B.n256 VSUBS 0.007399f
C297 B.n257 VSUBS 0.007399f
C298 B.n258 VSUBS 0.007399f
C299 B.n259 VSUBS 0.007399f
C300 B.n260 VSUBS 0.007399f
C301 B.n261 VSUBS 0.007399f
C302 B.n262 VSUBS 0.007399f
C303 B.n263 VSUBS 0.007399f
C304 B.n264 VSUBS 0.007399f
C305 B.n265 VSUBS 0.007399f
C306 B.n266 VSUBS 0.007399f
C307 B.n267 VSUBS 0.007399f
C308 B.n268 VSUBS 0.007399f
C309 B.n269 VSUBS 0.007399f
C310 B.n270 VSUBS 0.007399f
C311 B.n271 VSUBS 0.007399f
C312 B.n272 VSUBS 0.007399f
C313 B.n273 VSUBS 0.007399f
C314 B.n274 VSUBS 0.007399f
C315 B.n275 VSUBS 0.007399f
C316 B.n276 VSUBS 0.007399f
C317 B.n277 VSUBS 0.007399f
C318 B.n278 VSUBS 0.007399f
C319 B.n279 VSUBS 0.007399f
C320 B.n280 VSUBS 0.007399f
C321 B.n281 VSUBS 0.007399f
C322 B.n282 VSUBS 0.007399f
C323 B.n283 VSUBS 0.007399f
C324 B.n284 VSUBS 0.007399f
C325 B.n285 VSUBS 0.007399f
C326 B.n286 VSUBS 0.007399f
C327 B.n287 VSUBS 0.007399f
C328 B.n288 VSUBS 0.007399f
C329 B.n289 VSUBS 0.018366f
C330 B.n290 VSUBS 0.017539f
C331 B.n291 VSUBS 0.017539f
C332 B.n292 VSUBS 0.007399f
C333 B.n293 VSUBS 0.007399f
C334 B.n294 VSUBS 0.007399f
C335 B.n295 VSUBS 0.007399f
C336 B.n296 VSUBS 0.007399f
C337 B.n297 VSUBS 0.007399f
C338 B.n298 VSUBS 0.007399f
C339 B.n299 VSUBS 0.007399f
C340 B.n300 VSUBS 0.007399f
C341 B.n301 VSUBS 0.007399f
C342 B.n302 VSUBS 0.007399f
C343 B.n303 VSUBS 0.007399f
C344 B.n304 VSUBS 0.007399f
C345 B.n305 VSUBS 0.007399f
C346 B.n306 VSUBS 0.007399f
C347 B.n307 VSUBS 0.007399f
C348 B.n308 VSUBS 0.007399f
C349 B.n309 VSUBS 0.007399f
C350 B.n310 VSUBS 0.007399f
C351 B.n311 VSUBS 0.007399f
C352 B.n312 VSUBS 0.007399f
C353 B.n313 VSUBS 0.007399f
C354 B.n314 VSUBS 0.007399f
C355 B.n315 VSUBS 0.007399f
C356 B.n316 VSUBS 0.007399f
C357 B.n317 VSUBS 0.007399f
C358 B.n318 VSUBS 0.007399f
C359 B.n319 VSUBS 0.007399f
C360 B.n320 VSUBS 0.007399f
C361 B.n321 VSUBS 0.007399f
C362 B.n322 VSUBS 0.007399f
C363 B.n323 VSUBS 0.007399f
C364 B.n324 VSUBS 0.007399f
C365 B.n325 VSUBS 0.007399f
C366 B.n326 VSUBS 0.007399f
C367 B.n327 VSUBS 0.007399f
C368 B.n328 VSUBS 0.007399f
C369 B.n329 VSUBS 0.007399f
C370 B.n330 VSUBS 0.007399f
C371 B.n331 VSUBS 0.007399f
C372 B.n332 VSUBS 0.007399f
C373 B.n333 VSUBS 0.007399f
C374 B.n334 VSUBS 0.007399f
C375 B.n335 VSUBS 0.007399f
C376 B.n336 VSUBS 0.007399f
C377 B.n337 VSUBS 0.007399f
C378 B.n338 VSUBS 0.007399f
C379 B.n339 VSUBS 0.007399f
C380 B.n340 VSUBS 0.007399f
C381 B.n341 VSUBS 0.007399f
C382 B.n342 VSUBS 0.007399f
C383 B.n343 VSUBS 0.007399f
C384 B.n344 VSUBS 0.007399f
C385 B.n345 VSUBS 0.007399f
C386 B.n346 VSUBS 0.007399f
C387 B.n347 VSUBS 0.007399f
C388 B.n348 VSUBS 0.007399f
C389 B.n349 VSUBS 0.007399f
C390 B.n350 VSUBS 0.007399f
C391 B.n351 VSUBS 0.007399f
C392 B.n352 VSUBS 0.007399f
C393 B.n353 VSUBS 0.007399f
C394 B.n354 VSUBS 0.007399f
C395 B.n355 VSUBS 0.007399f
C396 B.n356 VSUBS 0.007399f
C397 B.n357 VSUBS 0.007399f
C398 B.n358 VSUBS 0.007399f
C399 B.n359 VSUBS 0.007399f
C400 B.n360 VSUBS 0.007399f
C401 B.n361 VSUBS 0.007399f
C402 B.n362 VSUBS 0.017539f
C403 B.n363 VSUBS 0.018366f
C404 B.n364 VSUBS 0.017539f
C405 B.n365 VSUBS 0.007399f
C406 B.n366 VSUBS 0.007399f
C407 B.n367 VSUBS 0.007399f
C408 B.n368 VSUBS 0.007399f
C409 B.n369 VSUBS 0.007399f
C410 B.n370 VSUBS 0.007399f
C411 B.n371 VSUBS 0.007399f
C412 B.n372 VSUBS 0.007399f
C413 B.n373 VSUBS 0.007399f
C414 B.n374 VSUBS 0.007399f
C415 B.n375 VSUBS 0.007399f
C416 B.n376 VSUBS 0.007399f
C417 B.n377 VSUBS 0.007399f
C418 B.n378 VSUBS 0.007399f
C419 B.n379 VSUBS 0.007399f
C420 B.n380 VSUBS 0.007399f
C421 B.n381 VSUBS 0.007399f
C422 B.n382 VSUBS 0.007399f
C423 B.n383 VSUBS 0.007399f
C424 B.n384 VSUBS 0.007399f
C425 B.n385 VSUBS 0.007399f
C426 B.n386 VSUBS 0.007399f
C427 B.n387 VSUBS 0.007399f
C428 B.n388 VSUBS 0.007399f
C429 B.n389 VSUBS 0.007399f
C430 B.n390 VSUBS 0.007399f
C431 B.n391 VSUBS 0.007399f
C432 B.n392 VSUBS 0.007399f
C433 B.n393 VSUBS 0.007399f
C434 B.n394 VSUBS 0.007399f
C435 B.n395 VSUBS 0.007399f
C436 B.n396 VSUBS 0.007399f
C437 B.n397 VSUBS 0.007399f
C438 B.n398 VSUBS 0.007399f
C439 B.n399 VSUBS 0.007399f
C440 B.n400 VSUBS 0.007399f
C441 B.n401 VSUBS 0.007399f
C442 B.n402 VSUBS 0.007399f
C443 B.n403 VSUBS 0.007399f
C444 B.n404 VSUBS 0.007399f
C445 B.n405 VSUBS 0.007399f
C446 B.n406 VSUBS 0.007399f
C447 B.n407 VSUBS 0.007399f
C448 B.n408 VSUBS 0.007399f
C449 B.n409 VSUBS 0.007399f
C450 B.n410 VSUBS 0.007399f
C451 B.n411 VSUBS 0.007399f
C452 B.n412 VSUBS 0.007399f
C453 B.n413 VSUBS 0.006963f
C454 B.n414 VSUBS 0.007399f
C455 B.n415 VSUBS 0.007399f
C456 B.n416 VSUBS 0.004135f
C457 B.n417 VSUBS 0.007399f
C458 B.n418 VSUBS 0.007399f
C459 B.n419 VSUBS 0.007399f
C460 B.n420 VSUBS 0.007399f
C461 B.n421 VSUBS 0.007399f
C462 B.n422 VSUBS 0.007399f
C463 B.n423 VSUBS 0.007399f
C464 B.n424 VSUBS 0.007399f
C465 B.n425 VSUBS 0.007399f
C466 B.n426 VSUBS 0.007399f
C467 B.n427 VSUBS 0.007399f
C468 B.n428 VSUBS 0.007399f
C469 B.n429 VSUBS 0.004135f
C470 B.n430 VSUBS 0.017142f
C471 B.n431 VSUBS 0.006963f
C472 B.n432 VSUBS 0.007399f
C473 B.n433 VSUBS 0.007399f
C474 B.n434 VSUBS 0.007399f
C475 B.n435 VSUBS 0.007399f
C476 B.n436 VSUBS 0.007399f
C477 B.n437 VSUBS 0.007399f
C478 B.n438 VSUBS 0.007399f
C479 B.n439 VSUBS 0.007399f
C480 B.n440 VSUBS 0.007399f
C481 B.n441 VSUBS 0.007399f
C482 B.n442 VSUBS 0.007399f
C483 B.n443 VSUBS 0.007399f
C484 B.n444 VSUBS 0.007399f
C485 B.n445 VSUBS 0.007399f
C486 B.n446 VSUBS 0.007399f
C487 B.n447 VSUBS 0.007399f
C488 B.n448 VSUBS 0.007399f
C489 B.n449 VSUBS 0.007399f
C490 B.n450 VSUBS 0.007399f
C491 B.n451 VSUBS 0.007399f
C492 B.n452 VSUBS 0.007399f
C493 B.n453 VSUBS 0.007399f
C494 B.n454 VSUBS 0.007399f
C495 B.n455 VSUBS 0.007399f
C496 B.n456 VSUBS 0.007399f
C497 B.n457 VSUBS 0.007399f
C498 B.n458 VSUBS 0.007399f
C499 B.n459 VSUBS 0.007399f
C500 B.n460 VSUBS 0.007399f
C501 B.n461 VSUBS 0.007399f
C502 B.n462 VSUBS 0.007399f
C503 B.n463 VSUBS 0.007399f
C504 B.n464 VSUBS 0.007399f
C505 B.n465 VSUBS 0.007399f
C506 B.n466 VSUBS 0.007399f
C507 B.n467 VSUBS 0.007399f
C508 B.n468 VSUBS 0.007399f
C509 B.n469 VSUBS 0.007399f
C510 B.n470 VSUBS 0.007399f
C511 B.n471 VSUBS 0.007399f
C512 B.n472 VSUBS 0.007399f
C513 B.n473 VSUBS 0.007399f
C514 B.n474 VSUBS 0.007399f
C515 B.n475 VSUBS 0.007399f
C516 B.n476 VSUBS 0.007399f
C517 B.n477 VSUBS 0.007399f
C518 B.n478 VSUBS 0.007399f
C519 B.n479 VSUBS 0.007399f
C520 B.n480 VSUBS 0.007399f
C521 B.n481 VSUBS 0.018366f
C522 B.n482 VSUBS 0.017539f
C523 B.n483 VSUBS 0.017539f
C524 B.n484 VSUBS 0.007399f
C525 B.n485 VSUBS 0.007399f
C526 B.n486 VSUBS 0.007399f
C527 B.n487 VSUBS 0.007399f
C528 B.n488 VSUBS 0.007399f
C529 B.n489 VSUBS 0.007399f
C530 B.n490 VSUBS 0.007399f
C531 B.n491 VSUBS 0.007399f
C532 B.n492 VSUBS 0.007399f
C533 B.n493 VSUBS 0.007399f
C534 B.n494 VSUBS 0.007399f
C535 B.n495 VSUBS 0.007399f
C536 B.n496 VSUBS 0.007399f
C537 B.n497 VSUBS 0.007399f
C538 B.n498 VSUBS 0.007399f
C539 B.n499 VSUBS 0.007399f
C540 B.n500 VSUBS 0.007399f
C541 B.n501 VSUBS 0.007399f
C542 B.n502 VSUBS 0.007399f
C543 B.n503 VSUBS 0.007399f
C544 B.n504 VSUBS 0.007399f
C545 B.n505 VSUBS 0.007399f
C546 B.n506 VSUBS 0.007399f
C547 B.n507 VSUBS 0.007399f
C548 B.n508 VSUBS 0.007399f
C549 B.n509 VSUBS 0.007399f
C550 B.n510 VSUBS 0.007399f
C551 B.n511 VSUBS 0.007399f
C552 B.n512 VSUBS 0.007399f
C553 B.n513 VSUBS 0.007399f
C554 B.n514 VSUBS 0.007399f
C555 B.n515 VSUBS 0.007399f
C556 B.n516 VSUBS 0.007399f
C557 B.n517 VSUBS 0.007399f
C558 B.n518 VSUBS 0.007399f
C559 B.n519 VSUBS 0.016753f
C560 VDD2.n0 VSUBS 0.025646f
C561 VDD2.n1 VSUBS 0.022472f
C562 VDD2.n2 VSUBS 0.012076f
C563 VDD2.n3 VSUBS 0.028542f
C564 VDD2.n4 VSUBS 0.012786f
C565 VDD2.n5 VSUBS 0.022472f
C566 VDD2.n6 VSUBS 0.012076f
C567 VDD2.n7 VSUBS 0.028542f
C568 VDD2.n8 VSUBS 0.012786f
C569 VDD2.n9 VSUBS 0.022472f
C570 VDD2.n10 VSUBS 0.012076f
C571 VDD2.n11 VSUBS 0.028542f
C572 VDD2.n12 VSUBS 0.012786f
C573 VDD2.n13 VSUBS 0.022472f
C574 VDD2.n14 VSUBS 0.012076f
C575 VDD2.n15 VSUBS 0.021407f
C576 VDD2.n16 VSUBS 0.018157f
C577 VDD2.t4 VSUBS 0.060852f
C578 VDD2.n17 VSUBS 0.122076f
C579 VDD2.n18 VSUBS 0.874707f
C580 VDD2.n19 VSUBS 0.012076f
C581 VDD2.n20 VSUBS 0.012786f
C582 VDD2.n21 VSUBS 0.028542f
C583 VDD2.n22 VSUBS 0.028542f
C584 VDD2.n23 VSUBS 0.012786f
C585 VDD2.n24 VSUBS 0.012076f
C586 VDD2.n25 VSUBS 0.022472f
C587 VDD2.n26 VSUBS 0.022472f
C588 VDD2.n27 VSUBS 0.012076f
C589 VDD2.n28 VSUBS 0.012786f
C590 VDD2.n29 VSUBS 0.028542f
C591 VDD2.n30 VSUBS 0.028542f
C592 VDD2.n31 VSUBS 0.012786f
C593 VDD2.n32 VSUBS 0.012076f
C594 VDD2.n33 VSUBS 0.022472f
C595 VDD2.n34 VSUBS 0.022472f
C596 VDD2.n35 VSUBS 0.012076f
C597 VDD2.n36 VSUBS 0.012786f
C598 VDD2.n37 VSUBS 0.028542f
C599 VDD2.n38 VSUBS 0.028542f
C600 VDD2.n39 VSUBS 0.012786f
C601 VDD2.n40 VSUBS 0.012076f
C602 VDD2.n41 VSUBS 0.022472f
C603 VDD2.n42 VSUBS 0.022472f
C604 VDD2.n43 VSUBS 0.012076f
C605 VDD2.n44 VSUBS 0.012786f
C606 VDD2.n45 VSUBS 0.028542f
C607 VDD2.n46 VSUBS 0.072347f
C608 VDD2.n47 VSUBS 0.012786f
C609 VDD2.n48 VSUBS 0.012076f
C610 VDD2.n49 VSUBS 0.049181f
C611 VDD2.n50 VSUBS 0.053733f
C612 VDD2.t5 VSUBS 0.16888f
C613 VDD2.t3 VSUBS 0.16888f
C614 VDD2.n51 VSUBS 1.24868f
C615 VDD2.n52 VSUBS 1.88928f
C616 VDD2.n53 VSUBS 0.025646f
C617 VDD2.n54 VSUBS 0.022472f
C618 VDD2.n55 VSUBS 0.012076f
C619 VDD2.n56 VSUBS 0.028542f
C620 VDD2.n57 VSUBS 0.012786f
C621 VDD2.n58 VSUBS 0.022472f
C622 VDD2.n59 VSUBS 0.012076f
C623 VDD2.n60 VSUBS 0.028542f
C624 VDD2.n61 VSUBS 0.012786f
C625 VDD2.n62 VSUBS 0.022472f
C626 VDD2.n63 VSUBS 0.012076f
C627 VDD2.n64 VSUBS 0.028542f
C628 VDD2.n65 VSUBS 0.012786f
C629 VDD2.n66 VSUBS 0.022472f
C630 VDD2.n67 VSUBS 0.012076f
C631 VDD2.n68 VSUBS 0.021407f
C632 VDD2.n69 VSUBS 0.018157f
C633 VDD2.t1 VSUBS 0.060852f
C634 VDD2.n70 VSUBS 0.122076f
C635 VDD2.n71 VSUBS 0.874707f
C636 VDD2.n72 VSUBS 0.012076f
C637 VDD2.n73 VSUBS 0.012786f
C638 VDD2.n74 VSUBS 0.028542f
C639 VDD2.n75 VSUBS 0.028542f
C640 VDD2.n76 VSUBS 0.012786f
C641 VDD2.n77 VSUBS 0.012076f
C642 VDD2.n78 VSUBS 0.022472f
C643 VDD2.n79 VSUBS 0.022472f
C644 VDD2.n80 VSUBS 0.012076f
C645 VDD2.n81 VSUBS 0.012786f
C646 VDD2.n82 VSUBS 0.028542f
C647 VDD2.n83 VSUBS 0.028542f
C648 VDD2.n84 VSUBS 0.012786f
C649 VDD2.n85 VSUBS 0.012076f
C650 VDD2.n86 VSUBS 0.022472f
C651 VDD2.n87 VSUBS 0.022472f
C652 VDD2.n88 VSUBS 0.012076f
C653 VDD2.n89 VSUBS 0.012786f
C654 VDD2.n90 VSUBS 0.028542f
C655 VDD2.n91 VSUBS 0.028542f
C656 VDD2.n92 VSUBS 0.012786f
C657 VDD2.n93 VSUBS 0.012076f
C658 VDD2.n94 VSUBS 0.022472f
C659 VDD2.n95 VSUBS 0.022472f
C660 VDD2.n96 VSUBS 0.012076f
C661 VDD2.n97 VSUBS 0.012786f
C662 VDD2.n98 VSUBS 0.028542f
C663 VDD2.n99 VSUBS 0.072347f
C664 VDD2.n100 VSUBS 0.012786f
C665 VDD2.n101 VSUBS 0.012076f
C666 VDD2.n102 VSUBS 0.049181f
C667 VDD2.n103 VSUBS 0.05198f
C668 VDD2.n104 VSUBS 1.74072f
C669 VDD2.t0 VSUBS 0.16888f
C670 VDD2.t2 VSUBS 0.16888f
C671 VDD2.n105 VSUBS 1.24866f
C672 VN.n0 VSUBS 0.272903f
C673 VN.t0 VSUBS 1.32854f
C674 VN.t1 VSUBS 1.45508f
C675 VN.n1 VSUBS 0.566145f
C676 VN.n2 VSUBS 0.58401f
C677 VN.n3 VSUBS 0.060121f
C678 VN.t2 VSUBS 1.40768f
C679 VN.n4 VSUBS 0.582656f
C680 VN.n5 VSUBS 0.046972f
C681 VN.n6 VSUBS 0.272903f
C682 VN.t5 VSUBS 1.32854f
C683 VN.t3 VSUBS 1.45508f
C684 VN.n7 VSUBS 0.566145f
C685 VN.n8 VSUBS 0.58401f
C686 VN.n9 VSUBS 0.060121f
C687 VN.t4 VSUBS 1.40768f
C688 VN.n10 VSUBS 0.582656f
C689 VN.n11 VSUBS 2.01378f
C690 VTAIL.t0 VSUBS 0.21909f
C691 VTAIL.t2 VSUBS 0.21909f
C692 VTAIL.n0 VSUBS 1.47027f
C693 VTAIL.n1 VSUBS 0.781165f
C694 VTAIL.n2 VSUBS 0.033271f
C695 VTAIL.n3 VSUBS 0.029153f
C696 VTAIL.n4 VSUBS 0.015666f
C697 VTAIL.n5 VSUBS 0.037028f
C698 VTAIL.n6 VSUBS 0.016587f
C699 VTAIL.n7 VSUBS 0.029153f
C700 VTAIL.n8 VSUBS 0.015666f
C701 VTAIL.n9 VSUBS 0.037028f
C702 VTAIL.n10 VSUBS 0.016587f
C703 VTAIL.n11 VSUBS 0.029153f
C704 VTAIL.n12 VSUBS 0.015666f
C705 VTAIL.n13 VSUBS 0.037028f
C706 VTAIL.n14 VSUBS 0.016587f
C707 VTAIL.n15 VSUBS 0.029153f
C708 VTAIL.n16 VSUBS 0.015666f
C709 VTAIL.n17 VSUBS 0.027771f
C710 VTAIL.n18 VSUBS 0.023556f
C711 VTAIL.t7 VSUBS 0.078944f
C712 VTAIL.n19 VSUBS 0.15837f
C713 VTAIL.n20 VSUBS 1.13477f
C714 VTAIL.n21 VSUBS 0.015666f
C715 VTAIL.n22 VSUBS 0.016587f
C716 VTAIL.n23 VSUBS 0.037028f
C717 VTAIL.n24 VSUBS 0.037028f
C718 VTAIL.n25 VSUBS 0.016587f
C719 VTAIL.n26 VSUBS 0.015666f
C720 VTAIL.n27 VSUBS 0.029153f
C721 VTAIL.n28 VSUBS 0.029153f
C722 VTAIL.n29 VSUBS 0.015666f
C723 VTAIL.n30 VSUBS 0.016587f
C724 VTAIL.n31 VSUBS 0.037028f
C725 VTAIL.n32 VSUBS 0.037028f
C726 VTAIL.n33 VSUBS 0.016587f
C727 VTAIL.n34 VSUBS 0.015666f
C728 VTAIL.n35 VSUBS 0.029153f
C729 VTAIL.n36 VSUBS 0.029153f
C730 VTAIL.n37 VSUBS 0.015666f
C731 VTAIL.n38 VSUBS 0.016587f
C732 VTAIL.n39 VSUBS 0.037028f
C733 VTAIL.n40 VSUBS 0.037028f
C734 VTAIL.n41 VSUBS 0.016587f
C735 VTAIL.n42 VSUBS 0.015666f
C736 VTAIL.n43 VSUBS 0.029153f
C737 VTAIL.n44 VSUBS 0.029153f
C738 VTAIL.n45 VSUBS 0.015666f
C739 VTAIL.n46 VSUBS 0.016587f
C740 VTAIL.n47 VSUBS 0.037028f
C741 VTAIL.n48 VSUBS 0.093856f
C742 VTAIL.n49 VSUBS 0.016587f
C743 VTAIL.n50 VSUBS 0.015666f
C744 VTAIL.n51 VSUBS 0.063802f
C745 VTAIL.n52 VSUBS 0.047274f
C746 VTAIL.n53 VSUBS 0.232217f
C747 VTAIL.t10 VSUBS 0.21909f
C748 VTAIL.t9 VSUBS 0.21909f
C749 VTAIL.n54 VSUBS 1.47027f
C750 VTAIL.n55 VSUBS 2.14552f
C751 VTAIL.t3 VSUBS 0.21909f
C752 VTAIL.t1 VSUBS 0.21909f
C753 VTAIL.n56 VSUBS 1.47028f
C754 VTAIL.n57 VSUBS 2.14551f
C755 VTAIL.n58 VSUBS 0.033271f
C756 VTAIL.n59 VSUBS 0.029153f
C757 VTAIL.n60 VSUBS 0.015666f
C758 VTAIL.n61 VSUBS 0.037028f
C759 VTAIL.n62 VSUBS 0.016587f
C760 VTAIL.n63 VSUBS 0.029153f
C761 VTAIL.n64 VSUBS 0.015666f
C762 VTAIL.n65 VSUBS 0.037028f
C763 VTAIL.n66 VSUBS 0.016587f
C764 VTAIL.n67 VSUBS 0.029153f
C765 VTAIL.n68 VSUBS 0.015666f
C766 VTAIL.n69 VSUBS 0.037028f
C767 VTAIL.n70 VSUBS 0.016587f
C768 VTAIL.n71 VSUBS 0.029153f
C769 VTAIL.n72 VSUBS 0.015666f
C770 VTAIL.n73 VSUBS 0.027771f
C771 VTAIL.n74 VSUBS 0.023556f
C772 VTAIL.t5 VSUBS 0.078944f
C773 VTAIL.n75 VSUBS 0.15837f
C774 VTAIL.n76 VSUBS 1.13477f
C775 VTAIL.n77 VSUBS 0.015666f
C776 VTAIL.n78 VSUBS 0.016587f
C777 VTAIL.n79 VSUBS 0.037028f
C778 VTAIL.n80 VSUBS 0.037028f
C779 VTAIL.n81 VSUBS 0.016587f
C780 VTAIL.n82 VSUBS 0.015666f
C781 VTAIL.n83 VSUBS 0.029153f
C782 VTAIL.n84 VSUBS 0.029153f
C783 VTAIL.n85 VSUBS 0.015666f
C784 VTAIL.n86 VSUBS 0.016587f
C785 VTAIL.n87 VSUBS 0.037028f
C786 VTAIL.n88 VSUBS 0.037028f
C787 VTAIL.n89 VSUBS 0.016587f
C788 VTAIL.n90 VSUBS 0.015666f
C789 VTAIL.n91 VSUBS 0.029153f
C790 VTAIL.n92 VSUBS 0.029153f
C791 VTAIL.n93 VSUBS 0.015666f
C792 VTAIL.n94 VSUBS 0.016587f
C793 VTAIL.n95 VSUBS 0.037028f
C794 VTAIL.n96 VSUBS 0.037028f
C795 VTAIL.n97 VSUBS 0.016587f
C796 VTAIL.n98 VSUBS 0.015666f
C797 VTAIL.n99 VSUBS 0.029153f
C798 VTAIL.n100 VSUBS 0.029153f
C799 VTAIL.n101 VSUBS 0.015666f
C800 VTAIL.n102 VSUBS 0.016587f
C801 VTAIL.n103 VSUBS 0.037028f
C802 VTAIL.n104 VSUBS 0.093856f
C803 VTAIL.n105 VSUBS 0.016587f
C804 VTAIL.n106 VSUBS 0.015666f
C805 VTAIL.n107 VSUBS 0.063802f
C806 VTAIL.n108 VSUBS 0.047274f
C807 VTAIL.n109 VSUBS 0.232217f
C808 VTAIL.t8 VSUBS 0.21909f
C809 VTAIL.t11 VSUBS 0.21909f
C810 VTAIL.n110 VSUBS 1.47028f
C811 VTAIL.n111 VSUBS 0.858292f
C812 VTAIL.n112 VSUBS 0.033271f
C813 VTAIL.n113 VSUBS 0.029153f
C814 VTAIL.n114 VSUBS 0.015666f
C815 VTAIL.n115 VSUBS 0.037028f
C816 VTAIL.n116 VSUBS 0.016587f
C817 VTAIL.n117 VSUBS 0.029153f
C818 VTAIL.n118 VSUBS 0.015666f
C819 VTAIL.n119 VSUBS 0.037028f
C820 VTAIL.n120 VSUBS 0.016587f
C821 VTAIL.n121 VSUBS 0.029153f
C822 VTAIL.n122 VSUBS 0.015666f
C823 VTAIL.n123 VSUBS 0.037028f
C824 VTAIL.n124 VSUBS 0.016587f
C825 VTAIL.n125 VSUBS 0.029153f
C826 VTAIL.n126 VSUBS 0.015666f
C827 VTAIL.n127 VSUBS 0.027771f
C828 VTAIL.n128 VSUBS 0.023556f
C829 VTAIL.t6 VSUBS 0.078944f
C830 VTAIL.n129 VSUBS 0.15837f
C831 VTAIL.n130 VSUBS 1.13477f
C832 VTAIL.n131 VSUBS 0.015666f
C833 VTAIL.n132 VSUBS 0.016587f
C834 VTAIL.n133 VSUBS 0.037028f
C835 VTAIL.n134 VSUBS 0.037028f
C836 VTAIL.n135 VSUBS 0.016587f
C837 VTAIL.n136 VSUBS 0.015666f
C838 VTAIL.n137 VSUBS 0.029153f
C839 VTAIL.n138 VSUBS 0.029153f
C840 VTAIL.n139 VSUBS 0.015666f
C841 VTAIL.n140 VSUBS 0.016587f
C842 VTAIL.n141 VSUBS 0.037028f
C843 VTAIL.n142 VSUBS 0.037028f
C844 VTAIL.n143 VSUBS 0.016587f
C845 VTAIL.n144 VSUBS 0.015666f
C846 VTAIL.n145 VSUBS 0.029153f
C847 VTAIL.n146 VSUBS 0.029153f
C848 VTAIL.n147 VSUBS 0.015666f
C849 VTAIL.n148 VSUBS 0.016587f
C850 VTAIL.n149 VSUBS 0.037028f
C851 VTAIL.n150 VSUBS 0.037028f
C852 VTAIL.n151 VSUBS 0.016587f
C853 VTAIL.n152 VSUBS 0.015666f
C854 VTAIL.n153 VSUBS 0.029153f
C855 VTAIL.n154 VSUBS 0.029153f
C856 VTAIL.n155 VSUBS 0.015666f
C857 VTAIL.n156 VSUBS 0.016587f
C858 VTAIL.n157 VSUBS 0.037028f
C859 VTAIL.n158 VSUBS 0.093856f
C860 VTAIL.n159 VSUBS 0.016587f
C861 VTAIL.n160 VSUBS 0.015666f
C862 VTAIL.n161 VSUBS 0.063802f
C863 VTAIL.n162 VSUBS 0.047274f
C864 VTAIL.n163 VSUBS 1.4093f
C865 VTAIL.n164 VSUBS 0.033271f
C866 VTAIL.n165 VSUBS 0.029153f
C867 VTAIL.n166 VSUBS 0.015666f
C868 VTAIL.n167 VSUBS 0.037028f
C869 VTAIL.n168 VSUBS 0.016587f
C870 VTAIL.n169 VSUBS 0.029153f
C871 VTAIL.n170 VSUBS 0.015666f
C872 VTAIL.n171 VSUBS 0.037028f
C873 VTAIL.n172 VSUBS 0.016587f
C874 VTAIL.n173 VSUBS 0.029153f
C875 VTAIL.n174 VSUBS 0.015666f
C876 VTAIL.n175 VSUBS 0.037028f
C877 VTAIL.n176 VSUBS 0.016587f
C878 VTAIL.n177 VSUBS 0.029153f
C879 VTAIL.n178 VSUBS 0.015666f
C880 VTAIL.n179 VSUBS 0.027771f
C881 VTAIL.n180 VSUBS 0.023556f
C882 VTAIL.t4 VSUBS 0.078944f
C883 VTAIL.n181 VSUBS 0.15837f
C884 VTAIL.n182 VSUBS 1.13477f
C885 VTAIL.n183 VSUBS 0.015666f
C886 VTAIL.n184 VSUBS 0.016587f
C887 VTAIL.n185 VSUBS 0.037028f
C888 VTAIL.n186 VSUBS 0.037028f
C889 VTAIL.n187 VSUBS 0.016587f
C890 VTAIL.n188 VSUBS 0.015666f
C891 VTAIL.n189 VSUBS 0.029153f
C892 VTAIL.n190 VSUBS 0.029153f
C893 VTAIL.n191 VSUBS 0.015666f
C894 VTAIL.n192 VSUBS 0.016587f
C895 VTAIL.n193 VSUBS 0.037028f
C896 VTAIL.n194 VSUBS 0.037028f
C897 VTAIL.n195 VSUBS 0.016587f
C898 VTAIL.n196 VSUBS 0.015666f
C899 VTAIL.n197 VSUBS 0.029153f
C900 VTAIL.n198 VSUBS 0.029153f
C901 VTAIL.n199 VSUBS 0.015666f
C902 VTAIL.n200 VSUBS 0.016587f
C903 VTAIL.n201 VSUBS 0.037028f
C904 VTAIL.n202 VSUBS 0.037028f
C905 VTAIL.n203 VSUBS 0.016587f
C906 VTAIL.n204 VSUBS 0.015666f
C907 VTAIL.n205 VSUBS 0.029153f
C908 VTAIL.n206 VSUBS 0.029153f
C909 VTAIL.n207 VSUBS 0.015666f
C910 VTAIL.n208 VSUBS 0.016587f
C911 VTAIL.n209 VSUBS 0.037028f
C912 VTAIL.n210 VSUBS 0.093856f
C913 VTAIL.n211 VSUBS 0.016587f
C914 VTAIL.n212 VSUBS 0.015666f
C915 VTAIL.n213 VSUBS 0.063802f
C916 VTAIL.n214 VSUBS 0.047274f
C917 VTAIL.n215 VSUBS 1.3763f
C918 VDD1.n0 VSUBS 0.025683f
C919 VDD1.n1 VSUBS 0.022505f
C920 VDD1.n2 VSUBS 0.012093f
C921 VDD1.n3 VSUBS 0.028584f
C922 VDD1.n4 VSUBS 0.012804f
C923 VDD1.n5 VSUBS 0.022505f
C924 VDD1.n6 VSUBS 0.012093f
C925 VDD1.n7 VSUBS 0.028584f
C926 VDD1.n8 VSUBS 0.012804f
C927 VDD1.n9 VSUBS 0.022505f
C928 VDD1.n10 VSUBS 0.012093f
C929 VDD1.n11 VSUBS 0.028584f
C930 VDD1.n12 VSUBS 0.012804f
C931 VDD1.n13 VSUBS 0.022505f
C932 VDD1.n14 VSUBS 0.012093f
C933 VDD1.n15 VSUBS 0.021438f
C934 VDD1.n16 VSUBS 0.018184f
C935 VDD1.t5 VSUBS 0.060941f
C936 VDD1.n17 VSUBS 0.122253f
C937 VDD1.n18 VSUBS 0.87598f
C938 VDD1.n19 VSUBS 0.012093f
C939 VDD1.n20 VSUBS 0.012804f
C940 VDD1.n21 VSUBS 0.028584f
C941 VDD1.n22 VSUBS 0.028584f
C942 VDD1.n23 VSUBS 0.012804f
C943 VDD1.n24 VSUBS 0.012093f
C944 VDD1.n25 VSUBS 0.022505f
C945 VDD1.n26 VSUBS 0.022505f
C946 VDD1.n27 VSUBS 0.012093f
C947 VDD1.n28 VSUBS 0.012804f
C948 VDD1.n29 VSUBS 0.028584f
C949 VDD1.n30 VSUBS 0.028584f
C950 VDD1.n31 VSUBS 0.012804f
C951 VDD1.n32 VSUBS 0.012093f
C952 VDD1.n33 VSUBS 0.022505f
C953 VDD1.n34 VSUBS 0.022505f
C954 VDD1.n35 VSUBS 0.012093f
C955 VDD1.n36 VSUBS 0.012804f
C956 VDD1.n37 VSUBS 0.028584f
C957 VDD1.n38 VSUBS 0.028584f
C958 VDD1.n39 VSUBS 0.012804f
C959 VDD1.n40 VSUBS 0.012093f
C960 VDD1.n41 VSUBS 0.022505f
C961 VDD1.n42 VSUBS 0.022505f
C962 VDD1.n43 VSUBS 0.012093f
C963 VDD1.n44 VSUBS 0.012804f
C964 VDD1.n45 VSUBS 0.028584f
C965 VDD1.n46 VSUBS 0.072452f
C966 VDD1.n47 VSUBS 0.012804f
C967 VDD1.n48 VSUBS 0.012093f
C968 VDD1.n49 VSUBS 0.049252f
C969 VDD1.n50 VSUBS 0.054196f
C970 VDD1.n51 VSUBS 0.025683f
C971 VDD1.n52 VSUBS 0.022505f
C972 VDD1.n53 VSUBS 0.012093f
C973 VDD1.n54 VSUBS 0.028584f
C974 VDD1.n55 VSUBS 0.012804f
C975 VDD1.n56 VSUBS 0.022505f
C976 VDD1.n57 VSUBS 0.012093f
C977 VDD1.n58 VSUBS 0.028584f
C978 VDD1.n59 VSUBS 0.012804f
C979 VDD1.n60 VSUBS 0.022505f
C980 VDD1.n61 VSUBS 0.012093f
C981 VDD1.n62 VSUBS 0.028584f
C982 VDD1.n63 VSUBS 0.012804f
C983 VDD1.n64 VSUBS 0.022505f
C984 VDD1.n65 VSUBS 0.012093f
C985 VDD1.n66 VSUBS 0.021438f
C986 VDD1.n67 VSUBS 0.018184f
C987 VDD1.t3 VSUBS 0.060941f
C988 VDD1.n68 VSUBS 0.122253f
C989 VDD1.n69 VSUBS 0.87598f
C990 VDD1.n70 VSUBS 0.012093f
C991 VDD1.n71 VSUBS 0.012804f
C992 VDD1.n72 VSUBS 0.028584f
C993 VDD1.n73 VSUBS 0.028584f
C994 VDD1.n74 VSUBS 0.012804f
C995 VDD1.n75 VSUBS 0.012093f
C996 VDD1.n76 VSUBS 0.022505f
C997 VDD1.n77 VSUBS 0.022505f
C998 VDD1.n78 VSUBS 0.012093f
C999 VDD1.n79 VSUBS 0.012804f
C1000 VDD1.n80 VSUBS 0.028584f
C1001 VDD1.n81 VSUBS 0.028584f
C1002 VDD1.n82 VSUBS 0.012804f
C1003 VDD1.n83 VSUBS 0.012093f
C1004 VDD1.n84 VSUBS 0.022505f
C1005 VDD1.n85 VSUBS 0.022505f
C1006 VDD1.n86 VSUBS 0.012093f
C1007 VDD1.n87 VSUBS 0.012804f
C1008 VDD1.n88 VSUBS 0.028584f
C1009 VDD1.n89 VSUBS 0.028584f
C1010 VDD1.n90 VSUBS 0.012804f
C1011 VDD1.n91 VSUBS 0.012093f
C1012 VDD1.n92 VSUBS 0.022505f
C1013 VDD1.n93 VSUBS 0.022505f
C1014 VDD1.n94 VSUBS 0.012093f
C1015 VDD1.n95 VSUBS 0.012804f
C1016 VDD1.n96 VSUBS 0.028584f
C1017 VDD1.n97 VSUBS 0.072452f
C1018 VDD1.n98 VSUBS 0.012804f
C1019 VDD1.n99 VSUBS 0.012093f
C1020 VDD1.n100 VSUBS 0.049252f
C1021 VDD1.n101 VSUBS 0.053811f
C1022 VDD1.t2 VSUBS 0.169126f
C1023 VDD1.t0 VSUBS 0.169126f
C1024 VDD1.n102 VSUBS 1.25049f
C1025 VDD1.n103 VSUBS 1.96739f
C1026 VDD1.t4 VSUBS 0.169126f
C1027 VDD1.t1 VSUBS 0.169126f
C1028 VDD1.n104 VSUBS 1.24887f
C1029 VDD1.n105 VSUBS 2.17005f
C1030 VP.n0 VSUBS 0.068425f
C1031 VP.t2 VSUBS 1.35832f
C1032 VP.n1 VSUBS 0.061469f
C1033 VP.n2 VSUBS 0.27902f
C1034 VP.t5 VSUBS 1.43923f
C1035 VP.t0 VSUBS 1.35832f
C1036 VP.t3 VSUBS 1.4877f
C1037 VP.n3 VSUBS 0.578835f
C1038 VP.n4 VSUBS 0.597101f
C1039 VP.n5 VSUBS 0.061469f
C1040 VP.n6 VSUBS 0.595717f
C1041 VP.n7 VSUBS 2.02999f
C1042 VP.t1 VSUBS 1.43923f
C1043 VP.n8 VSUBS 0.595717f
C1044 VP.n9 VSUBS 2.07523f
C1045 VP.n10 VSUBS 0.068425f
C1046 VP.n11 VSUBS 0.051279f
C1047 VP.n12 VSUBS 0.56479f
C1048 VP.n13 VSUBS 0.061469f
C1049 VP.t4 VSUBS 1.43923f
C1050 VP.n14 VSUBS 0.595717f
C1051 VP.n15 VSUBS 0.048025f
.ends

