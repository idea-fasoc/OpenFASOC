* NGSPICE file created from diff_pair_sample_1735.ext - technology: sky130A

.subckt diff_pair_sample_1735 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t7 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X1 B.t11 B.t9 B.t10 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=2.06
X2 VTAIL.t6 VP.t0 VDD1.t7 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=2.06
X3 B.t8 B.t6 B.t7 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=2.06
X4 VTAIL.t14 VN.t1 VDD2.t1 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=2.06
X5 VTAIL.t13 VN.t2 VDD2.t3 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X6 VDD2.t6 VN.t3 VTAIL.t12 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=2.06
X7 VTAIL.t3 VP.t1 VDD1.t6 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=2.06
X8 VTAIL.t1 VP.t2 VDD1.t5 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X9 VTAIL.t2 VP.t3 VDD1.t4 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X10 VDD2.t4 VN.t4 VTAIL.t11 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X11 VDD2.t0 VN.t5 VTAIL.t10 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X12 VDD2.t2 VN.t6 VTAIL.t9 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=2.06
X13 VDD1.t3 VP.t4 VTAIL.t5 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X14 VDD1.t2 VP.t5 VTAIL.t0 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=1.848 ps=11.53 w=11.2 l=2.06
X15 VDD1.t1 VP.t6 VTAIL.t7 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=2.06
X16 B.t5 B.t3 B.t4 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=2.06
X17 B.t2 B.t0 B.t1 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=0 ps=0 w=11.2 l=2.06
X18 VDD1.t0 VP.t7 VTAIL.t4 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=1.848 pd=11.53 as=4.368 ps=23.18 w=11.2 l=2.06
X19 VTAIL.t8 VN.t7 VDD2.t5 w_n3360_n3208# sky130_fd_pr__pfet_01v8 ad=4.368 pd=23.18 as=1.848 ps=11.53 w=11.2 l=2.06
R0 VN.n5 VN.t7 164.535
R1 VN.n28 VN.t3 164.535
R2 VN.n43 VN.n23 161.3
R3 VN.n42 VN.n41 161.3
R4 VN.n40 VN.n24 161.3
R5 VN.n39 VN.n38 161.3
R6 VN.n37 VN.n25 161.3
R7 VN.n35 VN.n34 161.3
R8 VN.n33 VN.n26 161.3
R9 VN.n32 VN.n31 161.3
R10 VN.n30 VN.n27 161.3
R11 VN.n20 VN.n0 161.3
R12 VN.n19 VN.n18 161.3
R13 VN.n17 VN.n1 161.3
R14 VN.n16 VN.n15 161.3
R15 VN.n14 VN.n2 161.3
R16 VN.n12 VN.n11 161.3
R17 VN.n10 VN.n3 161.3
R18 VN.n9 VN.n8 161.3
R19 VN.n7 VN.n4 161.3
R20 VN.n6 VN.t4 131.03
R21 VN.n13 VN.t2 131.03
R22 VN.n21 VN.t6 131.03
R23 VN.n29 VN.t0 131.03
R24 VN.n36 VN.t5 131.03
R25 VN.n44 VN.t1 131.03
R26 VN.n22 VN.n21 94.4317
R27 VN.n45 VN.n44 94.4317
R28 VN.n8 VN.n3 56.5617
R29 VN.n31 VN.n26 56.5617
R30 VN.n19 VN.n1 54.1398
R31 VN.n42 VN.n24 54.1398
R32 VN.n6 VN.n5 48.8225
R33 VN.n29 VN.n28 48.8225
R34 VN VN.n45 48.0285
R35 VN.n15 VN.n1 27.0143
R36 VN.n38 VN.n24 27.0143
R37 VN.n8 VN.n7 24.5923
R38 VN.n12 VN.n3 24.5923
R39 VN.n15 VN.n14 24.5923
R40 VN.n20 VN.n19 24.5923
R41 VN.n31 VN.n30 24.5923
R42 VN.n38 VN.n37 24.5923
R43 VN.n35 VN.n26 24.5923
R44 VN.n43 VN.n42 24.5923
R45 VN.n7 VN.n6 21.8872
R46 VN.n13 VN.n12 21.8872
R47 VN.n30 VN.n29 21.8872
R48 VN.n36 VN.n35 21.8872
R49 VN.n21 VN.n20 16.477
R50 VN.n44 VN.n43 16.477
R51 VN.n28 VN.n27 9.28418
R52 VN.n5 VN.n4 9.28418
R53 VN.n14 VN.n13 2.7056
R54 VN.n37 VN.n36 2.7056
R55 VN.n45 VN.n23 0.278335
R56 VN.n22 VN.n0 0.278335
R57 VN.n41 VN.n23 0.189894
R58 VN.n41 VN.n40 0.189894
R59 VN.n40 VN.n39 0.189894
R60 VN.n39 VN.n25 0.189894
R61 VN.n34 VN.n25 0.189894
R62 VN.n34 VN.n33 0.189894
R63 VN.n33 VN.n32 0.189894
R64 VN.n32 VN.n27 0.189894
R65 VN.n9 VN.n4 0.189894
R66 VN.n10 VN.n9 0.189894
R67 VN.n11 VN.n10 0.189894
R68 VN.n11 VN.n2 0.189894
R69 VN.n16 VN.n2 0.189894
R70 VN.n17 VN.n16 0.189894
R71 VN.n18 VN.n17 0.189894
R72 VN.n18 VN.n0 0.189894
R73 VN VN.n22 0.153485
R74 VDD2.n2 VDD2.n1 79.3827
R75 VDD2.n2 VDD2.n0 79.3827
R76 VDD2 VDD2.n5 79.3799
R77 VDD2.n4 VDD2.n3 78.4081
R78 VDD2.n4 VDD2.n2 42.642
R79 VDD2.n5 VDD2.t7 2.90273
R80 VDD2.n5 VDD2.t6 2.90273
R81 VDD2.n3 VDD2.t1 2.90273
R82 VDD2.n3 VDD2.t0 2.90273
R83 VDD2.n1 VDD2.t3 2.90273
R84 VDD2.n1 VDD2.t2 2.90273
R85 VDD2.n0 VDD2.t5 2.90273
R86 VDD2.n0 VDD2.t4 2.90273
R87 VDD2 VDD2.n4 1.08886
R88 VTAIL.n11 VTAIL.t6 64.6315
R89 VTAIL.n10 VTAIL.t12 64.6315
R90 VTAIL.n7 VTAIL.t14 64.6315
R91 VTAIL.n15 VTAIL.t9 64.6313
R92 VTAIL.n2 VTAIL.t8 64.6313
R93 VTAIL.n3 VTAIL.t7 64.6313
R94 VTAIL.n6 VTAIL.t3 64.6313
R95 VTAIL.n14 VTAIL.t4 64.6313
R96 VTAIL.n13 VTAIL.n12 61.7293
R97 VTAIL.n9 VTAIL.n8 61.7293
R98 VTAIL.n1 VTAIL.n0 61.729
R99 VTAIL.n5 VTAIL.n4 61.729
R100 VTAIL.n15 VTAIL.n14 24.0824
R101 VTAIL.n7 VTAIL.n6 24.0824
R102 VTAIL.n0 VTAIL.t11 2.90273
R103 VTAIL.n0 VTAIL.t13 2.90273
R104 VTAIL.n4 VTAIL.t5 2.90273
R105 VTAIL.n4 VTAIL.t1 2.90273
R106 VTAIL.n12 VTAIL.t0 2.90273
R107 VTAIL.n12 VTAIL.t2 2.90273
R108 VTAIL.n8 VTAIL.t10 2.90273
R109 VTAIL.n8 VTAIL.t15 2.90273
R110 VTAIL.n9 VTAIL.n7 2.06084
R111 VTAIL.n10 VTAIL.n9 2.06084
R112 VTAIL.n13 VTAIL.n11 2.06084
R113 VTAIL.n14 VTAIL.n13 2.06084
R114 VTAIL.n6 VTAIL.n5 2.06084
R115 VTAIL.n5 VTAIL.n3 2.06084
R116 VTAIL.n2 VTAIL.n1 2.06084
R117 VTAIL VTAIL.n15 2.00266
R118 VTAIL.n11 VTAIL.n10 0.470328
R119 VTAIL.n3 VTAIL.n2 0.470328
R120 VTAIL VTAIL.n1 0.0586897
R121 B.n513 B.n512 585
R122 B.n514 B.n71 585
R123 B.n516 B.n515 585
R124 B.n517 B.n70 585
R125 B.n519 B.n518 585
R126 B.n520 B.n69 585
R127 B.n522 B.n521 585
R128 B.n523 B.n68 585
R129 B.n525 B.n524 585
R130 B.n526 B.n67 585
R131 B.n528 B.n527 585
R132 B.n529 B.n66 585
R133 B.n531 B.n530 585
R134 B.n532 B.n65 585
R135 B.n534 B.n533 585
R136 B.n535 B.n64 585
R137 B.n537 B.n536 585
R138 B.n538 B.n63 585
R139 B.n540 B.n539 585
R140 B.n541 B.n62 585
R141 B.n543 B.n542 585
R142 B.n544 B.n61 585
R143 B.n546 B.n545 585
R144 B.n547 B.n60 585
R145 B.n549 B.n548 585
R146 B.n550 B.n59 585
R147 B.n552 B.n551 585
R148 B.n553 B.n58 585
R149 B.n555 B.n554 585
R150 B.n556 B.n57 585
R151 B.n558 B.n557 585
R152 B.n559 B.n56 585
R153 B.n561 B.n560 585
R154 B.n562 B.n55 585
R155 B.n564 B.n563 585
R156 B.n565 B.n54 585
R157 B.n567 B.n566 585
R158 B.n568 B.n53 585
R159 B.n570 B.n569 585
R160 B.n572 B.n571 585
R161 B.n573 B.n49 585
R162 B.n575 B.n574 585
R163 B.n576 B.n48 585
R164 B.n578 B.n577 585
R165 B.n579 B.n47 585
R166 B.n581 B.n580 585
R167 B.n582 B.n46 585
R168 B.n584 B.n583 585
R169 B.n585 B.n43 585
R170 B.n588 B.n587 585
R171 B.n589 B.n42 585
R172 B.n591 B.n590 585
R173 B.n592 B.n41 585
R174 B.n594 B.n593 585
R175 B.n595 B.n40 585
R176 B.n597 B.n596 585
R177 B.n598 B.n39 585
R178 B.n600 B.n599 585
R179 B.n601 B.n38 585
R180 B.n603 B.n602 585
R181 B.n604 B.n37 585
R182 B.n606 B.n605 585
R183 B.n607 B.n36 585
R184 B.n609 B.n608 585
R185 B.n610 B.n35 585
R186 B.n612 B.n611 585
R187 B.n613 B.n34 585
R188 B.n615 B.n614 585
R189 B.n616 B.n33 585
R190 B.n618 B.n617 585
R191 B.n619 B.n32 585
R192 B.n621 B.n620 585
R193 B.n622 B.n31 585
R194 B.n624 B.n623 585
R195 B.n625 B.n30 585
R196 B.n627 B.n626 585
R197 B.n628 B.n29 585
R198 B.n630 B.n629 585
R199 B.n631 B.n28 585
R200 B.n633 B.n632 585
R201 B.n634 B.n27 585
R202 B.n636 B.n635 585
R203 B.n637 B.n26 585
R204 B.n639 B.n638 585
R205 B.n640 B.n25 585
R206 B.n642 B.n641 585
R207 B.n643 B.n24 585
R208 B.n645 B.n644 585
R209 B.n511 B.n72 585
R210 B.n510 B.n509 585
R211 B.n508 B.n73 585
R212 B.n507 B.n506 585
R213 B.n505 B.n74 585
R214 B.n504 B.n503 585
R215 B.n502 B.n75 585
R216 B.n501 B.n500 585
R217 B.n499 B.n76 585
R218 B.n498 B.n497 585
R219 B.n496 B.n77 585
R220 B.n495 B.n494 585
R221 B.n493 B.n78 585
R222 B.n492 B.n491 585
R223 B.n490 B.n79 585
R224 B.n489 B.n488 585
R225 B.n487 B.n80 585
R226 B.n486 B.n485 585
R227 B.n484 B.n81 585
R228 B.n483 B.n482 585
R229 B.n481 B.n82 585
R230 B.n480 B.n479 585
R231 B.n478 B.n83 585
R232 B.n477 B.n476 585
R233 B.n475 B.n84 585
R234 B.n474 B.n473 585
R235 B.n472 B.n85 585
R236 B.n471 B.n470 585
R237 B.n469 B.n86 585
R238 B.n468 B.n467 585
R239 B.n466 B.n87 585
R240 B.n465 B.n464 585
R241 B.n463 B.n88 585
R242 B.n462 B.n461 585
R243 B.n460 B.n89 585
R244 B.n459 B.n458 585
R245 B.n457 B.n90 585
R246 B.n456 B.n455 585
R247 B.n454 B.n91 585
R248 B.n453 B.n452 585
R249 B.n451 B.n92 585
R250 B.n450 B.n449 585
R251 B.n448 B.n93 585
R252 B.n447 B.n446 585
R253 B.n445 B.n94 585
R254 B.n444 B.n443 585
R255 B.n442 B.n95 585
R256 B.n441 B.n440 585
R257 B.n439 B.n96 585
R258 B.n438 B.n437 585
R259 B.n436 B.n97 585
R260 B.n435 B.n434 585
R261 B.n433 B.n98 585
R262 B.n432 B.n431 585
R263 B.n430 B.n99 585
R264 B.n429 B.n428 585
R265 B.n427 B.n100 585
R266 B.n426 B.n425 585
R267 B.n424 B.n101 585
R268 B.n423 B.n422 585
R269 B.n421 B.n102 585
R270 B.n420 B.n419 585
R271 B.n418 B.n103 585
R272 B.n417 B.n416 585
R273 B.n415 B.n104 585
R274 B.n414 B.n413 585
R275 B.n412 B.n105 585
R276 B.n411 B.n410 585
R277 B.n409 B.n106 585
R278 B.n408 B.n407 585
R279 B.n406 B.n107 585
R280 B.n405 B.n404 585
R281 B.n403 B.n108 585
R282 B.n402 B.n401 585
R283 B.n400 B.n109 585
R284 B.n399 B.n398 585
R285 B.n397 B.n110 585
R286 B.n396 B.n395 585
R287 B.n394 B.n111 585
R288 B.n393 B.n392 585
R289 B.n391 B.n112 585
R290 B.n390 B.n389 585
R291 B.n388 B.n113 585
R292 B.n387 B.n386 585
R293 B.n385 B.n114 585
R294 B.n384 B.n383 585
R295 B.n382 B.n115 585
R296 B.n249 B.n248 585
R297 B.n250 B.n163 585
R298 B.n252 B.n251 585
R299 B.n253 B.n162 585
R300 B.n255 B.n254 585
R301 B.n256 B.n161 585
R302 B.n258 B.n257 585
R303 B.n259 B.n160 585
R304 B.n261 B.n260 585
R305 B.n262 B.n159 585
R306 B.n264 B.n263 585
R307 B.n265 B.n158 585
R308 B.n267 B.n266 585
R309 B.n268 B.n157 585
R310 B.n270 B.n269 585
R311 B.n271 B.n156 585
R312 B.n273 B.n272 585
R313 B.n274 B.n155 585
R314 B.n276 B.n275 585
R315 B.n277 B.n154 585
R316 B.n279 B.n278 585
R317 B.n280 B.n153 585
R318 B.n282 B.n281 585
R319 B.n283 B.n152 585
R320 B.n285 B.n284 585
R321 B.n286 B.n151 585
R322 B.n288 B.n287 585
R323 B.n289 B.n150 585
R324 B.n291 B.n290 585
R325 B.n292 B.n149 585
R326 B.n294 B.n293 585
R327 B.n295 B.n148 585
R328 B.n297 B.n296 585
R329 B.n298 B.n147 585
R330 B.n300 B.n299 585
R331 B.n301 B.n146 585
R332 B.n303 B.n302 585
R333 B.n304 B.n145 585
R334 B.n306 B.n305 585
R335 B.n308 B.n307 585
R336 B.n309 B.n141 585
R337 B.n311 B.n310 585
R338 B.n312 B.n140 585
R339 B.n314 B.n313 585
R340 B.n315 B.n139 585
R341 B.n317 B.n316 585
R342 B.n318 B.n138 585
R343 B.n320 B.n319 585
R344 B.n321 B.n135 585
R345 B.n324 B.n323 585
R346 B.n325 B.n134 585
R347 B.n327 B.n326 585
R348 B.n328 B.n133 585
R349 B.n330 B.n329 585
R350 B.n331 B.n132 585
R351 B.n333 B.n332 585
R352 B.n334 B.n131 585
R353 B.n336 B.n335 585
R354 B.n337 B.n130 585
R355 B.n339 B.n338 585
R356 B.n340 B.n129 585
R357 B.n342 B.n341 585
R358 B.n343 B.n128 585
R359 B.n345 B.n344 585
R360 B.n346 B.n127 585
R361 B.n348 B.n347 585
R362 B.n349 B.n126 585
R363 B.n351 B.n350 585
R364 B.n352 B.n125 585
R365 B.n354 B.n353 585
R366 B.n355 B.n124 585
R367 B.n357 B.n356 585
R368 B.n358 B.n123 585
R369 B.n360 B.n359 585
R370 B.n361 B.n122 585
R371 B.n363 B.n362 585
R372 B.n364 B.n121 585
R373 B.n366 B.n365 585
R374 B.n367 B.n120 585
R375 B.n369 B.n368 585
R376 B.n370 B.n119 585
R377 B.n372 B.n371 585
R378 B.n373 B.n118 585
R379 B.n375 B.n374 585
R380 B.n376 B.n117 585
R381 B.n378 B.n377 585
R382 B.n379 B.n116 585
R383 B.n381 B.n380 585
R384 B.n247 B.n164 585
R385 B.n246 B.n245 585
R386 B.n244 B.n165 585
R387 B.n243 B.n242 585
R388 B.n241 B.n166 585
R389 B.n240 B.n239 585
R390 B.n238 B.n167 585
R391 B.n237 B.n236 585
R392 B.n235 B.n168 585
R393 B.n234 B.n233 585
R394 B.n232 B.n169 585
R395 B.n231 B.n230 585
R396 B.n229 B.n170 585
R397 B.n228 B.n227 585
R398 B.n226 B.n171 585
R399 B.n225 B.n224 585
R400 B.n223 B.n172 585
R401 B.n222 B.n221 585
R402 B.n220 B.n173 585
R403 B.n219 B.n218 585
R404 B.n217 B.n174 585
R405 B.n216 B.n215 585
R406 B.n214 B.n175 585
R407 B.n213 B.n212 585
R408 B.n211 B.n176 585
R409 B.n210 B.n209 585
R410 B.n208 B.n177 585
R411 B.n207 B.n206 585
R412 B.n205 B.n178 585
R413 B.n204 B.n203 585
R414 B.n202 B.n179 585
R415 B.n201 B.n200 585
R416 B.n199 B.n180 585
R417 B.n198 B.n197 585
R418 B.n196 B.n181 585
R419 B.n195 B.n194 585
R420 B.n193 B.n182 585
R421 B.n192 B.n191 585
R422 B.n190 B.n183 585
R423 B.n189 B.n188 585
R424 B.n187 B.n184 585
R425 B.n186 B.n185 585
R426 B.n2 B.n0 585
R427 B.n709 B.n1 585
R428 B.n708 B.n707 585
R429 B.n706 B.n3 585
R430 B.n705 B.n704 585
R431 B.n703 B.n4 585
R432 B.n702 B.n701 585
R433 B.n700 B.n5 585
R434 B.n699 B.n698 585
R435 B.n697 B.n6 585
R436 B.n696 B.n695 585
R437 B.n694 B.n7 585
R438 B.n693 B.n692 585
R439 B.n691 B.n8 585
R440 B.n690 B.n689 585
R441 B.n688 B.n9 585
R442 B.n687 B.n686 585
R443 B.n685 B.n10 585
R444 B.n684 B.n683 585
R445 B.n682 B.n11 585
R446 B.n681 B.n680 585
R447 B.n679 B.n12 585
R448 B.n678 B.n677 585
R449 B.n676 B.n13 585
R450 B.n675 B.n674 585
R451 B.n673 B.n14 585
R452 B.n672 B.n671 585
R453 B.n670 B.n15 585
R454 B.n669 B.n668 585
R455 B.n667 B.n16 585
R456 B.n666 B.n665 585
R457 B.n664 B.n17 585
R458 B.n663 B.n662 585
R459 B.n661 B.n18 585
R460 B.n660 B.n659 585
R461 B.n658 B.n19 585
R462 B.n657 B.n656 585
R463 B.n655 B.n20 585
R464 B.n654 B.n653 585
R465 B.n652 B.n21 585
R466 B.n651 B.n650 585
R467 B.n649 B.n22 585
R468 B.n648 B.n647 585
R469 B.n646 B.n23 585
R470 B.n711 B.n710 585
R471 B.n248 B.n247 550.159
R472 B.n644 B.n23 550.159
R473 B.n380 B.n115 550.159
R474 B.n512 B.n511 550.159
R475 B.n136 B.t0 338.084
R476 B.n142 B.t6 338.084
R477 B.n44 B.t3 338.084
R478 B.n50 B.t9 338.084
R479 B.n247 B.n246 163.367
R480 B.n246 B.n165 163.367
R481 B.n242 B.n165 163.367
R482 B.n242 B.n241 163.367
R483 B.n241 B.n240 163.367
R484 B.n240 B.n167 163.367
R485 B.n236 B.n167 163.367
R486 B.n236 B.n235 163.367
R487 B.n235 B.n234 163.367
R488 B.n234 B.n169 163.367
R489 B.n230 B.n169 163.367
R490 B.n230 B.n229 163.367
R491 B.n229 B.n228 163.367
R492 B.n228 B.n171 163.367
R493 B.n224 B.n171 163.367
R494 B.n224 B.n223 163.367
R495 B.n223 B.n222 163.367
R496 B.n222 B.n173 163.367
R497 B.n218 B.n173 163.367
R498 B.n218 B.n217 163.367
R499 B.n217 B.n216 163.367
R500 B.n216 B.n175 163.367
R501 B.n212 B.n175 163.367
R502 B.n212 B.n211 163.367
R503 B.n211 B.n210 163.367
R504 B.n210 B.n177 163.367
R505 B.n206 B.n177 163.367
R506 B.n206 B.n205 163.367
R507 B.n205 B.n204 163.367
R508 B.n204 B.n179 163.367
R509 B.n200 B.n179 163.367
R510 B.n200 B.n199 163.367
R511 B.n199 B.n198 163.367
R512 B.n198 B.n181 163.367
R513 B.n194 B.n181 163.367
R514 B.n194 B.n193 163.367
R515 B.n193 B.n192 163.367
R516 B.n192 B.n183 163.367
R517 B.n188 B.n183 163.367
R518 B.n188 B.n187 163.367
R519 B.n187 B.n186 163.367
R520 B.n186 B.n2 163.367
R521 B.n710 B.n2 163.367
R522 B.n710 B.n709 163.367
R523 B.n709 B.n708 163.367
R524 B.n708 B.n3 163.367
R525 B.n704 B.n3 163.367
R526 B.n704 B.n703 163.367
R527 B.n703 B.n702 163.367
R528 B.n702 B.n5 163.367
R529 B.n698 B.n5 163.367
R530 B.n698 B.n697 163.367
R531 B.n697 B.n696 163.367
R532 B.n696 B.n7 163.367
R533 B.n692 B.n7 163.367
R534 B.n692 B.n691 163.367
R535 B.n691 B.n690 163.367
R536 B.n690 B.n9 163.367
R537 B.n686 B.n9 163.367
R538 B.n686 B.n685 163.367
R539 B.n685 B.n684 163.367
R540 B.n684 B.n11 163.367
R541 B.n680 B.n11 163.367
R542 B.n680 B.n679 163.367
R543 B.n679 B.n678 163.367
R544 B.n678 B.n13 163.367
R545 B.n674 B.n13 163.367
R546 B.n674 B.n673 163.367
R547 B.n673 B.n672 163.367
R548 B.n672 B.n15 163.367
R549 B.n668 B.n15 163.367
R550 B.n668 B.n667 163.367
R551 B.n667 B.n666 163.367
R552 B.n666 B.n17 163.367
R553 B.n662 B.n17 163.367
R554 B.n662 B.n661 163.367
R555 B.n661 B.n660 163.367
R556 B.n660 B.n19 163.367
R557 B.n656 B.n19 163.367
R558 B.n656 B.n655 163.367
R559 B.n655 B.n654 163.367
R560 B.n654 B.n21 163.367
R561 B.n650 B.n21 163.367
R562 B.n650 B.n649 163.367
R563 B.n649 B.n648 163.367
R564 B.n648 B.n23 163.367
R565 B.n248 B.n163 163.367
R566 B.n252 B.n163 163.367
R567 B.n253 B.n252 163.367
R568 B.n254 B.n253 163.367
R569 B.n254 B.n161 163.367
R570 B.n258 B.n161 163.367
R571 B.n259 B.n258 163.367
R572 B.n260 B.n259 163.367
R573 B.n260 B.n159 163.367
R574 B.n264 B.n159 163.367
R575 B.n265 B.n264 163.367
R576 B.n266 B.n265 163.367
R577 B.n266 B.n157 163.367
R578 B.n270 B.n157 163.367
R579 B.n271 B.n270 163.367
R580 B.n272 B.n271 163.367
R581 B.n272 B.n155 163.367
R582 B.n276 B.n155 163.367
R583 B.n277 B.n276 163.367
R584 B.n278 B.n277 163.367
R585 B.n278 B.n153 163.367
R586 B.n282 B.n153 163.367
R587 B.n283 B.n282 163.367
R588 B.n284 B.n283 163.367
R589 B.n284 B.n151 163.367
R590 B.n288 B.n151 163.367
R591 B.n289 B.n288 163.367
R592 B.n290 B.n289 163.367
R593 B.n290 B.n149 163.367
R594 B.n294 B.n149 163.367
R595 B.n295 B.n294 163.367
R596 B.n296 B.n295 163.367
R597 B.n296 B.n147 163.367
R598 B.n300 B.n147 163.367
R599 B.n301 B.n300 163.367
R600 B.n302 B.n301 163.367
R601 B.n302 B.n145 163.367
R602 B.n306 B.n145 163.367
R603 B.n307 B.n306 163.367
R604 B.n307 B.n141 163.367
R605 B.n311 B.n141 163.367
R606 B.n312 B.n311 163.367
R607 B.n313 B.n312 163.367
R608 B.n313 B.n139 163.367
R609 B.n317 B.n139 163.367
R610 B.n318 B.n317 163.367
R611 B.n319 B.n318 163.367
R612 B.n319 B.n135 163.367
R613 B.n324 B.n135 163.367
R614 B.n325 B.n324 163.367
R615 B.n326 B.n325 163.367
R616 B.n326 B.n133 163.367
R617 B.n330 B.n133 163.367
R618 B.n331 B.n330 163.367
R619 B.n332 B.n331 163.367
R620 B.n332 B.n131 163.367
R621 B.n336 B.n131 163.367
R622 B.n337 B.n336 163.367
R623 B.n338 B.n337 163.367
R624 B.n338 B.n129 163.367
R625 B.n342 B.n129 163.367
R626 B.n343 B.n342 163.367
R627 B.n344 B.n343 163.367
R628 B.n344 B.n127 163.367
R629 B.n348 B.n127 163.367
R630 B.n349 B.n348 163.367
R631 B.n350 B.n349 163.367
R632 B.n350 B.n125 163.367
R633 B.n354 B.n125 163.367
R634 B.n355 B.n354 163.367
R635 B.n356 B.n355 163.367
R636 B.n356 B.n123 163.367
R637 B.n360 B.n123 163.367
R638 B.n361 B.n360 163.367
R639 B.n362 B.n361 163.367
R640 B.n362 B.n121 163.367
R641 B.n366 B.n121 163.367
R642 B.n367 B.n366 163.367
R643 B.n368 B.n367 163.367
R644 B.n368 B.n119 163.367
R645 B.n372 B.n119 163.367
R646 B.n373 B.n372 163.367
R647 B.n374 B.n373 163.367
R648 B.n374 B.n117 163.367
R649 B.n378 B.n117 163.367
R650 B.n379 B.n378 163.367
R651 B.n380 B.n379 163.367
R652 B.n384 B.n115 163.367
R653 B.n385 B.n384 163.367
R654 B.n386 B.n385 163.367
R655 B.n386 B.n113 163.367
R656 B.n390 B.n113 163.367
R657 B.n391 B.n390 163.367
R658 B.n392 B.n391 163.367
R659 B.n392 B.n111 163.367
R660 B.n396 B.n111 163.367
R661 B.n397 B.n396 163.367
R662 B.n398 B.n397 163.367
R663 B.n398 B.n109 163.367
R664 B.n402 B.n109 163.367
R665 B.n403 B.n402 163.367
R666 B.n404 B.n403 163.367
R667 B.n404 B.n107 163.367
R668 B.n408 B.n107 163.367
R669 B.n409 B.n408 163.367
R670 B.n410 B.n409 163.367
R671 B.n410 B.n105 163.367
R672 B.n414 B.n105 163.367
R673 B.n415 B.n414 163.367
R674 B.n416 B.n415 163.367
R675 B.n416 B.n103 163.367
R676 B.n420 B.n103 163.367
R677 B.n421 B.n420 163.367
R678 B.n422 B.n421 163.367
R679 B.n422 B.n101 163.367
R680 B.n426 B.n101 163.367
R681 B.n427 B.n426 163.367
R682 B.n428 B.n427 163.367
R683 B.n428 B.n99 163.367
R684 B.n432 B.n99 163.367
R685 B.n433 B.n432 163.367
R686 B.n434 B.n433 163.367
R687 B.n434 B.n97 163.367
R688 B.n438 B.n97 163.367
R689 B.n439 B.n438 163.367
R690 B.n440 B.n439 163.367
R691 B.n440 B.n95 163.367
R692 B.n444 B.n95 163.367
R693 B.n445 B.n444 163.367
R694 B.n446 B.n445 163.367
R695 B.n446 B.n93 163.367
R696 B.n450 B.n93 163.367
R697 B.n451 B.n450 163.367
R698 B.n452 B.n451 163.367
R699 B.n452 B.n91 163.367
R700 B.n456 B.n91 163.367
R701 B.n457 B.n456 163.367
R702 B.n458 B.n457 163.367
R703 B.n458 B.n89 163.367
R704 B.n462 B.n89 163.367
R705 B.n463 B.n462 163.367
R706 B.n464 B.n463 163.367
R707 B.n464 B.n87 163.367
R708 B.n468 B.n87 163.367
R709 B.n469 B.n468 163.367
R710 B.n470 B.n469 163.367
R711 B.n470 B.n85 163.367
R712 B.n474 B.n85 163.367
R713 B.n475 B.n474 163.367
R714 B.n476 B.n475 163.367
R715 B.n476 B.n83 163.367
R716 B.n480 B.n83 163.367
R717 B.n481 B.n480 163.367
R718 B.n482 B.n481 163.367
R719 B.n482 B.n81 163.367
R720 B.n486 B.n81 163.367
R721 B.n487 B.n486 163.367
R722 B.n488 B.n487 163.367
R723 B.n488 B.n79 163.367
R724 B.n492 B.n79 163.367
R725 B.n493 B.n492 163.367
R726 B.n494 B.n493 163.367
R727 B.n494 B.n77 163.367
R728 B.n498 B.n77 163.367
R729 B.n499 B.n498 163.367
R730 B.n500 B.n499 163.367
R731 B.n500 B.n75 163.367
R732 B.n504 B.n75 163.367
R733 B.n505 B.n504 163.367
R734 B.n506 B.n505 163.367
R735 B.n506 B.n73 163.367
R736 B.n510 B.n73 163.367
R737 B.n511 B.n510 163.367
R738 B.n644 B.n643 163.367
R739 B.n643 B.n642 163.367
R740 B.n642 B.n25 163.367
R741 B.n638 B.n25 163.367
R742 B.n638 B.n637 163.367
R743 B.n637 B.n636 163.367
R744 B.n636 B.n27 163.367
R745 B.n632 B.n27 163.367
R746 B.n632 B.n631 163.367
R747 B.n631 B.n630 163.367
R748 B.n630 B.n29 163.367
R749 B.n626 B.n29 163.367
R750 B.n626 B.n625 163.367
R751 B.n625 B.n624 163.367
R752 B.n624 B.n31 163.367
R753 B.n620 B.n31 163.367
R754 B.n620 B.n619 163.367
R755 B.n619 B.n618 163.367
R756 B.n618 B.n33 163.367
R757 B.n614 B.n33 163.367
R758 B.n614 B.n613 163.367
R759 B.n613 B.n612 163.367
R760 B.n612 B.n35 163.367
R761 B.n608 B.n35 163.367
R762 B.n608 B.n607 163.367
R763 B.n607 B.n606 163.367
R764 B.n606 B.n37 163.367
R765 B.n602 B.n37 163.367
R766 B.n602 B.n601 163.367
R767 B.n601 B.n600 163.367
R768 B.n600 B.n39 163.367
R769 B.n596 B.n39 163.367
R770 B.n596 B.n595 163.367
R771 B.n595 B.n594 163.367
R772 B.n594 B.n41 163.367
R773 B.n590 B.n41 163.367
R774 B.n590 B.n589 163.367
R775 B.n589 B.n588 163.367
R776 B.n588 B.n43 163.367
R777 B.n583 B.n43 163.367
R778 B.n583 B.n582 163.367
R779 B.n582 B.n581 163.367
R780 B.n581 B.n47 163.367
R781 B.n577 B.n47 163.367
R782 B.n577 B.n576 163.367
R783 B.n576 B.n575 163.367
R784 B.n575 B.n49 163.367
R785 B.n571 B.n49 163.367
R786 B.n571 B.n570 163.367
R787 B.n570 B.n53 163.367
R788 B.n566 B.n53 163.367
R789 B.n566 B.n565 163.367
R790 B.n565 B.n564 163.367
R791 B.n564 B.n55 163.367
R792 B.n560 B.n55 163.367
R793 B.n560 B.n559 163.367
R794 B.n559 B.n558 163.367
R795 B.n558 B.n57 163.367
R796 B.n554 B.n57 163.367
R797 B.n554 B.n553 163.367
R798 B.n553 B.n552 163.367
R799 B.n552 B.n59 163.367
R800 B.n548 B.n59 163.367
R801 B.n548 B.n547 163.367
R802 B.n547 B.n546 163.367
R803 B.n546 B.n61 163.367
R804 B.n542 B.n61 163.367
R805 B.n542 B.n541 163.367
R806 B.n541 B.n540 163.367
R807 B.n540 B.n63 163.367
R808 B.n536 B.n63 163.367
R809 B.n536 B.n535 163.367
R810 B.n535 B.n534 163.367
R811 B.n534 B.n65 163.367
R812 B.n530 B.n65 163.367
R813 B.n530 B.n529 163.367
R814 B.n529 B.n528 163.367
R815 B.n528 B.n67 163.367
R816 B.n524 B.n67 163.367
R817 B.n524 B.n523 163.367
R818 B.n523 B.n522 163.367
R819 B.n522 B.n69 163.367
R820 B.n518 B.n69 163.367
R821 B.n518 B.n517 163.367
R822 B.n517 B.n516 163.367
R823 B.n516 B.n71 163.367
R824 B.n512 B.n71 163.367
R825 B.n136 B.t2 159.863
R826 B.n50 B.t10 159.863
R827 B.n142 B.t8 159.851
R828 B.n44 B.t4 159.851
R829 B.n137 B.t1 113.513
R830 B.n51 B.t11 113.513
R831 B.n143 B.t7 113.499
R832 B.n45 B.t5 113.499
R833 B.n322 B.n137 59.5399
R834 B.n144 B.n143 59.5399
R835 B.n586 B.n45 59.5399
R836 B.n52 B.n51 59.5399
R837 B.n137 B.n136 46.352
R838 B.n143 B.n142 46.352
R839 B.n45 B.n44 46.352
R840 B.n51 B.n50 46.352
R841 B.n513 B.n72 35.7468
R842 B.n646 B.n645 35.7468
R843 B.n382 B.n381 35.7468
R844 B.n249 B.n164 35.7468
R845 B B.n711 18.0485
R846 B.n645 B.n24 10.6151
R847 B.n641 B.n24 10.6151
R848 B.n641 B.n640 10.6151
R849 B.n640 B.n639 10.6151
R850 B.n639 B.n26 10.6151
R851 B.n635 B.n26 10.6151
R852 B.n635 B.n634 10.6151
R853 B.n634 B.n633 10.6151
R854 B.n633 B.n28 10.6151
R855 B.n629 B.n28 10.6151
R856 B.n629 B.n628 10.6151
R857 B.n628 B.n627 10.6151
R858 B.n627 B.n30 10.6151
R859 B.n623 B.n30 10.6151
R860 B.n623 B.n622 10.6151
R861 B.n622 B.n621 10.6151
R862 B.n621 B.n32 10.6151
R863 B.n617 B.n32 10.6151
R864 B.n617 B.n616 10.6151
R865 B.n616 B.n615 10.6151
R866 B.n615 B.n34 10.6151
R867 B.n611 B.n34 10.6151
R868 B.n611 B.n610 10.6151
R869 B.n610 B.n609 10.6151
R870 B.n609 B.n36 10.6151
R871 B.n605 B.n36 10.6151
R872 B.n605 B.n604 10.6151
R873 B.n604 B.n603 10.6151
R874 B.n603 B.n38 10.6151
R875 B.n599 B.n38 10.6151
R876 B.n599 B.n598 10.6151
R877 B.n598 B.n597 10.6151
R878 B.n597 B.n40 10.6151
R879 B.n593 B.n40 10.6151
R880 B.n593 B.n592 10.6151
R881 B.n592 B.n591 10.6151
R882 B.n591 B.n42 10.6151
R883 B.n587 B.n42 10.6151
R884 B.n585 B.n584 10.6151
R885 B.n584 B.n46 10.6151
R886 B.n580 B.n46 10.6151
R887 B.n580 B.n579 10.6151
R888 B.n579 B.n578 10.6151
R889 B.n578 B.n48 10.6151
R890 B.n574 B.n48 10.6151
R891 B.n574 B.n573 10.6151
R892 B.n573 B.n572 10.6151
R893 B.n569 B.n568 10.6151
R894 B.n568 B.n567 10.6151
R895 B.n567 B.n54 10.6151
R896 B.n563 B.n54 10.6151
R897 B.n563 B.n562 10.6151
R898 B.n562 B.n561 10.6151
R899 B.n561 B.n56 10.6151
R900 B.n557 B.n56 10.6151
R901 B.n557 B.n556 10.6151
R902 B.n556 B.n555 10.6151
R903 B.n555 B.n58 10.6151
R904 B.n551 B.n58 10.6151
R905 B.n551 B.n550 10.6151
R906 B.n550 B.n549 10.6151
R907 B.n549 B.n60 10.6151
R908 B.n545 B.n60 10.6151
R909 B.n545 B.n544 10.6151
R910 B.n544 B.n543 10.6151
R911 B.n543 B.n62 10.6151
R912 B.n539 B.n62 10.6151
R913 B.n539 B.n538 10.6151
R914 B.n538 B.n537 10.6151
R915 B.n537 B.n64 10.6151
R916 B.n533 B.n64 10.6151
R917 B.n533 B.n532 10.6151
R918 B.n532 B.n531 10.6151
R919 B.n531 B.n66 10.6151
R920 B.n527 B.n66 10.6151
R921 B.n527 B.n526 10.6151
R922 B.n526 B.n525 10.6151
R923 B.n525 B.n68 10.6151
R924 B.n521 B.n68 10.6151
R925 B.n521 B.n520 10.6151
R926 B.n520 B.n519 10.6151
R927 B.n519 B.n70 10.6151
R928 B.n515 B.n70 10.6151
R929 B.n515 B.n514 10.6151
R930 B.n514 B.n513 10.6151
R931 B.n383 B.n382 10.6151
R932 B.n383 B.n114 10.6151
R933 B.n387 B.n114 10.6151
R934 B.n388 B.n387 10.6151
R935 B.n389 B.n388 10.6151
R936 B.n389 B.n112 10.6151
R937 B.n393 B.n112 10.6151
R938 B.n394 B.n393 10.6151
R939 B.n395 B.n394 10.6151
R940 B.n395 B.n110 10.6151
R941 B.n399 B.n110 10.6151
R942 B.n400 B.n399 10.6151
R943 B.n401 B.n400 10.6151
R944 B.n401 B.n108 10.6151
R945 B.n405 B.n108 10.6151
R946 B.n406 B.n405 10.6151
R947 B.n407 B.n406 10.6151
R948 B.n407 B.n106 10.6151
R949 B.n411 B.n106 10.6151
R950 B.n412 B.n411 10.6151
R951 B.n413 B.n412 10.6151
R952 B.n413 B.n104 10.6151
R953 B.n417 B.n104 10.6151
R954 B.n418 B.n417 10.6151
R955 B.n419 B.n418 10.6151
R956 B.n419 B.n102 10.6151
R957 B.n423 B.n102 10.6151
R958 B.n424 B.n423 10.6151
R959 B.n425 B.n424 10.6151
R960 B.n425 B.n100 10.6151
R961 B.n429 B.n100 10.6151
R962 B.n430 B.n429 10.6151
R963 B.n431 B.n430 10.6151
R964 B.n431 B.n98 10.6151
R965 B.n435 B.n98 10.6151
R966 B.n436 B.n435 10.6151
R967 B.n437 B.n436 10.6151
R968 B.n437 B.n96 10.6151
R969 B.n441 B.n96 10.6151
R970 B.n442 B.n441 10.6151
R971 B.n443 B.n442 10.6151
R972 B.n443 B.n94 10.6151
R973 B.n447 B.n94 10.6151
R974 B.n448 B.n447 10.6151
R975 B.n449 B.n448 10.6151
R976 B.n449 B.n92 10.6151
R977 B.n453 B.n92 10.6151
R978 B.n454 B.n453 10.6151
R979 B.n455 B.n454 10.6151
R980 B.n455 B.n90 10.6151
R981 B.n459 B.n90 10.6151
R982 B.n460 B.n459 10.6151
R983 B.n461 B.n460 10.6151
R984 B.n461 B.n88 10.6151
R985 B.n465 B.n88 10.6151
R986 B.n466 B.n465 10.6151
R987 B.n467 B.n466 10.6151
R988 B.n467 B.n86 10.6151
R989 B.n471 B.n86 10.6151
R990 B.n472 B.n471 10.6151
R991 B.n473 B.n472 10.6151
R992 B.n473 B.n84 10.6151
R993 B.n477 B.n84 10.6151
R994 B.n478 B.n477 10.6151
R995 B.n479 B.n478 10.6151
R996 B.n479 B.n82 10.6151
R997 B.n483 B.n82 10.6151
R998 B.n484 B.n483 10.6151
R999 B.n485 B.n484 10.6151
R1000 B.n485 B.n80 10.6151
R1001 B.n489 B.n80 10.6151
R1002 B.n490 B.n489 10.6151
R1003 B.n491 B.n490 10.6151
R1004 B.n491 B.n78 10.6151
R1005 B.n495 B.n78 10.6151
R1006 B.n496 B.n495 10.6151
R1007 B.n497 B.n496 10.6151
R1008 B.n497 B.n76 10.6151
R1009 B.n501 B.n76 10.6151
R1010 B.n502 B.n501 10.6151
R1011 B.n503 B.n502 10.6151
R1012 B.n503 B.n74 10.6151
R1013 B.n507 B.n74 10.6151
R1014 B.n508 B.n507 10.6151
R1015 B.n509 B.n508 10.6151
R1016 B.n509 B.n72 10.6151
R1017 B.n250 B.n249 10.6151
R1018 B.n251 B.n250 10.6151
R1019 B.n251 B.n162 10.6151
R1020 B.n255 B.n162 10.6151
R1021 B.n256 B.n255 10.6151
R1022 B.n257 B.n256 10.6151
R1023 B.n257 B.n160 10.6151
R1024 B.n261 B.n160 10.6151
R1025 B.n262 B.n261 10.6151
R1026 B.n263 B.n262 10.6151
R1027 B.n263 B.n158 10.6151
R1028 B.n267 B.n158 10.6151
R1029 B.n268 B.n267 10.6151
R1030 B.n269 B.n268 10.6151
R1031 B.n269 B.n156 10.6151
R1032 B.n273 B.n156 10.6151
R1033 B.n274 B.n273 10.6151
R1034 B.n275 B.n274 10.6151
R1035 B.n275 B.n154 10.6151
R1036 B.n279 B.n154 10.6151
R1037 B.n280 B.n279 10.6151
R1038 B.n281 B.n280 10.6151
R1039 B.n281 B.n152 10.6151
R1040 B.n285 B.n152 10.6151
R1041 B.n286 B.n285 10.6151
R1042 B.n287 B.n286 10.6151
R1043 B.n287 B.n150 10.6151
R1044 B.n291 B.n150 10.6151
R1045 B.n292 B.n291 10.6151
R1046 B.n293 B.n292 10.6151
R1047 B.n293 B.n148 10.6151
R1048 B.n297 B.n148 10.6151
R1049 B.n298 B.n297 10.6151
R1050 B.n299 B.n298 10.6151
R1051 B.n299 B.n146 10.6151
R1052 B.n303 B.n146 10.6151
R1053 B.n304 B.n303 10.6151
R1054 B.n305 B.n304 10.6151
R1055 B.n309 B.n308 10.6151
R1056 B.n310 B.n309 10.6151
R1057 B.n310 B.n140 10.6151
R1058 B.n314 B.n140 10.6151
R1059 B.n315 B.n314 10.6151
R1060 B.n316 B.n315 10.6151
R1061 B.n316 B.n138 10.6151
R1062 B.n320 B.n138 10.6151
R1063 B.n321 B.n320 10.6151
R1064 B.n323 B.n134 10.6151
R1065 B.n327 B.n134 10.6151
R1066 B.n328 B.n327 10.6151
R1067 B.n329 B.n328 10.6151
R1068 B.n329 B.n132 10.6151
R1069 B.n333 B.n132 10.6151
R1070 B.n334 B.n333 10.6151
R1071 B.n335 B.n334 10.6151
R1072 B.n335 B.n130 10.6151
R1073 B.n339 B.n130 10.6151
R1074 B.n340 B.n339 10.6151
R1075 B.n341 B.n340 10.6151
R1076 B.n341 B.n128 10.6151
R1077 B.n345 B.n128 10.6151
R1078 B.n346 B.n345 10.6151
R1079 B.n347 B.n346 10.6151
R1080 B.n347 B.n126 10.6151
R1081 B.n351 B.n126 10.6151
R1082 B.n352 B.n351 10.6151
R1083 B.n353 B.n352 10.6151
R1084 B.n353 B.n124 10.6151
R1085 B.n357 B.n124 10.6151
R1086 B.n358 B.n357 10.6151
R1087 B.n359 B.n358 10.6151
R1088 B.n359 B.n122 10.6151
R1089 B.n363 B.n122 10.6151
R1090 B.n364 B.n363 10.6151
R1091 B.n365 B.n364 10.6151
R1092 B.n365 B.n120 10.6151
R1093 B.n369 B.n120 10.6151
R1094 B.n370 B.n369 10.6151
R1095 B.n371 B.n370 10.6151
R1096 B.n371 B.n118 10.6151
R1097 B.n375 B.n118 10.6151
R1098 B.n376 B.n375 10.6151
R1099 B.n377 B.n376 10.6151
R1100 B.n377 B.n116 10.6151
R1101 B.n381 B.n116 10.6151
R1102 B.n245 B.n164 10.6151
R1103 B.n245 B.n244 10.6151
R1104 B.n244 B.n243 10.6151
R1105 B.n243 B.n166 10.6151
R1106 B.n239 B.n166 10.6151
R1107 B.n239 B.n238 10.6151
R1108 B.n238 B.n237 10.6151
R1109 B.n237 B.n168 10.6151
R1110 B.n233 B.n168 10.6151
R1111 B.n233 B.n232 10.6151
R1112 B.n232 B.n231 10.6151
R1113 B.n231 B.n170 10.6151
R1114 B.n227 B.n170 10.6151
R1115 B.n227 B.n226 10.6151
R1116 B.n226 B.n225 10.6151
R1117 B.n225 B.n172 10.6151
R1118 B.n221 B.n172 10.6151
R1119 B.n221 B.n220 10.6151
R1120 B.n220 B.n219 10.6151
R1121 B.n219 B.n174 10.6151
R1122 B.n215 B.n174 10.6151
R1123 B.n215 B.n214 10.6151
R1124 B.n214 B.n213 10.6151
R1125 B.n213 B.n176 10.6151
R1126 B.n209 B.n176 10.6151
R1127 B.n209 B.n208 10.6151
R1128 B.n208 B.n207 10.6151
R1129 B.n207 B.n178 10.6151
R1130 B.n203 B.n178 10.6151
R1131 B.n203 B.n202 10.6151
R1132 B.n202 B.n201 10.6151
R1133 B.n201 B.n180 10.6151
R1134 B.n197 B.n180 10.6151
R1135 B.n197 B.n196 10.6151
R1136 B.n196 B.n195 10.6151
R1137 B.n195 B.n182 10.6151
R1138 B.n191 B.n182 10.6151
R1139 B.n191 B.n190 10.6151
R1140 B.n190 B.n189 10.6151
R1141 B.n189 B.n184 10.6151
R1142 B.n185 B.n184 10.6151
R1143 B.n185 B.n0 10.6151
R1144 B.n707 B.n1 10.6151
R1145 B.n707 B.n706 10.6151
R1146 B.n706 B.n705 10.6151
R1147 B.n705 B.n4 10.6151
R1148 B.n701 B.n4 10.6151
R1149 B.n701 B.n700 10.6151
R1150 B.n700 B.n699 10.6151
R1151 B.n699 B.n6 10.6151
R1152 B.n695 B.n6 10.6151
R1153 B.n695 B.n694 10.6151
R1154 B.n694 B.n693 10.6151
R1155 B.n693 B.n8 10.6151
R1156 B.n689 B.n8 10.6151
R1157 B.n689 B.n688 10.6151
R1158 B.n688 B.n687 10.6151
R1159 B.n687 B.n10 10.6151
R1160 B.n683 B.n10 10.6151
R1161 B.n683 B.n682 10.6151
R1162 B.n682 B.n681 10.6151
R1163 B.n681 B.n12 10.6151
R1164 B.n677 B.n12 10.6151
R1165 B.n677 B.n676 10.6151
R1166 B.n676 B.n675 10.6151
R1167 B.n675 B.n14 10.6151
R1168 B.n671 B.n14 10.6151
R1169 B.n671 B.n670 10.6151
R1170 B.n670 B.n669 10.6151
R1171 B.n669 B.n16 10.6151
R1172 B.n665 B.n16 10.6151
R1173 B.n665 B.n664 10.6151
R1174 B.n664 B.n663 10.6151
R1175 B.n663 B.n18 10.6151
R1176 B.n659 B.n18 10.6151
R1177 B.n659 B.n658 10.6151
R1178 B.n658 B.n657 10.6151
R1179 B.n657 B.n20 10.6151
R1180 B.n653 B.n20 10.6151
R1181 B.n653 B.n652 10.6151
R1182 B.n652 B.n651 10.6151
R1183 B.n651 B.n22 10.6151
R1184 B.n647 B.n22 10.6151
R1185 B.n647 B.n646 10.6151
R1186 B.n587 B.n586 9.36635
R1187 B.n569 B.n52 9.36635
R1188 B.n305 B.n144 9.36635
R1189 B.n323 B.n322 9.36635
R1190 B.n711 B.n0 2.81026
R1191 B.n711 B.n1 2.81026
R1192 B.n586 B.n585 1.24928
R1193 B.n572 B.n52 1.24928
R1194 B.n308 B.n144 1.24928
R1195 B.n322 B.n321 1.24928
R1196 VP.n13 VP.t0 164.535
R1197 VP.n15 VP.n12 161.3
R1198 VP.n17 VP.n16 161.3
R1199 VP.n18 VP.n11 161.3
R1200 VP.n20 VP.n19 161.3
R1201 VP.n22 VP.n10 161.3
R1202 VP.n24 VP.n23 161.3
R1203 VP.n25 VP.n9 161.3
R1204 VP.n27 VP.n26 161.3
R1205 VP.n28 VP.n8 161.3
R1206 VP.n54 VP.n0 161.3
R1207 VP.n53 VP.n52 161.3
R1208 VP.n51 VP.n1 161.3
R1209 VP.n50 VP.n49 161.3
R1210 VP.n48 VP.n2 161.3
R1211 VP.n46 VP.n45 161.3
R1212 VP.n44 VP.n3 161.3
R1213 VP.n43 VP.n42 161.3
R1214 VP.n41 VP.n4 161.3
R1215 VP.n39 VP.n38 161.3
R1216 VP.n37 VP.n5 161.3
R1217 VP.n36 VP.n35 161.3
R1218 VP.n34 VP.n6 161.3
R1219 VP.n33 VP.n32 161.3
R1220 VP.n7 VP.t1 131.03
R1221 VP.n40 VP.t4 131.03
R1222 VP.n47 VP.t2 131.03
R1223 VP.n55 VP.t6 131.03
R1224 VP.n29 VP.t7 131.03
R1225 VP.n21 VP.t3 131.03
R1226 VP.n14 VP.t5 131.03
R1227 VP.n31 VP.n7 94.4317
R1228 VP.n56 VP.n55 94.4317
R1229 VP.n30 VP.n29 94.4317
R1230 VP.n42 VP.n3 56.5617
R1231 VP.n16 VP.n11 56.5617
R1232 VP.n35 VP.n34 54.1398
R1233 VP.n53 VP.n1 54.1398
R1234 VP.n27 VP.n9 54.1398
R1235 VP.n14 VP.n13 48.8225
R1236 VP.n31 VP.n30 47.7497
R1237 VP.n35 VP.n5 27.0143
R1238 VP.n49 VP.n1 27.0143
R1239 VP.n23 VP.n9 27.0143
R1240 VP.n34 VP.n33 24.5923
R1241 VP.n39 VP.n5 24.5923
R1242 VP.n42 VP.n41 24.5923
R1243 VP.n46 VP.n3 24.5923
R1244 VP.n49 VP.n48 24.5923
R1245 VP.n54 VP.n53 24.5923
R1246 VP.n28 VP.n27 24.5923
R1247 VP.n20 VP.n11 24.5923
R1248 VP.n23 VP.n22 24.5923
R1249 VP.n16 VP.n15 24.5923
R1250 VP.n41 VP.n40 21.8872
R1251 VP.n47 VP.n46 21.8872
R1252 VP.n21 VP.n20 21.8872
R1253 VP.n15 VP.n14 21.8872
R1254 VP.n33 VP.n7 16.477
R1255 VP.n55 VP.n54 16.477
R1256 VP.n29 VP.n28 16.477
R1257 VP.n13 VP.n12 9.28418
R1258 VP.n40 VP.n39 2.7056
R1259 VP.n48 VP.n47 2.7056
R1260 VP.n22 VP.n21 2.7056
R1261 VP.n30 VP.n8 0.278335
R1262 VP.n32 VP.n31 0.278335
R1263 VP.n56 VP.n0 0.278335
R1264 VP.n17 VP.n12 0.189894
R1265 VP.n18 VP.n17 0.189894
R1266 VP.n19 VP.n18 0.189894
R1267 VP.n19 VP.n10 0.189894
R1268 VP.n24 VP.n10 0.189894
R1269 VP.n25 VP.n24 0.189894
R1270 VP.n26 VP.n25 0.189894
R1271 VP.n26 VP.n8 0.189894
R1272 VP.n32 VP.n6 0.189894
R1273 VP.n36 VP.n6 0.189894
R1274 VP.n37 VP.n36 0.189894
R1275 VP.n38 VP.n37 0.189894
R1276 VP.n38 VP.n4 0.189894
R1277 VP.n43 VP.n4 0.189894
R1278 VP.n44 VP.n43 0.189894
R1279 VP.n45 VP.n44 0.189894
R1280 VP.n45 VP.n2 0.189894
R1281 VP.n50 VP.n2 0.189894
R1282 VP.n51 VP.n50 0.189894
R1283 VP.n52 VP.n51 0.189894
R1284 VP.n52 VP.n0 0.189894
R1285 VP VP.n56 0.153485
R1286 VDD1 VDD1.n0 79.4964
R1287 VDD1.n3 VDD1.n2 79.3827
R1288 VDD1.n3 VDD1.n1 79.3827
R1289 VDD1.n5 VDD1.n4 78.4079
R1290 VDD1.n5 VDD1.n3 43.225
R1291 VDD1.n4 VDD1.t4 2.90273
R1292 VDD1.n4 VDD1.t0 2.90273
R1293 VDD1.n0 VDD1.t7 2.90273
R1294 VDD1.n0 VDD1.t2 2.90273
R1295 VDD1.n2 VDD1.t5 2.90273
R1296 VDD1.n2 VDD1.t1 2.90273
R1297 VDD1.n1 VDD1.t6 2.90273
R1298 VDD1.n1 VDD1.t3 2.90273
R1299 VDD1 VDD1.n5 0.972483
C0 B VDD1 1.46413f
C1 VTAIL VDD2 7.83029f
C2 B VDD2 1.54316f
C3 VDD1 w_n3360_n3208# 1.75757f
C4 w_n3360_n3208# VDD2 1.84963f
C5 VTAIL VP 8.0072f
C6 VN VTAIL 7.99309f
C7 B VP 1.81919f
C8 B VN 1.09352f
C9 VDD1 VDD2 1.49626f
C10 w_n3360_n3208# VP 7.10348f
C11 VN w_n3360_n3208# 6.66887f
C12 VDD1 VP 8.04827f
C13 VN VDD1 0.151066f
C14 B VTAIL 4.4669f
C15 VP VDD2 0.462523f
C16 VN VDD2 7.73794f
C17 VTAIL w_n3360_n3208# 3.99633f
C18 B w_n3360_n3208# 9.06442f
C19 VN VP 6.85193f
C20 VDD1 VTAIL 7.7795f
C21 VDD2 VSUBS 1.6125f
C22 VDD1 VSUBS 2.167579f
C23 VTAIL VSUBS 1.205143f
C24 VN VSUBS 6.028f
C25 VP VSUBS 3.006864f
C26 B VSUBS 4.330074f
C27 w_n3360_n3208# VSUBS 0.132854p
C28 VDD1.t7 VSUBS 0.218889f
C29 VDD1.t2 VSUBS 0.218889f
C30 VDD1.n0 VSUBS 1.70675f
C31 VDD1.t6 VSUBS 0.218889f
C32 VDD1.t3 VSUBS 0.218889f
C33 VDD1.n1 VSUBS 1.70564f
C34 VDD1.t5 VSUBS 0.218889f
C35 VDD1.t1 VSUBS 0.218889f
C36 VDD1.n2 VSUBS 1.70564f
C37 VDD1.n3 VSUBS 3.42244f
C38 VDD1.t4 VSUBS 0.218889f
C39 VDD1.t0 VSUBS 0.218889f
C40 VDD1.n4 VSUBS 1.69703f
C41 VDD1.n5 VSUBS 2.94737f
C42 VP.n0 VSUBS 0.045268f
C43 VP.t6 VSUBS 2.15414f
C44 VP.n1 VSUBS 0.037392f
C45 VP.n2 VSUBS 0.034338f
C46 VP.t2 VSUBS 2.15414f
C47 VP.n3 VSUBS 0.049915f
C48 VP.n4 VSUBS 0.034338f
C49 VP.t4 VSUBS 2.15414f
C50 VP.n5 VSUBS 0.066212f
C51 VP.n6 VSUBS 0.034338f
C52 VP.t1 VSUBS 2.15414f
C53 VP.n7 VSUBS 0.872433f
C54 VP.n8 VSUBS 0.045268f
C55 VP.t7 VSUBS 2.15414f
C56 VP.n9 VSUBS 0.037392f
C57 VP.n10 VSUBS 0.034338f
C58 VP.t3 VSUBS 2.15414f
C59 VP.n11 VSUBS 0.049915f
C60 VP.n12 VSUBS 0.287773f
C61 VP.t5 VSUBS 2.15414f
C62 VP.t0 VSUBS 2.34739f
C63 VP.n13 VSUBS 0.846373f
C64 VP.n14 VSUBS 0.868451f
C65 VP.n15 VSUBS 0.060218f
C66 VP.n16 VSUBS 0.049915f
C67 VP.n17 VSUBS 0.034338f
C68 VP.n18 VSUBS 0.034338f
C69 VP.n19 VSUBS 0.034338f
C70 VP.n20 VSUBS 0.060218f
C71 VP.n21 VSUBS 0.771508f
C72 VP.n22 VSUBS 0.035699f
C73 VP.n23 VSUBS 0.066212f
C74 VP.n24 VSUBS 0.034338f
C75 VP.n25 VSUBS 0.034338f
C76 VP.n26 VSUBS 0.034338f
C77 VP.n27 VSUBS 0.059902f
C78 VP.n28 VSUBS 0.053302f
C79 VP.n29 VSUBS 0.872433f
C80 VP.n30 VSUBS 1.77228f
C81 VP.n31 VSUBS 1.79821f
C82 VP.n32 VSUBS 0.045268f
C83 VP.n33 VSUBS 0.053302f
C84 VP.n34 VSUBS 0.059902f
C85 VP.n35 VSUBS 0.037392f
C86 VP.n36 VSUBS 0.034338f
C87 VP.n37 VSUBS 0.034338f
C88 VP.n38 VSUBS 0.034338f
C89 VP.n39 VSUBS 0.035699f
C90 VP.n40 VSUBS 0.771508f
C91 VP.n41 VSUBS 0.060218f
C92 VP.n42 VSUBS 0.049915f
C93 VP.n43 VSUBS 0.034338f
C94 VP.n44 VSUBS 0.034338f
C95 VP.n45 VSUBS 0.034338f
C96 VP.n46 VSUBS 0.060218f
C97 VP.n47 VSUBS 0.771508f
C98 VP.n48 VSUBS 0.035699f
C99 VP.n49 VSUBS 0.066212f
C100 VP.n50 VSUBS 0.034338f
C101 VP.n51 VSUBS 0.034338f
C102 VP.n52 VSUBS 0.034338f
C103 VP.n53 VSUBS 0.059902f
C104 VP.n54 VSUBS 0.053302f
C105 VP.n55 VSUBS 0.872433f
C106 VP.n56 VSUBS 0.045246f
C107 B.n0 VSUBS 0.004534f
C108 B.n1 VSUBS 0.004534f
C109 B.n2 VSUBS 0.007169f
C110 B.n3 VSUBS 0.007169f
C111 B.n4 VSUBS 0.007169f
C112 B.n5 VSUBS 0.007169f
C113 B.n6 VSUBS 0.007169f
C114 B.n7 VSUBS 0.007169f
C115 B.n8 VSUBS 0.007169f
C116 B.n9 VSUBS 0.007169f
C117 B.n10 VSUBS 0.007169f
C118 B.n11 VSUBS 0.007169f
C119 B.n12 VSUBS 0.007169f
C120 B.n13 VSUBS 0.007169f
C121 B.n14 VSUBS 0.007169f
C122 B.n15 VSUBS 0.007169f
C123 B.n16 VSUBS 0.007169f
C124 B.n17 VSUBS 0.007169f
C125 B.n18 VSUBS 0.007169f
C126 B.n19 VSUBS 0.007169f
C127 B.n20 VSUBS 0.007169f
C128 B.n21 VSUBS 0.007169f
C129 B.n22 VSUBS 0.007169f
C130 B.n23 VSUBS 0.017318f
C131 B.n24 VSUBS 0.007169f
C132 B.n25 VSUBS 0.007169f
C133 B.n26 VSUBS 0.007169f
C134 B.n27 VSUBS 0.007169f
C135 B.n28 VSUBS 0.007169f
C136 B.n29 VSUBS 0.007169f
C137 B.n30 VSUBS 0.007169f
C138 B.n31 VSUBS 0.007169f
C139 B.n32 VSUBS 0.007169f
C140 B.n33 VSUBS 0.007169f
C141 B.n34 VSUBS 0.007169f
C142 B.n35 VSUBS 0.007169f
C143 B.n36 VSUBS 0.007169f
C144 B.n37 VSUBS 0.007169f
C145 B.n38 VSUBS 0.007169f
C146 B.n39 VSUBS 0.007169f
C147 B.n40 VSUBS 0.007169f
C148 B.n41 VSUBS 0.007169f
C149 B.n42 VSUBS 0.007169f
C150 B.n43 VSUBS 0.007169f
C151 B.t5 VSUBS 0.37095f
C152 B.t4 VSUBS 0.388628f
C153 B.t3 VSUBS 1.06359f
C154 B.n44 VSUBS 0.192172f
C155 B.n45 VSUBS 0.071191f
C156 B.n46 VSUBS 0.007169f
C157 B.n47 VSUBS 0.007169f
C158 B.n48 VSUBS 0.007169f
C159 B.n49 VSUBS 0.007169f
C160 B.t11 VSUBS 0.370944f
C161 B.t10 VSUBS 0.388623f
C162 B.t9 VSUBS 1.06359f
C163 B.n50 VSUBS 0.192178f
C164 B.n51 VSUBS 0.071197f
C165 B.n52 VSUBS 0.016611f
C166 B.n53 VSUBS 0.007169f
C167 B.n54 VSUBS 0.007169f
C168 B.n55 VSUBS 0.007169f
C169 B.n56 VSUBS 0.007169f
C170 B.n57 VSUBS 0.007169f
C171 B.n58 VSUBS 0.007169f
C172 B.n59 VSUBS 0.007169f
C173 B.n60 VSUBS 0.007169f
C174 B.n61 VSUBS 0.007169f
C175 B.n62 VSUBS 0.007169f
C176 B.n63 VSUBS 0.007169f
C177 B.n64 VSUBS 0.007169f
C178 B.n65 VSUBS 0.007169f
C179 B.n66 VSUBS 0.007169f
C180 B.n67 VSUBS 0.007169f
C181 B.n68 VSUBS 0.007169f
C182 B.n69 VSUBS 0.007169f
C183 B.n70 VSUBS 0.007169f
C184 B.n71 VSUBS 0.007169f
C185 B.n72 VSUBS 0.018092f
C186 B.n73 VSUBS 0.007169f
C187 B.n74 VSUBS 0.007169f
C188 B.n75 VSUBS 0.007169f
C189 B.n76 VSUBS 0.007169f
C190 B.n77 VSUBS 0.007169f
C191 B.n78 VSUBS 0.007169f
C192 B.n79 VSUBS 0.007169f
C193 B.n80 VSUBS 0.007169f
C194 B.n81 VSUBS 0.007169f
C195 B.n82 VSUBS 0.007169f
C196 B.n83 VSUBS 0.007169f
C197 B.n84 VSUBS 0.007169f
C198 B.n85 VSUBS 0.007169f
C199 B.n86 VSUBS 0.007169f
C200 B.n87 VSUBS 0.007169f
C201 B.n88 VSUBS 0.007169f
C202 B.n89 VSUBS 0.007169f
C203 B.n90 VSUBS 0.007169f
C204 B.n91 VSUBS 0.007169f
C205 B.n92 VSUBS 0.007169f
C206 B.n93 VSUBS 0.007169f
C207 B.n94 VSUBS 0.007169f
C208 B.n95 VSUBS 0.007169f
C209 B.n96 VSUBS 0.007169f
C210 B.n97 VSUBS 0.007169f
C211 B.n98 VSUBS 0.007169f
C212 B.n99 VSUBS 0.007169f
C213 B.n100 VSUBS 0.007169f
C214 B.n101 VSUBS 0.007169f
C215 B.n102 VSUBS 0.007169f
C216 B.n103 VSUBS 0.007169f
C217 B.n104 VSUBS 0.007169f
C218 B.n105 VSUBS 0.007169f
C219 B.n106 VSUBS 0.007169f
C220 B.n107 VSUBS 0.007169f
C221 B.n108 VSUBS 0.007169f
C222 B.n109 VSUBS 0.007169f
C223 B.n110 VSUBS 0.007169f
C224 B.n111 VSUBS 0.007169f
C225 B.n112 VSUBS 0.007169f
C226 B.n113 VSUBS 0.007169f
C227 B.n114 VSUBS 0.007169f
C228 B.n115 VSUBS 0.017318f
C229 B.n116 VSUBS 0.007169f
C230 B.n117 VSUBS 0.007169f
C231 B.n118 VSUBS 0.007169f
C232 B.n119 VSUBS 0.007169f
C233 B.n120 VSUBS 0.007169f
C234 B.n121 VSUBS 0.007169f
C235 B.n122 VSUBS 0.007169f
C236 B.n123 VSUBS 0.007169f
C237 B.n124 VSUBS 0.007169f
C238 B.n125 VSUBS 0.007169f
C239 B.n126 VSUBS 0.007169f
C240 B.n127 VSUBS 0.007169f
C241 B.n128 VSUBS 0.007169f
C242 B.n129 VSUBS 0.007169f
C243 B.n130 VSUBS 0.007169f
C244 B.n131 VSUBS 0.007169f
C245 B.n132 VSUBS 0.007169f
C246 B.n133 VSUBS 0.007169f
C247 B.n134 VSUBS 0.007169f
C248 B.n135 VSUBS 0.007169f
C249 B.t1 VSUBS 0.370944f
C250 B.t2 VSUBS 0.388623f
C251 B.t0 VSUBS 1.06359f
C252 B.n136 VSUBS 0.192178f
C253 B.n137 VSUBS 0.071197f
C254 B.n138 VSUBS 0.007169f
C255 B.n139 VSUBS 0.007169f
C256 B.n140 VSUBS 0.007169f
C257 B.n141 VSUBS 0.007169f
C258 B.t7 VSUBS 0.37095f
C259 B.t8 VSUBS 0.388628f
C260 B.t6 VSUBS 1.06359f
C261 B.n142 VSUBS 0.192172f
C262 B.n143 VSUBS 0.071191f
C263 B.n144 VSUBS 0.016611f
C264 B.n145 VSUBS 0.007169f
C265 B.n146 VSUBS 0.007169f
C266 B.n147 VSUBS 0.007169f
C267 B.n148 VSUBS 0.007169f
C268 B.n149 VSUBS 0.007169f
C269 B.n150 VSUBS 0.007169f
C270 B.n151 VSUBS 0.007169f
C271 B.n152 VSUBS 0.007169f
C272 B.n153 VSUBS 0.007169f
C273 B.n154 VSUBS 0.007169f
C274 B.n155 VSUBS 0.007169f
C275 B.n156 VSUBS 0.007169f
C276 B.n157 VSUBS 0.007169f
C277 B.n158 VSUBS 0.007169f
C278 B.n159 VSUBS 0.007169f
C279 B.n160 VSUBS 0.007169f
C280 B.n161 VSUBS 0.007169f
C281 B.n162 VSUBS 0.007169f
C282 B.n163 VSUBS 0.007169f
C283 B.n164 VSUBS 0.017318f
C284 B.n165 VSUBS 0.007169f
C285 B.n166 VSUBS 0.007169f
C286 B.n167 VSUBS 0.007169f
C287 B.n168 VSUBS 0.007169f
C288 B.n169 VSUBS 0.007169f
C289 B.n170 VSUBS 0.007169f
C290 B.n171 VSUBS 0.007169f
C291 B.n172 VSUBS 0.007169f
C292 B.n173 VSUBS 0.007169f
C293 B.n174 VSUBS 0.007169f
C294 B.n175 VSUBS 0.007169f
C295 B.n176 VSUBS 0.007169f
C296 B.n177 VSUBS 0.007169f
C297 B.n178 VSUBS 0.007169f
C298 B.n179 VSUBS 0.007169f
C299 B.n180 VSUBS 0.007169f
C300 B.n181 VSUBS 0.007169f
C301 B.n182 VSUBS 0.007169f
C302 B.n183 VSUBS 0.007169f
C303 B.n184 VSUBS 0.007169f
C304 B.n185 VSUBS 0.007169f
C305 B.n186 VSUBS 0.007169f
C306 B.n187 VSUBS 0.007169f
C307 B.n188 VSUBS 0.007169f
C308 B.n189 VSUBS 0.007169f
C309 B.n190 VSUBS 0.007169f
C310 B.n191 VSUBS 0.007169f
C311 B.n192 VSUBS 0.007169f
C312 B.n193 VSUBS 0.007169f
C313 B.n194 VSUBS 0.007169f
C314 B.n195 VSUBS 0.007169f
C315 B.n196 VSUBS 0.007169f
C316 B.n197 VSUBS 0.007169f
C317 B.n198 VSUBS 0.007169f
C318 B.n199 VSUBS 0.007169f
C319 B.n200 VSUBS 0.007169f
C320 B.n201 VSUBS 0.007169f
C321 B.n202 VSUBS 0.007169f
C322 B.n203 VSUBS 0.007169f
C323 B.n204 VSUBS 0.007169f
C324 B.n205 VSUBS 0.007169f
C325 B.n206 VSUBS 0.007169f
C326 B.n207 VSUBS 0.007169f
C327 B.n208 VSUBS 0.007169f
C328 B.n209 VSUBS 0.007169f
C329 B.n210 VSUBS 0.007169f
C330 B.n211 VSUBS 0.007169f
C331 B.n212 VSUBS 0.007169f
C332 B.n213 VSUBS 0.007169f
C333 B.n214 VSUBS 0.007169f
C334 B.n215 VSUBS 0.007169f
C335 B.n216 VSUBS 0.007169f
C336 B.n217 VSUBS 0.007169f
C337 B.n218 VSUBS 0.007169f
C338 B.n219 VSUBS 0.007169f
C339 B.n220 VSUBS 0.007169f
C340 B.n221 VSUBS 0.007169f
C341 B.n222 VSUBS 0.007169f
C342 B.n223 VSUBS 0.007169f
C343 B.n224 VSUBS 0.007169f
C344 B.n225 VSUBS 0.007169f
C345 B.n226 VSUBS 0.007169f
C346 B.n227 VSUBS 0.007169f
C347 B.n228 VSUBS 0.007169f
C348 B.n229 VSUBS 0.007169f
C349 B.n230 VSUBS 0.007169f
C350 B.n231 VSUBS 0.007169f
C351 B.n232 VSUBS 0.007169f
C352 B.n233 VSUBS 0.007169f
C353 B.n234 VSUBS 0.007169f
C354 B.n235 VSUBS 0.007169f
C355 B.n236 VSUBS 0.007169f
C356 B.n237 VSUBS 0.007169f
C357 B.n238 VSUBS 0.007169f
C358 B.n239 VSUBS 0.007169f
C359 B.n240 VSUBS 0.007169f
C360 B.n241 VSUBS 0.007169f
C361 B.n242 VSUBS 0.007169f
C362 B.n243 VSUBS 0.007169f
C363 B.n244 VSUBS 0.007169f
C364 B.n245 VSUBS 0.007169f
C365 B.n246 VSUBS 0.007169f
C366 B.n247 VSUBS 0.017318f
C367 B.n248 VSUBS 0.018318f
C368 B.n249 VSUBS 0.018318f
C369 B.n250 VSUBS 0.007169f
C370 B.n251 VSUBS 0.007169f
C371 B.n252 VSUBS 0.007169f
C372 B.n253 VSUBS 0.007169f
C373 B.n254 VSUBS 0.007169f
C374 B.n255 VSUBS 0.007169f
C375 B.n256 VSUBS 0.007169f
C376 B.n257 VSUBS 0.007169f
C377 B.n258 VSUBS 0.007169f
C378 B.n259 VSUBS 0.007169f
C379 B.n260 VSUBS 0.007169f
C380 B.n261 VSUBS 0.007169f
C381 B.n262 VSUBS 0.007169f
C382 B.n263 VSUBS 0.007169f
C383 B.n264 VSUBS 0.007169f
C384 B.n265 VSUBS 0.007169f
C385 B.n266 VSUBS 0.007169f
C386 B.n267 VSUBS 0.007169f
C387 B.n268 VSUBS 0.007169f
C388 B.n269 VSUBS 0.007169f
C389 B.n270 VSUBS 0.007169f
C390 B.n271 VSUBS 0.007169f
C391 B.n272 VSUBS 0.007169f
C392 B.n273 VSUBS 0.007169f
C393 B.n274 VSUBS 0.007169f
C394 B.n275 VSUBS 0.007169f
C395 B.n276 VSUBS 0.007169f
C396 B.n277 VSUBS 0.007169f
C397 B.n278 VSUBS 0.007169f
C398 B.n279 VSUBS 0.007169f
C399 B.n280 VSUBS 0.007169f
C400 B.n281 VSUBS 0.007169f
C401 B.n282 VSUBS 0.007169f
C402 B.n283 VSUBS 0.007169f
C403 B.n284 VSUBS 0.007169f
C404 B.n285 VSUBS 0.007169f
C405 B.n286 VSUBS 0.007169f
C406 B.n287 VSUBS 0.007169f
C407 B.n288 VSUBS 0.007169f
C408 B.n289 VSUBS 0.007169f
C409 B.n290 VSUBS 0.007169f
C410 B.n291 VSUBS 0.007169f
C411 B.n292 VSUBS 0.007169f
C412 B.n293 VSUBS 0.007169f
C413 B.n294 VSUBS 0.007169f
C414 B.n295 VSUBS 0.007169f
C415 B.n296 VSUBS 0.007169f
C416 B.n297 VSUBS 0.007169f
C417 B.n298 VSUBS 0.007169f
C418 B.n299 VSUBS 0.007169f
C419 B.n300 VSUBS 0.007169f
C420 B.n301 VSUBS 0.007169f
C421 B.n302 VSUBS 0.007169f
C422 B.n303 VSUBS 0.007169f
C423 B.n304 VSUBS 0.007169f
C424 B.n305 VSUBS 0.006748f
C425 B.n306 VSUBS 0.007169f
C426 B.n307 VSUBS 0.007169f
C427 B.n308 VSUBS 0.004006f
C428 B.n309 VSUBS 0.007169f
C429 B.n310 VSUBS 0.007169f
C430 B.n311 VSUBS 0.007169f
C431 B.n312 VSUBS 0.007169f
C432 B.n313 VSUBS 0.007169f
C433 B.n314 VSUBS 0.007169f
C434 B.n315 VSUBS 0.007169f
C435 B.n316 VSUBS 0.007169f
C436 B.n317 VSUBS 0.007169f
C437 B.n318 VSUBS 0.007169f
C438 B.n319 VSUBS 0.007169f
C439 B.n320 VSUBS 0.007169f
C440 B.n321 VSUBS 0.004006f
C441 B.n322 VSUBS 0.016611f
C442 B.n323 VSUBS 0.006748f
C443 B.n324 VSUBS 0.007169f
C444 B.n325 VSUBS 0.007169f
C445 B.n326 VSUBS 0.007169f
C446 B.n327 VSUBS 0.007169f
C447 B.n328 VSUBS 0.007169f
C448 B.n329 VSUBS 0.007169f
C449 B.n330 VSUBS 0.007169f
C450 B.n331 VSUBS 0.007169f
C451 B.n332 VSUBS 0.007169f
C452 B.n333 VSUBS 0.007169f
C453 B.n334 VSUBS 0.007169f
C454 B.n335 VSUBS 0.007169f
C455 B.n336 VSUBS 0.007169f
C456 B.n337 VSUBS 0.007169f
C457 B.n338 VSUBS 0.007169f
C458 B.n339 VSUBS 0.007169f
C459 B.n340 VSUBS 0.007169f
C460 B.n341 VSUBS 0.007169f
C461 B.n342 VSUBS 0.007169f
C462 B.n343 VSUBS 0.007169f
C463 B.n344 VSUBS 0.007169f
C464 B.n345 VSUBS 0.007169f
C465 B.n346 VSUBS 0.007169f
C466 B.n347 VSUBS 0.007169f
C467 B.n348 VSUBS 0.007169f
C468 B.n349 VSUBS 0.007169f
C469 B.n350 VSUBS 0.007169f
C470 B.n351 VSUBS 0.007169f
C471 B.n352 VSUBS 0.007169f
C472 B.n353 VSUBS 0.007169f
C473 B.n354 VSUBS 0.007169f
C474 B.n355 VSUBS 0.007169f
C475 B.n356 VSUBS 0.007169f
C476 B.n357 VSUBS 0.007169f
C477 B.n358 VSUBS 0.007169f
C478 B.n359 VSUBS 0.007169f
C479 B.n360 VSUBS 0.007169f
C480 B.n361 VSUBS 0.007169f
C481 B.n362 VSUBS 0.007169f
C482 B.n363 VSUBS 0.007169f
C483 B.n364 VSUBS 0.007169f
C484 B.n365 VSUBS 0.007169f
C485 B.n366 VSUBS 0.007169f
C486 B.n367 VSUBS 0.007169f
C487 B.n368 VSUBS 0.007169f
C488 B.n369 VSUBS 0.007169f
C489 B.n370 VSUBS 0.007169f
C490 B.n371 VSUBS 0.007169f
C491 B.n372 VSUBS 0.007169f
C492 B.n373 VSUBS 0.007169f
C493 B.n374 VSUBS 0.007169f
C494 B.n375 VSUBS 0.007169f
C495 B.n376 VSUBS 0.007169f
C496 B.n377 VSUBS 0.007169f
C497 B.n378 VSUBS 0.007169f
C498 B.n379 VSUBS 0.007169f
C499 B.n380 VSUBS 0.018318f
C500 B.n381 VSUBS 0.018318f
C501 B.n382 VSUBS 0.017318f
C502 B.n383 VSUBS 0.007169f
C503 B.n384 VSUBS 0.007169f
C504 B.n385 VSUBS 0.007169f
C505 B.n386 VSUBS 0.007169f
C506 B.n387 VSUBS 0.007169f
C507 B.n388 VSUBS 0.007169f
C508 B.n389 VSUBS 0.007169f
C509 B.n390 VSUBS 0.007169f
C510 B.n391 VSUBS 0.007169f
C511 B.n392 VSUBS 0.007169f
C512 B.n393 VSUBS 0.007169f
C513 B.n394 VSUBS 0.007169f
C514 B.n395 VSUBS 0.007169f
C515 B.n396 VSUBS 0.007169f
C516 B.n397 VSUBS 0.007169f
C517 B.n398 VSUBS 0.007169f
C518 B.n399 VSUBS 0.007169f
C519 B.n400 VSUBS 0.007169f
C520 B.n401 VSUBS 0.007169f
C521 B.n402 VSUBS 0.007169f
C522 B.n403 VSUBS 0.007169f
C523 B.n404 VSUBS 0.007169f
C524 B.n405 VSUBS 0.007169f
C525 B.n406 VSUBS 0.007169f
C526 B.n407 VSUBS 0.007169f
C527 B.n408 VSUBS 0.007169f
C528 B.n409 VSUBS 0.007169f
C529 B.n410 VSUBS 0.007169f
C530 B.n411 VSUBS 0.007169f
C531 B.n412 VSUBS 0.007169f
C532 B.n413 VSUBS 0.007169f
C533 B.n414 VSUBS 0.007169f
C534 B.n415 VSUBS 0.007169f
C535 B.n416 VSUBS 0.007169f
C536 B.n417 VSUBS 0.007169f
C537 B.n418 VSUBS 0.007169f
C538 B.n419 VSUBS 0.007169f
C539 B.n420 VSUBS 0.007169f
C540 B.n421 VSUBS 0.007169f
C541 B.n422 VSUBS 0.007169f
C542 B.n423 VSUBS 0.007169f
C543 B.n424 VSUBS 0.007169f
C544 B.n425 VSUBS 0.007169f
C545 B.n426 VSUBS 0.007169f
C546 B.n427 VSUBS 0.007169f
C547 B.n428 VSUBS 0.007169f
C548 B.n429 VSUBS 0.007169f
C549 B.n430 VSUBS 0.007169f
C550 B.n431 VSUBS 0.007169f
C551 B.n432 VSUBS 0.007169f
C552 B.n433 VSUBS 0.007169f
C553 B.n434 VSUBS 0.007169f
C554 B.n435 VSUBS 0.007169f
C555 B.n436 VSUBS 0.007169f
C556 B.n437 VSUBS 0.007169f
C557 B.n438 VSUBS 0.007169f
C558 B.n439 VSUBS 0.007169f
C559 B.n440 VSUBS 0.007169f
C560 B.n441 VSUBS 0.007169f
C561 B.n442 VSUBS 0.007169f
C562 B.n443 VSUBS 0.007169f
C563 B.n444 VSUBS 0.007169f
C564 B.n445 VSUBS 0.007169f
C565 B.n446 VSUBS 0.007169f
C566 B.n447 VSUBS 0.007169f
C567 B.n448 VSUBS 0.007169f
C568 B.n449 VSUBS 0.007169f
C569 B.n450 VSUBS 0.007169f
C570 B.n451 VSUBS 0.007169f
C571 B.n452 VSUBS 0.007169f
C572 B.n453 VSUBS 0.007169f
C573 B.n454 VSUBS 0.007169f
C574 B.n455 VSUBS 0.007169f
C575 B.n456 VSUBS 0.007169f
C576 B.n457 VSUBS 0.007169f
C577 B.n458 VSUBS 0.007169f
C578 B.n459 VSUBS 0.007169f
C579 B.n460 VSUBS 0.007169f
C580 B.n461 VSUBS 0.007169f
C581 B.n462 VSUBS 0.007169f
C582 B.n463 VSUBS 0.007169f
C583 B.n464 VSUBS 0.007169f
C584 B.n465 VSUBS 0.007169f
C585 B.n466 VSUBS 0.007169f
C586 B.n467 VSUBS 0.007169f
C587 B.n468 VSUBS 0.007169f
C588 B.n469 VSUBS 0.007169f
C589 B.n470 VSUBS 0.007169f
C590 B.n471 VSUBS 0.007169f
C591 B.n472 VSUBS 0.007169f
C592 B.n473 VSUBS 0.007169f
C593 B.n474 VSUBS 0.007169f
C594 B.n475 VSUBS 0.007169f
C595 B.n476 VSUBS 0.007169f
C596 B.n477 VSUBS 0.007169f
C597 B.n478 VSUBS 0.007169f
C598 B.n479 VSUBS 0.007169f
C599 B.n480 VSUBS 0.007169f
C600 B.n481 VSUBS 0.007169f
C601 B.n482 VSUBS 0.007169f
C602 B.n483 VSUBS 0.007169f
C603 B.n484 VSUBS 0.007169f
C604 B.n485 VSUBS 0.007169f
C605 B.n486 VSUBS 0.007169f
C606 B.n487 VSUBS 0.007169f
C607 B.n488 VSUBS 0.007169f
C608 B.n489 VSUBS 0.007169f
C609 B.n490 VSUBS 0.007169f
C610 B.n491 VSUBS 0.007169f
C611 B.n492 VSUBS 0.007169f
C612 B.n493 VSUBS 0.007169f
C613 B.n494 VSUBS 0.007169f
C614 B.n495 VSUBS 0.007169f
C615 B.n496 VSUBS 0.007169f
C616 B.n497 VSUBS 0.007169f
C617 B.n498 VSUBS 0.007169f
C618 B.n499 VSUBS 0.007169f
C619 B.n500 VSUBS 0.007169f
C620 B.n501 VSUBS 0.007169f
C621 B.n502 VSUBS 0.007169f
C622 B.n503 VSUBS 0.007169f
C623 B.n504 VSUBS 0.007169f
C624 B.n505 VSUBS 0.007169f
C625 B.n506 VSUBS 0.007169f
C626 B.n507 VSUBS 0.007169f
C627 B.n508 VSUBS 0.007169f
C628 B.n509 VSUBS 0.007169f
C629 B.n510 VSUBS 0.007169f
C630 B.n511 VSUBS 0.017318f
C631 B.n512 VSUBS 0.018318f
C632 B.n513 VSUBS 0.017544f
C633 B.n514 VSUBS 0.007169f
C634 B.n515 VSUBS 0.007169f
C635 B.n516 VSUBS 0.007169f
C636 B.n517 VSUBS 0.007169f
C637 B.n518 VSUBS 0.007169f
C638 B.n519 VSUBS 0.007169f
C639 B.n520 VSUBS 0.007169f
C640 B.n521 VSUBS 0.007169f
C641 B.n522 VSUBS 0.007169f
C642 B.n523 VSUBS 0.007169f
C643 B.n524 VSUBS 0.007169f
C644 B.n525 VSUBS 0.007169f
C645 B.n526 VSUBS 0.007169f
C646 B.n527 VSUBS 0.007169f
C647 B.n528 VSUBS 0.007169f
C648 B.n529 VSUBS 0.007169f
C649 B.n530 VSUBS 0.007169f
C650 B.n531 VSUBS 0.007169f
C651 B.n532 VSUBS 0.007169f
C652 B.n533 VSUBS 0.007169f
C653 B.n534 VSUBS 0.007169f
C654 B.n535 VSUBS 0.007169f
C655 B.n536 VSUBS 0.007169f
C656 B.n537 VSUBS 0.007169f
C657 B.n538 VSUBS 0.007169f
C658 B.n539 VSUBS 0.007169f
C659 B.n540 VSUBS 0.007169f
C660 B.n541 VSUBS 0.007169f
C661 B.n542 VSUBS 0.007169f
C662 B.n543 VSUBS 0.007169f
C663 B.n544 VSUBS 0.007169f
C664 B.n545 VSUBS 0.007169f
C665 B.n546 VSUBS 0.007169f
C666 B.n547 VSUBS 0.007169f
C667 B.n548 VSUBS 0.007169f
C668 B.n549 VSUBS 0.007169f
C669 B.n550 VSUBS 0.007169f
C670 B.n551 VSUBS 0.007169f
C671 B.n552 VSUBS 0.007169f
C672 B.n553 VSUBS 0.007169f
C673 B.n554 VSUBS 0.007169f
C674 B.n555 VSUBS 0.007169f
C675 B.n556 VSUBS 0.007169f
C676 B.n557 VSUBS 0.007169f
C677 B.n558 VSUBS 0.007169f
C678 B.n559 VSUBS 0.007169f
C679 B.n560 VSUBS 0.007169f
C680 B.n561 VSUBS 0.007169f
C681 B.n562 VSUBS 0.007169f
C682 B.n563 VSUBS 0.007169f
C683 B.n564 VSUBS 0.007169f
C684 B.n565 VSUBS 0.007169f
C685 B.n566 VSUBS 0.007169f
C686 B.n567 VSUBS 0.007169f
C687 B.n568 VSUBS 0.007169f
C688 B.n569 VSUBS 0.006748f
C689 B.n570 VSUBS 0.007169f
C690 B.n571 VSUBS 0.007169f
C691 B.n572 VSUBS 0.004006f
C692 B.n573 VSUBS 0.007169f
C693 B.n574 VSUBS 0.007169f
C694 B.n575 VSUBS 0.007169f
C695 B.n576 VSUBS 0.007169f
C696 B.n577 VSUBS 0.007169f
C697 B.n578 VSUBS 0.007169f
C698 B.n579 VSUBS 0.007169f
C699 B.n580 VSUBS 0.007169f
C700 B.n581 VSUBS 0.007169f
C701 B.n582 VSUBS 0.007169f
C702 B.n583 VSUBS 0.007169f
C703 B.n584 VSUBS 0.007169f
C704 B.n585 VSUBS 0.004006f
C705 B.n586 VSUBS 0.016611f
C706 B.n587 VSUBS 0.006748f
C707 B.n588 VSUBS 0.007169f
C708 B.n589 VSUBS 0.007169f
C709 B.n590 VSUBS 0.007169f
C710 B.n591 VSUBS 0.007169f
C711 B.n592 VSUBS 0.007169f
C712 B.n593 VSUBS 0.007169f
C713 B.n594 VSUBS 0.007169f
C714 B.n595 VSUBS 0.007169f
C715 B.n596 VSUBS 0.007169f
C716 B.n597 VSUBS 0.007169f
C717 B.n598 VSUBS 0.007169f
C718 B.n599 VSUBS 0.007169f
C719 B.n600 VSUBS 0.007169f
C720 B.n601 VSUBS 0.007169f
C721 B.n602 VSUBS 0.007169f
C722 B.n603 VSUBS 0.007169f
C723 B.n604 VSUBS 0.007169f
C724 B.n605 VSUBS 0.007169f
C725 B.n606 VSUBS 0.007169f
C726 B.n607 VSUBS 0.007169f
C727 B.n608 VSUBS 0.007169f
C728 B.n609 VSUBS 0.007169f
C729 B.n610 VSUBS 0.007169f
C730 B.n611 VSUBS 0.007169f
C731 B.n612 VSUBS 0.007169f
C732 B.n613 VSUBS 0.007169f
C733 B.n614 VSUBS 0.007169f
C734 B.n615 VSUBS 0.007169f
C735 B.n616 VSUBS 0.007169f
C736 B.n617 VSUBS 0.007169f
C737 B.n618 VSUBS 0.007169f
C738 B.n619 VSUBS 0.007169f
C739 B.n620 VSUBS 0.007169f
C740 B.n621 VSUBS 0.007169f
C741 B.n622 VSUBS 0.007169f
C742 B.n623 VSUBS 0.007169f
C743 B.n624 VSUBS 0.007169f
C744 B.n625 VSUBS 0.007169f
C745 B.n626 VSUBS 0.007169f
C746 B.n627 VSUBS 0.007169f
C747 B.n628 VSUBS 0.007169f
C748 B.n629 VSUBS 0.007169f
C749 B.n630 VSUBS 0.007169f
C750 B.n631 VSUBS 0.007169f
C751 B.n632 VSUBS 0.007169f
C752 B.n633 VSUBS 0.007169f
C753 B.n634 VSUBS 0.007169f
C754 B.n635 VSUBS 0.007169f
C755 B.n636 VSUBS 0.007169f
C756 B.n637 VSUBS 0.007169f
C757 B.n638 VSUBS 0.007169f
C758 B.n639 VSUBS 0.007169f
C759 B.n640 VSUBS 0.007169f
C760 B.n641 VSUBS 0.007169f
C761 B.n642 VSUBS 0.007169f
C762 B.n643 VSUBS 0.007169f
C763 B.n644 VSUBS 0.018318f
C764 B.n645 VSUBS 0.018318f
C765 B.n646 VSUBS 0.017318f
C766 B.n647 VSUBS 0.007169f
C767 B.n648 VSUBS 0.007169f
C768 B.n649 VSUBS 0.007169f
C769 B.n650 VSUBS 0.007169f
C770 B.n651 VSUBS 0.007169f
C771 B.n652 VSUBS 0.007169f
C772 B.n653 VSUBS 0.007169f
C773 B.n654 VSUBS 0.007169f
C774 B.n655 VSUBS 0.007169f
C775 B.n656 VSUBS 0.007169f
C776 B.n657 VSUBS 0.007169f
C777 B.n658 VSUBS 0.007169f
C778 B.n659 VSUBS 0.007169f
C779 B.n660 VSUBS 0.007169f
C780 B.n661 VSUBS 0.007169f
C781 B.n662 VSUBS 0.007169f
C782 B.n663 VSUBS 0.007169f
C783 B.n664 VSUBS 0.007169f
C784 B.n665 VSUBS 0.007169f
C785 B.n666 VSUBS 0.007169f
C786 B.n667 VSUBS 0.007169f
C787 B.n668 VSUBS 0.007169f
C788 B.n669 VSUBS 0.007169f
C789 B.n670 VSUBS 0.007169f
C790 B.n671 VSUBS 0.007169f
C791 B.n672 VSUBS 0.007169f
C792 B.n673 VSUBS 0.007169f
C793 B.n674 VSUBS 0.007169f
C794 B.n675 VSUBS 0.007169f
C795 B.n676 VSUBS 0.007169f
C796 B.n677 VSUBS 0.007169f
C797 B.n678 VSUBS 0.007169f
C798 B.n679 VSUBS 0.007169f
C799 B.n680 VSUBS 0.007169f
C800 B.n681 VSUBS 0.007169f
C801 B.n682 VSUBS 0.007169f
C802 B.n683 VSUBS 0.007169f
C803 B.n684 VSUBS 0.007169f
C804 B.n685 VSUBS 0.007169f
C805 B.n686 VSUBS 0.007169f
C806 B.n687 VSUBS 0.007169f
C807 B.n688 VSUBS 0.007169f
C808 B.n689 VSUBS 0.007169f
C809 B.n690 VSUBS 0.007169f
C810 B.n691 VSUBS 0.007169f
C811 B.n692 VSUBS 0.007169f
C812 B.n693 VSUBS 0.007169f
C813 B.n694 VSUBS 0.007169f
C814 B.n695 VSUBS 0.007169f
C815 B.n696 VSUBS 0.007169f
C816 B.n697 VSUBS 0.007169f
C817 B.n698 VSUBS 0.007169f
C818 B.n699 VSUBS 0.007169f
C819 B.n700 VSUBS 0.007169f
C820 B.n701 VSUBS 0.007169f
C821 B.n702 VSUBS 0.007169f
C822 B.n703 VSUBS 0.007169f
C823 B.n704 VSUBS 0.007169f
C824 B.n705 VSUBS 0.007169f
C825 B.n706 VSUBS 0.007169f
C826 B.n707 VSUBS 0.007169f
C827 B.n708 VSUBS 0.007169f
C828 B.n709 VSUBS 0.007169f
C829 B.n710 VSUBS 0.007169f
C830 B.n711 VSUBS 0.016234f
C831 VTAIL.t11 VSUBS 0.220945f
C832 VTAIL.t13 VSUBS 0.220945f
C833 VTAIL.n0 VSUBS 1.59189f
C834 VTAIL.n1 VSUBS 0.71044f
C835 VTAIL.t8 VSUBS 2.10584f
C836 VTAIL.n2 VSUBS 0.832177f
C837 VTAIL.t7 VSUBS 2.10584f
C838 VTAIL.n3 VSUBS 0.832177f
C839 VTAIL.t5 VSUBS 0.220945f
C840 VTAIL.t1 VSUBS 0.220945f
C841 VTAIL.n4 VSUBS 1.59189f
C842 VTAIL.n5 VSUBS 0.871492f
C843 VTAIL.t3 VSUBS 2.10584f
C844 VTAIL.n6 VSUBS 2.07588f
C845 VTAIL.t14 VSUBS 2.10585f
C846 VTAIL.n7 VSUBS 2.07586f
C847 VTAIL.t10 VSUBS 0.220945f
C848 VTAIL.t15 VSUBS 0.220945f
C849 VTAIL.n8 VSUBS 1.59189f
C850 VTAIL.n9 VSUBS 0.871486f
C851 VTAIL.t12 VSUBS 2.10585f
C852 VTAIL.n10 VSUBS 0.832163f
C853 VTAIL.t6 VSUBS 2.10585f
C854 VTAIL.n11 VSUBS 0.832163f
C855 VTAIL.t0 VSUBS 0.220945f
C856 VTAIL.t2 VSUBS 0.220945f
C857 VTAIL.n12 VSUBS 1.59189f
C858 VTAIL.n13 VSUBS 0.871486f
C859 VTAIL.t4 VSUBS 2.10584f
C860 VTAIL.n14 VSUBS 2.07588f
C861 VTAIL.t9 VSUBS 2.10584f
C862 VTAIL.n15 VSUBS 2.0712f
C863 VDD2.t5 VSUBS 0.215982f
C864 VDD2.t4 VSUBS 0.215982f
C865 VDD2.n0 VSUBS 1.68298f
C866 VDD2.t3 VSUBS 0.215982f
C867 VDD2.t2 VSUBS 0.215982f
C868 VDD2.n1 VSUBS 1.68298f
C869 VDD2.n2 VSUBS 3.32581f
C870 VDD2.t1 VSUBS 0.215982f
C871 VDD2.t0 VSUBS 0.215982f
C872 VDD2.n3 VSUBS 1.67449f
C873 VDD2.n4 VSUBS 2.87841f
C874 VDD2.t7 VSUBS 0.215982f
C875 VDD2.t6 VSUBS 0.215982f
C876 VDD2.n5 VSUBS 1.68295f
C877 VN.n0 VSUBS 0.044141f
C878 VN.t6 VSUBS 2.1005f
C879 VN.n1 VSUBS 0.036461f
C880 VN.n2 VSUBS 0.033482f
C881 VN.t2 VSUBS 2.1005f
C882 VN.n3 VSUBS 0.048672f
C883 VN.n4 VSUBS 0.280606f
C884 VN.t4 VSUBS 2.1005f
C885 VN.t7 VSUBS 2.28893f
C886 VN.n5 VSUBS 0.825297f
C887 VN.n6 VSUBS 0.846824f
C888 VN.n7 VSUBS 0.058719f
C889 VN.n8 VSUBS 0.048672f
C890 VN.n9 VSUBS 0.033482f
C891 VN.n10 VSUBS 0.033482f
C892 VN.n11 VSUBS 0.033482f
C893 VN.n12 VSUBS 0.058719f
C894 VN.n13 VSUBS 0.752296f
C895 VN.n14 VSUBS 0.03481f
C896 VN.n15 VSUBS 0.064564f
C897 VN.n16 VSUBS 0.033482f
C898 VN.n17 VSUBS 0.033482f
C899 VN.n18 VSUBS 0.033482f
C900 VN.n19 VSUBS 0.05841f
C901 VN.n20 VSUBS 0.051975f
C902 VN.n21 VSUBS 0.850708f
C903 VN.n22 VSUBS 0.044119f
C904 VN.n23 VSUBS 0.044141f
C905 VN.t1 VSUBS 2.1005f
C906 VN.n24 VSUBS 0.036461f
C907 VN.n25 VSUBS 0.033482f
C908 VN.t5 VSUBS 2.1005f
C909 VN.n26 VSUBS 0.048672f
C910 VN.n27 VSUBS 0.280606f
C911 VN.t0 VSUBS 2.1005f
C912 VN.t3 VSUBS 2.28893f
C913 VN.n28 VSUBS 0.825297f
C914 VN.n29 VSUBS 0.846824f
C915 VN.n30 VSUBS 0.058719f
C916 VN.n31 VSUBS 0.048672f
C917 VN.n32 VSUBS 0.033482f
C918 VN.n33 VSUBS 0.033482f
C919 VN.n34 VSUBS 0.033482f
C920 VN.n35 VSUBS 0.058719f
C921 VN.n36 VSUBS 0.752296f
C922 VN.n37 VSUBS 0.03481f
C923 VN.n38 VSUBS 0.064564f
C924 VN.n39 VSUBS 0.033482f
C925 VN.n40 VSUBS 0.033482f
C926 VN.n41 VSUBS 0.033482f
C927 VN.n42 VSUBS 0.05841f
C928 VN.n43 VSUBS 0.051975f
C929 VN.n44 VSUBS 0.850708f
C930 VN.n45 VSUBS 1.74627f
.ends

