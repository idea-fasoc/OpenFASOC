* NGSPICE file created from diff_pair_sample_0217.ext - technology: sky130A

.subckt diff_pair_sample_0217 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0.90915 ps=5.84 w=5.51 l=3.18
X1 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0 ps=0 w=5.51 l=3.18
X2 VDD1.t1 VP.t1 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=0.90915 pd=5.84 as=2.1489 ps=11.8 w=5.51 l=3.18
X3 VTAIL.t5 VP.t2 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0.90915 ps=5.84 w=5.51 l=3.18
X4 VDD2.t3 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.90915 pd=5.84 as=2.1489 ps=11.8 w=5.51 l=3.18
X5 VDD1.t0 VP.t3 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=0.90915 pd=5.84 as=2.1489 ps=11.8 w=5.51 l=3.18
X6 VDD2.t2 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.90915 pd=5.84 as=2.1489 ps=11.8 w=5.51 l=3.18
X7 VTAIL.t2 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0.90915 ps=5.84 w=5.51 l=3.18
X8 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0 ps=0 w=5.51 l=3.18
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0 ps=0 w=5.51 l=3.18
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0 ps=0 w=5.51 l=3.18
X11 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1489 pd=11.8 as=0.90915 ps=5.84 w=5.51 l=3.18
R0 VP.n17 VP.n16 161.3
R1 VP.n15 VP.n1 161.3
R2 VP.n14 VP.n13 161.3
R3 VP.n12 VP.n2 161.3
R4 VP.n11 VP.n10 161.3
R5 VP.n9 VP.n3 161.3
R6 VP.n8 VP.n7 161.3
R7 VP.n6 VP.n4 77.5892
R8 VP.n18 VP.n0 77.5892
R9 VP.n5 VP.t0 76.3397
R10 VP.n5 VP.t1 75.2492
R11 VP.n6 VP.n5 45.8061
R12 VP.n4 VP.t2 41.7587
R13 VP.n0 VP.t3 41.7587
R14 VP.n10 VP.n2 40.4934
R15 VP.n14 VP.n2 40.4934
R16 VP.n9 VP.n8 24.4675
R17 VP.n10 VP.n9 24.4675
R18 VP.n15 VP.n14 24.4675
R19 VP.n16 VP.n15 24.4675
R20 VP.n8 VP.n4 12.4787
R21 VP.n16 VP.n0 12.4787
R22 VP.n7 VP.n6 0.354971
R23 VP.n18 VP.n17 0.354971
R24 VP VP.n18 0.26696
R25 VP.n7 VP.n3 0.189894
R26 VP.n11 VP.n3 0.189894
R27 VP.n12 VP.n11 0.189894
R28 VP.n13 VP.n12 0.189894
R29 VP.n13 VP.n1 0.189894
R30 VP.n17 VP.n1 0.189894
R31 VDD1 VDD1.n1 109.495
R32 VDD1 VDD1.n0 71.4846
R33 VDD1.n0 VDD1.t2 3.59397
R34 VDD1.n0 VDD1.t1 3.59397
R35 VDD1.n1 VDD1.t3 3.59397
R36 VDD1.n1 VDD1.t0 3.59397
R37 VTAIL.n5 VTAIL.t7 58.342
R38 VTAIL.n4 VTAIL.t1 58.342
R39 VTAIL.n3 VTAIL.t3 58.342
R40 VTAIL.n6 VTAIL.t6 58.3411
R41 VTAIL.n7 VTAIL.t0 58.341
R42 VTAIL.n0 VTAIL.t2 58.341
R43 VTAIL.n1 VTAIL.t4 58.341
R44 VTAIL.n2 VTAIL.t5 58.341
R45 VTAIL.n7 VTAIL.n6 20.1427
R46 VTAIL.n3 VTAIL.n2 20.1427
R47 VTAIL.n4 VTAIL.n3 3.02636
R48 VTAIL.n6 VTAIL.n5 3.02636
R49 VTAIL.n2 VTAIL.n1 3.02636
R50 VTAIL VTAIL.n0 1.57162
R51 VTAIL VTAIL.n7 1.45524
R52 VTAIL.n5 VTAIL.n4 0.470328
R53 VTAIL.n1 VTAIL.n0 0.470328
R54 B.n598 B.n597 585
R55 B.n599 B.n598 585
R56 B.n211 B.n101 585
R57 B.n210 B.n209 585
R58 B.n208 B.n207 585
R59 B.n206 B.n205 585
R60 B.n204 B.n203 585
R61 B.n202 B.n201 585
R62 B.n200 B.n199 585
R63 B.n198 B.n197 585
R64 B.n196 B.n195 585
R65 B.n194 B.n193 585
R66 B.n192 B.n191 585
R67 B.n190 B.n189 585
R68 B.n188 B.n187 585
R69 B.n186 B.n185 585
R70 B.n184 B.n183 585
R71 B.n182 B.n181 585
R72 B.n180 B.n179 585
R73 B.n178 B.n177 585
R74 B.n176 B.n175 585
R75 B.n174 B.n173 585
R76 B.n172 B.n171 585
R77 B.n170 B.n169 585
R78 B.n168 B.n167 585
R79 B.n166 B.n165 585
R80 B.n164 B.n163 585
R81 B.n162 B.n161 585
R82 B.n160 B.n159 585
R83 B.n158 B.n157 585
R84 B.n156 B.n155 585
R85 B.n154 B.n153 585
R86 B.n152 B.n151 585
R87 B.n149 B.n148 585
R88 B.n147 B.n146 585
R89 B.n145 B.n144 585
R90 B.n143 B.n142 585
R91 B.n141 B.n140 585
R92 B.n139 B.n138 585
R93 B.n137 B.n136 585
R94 B.n135 B.n134 585
R95 B.n133 B.n132 585
R96 B.n131 B.n130 585
R97 B.n129 B.n128 585
R98 B.n127 B.n126 585
R99 B.n125 B.n124 585
R100 B.n123 B.n122 585
R101 B.n121 B.n120 585
R102 B.n119 B.n118 585
R103 B.n117 B.n116 585
R104 B.n115 B.n114 585
R105 B.n113 B.n112 585
R106 B.n111 B.n110 585
R107 B.n109 B.n108 585
R108 B.n74 B.n73 585
R109 B.n602 B.n601 585
R110 B.n596 B.n102 585
R111 B.n102 B.n71 585
R112 B.n595 B.n70 585
R113 B.n606 B.n70 585
R114 B.n594 B.n69 585
R115 B.n607 B.n69 585
R116 B.n593 B.n68 585
R117 B.n608 B.n68 585
R118 B.n592 B.n591 585
R119 B.n591 B.n64 585
R120 B.n590 B.n63 585
R121 B.n614 B.n63 585
R122 B.n589 B.n62 585
R123 B.n615 B.n62 585
R124 B.n588 B.n61 585
R125 B.n616 B.n61 585
R126 B.n587 B.n586 585
R127 B.n586 B.n60 585
R128 B.n585 B.n56 585
R129 B.n622 B.n56 585
R130 B.n584 B.n55 585
R131 B.n623 B.n55 585
R132 B.n583 B.n54 585
R133 B.n624 B.n54 585
R134 B.n582 B.n581 585
R135 B.n581 B.n50 585
R136 B.n580 B.n49 585
R137 B.n630 B.n49 585
R138 B.n579 B.n48 585
R139 B.n631 B.n48 585
R140 B.n578 B.n47 585
R141 B.n632 B.n47 585
R142 B.n577 B.n576 585
R143 B.n576 B.n43 585
R144 B.n575 B.n42 585
R145 B.n638 B.n42 585
R146 B.n574 B.n41 585
R147 B.n639 B.n41 585
R148 B.n573 B.n40 585
R149 B.n640 B.n40 585
R150 B.n572 B.n571 585
R151 B.n571 B.n36 585
R152 B.n570 B.n35 585
R153 B.n646 B.n35 585
R154 B.n569 B.n34 585
R155 B.n647 B.n34 585
R156 B.n568 B.n33 585
R157 B.n648 B.n33 585
R158 B.n567 B.n566 585
R159 B.n566 B.n29 585
R160 B.n565 B.n28 585
R161 B.n654 B.n28 585
R162 B.n564 B.n27 585
R163 B.n655 B.n27 585
R164 B.n563 B.n26 585
R165 B.n656 B.n26 585
R166 B.n562 B.n561 585
R167 B.n561 B.n22 585
R168 B.n560 B.n21 585
R169 B.n662 B.n21 585
R170 B.n559 B.n20 585
R171 B.n663 B.n20 585
R172 B.n558 B.n19 585
R173 B.n664 B.n19 585
R174 B.n557 B.n556 585
R175 B.n556 B.n18 585
R176 B.n555 B.n14 585
R177 B.n670 B.n14 585
R178 B.n554 B.n13 585
R179 B.n671 B.n13 585
R180 B.n553 B.n12 585
R181 B.n672 B.n12 585
R182 B.n552 B.n551 585
R183 B.n551 B.n8 585
R184 B.n550 B.n7 585
R185 B.n678 B.n7 585
R186 B.n549 B.n6 585
R187 B.n679 B.n6 585
R188 B.n548 B.n5 585
R189 B.n680 B.n5 585
R190 B.n547 B.n546 585
R191 B.n546 B.n4 585
R192 B.n545 B.n212 585
R193 B.n545 B.n544 585
R194 B.n535 B.n213 585
R195 B.n214 B.n213 585
R196 B.n537 B.n536 585
R197 B.n538 B.n537 585
R198 B.n534 B.n219 585
R199 B.n219 B.n218 585
R200 B.n533 B.n532 585
R201 B.n532 B.n531 585
R202 B.n221 B.n220 585
R203 B.n524 B.n221 585
R204 B.n523 B.n522 585
R205 B.n525 B.n523 585
R206 B.n521 B.n226 585
R207 B.n226 B.n225 585
R208 B.n520 B.n519 585
R209 B.n519 B.n518 585
R210 B.n228 B.n227 585
R211 B.n229 B.n228 585
R212 B.n511 B.n510 585
R213 B.n512 B.n511 585
R214 B.n509 B.n234 585
R215 B.n234 B.n233 585
R216 B.n508 B.n507 585
R217 B.n507 B.n506 585
R218 B.n236 B.n235 585
R219 B.n237 B.n236 585
R220 B.n499 B.n498 585
R221 B.n500 B.n499 585
R222 B.n497 B.n242 585
R223 B.n242 B.n241 585
R224 B.n496 B.n495 585
R225 B.n495 B.n494 585
R226 B.n244 B.n243 585
R227 B.n245 B.n244 585
R228 B.n487 B.n486 585
R229 B.n488 B.n487 585
R230 B.n485 B.n250 585
R231 B.n250 B.n249 585
R232 B.n484 B.n483 585
R233 B.n483 B.n482 585
R234 B.n252 B.n251 585
R235 B.n253 B.n252 585
R236 B.n475 B.n474 585
R237 B.n476 B.n475 585
R238 B.n473 B.n258 585
R239 B.n258 B.n257 585
R240 B.n472 B.n471 585
R241 B.n471 B.n470 585
R242 B.n260 B.n259 585
R243 B.n261 B.n260 585
R244 B.n463 B.n462 585
R245 B.n464 B.n463 585
R246 B.n461 B.n266 585
R247 B.n266 B.n265 585
R248 B.n460 B.n459 585
R249 B.n459 B.n458 585
R250 B.n268 B.n267 585
R251 B.n451 B.n268 585
R252 B.n450 B.n449 585
R253 B.n452 B.n450 585
R254 B.n448 B.n273 585
R255 B.n273 B.n272 585
R256 B.n447 B.n446 585
R257 B.n446 B.n445 585
R258 B.n275 B.n274 585
R259 B.n276 B.n275 585
R260 B.n438 B.n437 585
R261 B.n439 B.n438 585
R262 B.n436 B.n281 585
R263 B.n281 B.n280 585
R264 B.n435 B.n434 585
R265 B.n434 B.n433 585
R266 B.n283 B.n282 585
R267 B.n284 B.n283 585
R268 B.n429 B.n428 585
R269 B.n287 B.n286 585
R270 B.n425 B.n424 585
R271 B.n426 B.n425 585
R272 B.n423 B.n314 585
R273 B.n422 B.n421 585
R274 B.n420 B.n419 585
R275 B.n418 B.n417 585
R276 B.n416 B.n415 585
R277 B.n414 B.n413 585
R278 B.n412 B.n411 585
R279 B.n410 B.n409 585
R280 B.n408 B.n407 585
R281 B.n406 B.n405 585
R282 B.n404 B.n403 585
R283 B.n402 B.n401 585
R284 B.n400 B.n399 585
R285 B.n398 B.n397 585
R286 B.n396 B.n395 585
R287 B.n394 B.n393 585
R288 B.n392 B.n391 585
R289 B.n390 B.n389 585
R290 B.n388 B.n387 585
R291 B.n386 B.n385 585
R292 B.n384 B.n383 585
R293 B.n382 B.n381 585
R294 B.n380 B.n379 585
R295 B.n378 B.n377 585
R296 B.n376 B.n375 585
R297 B.n374 B.n373 585
R298 B.n372 B.n371 585
R299 B.n370 B.n369 585
R300 B.n368 B.n367 585
R301 B.n365 B.n364 585
R302 B.n363 B.n362 585
R303 B.n361 B.n360 585
R304 B.n359 B.n358 585
R305 B.n357 B.n356 585
R306 B.n355 B.n354 585
R307 B.n353 B.n352 585
R308 B.n351 B.n350 585
R309 B.n349 B.n348 585
R310 B.n347 B.n346 585
R311 B.n345 B.n344 585
R312 B.n343 B.n342 585
R313 B.n341 B.n340 585
R314 B.n339 B.n338 585
R315 B.n337 B.n336 585
R316 B.n335 B.n334 585
R317 B.n333 B.n332 585
R318 B.n331 B.n330 585
R319 B.n329 B.n328 585
R320 B.n327 B.n326 585
R321 B.n325 B.n324 585
R322 B.n323 B.n322 585
R323 B.n321 B.n320 585
R324 B.n430 B.n285 585
R325 B.n285 B.n284 585
R326 B.n432 B.n431 585
R327 B.n433 B.n432 585
R328 B.n279 B.n278 585
R329 B.n280 B.n279 585
R330 B.n441 B.n440 585
R331 B.n440 B.n439 585
R332 B.n442 B.n277 585
R333 B.n277 B.n276 585
R334 B.n444 B.n443 585
R335 B.n445 B.n444 585
R336 B.n271 B.n270 585
R337 B.n272 B.n271 585
R338 B.n454 B.n453 585
R339 B.n453 B.n452 585
R340 B.n455 B.n269 585
R341 B.n451 B.n269 585
R342 B.n457 B.n456 585
R343 B.n458 B.n457 585
R344 B.n264 B.n263 585
R345 B.n265 B.n264 585
R346 B.n466 B.n465 585
R347 B.n465 B.n464 585
R348 B.n467 B.n262 585
R349 B.n262 B.n261 585
R350 B.n469 B.n468 585
R351 B.n470 B.n469 585
R352 B.n256 B.n255 585
R353 B.n257 B.n256 585
R354 B.n478 B.n477 585
R355 B.n477 B.n476 585
R356 B.n479 B.n254 585
R357 B.n254 B.n253 585
R358 B.n481 B.n480 585
R359 B.n482 B.n481 585
R360 B.n248 B.n247 585
R361 B.n249 B.n248 585
R362 B.n490 B.n489 585
R363 B.n489 B.n488 585
R364 B.n491 B.n246 585
R365 B.n246 B.n245 585
R366 B.n493 B.n492 585
R367 B.n494 B.n493 585
R368 B.n240 B.n239 585
R369 B.n241 B.n240 585
R370 B.n502 B.n501 585
R371 B.n501 B.n500 585
R372 B.n503 B.n238 585
R373 B.n238 B.n237 585
R374 B.n505 B.n504 585
R375 B.n506 B.n505 585
R376 B.n232 B.n231 585
R377 B.n233 B.n232 585
R378 B.n514 B.n513 585
R379 B.n513 B.n512 585
R380 B.n515 B.n230 585
R381 B.n230 B.n229 585
R382 B.n517 B.n516 585
R383 B.n518 B.n517 585
R384 B.n224 B.n223 585
R385 B.n225 B.n224 585
R386 B.n527 B.n526 585
R387 B.n526 B.n525 585
R388 B.n528 B.n222 585
R389 B.n524 B.n222 585
R390 B.n530 B.n529 585
R391 B.n531 B.n530 585
R392 B.n217 B.n216 585
R393 B.n218 B.n217 585
R394 B.n540 B.n539 585
R395 B.n539 B.n538 585
R396 B.n541 B.n215 585
R397 B.n215 B.n214 585
R398 B.n543 B.n542 585
R399 B.n544 B.n543 585
R400 B.n2 B.n0 585
R401 B.n4 B.n2 585
R402 B.n3 B.n1 585
R403 B.n679 B.n3 585
R404 B.n677 B.n676 585
R405 B.n678 B.n677 585
R406 B.n675 B.n9 585
R407 B.n9 B.n8 585
R408 B.n674 B.n673 585
R409 B.n673 B.n672 585
R410 B.n11 B.n10 585
R411 B.n671 B.n11 585
R412 B.n669 B.n668 585
R413 B.n670 B.n669 585
R414 B.n667 B.n15 585
R415 B.n18 B.n15 585
R416 B.n666 B.n665 585
R417 B.n665 B.n664 585
R418 B.n17 B.n16 585
R419 B.n663 B.n17 585
R420 B.n661 B.n660 585
R421 B.n662 B.n661 585
R422 B.n659 B.n23 585
R423 B.n23 B.n22 585
R424 B.n658 B.n657 585
R425 B.n657 B.n656 585
R426 B.n25 B.n24 585
R427 B.n655 B.n25 585
R428 B.n653 B.n652 585
R429 B.n654 B.n653 585
R430 B.n651 B.n30 585
R431 B.n30 B.n29 585
R432 B.n650 B.n649 585
R433 B.n649 B.n648 585
R434 B.n32 B.n31 585
R435 B.n647 B.n32 585
R436 B.n645 B.n644 585
R437 B.n646 B.n645 585
R438 B.n643 B.n37 585
R439 B.n37 B.n36 585
R440 B.n642 B.n641 585
R441 B.n641 B.n640 585
R442 B.n39 B.n38 585
R443 B.n639 B.n39 585
R444 B.n637 B.n636 585
R445 B.n638 B.n637 585
R446 B.n635 B.n44 585
R447 B.n44 B.n43 585
R448 B.n634 B.n633 585
R449 B.n633 B.n632 585
R450 B.n46 B.n45 585
R451 B.n631 B.n46 585
R452 B.n629 B.n628 585
R453 B.n630 B.n629 585
R454 B.n627 B.n51 585
R455 B.n51 B.n50 585
R456 B.n626 B.n625 585
R457 B.n625 B.n624 585
R458 B.n53 B.n52 585
R459 B.n623 B.n53 585
R460 B.n621 B.n620 585
R461 B.n622 B.n621 585
R462 B.n619 B.n57 585
R463 B.n60 B.n57 585
R464 B.n618 B.n617 585
R465 B.n617 B.n616 585
R466 B.n59 B.n58 585
R467 B.n615 B.n59 585
R468 B.n613 B.n612 585
R469 B.n614 B.n613 585
R470 B.n611 B.n65 585
R471 B.n65 B.n64 585
R472 B.n610 B.n609 585
R473 B.n609 B.n608 585
R474 B.n67 B.n66 585
R475 B.n607 B.n67 585
R476 B.n605 B.n604 585
R477 B.n606 B.n605 585
R478 B.n603 B.n72 585
R479 B.n72 B.n71 585
R480 B.n682 B.n681 585
R481 B.n681 B.n680 585
R482 B.n428 B.n285 482.89
R483 B.n601 B.n72 482.89
R484 B.n320 B.n283 482.89
R485 B.n598 B.n102 482.89
R486 B.n599 B.n100 256.663
R487 B.n599 B.n99 256.663
R488 B.n599 B.n98 256.663
R489 B.n599 B.n97 256.663
R490 B.n599 B.n96 256.663
R491 B.n599 B.n95 256.663
R492 B.n599 B.n94 256.663
R493 B.n599 B.n93 256.663
R494 B.n599 B.n92 256.663
R495 B.n599 B.n91 256.663
R496 B.n599 B.n90 256.663
R497 B.n599 B.n89 256.663
R498 B.n599 B.n88 256.663
R499 B.n599 B.n87 256.663
R500 B.n599 B.n86 256.663
R501 B.n599 B.n85 256.663
R502 B.n599 B.n84 256.663
R503 B.n599 B.n83 256.663
R504 B.n599 B.n82 256.663
R505 B.n599 B.n81 256.663
R506 B.n599 B.n80 256.663
R507 B.n599 B.n79 256.663
R508 B.n599 B.n78 256.663
R509 B.n599 B.n77 256.663
R510 B.n599 B.n76 256.663
R511 B.n599 B.n75 256.663
R512 B.n600 B.n599 256.663
R513 B.n427 B.n426 256.663
R514 B.n426 B.n288 256.663
R515 B.n426 B.n289 256.663
R516 B.n426 B.n290 256.663
R517 B.n426 B.n291 256.663
R518 B.n426 B.n292 256.663
R519 B.n426 B.n293 256.663
R520 B.n426 B.n294 256.663
R521 B.n426 B.n295 256.663
R522 B.n426 B.n296 256.663
R523 B.n426 B.n297 256.663
R524 B.n426 B.n298 256.663
R525 B.n426 B.n299 256.663
R526 B.n426 B.n300 256.663
R527 B.n426 B.n301 256.663
R528 B.n426 B.n302 256.663
R529 B.n426 B.n303 256.663
R530 B.n426 B.n304 256.663
R531 B.n426 B.n305 256.663
R532 B.n426 B.n306 256.663
R533 B.n426 B.n307 256.663
R534 B.n426 B.n308 256.663
R535 B.n426 B.n309 256.663
R536 B.n426 B.n310 256.663
R537 B.n426 B.n311 256.663
R538 B.n426 B.n312 256.663
R539 B.n426 B.n313 256.663
R540 B.n318 B.t4 250.54
R541 B.n315 B.t8 250.54
R542 B.n106 B.t11 250.54
R543 B.n103 B.t15 250.54
R544 B.n432 B.n285 163.367
R545 B.n432 B.n279 163.367
R546 B.n440 B.n279 163.367
R547 B.n440 B.n277 163.367
R548 B.n444 B.n277 163.367
R549 B.n444 B.n271 163.367
R550 B.n453 B.n271 163.367
R551 B.n453 B.n269 163.367
R552 B.n457 B.n269 163.367
R553 B.n457 B.n264 163.367
R554 B.n465 B.n264 163.367
R555 B.n465 B.n262 163.367
R556 B.n469 B.n262 163.367
R557 B.n469 B.n256 163.367
R558 B.n477 B.n256 163.367
R559 B.n477 B.n254 163.367
R560 B.n481 B.n254 163.367
R561 B.n481 B.n248 163.367
R562 B.n489 B.n248 163.367
R563 B.n489 B.n246 163.367
R564 B.n493 B.n246 163.367
R565 B.n493 B.n240 163.367
R566 B.n501 B.n240 163.367
R567 B.n501 B.n238 163.367
R568 B.n505 B.n238 163.367
R569 B.n505 B.n232 163.367
R570 B.n513 B.n232 163.367
R571 B.n513 B.n230 163.367
R572 B.n517 B.n230 163.367
R573 B.n517 B.n224 163.367
R574 B.n526 B.n224 163.367
R575 B.n526 B.n222 163.367
R576 B.n530 B.n222 163.367
R577 B.n530 B.n217 163.367
R578 B.n539 B.n217 163.367
R579 B.n539 B.n215 163.367
R580 B.n543 B.n215 163.367
R581 B.n543 B.n2 163.367
R582 B.n681 B.n2 163.367
R583 B.n681 B.n3 163.367
R584 B.n677 B.n3 163.367
R585 B.n677 B.n9 163.367
R586 B.n673 B.n9 163.367
R587 B.n673 B.n11 163.367
R588 B.n669 B.n11 163.367
R589 B.n669 B.n15 163.367
R590 B.n665 B.n15 163.367
R591 B.n665 B.n17 163.367
R592 B.n661 B.n17 163.367
R593 B.n661 B.n23 163.367
R594 B.n657 B.n23 163.367
R595 B.n657 B.n25 163.367
R596 B.n653 B.n25 163.367
R597 B.n653 B.n30 163.367
R598 B.n649 B.n30 163.367
R599 B.n649 B.n32 163.367
R600 B.n645 B.n32 163.367
R601 B.n645 B.n37 163.367
R602 B.n641 B.n37 163.367
R603 B.n641 B.n39 163.367
R604 B.n637 B.n39 163.367
R605 B.n637 B.n44 163.367
R606 B.n633 B.n44 163.367
R607 B.n633 B.n46 163.367
R608 B.n629 B.n46 163.367
R609 B.n629 B.n51 163.367
R610 B.n625 B.n51 163.367
R611 B.n625 B.n53 163.367
R612 B.n621 B.n53 163.367
R613 B.n621 B.n57 163.367
R614 B.n617 B.n57 163.367
R615 B.n617 B.n59 163.367
R616 B.n613 B.n59 163.367
R617 B.n613 B.n65 163.367
R618 B.n609 B.n65 163.367
R619 B.n609 B.n67 163.367
R620 B.n605 B.n67 163.367
R621 B.n605 B.n72 163.367
R622 B.n425 B.n287 163.367
R623 B.n425 B.n314 163.367
R624 B.n421 B.n420 163.367
R625 B.n417 B.n416 163.367
R626 B.n413 B.n412 163.367
R627 B.n409 B.n408 163.367
R628 B.n405 B.n404 163.367
R629 B.n401 B.n400 163.367
R630 B.n397 B.n396 163.367
R631 B.n393 B.n392 163.367
R632 B.n389 B.n388 163.367
R633 B.n385 B.n384 163.367
R634 B.n381 B.n380 163.367
R635 B.n377 B.n376 163.367
R636 B.n373 B.n372 163.367
R637 B.n369 B.n368 163.367
R638 B.n364 B.n363 163.367
R639 B.n360 B.n359 163.367
R640 B.n356 B.n355 163.367
R641 B.n352 B.n351 163.367
R642 B.n348 B.n347 163.367
R643 B.n344 B.n343 163.367
R644 B.n340 B.n339 163.367
R645 B.n336 B.n335 163.367
R646 B.n332 B.n331 163.367
R647 B.n328 B.n327 163.367
R648 B.n324 B.n323 163.367
R649 B.n434 B.n283 163.367
R650 B.n434 B.n281 163.367
R651 B.n438 B.n281 163.367
R652 B.n438 B.n275 163.367
R653 B.n446 B.n275 163.367
R654 B.n446 B.n273 163.367
R655 B.n450 B.n273 163.367
R656 B.n450 B.n268 163.367
R657 B.n459 B.n268 163.367
R658 B.n459 B.n266 163.367
R659 B.n463 B.n266 163.367
R660 B.n463 B.n260 163.367
R661 B.n471 B.n260 163.367
R662 B.n471 B.n258 163.367
R663 B.n475 B.n258 163.367
R664 B.n475 B.n252 163.367
R665 B.n483 B.n252 163.367
R666 B.n483 B.n250 163.367
R667 B.n487 B.n250 163.367
R668 B.n487 B.n244 163.367
R669 B.n495 B.n244 163.367
R670 B.n495 B.n242 163.367
R671 B.n499 B.n242 163.367
R672 B.n499 B.n236 163.367
R673 B.n507 B.n236 163.367
R674 B.n507 B.n234 163.367
R675 B.n511 B.n234 163.367
R676 B.n511 B.n228 163.367
R677 B.n519 B.n228 163.367
R678 B.n519 B.n226 163.367
R679 B.n523 B.n226 163.367
R680 B.n523 B.n221 163.367
R681 B.n532 B.n221 163.367
R682 B.n532 B.n219 163.367
R683 B.n537 B.n219 163.367
R684 B.n537 B.n213 163.367
R685 B.n545 B.n213 163.367
R686 B.n546 B.n545 163.367
R687 B.n546 B.n5 163.367
R688 B.n6 B.n5 163.367
R689 B.n7 B.n6 163.367
R690 B.n551 B.n7 163.367
R691 B.n551 B.n12 163.367
R692 B.n13 B.n12 163.367
R693 B.n14 B.n13 163.367
R694 B.n556 B.n14 163.367
R695 B.n556 B.n19 163.367
R696 B.n20 B.n19 163.367
R697 B.n21 B.n20 163.367
R698 B.n561 B.n21 163.367
R699 B.n561 B.n26 163.367
R700 B.n27 B.n26 163.367
R701 B.n28 B.n27 163.367
R702 B.n566 B.n28 163.367
R703 B.n566 B.n33 163.367
R704 B.n34 B.n33 163.367
R705 B.n35 B.n34 163.367
R706 B.n571 B.n35 163.367
R707 B.n571 B.n40 163.367
R708 B.n41 B.n40 163.367
R709 B.n42 B.n41 163.367
R710 B.n576 B.n42 163.367
R711 B.n576 B.n47 163.367
R712 B.n48 B.n47 163.367
R713 B.n49 B.n48 163.367
R714 B.n581 B.n49 163.367
R715 B.n581 B.n54 163.367
R716 B.n55 B.n54 163.367
R717 B.n56 B.n55 163.367
R718 B.n586 B.n56 163.367
R719 B.n586 B.n61 163.367
R720 B.n62 B.n61 163.367
R721 B.n63 B.n62 163.367
R722 B.n591 B.n63 163.367
R723 B.n591 B.n68 163.367
R724 B.n69 B.n68 163.367
R725 B.n70 B.n69 163.367
R726 B.n102 B.n70 163.367
R727 B.n108 B.n74 163.367
R728 B.n112 B.n111 163.367
R729 B.n116 B.n115 163.367
R730 B.n120 B.n119 163.367
R731 B.n124 B.n123 163.367
R732 B.n128 B.n127 163.367
R733 B.n132 B.n131 163.367
R734 B.n136 B.n135 163.367
R735 B.n140 B.n139 163.367
R736 B.n144 B.n143 163.367
R737 B.n148 B.n147 163.367
R738 B.n153 B.n152 163.367
R739 B.n157 B.n156 163.367
R740 B.n161 B.n160 163.367
R741 B.n165 B.n164 163.367
R742 B.n169 B.n168 163.367
R743 B.n173 B.n172 163.367
R744 B.n177 B.n176 163.367
R745 B.n181 B.n180 163.367
R746 B.n185 B.n184 163.367
R747 B.n189 B.n188 163.367
R748 B.n193 B.n192 163.367
R749 B.n197 B.n196 163.367
R750 B.n201 B.n200 163.367
R751 B.n205 B.n204 163.367
R752 B.n209 B.n208 163.367
R753 B.n598 B.n101 163.367
R754 B.n318 B.t7 139.189
R755 B.n103 B.t16 139.189
R756 B.n315 B.t10 139.183
R757 B.n106 B.t13 139.183
R758 B.n426 B.n284 131.572
R759 B.n599 B.n71 131.572
R760 B.n428 B.n427 71.676
R761 B.n314 B.n288 71.676
R762 B.n420 B.n289 71.676
R763 B.n416 B.n290 71.676
R764 B.n412 B.n291 71.676
R765 B.n408 B.n292 71.676
R766 B.n404 B.n293 71.676
R767 B.n400 B.n294 71.676
R768 B.n396 B.n295 71.676
R769 B.n392 B.n296 71.676
R770 B.n388 B.n297 71.676
R771 B.n384 B.n298 71.676
R772 B.n380 B.n299 71.676
R773 B.n376 B.n300 71.676
R774 B.n372 B.n301 71.676
R775 B.n368 B.n302 71.676
R776 B.n363 B.n303 71.676
R777 B.n359 B.n304 71.676
R778 B.n355 B.n305 71.676
R779 B.n351 B.n306 71.676
R780 B.n347 B.n307 71.676
R781 B.n343 B.n308 71.676
R782 B.n339 B.n309 71.676
R783 B.n335 B.n310 71.676
R784 B.n331 B.n311 71.676
R785 B.n327 B.n312 71.676
R786 B.n323 B.n313 71.676
R787 B.n601 B.n600 71.676
R788 B.n108 B.n75 71.676
R789 B.n112 B.n76 71.676
R790 B.n116 B.n77 71.676
R791 B.n120 B.n78 71.676
R792 B.n124 B.n79 71.676
R793 B.n128 B.n80 71.676
R794 B.n132 B.n81 71.676
R795 B.n136 B.n82 71.676
R796 B.n140 B.n83 71.676
R797 B.n144 B.n84 71.676
R798 B.n148 B.n85 71.676
R799 B.n153 B.n86 71.676
R800 B.n157 B.n87 71.676
R801 B.n161 B.n88 71.676
R802 B.n165 B.n89 71.676
R803 B.n169 B.n90 71.676
R804 B.n173 B.n91 71.676
R805 B.n177 B.n92 71.676
R806 B.n181 B.n93 71.676
R807 B.n185 B.n94 71.676
R808 B.n189 B.n95 71.676
R809 B.n193 B.n96 71.676
R810 B.n197 B.n97 71.676
R811 B.n201 B.n98 71.676
R812 B.n205 B.n99 71.676
R813 B.n209 B.n100 71.676
R814 B.n101 B.n100 71.676
R815 B.n208 B.n99 71.676
R816 B.n204 B.n98 71.676
R817 B.n200 B.n97 71.676
R818 B.n196 B.n96 71.676
R819 B.n192 B.n95 71.676
R820 B.n188 B.n94 71.676
R821 B.n184 B.n93 71.676
R822 B.n180 B.n92 71.676
R823 B.n176 B.n91 71.676
R824 B.n172 B.n90 71.676
R825 B.n168 B.n89 71.676
R826 B.n164 B.n88 71.676
R827 B.n160 B.n87 71.676
R828 B.n156 B.n86 71.676
R829 B.n152 B.n85 71.676
R830 B.n147 B.n84 71.676
R831 B.n143 B.n83 71.676
R832 B.n139 B.n82 71.676
R833 B.n135 B.n81 71.676
R834 B.n131 B.n80 71.676
R835 B.n127 B.n79 71.676
R836 B.n123 B.n78 71.676
R837 B.n119 B.n77 71.676
R838 B.n115 B.n76 71.676
R839 B.n111 B.n75 71.676
R840 B.n600 B.n74 71.676
R841 B.n427 B.n287 71.676
R842 B.n421 B.n288 71.676
R843 B.n417 B.n289 71.676
R844 B.n413 B.n290 71.676
R845 B.n409 B.n291 71.676
R846 B.n405 B.n292 71.676
R847 B.n401 B.n293 71.676
R848 B.n397 B.n294 71.676
R849 B.n393 B.n295 71.676
R850 B.n389 B.n296 71.676
R851 B.n385 B.n297 71.676
R852 B.n381 B.n298 71.676
R853 B.n377 B.n299 71.676
R854 B.n373 B.n300 71.676
R855 B.n369 B.n301 71.676
R856 B.n364 B.n302 71.676
R857 B.n360 B.n303 71.676
R858 B.n356 B.n304 71.676
R859 B.n352 B.n305 71.676
R860 B.n348 B.n306 71.676
R861 B.n344 B.n307 71.676
R862 B.n340 B.n308 71.676
R863 B.n336 B.n309 71.676
R864 B.n332 B.n310 71.676
R865 B.n328 B.n311 71.676
R866 B.n324 B.n312 71.676
R867 B.n320 B.n313 71.676
R868 B.n319 B.t6 71.1154
R869 B.n104 B.t17 71.1154
R870 B.n316 B.t9 71.1096
R871 B.n107 B.t14 71.1096
R872 B.n433 B.n284 69.3561
R873 B.n433 B.n280 69.3561
R874 B.n439 B.n280 69.3561
R875 B.n439 B.n276 69.3561
R876 B.n445 B.n276 69.3561
R877 B.n445 B.n272 69.3561
R878 B.n452 B.n272 69.3561
R879 B.n452 B.n451 69.3561
R880 B.n458 B.n265 69.3561
R881 B.n464 B.n265 69.3561
R882 B.n464 B.n261 69.3561
R883 B.n470 B.n261 69.3561
R884 B.n470 B.n257 69.3561
R885 B.n476 B.n257 69.3561
R886 B.n476 B.n253 69.3561
R887 B.n482 B.n253 69.3561
R888 B.n482 B.n249 69.3561
R889 B.n488 B.n249 69.3561
R890 B.n488 B.n245 69.3561
R891 B.n494 B.n245 69.3561
R892 B.n500 B.n241 69.3561
R893 B.n500 B.n237 69.3561
R894 B.n506 B.n237 69.3561
R895 B.n506 B.n233 69.3561
R896 B.n512 B.n233 69.3561
R897 B.n512 B.n229 69.3561
R898 B.n518 B.n229 69.3561
R899 B.n518 B.n225 69.3561
R900 B.n525 B.n225 69.3561
R901 B.n525 B.n524 69.3561
R902 B.n531 B.n218 69.3561
R903 B.n538 B.n218 69.3561
R904 B.n538 B.n214 69.3561
R905 B.n544 B.n214 69.3561
R906 B.n544 B.n4 69.3561
R907 B.n680 B.n4 69.3561
R908 B.n680 B.n679 69.3561
R909 B.n679 B.n678 69.3561
R910 B.n678 B.n8 69.3561
R911 B.n672 B.n8 69.3561
R912 B.n672 B.n671 69.3561
R913 B.n671 B.n670 69.3561
R914 B.n664 B.n18 69.3561
R915 B.n664 B.n663 69.3561
R916 B.n663 B.n662 69.3561
R917 B.n662 B.n22 69.3561
R918 B.n656 B.n22 69.3561
R919 B.n656 B.n655 69.3561
R920 B.n655 B.n654 69.3561
R921 B.n654 B.n29 69.3561
R922 B.n648 B.n29 69.3561
R923 B.n648 B.n647 69.3561
R924 B.n646 B.n36 69.3561
R925 B.n640 B.n36 69.3561
R926 B.n640 B.n639 69.3561
R927 B.n639 B.n638 69.3561
R928 B.n638 B.n43 69.3561
R929 B.n632 B.n43 69.3561
R930 B.n632 B.n631 69.3561
R931 B.n631 B.n630 69.3561
R932 B.n630 B.n50 69.3561
R933 B.n624 B.n50 69.3561
R934 B.n624 B.n623 69.3561
R935 B.n623 B.n622 69.3561
R936 B.n616 B.n60 69.3561
R937 B.n616 B.n615 69.3561
R938 B.n615 B.n614 69.3561
R939 B.n614 B.n64 69.3561
R940 B.n608 B.n64 69.3561
R941 B.n608 B.n607 69.3561
R942 B.n607 B.n606 69.3561
R943 B.n606 B.n71 69.3561
R944 B.n319 B.n318 68.0732
R945 B.n316 B.n315 68.0732
R946 B.n107 B.n106 68.0732
R947 B.n104 B.n103 68.0732
R948 B.n494 B.t3 63.2365
R949 B.t0 B.n646 63.2365
R950 B.n366 B.n319 59.5399
R951 B.n317 B.n316 59.5399
R952 B.n150 B.n107 59.5399
R953 B.n105 B.n104 59.5399
R954 B.n531 B.t1 53.0371
R955 B.n670 B.t2 53.0371
R956 B.n458 B.t5 42.8378
R957 B.n622 B.t12 42.8378
R958 B.n603 B.n602 31.3761
R959 B.n597 B.n596 31.3761
R960 B.n321 B.n282 31.3761
R961 B.n430 B.n429 31.3761
R962 B.n451 B.t5 26.5188
R963 B.n60 B.t12 26.5188
R964 B B.n682 18.0485
R965 B.n524 B.t1 16.3195
R966 B.n18 B.t2 16.3195
R967 B.n602 B.n73 10.6151
R968 B.n109 B.n73 10.6151
R969 B.n110 B.n109 10.6151
R970 B.n113 B.n110 10.6151
R971 B.n114 B.n113 10.6151
R972 B.n117 B.n114 10.6151
R973 B.n118 B.n117 10.6151
R974 B.n121 B.n118 10.6151
R975 B.n122 B.n121 10.6151
R976 B.n125 B.n122 10.6151
R977 B.n126 B.n125 10.6151
R978 B.n129 B.n126 10.6151
R979 B.n130 B.n129 10.6151
R980 B.n133 B.n130 10.6151
R981 B.n134 B.n133 10.6151
R982 B.n137 B.n134 10.6151
R983 B.n138 B.n137 10.6151
R984 B.n141 B.n138 10.6151
R985 B.n142 B.n141 10.6151
R986 B.n145 B.n142 10.6151
R987 B.n146 B.n145 10.6151
R988 B.n149 B.n146 10.6151
R989 B.n154 B.n151 10.6151
R990 B.n155 B.n154 10.6151
R991 B.n158 B.n155 10.6151
R992 B.n159 B.n158 10.6151
R993 B.n162 B.n159 10.6151
R994 B.n163 B.n162 10.6151
R995 B.n166 B.n163 10.6151
R996 B.n167 B.n166 10.6151
R997 B.n171 B.n170 10.6151
R998 B.n174 B.n171 10.6151
R999 B.n175 B.n174 10.6151
R1000 B.n178 B.n175 10.6151
R1001 B.n179 B.n178 10.6151
R1002 B.n182 B.n179 10.6151
R1003 B.n183 B.n182 10.6151
R1004 B.n186 B.n183 10.6151
R1005 B.n187 B.n186 10.6151
R1006 B.n190 B.n187 10.6151
R1007 B.n191 B.n190 10.6151
R1008 B.n194 B.n191 10.6151
R1009 B.n195 B.n194 10.6151
R1010 B.n198 B.n195 10.6151
R1011 B.n199 B.n198 10.6151
R1012 B.n202 B.n199 10.6151
R1013 B.n203 B.n202 10.6151
R1014 B.n206 B.n203 10.6151
R1015 B.n207 B.n206 10.6151
R1016 B.n210 B.n207 10.6151
R1017 B.n211 B.n210 10.6151
R1018 B.n597 B.n211 10.6151
R1019 B.n435 B.n282 10.6151
R1020 B.n436 B.n435 10.6151
R1021 B.n437 B.n436 10.6151
R1022 B.n437 B.n274 10.6151
R1023 B.n447 B.n274 10.6151
R1024 B.n448 B.n447 10.6151
R1025 B.n449 B.n448 10.6151
R1026 B.n449 B.n267 10.6151
R1027 B.n460 B.n267 10.6151
R1028 B.n461 B.n460 10.6151
R1029 B.n462 B.n461 10.6151
R1030 B.n462 B.n259 10.6151
R1031 B.n472 B.n259 10.6151
R1032 B.n473 B.n472 10.6151
R1033 B.n474 B.n473 10.6151
R1034 B.n474 B.n251 10.6151
R1035 B.n484 B.n251 10.6151
R1036 B.n485 B.n484 10.6151
R1037 B.n486 B.n485 10.6151
R1038 B.n486 B.n243 10.6151
R1039 B.n496 B.n243 10.6151
R1040 B.n497 B.n496 10.6151
R1041 B.n498 B.n497 10.6151
R1042 B.n498 B.n235 10.6151
R1043 B.n508 B.n235 10.6151
R1044 B.n509 B.n508 10.6151
R1045 B.n510 B.n509 10.6151
R1046 B.n510 B.n227 10.6151
R1047 B.n520 B.n227 10.6151
R1048 B.n521 B.n520 10.6151
R1049 B.n522 B.n521 10.6151
R1050 B.n522 B.n220 10.6151
R1051 B.n533 B.n220 10.6151
R1052 B.n534 B.n533 10.6151
R1053 B.n536 B.n534 10.6151
R1054 B.n536 B.n535 10.6151
R1055 B.n535 B.n212 10.6151
R1056 B.n547 B.n212 10.6151
R1057 B.n548 B.n547 10.6151
R1058 B.n549 B.n548 10.6151
R1059 B.n550 B.n549 10.6151
R1060 B.n552 B.n550 10.6151
R1061 B.n553 B.n552 10.6151
R1062 B.n554 B.n553 10.6151
R1063 B.n555 B.n554 10.6151
R1064 B.n557 B.n555 10.6151
R1065 B.n558 B.n557 10.6151
R1066 B.n559 B.n558 10.6151
R1067 B.n560 B.n559 10.6151
R1068 B.n562 B.n560 10.6151
R1069 B.n563 B.n562 10.6151
R1070 B.n564 B.n563 10.6151
R1071 B.n565 B.n564 10.6151
R1072 B.n567 B.n565 10.6151
R1073 B.n568 B.n567 10.6151
R1074 B.n569 B.n568 10.6151
R1075 B.n570 B.n569 10.6151
R1076 B.n572 B.n570 10.6151
R1077 B.n573 B.n572 10.6151
R1078 B.n574 B.n573 10.6151
R1079 B.n575 B.n574 10.6151
R1080 B.n577 B.n575 10.6151
R1081 B.n578 B.n577 10.6151
R1082 B.n579 B.n578 10.6151
R1083 B.n580 B.n579 10.6151
R1084 B.n582 B.n580 10.6151
R1085 B.n583 B.n582 10.6151
R1086 B.n584 B.n583 10.6151
R1087 B.n585 B.n584 10.6151
R1088 B.n587 B.n585 10.6151
R1089 B.n588 B.n587 10.6151
R1090 B.n589 B.n588 10.6151
R1091 B.n590 B.n589 10.6151
R1092 B.n592 B.n590 10.6151
R1093 B.n593 B.n592 10.6151
R1094 B.n594 B.n593 10.6151
R1095 B.n595 B.n594 10.6151
R1096 B.n596 B.n595 10.6151
R1097 B.n429 B.n286 10.6151
R1098 B.n424 B.n286 10.6151
R1099 B.n424 B.n423 10.6151
R1100 B.n423 B.n422 10.6151
R1101 B.n422 B.n419 10.6151
R1102 B.n419 B.n418 10.6151
R1103 B.n418 B.n415 10.6151
R1104 B.n415 B.n414 10.6151
R1105 B.n414 B.n411 10.6151
R1106 B.n411 B.n410 10.6151
R1107 B.n410 B.n407 10.6151
R1108 B.n407 B.n406 10.6151
R1109 B.n406 B.n403 10.6151
R1110 B.n403 B.n402 10.6151
R1111 B.n402 B.n399 10.6151
R1112 B.n399 B.n398 10.6151
R1113 B.n398 B.n395 10.6151
R1114 B.n395 B.n394 10.6151
R1115 B.n394 B.n391 10.6151
R1116 B.n391 B.n390 10.6151
R1117 B.n390 B.n387 10.6151
R1118 B.n387 B.n386 10.6151
R1119 B.n383 B.n382 10.6151
R1120 B.n382 B.n379 10.6151
R1121 B.n379 B.n378 10.6151
R1122 B.n378 B.n375 10.6151
R1123 B.n375 B.n374 10.6151
R1124 B.n374 B.n371 10.6151
R1125 B.n371 B.n370 10.6151
R1126 B.n370 B.n367 10.6151
R1127 B.n365 B.n362 10.6151
R1128 B.n362 B.n361 10.6151
R1129 B.n361 B.n358 10.6151
R1130 B.n358 B.n357 10.6151
R1131 B.n357 B.n354 10.6151
R1132 B.n354 B.n353 10.6151
R1133 B.n353 B.n350 10.6151
R1134 B.n350 B.n349 10.6151
R1135 B.n349 B.n346 10.6151
R1136 B.n346 B.n345 10.6151
R1137 B.n345 B.n342 10.6151
R1138 B.n342 B.n341 10.6151
R1139 B.n341 B.n338 10.6151
R1140 B.n338 B.n337 10.6151
R1141 B.n337 B.n334 10.6151
R1142 B.n334 B.n333 10.6151
R1143 B.n333 B.n330 10.6151
R1144 B.n330 B.n329 10.6151
R1145 B.n329 B.n326 10.6151
R1146 B.n326 B.n325 10.6151
R1147 B.n325 B.n322 10.6151
R1148 B.n322 B.n321 10.6151
R1149 B.n431 B.n430 10.6151
R1150 B.n431 B.n278 10.6151
R1151 B.n441 B.n278 10.6151
R1152 B.n442 B.n441 10.6151
R1153 B.n443 B.n442 10.6151
R1154 B.n443 B.n270 10.6151
R1155 B.n454 B.n270 10.6151
R1156 B.n455 B.n454 10.6151
R1157 B.n456 B.n455 10.6151
R1158 B.n456 B.n263 10.6151
R1159 B.n466 B.n263 10.6151
R1160 B.n467 B.n466 10.6151
R1161 B.n468 B.n467 10.6151
R1162 B.n468 B.n255 10.6151
R1163 B.n478 B.n255 10.6151
R1164 B.n479 B.n478 10.6151
R1165 B.n480 B.n479 10.6151
R1166 B.n480 B.n247 10.6151
R1167 B.n490 B.n247 10.6151
R1168 B.n491 B.n490 10.6151
R1169 B.n492 B.n491 10.6151
R1170 B.n492 B.n239 10.6151
R1171 B.n502 B.n239 10.6151
R1172 B.n503 B.n502 10.6151
R1173 B.n504 B.n503 10.6151
R1174 B.n504 B.n231 10.6151
R1175 B.n514 B.n231 10.6151
R1176 B.n515 B.n514 10.6151
R1177 B.n516 B.n515 10.6151
R1178 B.n516 B.n223 10.6151
R1179 B.n527 B.n223 10.6151
R1180 B.n528 B.n527 10.6151
R1181 B.n529 B.n528 10.6151
R1182 B.n529 B.n216 10.6151
R1183 B.n540 B.n216 10.6151
R1184 B.n541 B.n540 10.6151
R1185 B.n542 B.n541 10.6151
R1186 B.n542 B.n0 10.6151
R1187 B.n676 B.n1 10.6151
R1188 B.n676 B.n675 10.6151
R1189 B.n675 B.n674 10.6151
R1190 B.n674 B.n10 10.6151
R1191 B.n668 B.n10 10.6151
R1192 B.n668 B.n667 10.6151
R1193 B.n667 B.n666 10.6151
R1194 B.n666 B.n16 10.6151
R1195 B.n660 B.n16 10.6151
R1196 B.n660 B.n659 10.6151
R1197 B.n659 B.n658 10.6151
R1198 B.n658 B.n24 10.6151
R1199 B.n652 B.n24 10.6151
R1200 B.n652 B.n651 10.6151
R1201 B.n651 B.n650 10.6151
R1202 B.n650 B.n31 10.6151
R1203 B.n644 B.n31 10.6151
R1204 B.n644 B.n643 10.6151
R1205 B.n643 B.n642 10.6151
R1206 B.n642 B.n38 10.6151
R1207 B.n636 B.n38 10.6151
R1208 B.n636 B.n635 10.6151
R1209 B.n635 B.n634 10.6151
R1210 B.n634 B.n45 10.6151
R1211 B.n628 B.n45 10.6151
R1212 B.n628 B.n627 10.6151
R1213 B.n627 B.n626 10.6151
R1214 B.n626 B.n52 10.6151
R1215 B.n620 B.n52 10.6151
R1216 B.n620 B.n619 10.6151
R1217 B.n619 B.n618 10.6151
R1218 B.n618 B.n58 10.6151
R1219 B.n612 B.n58 10.6151
R1220 B.n612 B.n611 10.6151
R1221 B.n611 B.n610 10.6151
R1222 B.n610 B.n66 10.6151
R1223 B.n604 B.n66 10.6151
R1224 B.n604 B.n603 10.6151
R1225 B.n151 B.n150 6.5566
R1226 B.n167 B.n105 6.5566
R1227 B.n383 B.n317 6.5566
R1228 B.n367 B.n366 6.5566
R1229 B.t3 B.n241 6.12011
R1230 B.n647 B.t0 6.12011
R1231 B.n150 B.n149 4.05904
R1232 B.n170 B.n105 4.05904
R1233 B.n386 B.n317 4.05904
R1234 B.n366 B.n365 4.05904
R1235 B.n682 B.n0 2.81026
R1236 B.n682 B.n1 2.81026
R1237 VN.n0 VN.t2 76.3399
R1238 VN.n1 VN.t1 76.3399
R1239 VN.n0 VN.t0 75.2492
R1240 VN.n1 VN.t3 75.2492
R1241 VN VN.n1 45.9715
R1242 VN VN.n0 2.64952
R1243 VDD2.n2 VDD2.n0 108.969
R1244 VDD2.n2 VDD2.n1 71.4264
R1245 VDD2.n1 VDD2.t0 3.59397
R1246 VDD2.n1 VDD2.t2 3.59397
R1247 VDD2.n0 VDD2.t1 3.59397
R1248 VDD2.n0 VDD2.t3 3.59397
R1249 VDD2 VDD2.n2 0.0586897
C0 VP VDD2 0.431056f
C1 VTAIL VP 2.88279f
C2 VN VDD1 0.149368f
C3 VDD2 VN 2.43689f
C4 VDD2 VDD1 1.16766f
C5 VTAIL VN 2.86868f
C6 VP VN 5.41131f
C7 VTAIL VDD1 4.10636f
C8 VP VDD1 2.71769f
C9 VTAIL VDD2 4.16446f
C10 VDD2 B 3.5921f
C11 VDD1 B 7.35412f
C12 VTAIL B 6.180125f
C13 VN B 11.27217f
C14 VP B 9.598896f
C15 VDD2.t1 B 0.122608f
C16 VDD2.t3 B 0.122608f
C17 VDD2.n0 B 1.48111f
C18 VDD2.t0 B 0.122608f
C19 VDD2.t2 B 0.122608f
C20 VDD2.n1 B 1.02383f
C21 VDD2.n2 B 3.32401f
C22 VN.t0 B 1.48354f
C23 VN.t2 B 1.49256f
C24 VN.n0 B 0.896601f
C25 VN.t3 B 1.48354f
C26 VN.t1 B 1.49256f
C27 VN.n1 B 2.27859f
C28 VTAIL.t2 B 0.907382f
C29 VTAIL.n0 B 0.369115f
C30 VTAIL.t4 B 0.907382f
C31 VTAIL.n1 B 0.467099f
C32 VTAIL.t5 B 0.907382f
C33 VTAIL.n2 B 1.24314f
C34 VTAIL.t3 B 0.907382f
C35 VTAIL.n3 B 1.24314f
C36 VTAIL.t1 B 0.907382f
C37 VTAIL.n4 B 0.467098f
C38 VTAIL.t7 B 0.907382f
C39 VTAIL.n5 B 0.467098f
C40 VTAIL.t6 B 0.907378f
C41 VTAIL.n6 B 1.24314f
C42 VTAIL.t0 B 0.907382f
C43 VTAIL.n7 B 1.13731f
C44 VDD1.t2 B 0.124364f
C45 VDD1.t1 B 0.124364f
C46 VDD1.n0 B 1.03891f
C47 VDD1.t3 B 0.124364f
C48 VDD1.t0 B 0.124364f
C49 VDD1.n1 B 1.52644f
C50 VP.t3 B 1.24039f
C51 VP.n0 B 0.563567f
C52 VP.n1 B 0.026887f
C53 VP.n2 B 0.021736f
C54 VP.n3 B 0.026887f
C55 VP.t2 B 1.24039f
C56 VP.n4 B 0.563567f
C57 VP.t0 B 1.53967f
C58 VP.t1 B 1.53038f
C59 VP.n5 B 2.33925f
C60 VP.n6 B 1.3411f
C61 VP.n7 B 0.043395f
C62 VP.n8 B 0.037986f
C63 VP.n9 B 0.05011f
C64 VP.n10 B 0.053437f
C65 VP.n11 B 0.026887f
C66 VP.n12 B 0.026887f
C67 VP.n13 B 0.026887f
C68 VP.n14 B 0.053437f
C69 VP.n15 B 0.05011f
C70 VP.n16 B 0.037986f
C71 VP.n17 B 0.043395f
C72 VP.n18 B 0.065915f
.ends

