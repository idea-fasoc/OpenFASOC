* NGSPICE file created from diff_pair_sample_1663.ext - technology: sky130A

.subckt diff_pair_sample_1663 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t9 VN.t0 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=2.44035 ps=15.12 w=14.79 l=1.41
X1 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=0 ps=0 w=14.79 l=1.41
X2 VDD2.t1 VN.t1 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=5.7681 ps=30.36 w=14.79 l=1.41
X3 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=0 ps=0 w=14.79 l=1.41
X4 VDD1.t5 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=2.44035 ps=15.12 w=14.79 l=1.41
X5 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=2.44035 ps=15.12 w=14.79 l=1.41
X6 VDD2.t2 VN.t2 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=2.44035 ps=15.12 w=14.79 l=1.41
X7 VDD1.t3 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=5.7681 ps=30.36 w=14.79 l=1.41
X8 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=0 ps=0 w=14.79 l=1.41
X9 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=0 ps=0 w=14.79 l=1.41
X10 VDD1.t2 VP.t3 VTAIL.t11 B.t4 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=5.7681 ps=30.36 w=14.79 l=1.41
X11 VDD2.t5 VN.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=5.7681 ps=30.36 w=14.79 l=1.41
X12 VTAIL.t5 VN.t4 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=2.44035 ps=15.12 w=14.79 l=1.41
X13 VTAIL.t10 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=2.44035 ps=15.12 w=14.79 l=1.41
X14 VDD2.t0 VN.t5 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7681 pd=30.36 as=2.44035 ps=15.12 w=14.79 l=1.41
X15 VTAIL.t1 VP.t5 VDD1.t0 B.t1 sky130_fd_pr__nfet_01v8 ad=2.44035 pd=15.12 as=2.44035 ps=15.12 w=14.79 l=1.41
R0 VN.n3 VN.t2 287.901
R1 VN.n13 VN.t3 287.901
R2 VN.n2 VN.t4 252.794
R3 VN.n8 VN.t1 252.794
R4 VN.n12 VN.t0 252.794
R5 VN.n18 VN.t5 252.794
R6 VN.n9 VN.n8 174.024
R7 VN.n19 VN.n18 174.024
R8 VN.n17 VN.n10 161.3
R9 VN.n16 VN.n15 161.3
R10 VN.n14 VN.n11 161.3
R11 VN.n7 VN.n0 161.3
R12 VN.n6 VN.n5 161.3
R13 VN.n4 VN.n1 161.3
R14 VN.n6 VN.n1 53.1199
R15 VN.n16 VN.n11 53.1199
R16 VN VN.n19 46.4342
R17 VN.n3 VN.n2 41.8164
R18 VN.n13 VN.n12 41.8164
R19 VN.n7 VN.n6 27.8669
R20 VN.n17 VN.n16 27.8669
R21 VN.n2 VN.n1 24.4675
R22 VN.n12 VN.n11 24.4675
R23 VN.n14 VN.n13 17.5844
R24 VN.n4 VN.n3 17.5844
R25 VN.n8 VN.n7 11.7447
R26 VN.n18 VN.n17 11.7447
R27 VN.n19 VN.n10 0.189894
R28 VN.n15 VN.n10 0.189894
R29 VN.n15 VN.n14 0.189894
R30 VN.n5 VN.n4 0.189894
R31 VN.n5 VN.n0 0.189894
R32 VN.n9 VN.n0 0.189894
R33 VN VN.n9 0.0516364
R34 VDD2.n159 VDD2.n83 289.615
R35 VDD2.n76 VDD2.n0 289.615
R36 VDD2.n160 VDD2.n159 185
R37 VDD2.n158 VDD2.n157 185
R38 VDD2.n156 VDD2.n86 185
R39 VDD2.n90 VDD2.n87 185
R40 VDD2.n151 VDD2.n150 185
R41 VDD2.n149 VDD2.n148 185
R42 VDD2.n92 VDD2.n91 185
R43 VDD2.n143 VDD2.n142 185
R44 VDD2.n141 VDD2.n140 185
R45 VDD2.n96 VDD2.n95 185
R46 VDD2.n135 VDD2.n134 185
R47 VDD2.n133 VDD2.n132 185
R48 VDD2.n100 VDD2.n99 185
R49 VDD2.n127 VDD2.n126 185
R50 VDD2.n125 VDD2.n124 185
R51 VDD2.n104 VDD2.n103 185
R52 VDD2.n119 VDD2.n118 185
R53 VDD2.n117 VDD2.n116 185
R54 VDD2.n108 VDD2.n107 185
R55 VDD2.n111 VDD2.n110 185
R56 VDD2.n27 VDD2.n26 185
R57 VDD2.n24 VDD2.n23 185
R58 VDD2.n33 VDD2.n32 185
R59 VDD2.n35 VDD2.n34 185
R60 VDD2.n20 VDD2.n19 185
R61 VDD2.n41 VDD2.n40 185
R62 VDD2.n43 VDD2.n42 185
R63 VDD2.n16 VDD2.n15 185
R64 VDD2.n49 VDD2.n48 185
R65 VDD2.n51 VDD2.n50 185
R66 VDD2.n12 VDD2.n11 185
R67 VDD2.n57 VDD2.n56 185
R68 VDD2.n59 VDD2.n58 185
R69 VDD2.n8 VDD2.n7 185
R70 VDD2.n65 VDD2.n64 185
R71 VDD2.n68 VDD2.n67 185
R72 VDD2.n66 VDD2.n4 185
R73 VDD2.n73 VDD2.n3 185
R74 VDD2.n75 VDD2.n74 185
R75 VDD2.n77 VDD2.n76 185
R76 VDD2.t0 VDD2.n109 147.659
R77 VDD2.t2 VDD2.n25 147.659
R78 VDD2.n159 VDD2.n158 104.615
R79 VDD2.n158 VDD2.n86 104.615
R80 VDD2.n90 VDD2.n86 104.615
R81 VDD2.n150 VDD2.n90 104.615
R82 VDD2.n150 VDD2.n149 104.615
R83 VDD2.n149 VDD2.n91 104.615
R84 VDD2.n142 VDD2.n91 104.615
R85 VDD2.n142 VDD2.n141 104.615
R86 VDD2.n141 VDD2.n95 104.615
R87 VDD2.n134 VDD2.n95 104.615
R88 VDD2.n134 VDD2.n133 104.615
R89 VDD2.n133 VDD2.n99 104.615
R90 VDD2.n126 VDD2.n99 104.615
R91 VDD2.n126 VDD2.n125 104.615
R92 VDD2.n125 VDD2.n103 104.615
R93 VDD2.n118 VDD2.n103 104.615
R94 VDD2.n118 VDD2.n117 104.615
R95 VDD2.n117 VDD2.n107 104.615
R96 VDD2.n110 VDD2.n107 104.615
R97 VDD2.n26 VDD2.n23 104.615
R98 VDD2.n33 VDD2.n23 104.615
R99 VDD2.n34 VDD2.n33 104.615
R100 VDD2.n34 VDD2.n19 104.615
R101 VDD2.n41 VDD2.n19 104.615
R102 VDD2.n42 VDD2.n41 104.615
R103 VDD2.n42 VDD2.n15 104.615
R104 VDD2.n49 VDD2.n15 104.615
R105 VDD2.n50 VDD2.n49 104.615
R106 VDD2.n50 VDD2.n11 104.615
R107 VDD2.n57 VDD2.n11 104.615
R108 VDD2.n58 VDD2.n57 104.615
R109 VDD2.n58 VDD2.n7 104.615
R110 VDD2.n65 VDD2.n7 104.615
R111 VDD2.n67 VDD2.n65 104.615
R112 VDD2.n67 VDD2.n66 104.615
R113 VDD2.n66 VDD2.n3 104.615
R114 VDD2.n75 VDD2.n3 104.615
R115 VDD2.n76 VDD2.n75 104.615
R116 VDD2.n82 VDD2.n81 64.1497
R117 VDD2 VDD2.n165 64.1468
R118 VDD2.n82 VDD2.n80 52.8429
R119 VDD2.n110 VDD2.t0 52.3082
R120 VDD2.n26 VDD2.t2 52.3082
R121 VDD2.n164 VDD2.n163 51.7732
R122 VDD2.n164 VDD2.n82 41.3403
R123 VDD2.n111 VDD2.n109 15.6677
R124 VDD2.n27 VDD2.n25 15.6677
R125 VDD2.n157 VDD2.n156 13.1884
R126 VDD2.n74 VDD2.n73 13.1884
R127 VDD2.n160 VDD2.n85 12.8005
R128 VDD2.n155 VDD2.n87 12.8005
R129 VDD2.n112 VDD2.n108 12.8005
R130 VDD2.n28 VDD2.n24 12.8005
R131 VDD2.n72 VDD2.n4 12.8005
R132 VDD2.n77 VDD2.n2 12.8005
R133 VDD2.n161 VDD2.n83 12.0247
R134 VDD2.n152 VDD2.n151 12.0247
R135 VDD2.n116 VDD2.n115 12.0247
R136 VDD2.n32 VDD2.n31 12.0247
R137 VDD2.n69 VDD2.n68 12.0247
R138 VDD2.n78 VDD2.n0 12.0247
R139 VDD2.n148 VDD2.n89 11.249
R140 VDD2.n119 VDD2.n106 11.249
R141 VDD2.n35 VDD2.n22 11.249
R142 VDD2.n64 VDD2.n6 11.249
R143 VDD2.n147 VDD2.n92 10.4732
R144 VDD2.n120 VDD2.n104 10.4732
R145 VDD2.n36 VDD2.n20 10.4732
R146 VDD2.n63 VDD2.n8 10.4732
R147 VDD2.n144 VDD2.n143 9.69747
R148 VDD2.n124 VDD2.n123 9.69747
R149 VDD2.n40 VDD2.n39 9.69747
R150 VDD2.n60 VDD2.n59 9.69747
R151 VDD2.n163 VDD2.n162 9.45567
R152 VDD2.n80 VDD2.n79 9.45567
R153 VDD2.n137 VDD2.n136 9.3005
R154 VDD2.n139 VDD2.n138 9.3005
R155 VDD2.n94 VDD2.n93 9.3005
R156 VDD2.n145 VDD2.n144 9.3005
R157 VDD2.n147 VDD2.n146 9.3005
R158 VDD2.n89 VDD2.n88 9.3005
R159 VDD2.n153 VDD2.n152 9.3005
R160 VDD2.n155 VDD2.n154 9.3005
R161 VDD2.n162 VDD2.n161 9.3005
R162 VDD2.n85 VDD2.n84 9.3005
R163 VDD2.n98 VDD2.n97 9.3005
R164 VDD2.n131 VDD2.n130 9.3005
R165 VDD2.n129 VDD2.n128 9.3005
R166 VDD2.n102 VDD2.n101 9.3005
R167 VDD2.n123 VDD2.n122 9.3005
R168 VDD2.n121 VDD2.n120 9.3005
R169 VDD2.n106 VDD2.n105 9.3005
R170 VDD2.n115 VDD2.n114 9.3005
R171 VDD2.n113 VDD2.n112 9.3005
R172 VDD2.n79 VDD2.n78 9.3005
R173 VDD2.n2 VDD2.n1 9.3005
R174 VDD2.n47 VDD2.n46 9.3005
R175 VDD2.n45 VDD2.n44 9.3005
R176 VDD2.n18 VDD2.n17 9.3005
R177 VDD2.n39 VDD2.n38 9.3005
R178 VDD2.n37 VDD2.n36 9.3005
R179 VDD2.n22 VDD2.n21 9.3005
R180 VDD2.n31 VDD2.n30 9.3005
R181 VDD2.n29 VDD2.n28 9.3005
R182 VDD2.n14 VDD2.n13 9.3005
R183 VDD2.n53 VDD2.n52 9.3005
R184 VDD2.n55 VDD2.n54 9.3005
R185 VDD2.n10 VDD2.n9 9.3005
R186 VDD2.n61 VDD2.n60 9.3005
R187 VDD2.n63 VDD2.n62 9.3005
R188 VDD2.n6 VDD2.n5 9.3005
R189 VDD2.n70 VDD2.n69 9.3005
R190 VDD2.n72 VDD2.n71 9.3005
R191 VDD2.n140 VDD2.n94 8.92171
R192 VDD2.n127 VDD2.n102 8.92171
R193 VDD2.n43 VDD2.n18 8.92171
R194 VDD2.n56 VDD2.n10 8.92171
R195 VDD2.n139 VDD2.n96 8.14595
R196 VDD2.n128 VDD2.n100 8.14595
R197 VDD2.n44 VDD2.n16 8.14595
R198 VDD2.n55 VDD2.n12 8.14595
R199 VDD2.n136 VDD2.n135 7.3702
R200 VDD2.n132 VDD2.n131 7.3702
R201 VDD2.n48 VDD2.n47 7.3702
R202 VDD2.n52 VDD2.n51 7.3702
R203 VDD2.n135 VDD2.n98 6.59444
R204 VDD2.n132 VDD2.n98 6.59444
R205 VDD2.n48 VDD2.n14 6.59444
R206 VDD2.n51 VDD2.n14 6.59444
R207 VDD2.n136 VDD2.n96 5.81868
R208 VDD2.n131 VDD2.n100 5.81868
R209 VDD2.n47 VDD2.n16 5.81868
R210 VDD2.n52 VDD2.n12 5.81868
R211 VDD2.n140 VDD2.n139 5.04292
R212 VDD2.n128 VDD2.n127 5.04292
R213 VDD2.n44 VDD2.n43 5.04292
R214 VDD2.n56 VDD2.n55 5.04292
R215 VDD2.n113 VDD2.n109 4.38563
R216 VDD2.n29 VDD2.n25 4.38563
R217 VDD2.n143 VDD2.n94 4.26717
R218 VDD2.n124 VDD2.n102 4.26717
R219 VDD2.n40 VDD2.n18 4.26717
R220 VDD2.n59 VDD2.n10 4.26717
R221 VDD2.n144 VDD2.n92 3.49141
R222 VDD2.n123 VDD2.n104 3.49141
R223 VDD2.n39 VDD2.n20 3.49141
R224 VDD2.n60 VDD2.n8 3.49141
R225 VDD2.n148 VDD2.n147 2.71565
R226 VDD2.n120 VDD2.n119 2.71565
R227 VDD2.n36 VDD2.n35 2.71565
R228 VDD2.n64 VDD2.n63 2.71565
R229 VDD2.n163 VDD2.n83 1.93989
R230 VDD2.n151 VDD2.n89 1.93989
R231 VDD2.n116 VDD2.n106 1.93989
R232 VDD2.n32 VDD2.n22 1.93989
R233 VDD2.n68 VDD2.n6 1.93989
R234 VDD2.n80 VDD2.n0 1.93989
R235 VDD2.n165 VDD2.t3 1.33924
R236 VDD2.n165 VDD2.t5 1.33924
R237 VDD2.n81 VDD2.t4 1.33924
R238 VDD2.n81 VDD2.t1 1.33924
R239 VDD2 VDD2.n164 1.18369
R240 VDD2.n161 VDD2.n160 1.16414
R241 VDD2.n152 VDD2.n87 1.16414
R242 VDD2.n115 VDD2.n108 1.16414
R243 VDD2.n31 VDD2.n24 1.16414
R244 VDD2.n69 VDD2.n4 1.16414
R245 VDD2.n78 VDD2.n77 1.16414
R246 VDD2.n157 VDD2.n85 0.388379
R247 VDD2.n156 VDD2.n155 0.388379
R248 VDD2.n112 VDD2.n111 0.388379
R249 VDD2.n28 VDD2.n27 0.388379
R250 VDD2.n73 VDD2.n72 0.388379
R251 VDD2.n74 VDD2.n2 0.388379
R252 VDD2.n162 VDD2.n84 0.155672
R253 VDD2.n154 VDD2.n84 0.155672
R254 VDD2.n154 VDD2.n153 0.155672
R255 VDD2.n153 VDD2.n88 0.155672
R256 VDD2.n146 VDD2.n88 0.155672
R257 VDD2.n146 VDD2.n145 0.155672
R258 VDD2.n145 VDD2.n93 0.155672
R259 VDD2.n138 VDD2.n93 0.155672
R260 VDD2.n138 VDD2.n137 0.155672
R261 VDD2.n137 VDD2.n97 0.155672
R262 VDD2.n130 VDD2.n97 0.155672
R263 VDD2.n130 VDD2.n129 0.155672
R264 VDD2.n129 VDD2.n101 0.155672
R265 VDD2.n122 VDD2.n101 0.155672
R266 VDD2.n122 VDD2.n121 0.155672
R267 VDD2.n121 VDD2.n105 0.155672
R268 VDD2.n114 VDD2.n105 0.155672
R269 VDD2.n114 VDD2.n113 0.155672
R270 VDD2.n30 VDD2.n29 0.155672
R271 VDD2.n30 VDD2.n21 0.155672
R272 VDD2.n37 VDD2.n21 0.155672
R273 VDD2.n38 VDD2.n37 0.155672
R274 VDD2.n38 VDD2.n17 0.155672
R275 VDD2.n45 VDD2.n17 0.155672
R276 VDD2.n46 VDD2.n45 0.155672
R277 VDD2.n46 VDD2.n13 0.155672
R278 VDD2.n53 VDD2.n13 0.155672
R279 VDD2.n54 VDD2.n53 0.155672
R280 VDD2.n54 VDD2.n9 0.155672
R281 VDD2.n61 VDD2.n9 0.155672
R282 VDD2.n62 VDD2.n61 0.155672
R283 VDD2.n62 VDD2.n5 0.155672
R284 VDD2.n70 VDD2.n5 0.155672
R285 VDD2.n71 VDD2.n70 0.155672
R286 VDD2.n71 VDD2.n1 0.155672
R287 VDD2.n79 VDD2.n1 0.155672
R288 VTAIL.n330 VTAIL.n254 289.615
R289 VTAIL.n78 VTAIL.n2 289.615
R290 VTAIL.n248 VTAIL.n172 289.615
R291 VTAIL.n164 VTAIL.n88 289.615
R292 VTAIL.n281 VTAIL.n280 185
R293 VTAIL.n278 VTAIL.n277 185
R294 VTAIL.n287 VTAIL.n286 185
R295 VTAIL.n289 VTAIL.n288 185
R296 VTAIL.n274 VTAIL.n273 185
R297 VTAIL.n295 VTAIL.n294 185
R298 VTAIL.n297 VTAIL.n296 185
R299 VTAIL.n270 VTAIL.n269 185
R300 VTAIL.n303 VTAIL.n302 185
R301 VTAIL.n305 VTAIL.n304 185
R302 VTAIL.n266 VTAIL.n265 185
R303 VTAIL.n311 VTAIL.n310 185
R304 VTAIL.n313 VTAIL.n312 185
R305 VTAIL.n262 VTAIL.n261 185
R306 VTAIL.n319 VTAIL.n318 185
R307 VTAIL.n322 VTAIL.n321 185
R308 VTAIL.n320 VTAIL.n258 185
R309 VTAIL.n327 VTAIL.n257 185
R310 VTAIL.n329 VTAIL.n328 185
R311 VTAIL.n331 VTAIL.n330 185
R312 VTAIL.n29 VTAIL.n28 185
R313 VTAIL.n26 VTAIL.n25 185
R314 VTAIL.n35 VTAIL.n34 185
R315 VTAIL.n37 VTAIL.n36 185
R316 VTAIL.n22 VTAIL.n21 185
R317 VTAIL.n43 VTAIL.n42 185
R318 VTAIL.n45 VTAIL.n44 185
R319 VTAIL.n18 VTAIL.n17 185
R320 VTAIL.n51 VTAIL.n50 185
R321 VTAIL.n53 VTAIL.n52 185
R322 VTAIL.n14 VTAIL.n13 185
R323 VTAIL.n59 VTAIL.n58 185
R324 VTAIL.n61 VTAIL.n60 185
R325 VTAIL.n10 VTAIL.n9 185
R326 VTAIL.n67 VTAIL.n66 185
R327 VTAIL.n70 VTAIL.n69 185
R328 VTAIL.n68 VTAIL.n6 185
R329 VTAIL.n75 VTAIL.n5 185
R330 VTAIL.n77 VTAIL.n76 185
R331 VTAIL.n79 VTAIL.n78 185
R332 VTAIL.n249 VTAIL.n248 185
R333 VTAIL.n247 VTAIL.n246 185
R334 VTAIL.n245 VTAIL.n175 185
R335 VTAIL.n179 VTAIL.n176 185
R336 VTAIL.n240 VTAIL.n239 185
R337 VTAIL.n238 VTAIL.n237 185
R338 VTAIL.n181 VTAIL.n180 185
R339 VTAIL.n232 VTAIL.n231 185
R340 VTAIL.n230 VTAIL.n229 185
R341 VTAIL.n185 VTAIL.n184 185
R342 VTAIL.n224 VTAIL.n223 185
R343 VTAIL.n222 VTAIL.n221 185
R344 VTAIL.n189 VTAIL.n188 185
R345 VTAIL.n216 VTAIL.n215 185
R346 VTAIL.n214 VTAIL.n213 185
R347 VTAIL.n193 VTAIL.n192 185
R348 VTAIL.n208 VTAIL.n207 185
R349 VTAIL.n206 VTAIL.n205 185
R350 VTAIL.n197 VTAIL.n196 185
R351 VTAIL.n200 VTAIL.n199 185
R352 VTAIL.n165 VTAIL.n164 185
R353 VTAIL.n163 VTAIL.n162 185
R354 VTAIL.n161 VTAIL.n91 185
R355 VTAIL.n95 VTAIL.n92 185
R356 VTAIL.n156 VTAIL.n155 185
R357 VTAIL.n154 VTAIL.n153 185
R358 VTAIL.n97 VTAIL.n96 185
R359 VTAIL.n148 VTAIL.n147 185
R360 VTAIL.n146 VTAIL.n145 185
R361 VTAIL.n101 VTAIL.n100 185
R362 VTAIL.n140 VTAIL.n139 185
R363 VTAIL.n138 VTAIL.n137 185
R364 VTAIL.n105 VTAIL.n104 185
R365 VTAIL.n132 VTAIL.n131 185
R366 VTAIL.n130 VTAIL.n129 185
R367 VTAIL.n109 VTAIL.n108 185
R368 VTAIL.n124 VTAIL.n123 185
R369 VTAIL.n122 VTAIL.n121 185
R370 VTAIL.n113 VTAIL.n112 185
R371 VTAIL.n116 VTAIL.n115 185
R372 VTAIL.t11 VTAIL.n198 147.659
R373 VTAIL.t6 VTAIL.n114 147.659
R374 VTAIL.t8 VTAIL.n279 147.659
R375 VTAIL.t2 VTAIL.n27 147.659
R376 VTAIL.n280 VTAIL.n277 104.615
R377 VTAIL.n287 VTAIL.n277 104.615
R378 VTAIL.n288 VTAIL.n287 104.615
R379 VTAIL.n288 VTAIL.n273 104.615
R380 VTAIL.n295 VTAIL.n273 104.615
R381 VTAIL.n296 VTAIL.n295 104.615
R382 VTAIL.n296 VTAIL.n269 104.615
R383 VTAIL.n303 VTAIL.n269 104.615
R384 VTAIL.n304 VTAIL.n303 104.615
R385 VTAIL.n304 VTAIL.n265 104.615
R386 VTAIL.n311 VTAIL.n265 104.615
R387 VTAIL.n312 VTAIL.n311 104.615
R388 VTAIL.n312 VTAIL.n261 104.615
R389 VTAIL.n319 VTAIL.n261 104.615
R390 VTAIL.n321 VTAIL.n319 104.615
R391 VTAIL.n321 VTAIL.n320 104.615
R392 VTAIL.n320 VTAIL.n257 104.615
R393 VTAIL.n329 VTAIL.n257 104.615
R394 VTAIL.n330 VTAIL.n329 104.615
R395 VTAIL.n28 VTAIL.n25 104.615
R396 VTAIL.n35 VTAIL.n25 104.615
R397 VTAIL.n36 VTAIL.n35 104.615
R398 VTAIL.n36 VTAIL.n21 104.615
R399 VTAIL.n43 VTAIL.n21 104.615
R400 VTAIL.n44 VTAIL.n43 104.615
R401 VTAIL.n44 VTAIL.n17 104.615
R402 VTAIL.n51 VTAIL.n17 104.615
R403 VTAIL.n52 VTAIL.n51 104.615
R404 VTAIL.n52 VTAIL.n13 104.615
R405 VTAIL.n59 VTAIL.n13 104.615
R406 VTAIL.n60 VTAIL.n59 104.615
R407 VTAIL.n60 VTAIL.n9 104.615
R408 VTAIL.n67 VTAIL.n9 104.615
R409 VTAIL.n69 VTAIL.n67 104.615
R410 VTAIL.n69 VTAIL.n68 104.615
R411 VTAIL.n68 VTAIL.n5 104.615
R412 VTAIL.n77 VTAIL.n5 104.615
R413 VTAIL.n78 VTAIL.n77 104.615
R414 VTAIL.n248 VTAIL.n247 104.615
R415 VTAIL.n247 VTAIL.n175 104.615
R416 VTAIL.n179 VTAIL.n175 104.615
R417 VTAIL.n239 VTAIL.n179 104.615
R418 VTAIL.n239 VTAIL.n238 104.615
R419 VTAIL.n238 VTAIL.n180 104.615
R420 VTAIL.n231 VTAIL.n180 104.615
R421 VTAIL.n231 VTAIL.n230 104.615
R422 VTAIL.n230 VTAIL.n184 104.615
R423 VTAIL.n223 VTAIL.n184 104.615
R424 VTAIL.n223 VTAIL.n222 104.615
R425 VTAIL.n222 VTAIL.n188 104.615
R426 VTAIL.n215 VTAIL.n188 104.615
R427 VTAIL.n215 VTAIL.n214 104.615
R428 VTAIL.n214 VTAIL.n192 104.615
R429 VTAIL.n207 VTAIL.n192 104.615
R430 VTAIL.n207 VTAIL.n206 104.615
R431 VTAIL.n206 VTAIL.n196 104.615
R432 VTAIL.n199 VTAIL.n196 104.615
R433 VTAIL.n164 VTAIL.n163 104.615
R434 VTAIL.n163 VTAIL.n91 104.615
R435 VTAIL.n95 VTAIL.n91 104.615
R436 VTAIL.n155 VTAIL.n95 104.615
R437 VTAIL.n155 VTAIL.n154 104.615
R438 VTAIL.n154 VTAIL.n96 104.615
R439 VTAIL.n147 VTAIL.n96 104.615
R440 VTAIL.n147 VTAIL.n146 104.615
R441 VTAIL.n146 VTAIL.n100 104.615
R442 VTAIL.n139 VTAIL.n100 104.615
R443 VTAIL.n139 VTAIL.n138 104.615
R444 VTAIL.n138 VTAIL.n104 104.615
R445 VTAIL.n131 VTAIL.n104 104.615
R446 VTAIL.n131 VTAIL.n130 104.615
R447 VTAIL.n130 VTAIL.n108 104.615
R448 VTAIL.n123 VTAIL.n108 104.615
R449 VTAIL.n123 VTAIL.n122 104.615
R450 VTAIL.n122 VTAIL.n112 104.615
R451 VTAIL.n115 VTAIL.n112 104.615
R452 VTAIL.n280 VTAIL.t8 52.3082
R453 VTAIL.n28 VTAIL.t2 52.3082
R454 VTAIL.n199 VTAIL.t11 52.3082
R455 VTAIL.n115 VTAIL.t6 52.3082
R456 VTAIL.n171 VTAIL.n170 47.1514
R457 VTAIL.n87 VTAIL.n86 47.1514
R458 VTAIL.n1 VTAIL.n0 47.1512
R459 VTAIL.n85 VTAIL.n84 47.1512
R460 VTAIL.n335 VTAIL.n334 35.0944
R461 VTAIL.n83 VTAIL.n82 35.0944
R462 VTAIL.n253 VTAIL.n252 35.0944
R463 VTAIL.n169 VTAIL.n168 35.0944
R464 VTAIL.n87 VTAIL.n85 28.1169
R465 VTAIL.n335 VTAIL.n253 26.6169
R466 VTAIL.n281 VTAIL.n279 15.6677
R467 VTAIL.n29 VTAIL.n27 15.6677
R468 VTAIL.n200 VTAIL.n198 15.6677
R469 VTAIL.n116 VTAIL.n114 15.6677
R470 VTAIL.n328 VTAIL.n327 13.1884
R471 VTAIL.n76 VTAIL.n75 13.1884
R472 VTAIL.n246 VTAIL.n245 13.1884
R473 VTAIL.n162 VTAIL.n161 13.1884
R474 VTAIL.n282 VTAIL.n278 12.8005
R475 VTAIL.n326 VTAIL.n258 12.8005
R476 VTAIL.n331 VTAIL.n256 12.8005
R477 VTAIL.n30 VTAIL.n26 12.8005
R478 VTAIL.n74 VTAIL.n6 12.8005
R479 VTAIL.n79 VTAIL.n4 12.8005
R480 VTAIL.n249 VTAIL.n174 12.8005
R481 VTAIL.n244 VTAIL.n176 12.8005
R482 VTAIL.n201 VTAIL.n197 12.8005
R483 VTAIL.n165 VTAIL.n90 12.8005
R484 VTAIL.n160 VTAIL.n92 12.8005
R485 VTAIL.n117 VTAIL.n113 12.8005
R486 VTAIL.n286 VTAIL.n285 12.0247
R487 VTAIL.n323 VTAIL.n322 12.0247
R488 VTAIL.n332 VTAIL.n254 12.0247
R489 VTAIL.n34 VTAIL.n33 12.0247
R490 VTAIL.n71 VTAIL.n70 12.0247
R491 VTAIL.n80 VTAIL.n2 12.0247
R492 VTAIL.n250 VTAIL.n172 12.0247
R493 VTAIL.n241 VTAIL.n240 12.0247
R494 VTAIL.n205 VTAIL.n204 12.0247
R495 VTAIL.n166 VTAIL.n88 12.0247
R496 VTAIL.n157 VTAIL.n156 12.0247
R497 VTAIL.n121 VTAIL.n120 12.0247
R498 VTAIL.n289 VTAIL.n276 11.249
R499 VTAIL.n318 VTAIL.n260 11.249
R500 VTAIL.n37 VTAIL.n24 11.249
R501 VTAIL.n66 VTAIL.n8 11.249
R502 VTAIL.n237 VTAIL.n178 11.249
R503 VTAIL.n208 VTAIL.n195 11.249
R504 VTAIL.n153 VTAIL.n94 11.249
R505 VTAIL.n124 VTAIL.n111 11.249
R506 VTAIL.n290 VTAIL.n274 10.4732
R507 VTAIL.n317 VTAIL.n262 10.4732
R508 VTAIL.n38 VTAIL.n22 10.4732
R509 VTAIL.n65 VTAIL.n10 10.4732
R510 VTAIL.n236 VTAIL.n181 10.4732
R511 VTAIL.n209 VTAIL.n193 10.4732
R512 VTAIL.n152 VTAIL.n97 10.4732
R513 VTAIL.n125 VTAIL.n109 10.4732
R514 VTAIL.n294 VTAIL.n293 9.69747
R515 VTAIL.n314 VTAIL.n313 9.69747
R516 VTAIL.n42 VTAIL.n41 9.69747
R517 VTAIL.n62 VTAIL.n61 9.69747
R518 VTAIL.n233 VTAIL.n232 9.69747
R519 VTAIL.n213 VTAIL.n212 9.69747
R520 VTAIL.n149 VTAIL.n148 9.69747
R521 VTAIL.n129 VTAIL.n128 9.69747
R522 VTAIL.n334 VTAIL.n333 9.45567
R523 VTAIL.n82 VTAIL.n81 9.45567
R524 VTAIL.n252 VTAIL.n251 9.45567
R525 VTAIL.n168 VTAIL.n167 9.45567
R526 VTAIL.n333 VTAIL.n332 9.3005
R527 VTAIL.n256 VTAIL.n255 9.3005
R528 VTAIL.n301 VTAIL.n300 9.3005
R529 VTAIL.n299 VTAIL.n298 9.3005
R530 VTAIL.n272 VTAIL.n271 9.3005
R531 VTAIL.n293 VTAIL.n292 9.3005
R532 VTAIL.n291 VTAIL.n290 9.3005
R533 VTAIL.n276 VTAIL.n275 9.3005
R534 VTAIL.n285 VTAIL.n284 9.3005
R535 VTAIL.n283 VTAIL.n282 9.3005
R536 VTAIL.n268 VTAIL.n267 9.3005
R537 VTAIL.n307 VTAIL.n306 9.3005
R538 VTAIL.n309 VTAIL.n308 9.3005
R539 VTAIL.n264 VTAIL.n263 9.3005
R540 VTAIL.n315 VTAIL.n314 9.3005
R541 VTAIL.n317 VTAIL.n316 9.3005
R542 VTAIL.n260 VTAIL.n259 9.3005
R543 VTAIL.n324 VTAIL.n323 9.3005
R544 VTAIL.n326 VTAIL.n325 9.3005
R545 VTAIL.n81 VTAIL.n80 9.3005
R546 VTAIL.n4 VTAIL.n3 9.3005
R547 VTAIL.n49 VTAIL.n48 9.3005
R548 VTAIL.n47 VTAIL.n46 9.3005
R549 VTAIL.n20 VTAIL.n19 9.3005
R550 VTAIL.n41 VTAIL.n40 9.3005
R551 VTAIL.n39 VTAIL.n38 9.3005
R552 VTAIL.n24 VTAIL.n23 9.3005
R553 VTAIL.n33 VTAIL.n32 9.3005
R554 VTAIL.n31 VTAIL.n30 9.3005
R555 VTAIL.n16 VTAIL.n15 9.3005
R556 VTAIL.n55 VTAIL.n54 9.3005
R557 VTAIL.n57 VTAIL.n56 9.3005
R558 VTAIL.n12 VTAIL.n11 9.3005
R559 VTAIL.n63 VTAIL.n62 9.3005
R560 VTAIL.n65 VTAIL.n64 9.3005
R561 VTAIL.n8 VTAIL.n7 9.3005
R562 VTAIL.n72 VTAIL.n71 9.3005
R563 VTAIL.n74 VTAIL.n73 9.3005
R564 VTAIL.n226 VTAIL.n225 9.3005
R565 VTAIL.n228 VTAIL.n227 9.3005
R566 VTAIL.n183 VTAIL.n182 9.3005
R567 VTAIL.n234 VTAIL.n233 9.3005
R568 VTAIL.n236 VTAIL.n235 9.3005
R569 VTAIL.n178 VTAIL.n177 9.3005
R570 VTAIL.n242 VTAIL.n241 9.3005
R571 VTAIL.n244 VTAIL.n243 9.3005
R572 VTAIL.n251 VTAIL.n250 9.3005
R573 VTAIL.n174 VTAIL.n173 9.3005
R574 VTAIL.n187 VTAIL.n186 9.3005
R575 VTAIL.n220 VTAIL.n219 9.3005
R576 VTAIL.n218 VTAIL.n217 9.3005
R577 VTAIL.n191 VTAIL.n190 9.3005
R578 VTAIL.n212 VTAIL.n211 9.3005
R579 VTAIL.n210 VTAIL.n209 9.3005
R580 VTAIL.n195 VTAIL.n194 9.3005
R581 VTAIL.n204 VTAIL.n203 9.3005
R582 VTAIL.n202 VTAIL.n201 9.3005
R583 VTAIL.n142 VTAIL.n141 9.3005
R584 VTAIL.n144 VTAIL.n143 9.3005
R585 VTAIL.n99 VTAIL.n98 9.3005
R586 VTAIL.n150 VTAIL.n149 9.3005
R587 VTAIL.n152 VTAIL.n151 9.3005
R588 VTAIL.n94 VTAIL.n93 9.3005
R589 VTAIL.n158 VTAIL.n157 9.3005
R590 VTAIL.n160 VTAIL.n159 9.3005
R591 VTAIL.n167 VTAIL.n166 9.3005
R592 VTAIL.n90 VTAIL.n89 9.3005
R593 VTAIL.n103 VTAIL.n102 9.3005
R594 VTAIL.n136 VTAIL.n135 9.3005
R595 VTAIL.n134 VTAIL.n133 9.3005
R596 VTAIL.n107 VTAIL.n106 9.3005
R597 VTAIL.n128 VTAIL.n127 9.3005
R598 VTAIL.n126 VTAIL.n125 9.3005
R599 VTAIL.n111 VTAIL.n110 9.3005
R600 VTAIL.n120 VTAIL.n119 9.3005
R601 VTAIL.n118 VTAIL.n117 9.3005
R602 VTAIL.n297 VTAIL.n272 8.92171
R603 VTAIL.n310 VTAIL.n264 8.92171
R604 VTAIL.n45 VTAIL.n20 8.92171
R605 VTAIL.n58 VTAIL.n12 8.92171
R606 VTAIL.n229 VTAIL.n183 8.92171
R607 VTAIL.n216 VTAIL.n191 8.92171
R608 VTAIL.n145 VTAIL.n99 8.92171
R609 VTAIL.n132 VTAIL.n107 8.92171
R610 VTAIL.n298 VTAIL.n270 8.14595
R611 VTAIL.n309 VTAIL.n266 8.14595
R612 VTAIL.n46 VTAIL.n18 8.14595
R613 VTAIL.n57 VTAIL.n14 8.14595
R614 VTAIL.n228 VTAIL.n185 8.14595
R615 VTAIL.n217 VTAIL.n189 8.14595
R616 VTAIL.n144 VTAIL.n101 8.14595
R617 VTAIL.n133 VTAIL.n105 8.14595
R618 VTAIL.n302 VTAIL.n301 7.3702
R619 VTAIL.n306 VTAIL.n305 7.3702
R620 VTAIL.n50 VTAIL.n49 7.3702
R621 VTAIL.n54 VTAIL.n53 7.3702
R622 VTAIL.n225 VTAIL.n224 7.3702
R623 VTAIL.n221 VTAIL.n220 7.3702
R624 VTAIL.n141 VTAIL.n140 7.3702
R625 VTAIL.n137 VTAIL.n136 7.3702
R626 VTAIL.n302 VTAIL.n268 6.59444
R627 VTAIL.n305 VTAIL.n268 6.59444
R628 VTAIL.n50 VTAIL.n16 6.59444
R629 VTAIL.n53 VTAIL.n16 6.59444
R630 VTAIL.n224 VTAIL.n187 6.59444
R631 VTAIL.n221 VTAIL.n187 6.59444
R632 VTAIL.n140 VTAIL.n103 6.59444
R633 VTAIL.n137 VTAIL.n103 6.59444
R634 VTAIL.n301 VTAIL.n270 5.81868
R635 VTAIL.n306 VTAIL.n266 5.81868
R636 VTAIL.n49 VTAIL.n18 5.81868
R637 VTAIL.n54 VTAIL.n14 5.81868
R638 VTAIL.n225 VTAIL.n185 5.81868
R639 VTAIL.n220 VTAIL.n189 5.81868
R640 VTAIL.n141 VTAIL.n101 5.81868
R641 VTAIL.n136 VTAIL.n105 5.81868
R642 VTAIL.n298 VTAIL.n297 5.04292
R643 VTAIL.n310 VTAIL.n309 5.04292
R644 VTAIL.n46 VTAIL.n45 5.04292
R645 VTAIL.n58 VTAIL.n57 5.04292
R646 VTAIL.n229 VTAIL.n228 5.04292
R647 VTAIL.n217 VTAIL.n216 5.04292
R648 VTAIL.n145 VTAIL.n144 5.04292
R649 VTAIL.n133 VTAIL.n132 5.04292
R650 VTAIL.n202 VTAIL.n198 4.38563
R651 VTAIL.n118 VTAIL.n114 4.38563
R652 VTAIL.n283 VTAIL.n279 4.38563
R653 VTAIL.n31 VTAIL.n27 4.38563
R654 VTAIL.n294 VTAIL.n272 4.26717
R655 VTAIL.n313 VTAIL.n264 4.26717
R656 VTAIL.n42 VTAIL.n20 4.26717
R657 VTAIL.n61 VTAIL.n12 4.26717
R658 VTAIL.n232 VTAIL.n183 4.26717
R659 VTAIL.n213 VTAIL.n191 4.26717
R660 VTAIL.n148 VTAIL.n99 4.26717
R661 VTAIL.n129 VTAIL.n107 4.26717
R662 VTAIL.n293 VTAIL.n274 3.49141
R663 VTAIL.n314 VTAIL.n262 3.49141
R664 VTAIL.n41 VTAIL.n22 3.49141
R665 VTAIL.n62 VTAIL.n10 3.49141
R666 VTAIL.n233 VTAIL.n181 3.49141
R667 VTAIL.n212 VTAIL.n193 3.49141
R668 VTAIL.n149 VTAIL.n97 3.49141
R669 VTAIL.n128 VTAIL.n109 3.49141
R670 VTAIL.n290 VTAIL.n289 2.71565
R671 VTAIL.n318 VTAIL.n317 2.71565
R672 VTAIL.n38 VTAIL.n37 2.71565
R673 VTAIL.n66 VTAIL.n65 2.71565
R674 VTAIL.n237 VTAIL.n236 2.71565
R675 VTAIL.n209 VTAIL.n208 2.71565
R676 VTAIL.n153 VTAIL.n152 2.71565
R677 VTAIL.n125 VTAIL.n124 2.71565
R678 VTAIL.n286 VTAIL.n276 1.93989
R679 VTAIL.n322 VTAIL.n260 1.93989
R680 VTAIL.n334 VTAIL.n254 1.93989
R681 VTAIL.n34 VTAIL.n24 1.93989
R682 VTAIL.n70 VTAIL.n8 1.93989
R683 VTAIL.n82 VTAIL.n2 1.93989
R684 VTAIL.n252 VTAIL.n172 1.93989
R685 VTAIL.n240 VTAIL.n178 1.93989
R686 VTAIL.n205 VTAIL.n195 1.93989
R687 VTAIL.n168 VTAIL.n88 1.93989
R688 VTAIL.n156 VTAIL.n94 1.93989
R689 VTAIL.n121 VTAIL.n111 1.93989
R690 VTAIL.n169 VTAIL.n87 1.5005
R691 VTAIL.n253 VTAIL.n171 1.5005
R692 VTAIL.n85 VTAIL.n83 1.5005
R693 VTAIL.n0 VTAIL.t7 1.33924
R694 VTAIL.n0 VTAIL.t5 1.33924
R695 VTAIL.n84 VTAIL.t3 1.33924
R696 VTAIL.n84 VTAIL.t10 1.33924
R697 VTAIL.n170 VTAIL.t0 1.33924
R698 VTAIL.n170 VTAIL.t1 1.33924
R699 VTAIL.n86 VTAIL.t4 1.33924
R700 VTAIL.n86 VTAIL.t9 1.33924
R701 VTAIL.n171 VTAIL.n169 1.22033
R702 VTAIL.n83 VTAIL.n1 1.22033
R703 VTAIL.n285 VTAIL.n278 1.16414
R704 VTAIL.n323 VTAIL.n258 1.16414
R705 VTAIL.n332 VTAIL.n331 1.16414
R706 VTAIL.n33 VTAIL.n26 1.16414
R707 VTAIL.n71 VTAIL.n6 1.16414
R708 VTAIL.n80 VTAIL.n79 1.16414
R709 VTAIL.n250 VTAIL.n249 1.16414
R710 VTAIL.n241 VTAIL.n176 1.16414
R711 VTAIL.n204 VTAIL.n197 1.16414
R712 VTAIL.n166 VTAIL.n165 1.16414
R713 VTAIL.n157 VTAIL.n92 1.16414
R714 VTAIL.n120 VTAIL.n113 1.16414
R715 VTAIL VTAIL.n335 1.06731
R716 VTAIL VTAIL.n1 0.43369
R717 VTAIL.n282 VTAIL.n281 0.388379
R718 VTAIL.n327 VTAIL.n326 0.388379
R719 VTAIL.n328 VTAIL.n256 0.388379
R720 VTAIL.n30 VTAIL.n29 0.388379
R721 VTAIL.n75 VTAIL.n74 0.388379
R722 VTAIL.n76 VTAIL.n4 0.388379
R723 VTAIL.n246 VTAIL.n174 0.388379
R724 VTAIL.n245 VTAIL.n244 0.388379
R725 VTAIL.n201 VTAIL.n200 0.388379
R726 VTAIL.n162 VTAIL.n90 0.388379
R727 VTAIL.n161 VTAIL.n160 0.388379
R728 VTAIL.n117 VTAIL.n116 0.388379
R729 VTAIL.n284 VTAIL.n283 0.155672
R730 VTAIL.n284 VTAIL.n275 0.155672
R731 VTAIL.n291 VTAIL.n275 0.155672
R732 VTAIL.n292 VTAIL.n291 0.155672
R733 VTAIL.n292 VTAIL.n271 0.155672
R734 VTAIL.n299 VTAIL.n271 0.155672
R735 VTAIL.n300 VTAIL.n299 0.155672
R736 VTAIL.n300 VTAIL.n267 0.155672
R737 VTAIL.n307 VTAIL.n267 0.155672
R738 VTAIL.n308 VTAIL.n307 0.155672
R739 VTAIL.n308 VTAIL.n263 0.155672
R740 VTAIL.n315 VTAIL.n263 0.155672
R741 VTAIL.n316 VTAIL.n315 0.155672
R742 VTAIL.n316 VTAIL.n259 0.155672
R743 VTAIL.n324 VTAIL.n259 0.155672
R744 VTAIL.n325 VTAIL.n324 0.155672
R745 VTAIL.n325 VTAIL.n255 0.155672
R746 VTAIL.n333 VTAIL.n255 0.155672
R747 VTAIL.n32 VTAIL.n31 0.155672
R748 VTAIL.n32 VTAIL.n23 0.155672
R749 VTAIL.n39 VTAIL.n23 0.155672
R750 VTAIL.n40 VTAIL.n39 0.155672
R751 VTAIL.n40 VTAIL.n19 0.155672
R752 VTAIL.n47 VTAIL.n19 0.155672
R753 VTAIL.n48 VTAIL.n47 0.155672
R754 VTAIL.n48 VTAIL.n15 0.155672
R755 VTAIL.n55 VTAIL.n15 0.155672
R756 VTAIL.n56 VTAIL.n55 0.155672
R757 VTAIL.n56 VTAIL.n11 0.155672
R758 VTAIL.n63 VTAIL.n11 0.155672
R759 VTAIL.n64 VTAIL.n63 0.155672
R760 VTAIL.n64 VTAIL.n7 0.155672
R761 VTAIL.n72 VTAIL.n7 0.155672
R762 VTAIL.n73 VTAIL.n72 0.155672
R763 VTAIL.n73 VTAIL.n3 0.155672
R764 VTAIL.n81 VTAIL.n3 0.155672
R765 VTAIL.n251 VTAIL.n173 0.155672
R766 VTAIL.n243 VTAIL.n173 0.155672
R767 VTAIL.n243 VTAIL.n242 0.155672
R768 VTAIL.n242 VTAIL.n177 0.155672
R769 VTAIL.n235 VTAIL.n177 0.155672
R770 VTAIL.n235 VTAIL.n234 0.155672
R771 VTAIL.n234 VTAIL.n182 0.155672
R772 VTAIL.n227 VTAIL.n182 0.155672
R773 VTAIL.n227 VTAIL.n226 0.155672
R774 VTAIL.n226 VTAIL.n186 0.155672
R775 VTAIL.n219 VTAIL.n186 0.155672
R776 VTAIL.n219 VTAIL.n218 0.155672
R777 VTAIL.n218 VTAIL.n190 0.155672
R778 VTAIL.n211 VTAIL.n190 0.155672
R779 VTAIL.n211 VTAIL.n210 0.155672
R780 VTAIL.n210 VTAIL.n194 0.155672
R781 VTAIL.n203 VTAIL.n194 0.155672
R782 VTAIL.n203 VTAIL.n202 0.155672
R783 VTAIL.n167 VTAIL.n89 0.155672
R784 VTAIL.n159 VTAIL.n89 0.155672
R785 VTAIL.n159 VTAIL.n158 0.155672
R786 VTAIL.n158 VTAIL.n93 0.155672
R787 VTAIL.n151 VTAIL.n93 0.155672
R788 VTAIL.n151 VTAIL.n150 0.155672
R789 VTAIL.n150 VTAIL.n98 0.155672
R790 VTAIL.n143 VTAIL.n98 0.155672
R791 VTAIL.n143 VTAIL.n142 0.155672
R792 VTAIL.n142 VTAIL.n102 0.155672
R793 VTAIL.n135 VTAIL.n102 0.155672
R794 VTAIL.n135 VTAIL.n134 0.155672
R795 VTAIL.n134 VTAIL.n106 0.155672
R796 VTAIL.n127 VTAIL.n106 0.155672
R797 VTAIL.n127 VTAIL.n126 0.155672
R798 VTAIL.n126 VTAIL.n110 0.155672
R799 VTAIL.n119 VTAIL.n110 0.155672
R800 VTAIL.n119 VTAIL.n118 0.155672
R801 B.n785 B.n784 585
R802 B.n786 B.n785 585
R803 B.n328 B.n109 585
R804 B.n327 B.n326 585
R805 B.n325 B.n324 585
R806 B.n323 B.n322 585
R807 B.n321 B.n320 585
R808 B.n319 B.n318 585
R809 B.n317 B.n316 585
R810 B.n315 B.n314 585
R811 B.n313 B.n312 585
R812 B.n311 B.n310 585
R813 B.n309 B.n308 585
R814 B.n307 B.n306 585
R815 B.n305 B.n304 585
R816 B.n303 B.n302 585
R817 B.n301 B.n300 585
R818 B.n299 B.n298 585
R819 B.n297 B.n296 585
R820 B.n295 B.n294 585
R821 B.n293 B.n292 585
R822 B.n291 B.n290 585
R823 B.n289 B.n288 585
R824 B.n287 B.n286 585
R825 B.n285 B.n284 585
R826 B.n283 B.n282 585
R827 B.n281 B.n280 585
R828 B.n279 B.n278 585
R829 B.n277 B.n276 585
R830 B.n275 B.n274 585
R831 B.n273 B.n272 585
R832 B.n271 B.n270 585
R833 B.n269 B.n268 585
R834 B.n267 B.n266 585
R835 B.n265 B.n264 585
R836 B.n263 B.n262 585
R837 B.n261 B.n260 585
R838 B.n259 B.n258 585
R839 B.n257 B.n256 585
R840 B.n255 B.n254 585
R841 B.n253 B.n252 585
R842 B.n251 B.n250 585
R843 B.n249 B.n248 585
R844 B.n247 B.n246 585
R845 B.n245 B.n244 585
R846 B.n243 B.n242 585
R847 B.n241 B.n240 585
R848 B.n239 B.n238 585
R849 B.n237 B.n236 585
R850 B.n235 B.n234 585
R851 B.n233 B.n232 585
R852 B.n230 B.n229 585
R853 B.n228 B.n227 585
R854 B.n226 B.n225 585
R855 B.n224 B.n223 585
R856 B.n222 B.n221 585
R857 B.n220 B.n219 585
R858 B.n218 B.n217 585
R859 B.n216 B.n215 585
R860 B.n214 B.n213 585
R861 B.n212 B.n211 585
R862 B.n210 B.n209 585
R863 B.n208 B.n207 585
R864 B.n206 B.n205 585
R865 B.n204 B.n203 585
R866 B.n202 B.n201 585
R867 B.n200 B.n199 585
R868 B.n198 B.n197 585
R869 B.n196 B.n195 585
R870 B.n194 B.n193 585
R871 B.n192 B.n191 585
R872 B.n190 B.n189 585
R873 B.n188 B.n187 585
R874 B.n186 B.n185 585
R875 B.n184 B.n183 585
R876 B.n182 B.n181 585
R877 B.n180 B.n179 585
R878 B.n178 B.n177 585
R879 B.n176 B.n175 585
R880 B.n174 B.n173 585
R881 B.n172 B.n171 585
R882 B.n170 B.n169 585
R883 B.n168 B.n167 585
R884 B.n166 B.n165 585
R885 B.n164 B.n163 585
R886 B.n162 B.n161 585
R887 B.n160 B.n159 585
R888 B.n158 B.n157 585
R889 B.n156 B.n155 585
R890 B.n154 B.n153 585
R891 B.n152 B.n151 585
R892 B.n150 B.n149 585
R893 B.n148 B.n147 585
R894 B.n146 B.n145 585
R895 B.n144 B.n143 585
R896 B.n142 B.n141 585
R897 B.n140 B.n139 585
R898 B.n138 B.n137 585
R899 B.n136 B.n135 585
R900 B.n134 B.n133 585
R901 B.n132 B.n131 585
R902 B.n130 B.n129 585
R903 B.n128 B.n127 585
R904 B.n126 B.n125 585
R905 B.n124 B.n123 585
R906 B.n122 B.n121 585
R907 B.n120 B.n119 585
R908 B.n118 B.n117 585
R909 B.n116 B.n115 585
R910 B.n53 B.n52 585
R911 B.n783 B.n54 585
R912 B.n787 B.n54 585
R913 B.n782 B.n781 585
R914 B.n781 B.n50 585
R915 B.n780 B.n49 585
R916 B.n793 B.n49 585
R917 B.n779 B.n48 585
R918 B.n794 B.n48 585
R919 B.n778 B.n47 585
R920 B.n795 B.n47 585
R921 B.n777 B.n776 585
R922 B.n776 B.n46 585
R923 B.n775 B.n42 585
R924 B.n801 B.n42 585
R925 B.n774 B.n41 585
R926 B.n802 B.n41 585
R927 B.n773 B.n40 585
R928 B.n803 B.n40 585
R929 B.n772 B.n771 585
R930 B.n771 B.n36 585
R931 B.n770 B.n35 585
R932 B.n809 B.n35 585
R933 B.n769 B.n34 585
R934 B.n810 B.n34 585
R935 B.n768 B.n33 585
R936 B.n811 B.n33 585
R937 B.n767 B.n766 585
R938 B.n766 B.n29 585
R939 B.n765 B.n28 585
R940 B.n817 B.n28 585
R941 B.n764 B.n27 585
R942 B.n818 B.n27 585
R943 B.n763 B.n26 585
R944 B.n819 B.n26 585
R945 B.n762 B.n761 585
R946 B.n761 B.n22 585
R947 B.n760 B.n21 585
R948 B.n825 B.n21 585
R949 B.n759 B.n20 585
R950 B.n826 B.n20 585
R951 B.n758 B.n19 585
R952 B.n827 B.n19 585
R953 B.n757 B.n756 585
R954 B.n756 B.n15 585
R955 B.n755 B.n14 585
R956 B.n833 B.n14 585
R957 B.n754 B.n13 585
R958 B.n834 B.n13 585
R959 B.n753 B.n12 585
R960 B.n835 B.n12 585
R961 B.n752 B.n751 585
R962 B.n751 B.n750 585
R963 B.n749 B.n748 585
R964 B.n749 B.n8 585
R965 B.n747 B.n7 585
R966 B.n842 B.n7 585
R967 B.n746 B.n6 585
R968 B.n843 B.n6 585
R969 B.n745 B.n5 585
R970 B.n844 B.n5 585
R971 B.n744 B.n743 585
R972 B.n743 B.n4 585
R973 B.n742 B.n329 585
R974 B.n742 B.n741 585
R975 B.n732 B.n330 585
R976 B.n331 B.n330 585
R977 B.n734 B.n733 585
R978 B.n735 B.n734 585
R979 B.n731 B.n336 585
R980 B.n336 B.n335 585
R981 B.n730 B.n729 585
R982 B.n729 B.n728 585
R983 B.n338 B.n337 585
R984 B.n339 B.n338 585
R985 B.n721 B.n720 585
R986 B.n722 B.n721 585
R987 B.n719 B.n343 585
R988 B.n347 B.n343 585
R989 B.n718 B.n717 585
R990 B.n717 B.n716 585
R991 B.n345 B.n344 585
R992 B.n346 B.n345 585
R993 B.n709 B.n708 585
R994 B.n710 B.n709 585
R995 B.n707 B.n352 585
R996 B.n352 B.n351 585
R997 B.n706 B.n705 585
R998 B.n705 B.n704 585
R999 B.n354 B.n353 585
R1000 B.n355 B.n354 585
R1001 B.n697 B.n696 585
R1002 B.n698 B.n697 585
R1003 B.n695 B.n360 585
R1004 B.n360 B.n359 585
R1005 B.n694 B.n693 585
R1006 B.n693 B.n692 585
R1007 B.n362 B.n361 585
R1008 B.n363 B.n362 585
R1009 B.n685 B.n684 585
R1010 B.n686 B.n685 585
R1011 B.n683 B.n368 585
R1012 B.n368 B.n367 585
R1013 B.n682 B.n681 585
R1014 B.n681 B.n680 585
R1015 B.n370 B.n369 585
R1016 B.n673 B.n370 585
R1017 B.n672 B.n671 585
R1018 B.n674 B.n672 585
R1019 B.n670 B.n375 585
R1020 B.n375 B.n374 585
R1021 B.n669 B.n668 585
R1022 B.n668 B.n667 585
R1023 B.n377 B.n376 585
R1024 B.n378 B.n377 585
R1025 B.n660 B.n659 585
R1026 B.n661 B.n660 585
R1027 B.n381 B.n380 585
R1028 B.n442 B.n440 585
R1029 B.n443 B.n439 585
R1030 B.n443 B.n382 585
R1031 B.n446 B.n445 585
R1032 B.n447 B.n438 585
R1033 B.n449 B.n448 585
R1034 B.n451 B.n437 585
R1035 B.n454 B.n453 585
R1036 B.n455 B.n436 585
R1037 B.n457 B.n456 585
R1038 B.n459 B.n435 585
R1039 B.n462 B.n461 585
R1040 B.n463 B.n434 585
R1041 B.n465 B.n464 585
R1042 B.n467 B.n433 585
R1043 B.n470 B.n469 585
R1044 B.n471 B.n432 585
R1045 B.n473 B.n472 585
R1046 B.n475 B.n431 585
R1047 B.n478 B.n477 585
R1048 B.n479 B.n430 585
R1049 B.n481 B.n480 585
R1050 B.n483 B.n429 585
R1051 B.n486 B.n485 585
R1052 B.n487 B.n428 585
R1053 B.n489 B.n488 585
R1054 B.n491 B.n427 585
R1055 B.n494 B.n493 585
R1056 B.n495 B.n426 585
R1057 B.n497 B.n496 585
R1058 B.n499 B.n425 585
R1059 B.n502 B.n501 585
R1060 B.n503 B.n424 585
R1061 B.n505 B.n504 585
R1062 B.n507 B.n423 585
R1063 B.n510 B.n509 585
R1064 B.n511 B.n422 585
R1065 B.n513 B.n512 585
R1066 B.n515 B.n421 585
R1067 B.n518 B.n517 585
R1068 B.n519 B.n420 585
R1069 B.n521 B.n520 585
R1070 B.n523 B.n419 585
R1071 B.n526 B.n525 585
R1072 B.n527 B.n418 585
R1073 B.n529 B.n528 585
R1074 B.n531 B.n417 585
R1075 B.n534 B.n533 585
R1076 B.n535 B.n416 585
R1077 B.n540 B.n539 585
R1078 B.n542 B.n415 585
R1079 B.n545 B.n544 585
R1080 B.n546 B.n414 585
R1081 B.n548 B.n547 585
R1082 B.n550 B.n413 585
R1083 B.n553 B.n552 585
R1084 B.n554 B.n412 585
R1085 B.n556 B.n555 585
R1086 B.n558 B.n411 585
R1087 B.n561 B.n560 585
R1088 B.n562 B.n407 585
R1089 B.n564 B.n563 585
R1090 B.n566 B.n406 585
R1091 B.n569 B.n568 585
R1092 B.n570 B.n405 585
R1093 B.n572 B.n571 585
R1094 B.n574 B.n404 585
R1095 B.n577 B.n576 585
R1096 B.n578 B.n403 585
R1097 B.n580 B.n579 585
R1098 B.n582 B.n402 585
R1099 B.n585 B.n584 585
R1100 B.n586 B.n401 585
R1101 B.n588 B.n587 585
R1102 B.n590 B.n400 585
R1103 B.n593 B.n592 585
R1104 B.n594 B.n399 585
R1105 B.n596 B.n595 585
R1106 B.n598 B.n398 585
R1107 B.n601 B.n600 585
R1108 B.n602 B.n397 585
R1109 B.n604 B.n603 585
R1110 B.n606 B.n396 585
R1111 B.n609 B.n608 585
R1112 B.n610 B.n395 585
R1113 B.n612 B.n611 585
R1114 B.n614 B.n394 585
R1115 B.n617 B.n616 585
R1116 B.n618 B.n393 585
R1117 B.n620 B.n619 585
R1118 B.n622 B.n392 585
R1119 B.n625 B.n624 585
R1120 B.n626 B.n391 585
R1121 B.n628 B.n627 585
R1122 B.n630 B.n390 585
R1123 B.n633 B.n632 585
R1124 B.n634 B.n389 585
R1125 B.n636 B.n635 585
R1126 B.n638 B.n388 585
R1127 B.n641 B.n640 585
R1128 B.n642 B.n387 585
R1129 B.n644 B.n643 585
R1130 B.n646 B.n386 585
R1131 B.n649 B.n648 585
R1132 B.n650 B.n385 585
R1133 B.n652 B.n651 585
R1134 B.n654 B.n384 585
R1135 B.n657 B.n656 585
R1136 B.n658 B.n383 585
R1137 B.n663 B.n662 585
R1138 B.n662 B.n661 585
R1139 B.n664 B.n379 585
R1140 B.n379 B.n378 585
R1141 B.n666 B.n665 585
R1142 B.n667 B.n666 585
R1143 B.n373 B.n372 585
R1144 B.n374 B.n373 585
R1145 B.n676 B.n675 585
R1146 B.n675 B.n674 585
R1147 B.n677 B.n371 585
R1148 B.n673 B.n371 585
R1149 B.n679 B.n678 585
R1150 B.n680 B.n679 585
R1151 B.n366 B.n365 585
R1152 B.n367 B.n366 585
R1153 B.n688 B.n687 585
R1154 B.n687 B.n686 585
R1155 B.n689 B.n364 585
R1156 B.n364 B.n363 585
R1157 B.n691 B.n690 585
R1158 B.n692 B.n691 585
R1159 B.n358 B.n357 585
R1160 B.n359 B.n358 585
R1161 B.n700 B.n699 585
R1162 B.n699 B.n698 585
R1163 B.n701 B.n356 585
R1164 B.n356 B.n355 585
R1165 B.n703 B.n702 585
R1166 B.n704 B.n703 585
R1167 B.n350 B.n349 585
R1168 B.n351 B.n350 585
R1169 B.n712 B.n711 585
R1170 B.n711 B.n710 585
R1171 B.n713 B.n348 585
R1172 B.n348 B.n346 585
R1173 B.n715 B.n714 585
R1174 B.n716 B.n715 585
R1175 B.n342 B.n341 585
R1176 B.n347 B.n342 585
R1177 B.n724 B.n723 585
R1178 B.n723 B.n722 585
R1179 B.n725 B.n340 585
R1180 B.n340 B.n339 585
R1181 B.n727 B.n726 585
R1182 B.n728 B.n727 585
R1183 B.n334 B.n333 585
R1184 B.n335 B.n334 585
R1185 B.n737 B.n736 585
R1186 B.n736 B.n735 585
R1187 B.n738 B.n332 585
R1188 B.n332 B.n331 585
R1189 B.n740 B.n739 585
R1190 B.n741 B.n740 585
R1191 B.n3 B.n0 585
R1192 B.n4 B.n3 585
R1193 B.n841 B.n1 585
R1194 B.n842 B.n841 585
R1195 B.n840 B.n839 585
R1196 B.n840 B.n8 585
R1197 B.n838 B.n9 585
R1198 B.n750 B.n9 585
R1199 B.n837 B.n836 585
R1200 B.n836 B.n835 585
R1201 B.n11 B.n10 585
R1202 B.n834 B.n11 585
R1203 B.n832 B.n831 585
R1204 B.n833 B.n832 585
R1205 B.n830 B.n16 585
R1206 B.n16 B.n15 585
R1207 B.n829 B.n828 585
R1208 B.n828 B.n827 585
R1209 B.n18 B.n17 585
R1210 B.n826 B.n18 585
R1211 B.n824 B.n823 585
R1212 B.n825 B.n824 585
R1213 B.n822 B.n23 585
R1214 B.n23 B.n22 585
R1215 B.n821 B.n820 585
R1216 B.n820 B.n819 585
R1217 B.n25 B.n24 585
R1218 B.n818 B.n25 585
R1219 B.n816 B.n815 585
R1220 B.n817 B.n816 585
R1221 B.n814 B.n30 585
R1222 B.n30 B.n29 585
R1223 B.n813 B.n812 585
R1224 B.n812 B.n811 585
R1225 B.n32 B.n31 585
R1226 B.n810 B.n32 585
R1227 B.n808 B.n807 585
R1228 B.n809 B.n808 585
R1229 B.n806 B.n37 585
R1230 B.n37 B.n36 585
R1231 B.n805 B.n804 585
R1232 B.n804 B.n803 585
R1233 B.n39 B.n38 585
R1234 B.n802 B.n39 585
R1235 B.n800 B.n799 585
R1236 B.n801 B.n800 585
R1237 B.n798 B.n43 585
R1238 B.n46 B.n43 585
R1239 B.n797 B.n796 585
R1240 B.n796 B.n795 585
R1241 B.n45 B.n44 585
R1242 B.n794 B.n45 585
R1243 B.n792 B.n791 585
R1244 B.n793 B.n792 585
R1245 B.n790 B.n51 585
R1246 B.n51 B.n50 585
R1247 B.n789 B.n788 585
R1248 B.n788 B.n787 585
R1249 B.n845 B.n844 585
R1250 B.n843 B.n2 585
R1251 B.n788 B.n53 530.939
R1252 B.n785 B.n54 530.939
R1253 B.n660 B.n383 530.939
R1254 B.n662 B.n381 530.939
R1255 B.n112 B.t6 457.882
R1256 B.n110 B.t14 457.882
R1257 B.n408 B.t10 457.882
R1258 B.n536 B.t17 457.882
R1259 B.n112 B.t8 363.961
R1260 B.n110 B.t15 363.961
R1261 B.n408 B.t13 363.961
R1262 B.n536 B.t19 363.961
R1263 B.n111 B.t16 330.216
R1264 B.n409 B.t12 330.216
R1265 B.n113 B.t9 330.216
R1266 B.n537 B.t18 330.216
R1267 B.n786 B.n108 256.663
R1268 B.n786 B.n107 256.663
R1269 B.n786 B.n106 256.663
R1270 B.n786 B.n105 256.663
R1271 B.n786 B.n104 256.663
R1272 B.n786 B.n103 256.663
R1273 B.n786 B.n102 256.663
R1274 B.n786 B.n101 256.663
R1275 B.n786 B.n100 256.663
R1276 B.n786 B.n99 256.663
R1277 B.n786 B.n98 256.663
R1278 B.n786 B.n97 256.663
R1279 B.n786 B.n96 256.663
R1280 B.n786 B.n95 256.663
R1281 B.n786 B.n94 256.663
R1282 B.n786 B.n93 256.663
R1283 B.n786 B.n92 256.663
R1284 B.n786 B.n91 256.663
R1285 B.n786 B.n90 256.663
R1286 B.n786 B.n89 256.663
R1287 B.n786 B.n88 256.663
R1288 B.n786 B.n87 256.663
R1289 B.n786 B.n86 256.663
R1290 B.n786 B.n85 256.663
R1291 B.n786 B.n84 256.663
R1292 B.n786 B.n83 256.663
R1293 B.n786 B.n82 256.663
R1294 B.n786 B.n81 256.663
R1295 B.n786 B.n80 256.663
R1296 B.n786 B.n79 256.663
R1297 B.n786 B.n78 256.663
R1298 B.n786 B.n77 256.663
R1299 B.n786 B.n76 256.663
R1300 B.n786 B.n75 256.663
R1301 B.n786 B.n74 256.663
R1302 B.n786 B.n73 256.663
R1303 B.n786 B.n72 256.663
R1304 B.n786 B.n71 256.663
R1305 B.n786 B.n70 256.663
R1306 B.n786 B.n69 256.663
R1307 B.n786 B.n68 256.663
R1308 B.n786 B.n67 256.663
R1309 B.n786 B.n66 256.663
R1310 B.n786 B.n65 256.663
R1311 B.n786 B.n64 256.663
R1312 B.n786 B.n63 256.663
R1313 B.n786 B.n62 256.663
R1314 B.n786 B.n61 256.663
R1315 B.n786 B.n60 256.663
R1316 B.n786 B.n59 256.663
R1317 B.n786 B.n58 256.663
R1318 B.n786 B.n57 256.663
R1319 B.n786 B.n56 256.663
R1320 B.n786 B.n55 256.663
R1321 B.n441 B.n382 256.663
R1322 B.n444 B.n382 256.663
R1323 B.n450 B.n382 256.663
R1324 B.n452 B.n382 256.663
R1325 B.n458 B.n382 256.663
R1326 B.n460 B.n382 256.663
R1327 B.n466 B.n382 256.663
R1328 B.n468 B.n382 256.663
R1329 B.n474 B.n382 256.663
R1330 B.n476 B.n382 256.663
R1331 B.n482 B.n382 256.663
R1332 B.n484 B.n382 256.663
R1333 B.n490 B.n382 256.663
R1334 B.n492 B.n382 256.663
R1335 B.n498 B.n382 256.663
R1336 B.n500 B.n382 256.663
R1337 B.n506 B.n382 256.663
R1338 B.n508 B.n382 256.663
R1339 B.n514 B.n382 256.663
R1340 B.n516 B.n382 256.663
R1341 B.n522 B.n382 256.663
R1342 B.n524 B.n382 256.663
R1343 B.n530 B.n382 256.663
R1344 B.n532 B.n382 256.663
R1345 B.n541 B.n382 256.663
R1346 B.n543 B.n382 256.663
R1347 B.n549 B.n382 256.663
R1348 B.n551 B.n382 256.663
R1349 B.n557 B.n382 256.663
R1350 B.n559 B.n382 256.663
R1351 B.n565 B.n382 256.663
R1352 B.n567 B.n382 256.663
R1353 B.n573 B.n382 256.663
R1354 B.n575 B.n382 256.663
R1355 B.n581 B.n382 256.663
R1356 B.n583 B.n382 256.663
R1357 B.n589 B.n382 256.663
R1358 B.n591 B.n382 256.663
R1359 B.n597 B.n382 256.663
R1360 B.n599 B.n382 256.663
R1361 B.n605 B.n382 256.663
R1362 B.n607 B.n382 256.663
R1363 B.n613 B.n382 256.663
R1364 B.n615 B.n382 256.663
R1365 B.n621 B.n382 256.663
R1366 B.n623 B.n382 256.663
R1367 B.n629 B.n382 256.663
R1368 B.n631 B.n382 256.663
R1369 B.n637 B.n382 256.663
R1370 B.n639 B.n382 256.663
R1371 B.n645 B.n382 256.663
R1372 B.n647 B.n382 256.663
R1373 B.n653 B.n382 256.663
R1374 B.n655 B.n382 256.663
R1375 B.n847 B.n846 256.663
R1376 B.n117 B.n116 163.367
R1377 B.n121 B.n120 163.367
R1378 B.n125 B.n124 163.367
R1379 B.n129 B.n128 163.367
R1380 B.n133 B.n132 163.367
R1381 B.n137 B.n136 163.367
R1382 B.n141 B.n140 163.367
R1383 B.n145 B.n144 163.367
R1384 B.n149 B.n148 163.367
R1385 B.n153 B.n152 163.367
R1386 B.n157 B.n156 163.367
R1387 B.n161 B.n160 163.367
R1388 B.n165 B.n164 163.367
R1389 B.n169 B.n168 163.367
R1390 B.n173 B.n172 163.367
R1391 B.n177 B.n176 163.367
R1392 B.n181 B.n180 163.367
R1393 B.n185 B.n184 163.367
R1394 B.n189 B.n188 163.367
R1395 B.n193 B.n192 163.367
R1396 B.n197 B.n196 163.367
R1397 B.n201 B.n200 163.367
R1398 B.n205 B.n204 163.367
R1399 B.n209 B.n208 163.367
R1400 B.n213 B.n212 163.367
R1401 B.n217 B.n216 163.367
R1402 B.n221 B.n220 163.367
R1403 B.n225 B.n224 163.367
R1404 B.n229 B.n228 163.367
R1405 B.n234 B.n233 163.367
R1406 B.n238 B.n237 163.367
R1407 B.n242 B.n241 163.367
R1408 B.n246 B.n245 163.367
R1409 B.n250 B.n249 163.367
R1410 B.n254 B.n253 163.367
R1411 B.n258 B.n257 163.367
R1412 B.n262 B.n261 163.367
R1413 B.n266 B.n265 163.367
R1414 B.n270 B.n269 163.367
R1415 B.n274 B.n273 163.367
R1416 B.n278 B.n277 163.367
R1417 B.n282 B.n281 163.367
R1418 B.n286 B.n285 163.367
R1419 B.n290 B.n289 163.367
R1420 B.n294 B.n293 163.367
R1421 B.n298 B.n297 163.367
R1422 B.n302 B.n301 163.367
R1423 B.n306 B.n305 163.367
R1424 B.n310 B.n309 163.367
R1425 B.n314 B.n313 163.367
R1426 B.n318 B.n317 163.367
R1427 B.n322 B.n321 163.367
R1428 B.n326 B.n325 163.367
R1429 B.n785 B.n109 163.367
R1430 B.n660 B.n377 163.367
R1431 B.n668 B.n377 163.367
R1432 B.n668 B.n375 163.367
R1433 B.n672 B.n375 163.367
R1434 B.n672 B.n370 163.367
R1435 B.n681 B.n370 163.367
R1436 B.n681 B.n368 163.367
R1437 B.n685 B.n368 163.367
R1438 B.n685 B.n362 163.367
R1439 B.n693 B.n362 163.367
R1440 B.n693 B.n360 163.367
R1441 B.n697 B.n360 163.367
R1442 B.n697 B.n354 163.367
R1443 B.n705 B.n354 163.367
R1444 B.n705 B.n352 163.367
R1445 B.n709 B.n352 163.367
R1446 B.n709 B.n345 163.367
R1447 B.n717 B.n345 163.367
R1448 B.n717 B.n343 163.367
R1449 B.n721 B.n343 163.367
R1450 B.n721 B.n338 163.367
R1451 B.n729 B.n338 163.367
R1452 B.n729 B.n336 163.367
R1453 B.n734 B.n336 163.367
R1454 B.n734 B.n330 163.367
R1455 B.n742 B.n330 163.367
R1456 B.n743 B.n742 163.367
R1457 B.n743 B.n5 163.367
R1458 B.n6 B.n5 163.367
R1459 B.n7 B.n6 163.367
R1460 B.n749 B.n7 163.367
R1461 B.n751 B.n749 163.367
R1462 B.n751 B.n12 163.367
R1463 B.n13 B.n12 163.367
R1464 B.n14 B.n13 163.367
R1465 B.n756 B.n14 163.367
R1466 B.n756 B.n19 163.367
R1467 B.n20 B.n19 163.367
R1468 B.n21 B.n20 163.367
R1469 B.n761 B.n21 163.367
R1470 B.n761 B.n26 163.367
R1471 B.n27 B.n26 163.367
R1472 B.n28 B.n27 163.367
R1473 B.n766 B.n28 163.367
R1474 B.n766 B.n33 163.367
R1475 B.n34 B.n33 163.367
R1476 B.n35 B.n34 163.367
R1477 B.n771 B.n35 163.367
R1478 B.n771 B.n40 163.367
R1479 B.n41 B.n40 163.367
R1480 B.n42 B.n41 163.367
R1481 B.n776 B.n42 163.367
R1482 B.n776 B.n47 163.367
R1483 B.n48 B.n47 163.367
R1484 B.n49 B.n48 163.367
R1485 B.n781 B.n49 163.367
R1486 B.n781 B.n54 163.367
R1487 B.n443 B.n442 163.367
R1488 B.n445 B.n443 163.367
R1489 B.n449 B.n438 163.367
R1490 B.n453 B.n451 163.367
R1491 B.n457 B.n436 163.367
R1492 B.n461 B.n459 163.367
R1493 B.n465 B.n434 163.367
R1494 B.n469 B.n467 163.367
R1495 B.n473 B.n432 163.367
R1496 B.n477 B.n475 163.367
R1497 B.n481 B.n430 163.367
R1498 B.n485 B.n483 163.367
R1499 B.n489 B.n428 163.367
R1500 B.n493 B.n491 163.367
R1501 B.n497 B.n426 163.367
R1502 B.n501 B.n499 163.367
R1503 B.n505 B.n424 163.367
R1504 B.n509 B.n507 163.367
R1505 B.n513 B.n422 163.367
R1506 B.n517 B.n515 163.367
R1507 B.n521 B.n420 163.367
R1508 B.n525 B.n523 163.367
R1509 B.n529 B.n418 163.367
R1510 B.n533 B.n531 163.367
R1511 B.n540 B.n416 163.367
R1512 B.n544 B.n542 163.367
R1513 B.n548 B.n414 163.367
R1514 B.n552 B.n550 163.367
R1515 B.n556 B.n412 163.367
R1516 B.n560 B.n558 163.367
R1517 B.n564 B.n407 163.367
R1518 B.n568 B.n566 163.367
R1519 B.n572 B.n405 163.367
R1520 B.n576 B.n574 163.367
R1521 B.n580 B.n403 163.367
R1522 B.n584 B.n582 163.367
R1523 B.n588 B.n401 163.367
R1524 B.n592 B.n590 163.367
R1525 B.n596 B.n399 163.367
R1526 B.n600 B.n598 163.367
R1527 B.n604 B.n397 163.367
R1528 B.n608 B.n606 163.367
R1529 B.n612 B.n395 163.367
R1530 B.n616 B.n614 163.367
R1531 B.n620 B.n393 163.367
R1532 B.n624 B.n622 163.367
R1533 B.n628 B.n391 163.367
R1534 B.n632 B.n630 163.367
R1535 B.n636 B.n389 163.367
R1536 B.n640 B.n638 163.367
R1537 B.n644 B.n387 163.367
R1538 B.n648 B.n646 163.367
R1539 B.n652 B.n385 163.367
R1540 B.n656 B.n654 163.367
R1541 B.n662 B.n379 163.367
R1542 B.n666 B.n379 163.367
R1543 B.n666 B.n373 163.367
R1544 B.n675 B.n373 163.367
R1545 B.n675 B.n371 163.367
R1546 B.n679 B.n371 163.367
R1547 B.n679 B.n366 163.367
R1548 B.n687 B.n366 163.367
R1549 B.n687 B.n364 163.367
R1550 B.n691 B.n364 163.367
R1551 B.n691 B.n358 163.367
R1552 B.n699 B.n358 163.367
R1553 B.n699 B.n356 163.367
R1554 B.n703 B.n356 163.367
R1555 B.n703 B.n350 163.367
R1556 B.n711 B.n350 163.367
R1557 B.n711 B.n348 163.367
R1558 B.n715 B.n348 163.367
R1559 B.n715 B.n342 163.367
R1560 B.n723 B.n342 163.367
R1561 B.n723 B.n340 163.367
R1562 B.n727 B.n340 163.367
R1563 B.n727 B.n334 163.367
R1564 B.n736 B.n334 163.367
R1565 B.n736 B.n332 163.367
R1566 B.n740 B.n332 163.367
R1567 B.n740 B.n3 163.367
R1568 B.n845 B.n3 163.367
R1569 B.n841 B.n2 163.367
R1570 B.n841 B.n840 163.367
R1571 B.n840 B.n9 163.367
R1572 B.n836 B.n9 163.367
R1573 B.n836 B.n11 163.367
R1574 B.n832 B.n11 163.367
R1575 B.n832 B.n16 163.367
R1576 B.n828 B.n16 163.367
R1577 B.n828 B.n18 163.367
R1578 B.n824 B.n18 163.367
R1579 B.n824 B.n23 163.367
R1580 B.n820 B.n23 163.367
R1581 B.n820 B.n25 163.367
R1582 B.n816 B.n25 163.367
R1583 B.n816 B.n30 163.367
R1584 B.n812 B.n30 163.367
R1585 B.n812 B.n32 163.367
R1586 B.n808 B.n32 163.367
R1587 B.n808 B.n37 163.367
R1588 B.n804 B.n37 163.367
R1589 B.n804 B.n39 163.367
R1590 B.n800 B.n39 163.367
R1591 B.n800 B.n43 163.367
R1592 B.n796 B.n43 163.367
R1593 B.n796 B.n45 163.367
R1594 B.n792 B.n45 163.367
R1595 B.n792 B.n51 163.367
R1596 B.n788 B.n51 163.367
R1597 B.n55 B.n53 71.676
R1598 B.n117 B.n56 71.676
R1599 B.n121 B.n57 71.676
R1600 B.n125 B.n58 71.676
R1601 B.n129 B.n59 71.676
R1602 B.n133 B.n60 71.676
R1603 B.n137 B.n61 71.676
R1604 B.n141 B.n62 71.676
R1605 B.n145 B.n63 71.676
R1606 B.n149 B.n64 71.676
R1607 B.n153 B.n65 71.676
R1608 B.n157 B.n66 71.676
R1609 B.n161 B.n67 71.676
R1610 B.n165 B.n68 71.676
R1611 B.n169 B.n69 71.676
R1612 B.n173 B.n70 71.676
R1613 B.n177 B.n71 71.676
R1614 B.n181 B.n72 71.676
R1615 B.n185 B.n73 71.676
R1616 B.n189 B.n74 71.676
R1617 B.n193 B.n75 71.676
R1618 B.n197 B.n76 71.676
R1619 B.n201 B.n77 71.676
R1620 B.n205 B.n78 71.676
R1621 B.n209 B.n79 71.676
R1622 B.n213 B.n80 71.676
R1623 B.n217 B.n81 71.676
R1624 B.n221 B.n82 71.676
R1625 B.n225 B.n83 71.676
R1626 B.n229 B.n84 71.676
R1627 B.n234 B.n85 71.676
R1628 B.n238 B.n86 71.676
R1629 B.n242 B.n87 71.676
R1630 B.n246 B.n88 71.676
R1631 B.n250 B.n89 71.676
R1632 B.n254 B.n90 71.676
R1633 B.n258 B.n91 71.676
R1634 B.n262 B.n92 71.676
R1635 B.n266 B.n93 71.676
R1636 B.n270 B.n94 71.676
R1637 B.n274 B.n95 71.676
R1638 B.n278 B.n96 71.676
R1639 B.n282 B.n97 71.676
R1640 B.n286 B.n98 71.676
R1641 B.n290 B.n99 71.676
R1642 B.n294 B.n100 71.676
R1643 B.n298 B.n101 71.676
R1644 B.n302 B.n102 71.676
R1645 B.n306 B.n103 71.676
R1646 B.n310 B.n104 71.676
R1647 B.n314 B.n105 71.676
R1648 B.n318 B.n106 71.676
R1649 B.n322 B.n107 71.676
R1650 B.n326 B.n108 71.676
R1651 B.n109 B.n108 71.676
R1652 B.n325 B.n107 71.676
R1653 B.n321 B.n106 71.676
R1654 B.n317 B.n105 71.676
R1655 B.n313 B.n104 71.676
R1656 B.n309 B.n103 71.676
R1657 B.n305 B.n102 71.676
R1658 B.n301 B.n101 71.676
R1659 B.n297 B.n100 71.676
R1660 B.n293 B.n99 71.676
R1661 B.n289 B.n98 71.676
R1662 B.n285 B.n97 71.676
R1663 B.n281 B.n96 71.676
R1664 B.n277 B.n95 71.676
R1665 B.n273 B.n94 71.676
R1666 B.n269 B.n93 71.676
R1667 B.n265 B.n92 71.676
R1668 B.n261 B.n91 71.676
R1669 B.n257 B.n90 71.676
R1670 B.n253 B.n89 71.676
R1671 B.n249 B.n88 71.676
R1672 B.n245 B.n87 71.676
R1673 B.n241 B.n86 71.676
R1674 B.n237 B.n85 71.676
R1675 B.n233 B.n84 71.676
R1676 B.n228 B.n83 71.676
R1677 B.n224 B.n82 71.676
R1678 B.n220 B.n81 71.676
R1679 B.n216 B.n80 71.676
R1680 B.n212 B.n79 71.676
R1681 B.n208 B.n78 71.676
R1682 B.n204 B.n77 71.676
R1683 B.n200 B.n76 71.676
R1684 B.n196 B.n75 71.676
R1685 B.n192 B.n74 71.676
R1686 B.n188 B.n73 71.676
R1687 B.n184 B.n72 71.676
R1688 B.n180 B.n71 71.676
R1689 B.n176 B.n70 71.676
R1690 B.n172 B.n69 71.676
R1691 B.n168 B.n68 71.676
R1692 B.n164 B.n67 71.676
R1693 B.n160 B.n66 71.676
R1694 B.n156 B.n65 71.676
R1695 B.n152 B.n64 71.676
R1696 B.n148 B.n63 71.676
R1697 B.n144 B.n62 71.676
R1698 B.n140 B.n61 71.676
R1699 B.n136 B.n60 71.676
R1700 B.n132 B.n59 71.676
R1701 B.n128 B.n58 71.676
R1702 B.n124 B.n57 71.676
R1703 B.n120 B.n56 71.676
R1704 B.n116 B.n55 71.676
R1705 B.n441 B.n381 71.676
R1706 B.n445 B.n444 71.676
R1707 B.n450 B.n449 71.676
R1708 B.n453 B.n452 71.676
R1709 B.n458 B.n457 71.676
R1710 B.n461 B.n460 71.676
R1711 B.n466 B.n465 71.676
R1712 B.n469 B.n468 71.676
R1713 B.n474 B.n473 71.676
R1714 B.n477 B.n476 71.676
R1715 B.n482 B.n481 71.676
R1716 B.n485 B.n484 71.676
R1717 B.n490 B.n489 71.676
R1718 B.n493 B.n492 71.676
R1719 B.n498 B.n497 71.676
R1720 B.n501 B.n500 71.676
R1721 B.n506 B.n505 71.676
R1722 B.n509 B.n508 71.676
R1723 B.n514 B.n513 71.676
R1724 B.n517 B.n516 71.676
R1725 B.n522 B.n521 71.676
R1726 B.n525 B.n524 71.676
R1727 B.n530 B.n529 71.676
R1728 B.n533 B.n532 71.676
R1729 B.n541 B.n540 71.676
R1730 B.n544 B.n543 71.676
R1731 B.n549 B.n548 71.676
R1732 B.n552 B.n551 71.676
R1733 B.n557 B.n556 71.676
R1734 B.n560 B.n559 71.676
R1735 B.n565 B.n564 71.676
R1736 B.n568 B.n567 71.676
R1737 B.n573 B.n572 71.676
R1738 B.n576 B.n575 71.676
R1739 B.n581 B.n580 71.676
R1740 B.n584 B.n583 71.676
R1741 B.n589 B.n588 71.676
R1742 B.n592 B.n591 71.676
R1743 B.n597 B.n596 71.676
R1744 B.n600 B.n599 71.676
R1745 B.n605 B.n604 71.676
R1746 B.n608 B.n607 71.676
R1747 B.n613 B.n612 71.676
R1748 B.n616 B.n615 71.676
R1749 B.n621 B.n620 71.676
R1750 B.n624 B.n623 71.676
R1751 B.n629 B.n628 71.676
R1752 B.n632 B.n631 71.676
R1753 B.n637 B.n636 71.676
R1754 B.n640 B.n639 71.676
R1755 B.n645 B.n644 71.676
R1756 B.n648 B.n647 71.676
R1757 B.n653 B.n652 71.676
R1758 B.n656 B.n655 71.676
R1759 B.n442 B.n441 71.676
R1760 B.n444 B.n438 71.676
R1761 B.n451 B.n450 71.676
R1762 B.n452 B.n436 71.676
R1763 B.n459 B.n458 71.676
R1764 B.n460 B.n434 71.676
R1765 B.n467 B.n466 71.676
R1766 B.n468 B.n432 71.676
R1767 B.n475 B.n474 71.676
R1768 B.n476 B.n430 71.676
R1769 B.n483 B.n482 71.676
R1770 B.n484 B.n428 71.676
R1771 B.n491 B.n490 71.676
R1772 B.n492 B.n426 71.676
R1773 B.n499 B.n498 71.676
R1774 B.n500 B.n424 71.676
R1775 B.n507 B.n506 71.676
R1776 B.n508 B.n422 71.676
R1777 B.n515 B.n514 71.676
R1778 B.n516 B.n420 71.676
R1779 B.n523 B.n522 71.676
R1780 B.n524 B.n418 71.676
R1781 B.n531 B.n530 71.676
R1782 B.n532 B.n416 71.676
R1783 B.n542 B.n541 71.676
R1784 B.n543 B.n414 71.676
R1785 B.n550 B.n549 71.676
R1786 B.n551 B.n412 71.676
R1787 B.n558 B.n557 71.676
R1788 B.n559 B.n407 71.676
R1789 B.n566 B.n565 71.676
R1790 B.n567 B.n405 71.676
R1791 B.n574 B.n573 71.676
R1792 B.n575 B.n403 71.676
R1793 B.n582 B.n581 71.676
R1794 B.n583 B.n401 71.676
R1795 B.n590 B.n589 71.676
R1796 B.n591 B.n399 71.676
R1797 B.n598 B.n597 71.676
R1798 B.n599 B.n397 71.676
R1799 B.n606 B.n605 71.676
R1800 B.n607 B.n395 71.676
R1801 B.n614 B.n613 71.676
R1802 B.n615 B.n393 71.676
R1803 B.n622 B.n621 71.676
R1804 B.n623 B.n391 71.676
R1805 B.n630 B.n629 71.676
R1806 B.n631 B.n389 71.676
R1807 B.n638 B.n637 71.676
R1808 B.n639 B.n387 71.676
R1809 B.n646 B.n645 71.676
R1810 B.n647 B.n385 71.676
R1811 B.n654 B.n653 71.676
R1812 B.n655 B.n383 71.676
R1813 B.n846 B.n845 71.676
R1814 B.n846 B.n2 71.676
R1815 B.n661 B.n382 70.7207
R1816 B.n787 B.n786 70.7207
R1817 B.n114 B.n113 59.5399
R1818 B.n231 B.n111 59.5399
R1819 B.n410 B.n409 59.5399
R1820 B.n538 B.n537 59.5399
R1821 B.n661 B.n378 37.2793
R1822 B.n667 B.n378 37.2793
R1823 B.n667 B.n374 37.2793
R1824 B.n674 B.n374 37.2793
R1825 B.n674 B.n673 37.2793
R1826 B.n680 B.n367 37.2793
R1827 B.n686 B.n367 37.2793
R1828 B.n686 B.n363 37.2793
R1829 B.n692 B.n363 37.2793
R1830 B.n692 B.n359 37.2793
R1831 B.n698 B.n359 37.2793
R1832 B.n698 B.n355 37.2793
R1833 B.n704 B.n355 37.2793
R1834 B.n710 B.n351 37.2793
R1835 B.n710 B.n346 37.2793
R1836 B.n716 B.n346 37.2793
R1837 B.n716 B.n347 37.2793
R1838 B.n722 B.n339 37.2793
R1839 B.n728 B.n339 37.2793
R1840 B.n728 B.n335 37.2793
R1841 B.n735 B.n335 37.2793
R1842 B.n741 B.n331 37.2793
R1843 B.n741 B.n4 37.2793
R1844 B.n844 B.n4 37.2793
R1845 B.n844 B.n843 37.2793
R1846 B.n843 B.n842 37.2793
R1847 B.n842 B.n8 37.2793
R1848 B.n750 B.n8 37.2793
R1849 B.n835 B.n834 37.2793
R1850 B.n834 B.n833 37.2793
R1851 B.n833 B.n15 37.2793
R1852 B.n827 B.n15 37.2793
R1853 B.n826 B.n825 37.2793
R1854 B.n825 B.n22 37.2793
R1855 B.n819 B.n22 37.2793
R1856 B.n819 B.n818 37.2793
R1857 B.n817 B.n29 37.2793
R1858 B.n811 B.n29 37.2793
R1859 B.n811 B.n810 37.2793
R1860 B.n810 B.n809 37.2793
R1861 B.n809 B.n36 37.2793
R1862 B.n803 B.n36 37.2793
R1863 B.n803 B.n802 37.2793
R1864 B.n802 B.n801 37.2793
R1865 B.n795 B.n46 37.2793
R1866 B.n795 B.n794 37.2793
R1867 B.n794 B.n793 37.2793
R1868 B.n793 B.n50 37.2793
R1869 B.n787 B.n50 37.2793
R1870 B.n663 B.n380 34.4981
R1871 B.n659 B.n658 34.4981
R1872 B.n784 B.n783 34.4981
R1873 B.n789 B.n52 34.4981
R1874 B.n113 B.n112 33.746
R1875 B.n111 B.n110 33.746
R1876 B.n409 B.n408 33.746
R1877 B.n537 B.n536 33.746
R1878 B.t3 B.n351 33.4418
R1879 B.n818 B.t4 33.4418
R1880 B.n673 B.t11 29.0561
R1881 B.n722 B.t5 29.0561
R1882 B.n827 B.t1 29.0561
R1883 B.n46 B.t7 29.0561
R1884 B.t2 B.n331 24.6703
R1885 B.n750 B.t0 24.6703
R1886 B B.n847 18.0485
R1887 B.n735 B.t2 12.6095
R1888 B.n835 B.t0 12.6095
R1889 B.n664 B.n663 10.6151
R1890 B.n665 B.n664 10.6151
R1891 B.n665 B.n372 10.6151
R1892 B.n676 B.n372 10.6151
R1893 B.n677 B.n676 10.6151
R1894 B.n678 B.n677 10.6151
R1895 B.n678 B.n365 10.6151
R1896 B.n688 B.n365 10.6151
R1897 B.n689 B.n688 10.6151
R1898 B.n690 B.n689 10.6151
R1899 B.n690 B.n357 10.6151
R1900 B.n700 B.n357 10.6151
R1901 B.n701 B.n700 10.6151
R1902 B.n702 B.n701 10.6151
R1903 B.n702 B.n349 10.6151
R1904 B.n712 B.n349 10.6151
R1905 B.n713 B.n712 10.6151
R1906 B.n714 B.n713 10.6151
R1907 B.n714 B.n341 10.6151
R1908 B.n724 B.n341 10.6151
R1909 B.n725 B.n724 10.6151
R1910 B.n726 B.n725 10.6151
R1911 B.n726 B.n333 10.6151
R1912 B.n737 B.n333 10.6151
R1913 B.n738 B.n737 10.6151
R1914 B.n739 B.n738 10.6151
R1915 B.n739 B.n0 10.6151
R1916 B.n440 B.n380 10.6151
R1917 B.n440 B.n439 10.6151
R1918 B.n446 B.n439 10.6151
R1919 B.n447 B.n446 10.6151
R1920 B.n448 B.n447 10.6151
R1921 B.n448 B.n437 10.6151
R1922 B.n454 B.n437 10.6151
R1923 B.n455 B.n454 10.6151
R1924 B.n456 B.n455 10.6151
R1925 B.n456 B.n435 10.6151
R1926 B.n462 B.n435 10.6151
R1927 B.n463 B.n462 10.6151
R1928 B.n464 B.n463 10.6151
R1929 B.n464 B.n433 10.6151
R1930 B.n470 B.n433 10.6151
R1931 B.n471 B.n470 10.6151
R1932 B.n472 B.n471 10.6151
R1933 B.n472 B.n431 10.6151
R1934 B.n478 B.n431 10.6151
R1935 B.n479 B.n478 10.6151
R1936 B.n480 B.n479 10.6151
R1937 B.n480 B.n429 10.6151
R1938 B.n486 B.n429 10.6151
R1939 B.n487 B.n486 10.6151
R1940 B.n488 B.n487 10.6151
R1941 B.n488 B.n427 10.6151
R1942 B.n494 B.n427 10.6151
R1943 B.n495 B.n494 10.6151
R1944 B.n496 B.n495 10.6151
R1945 B.n496 B.n425 10.6151
R1946 B.n502 B.n425 10.6151
R1947 B.n503 B.n502 10.6151
R1948 B.n504 B.n503 10.6151
R1949 B.n504 B.n423 10.6151
R1950 B.n510 B.n423 10.6151
R1951 B.n511 B.n510 10.6151
R1952 B.n512 B.n511 10.6151
R1953 B.n512 B.n421 10.6151
R1954 B.n518 B.n421 10.6151
R1955 B.n519 B.n518 10.6151
R1956 B.n520 B.n519 10.6151
R1957 B.n520 B.n419 10.6151
R1958 B.n526 B.n419 10.6151
R1959 B.n527 B.n526 10.6151
R1960 B.n528 B.n527 10.6151
R1961 B.n528 B.n417 10.6151
R1962 B.n534 B.n417 10.6151
R1963 B.n535 B.n534 10.6151
R1964 B.n539 B.n535 10.6151
R1965 B.n545 B.n415 10.6151
R1966 B.n546 B.n545 10.6151
R1967 B.n547 B.n546 10.6151
R1968 B.n547 B.n413 10.6151
R1969 B.n553 B.n413 10.6151
R1970 B.n554 B.n553 10.6151
R1971 B.n555 B.n554 10.6151
R1972 B.n555 B.n411 10.6151
R1973 B.n562 B.n561 10.6151
R1974 B.n563 B.n562 10.6151
R1975 B.n563 B.n406 10.6151
R1976 B.n569 B.n406 10.6151
R1977 B.n570 B.n569 10.6151
R1978 B.n571 B.n570 10.6151
R1979 B.n571 B.n404 10.6151
R1980 B.n577 B.n404 10.6151
R1981 B.n578 B.n577 10.6151
R1982 B.n579 B.n578 10.6151
R1983 B.n579 B.n402 10.6151
R1984 B.n585 B.n402 10.6151
R1985 B.n586 B.n585 10.6151
R1986 B.n587 B.n586 10.6151
R1987 B.n587 B.n400 10.6151
R1988 B.n593 B.n400 10.6151
R1989 B.n594 B.n593 10.6151
R1990 B.n595 B.n594 10.6151
R1991 B.n595 B.n398 10.6151
R1992 B.n601 B.n398 10.6151
R1993 B.n602 B.n601 10.6151
R1994 B.n603 B.n602 10.6151
R1995 B.n603 B.n396 10.6151
R1996 B.n609 B.n396 10.6151
R1997 B.n610 B.n609 10.6151
R1998 B.n611 B.n610 10.6151
R1999 B.n611 B.n394 10.6151
R2000 B.n617 B.n394 10.6151
R2001 B.n618 B.n617 10.6151
R2002 B.n619 B.n618 10.6151
R2003 B.n619 B.n392 10.6151
R2004 B.n625 B.n392 10.6151
R2005 B.n626 B.n625 10.6151
R2006 B.n627 B.n626 10.6151
R2007 B.n627 B.n390 10.6151
R2008 B.n633 B.n390 10.6151
R2009 B.n634 B.n633 10.6151
R2010 B.n635 B.n634 10.6151
R2011 B.n635 B.n388 10.6151
R2012 B.n641 B.n388 10.6151
R2013 B.n642 B.n641 10.6151
R2014 B.n643 B.n642 10.6151
R2015 B.n643 B.n386 10.6151
R2016 B.n649 B.n386 10.6151
R2017 B.n650 B.n649 10.6151
R2018 B.n651 B.n650 10.6151
R2019 B.n651 B.n384 10.6151
R2020 B.n657 B.n384 10.6151
R2021 B.n658 B.n657 10.6151
R2022 B.n659 B.n376 10.6151
R2023 B.n669 B.n376 10.6151
R2024 B.n670 B.n669 10.6151
R2025 B.n671 B.n670 10.6151
R2026 B.n671 B.n369 10.6151
R2027 B.n682 B.n369 10.6151
R2028 B.n683 B.n682 10.6151
R2029 B.n684 B.n683 10.6151
R2030 B.n684 B.n361 10.6151
R2031 B.n694 B.n361 10.6151
R2032 B.n695 B.n694 10.6151
R2033 B.n696 B.n695 10.6151
R2034 B.n696 B.n353 10.6151
R2035 B.n706 B.n353 10.6151
R2036 B.n707 B.n706 10.6151
R2037 B.n708 B.n707 10.6151
R2038 B.n708 B.n344 10.6151
R2039 B.n718 B.n344 10.6151
R2040 B.n719 B.n718 10.6151
R2041 B.n720 B.n719 10.6151
R2042 B.n720 B.n337 10.6151
R2043 B.n730 B.n337 10.6151
R2044 B.n731 B.n730 10.6151
R2045 B.n733 B.n731 10.6151
R2046 B.n733 B.n732 10.6151
R2047 B.n732 B.n329 10.6151
R2048 B.n744 B.n329 10.6151
R2049 B.n745 B.n744 10.6151
R2050 B.n746 B.n745 10.6151
R2051 B.n747 B.n746 10.6151
R2052 B.n748 B.n747 10.6151
R2053 B.n752 B.n748 10.6151
R2054 B.n753 B.n752 10.6151
R2055 B.n754 B.n753 10.6151
R2056 B.n755 B.n754 10.6151
R2057 B.n757 B.n755 10.6151
R2058 B.n758 B.n757 10.6151
R2059 B.n759 B.n758 10.6151
R2060 B.n760 B.n759 10.6151
R2061 B.n762 B.n760 10.6151
R2062 B.n763 B.n762 10.6151
R2063 B.n764 B.n763 10.6151
R2064 B.n765 B.n764 10.6151
R2065 B.n767 B.n765 10.6151
R2066 B.n768 B.n767 10.6151
R2067 B.n769 B.n768 10.6151
R2068 B.n770 B.n769 10.6151
R2069 B.n772 B.n770 10.6151
R2070 B.n773 B.n772 10.6151
R2071 B.n774 B.n773 10.6151
R2072 B.n775 B.n774 10.6151
R2073 B.n777 B.n775 10.6151
R2074 B.n778 B.n777 10.6151
R2075 B.n779 B.n778 10.6151
R2076 B.n780 B.n779 10.6151
R2077 B.n782 B.n780 10.6151
R2078 B.n783 B.n782 10.6151
R2079 B.n839 B.n1 10.6151
R2080 B.n839 B.n838 10.6151
R2081 B.n838 B.n837 10.6151
R2082 B.n837 B.n10 10.6151
R2083 B.n831 B.n10 10.6151
R2084 B.n831 B.n830 10.6151
R2085 B.n830 B.n829 10.6151
R2086 B.n829 B.n17 10.6151
R2087 B.n823 B.n17 10.6151
R2088 B.n823 B.n822 10.6151
R2089 B.n822 B.n821 10.6151
R2090 B.n821 B.n24 10.6151
R2091 B.n815 B.n24 10.6151
R2092 B.n815 B.n814 10.6151
R2093 B.n814 B.n813 10.6151
R2094 B.n813 B.n31 10.6151
R2095 B.n807 B.n31 10.6151
R2096 B.n807 B.n806 10.6151
R2097 B.n806 B.n805 10.6151
R2098 B.n805 B.n38 10.6151
R2099 B.n799 B.n38 10.6151
R2100 B.n799 B.n798 10.6151
R2101 B.n798 B.n797 10.6151
R2102 B.n797 B.n44 10.6151
R2103 B.n791 B.n44 10.6151
R2104 B.n791 B.n790 10.6151
R2105 B.n790 B.n789 10.6151
R2106 B.n115 B.n52 10.6151
R2107 B.n118 B.n115 10.6151
R2108 B.n119 B.n118 10.6151
R2109 B.n122 B.n119 10.6151
R2110 B.n123 B.n122 10.6151
R2111 B.n126 B.n123 10.6151
R2112 B.n127 B.n126 10.6151
R2113 B.n130 B.n127 10.6151
R2114 B.n131 B.n130 10.6151
R2115 B.n134 B.n131 10.6151
R2116 B.n135 B.n134 10.6151
R2117 B.n138 B.n135 10.6151
R2118 B.n139 B.n138 10.6151
R2119 B.n142 B.n139 10.6151
R2120 B.n143 B.n142 10.6151
R2121 B.n146 B.n143 10.6151
R2122 B.n147 B.n146 10.6151
R2123 B.n150 B.n147 10.6151
R2124 B.n151 B.n150 10.6151
R2125 B.n154 B.n151 10.6151
R2126 B.n155 B.n154 10.6151
R2127 B.n158 B.n155 10.6151
R2128 B.n159 B.n158 10.6151
R2129 B.n162 B.n159 10.6151
R2130 B.n163 B.n162 10.6151
R2131 B.n166 B.n163 10.6151
R2132 B.n167 B.n166 10.6151
R2133 B.n170 B.n167 10.6151
R2134 B.n171 B.n170 10.6151
R2135 B.n174 B.n171 10.6151
R2136 B.n175 B.n174 10.6151
R2137 B.n178 B.n175 10.6151
R2138 B.n179 B.n178 10.6151
R2139 B.n182 B.n179 10.6151
R2140 B.n183 B.n182 10.6151
R2141 B.n186 B.n183 10.6151
R2142 B.n187 B.n186 10.6151
R2143 B.n190 B.n187 10.6151
R2144 B.n191 B.n190 10.6151
R2145 B.n194 B.n191 10.6151
R2146 B.n195 B.n194 10.6151
R2147 B.n198 B.n195 10.6151
R2148 B.n199 B.n198 10.6151
R2149 B.n202 B.n199 10.6151
R2150 B.n203 B.n202 10.6151
R2151 B.n206 B.n203 10.6151
R2152 B.n207 B.n206 10.6151
R2153 B.n210 B.n207 10.6151
R2154 B.n211 B.n210 10.6151
R2155 B.n215 B.n214 10.6151
R2156 B.n218 B.n215 10.6151
R2157 B.n219 B.n218 10.6151
R2158 B.n222 B.n219 10.6151
R2159 B.n223 B.n222 10.6151
R2160 B.n226 B.n223 10.6151
R2161 B.n227 B.n226 10.6151
R2162 B.n230 B.n227 10.6151
R2163 B.n235 B.n232 10.6151
R2164 B.n236 B.n235 10.6151
R2165 B.n239 B.n236 10.6151
R2166 B.n240 B.n239 10.6151
R2167 B.n243 B.n240 10.6151
R2168 B.n244 B.n243 10.6151
R2169 B.n247 B.n244 10.6151
R2170 B.n248 B.n247 10.6151
R2171 B.n251 B.n248 10.6151
R2172 B.n252 B.n251 10.6151
R2173 B.n255 B.n252 10.6151
R2174 B.n256 B.n255 10.6151
R2175 B.n259 B.n256 10.6151
R2176 B.n260 B.n259 10.6151
R2177 B.n263 B.n260 10.6151
R2178 B.n264 B.n263 10.6151
R2179 B.n267 B.n264 10.6151
R2180 B.n268 B.n267 10.6151
R2181 B.n271 B.n268 10.6151
R2182 B.n272 B.n271 10.6151
R2183 B.n275 B.n272 10.6151
R2184 B.n276 B.n275 10.6151
R2185 B.n279 B.n276 10.6151
R2186 B.n280 B.n279 10.6151
R2187 B.n283 B.n280 10.6151
R2188 B.n284 B.n283 10.6151
R2189 B.n287 B.n284 10.6151
R2190 B.n288 B.n287 10.6151
R2191 B.n291 B.n288 10.6151
R2192 B.n292 B.n291 10.6151
R2193 B.n295 B.n292 10.6151
R2194 B.n296 B.n295 10.6151
R2195 B.n299 B.n296 10.6151
R2196 B.n300 B.n299 10.6151
R2197 B.n303 B.n300 10.6151
R2198 B.n304 B.n303 10.6151
R2199 B.n307 B.n304 10.6151
R2200 B.n308 B.n307 10.6151
R2201 B.n311 B.n308 10.6151
R2202 B.n312 B.n311 10.6151
R2203 B.n315 B.n312 10.6151
R2204 B.n316 B.n315 10.6151
R2205 B.n319 B.n316 10.6151
R2206 B.n320 B.n319 10.6151
R2207 B.n323 B.n320 10.6151
R2208 B.n324 B.n323 10.6151
R2209 B.n327 B.n324 10.6151
R2210 B.n328 B.n327 10.6151
R2211 B.n784 B.n328 10.6151
R2212 B.n680 B.t11 8.22377
R2213 B.n347 B.t5 8.22377
R2214 B.t1 B.n826 8.22377
R2215 B.n801 B.t7 8.22377
R2216 B.n847 B.n0 8.11757
R2217 B.n847 B.n1 8.11757
R2218 B.n538 B.n415 6.5566
R2219 B.n411 B.n410 6.5566
R2220 B.n214 B.n114 6.5566
R2221 B.n231 B.n230 6.5566
R2222 B.n539 B.n538 4.05904
R2223 B.n561 B.n410 4.05904
R2224 B.n211 B.n114 4.05904
R2225 B.n232 B.n231 4.05904
R2226 B.n704 B.t3 3.83803
R2227 B.t4 B.n817 3.83803
R2228 VP.n7 VP.t1 287.901
R2229 VP.n20 VP.t4 252.794
R2230 VP.n14 VP.t0 252.794
R2231 VP.n26 VP.t2 252.794
R2232 VP.n6 VP.t5 252.794
R2233 VP.n12 VP.t3 252.794
R2234 VP.n15 VP.n14 174.024
R2235 VP.n27 VP.n26 174.024
R2236 VP.n13 VP.n12 174.024
R2237 VP.n8 VP.n5 161.3
R2238 VP.n10 VP.n9 161.3
R2239 VP.n11 VP.n4 161.3
R2240 VP.n25 VP.n0 161.3
R2241 VP.n24 VP.n23 161.3
R2242 VP.n22 VP.n1 161.3
R2243 VP.n21 VP.n20 161.3
R2244 VP.n19 VP.n2 161.3
R2245 VP.n18 VP.n17 161.3
R2246 VP.n16 VP.n3 161.3
R2247 VP.n19 VP.n18 53.1199
R2248 VP.n24 VP.n1 53.1199
R2249 VP.n10 VP.n5 53.1199
R2250 VP.n15 VP.n13 46.0535
R2251 VP.n7 VP.n6 41.8164
R2252 VP.n18 VP.n3 27.8669
R2253 VP.n25 VP.n24 27.8669
R2254 VP.n11 VP.n10 27.8669
R2255 VP.n20 VP.n19 24.4675
R2256 VP.n20 VP.n1 24.4675
R2257 VP.n6 VP.n5 24.4675
R2258 VP.n8 VP.n7 17.5844
R2259 VP.n14 VP.n3 11.7447
R2260 VP.n26 VP.n25 11.7447
R2261 VP.n12 VP.n11 11.7447
R2262 VP.n9 VP.n8 0.189894
R2263 VP.n9 VP.n4 0.189894
R2264 VP.n13 VP.n4 0.189894
R2265 VP.n16 VP.n15 0.189894
R2266 VP.n17 VP.n16 0.189894
R2267 VP.n17 VP.n2 0.189894
R2268 VP.n21 VP.n2 0.189894
R2269 VP.n22 VP.n21 0.189894
R2270 VP.n23 VP.n22 0.189894
R2271 VP.n23 VP.n0 0.189894
R2272 VP.n27 VP.n0 0.189894
R2273 VP VP.n27 0.0516364
R2274 VDD1.n76 VDD1.n0 289.615
R2275 VDD1.n157 VDD1.n81 289.615
R2276 VDD1.n77 VDD1.n76 185
R2277 VDD1.n75 VDD1.n74 185
R2278 VDD1.n73 VDD1.n3 185
R2279 VDD1.n7 VDD1.n4 185
R2280 VDD1.n68 VDD1.n67 185
R2281 VDD1.n66 VDD1.n65 185
R2282 VDD1.n9 VDD1.n8 185
R2283 VDD1.n60 VDD1.n59 185
R2284 VDD1.n58 VDD1.n57 185
R2285 VDD1.n13 VDD1.n12 185
R2286 VDD1.n52 VDD1.n51 185
R2287 VDD1.n50 VDD1.n49 185
R2288 VDD1.n17 VDD1.n16 185
R2289 VDD1.n44 VDD1.n43 185
R2290 VDD1.n42 VDD1.n41 185
R2291 VDD1.n21 VDD1.n20 185
R2292 VDD1.n36 VDD1.n35 185
R2293 VDD1.n34 VDD1.n33 185
R2294 VDD1.n25 VDD1.n24 185
R2295 VDD1.n28 VDD1.n27 185
R2296 VDD1.n108 VDD1.n107 185
R2297 VDD1.n105 VDD1.n104 185
R2298 VDD1.n114 VDD1.n113 185
R2299 VDD1.n116 VDD1.n115 185
R2300 VDD1.n101 VDD1.n100 185
R2301 VDD1.n122 VDD1.n121 185
R2302 VDD1.n124 VDD1.n123 185
R2303 VDD1.n97 VDD1.n96 185
R2304 VDD1.n130 VDD1.n129 185
R2305 VDD1.n132 VDD1.n131 185
R2306 VDD1.n93 VDD1.n92 185
R2307 VDD1.n138 VDD1.n137 185
R2308 VDD1.n140 VDD1.n139 185
R2309 VDD1.n89 VDD1.n88 185
R2310 VDD1.n146 VDD1.n145 185
R2311 VDD1.n149 VDD1.n148 185
R2312 VDD1.n147 VDD1.n85 185
R2313 VDD1.n154 VDD1.n84 185
R2314 VDD1.n156 VDD1.n155 185
R2315 VDD1.n158 VDD1.n157 185
R2316 VDD1.t4 VDD1.n26 147.659
R2317 VDD1.t5 VDD1.n106 147.659
R2318 VDD1.n76 VDD1.n75 104.615
R2319 VDD1.n75 VDD1.n3 104.615
R2320 VDD1.n7 VDD1.n3 104.615
R2321 VDD1.n67 VDD1.n7 104.615
R2322 VDD1.n67 VDD1.n66 104.615
R2323 VDD1.n66 VDD1.n8 104.615
R2324 VDD1.n59 VDD1.n8 104.615
R2325 VDD1.n59 VDD1.n58 104.615
R2326 VDD1.n58 VDD1.n12 104.615
R2327 VDD1.n51 VDD1.n12 104.615
R2328 VDD1.n51 VDD1.n50 104.615
R2329 VDD1.n50 VDD1.n16 104.615
R2330 VDD1.n43 VDD1.n16 104.615
R2331 VDD1.n43 VDD1.n42 104.615
R2332 VDD1.n42 VDD1.n20 104.615
R2333 VDD1.n35 VDD1.n20 104.615
R2334 VDD1.n35 VDD1.n34 104.615
R2335 VDD1.n34 VDD1.n24 104.615
R2336 VDD1.n27 VDD1.n24 104.615
R2337 VDD1.n107 VDD1.n104 104.615
R2338 VDD1.n114 VDD1.n104 104.615
R2339 VDD1.n115 VDD1.n114 104.615
R2340 VDD1.n115 VDD1.n100 104.615
R2341 VDD1.n122 VDD1.n100 104.615
R2342 VDD1.n123 VDD1.n122 104.615
R2343 VDD1.n123 VDD1.n96 104.615
R2344 VDD1.n130 VDD1.n96 104.615
R2345 VDD1.n131 VDD1.n130 104.615
R2346 VDD1.n131 VDD1.n92 104.615
R2347 VDD1.n138 VDD1.n92 104.615
R2348 VDD1.n139 VDD1.n138 104.615
R2349 VDD1.n139 VDD1.n88 104.615
R2350 VDD1.n146 VDD1.n88 104.615
R2351 VDD1.n148 VDD1.n146 104.615
R2352 VDD1.n148 VDD1.n147 104.615
R2353 VDD1.n147 VDD1.n84 104.615
R2354 VDD1.n156 VDD1.n84 104.615
R2355 VDD1.n157 VDD1.n156 104.615
R2356 VDD1.n163 VDD1.n162 64.1497
R2357 VDD1.n165 VDD1.n164 63.83
R2358 VDD1 VDD1.n80 52.9564
R2359 VDD1.n163 VDD1.n161 52.8429
R2360 VDD1.n27 VDD1.t4 52.3082
R2361 VDD1.n107 VDD1.t5 52.3082
R2362 VDD1.n165 VDD1.n163 42.6733
R2363 VDD1.n28 VDD1.n26 15.6677
R2364 VDD1.n108 VDD1.n106 15.6677
R2365 VDD1.n74 VDD1.n73 13.1884
R2366 VDD1.n155 VDD1.n154 13.1884
R2367 VDD1.n77 VDD1.n2 12.8005
R2368 VDD1.n72 VDD1.n4 12.8005
R2369 VDD1.n29 VDD1.n25 12.8005
R2370 VDD1.n109 VDD1.n105 12.8005
R2371 VDD1.n153 VDD1.n85 12.8005
R2372 VDD1.n158 VDD1.n83 12.8005
R2373 VDD1.n78 VDD1.n0 12.0247
R2374 VDD1.n69 VDD1.n68 12.0247
R2375 VDD1.n33 VDD1.n32 12.0247
R2376 VDD1.n113 VDD1.n112 12.0247
R2377 VDD1.n150 VDD1.n149 12.0247
R2378 VDD1.n159 VDD1.n81 12.0247
R2379 VDD1.n65 VDD1.n6 11.249
R2380 VDD1.n36 VDD1.n23 11.249
R2381 VDD1.n116 VDD1.n103 11.249
R2382 VDD1.n145 VDD1.n87 11.249
R2383 VDD1.n64 VDD1.n9 10.4732
R2384 VDD1.n37 VDD1.n21 10.4732
R2385 VDD1.n117 VDD1.n101 10.4732
R2386 VDD1.n144 VDD1.n89 10.4732
R2387 VDD1.n61 VDD1.n60 9.69747
R2388 VDD1.n41 VDD1.n40 9.69747
R2389 VDD1.n121 VDD1.n120 9.69747
R2390 VDD1.n141 VDD1.n140 9.69747
R2391 VDD1.n80 VDD1.n79 9.45567
R2392 VDD1.n161 VDD1.n160 9.45567
R2393 VDD1.n54 VDD1.n53 9.3005
R2394 VDD1.n56 VDD1.n55 9.3005
R2395 VDD1.n11 VDD1.n10 9.3005
R2396 VDD1.n62 VDD1.n61 9.3005
R2397 VDD1.n64 VDD1.n63 9.3005
R2398 VDD1.n6 VDD1.n5 9.3005
R2399 VDD1.n70 VDD1.n69 9.3005
R2400 VDD1.n72 VDD1.n71 9.3005
R2401 VDD1.n79 VDD1.n78 9.3005
R2402 VDD1.n2 VDD1.n1 9.3005
R2403 VDD1.n15 VDD1.n14 9.3005
R2404 VDD1.n48 VDD1.n47 9.3005
R2405 VDD1.n46 VDD1.n45 9.3005
R2406 VDD1.n19 VDD1.n18 9.3005
R2407 VDD1.n40 VDD1.n39 9.3005
R2408 VDD1.n38 VDD1.n37 9.3005
R2409 VDD1.n23 VDD1.n22 9.3005
R2410 VDD1.n32 VDD1.n31 9.3005
R2411 VDD1.n30 VDD1.n29 9.3005
R2412 VDD1.n160 VDD1.n159 9.3005
R2413 VDD1.n83 VDD1.n82 9.3005
R2414 VDD1.n128 VDD1.n127 9.3005
R2415 VDD1.n126 VDD1.n125 9.3005
R2416 VDD1.n99 VDD1.n98 9.3005
R2417 VDD1.n120 VDD1.n119 9.3005
R2418 VDD1.n118 VDD1.n117 9.3005
R2419 VDD1.n103 VDD1.n102 9.3005
R2420 VDD1.n112 VDD1.n111 9.3005
R2421 VDD1.n110 VDD1.n109 9.3005
R2422 VDD1.n95 VDD1.n94 9.3005
R2423 VDD1.n134 VDD1.n133 9.3005
R2424 VDD1.n136 VDD1.n135 9.3005
R2425 VDD1.n91 VDD1.n90 9.3005
R2426 VDD1.n142 VDD1.n141 9.3005
R2427 VDD1.n144 VDD1.n143 9.3005
R2428 VDD1.n87 VDD1.n86 9.3005
R2429 VDD1.n151 VDD1.n150 9.3005
R2430 VDD1.n153 VDD1.n152 9.3005
R2431 VDD1.n57 VDD1.n11 8.92171
R2432 VDD1.n44 VDD1.n19 8.92171
R2433 VDD1.n124 VDD1.n99 8.92171
R2434 VDD1.n137 VDD1.n91 8.92171
R2435 VDD1.n56 VDD1.n13 8.14595
R2436 VDD1.n45 VDD1.n17 8.14595
R2437 VDD1.n125 VDD1.n97 8.14595
R2438 VDD1.n136 VDD1.n93 8.14595
R2439 VDD1.n53 VDD1.n52 7.3702
R2440 VDD1.n49 VDD1.n48 7.3702
R2441 VDD1.n129 VDD1.n128 7.3702
R2442 VDD1.n133 VDD1.n132 7.3702
R2443 VDD1.n52 VDD1.n15 6.59444
R2444 VDD1.n49 VDD1.n15 6.59444
R2445 VDD1.n129 VDD1.n95 6.59444
R2446 VDD1.n132 VDD1.n95 6.59444
R2447 VDD1.n53 VDD1.n13 5.81868
R2448 VDD1.n48 VDD1.n17 5.81868
R2449 VDD1.n128 VDD1.n97 5.81868
R2450 VDD1.n133 VDD1.n93 5.81868
R2451 VDD1.n57 VDD1.n56 5.04292
R2452 VDD1.n45 VDD1.n44 5.04292
R2453 VDD1.n125 VDD1.n124 5.04292
R2454 VDD1.n137 VDD1.n136 5.04292
R2455 VDD1.n30 VDD1.n26 4.38563
R2456 VDD1.n110 VDD1.n106 4.38563
R2457 VDD1.n60 VDD1.n11 4.26717
R2458 VDD1.n41 VDD1.n19 4.26717
R2459 VDD1.n121 VDD1.n99 4.26717
R2460 VDD1.n140 VDD1.n91 4.26717
R2461 VDD1.n61 VDD1.n9 3.49141
R2462 VDD1.n40 VDD1.n21 3.49141
R2463 VDD1.n120 VDD1.n101 3.49141
R2464 VDD1.n141 VDD1.n89 3.49141
R2465 VDD1.n65 VDD1.n64 2.71565
R2466 VDD1.n37 VDD1.n36 2.71565
R2467 VDD1.n117 VDD1.n116 2.71565
R2468 VDD1.n145 VDD1.n144 2.71565
R2469 VDD1.n80 VDD1.n0 1.93989
R2470 VDD1.n68 VDD1.n6 1.93989
R2471 VDD1.n33 VDD1.n23 1.93989
R2472 VDD1.n113 VDD1.n103 1.93989
R2473 VDD1.n149 VDD1.n87 1.93989
R2474 VDD1.n161 VDD1.n81 1.93989
R2475 VDD1.n164 VDD1.t0 1.33924
R2476 VDD1.n164 VDD1.t2 1.33924
R2477 VDD1.n162 VDD1.t1 1.33924
R2478 VDD1.n162 VDD1.t3 1.33924
R2479 VDD1.n78 VDD1.n77 1.16414
R2480 VDD1.n69 VDD1.n4 1.16414
R2481 VDD1.n32 VDD1.n25 1.16414
R2482 VDD1.n112 VDD1.n105 1.16414
R2483 VDD1.n150 VDD1.n85 1.16414
R2484 VDD1.n159 VDD1.n158 1.16414
R2485 VDD1.n74 VDD1.n2 0.388379
R2486 VDD1.n73 VDD1.n72 0.388379
R2487 VDD1.n29 VDD1.n28 0.388379
R2488 VDD1.n109 VDD1.n108 0.388379
R2489 VDD1.n154 VDD1.n153 0.388379
R2490 VDD1.n155 VDD1.n83 0.388379
R2491 VDD1 VDD1.n165 0.31731
R2492 VDD1.n79 VDD1.n1 0.155672
R2493 VDD1.n71 VDD1.n1 0.155672
R2494 VDD1.n71 VDD1.n70 0.155672
R2495 VDD1.n70 VDD1.n5 0.155672
R2496 VDD1.n63 VDD1.n5 0.155672
R2497 VDD1.n63 VDD1.n62 0.155672
R2498 VDD1.n62 VDD1.n10 0.155672
R2499 VDD1.n55 VDD1.n10 0.155672
R2500 VDD1.n55 VDD1.n54 0.155672
R2501 VDD1.n54 VDD1.n14 0.155672
R2502 VDD1.n47 VDD1.n14 0.155672
R2503 VDD1.n47 VDD1.n46 0.155672
R2504 VDD1.n46 VDD1.n18 0.155672
R2505 VDD1.n39 VDD1.n18 0.155672
R2506 VDD1.n39 VDD1.n38 0.155672
R2507 VDD1.n38 VDD1.n22 0.155672
R2508 VDD1.n31 VDD1.n22 0.155672
R2509 VDD1.n31 VDD1.n30 0.155672
R2510 VDD1.n111 VDD1.n110 0.155672
R2511 VDD1.n111 VDD1.n102 0.155672
R2512 VDD1.n118 VDD1.n102 0.155672
R2513 VDD1.n119 VDD1.n118 0.155672
R2514 VDD1.n119 VDD1.n98 0.155672
R2515 VDD1.n126 VDD1.n98 0.155672
R2516 VDD1.n127 VDD1.n126 0.155672
R2517 VDD1.n127 VDD1.n94 0.155672
R2518 VDD1.n134 VDD1.n94 0.155672
R2519 VDD1.n135 VDD1.n134 0.155672
R2520 VDD1.n135 VDD1.n90 0.155672
R2521 VDD1.n142 VDD1.n90 0.155672
R2522 VDD1.n143 VDD1.n142 0.155672
R2523 VDD1.n143 VDD1.n86 0.155672
R2524 VDD1.n151 VDD1.n86 0.155672
R2525 VDD1.n152 VDD1.n151 0.155672
R2526 VDD1.n152 VDD1.n82 0.155672
R2527 VDD1.n160 VDD1.n82 0.155672
C0 VN VTAIL 6.79474f
C1 VTAIL VDD1 9.39954f
C2 VN VDD1 0.149107f
C3 VTAIL VDD2 9.43944f
C4 VP VTAIL 6.80925f
C5 VN VDD2 7.02215f
C6 VP VN 6.28696f
C7 VDD1 VDD2 0.973764f
C8 VP VDD1 7.226439f
C9 VP VDD2 0.357894f
C10 VDD2 B 5.537411f
C11 VDD1 B 5.609575f
C12 VTAIL B 8.037611f
C13 VN B 9.81487f
C14 VP B 8.091546f
C15 VDD1.n0 B 0.029938f
C16 VDD1.n1 B 0.021823f
C17 VDD1.n2 B 0.011727f
C18 VDD1.n3 B 0.027718f
C19 VDD1.n4 B 0.012417f
C20 VDD1.n5 B 0.021823f
C21 VDD1.n6 B 0.011727f
C22 VDD1.n7 B 0.027718f
C23 VDD1.n8 B 0.027718f
C24 VDD1.n9 B 0.012417f
C25 VDD1.n10 B 0.021823f
C26 VDD1.n11 B 0.011727f
C27 VDD1.n12 B 0.027718f
C28 VDD1.n13 B 0.012417f
C29 VDD1.n14 B 0.021823f
C30 VDD1.n15 B 0.011727f
C31 VDD1.n16 B 0.027718f
C32 VDD1.n17 B 0.012417f
C33 VDD1.n18 B 0.021823f
C34 VDD1.n19 B 0.011727f
C35 VDD1.n20 B 0.027718f
C36 VDD1.n21 B 0.012417f
C37 VDD1.n22 B 0.021823f
C38 VDD1.n23 B 0.011727f
C39 VDD1.n24 B 0.027718f
C40 VDD1.n25 B 0.012417f
C41 VDD1.n26 B 0.141185f
C42 VDD1.t4 B 0.045687f
C43 VDD1.n27 B 0.020788f
C44 VDD1.n28 B 0.016374f
C45 VDD1.n29 B 0.011727f
C46 VDD1.n30 B 1.39883f
C47 VDD1.n31 B 0.021823f
C48 VDD1.n32 B 0.011727f
C49 VDD1.n33 B 0.012417f
C50 VDD1.n34 B 0.027718f
C51 VDD1.n35 B 0.027718f
C52 VDD1.n36 B 0.012417f
C53 VDD1.n37 B 0.011727f
C54 VDD1.n38 B 0.021823f
C55 VDD1.n39 B 0.021823f
C56 VDD1.n40 B 0.011727f
C57 VDD1.n41 B 0.012417f
C58 VDD1.n42 B 0.027718f
C59 VDD1.n43 B 0.027718f
C60 VDD1.n44 B 0.012417f
C61 VDD1.n45 B 0.011727f
C62 VDD1.n46 B 0.021823f
C63 VDD1.n47 B 0.021823f
C64 VDD1.n48 B 0.011727f
C65 VDD1.n49 B 0.012417f
C66 VDD1.n50 B 0.027718f
C67 VDD1.n51 B 0.027718f
C68 VDD1.n52 B 0.012417f
C69 VDD1.n53 B 0.011727f
C70 VDD1.n54 B 0.021823f
C71 VDD1.n55 B 0.021823f
C72 VDD1.n56 B 0.011727f
C73 VDD1.n57 B 0.012417f
C74 VDD1.n58 B 0.027718f
C75 VDD1.n59 B 0.027718f
C76 VDD1.n60 B 0.012417f
C77 VDD1.n61 B 0.011727f
C78 VDD1.n62 B 0.021823f
C79 VDD1.n63 B 0.021823f
C80 VDD1.n64 B 0.011727f
C81 VDD1.n65 B 0.012417f
C82 VDD1.n66 B 0.027718f
C83 VDD1.n67 B 0.027718f
C84 VDD1.n68 B 0.012417f
C85 VDD1.n69 B 0.011727f
C86 VDD1.n70 B 0.021823f
C87 VDD1.n71 B 0.021823f
C88 VDD1.n72 B 0.011727f
C89 VDD1.n73 B 0.012072f
C90 VDD1.n74 B 0.012072f
C91 VDD1.n75 B 0.027718f
C92 VDD1.n76 B 0.058702f
C93 VDD1.n77 B 0.012417f
C94 VDD1.n78 B 0.011727f
C95 VDD1.n79 B 0.054915f
C96 VDD1.n80 B 0.050736f
C97 VDD1.n81 B 0.029938f
C98 VDD1.n82 B 0.021823f
C99 VDD1.n83 B 0.011727f
C100 VDD1.n84 B 0.027718f
C101 VDD1.n85 B 0.012417f
C102 VDD1.n86 B 0.021823f
C103 VDD1.n87 B 0.011727f
C104 VDD1.n88 B 0.027718f
C105 VDD1.n89 B 0.012417f
C106 VDD1.n90 B 0.021823f
C107 VDD1.n91 B 0.011727f
C108 VDD1.n92 B 0.027718f
C109 VDD1.n93 B 0.012417f
C110 VDD1.n94 B 0.021823f
C111 VDD1.n95 B 0.011727f
C112 VDD1.n96 B 0.027718f
C113 VDD1.n97 B 0.012417f
C114 VDD1.n98 B 0.021823f
C115 VDD1.n99 B 0.011727f
C116 VDD1.n100 B 0.027718f
C117 VDD1.n101 B 0.012417f
C118 VDD1.n102 B 0.021823f
C119 VDD1.n103 B 0.011727f
C120 VDD1.n104 B 0.027718f
C121 VDD1.n105 B 0.012417f
C122 VDD1.n106 B 0.141185f
C123 VDD1.t5 B 0.045687f
C124 VDD1.n107 B 0.020788f
C125 VDD1.n108 B 0.016374f
C126 VDD1.n109 B 0.011727f
C127 VDD1.n110 B 1.39883f
C128 VDD1.n111 B 0.021823f
C129 VDD1.n112 B 0.011727f
C130 VDD1.n113 B 0.012417f
C131 VDD1.n114 B 0.027718f
C132 VDD1.n115 B 0.027718f
C133 VDD1.n116 B 0.012417f
C134 VDD1.n117 B 0.011727f
C135 VDD1.n118 B 0.021823f
C136 VDD1.n119 B 0.021823f
C137 VDD1.n120 B 0.011727f
C138 VDD1.n121 B 0.012417f
C139 VDD1.n122 B 0.027718f
C140 VDD1.n123 B 0.027718f
C141 VDD1.n124 B 0.012417f
C142 VDD1.n125 B 0.011727f
C143 VDD1.n126 B 0.021823f
C144 VDD1.n127 B 0.021823f
C145 VDD1.n128 B 0.011727f
C146 VDD1.n129 B 0.012417f
C147 VDD1.n130 B 0.027718f
C148 VDD1.n131 B 0.027718f
C149 VDD1.n132 B 0.012417f
C150 VDD1.n133 B 0.011727f
C151 VDD1.n134 B 0.021823f
C152 VDD1.n135 B 0.021823f
C153 VDD1.n136 B 0.011727f
C154 VDD1.n137 B 0.012417f
C155 VDD1.n138 B 0.027718f
C156 VDD1.n139 B 0.027718f
C157 VDD1.n140 B 0.012417f
C158 VDD1.n141 B 0.011727f
C159 VDD1.n142 B 0.021823f
C160 VDD1.n143 B 0.021823f
C161 VDD1.n144 B 0.011727f
C162 VDD1.n145 B 0.012417f
C163 VDD1.n146 B 0.027718f
C164 VDD1.n147 B 0.027718f
C165 VDD1.n148 B 0.027718f
C166 VDD1.n149 B 0.012417f
C167 VDD1.n150 B 0.011727f
C168 VDD1.n151 B 0.021823f
C169 VDD1.n152 B 0.021823f
C170 VDD1.n153 B 0.011727f
C171 VDD1.n154 B 0.012072f
C172 VDD1.n155 B 0.012072f
C173 VDD1.n156 B 0.027718f
C174 VDD1.n157 B 0.058702f
C175 VDD1.n158 B 0.012417f
C176 VDD1.n159 B 0.011727f
C177 VDD1.n160 B 0.054915f
C178 VDD1.n161 B 0.050315f
C179 VDD1.t1 B 0.255056f
C180 VDD1.t3 B 0.255056f
C181 VDD1.n162 B 2.30819f
C182 VDD1.n163 B 2.11938f
C183 VDD1.t0 B 0.255056f
C184 VDD1.t2 B 0.255056f
C185 VDD1.n164 B 2.30662f
C186 VDD1.n165 B 2.32543f
C187 VP.n0 B 0.033503f
C188 VP.t2 B 1.91389f
C189 VP.n1 B 0.059446f
C190 VP.n2 B 0.033503f
C191 VP.t4 B 1.91389f
C192 VP.n3 B 0.049644f
C193 VP.n4 B 0.033503f
C194 VP.t3 B 1.91389f
C195 VP.n5 B 0.059446f
C196 VP.t1 B 2.01242f
C197 VP.t5 B 1.91389f
C198 VP.n6 B 0.759859f
C199 VP.n7 B 0.754535f
C200 VP.n8 B 0.210688f
C201 VP.n9 B 0.033503f
C202 VP.n10 B 0.03514f
C203 VP.n11 B 0.049644f
C204 VP.n12 B 0.749949f
C205 VP.n13 B 1.61047f
C206 VP.t0 B 1.91389f
C207 VP.n14 B 0.749949f
C208 VP.n15 B 1.63662f
C209 VP.n16 B 0.033503f
C210 VP.n17 B 0.033503f
C211 VP.n18 B 0.03514f
C212 VP.n19 B 0.059446f
C213 VP.n20 B 0.715114f
C214 VP.n21 B 0.033503f
C215 VP.n22 B 0.033503f
C216 VP.n23 B 0.033503f
C217 VP.n24 B 0.03514f
C218 VP.n25 B 0.049644f
C219 VP.n26 B 0.749949f
C220 VP.n27 B 0.031205f
C221 VTAIL.t7 B 0.266259f
C222 VTAIL.t5 B 0.266259f
C223 VTAIL.n0 B 2.34456f
C224 VTAIL.n1 B 0.337283f
C225 VTAIL.n2 B 0.031253f
C226 VTAIL.n3 B 0.022782f
C227 VTAIL.n4 B 0.012242f
C228 VTAIL.n5 B 0.028935f
C229 VTAIL.n6 B 0.012962f
C230 VTAIL.n7 B 0.022782f
C231 VTAIL.n8 B 0.012242f
C232 VTAIL.n9 B 0.028935f
C233 VTAIL.n10 B 0.012962f
C234 VTAIL.n11 B 0.022782f
C235 VTAIL.n12 B 0.012242f
C236 VTAIL.n13 B 0.028935f
C237 VTAIL.n14 B 0.012962f
C238 VTAIL.n15 B 0.022782f
C239 VTAIL.n16 B 0.012242f
C240 VTAIL.n17 B 0.028935f
C241 VTAIL.n18 B 0.012962f
C242 VTAIL.n19 B 0.022782f
C243 VTAIL.n20 B 0.012242f
C244 VTAIL.n21 B 0.028935f
C245 VTAIL.n22 B 0.012962f
C246 VTAIL.n23 B 0.022782f
C247 VTAIL.n24 B 0.012242f
C248 VTAIL.n25 B 0.028935f
C249 VTAIL.n26 B 0.012962f
C250 VTAIL.n27 B 0.147386f
C251 VTAIL.t2 B 0.047694f
C252 VTAIL.n28 B 0.021701f
C253 VTAIL.n29 B 0.017093f
C254 VTAIL.n30 B 0.012242f
C255 VTAIL.n31 B 1.46027f
C256 VTAIL.n32 B 0.022782f
C257 VTAIL.n33 B 0.012242f
C258 VTAIL.n34 B 0.012962f
C259 VTAIL.n35 B 0.028935f
C260 VTAIL.n36 B 0.028935f
C261 VTAIL.n37 B 0.012962f
C262 VTAIL.n38 B 0.012242f
C263 VTAIL.n39 B 0.022782f
C264 VTAIL.n40 B 0.022782f
C265 VTAIL.n41 B 0.012242f
C266 VTAIL.n42 B 0.012962f
C267 VTAIL.n43 B 0.028935f
C268 VTAIL.n44 B 0.028935f
C269 VTAIL.n45 B 0.012962f
C270 VTAIL.n46 B 0.012242f
C271 VTAIL.n47 B 0.022782f
C272 VTAIL.n48 B 0.022782f
C273 VTAIL.n49 B 0.012242f
C274 VTAIL.n50 B 0.012962f
C275 VTAIL.n51 B 0.028935f
C276 VTAIL.n52 B 0.028935f
C277 VTAIL.n53 B 0.012962f
C278 VTAIL.n54 B 0.012242f
C279 VTAIL.n55 B 0.022782f
C280 VTAIL.n56 B 0.022782f
C281 VTAIL.n57 B 0.012242f
C282 VTAIL.n58 B 0.012962f
C283 VTAIL.n59 B 0.028935f
C284 VTAIL.n60 B 0.028935f
C285 VTAIL.n61 B 0.012962f
C286 VTAIL.n62 B 0.012242f
C287 VTAIL.n63 B 0.022782f
C288 VTAIL.n64 B 0.022782f
C289 VTAIL.n65 B 0.012242f
C290 VTAIL.n66 B 0.012962f
C291 VTAIL.n67 B 0.028935f
C292 VTAIL.n68 B 0.028935f
C293 VTAIL.n69 B 0.028935f
C294 VTAIL.n70 B 0.012962f
C295 VTAIL.n71 B 0.012242f
C296 VTAIL.n72 B 0.022782f
C297 VTAIL.n73 B 0.022782f
C298 VTAIL.n74 B 0.012242f
C299 VTAIL.n75 B 0.012602f
C300 VTAIL.n76 B 0.012602f
C301 VTAIL.n77 B 0.028935f
C302 VTAIL.n78 B 0.061281f
C303 VTAIL.n79 B 0.012962f
C304 VTAIL.n80 B 0.012242f
C305 VTAIL.n81 B 0.057327f
C306 VTAIL.n82 B 0.034287f
C307 VTAIL.n83 B 0.221752f
C308 VTAIL.t3 B 0.266259f
C309 VTAIL.t10 B 0.266259f
C310 VTAIL.n84 B 2.34456f
C311 VTAIL.n85 B 1.79167f
C312 VTAIL.t4 B 0.266259f
C313 VTAIL.t9 B 0.266259f
C314 VTAIL.n86 B 2.34457f
C315 VTAIL.n87 B 1.79166f
C316 VTAIL.n88 B 0.031253f
C317 VTAIL.n89 B 0.022782f
C318 VTAIL.n90 B 0.012242f
C319 VTAIL.n91 B 0.028935f
C320 VTAIL.n92 B 0.012962f
C321 VTAIL.n93 B 0.022782f
C322 VTAIL.n94 B 0.012242f
C323 VTAIL.n95 B 0.028935f
C324 VTAIL.n96 B 0.028935f
C325 VTAIL.n97 B 0.012962f
C326 VTAIL.n98 B 0.022782f
C327 VTAIL.n99 B 0.012242f
C328 VTAIL.n100 B 0.028935f
C329 VTAIL.n101 B 0.012962f
C330 VTAIL.n102 B 0.022782f
C331 VTAIL.n103 B 0.012242f
C332 VTAIL.n104 B 0.028935f
C333 VTAIL.n105 B 0.012962f
C334 VTAIL.n106 B 0.022782f
C335 VTAIL.n107 B 0.012242f
C336 VTAIL.n108 B 0.028935f
C337 VTAIL.n109 B 0.012962f
C338 VTAIL.n110 B 0.022782f
C339 VTAIL.n111 B 0.012242f
C340 VTAIL.n112 B 0.028935f
C341 VTAIL.n113 B 0.012962f
C342 VTAIL.n114 B 0.147386f
C343 VTAIL.t6 B 0.047694f
C344 VTAIL.n115 B 0.021701f
C345 VTAIL.n116 B 0.017093f
C346 VTAIL.n117 B 0.012242f
C347 VTAIL.n118 B 1.46027f
C348 VTAIL.n119 B 0.022782f
C349 VTAIL.n120 B 0.012242f
C350 VTAIL.n121 B 0.012962f
C351 VTAIL.n122 B 0.028935f
C352 VTAIL.n123 B 0.028935f
C353 VTAIL.n124 B 0.012962f
C354 VTAIL.n125 B 0.012242f
C355 VTAIL.n126 B 0.022782f
C356 VTAIL.n127 B 0.022782f
C357 VTAIL.n128 B 0.012242f
C358 VTAIL.n129 B 0.012962f
C359 VTAIL.n130 B 0.028935f
C360 VTAIL.n131 B 0.028935f
C361 VTAIL.n132 B 0.012962f
C362 VTAIL.n133 B 0.012242f
C363 VTAIL.n134 B 0.022782f
C364 VTAIL.n135 B 0.022782f
C365 VTAIL.n136 B 0.012242f
C366 VTAIL.n137 B 0.012962f
C367 VTAIL.n138 B 0.028935f
C368 VTAIL.n139 B 0.028935f
C369 VTAIL.n140 B 0.012962f
C370 VTAIL.n141 B 0.012242f
C371 VTAIL.n142 B 0.022782f
C372 VTAIL.n143 B 0.022782f
C373 VTAIL.n144 B 0.012242f
C374 VTAIL.n145 B 0.012962f
C375 VTAIL.n146 B 0.028935f
C376 VTAIL.n147 B 0.028935f
C377 VTAIL.n148 B 0.012962f
C378 VTAIL.n149 B 0.012242f
C379 VTAIL.n150 B 0.022782f
C380 VTAIL.n151 B 0.022782f
C381 VTAIL.n152 B 0.012242f
C382 VTAIL.n153 B 0.012962f
C383 VTAIL.n154 B 0.028935f
C384 VTAIL.n155 B 0.028935f
C385 VTAIL.n156 B 0.012962f
C386 VTAIL.n157 B 0.012242f
C387 VTAIL.n158 B 0.022782f
C388 VTAIL.n159 B 0.022782f
C389 VTAIL.n160 B 0.012242f
C390 VTAIL.n161 B 0.012602f
C391 VTAIL.n162 B 0.012602f
C392 VTAIL.n163 B 0.028935f
C393 VTAIL.n164 B 0.061281f
C394 VTAIL.n165 B 0.012962f
C395 VTAIL.n166 B 0.012242f
C396 VTAIL.n167 B 0.057327f
C397 VTAIL.n168 B 0.034287f
C398 VTAIL.n169 B 0.221752f
C399 VTAIL.t0 B 0.266259f
C400 VTAIL.t1 B 0.266259f
C401 VTAIL.n170 B 2.34457f
C402 VTAIL.n171 B 0.415584f
C403 VTAIL.n172 B 0.031253f
C404 VTAIL.n173 B 0.022782f
C405 VTAIL.n174 B 0.012242f
C406 VTAIL.n175 B 0.028935f
C407 VTAIL.n176 B 0.012962f
C408 VTAIL.n177 B 0.022782f
C409 VTAIL.n178 B 0.012242f
C410 VTAIL.n179 B 0.028935f
C411 VTAIL.n180 B 0.028935f
C412 VTAIL.n181 B 0.012962f
C413 VTAIL.n182 B 0.022782f
C414 VTAIL.n183 B 0.012242f
C415 VTAIL.n184 B 0.028935f
C416 VTAIL.n185 B 0.012962f
C417 VTAIL.n186 B 0.022782f
C418 VTAIL.n187 B 0.012242f
C419 VTAIL.n188 B 0.028935f
C420 VTAIL.n189 B 0.012962f
C421 VTAIL.n190 B 0.022782f
C422 VTAIL.n191 B 0.012242f
C423 VTAIL.n192 B 0.028935f
C424 VTAIL.n193 B 0.012962f
C425 VTAIL.n194 B 0.022782f
C426 VTAIL.n195 B 0.012242f
C427 VTAIL.n196 B 0.028935f
C428 VTAIL.n197 B 0.012962f
C429 VTAIL.n198 B 0.147386f
C430 VTAIL.t11 B 0.047694f
C431 VTAIL.n199 B 0.021701f
C432 VTAIL.n200 B 0.017093f
C433 VTAIL.n201 B 0.012242f
C434 VTAIL.n202 B 1.46027f
C435 VTAIL.n203 B 0.022782f
C436 VTAIL.n204 B 0.012242f
C437 VTAIL.n205 B 0.012962f
C438 VTAIL.n206 B 0.028935f
C439 VTAIL.n207 B 0.028935f
C440 VTAIL.n208 B 0.012962f
C441 VTAIL.n209 B 0.012242f
C442 VTAIL.n210 B 0.022782f
C443 VTAIL.n211 B 0.022782f
C444 VTAIL.n212 B 0.012242f
C445 VTAIL.n213 B 0.012962f
C446 VTAIL.n214 B 0.028935f
C447 VTAIL.n215 B 0.028935f
C448 VTAIL.n216 B 0.012962f
C449 VTAIL.n217 B 0.012242f
C450 VTAIL.n218 B 0.022782f
C451 VTAIL.n219 B 0.022782f
C452 VTAIL.n220 B 0.012242f
C453 VTAIL.n221 B 0.012962f
C454 VTAIL.n222 B 0.028935f
C455 VTAIL.n223 B 0.028935f
C456 VTAIL.n224 B 0.012962f
C457 VTAIL.n225 B 0.012242f
C458 VTAIL.n226 B 0.022782f
C459 VTAIL.n227 B 0.022782f
C460 VTAIL.n228 B 0.012242f
C461 VTAIL.n229 B 0.012962f
C462 VTAIL.n230 B 0.028935f
C463 VTAIL.n231 B 0.028935f
C464 VTAIL.n232 B 0.012962f
C465 VTAIL.n233 B 0.012242f
C466 VTAIL.n234 B 0.022782f
C467 VTAIL.n235 B 0.022782f
C468 VTAIL.n236 B 0.012242f
C469 VTAIL.n237 B 0.012962f
C470 VTAIL.n238 B 0.028935f
C471 VTAIL.n239 B 0.028935f
C472 VTAIL.n240 B 0.012962f
C473 VTAIL.n241 B 0.012242f
C474 VTAIL.n242 B 0.022782f
C475 VTAIL.n243 B 0.022782f
C476 VTAIL.n244 B 0.012242f
C477 VTAIL.n245 B 0.012602f
C478 VTAIL.n246 B 0.012602f
C479 VTAIL.n247 B 0.028935f
C480 VTAIL.n248 B 0.061281f
C481 VTAIL.n249 B 0.012962f
C482 VTAIL.n250 B 0.012242f
C483 VTAIL.n251 B 0.057327f
C484 VTAIL.n252 B 0.034287f
C485 VTAIL.n253 B 1.48772f
C486 VTAIL.n254 B 0.031253f
C487 VTAIL.n255 B 0.022782f
C488 VTAIL.n256 B 0.012242f
C489 VTAIL.n257 B 0.028935f
C490 VTAIL.n258 B 0.012962f
C491 VTAIL.n259 B 0.022782f
C492 VTAIL.n260 B 0.012242f
C493 VTAIL.n261 B 0.028935f
C494 VTAIL.n262 B 0.012962f
C495 VTAIL.n263 B 0.022782f
C496 VTAIL.n264 B 0.012242f
C497 VTAIL.n265 B 0.028935f
C498 VTAIL.n266 B 0.012962f
C499 VTAIL.n267 B 0.022782f
C500 VTAIL.n268 B 0.012242f
C501 VTAIL.n269 B 0.028935f
C502 VTAIL.n270 B 0.012962f
C503 VTAIL.n271 B 0.022782f
C504 VTAIL.n272 B 0.012242f
C505 VTAIL.n273 B 0.028935f
C506 VTAIL.n274 B 0.012962f
C507 VTAIL.n275 B 0.022782f
C508 VTAIL.n276 B 0.012242f
C509 VTAIL.n277 B 0.028935f
C510 VTAIL.n278 B 0.012962f
C511 VTAIL.n279 B 0.147386f
C512 VTAIL.t8 B 0.047694f
C513 VTAIL.n280 B 0.021701f
C514 VTAIL.n281 B 0.017093f
C515 VTAIL.n282 B 0.012242f
C516 VTAIL.n283 B 1.46027f
C517 VTAIL.n284 B 0.022782f
C518 VTAIL.n285 B 0.012242f
C519 VTAIL.n286 B 0.012962f
C520 VTAIL.n287 B 0.028935f
C521 VTAIL.n288 B 0.028935f
C522 VTAIL.n289 B 0.012962f
C523 VTAIL.n290 B 0.012242f
C524 VTAIL.n291 B 0.022782f
C525 VTAIL.n292 B 0.022782f
C526 VTAIL.n293 B 0.012242f
C527 VTAIL.n294 B 0.012962f
C528 VTAIL.n295 B 0.028935f
C529 VTAIL.n296 B 0.028935f
C530 VTAIL.n297 B 0.012962f
C531 VTAIL.n298 B 0.012242f
C532 VTAIL.n299 B 0.022782f
C533 VTAIL.n300 B 0.022782f
C534 VTAIL.n301 B 0.012242f
C535 VTAIL.n302 B 0.012962f
C536 VTAIL.n303 B 0.028935f
C537 VTAIL.n304 B 0.028935f
C538 VTAIL.n305 B 0.012962f
C539 VTAIL.n306 B 0.012242f
C540 VTAIL.n307 B 0.022782f
C541 VTAIL.n308 B 0.022782f
C542 VTAIL.n309 B 0.012242f
C543 VTAIL.n310 B 0.012962f
C544 VTAIL.n311 B 0.028935f
C545 VTAIL.n312 B 0.028935f
C546 VTAIL.n313 B 0.012962f
C547 VTAIL.n314 B 0.012242f
C548 VTAIL.n315 B 0.022782f
C549 VTAIL.n316 B 0.022782f
C550 VTAIL.n317 B 0.012242f
C551 VTAIL.n318 B 0.012962f
C552 VTAIL.n319 B 0.028935f
C553 VTAIL.n320 B 0.028935f
C554 VTAIL.n321 B 0.028935f
C555 VTAIL.n322 B 0.012962f
C556 VTAIL.n323 B 0.012242f
C557 VTAIL.n324 B 0.022782f
C558 VTAIL.n325 B 0.022782f
C559 VTAIL.n326 B 0.012242f
C560 VTAIL.n327 B 0.012602f
C561 VTAIL.n328 B 0.012602f
C562 VTAIL.n329 B 0.028935f
C563 VTAIL.n330 B 0.061281f
C564 VTAIL.n331 B 0.012962f
C565 VTAIL.n332 B 0.012242f
C566 VTAIL.n333 B 0.057327f
C567 VTAIL.n334 B 0.034287f
C568 VTAIL.n335 B 1.45592f
C569 VDD2.n0 B 0.029721f
C570 VDD2.n1 B 0.021665f
C571 VDD2.n2 B 0.011642f
C572 VDD2.n3 B 0.027517f
C573 VDD2.n4 B 0.012327f
C574 VDD2.n5 B 0.021665f
C575 VDD2.n6 B 0.011642f
C576 VDD2.n7 B 0.027517f
C577 VDD2.n8 B 0.012327f
C578 VDD2.n9 B 0.021665f
C579 VDD2.n10 B 0.011642f
C580 VDD2.n11 B 0.027517f
C581 VDD2.n12 B 0.012327f
C582 VDD2.n13 B 0.021665f
C583 VDD2.n14 B 0.011642f
C584 VDD2.n15 B 0.027517f
C585 VDD2.n16 B 0.012327f
C586 VDD2.n17 B 0.021665f
C587 VDD2.n18 B 0.011642f
C588 VDD2.n19 B 0.027517f
C589 VDD2.n20 B 0.012327f
C590 VDD2.n21 B 0.021665f
C591 VDD2.n22 B 0.011642f
C592 VDD2.n23 B 0.027517f
C593 VDD2.n24 B 0.012327f
C594 VDD2.n25 B 0.140164f
C595 VDD2.t2 B 0.045357f
C596 VDD2.n26 B 0.020638f
C597 VDD2.n27 B 0.016255f
C598 VDD2.n28 B 0.011642f
C599 VDD2.n29 B 1.38872f
C600 VDD2.n30 B 0.021665f
C601 VDD2.n31 B 0.011642f
C602 VDD2.n32 B 0.012327f
C603 VDD2.n33 B 0.027517f
C604 VDD2.n34 B 0.027517f
C605 VDD2.n35 B 0.012327f
C606 VDD2.n36 B 0.011642f
C607 VDD2.n37 B 0.021665f
C608 VDD2.n38 B 0.021665f
C609 VDD2.n39 B 0.011642f
C610 VDD2.n40 B 0.012327f
C611 VDD2.n41 B 0.027517f
C612 VDD2.n42 B 0.027517f
C613 VDD2.n43 B 0.012327f
C614 VDD2.n44 B 0.011642f
C615 VDD2.n45 B 0.021665f
C616 VDD2.n46 B 0.021665f
C617 VDD2.n47 B 0.011642f
C618 VDD2.n48 B 0.012327f
C619 VDD2.n49 B 0.027517f
C620 VDD2.n50 B 0.027517f
C621 VDD2.n51 B 0.012327f
C622 VDD2.n52 B 0.011642f
C623 VDD2.n53 B 0.021665f
C624 VDD2.n54 B 0.021665f
C625 VDD2.n55 B 0.011642f
C626 VDD2.n56 B 0.012327f
C627 VDD2.n57 B 0.027517f
C628 VDD2.n58 B 0.027517f
C629 VDD2.n59 B 0.012327f
C630 VDD2.n60 B 0.011642f
C631 VDD2.n61 B 0.021665f
C632 VDD2.n62 B 0.021665f
C633 VDD2.n63 B 0.011642f
C634 VDD2.n64 B 0.012327f
C635 VDD2.n65 B 0.027517f
C636 VDD2.n66 B 0.027517f
C637 VDD2.n67 B 0.027517f
C638 VDD2.n68 B 0.012327f
C639 VDD2.n69 B 0.011642f
C640 VDD2.n70 B 0.021665f
C641 VDD2.n71 B 0.021665f
C642 VDD2.n72 B 0.011642f
C643 VDD2.n73 B 0.011984f
C644 VDD2.n74 B 0.011984f
C645 VDD2.n75 B 0.027517f
C646 VDD2.n76 B 0.058278f
C647 VDD2.n77 B 0.012327f
C648 VDD2.n78 B 0.011642f
C649 VDD2.n79 B 0.054518f
C650 VDD2.n80 B 0.049952f
C651 VDD2.t4 B 0.253212f
C652 VDD2.t1 B 0.253212f
C653 VDD2.n81 B 2.2915f
C654 VDD2.n82 B 2.02139f
C655 VDD2.n83 B 0.029721f
C656 VDD2.n84 B 0.021665f
C657 VDD2.n85 B 0.011642f
C658 VDD2.n86 B 0.027517f
C659 VDD2.n87 B 0.012327f
C660 VDD2.n88 B 0.021665f
C661 VDD2.n89 B 0.011642f
C662 VDD2.n90 B 0.027517f
C663 VDD2.n91 B 0.027517f
C664 VDD2.n92 B 0.012327f
C665 VDD2.n93 B 0.021665f
C666 VDD2.n94 B 0.011642f
C667 VDD2.n95 B 0.027517f
C668 VDD2.n96 B 0.012327f
C669 VDD2.n97 B 0.021665f
C670 VDD2.n98 B 0.011642f
C671 VDD2.n99 B 0.027517f
C672 VDD2.n100 B 0.012327f
C673 VDD2.n101 B 0.021665f
C674 VDD2.n102 B 0.011642f
C675 VDD2.n103 B 0.027517f
C676 VDD2.n104 B 0.012327f
C677 VDD2.n105 B 0.021665f
C678 VDD2.n106 B 0.011642f
C679 VDD2.n107 B 0.027517f
C680 VDD2.n108 B 0.012327f
C681 VDD2.n109 B 0.140164f
C682 VDD2.t0 B 0.045357f
C683 VDD2.n110 B 0.020638f
C684 VDD2.n111 B 0.016255f
C685 VDD2.n112 B 0.011642f
C686 VDD2.n113 B 1.38872f
C687 VDD2.n114 B 0.021665f
C688 VDD2.n115 B 0.011642f
C689 VDD2.n116 B 0.012327f
C690 VDD2.n117 B 0.027517f
C691 VDD2.n118 B 0.027517f
C692 VDD2.n119 B 0.012327f
C693 VDD2.n120 B 0.011642f
C694 VDD2.n121 B 0.021665f
C695 VDD2.n122 B 0.021665f
C696 VDD2.n123 B 0.011642f
C697 VDD2.n124 B 0.012327f
C698 VDD2.n125 B 0.027517f
C699 VDD2.n126 B 0.027517f
C700 VDD2.n127 B 0.012327f
C701 VDD2.n128 B 0.011642f
C702 VDD2.n129 B 0.021665f
C703 VDD2.n130 B 0.021665f
C704 VDD2.n131 B 0.011642f
C705 VDD2.n132 B 0.012327f
C706 VDD2.n133 B 0.027517f
C707 VDD2.n134 B 0.027517f
C708 VDD2.n135 B 0.012327f
C709 VDD2.n136 B 0.011642f
C710 VDD2.n137 B 0.021665f
C711 VDD2.n138 B 0.021665f
C712 VDD2.n139 B 0.011642f
C713 VDD2.n140 B 0.012327f
C714 VDD2.n141 B 0.027517f
C715 VDD2.n142 B 0.027517f
C716 VDD2.n143 B 0.012327f
C717 VDD2.n144 B 0.011642f
C718 VDD2.n145 B 0.021665f
C719 VDD2.n146 B 0.021665f
C720 VDD2.n147 B 0.011642f
C721 VDD2.n148 B 0.012327f
C722 VDD2.n149 B 0.027517f
C723 VDD2.n150 B 0.027517f
C724 VDD2.n151 B 0.012327f
C725 VDD2.n152 B 0.011642f
C726 VDD2.n153 B 0.021665f
C727 VDD2.n154 B 0.021665f
C728 VDD2.n155 B 0.011642f
C729 VDD2.n156 B 0.011984f
C730 VDD2.n157 B 0.011984f
C731 VDD2.n158 B 0.027517f
C732 VDD2.n159 B 0.058278f
C733 VDD2.n160 B 0.012327f
C734 VDD2.n161 B 0.011642f
C735 VDD2.n162 B 0.054518f
C736 VDD2.n163 B 0.047535f
C737 VDD2.n164 B 2.12804f
C738 VDD2.t3 B 0.253212f
C739 VDD2.t5 B 0.253212f
C740 VDD2.n165 B 2.29148f
C741 VN.n0 B 0.033096f
C742 VN.t1 B 1.89065f
C743 VN.n1 B 0.058724f
C744 VN.t2 B 1.98798f
C745 VN.t4 B 1.89065f
C746 VN.n2 B 0.750631f
C747 VN.n3 B 0.745372f
C748 VN.n4 B 0.208129f
C749 VN.n5 B 0.033096f
C750 VN.n6 B 0.034713f
C751 VN.n7 B 0.049041f
C752 VN.n8 B 0.740842f
C753 VN.n9 B 0.030826f
C754 VN.n10 B 0.033096f
C755 VN.t5 B 1.89065f
C756 VN.n11 B 0.058724f
C757 VN.t3 B 1.98798f
C758 VN.t0 B 1.89065f
C759 VN.n12 B 0.750631f
C760 VN.n13 B 0.745372f
C761 VN.n14 B 0.208129f
C762 VN.n15 B 0.033096f
C763 VN.n16 B 0.034713f
C764 VN.n17 B 0.049041f
C765 VN.n18 B 0.740842f
C766 VN.n19 B 1.61252f
.ends

