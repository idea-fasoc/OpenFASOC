* NGSPICE file created from diff_pair_sample_1695.ext - technology: sky130A

.subckt diff_pair_sample_1695 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VN.t0 VDD2.t3 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=1.56255 ps=9.8 w=9.47 l=1.41
X1 VDD1.t7 VP.t0 VTAIL.t2 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=3.6933 ps=19.72 w=9.47 l=1.41
X2 VDD2.t2 VN.t1 VTAIL.t14 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
X3 VTAIL.t13 VN.t2 VDD2.t7 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=1.56255 ps=9.8 w=9.47 l=1.41
X4 B.t11 B.t9 B.t10 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=0 ps=0 w=9.47 l=1.41
X5 VTAIL.t1 VP.t1 VDD1.t6 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=1.56255 ps=9.8 w=9.47 l=1.41
X6 VTAIL.t4 VP.t2 VDD1.t5 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
X7 B.t8 B.t6 B.t7 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=0 ps=0 w=9.47 l=1.41
X8 VDD2.t5 VN.t3 VTAIL.t12 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=3.6933 ps=19.72 w=9.47 l=1.41
X9 VTAIL.t6 VP.t3 VDD1.t4 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
X10 B.t5 B.t3 B.t4 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=0 ps=0 w=9.47 l=1.41
X11 VDD2.t1 VN.t4 VTAIL.t11 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
X12 VDD1.t3 VP.t4 VTAIL.t3 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
X13 VTAIL.t10 VN.t5 VDD2.t6 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
X14 VTAIL.t9 VN.t6 VDD2.t0 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
X15 B.t2 B.t0 B.t1 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=0 ps=0 w=9.47 l=1.41
X16 VDD1.t2 VP.t5 VTAIL.t5 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=3.6933 ps=19.72 w=9.47 l=1.41
X17 VTAIL.t7 VP.t6 VDD1.t1 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=3.6933 pd=19.72 as=1.56255 ps=9.8 w=9.47 l=1.41
X18 VDD2.t4 VN.t7 VTAIL.t8 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=3.6933 ps=19.72 w=9.47 l=1.41
X19 VDD1.t0 VP.t7 VTAIL.t0 w_n2710_n2862# sky130_fd_pr__pfet_01v8 ad=1.56255 pd=9.8 as=1.56255 ps=9.8 w=9.47 l=1.41
R0 VN.n5 VN.t0 193.107
R1 VN.n24 VN.t3 193.107
R2 VN.n18 VN.n17 180.385
R3 VN.n37 VN.n36 180.385
R4 VN.n4 VN.t1 161.863
R5 VN.n10 VN.t5 161.863
R6 VN.n17 VN.t7 161.863
R7 VN.n23 VN.t6 161.863
R8 VN.n29 VN.t4 161.863
R9 VN.n36 VN.t2 161.863
R10 VN.n35 VN.n19 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n32 VN.n20 161.3
R13 VN.n31 VN.n30 161.3
R14 VN.n28 VN.n21 161.3
R15 VN.n27 VN.n26 161.3
R16 VN.n25 VN.n22 161.3
R17 VN.n16 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n15 VN.n1 56.5193
R25 VN.n34 VN.n20 56.5193
R26 VN.n5 VN.n4 47.8106
R27 VN.n24 VN.n23 47.8106
R28 VN VN.n37 43.6236
R29 VN.n8 VN.n3 40.4934
R30 VN.n9 VN.n8 40.4934
R31 VN.n27 VN.n22 40.4934
R32 VN.n28 VN.n27 40.4934
R33 VN.n11 VN.n1 24.4675
R34 VN.n16 VN.n15 24.4675
R35 VN.n30 VN.n20 24.4675
R36 VN.n35 VN.n34 24.4675
R37 VN.n25 VN.n24 18.2406
R38 VN.n6 VN.n5 18.2406
R39 VN.n4 VN.n3 18.1061
R40 VN.n10 VN.n9 18.1061
R41 VN.n23 VN.n22 18.1061
R42 VN.n29 VN.n28 18.1061
R43 VN.n11 VN.n10 6.36192
R44 VN.n30 VN.n29 6.36192
R45 VN.n17 VN.n16 5.38324
R46 VN.n36 VN.n35 5.38324
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n26 VN.n21 0.189894
R53 VN.n26 VN.n25 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VDD2.n2 VDD2.n1 83.736
R63 VDD2.n2 VDD2.n0 83.736
R64 VDD2 VDD2.n5 83.7331
R65 VDD2.n4 VDD2.n3 83.0415
R66 VDD2.n4 VDD2.n2 38.6291
R67 VDD2.n5 VDD2.t0 3.43292
R68 VDD2.n5 VDD2.t5 3.43292
R69 VDD2.n3 VDD2.t7 3.43292
R70 VDD2.n3 VDD2.t1 3.43292
R71 VDD2.n1 VDD2.t6 3.43292
R72 VDD2.n1 VDD2.t4 3.43292
R73 VDD2.n0 VDD2.t3 3.43292
R74 VDD2.n0 VDD2.t2 3.43292
R75 VDD2 VDD2.n4 0.80869
R76 VTAIL.n402 VTAIL.n358 756.745
R77 VTAIL.n46 VTAIL.n2 756.745
R78 VTAIL.n96 VTAIL.n52 756.745
R79 VTAIL.n148 VTAIL.n104 756.745
R80 VTAIL.n352 VTAIL.n308 756.745
R81 VTAIL.n300 VTAIL.n256 756.745
R82 VTAIL.n250 VTAIL.n206 756.745
R83 VTAIL.n198 VTAIL.n154 756.745
R84 VTAIL.n375 VTAIL.n374 585
R85 VTAIL.n377 VTAIL.n376 585
R86 VTAIL.n370 VTAIL.n369 585
R87 VTAIL.n383 VTAIL.n382 585
R88 VTAIL.n385 VTAIL.n384 585
R89 VTAIL.n366 VTAIL.n365 585
R90 VTAIL.n392 VTAIL.n391 585
R91 VTAIL.n393 VTAIL.n364 585
R92 VTAIL.n395 VTAIL.n394 585
R93 VTAIL.n362 VTAIL.n361 585
R94 VTAIL.n401 VTAIL.n400 585
R95 VTAIL.n403 VTAIL.n402 585
R96 VTAIL.n19 VTAIL.n18 585
R97 VTAIL.n21 VTAIL.n20 585
R98 VTAIL.n14 VTAIL.n13 585
R99 VTAIL.n27 VTAIL.n26 585
R100 VTAIL.n29 VTAIL.n28 585
R101 VTAIL.n10 VTAIL.n9 585
R102 VTAIL.n36 VTAIL.n35 585
R103 VTAIL.n37 VTAIL.n8 585
R104 VTAIL.n39 VTAIL.n38 585
R105 VTAIL.n6 VTAIL.n5 585
R106 VTAIL.n45 VTAIL.n44 585
R107 VTAIL.n47 VTAIL.n46 585
R108 VTAIL.n69 VTAIL.n68 585
R109 VTAIL.n71 VTAIL.n70 585
R110 VTAIL.n64 VTAIL.n63 585
R111 VTAIL.n77 VTAIL.n76 585
R112 VTAIL.n79 VTAIL.n78 585
R113 VTAIL.n60 VTAIL.n59 585
R114 VTAIL.n86 VTAIL.n85 585
R115 VTAIL.n87 VTAIL.n58 585
R116 VTAIL.n89 VTAIL.n88 585
R117 VTAIL.n56 VTAIL.n55 585
R118 VTAIL.n95 VTAIL.n94 585
R119 VTAIL.n97 VTAIL.n96 585
R120 VTAIL.n121 VTAIL.n120 585
R121 VTAIL.n123 VTAIL.n122 585
R122 VTAIL.n116 VTAIL.n115 585
R123 VTAIL.n129 VTAIL.n128 585
R124 VTAIL.n131 VTAIL.n130 585
R125 VTAIL.n112 VTAIL.n111 585
R126 VTAIL.n138 VTAIL.n137 585
R127 VTAIL.n139 VTAIL.n110 585
R128 VTAIL.n141 VTAIL.n140 585
R129 VTAIL.n108 VTAIL.n107 585
R130 VTAIL.n147 VTAIL.n146 585
R131 VTAIL.n149 VTAIL.n148 585
R132 VTAIL.n353 VTAIL.n352 585
R133 VTAIL.n351 VTAIL.n350 585
R134 VTAIL.n312 VTAIL.n311 585
R135 VTAIL.n316 VTAIL.n314 585
R136 VTAIL.n345 VTAIL.n344 585
R137 VTAIL.n343 VTAIL.n342 585
R138 VTAIL.n318 VTAIL.n317 585
R139 VTAIL.n337 VTAIL.n336 585
R140 VTAIL.n335 VTAIL.n334 585
R141 VTAIL.n322 VTAIL.n321 585
R142 VTAIL.n329 VTAIL.n328 585
R143 VTAIL.n327 VTAIL.n326 585
R144 VTAIL.n301 VTAIL.n300 585
R145 VTAIL.n299 VTAIL.n298 585
R146 VTAIL.n260 VTAIL.n259 585
R147 VTAIL.n264 VTAIL.n262 585
R148 VTAIL.n293 VTAIL.n292 585
R149 VTAIL.n291 VTAIL.n290 585
R150 VTAIL.n266 VTAIL.n265 585
R151 VTAIL.n285 VTAIL.n284 585
R152 VTAIL.n283 VTAIL.n282 585
R153 VTAIL.n270 VTAIL.n269 585
R154 VTAIL.n277 VTAIL.n276 585
R155 VTAIL.n275 VTAIL.n274 585
R156 VTAIL.n251 VTAIL.n250 585
R157 VTAIL.n249 VTAIL.n248 585
R158 VTAIL.n210 VTAIL.n209 585
R159 VTAIL.n214 VTAIL.n212 585
R160 VTAIL.n243 VTAIL.n242 585
R161 VTAIL.n241 VTAIL.n240 585
R162 VTAIL.n216 VTAIL.n215 585
R163 VTAIL.n235 VTAIL.n234 585
R164 VTAIL.n233 VTAIL.n232 585
R165 VTAIL.n220 VTAIL.n219 585
R166 VTAIL.n227 VTAIL.n226 585
R167 VTAIL.n225 VTAIL.n224 585
R168 VTAIL.n199 VTAIL.n198 585
R169 VTAIL.n197 VTAIL.n196 585
R170 VTAIL.n158 VTAIL.n157 585
R171 VTAIL.n162 VTAIL.n160 585
R172 VTAIL.n191 VTAIL.n190 585
R173 VTAIL.n189 VTAIL.n188 585
R174 VTAIL.n164 VTAIL.n163 585
R175 VTAIL.n183 VTAIL.n182 585
R176 VTAIL.n181 VTAIL.n180 585
R177 VTAIL.n168 VTAIL.n167 585
R178 VTAIL.n175 VTAIL.n174 585
R179 VTAIL.n173 VTAIL.n172 585
R180 VTAIL.n373 VTAIL.t8 329.038
R181 VTAIL.n17 VTAIL.t15 329.038
R182 VTAIL.n67 VTAIL.t2 329.038
R183 VTAIL.n119 VTAIL.t7 329.038
R184 VTAIL.n325 VTAIL.t5 329.038
R185 VTAIL.n273 VTAIL.t1 329.038
R186 VTAIL.n223 VTAIL.t12 329.038
R187 VTAIL.n171 VTAIL.t13 329.038
R188 VTAIL.n376 VTAIL.n375 171.744
R189 VTAIL.n376 VTAIL.n369 171.744
R190 VTAIL.n383 VTAIL.n369 171.744
R191 VTAIL.n384 VTAIL.n383 171.744
R192 VTAIL.n384 VTAIL.n365 171.744
R193 VTAIL.n392 VTAIL.n365 171.744
R194 VTAIL.n393 VTAIL.n392 171.744
R195 VTAIL.n394 VTAIL.n393 171.744
R196 VTAIL.n394 VTAIL.n361 171.744
R197 VTAIL.n401 VTAIL.n361 171.744
R198 VTAIL.n402 VTAIL.n401 171.744
R199 VTAIL.n20 VTAIL.n19 171.744
R200 VTAIL.n20 VTAIL.n13 171.744
R201 VTAIL.n27 VTAIL.n13 171.744
R202 VTAIL.n28 VTAIL.n27 171.744
R203 VTAIL.n28 VTAIL.n9 171.744
R204 VTAIL.n36 VTAIL.n9 171.744
R205 VTAIL.n37 VTAIL.n36 171.744
R206 VTAIL.n38 VTAIL.n37 171.744
R207 VTAIL.n38 VTAIL.n5 171.744
R208 VTAIL.n45 VTAIL.n5 171.744
R209 VTAIL.n46 VTAIL.n45 171.744
R210 VTAIL.n70 VTAIL.n69 171.744
R211 VTAIL.n70 VTAIL.n63 171.744
R212 VTAIL.n77 VTAIL.n63 171.744
R213 VTAIL.n78 VTAIL.n77 171.744
R214 VTAIL.n78 VTAIL.n59 171.744
R215 VTAIL.n86 VTAIL.n59 171.744
R216 VTAIL.n87 VTAIL.n86 171.744
R217 VTAIL.n88 VTAIL.n87 171.744
R218 VTAIL.n88 VTAIL.n55 171.744
R219 VTAIL.n95 VTAIL.n55 171.744
R220 VTAIL.n96 VTAIL.n95 171.744
R221 VTAIL.n122 VTAIL.n121 171.744
R222 VTAIL.n122 VTAIL.n115 171.744
R223 VTAIL.n129 VTAIL.n115 171.744
R224 VTAIL.n130 VTAIL.n129 171.744
R225 VTAIL.n130 VTAIL.n111 171.744
R226 VTAIL.n138 VTAIL.n111 171.744
R227 VTAIL.n139 VTAIL.n138 171.744
R228 VTAIL.n140 VTAIL.n139 171.744
R229 VTAIL.n140 VTAIL.n107 171.744
R230 VTAIL.n147 VTAIL.n107 171.744
R231 VTAIL.n148 VTAIL.n147 171.744
R232 VTAIL.n352 VTAIL.n351 171.744
R233 VTAIL.n351 VTAIL.n311 171.744
R234 VTAIL.n316 VTAIL.n311 171.744
R235 VTAIL.n344 VTAIL.n316 171.744
R236 VTAIL.n344 VTAIL.n343 171.744
R237 VTAIL.n343 VTAIL.n317 171.744
R238 VTAIL.n336 VTAIL.n317 171.744
R239 VTAIL.n336 VTAIL.n335 171.744
R240 VTAIL.n335 VTAIL.n321 171.744
R241 VTAIL.n328 VTAIL.n321 171.744
R242 VTAIL.n328 VTAIL.n327 171.744
R243 VTAIL.n300 VTAIL.n299 171.744
R244 VTAIL.n299 VTAIL.n259 171.744
R245 VTAIL.n264 VTAIL.n259 171.744
R246 VTAIL.n292 VTAIL.n264 171.744
R247 VTAIL.n292 VTAIL.n291 171.744
R248 VTAIL.n291 VTAIL.n265 171.744
R249 VTAIL.n284 VTAIL.n265 171.744
R250 VTAIL.n284 VTAIL.n283 171.744
R251 VTAIL.n283 VTAIL.n269 171.744
R252 VTAIL.n276 VTAIL.n269 171.744
R253 VTAIL.n276 VTAIL.n275 171.744
R254 VTAIL.n250 VTAIL.n249 171.744
R255 VTAIL.n249 VTAIL.n209 171.744
R256 VTAIL.n214 VTAIL.n209 171.744
R257 VTAIL.n242 VTAIL.n214 171.744
R258 VTAIL.n242 VTAIL.n241 171.744
R259 VTAIL.n241 VTAIL.n215 171.744
R260 VTAIL.n234 VTAIL.n215 171.744
R261 VTAIL.n234 VTAIL.n233 171.744
R262 VTAIL.n233 VTAIL.n219 171.744
R263 VTAIL.n226 VTAIL.n219 171.744
R264 VTAIL.n226 VTAIL.n225 171.744
R265 VTAIL.n198 VTAIL.n197 171.744
R266 VTAIL.n197 VTAIL.n157 171.744
R267 VTAIL.n162 VTAIL.n157 171.744
R268 VTAIL.n190 VTAIL.n162 171.744
R269 VTAIL.n190 VTAIL.n189 171.744
R270 VTAIL.n189 VTAIL.n163 171.744
R271 VTAIL.n182 VTAIL.n163 171.744
R272 VTAIL.n182 VTAIL.n181 171.744
R273 VTAIL.n181 VTAIL.n167 171.744
R274 VTAIL.n174 VTAIL.n167 171.744
R275 VTAIL.n174 VTAIL.n173 171.744
R276 VTAIL.n375 VTAIL.t8 85.8723
R277 VTAIL.n19 VTAIL.t15 85.8723
R278 VTAIL.n69 VTAIL.t2 85.8723
R279 VTAIL.n121 VTAIL.t7 85.8723
R280 VTAIL.n327 VTAIL.t5 85.8723
R281 VTAIL.n275 VTAIL.t1 85.8723
R282 VTAIL.n225 VTAIL.t12 85.8723
R283 VTAIL.n173 VTAIL.t13 85.8723
R284 VTAIL.n307 VTAIL.n306 66.3627
R285 VTAIL.n205 VTAIL.n204 66.3627
R286 VTAIL.n1 VTAIL.n0 66.3625
R287 VTAIL.n103 VTAIL.n102 66.3625
R288 VTAIL.n407 VTAIL.n406 36.646
R289 VTAIL.n51 VTAIL.n50 36.646
R290 VTAIL.n101 VTAIL.n100 36.646
R291 VTAIL.n153 VTAIL.n152 36.646
R292 VTAIL.n357 VTAIL.n356 36.646
R293 VTAIL.n305 VTAIL.n304 36.646
R294 VTAIL.n255 VTAIL.n254 36.646
R295 VTAIL.n203 VTAIL.n202 36.646
R296 VTAIL.n407 VTAIL.n357 22.0307
R297 VTAIL.n203 VTAIL.n153 22.0307
R298 VTAIL.n395 VTAIL.n362 13.1884
R299 VTAIL.n39 VTAIL.n6 13.1884
R300 VTAIL.n89 VTAIL.n56 13.1884
R301 VTAIL.n141 VTAIL.n108 13.1884
R302 VTAIL.n314 VTAIL.n312 13.1884
R303 VTAIL.n262 VTAIL.n260 13.1884
R304 VTAIL.n212 VTAIL.n210 13.1884
R305 VTAIL.n160 VTAIL.n158 13.1884
R306 VTAIL.n396 VTAIL.n364 12.8005
R307 VTAIL.n400 VTAIL.n399 12.8005
R308 VTAIL.n40 VTAIL.n8 12.8005
R309 VTAIL.n44 VTAIL.n43 12.8005
R310 VTAIL.n90 VTAIL.n58 12.8005
R311 VTAIL.n94 VTAIL.n93 12.8005
R312 VTAIL.n142 VTAIL.n110 12.8005
R313 VTAIL.n146 VTAIL.n145 12.8005
R314 VTAIL.n350 VTAIL.n349 12.8005
R315 VTAIL.n346 VTAIL.n345 12.8005
R316 VTAIL.n298 VTAIL.n297 12.8005
R317 VTAIL.n294 VTAIL.n293 12.8005
R318 VTAIL.n248 VTAIL.n247 12.8005
R319 VTAIL.n244 VTAIL.n243 12.8005
R320 VTAIL.n196 VTAIL.n195 12.8005
R321 VTAIL.n192 VTAIL.n191 12.8005
R322 VTAIL.n391 VTAIL.n390 12.0247
R323 VTAIL.n403 VTAIL.n360 12.0247
R324 VTAIL.n35 VTAIL.n34 12.0247
R325 VTAIL.n47 VTAIL.n4 12.0247
R326 VTAIL.n85 VTAIL.n84 12.0247
R327 VTAIL.n97 VTAIL.n54 12.0247
R328 VTAIL.n137 VTAIL.n136 12.0247
R329 VTAIL.n149 VTAIL.n106 12.0247
R330 VTAIL.n353 VTAIL.n310 12.0247
R331 VTAIL.n342 VTAIL.n315 12.0247
R332 VTAIL.n301 VTAIL.n258 12.0247
R333 VTAIL.n290 VTAIL.n263 12.0247
R334 VTAIL.n251 VTAIL.n208 12.0247
R335 VTAIL.n240 VTAIL.n213 12.0247
R336 VTAIL.n199 VTAIL.n156 12.0247
R337 VTAIL.n188 VTAIL.n161 12.0247
R338 VTAIL.n389 VTAIL.n366 11.249
R339 VTAIL.n404 VTAIL.n358 11.249
R340 VTAIL.n33 VTAIL.n10 11.249
R341 VTAIL.n48 VTAIL.n2 11.249
R342 VTAIL.n83 VTAIL.n60 11.249
R343 VTAIL.n98 VTAIL.n52 11.249
R344 VTAIL.n135 VTAIL.n112 11.249
R345 VTAIL.n150 VTAIL.n104 11.249
R346 VTAIL.n354 VTAIL.n308 11.249
R347 VTAIL.n341 VTAIL.n318 11.249
R348 VTAIL.n302 VTAIL.n256 11.249
R349 VTAIL.n289 VTAIL.n266 11.249
R350 VTAIL.n252 VTAIL.n206 11.249
R351 VTAIL.n239 VTAIL.n216 11.249
R352 VTAIL.n200 VTAIL.n154 11.249
R353 VTAIL.n187 VTAIL.n164 11.249
R354 VTAIL.n374 VTAIL.n373 10.7239
R355 VTAIL.n18 VTAIL.n17 10.7239
R356 VTAIL.n68 VTAIL.n67 10.7239
R357 VTAIL.n120 VTAIL.n119 10.7239
R358 VTAIL.n326 VTAIL.n325 10.7239
R359 VTAIL.n274 VTAIL.n273 10.7239
R360 VTAIL.n224 VTAIL.n223 10.7239
R361 VTAIL.n172 VTAIL.n171 10.7239
R362 VTAIL.n386 VTAIL.n385 10.4732
R363 VTAIL.n30 VTAIL.n29 10.4732
R364 VTAIL.n80 VTAIL.n79 10.4732
R365 VTAIL.n132 VTAIL.n131 10.4732
R366 VTAIL.n338 VTAIL.n337 10.4732
R367 VTAIL.n286 VTAIL.n285 10.4732
R368 VTAIL.n236 VTAIL.n235 10.4732
R369 VTAIL.n184 VTAIL.n183 10.4732
R370 VTAIL.n382 VTAIL.n368 9.69747
R371 VTAIL.n26 VTAIL.n12 9.69747
R372 VTAIL.n76 VTAIL.n62 9.69747
R373 VTAIL.n128 VTAIL.n114 9.69747
R374 VTAIL.n334 VTAIL.n320 9.69747
R375 VTAIL.n282 VTAIL.n268 9.69747
R376 VTAIL.n232 VTAIL.n218 9.69747
R377 VTAIL.n180 VTAIL.n166 9.69747
R378 VTAIL.n406 VTAIL.n405 9.45567
R379 VTAIL.n50 VTAIL.n49 9.45567
R380 VTAIL.n100 VTAIL.n99 9.45567
R381 VTAIL.n152 VTAIL.n151 9.45567
R382 VTAIL.n356 VTAIL.n355 9.45567
R383 VTAIL.n304 VTAIL.n303 9.45567
R384 VTAIL.n254 VTAIL.n253 9.45567
R385 VTAIL.n202 VTAIL.n201 9.45567
R386 VTAIL.n405 VTAIL.n404 9.3005
R387 VTAIL.n360 VTAIL.n359 9.3005
R388 VTAIL.n399 VTAIL.n398 9.3005
R389 VTAIL.n372 VTAIL.n371 9.3005
R390 VTAIL.n379 VTAIL.n378 9.3005
R391 VTAIL.n381 VTAIL.n380 9.3005
R392 VTAIL.n368 VTAIL.n367 9.3005
R393 VTAIL.n387 VTAIL.n386 9.3005
R394 VTAIL.n389 VTAIL.n388 9.3005
R395 VTAIL.n390 VTAIL.n363 9.3005
R396 VTAIL.n397 VTAIL.n396 9.3005
R397 VTAIL.n49 VTAIL.n48 9.3005
R398 VTAIL.n4 VTAIL.n3 9.3005
R399 VTAIL.n43 VTAIL.n42 9.3005
R400 VTAIL.n16 VTAIL.n15 9.3005
R401 VTAIL.n23 VTAIL.n22 9.3005
R402 VTAIL.n25 VTAIL.n24 9.3005
R403 VTAIL.n12 VTAIL.n11 9.3005
R404 VTAIL.n31 VTAIL.n30 9.3005
R405 VTAIL.n33 VTAIL.n32 9.3005
R406 VTAIL.n34 VTAIL.n7 9.3005
R407 VTAIL.n41 VTAIL.n40 9.3005
R408 VTAIL.n99 VTAIL.n98 9.3005
R409 VTAIL.n54 VTAIL.n53 9.3005
R410 VTAIL.n93 VTAIL.n92 9.3005
R411 VTAIL.n66 VTAIL.n65 9.3005
R412 VTAIL.n73 VTAIL.n72 9.3005
R413 VTAIL.n75 VTAIL.n74 9.3005
R414 VTAIL.n62 VTAIL.n61 9.3005
R415 VTAIL.n81 VTAIL.n80 9.3005
R416 VTAIL.n83 VTAIL.n82 9.3005
R417 VTAIL.n84 VTAIL.n57 9.3005
R418 VTAIL.n91 VTAIL.n90 9.3005
R419 VTAIL.n151 VTAIL.n150 9.3005
R420 VTAIL.n106 VTAIL.n105 9.3005
R421 VTAIL.n145 VTAIL.n144 9.3005
R422 VTAIL.n118 VTAIL.n117 9.3005
R423 VTAIL.n125 VTAIL.n124 9.3005
R424 VTAIL.n127 VTAIL.n126 9.3005
R425 VTAIL.n114 VTAIL.n113 9.3005
R426 VTAIL.n133 VTAIL.n132 9.3005
R427 VTAIL.n135 VTAIL.n134 9.3005
R428 VTAIL.n136 VTAIL.n109 9.3005
R429 VTAIL.n143 VTAIL.n142 9.3005
R430 VTAIL.n324 VTAIL.n323 9.3005
R431 VTAIL.n331 VTAIL.n330 9.3005
R432 VTAIL.n333 VTAIL.n332 9.3005
R433 VTAIL.n320 VTAIL.n319 9.3005
R434 VTAIL.n339 VTAIL.n338 9.3005
R435 VTAIL.n341 VTAIL.n340 9.3005
R436 VTAIL.n315 VTAIL.n313 9.3005
R437 VTAIL.n347 VTAIL.n346 9.3005
R438 VTAIL.n355 VTAIL.n354 9.3005
R439 VTAIL.n310 VTAIL.n309 9.3005
R440 VTAIL.n349 VTAIL.n348 9.3005
R441 VTAIL.n272 VTAIL.n271 9.3005
R442 VTAIL.n279 VTAIL.n278 9.3005
R443 VTAIL.n281 VTAIL.n280 9.3005
R444 VTAIL.n268 VTAIL.n267 9.3005
R445 VTAIL.n287 VTAIL.n286 9.3005
R446 VTAIL.n289 VTAIL.n288 9.3005
R447 VTAIL.n263 VTAIL.n261 9.3005
R448 VTAIL.n295 VTAIL.n294 9.3005
R449 VTAIL.n303 VTAIL.n302 9.3005
R450 VTAIL.n258 VTAIL.n257 9.3005
R451 VTAIL.n297 VTAIL.n296 9.3005
R452 VTAIL.n222 VTAIL.n221 9.3005
R453 VTAIL.n229 VTAIL.n228 9.3005
R454 VTAIL.n231 VTAIL.n230 9.3005
R455 VTAIL.n218 VTAIL.n217 9.3005
R456 VTAIL.n237 VTAIL.n236 9.3005
R457 VTAIL.n239 VTAIL.n238 9.3005
R458 VTAIL.n213 VTAIL.n211 9.3005
R459 VTAIL.n245 VTAIL.n244 9.3005
R460 VTAIL.n253 VTAIL.n252 9.3005
R461 VTAIL.n208 VTAIL.n207 9.3005
R462 VTAIL.n247 VTAIL.n246 9.3005
R463 VTAIL.n170 VTAIL.n169 9.3005
R464 VTAIL.n177 VTAIL.n176 9.3005
R465 VTAIL.n179 VTAIL.n178 9.3005
R466 VTAIL.n166 VTAIL.n165 9.3005
R467 VTAIL.n185 VTAIL.n184 9.3005
R468 VTAIL.n187 VTAIL.n186 9.3005
R469 VTAIL.n161 VTAIL.n159 9.3005
R470 VTAIL.n193 VTAIL.n192 9.3005
R471 VTAIL.n201 VTAIL.n200 9.3005
R472 VTAIL.n156 VTAIL.n155 9.3005
R473 VTAIL.n195 VTAIL.n194 9.3005
R474 VTAIL.n381 VTAIL.n370 8.92171
R475 VTAIL.n25 VTAIL.n14 8.92171
R476 VTAIL.n75 VTAIL.n64 8.92171
R477 VTAIL.n127 VTAIL.n116 8.92171
R478 VTAIL.n333 VTAIL.n322 8.92171
R479 VTAIL.n281 VTAIL.n270 8.92171
R480 VTAIL.n231 VTAIL.n220 8.92171
R481 VTAIL.n179 VTAIL.n168 8.92171
R482 VTAIL.n378 VTAIL.n377 8.14595
R483 VTAIL.n22 VTAIL.n21 8.14595
R484 VTAIL.n72 VTAIL.n71 8.14595
R485 VTAIL.n124 VTAIL.n123 8.14595
R486 VTAIL.n330 VTAIL.n329 8.14595
R487 VTAIL.n278 VTAIL.n277 8.14595
R488 VTAIL.n228 VTAIL.n227 8.14595
R489 VTAIL.n176 VTAIL.n175 8.14595
R490 VTAIL.n374 VTAIL.n372 7.3702
R491 VTAIL.n18 VTAIL.n16 7.3702
R492 VTAIL.n68 VTAIL.n66 7.3702
R493 VTAIL.n120 VTAIL.n118 7.3702
R494 VTAIL.n326 VTAIL.n324 7.3702
R495 VTAIL.n274 VTAIL.n272 7.3702
R496 VTAIL.n224 VTAIL.n222 7.3702
R497 VTAIL.n172 VTAIL.n170 7.3702
R498 VTAIL.n377 VTAIL.n372 5.81868
R499 VTAIL.n21 VTAIL.n16 5.81868
R500 VTAIL.n71 VTAIL.n66 5.81868
R501 VTAIL.n123 VTAIL.n118 5.81868
R502 VTAIL.n329 VTAIL.n324 5.81868
R503 VTAIL.n277 VTAIL.n272 5.81868
R504 VTAIL.n227 VTAIL.n222 5.81868
R505 VTAIL.n175 VTAIL.n170 5.81868
R506 VTAIL.n378 VTAIL.n370 5.04292
R507 VTAIL.n22 VTAIL.n14 5.04292
R508 VTAIL.n72 VTAIL.n64 5.04292
R509 VTAIL.n124 VTAIL.n116 5.04292
R510 VTAIL.n330 VTAIL.n322 5.04292
R511 VTAIL.n278 VTAIL.n270 5.04292
R512 VTAIL.n228 VTAIL.n220 5.04292
R513 VTAIL.n176 VTAIL.n168 5.04292
R514 VTAIL.n382 VTAIL.n381 4.26717
R515 VTAIL.n26 VTAIL.n25 4.26717
R516 VTAIL.n76 VTAIL.n75 4.26717
R517 VTAIL.n128 VTAIL.n127 4.26717
R518 VTAIL.n334 VTAIL.n333 4.26717
R519 VTAIL.n282 VTAIL.n281 4.26717
R520 VTAIL.n232 VTAIL.n231 4.26717
R521 VTAIL.n180 VTAIL.n179 4.26717
R522 VTAIL.n385 VTAIL.n368 3.49141
R523 VTAIL.n29 VTAIL.n12 3.49141
R524 VTAIL.n79 VTAIL.n62 3.49141
R525 VTAIL.n131 VTAIL.n114 3.49141
R526 VTAIL.n337 VTAIL.n320 3.49141
R527 VTAIL.n285 VTAIL.n268 3.49141
R528 VTAIL.n235 VTAIL.n218 3.49141
R529 VTAIL.n183 VTAIL.n166 3.49141
R530 VTAIL.n0 VTAIL.t14 3.43292
R531 VTAIL.n0 VTAIL.t10 3.43292
R532 VTAIL.n102 VTAIL.t0 3.43292
R533 VTAIL.n102 VTAIL.t4 3.43292
R534 VTAIL.n306 VTAIL.t3 3.43292
R535 VTAIL.n306 VTAIL.t6 3.43292
R536 VTAIL.n204 VTAIL.t11 3.43292
R537 VTAIL.n204 VTAIL.t9 3.43292
R538 VTAIL.n386 VTAIL.n366 2.71565
R539 VTAIL.n406 VTAIL.n358 2.71565
R540 VTAIL.n30 VTAIL.n10 2.71565
R541 VTAIL.n50 VTAIL.n2 2.71565
R542 VTAIL.n80 VTAIL.n60 2.71565
R543 VTAIL.n100 VTAIL.n52 2.71565
R544 VTAIL.n132 VTAIL.n112 2.71565
R545 VTAIL.n152 VTAIL.n104 2.71565
R546 VTAIL.n356 VTAIL.n308 2.71565
R547 VTAIL.n338 VTAIL.n318 2.71565
R548 VTAIL.n304 VTAIL.n256 2.71565
R549 VTAIL.n286 VTAIL.n266 2.71565
R550 VTAIL.n254 VTAIL.n206 2.71565
R551 VTAIL.n236 VTAIL.n216 2.71565
R552 VTAIL.n202 VTAIL.n154 2.71565
R553 VTAIL.n184 VTAIL.n164 2.71565
R554 VTAIL.n373 VTAIL.n371 2.41283
R555 VTAIL.n17 VTAIL.n15 2.41283
R556 VTAIL.n67 VTAIL.n65 2.41283
R557 VTAIL.n119 VTAIL.n117 2.41283
R558 VTAIL.n325 VTAIL.n323 2.41283
R559 VTAIL.n273 VTAIL.n271 2.41283
R560 VTAIL.n223 VTAIL.n221 2.41283
R561 VTAIL.n171 VTAIL.n169 2.41283
R562 VTAIL.n391 VTAIL.n389 1.93989
R563 VTAIL.n404 VTAIL.n403 1.93989
R564 VTAIL.n35 VTAIL.n33 1.93989
R565 VTAIL.n48 VTAIL.n47 1.93989
R566 VTAIL.n85 VTAIL.n83 1.93989
R567 VTAIL.n98 VTAIL.n97 1.93989
R568 VTAIL.n137 VTAIL.n135 1.93989
R569 VTAIL.n150 VTAIL.n149 1.93989
R570 VTAIL.n354 VTAIL.n353 1.93989
R571 VTAIL.n342 VTAIL.n341 1.93989
R572 VTAIL.n302 VTAIL.n301 1.93989
R573 VTAIL.n290 VTAIL.n289 1.93989
R574 VTAIL.n252 VTAIL.n251 1.93989
R575 VTAIL.n240 VTAIL.n239 1.93989
R576 VTAIL.n200 VTAIL.n199 1.93989
R577 VTAIL.n188 VTAIL.n187 1.93989
R578 VTAIL.n205 VTAIL.n203 1.5005
R579 VTAIL.n255 VTAIL.n205 1.5005
R580 VTAIL.n307 VTAIL.n305 1.5005
R581 VTAIL.n357 VTAIL.n307 1.5005
R582 VTAIL.n153 VTAIL.n103 1.5005
R583 VTAIL.n103 VTAIL.n101 1.5005
R584 VTAIL.n51 VTAIL.n1 1.5005
R585 VTAIL VTAIL.n407 1.44231
R586 VTAIL.n390 VTAIL.n364 1.16414
R587 VTAIL.n400 VTAIL.n360 1.16414
R588 VTAIL.n34 VTAIL.n8 1.16414
R589 VTAIL.n44 VTAIL.n4 1.16414
R590 VTAIL.n84 VTAIL.n58 1.16414
R591 VTAIL.n94 VTAIL.n54 1.16414
R592 VTAIL.n136 VTAIL.n110 1.16414
R593 VTAIL.n146 VTAIL.n106 1.16414
R594 VTAIL.n350 VTAIL.n310 1.16414
R595 VTAIL.n345 VTAIL.n315 1.16414
R596 VTAIL.n298 VTAIL.n258 1.16414
R597 VTAIL.n293 VTAIL.n263 1.16414
R598 VTAIL.n248 VTAIL.n208 1.16414
R599 VTAIL.n243 VTAIL.n213 1.16414
R600 VTAIL.n196 VTAIL.n156 1.16414
R601 VTAIL.n191 VTAIL.n161 1.16414
R602 VTAIL.n305 VTAIL.n255 0.470328
R603 VTAIL.n101 VTAIL.n51 0.470328
R604 VTAIL.n396 VTAIL.n395 0.388379
R605 VTAIL.n399 VTAIL.n362 0.388379
R606 VTAIL.n40 VTAIL.n39 0.388379
R607 VTAIL.n43 VTAIL.n6 0.388379
R608 VTAIL.n90 VTAIL.n89 0.388379
R609 VTAIL.n93 VTAIL.n56 0.388379
R610 VTAIL.n142 VTAIL.n141 0.388379
R611 VTAIL.n145 VTAIL.n108 0.388379
R612 VTAIL.n349 VTAIL.n312 0.388379
R613 VTAIL.n346 VTAIL.n314 0.388379
R614 VTAIL.n297 VTAIL.n260 0.388379
R615 VTAIL.n294 VTAIL.n262 0.388379
R616 VTAIL.n247 VTAIL.n210 0.388379
R617 VTAIL.n244 VTAIL.n212 0.388379
R618 VTAIL.n195 VTAIL.n158 0.388379
R619 VTAIL.n192 VTAIL.n160 0.388379
R620 VTAIL.n379 VTAIL.n371 0.155672
R621 VTAIL.n380 VTAIL.n379 0.155672
R622 VTAIL.n380 VTAIL.n367 0.155672
R623 VTAIL.n387 VTAIL.n367 0.155672
R624 VTAIL.n388 VTAIL.n387 0.155672
R625 VTAIL.n388 VTAIL.n363 0.155672
R626 VTAIL.n397 VTAIL.n363 0.155672
R627 VTAIL.n398 VTAIL.n397 0.155672
R628 VTAIL.n398 VTAIL.n359 0.155672
R629 VTAIL.n405 VTAIL.n359 0.155672
R630 VTAIL.n23 VTAIL.n15 0.155672
R631 VTAIL.n24 VTAIL.n23 0.155672
R632 VTAIL.n24 VTAIL.n11 0.155672
R633 VTAIL.n31 VTAIL.n11 0.155672
R634 VTAIL.n32 VTAIL.n31 0.155672
R635 VTAIL.n32 VTAIL.n7 0.155672
R636 VTAIL.n41 VTAIL.n7 0.155672
R637 VTAIL.n42 VTAIL.n41 0.155672
R638 VTAIL.n42 VTAIL.n3 0.155672
R639 VTAIL.n49 VTAIL.n3 0.155672
R640 VTAIL.n73 VTAIL.n65 0.155672
R641 VTAIL.n74 VTAIL.n73 0.155672
R642 VTAIL.n74 VTAIL.n61 0.155672
R643 VTAIL.n81 VTAIL.n61 0.155672
R644 VTAIL.n82 VTAIL.n81 0.155672
R645 VTAIL.n82 VTAIL.n57 0.155672
R646 VTAIL.n91 VTAIL.n57 0.155672
R647 VTAIL.n92 VTAIL.n91 0.155672
R648 VTAIL.n92 VTAIL.n53 0.155672
R649 VTAIL.n99 VTAIL.n53 0.155672
R650 VTAIL.n125 VTAIL.n117 0.155672
R651 VTAIL.n126 VTAIL.n125 0.155672
R652 VTAIL.n126 VTAIL.n113 0.155672
R653 VTAIL.n133 VTAIL.n113 0.155672
R654 VTAIL.n134 VTAIL.n133 0.155672
R655 VTAIL.n134 VTAIL.n109 0.155672
R656 VTAIL.n143 VTAIL.n109 0.155672
R657 VTAIL.n144 VTAIL.n143 0.155672
R658 VTAIL.n144 VTAIL.n105 0.155672
R659 VTAIL.n151 VTAIL.n105 0.155672
R660 VTAIL.n355 VTAIL.n309 0.155672
R661 VTAIL.n348 VTAIL.n309 0.155672
R662 VTAIL.n348 VTAIL.n347 0.155672
R663 VTAIL.n347 VTAIL.n313 0.155672
R664 VTAIL.n340 VTAIL.n313 0.155672
R665 VTAIL.n340 VTAIL.n339 0.155672
R666 VTAIL.n339 VTAIL.n319 0.155672
R667 VTAIL.n332 VTAIL.n319 0.155672
R668 VTAIL.n332 VTAIL.n331 0.155672
R669 VTAIL.n331 VTAIL.n323 0.155672
R670 VTAIL.n303 VTAIL.n257 0.155672
R671 VTAIL.n296 VTAIL.n257 0.155672
R672 VTAIL.n296 VTAIL.n295 0.155672
R673 VTAIL.n295 VTAIL.n261 0.155672
R674 VTAIL.n288 VTAIL.n261 0.155672
R675 VTAIL.n288 VTAIL.n287 0.155672
R676 VTAIL.n287 VTAIL.n267 0.155672
R677 VTAIL.n280 VTAIL.n267 0.155672
R678 VTAIL.n280 VTAIL.n279 0.155672
R679 VTAIL.n279 VTAIL.n271 0.155672
R680 VTAIL.n253 VTAIL.n207 0.155672
R681 VTAIL.n246 VTAIL.n207 0.155672
R682 VTAIL.n246 VTAIL.n245 0.155672
R683 VTAIL.n245 VTAIL.n211 0.155672
R684 VTAIL.n238 VTAIL.n211 0.155672
R685 VTAIL.n238 VTAIL.n237 0.155672
R686 VTAIL.n237 VTAIL.n217 0.155672
R687 VTAIL.n230 VTAIL.n217 0.155672
R688 VTAIL.n230 VTAIL.n229 0.155672
R689 VTAIL.n229 VTAIL.n221 0.155672
R690 VTAIL.n201 VTAIL.n155 0.155672
R691 VTAIL.n194 VTAIL.n155 0.155672
R692 VTAIL.n194 VTAIL.n193 0.155672
R693 VTAIL.n193 VTAIL.n159 0.155672
R694 VTAIL.n186 VTAIL.n159 0.155672
R695 VTAIL.n186 VTAIL.n185 0.155672
R696 VTAIL.n185 VTAIL.n165 0.155672
R697 VTAIL.n178 VTAIL.n165 0.155672
R698 VTAIL.n178 VTAIL.n177 0.155672
R699 VTAIL.n177 VTAIL.n169 0.155672
R700 VTAIL VTAIL.n1 0.0586897
R701 VP.n11 VP.t1 193.107
R702 VP.n26 VP.n25 180.385
R703 VP.n46 VP.n45 180.385
R704 VP.n24 VP.n23 180.385
R705 VP.n25 VP.t6 161.863
R706 VP.n31 VP.t7 161.863
R707 VP.n38 VP.t2 161.863
R708 VP.n45 VP.t0 161.863
R709 VP.n23 VP.t5 161.863
R710 VP.n16 VP.t3 161.863
R711 VP.n10 VP.t4 161.863
R712 VP.n12 VP.n9 161.3
R713 VP.n14 VP.n13 161.3
R714 VP.n15 VP.n8 161.3
R715 VP.n18 VP.n17 161.3
R716 VP.n19 VP.n7 161.3
R717 VP.n21 VP.n20 161.3
R718 VP.n22 VP.n6 161.3
R719 VP.n44 VP.n0 161.3
R720 VP.n43 VP.n42 161.3
R721 VP.n41 VP.n1 161.3
R722 VP.n40 VP.n39 161.3
R723 VP.n37 VP.n2 161.3
R724 VP.n36 VP.n35 161.3
R725 VP.n34 VP.n3 161.3
R726 VP.n33 VP.n32 161.3
R727 VP.n30 VP.n4 161.3
R728 VP.n29 VP.n28 161.3
R729 VP.n27 VP.n5 161.3
R730 VP.n30 VP.n29 56.5193
R731 VP.n43 VP.n1 56.5193
R732 VP.n21 VP.n7 56.5193
R733 VP.n11 VP.n10 47.8106
R734 VP.n26 VP.n24 43.2429
R735 VP.n36 VP.n3 40.4934
R736 VP.n37 VP.n36 40.4934
R737 VP.n15 VP.n14 40.4934
R738 VP.n14 VP.n9 40.4934
R739 VP.n29 VP.n5 24.4675
R740 VP.n32 VP.n30 24.4675
R741 VP.n39 VP.n1 24.4675
R742 VP.n44 VP.n43 24.4675
R743 VP.n22 VP.n21 24.4675
R744 VP.n17 VP.n7 24.4675
R745 VP.n12 VP.n11 18.2406
R746 VP.n31 VP.n3 18.1061
R747 VP.n38 VP.n37 18.1061
R748 VP.n16 VP.n15 18.1061
R749 VP.n10 VP.n9 18.1061
R750 VP.n32 VP.n31 6.36192
R751 VP.n39 VP.n38 6.36192
R752 VP.n17 VP.n16 6.36192
R753 VP.n25 VP.n5 5.38324
R754 VP.n45 VP.n44 5.38324
R755 VP.n23 VP.n22 5.38324
R756 VP.n13 VP.n12 0.189894
R757 VP.n13 VP.n8 0.189894
R758 VP.n18 VP.n8 0.189894
R759 VP.n19 VP.n18 0.189894
R760 VP.n20 VP.n19 0.189894
R761 VP.n20 VP.n6 0.189894
R762 VP.n24 VP.n6 0.189894
R763 VP.n27 VP.n26 0.189894
R764 VP.n28 VP.n27 0.189894
R765 VP.n28 VP.n4 0.189894
R766 VP.n33 VP.n4 0.189894
R767 VP.n34 VP.n33 0.189894
R768 VP.n35 VP.n34 0.189894
R769 VP.n35 VP.n2 0.189894
R770 VP.n40 VP.n2 0.189894
R771 VP.n41 VP.n40 0.189894
R772 VP.n42 VP.n41 0.189894
R773 VP.n42 VP.n0 0.189894
R774 VP.n46 VP.n0 0.189894
R775 VP VP.n46 0.0516364
R776 VDD1 VDD1.n0 83.8497
R777 VDD1.n3 VDD1.n2 83.736
R778 VDD1.n3 VDD1.n1 83.736
R779 VDD1.n5 VDD1.n4 83.0413
R780 VDD1.n5 VDD1.n3 39.2121
R781 VDD1.n4 VDD1.t4 3.43292
R782 VDD1.n4 VDD1.t2 3.43292
R783 VDD1.n0 VDD1.t6 3.43292
R784 VDD1.n0 VDD1.t3 3.43292
R785 VDD1.n2 VDD1.t5 3.43292
R786 VDD1.n2 VDD1.t7 3.43292
R787 VDD1.n1 VDD1.t1 3.43292
R788 VDD1.n1 VDD1.t0 3.43292
R789 VDD1 VDD1.n5 0.69231
R790 B.n322 B.n321 585
R791 B.n320 B.n97 585
R792 B.n319 B.n318 585
R793 B.n317 B.n98 585
R794 B.n316 B.n315 585
R795 B.n314 B.n99 585
R796 B.n313 B.n312 585
R797 B.n311 B.n100 585
R798 B.n310 B.n309 585
R799 B.n308 B.n101 585
R800 B.n307 B.n306 585
R801 B.n305 B.n102 585
R802 B.n304 B.n303 585
R803 B.n302 B.n103 585
R804 B.n301 B.n300 585
R805 B.n299 B.n104 585
R806 B.n298 B.n297 585
R807 B.n296 B.n105 585
R808 B.n295 B.n294 585
R809 B.n293 B.n106 585
R810 B.n292 B.n291 585
R811 B.n290 B.n107 585
R812 B.n289 B.n288 585
R813 B.n287 B.n108 585
R814 B.n286 B.n285 585
R815 B.n284 B.n109 585
R816 B.n283 B.n282 585
R817 B.n281 B.n110 585
R818 B.n280 B.n279 585
R819 B.n278 B.n111 585
R820 B.n277 B.n276 585
R821 B.n275 B.n112 585
R822 B.n274 B.n273 585
R823 B.n272 B.n113 585
R824 B.n271 B.n270 585
R825 B.n266 B.n114 585
R826 B.n265 B.n264 585
R827 B.n263 B.n115 585
R828 B.n262 B.n261 585
R829 B.n260 B.n116 585
R830 B.n259 B.n258 585
R831 B.n257 B.n117 585
R832 B.n256 B.n255 585
R833 B.n254 B.n118 585
R834 B.n252 B.n251 585
R835 B.n250 B.n121 585
R836 B.n249 B.n248 585
R837 B.n247 B.n122 585
R838 B.n246 B.n245 585
R839 B.n244 B.n123 585
R840 B.n243 B.n242 585
R841 B.n241 B.n124 585
R842 B.n240 B.n239 585
R843 B.n238 B.n125 585
R844 B.n237 B.n236 585
R845 B.n235 B.n126 585
R846 B.n234 B.n233 585
R847 B.n232 B.n127 585
R848 B.n231 B.n230 585
R849 B.n229 B.n128 585
R850 B.n228 B.n227 585
R851 B.n226 B.n129 585
R852 B.n225 B.n224 585
R853 B.n223 B.n130 585
R854 B.n222 B.n221 585
R855 B.n220 B.n131 585
R856 B.n219 B.n218 585
R857 B.n217 B.n132 585
R858 B.n216 B.n215 585
R859 B.n214 B.n133 585
R860 B.n213 B.n212 585
R861 B.n211 B.n134 585
R862 B.n210 B.n209 585
R863 B.n208 B.n135 585
R864 B.n207 B.n206 585
R865 B.n205 B.n136 585
R866 B.n204 B.n203 585
R867 B.n202 B.n137 585
R868 B.n323 B.n96 585
R869 B.n325 B.n324 585
R870 B.n326 B.n95 585
R871 B.n328 B.n327 585
R872 B.n329 B.n94 585
R873 B.n331 B.n330 585
R874 B.n332 B.n93 585
R875 B.n334 B.n333 585
R876 B.n335 B.n92 585
R877 B.n337 B.n336 585
R878 B.n338 B.n91 585
R879 B.n340 B.n339 585
R880 B.n341 B.n90 585
R881 B.n343 B.n342 585
R882 B.n344 B.n89 585
R883 B.n346 B.n345 585
R884 B.n347 B.n88 585
R885 B.n349 B.n348 585
R886 B.n350 B.n87 585
R887 B.n352 B.n351 585
R888 B.n353 B.n86 585
R889 B.n355 B.n354 585
R890 B.n356 B.n85 585
R891 B.n358 B.n357 585
R892 B.n359 B.n84 585
R893 B.n361 B.n360 585
R894 B.n362 B.n83 585
R895 B.n364 B.n363 585
R896 B.n365 B.n82 585
R897 B.n367 B.n366 585
R898 B.n368 B.n81 585
R899 B.n370 B.n369 585
R900 B.n371 B.n80 585
R901 B.n373 B.n372 585
R902 B.n374 B.n79 585
R903 B.n376 B.n375 585
R904 B.n377 B.n78 585
R905 B.n379 B.n378 585
R906 B.n380 B.n77 585
R907 B.n382 B.n381 585
R908 B.n383 B.n76 585
R909 B.n385 B.n384 585
R910 B.n386 B.n75 585
R911 B.n388 B.n387 585
R912 B.n389 B.n74 585
R913 B.n391 B.n390 585
R914 B.n392 B.n73 585
R915 B.n394 B.n393 585
R916 B.n395 B.n72 585
R917 B.n397 B.n396 585
R918 B.n398 B.n71 585
R919 B.n400 B.n399 585
R920 B.n401 B.n70 585
R921 B.n403 B.n402 585
R922 B.n404 B.n69 585
R923 B.n406 B.n405 585
R924 B.n407 B.n68 585
R925 B.n409 B.n408 585
R926 B.n410 B.n67 585
R927 B.n412 B.n411 585
R928 B.n413 B.n66 585
R929 B.n415 B.n414 585
R930 B.n416 B.n65 585
R931 B.n418 B.n417 585
R932 B.n419 B.n64 585
R933 B.n421 B.n420 585
R934 B.n422 B.n63 585
R935 B.n424 B.n423 585
R936 B.n542 B.n541 585
R937 B.n540 B.n19 585
R938 B.n539 B.n538 585
R939 B.n537 B.n20 585
R940 B.n536 B.n535 585
R941 B.n534 B.n21 585
R942 B.n533 B.n532 585
R943 B.n531 B.n22 585
R944 B.n530 B.n529 585
R945 B.n528 B.n23 585
R946 B.n527 B.n526 585
R947 B.n525 B.n24 585
R948 B.n524 B.n523 585
R949 B.n522 B.n25 585
R950 B.n521 B.n520 585
R951 B.n519 B.n26 585
R952 B.n518 B.n517 585
R953 B.n516 B.n27 585
R954 B.n515 B.n514 585
R955 B.n513 B.n28 585
R956 B.n512 B.n511 585
R957 B.n510 B.n29 585
R958 B.n509 B.n508 585
R959 B.n507 B.n30 585
R960 B.n506 B.n505 585
R961 B.n504 B.n31 585
R962 B.n503 B.n502 585
R963 B.n501 B.n32 585
R964 B.n500 B.n499 585
R965 B.n498 B.n33 585
R966 B.n497 B.n496 585
R967 B.n495 B.n34 585
R968 B.n494 B.n493 585
R969 B.n492 B.n35 585
R970 B.n490 B.n489 585
R971 B.n488 B.n38 585
R972 B.n487 B.n486 585
R973 B.n485 B.n39 585
R974 B.n484 B.n483 585
R975 B.n482 B.n40 585
R976 B.n481 B.n480 585
R977 B.n479 B.n41 585
R978 B.n478 B.n477 585
R979 B.n476 B.n42 585
R980 B.n475 B.n474 585
R981 B.n473 B.n43 585
R982 B.n472 B.n471 585
R983 B.n470 B.n47 585
R984 B.n469 B.n468 585
R985 B.n467 B.n48 585
R986 B.n466 B.n465 585
R987 B.n464 B.n49 585
R988 B.n463 B.n462 585
R989 B.n461 B.n50 585
R990 B.n460 B.n459 585
R991 B.n458 B.n51 585
R992 B.n457 B.n456 585
R993 B.n455 B.n52 585
R994 B.n454 B.n453 585
R995 B.n452 B.n53 585
R996 B.n451 B.n450 585
R997 B.n449 B.n54 585
R998 B.n448 B.n447 585
R999 B.n446 B.n55 585
R1000 B.n445 B.n444 585
R1001 B.n443 B.n56 585
R1002 B.n442 B.n441 585
R1003 B.n440 B.n57 585
R1004 B.n439 B.n438 585
R1005 B.n437 B.n58 585
R1006 B.n436 B.n435 585
R1007 B.n434 B.n59 585
R1008 B.n433 B.n432 585
R1009 B.n431 B.n60 585
R1010 B.n430 B.n429 585
R1011 B.n428 B.n61 585
R1012 B.n427 B.n426 585
R1013 B.n425 B.n62 585
R1014 B.n543 B.n18 585
R1015 B.n545 B.n544 585
R1016 B.n546 B.n17 585
R1017 B.n548 B.n547 585
R1018 B.n549 B.n16 585
R1019 B.n551 B.n550 585
R1020 B.n552 B.n15 585
R1021 B.n554 B.n553 585
R1022 B.n555 B.n14 585
R1023 B.n557 B.n556 585
R1024 B.n558 B.n13 585
R1025 B.n560 B.n559 585
R1026 B.n561 B.n12 585
R1027 B.n563 B.n562 585
R1028 B.n564 B.n11 585
R1029 B.n566 B.n565 585
R1030 B.n567 B.n10 585
R1031 B.n569 B.n568 585
R1032 B.n570 B.n9 585
R1033 B.n572 B.n571 585
R1034 B.n573 B.n8 585
R1035 B.n575 B.n574 585
R1036 B.n576 B.n7 585
R1037 B.n578 B.n577 585
R1038 B.n579 B.n6 585
R1039 B.n581 B.n580 585
R1040 B.n582 B.n5 585
R1041 B.n584 B.n583 585
R1042 B.n585 B.n4 585
R1043 B.n587 B.n586 585
R1044 B.n588 B.n3 585
R1045 B.n590 B.n589 585
R1046 B.n591 B.n0 585
R1047 B.n2 B.n1 585
R1048 B.n154 B.n153 585
R1049 B.n156 B.n155 585
R1050 B.n157 B.n152 585
R1051 B.n159 B.n158 585
R1052 B.n160 B.n151 585
R1053 B.n162 B.n161 585
R1054 B.n163 B.n150 585
R1055 B.n165 B.n164 585
R1056 B.n166 B.n149 585
R1057 B.n168 B.n167 585
R1058 B.n169 B.n148 585
R1059 B.n171 B.n170 585
R1060 B.n172 B.n147 585
R1061 B.n174 B.n173 585
R1062 B.n175 B.n146 585
R1063 B.n177 B.n176 585
R1064 B.n178 B.n145 585
R1065 B.n180 B.n179 585
R1066 B.n181 B.n144 585
R1067 B.n183 B.n182 585
R1068 B.n184 B.n143 585
R1069 B.n186 B.n185 585
R1070 B.n187 B.n142 585
R1071 B.n189 B.n188 585
R1072 B.n190 B.n141 585
R1073 B.n192 B.n191 585
R1074 B.n193 B.n140 585
R1075 B.n195 B.n194 585
R1076 B.n196 B.n139 585
R1077 B.n198 B.n197 585
R1078 B.n199 B.n138 585
R1079 B.n201 B.n200 585
R1080 B.n202 B.n201 526.135
R1081 B.n321 B.n96 526.135
R1082 B.n423 B.n62 526.135
R1083 B.n543 B.n542 526.135
R1084 B.n119 B.t0 366.952
R1085 B.n267 B.t9 366.952
R1086 B.n44 B.t6 366.952
R1087 B.n36 B.t3 366.952
R1088 B.n267 B.t10 363.997
R1089 B.n44 B.t8 363.997
R1090 B.n119 B.t1 363.997
R1091 B.n36 B.t5 363.997
R1092 B.n268 B.t11 330.252
R1093 B.n45 B.t7 330.252
R1094 B.n120 B.t2 330.252
R1095 B.n37 B.t4 330.252
R1096 B.n593 B.n592 256.663
R1097 B.n592 B.n591 235.042
R1098 B.n592 B.n2 235.042
R1099 B.n203 B.n202 163.367
R1100 B.n203 B.n136 163.367
R1101 B.n207 B.n136 163.367
R1102 B.n208 B.n207 163.367
R1103 B.n209 B.n208 163.367
R1104 B.n209 B.n134 163.367
R1105 B.n213 B.n134 163.367
R1106 B.n214 B.n213 163.367
R1107 B.n215 B.n214 163.367
R1108 B.n215 B.n132 163.367
R1109 B.n219 B.n132 163.367
R1110 B.n220 B.n219 163.367
R1111 B.n221 B.n220 163.367
R1112 B.n221 B.n130 163.367
R1113 B.n225 B.n130 163.367
R1114 B.n226 B.n225 163.367
R1115 B.n227 B.n226 163.367
R1116 B.n227 B.n128 163.367
R1117 B.n231 B.n128 163.367
R1118 B.n232 B.n231 163.367
R1119 B.n233 B.n232 163.367
R1120 B.n233 B.n126 163.367
R1121 B.n237 B.n126 163.367
R1122 B.n238 B.n237 163.367
R1123 B.n239 B.n238 163.367
R1124 B.n239 B.n124 163.367
R1125 B.n243 B.n124 163.367
R1126 B.n244 B.n243 163.367
R1127 B.n245 B.n244 163.367
R1128 B.n245 B.n122 163.367
R1129 B.n249 B.n122 163.367
R1130 B.n250 B.n249 163.367
R1131 B.n251 B.n250 163.367
R1132 B.n251 B.n118 163.367
R1133 B.n256 B.n118 163.367
R1134 B.n257 B.n256 163.367
R1135 B.n258 B.n257 163.367
R1136 B.n258 B.n116 163.367
R1137 B.n262 B.n116 163.367
R1138 B.n263 B.n262 163.367
R1139 B.n264 B.n263 163.367
R1140 B.n264 B.n114 163.367
R1141 B.n271 B.n114 163.367
R1142 B.n272 B.n271 163.367
R1143 B.n273 B.n272 163.367
R1144 B.n273 B.n112 163.367
R1145 B.n277 B.n112 163.367
R1146 B.n278 B.n277 163.367
R1147 B.n279 B.n278 163.367
R1148 B.n279 B.n110 163.367
R1149 B.n283 B.n110 163.367
R1150 B.n284 B.n283 163.367
R1151 B.n285 B.n284 163.367
R1152 B.n285 B.n108 163.367
R1153 B.n289 B.n108 163.367
R1154 B.n290 B.n289 163.367
R1155 B.n291 B.n290 163.367
R1156 B.n291 B.n106 163.367
R1157 B.n295 B.n106 163.367
R1158 B.n296 B.n295 163.367
R1159 B.n297 B.n296 163.367
R1160 B.n297 B.n104 163.367
R1161 B.n301 B.n104 163.367
R1162 B.n302 B.n301 163.367
R1163 B.n303 B.n302 163.367
R1164 B.n303 B.n102 163.367
R1165 B.n307 B.n102 163.367
R1166 B.n308 B.n307 163.367
R1167 B.n309 B.n308 163.367
R1168 B.n309 B.n100 163.367
R1169 B.n313 B.n100 163.367
R1170 B.n314 B.n313 163.367
R1171 B.n315 B.n314 163.367
R1172 B.n315 B.n98 163.367
R1173 B.n319 B.n98 163.367
R1174 B.n320 B.n319 163.367
R1175 B.n321 B.n320 163.367
R1176 B.n423 B.n422 163.367
R1177 B.n422 B.n421 163.367
R1178 B.n421 B.n64 163.367
R1179 B.n417 B.n64 163.367
R1180 B.n417 B.n416 163.367
R1181 B.n416 B.n415 163.367
R1182 B.n415 B.n66 163.367
R1183 B.n411 B.n66 163.367
R1184 B.n411 B.n410 163.367
R1185 B.n410 B.n409 163.367
R1186 B.n409 B.n68 163.367
R1187 B.n405 B.n68 163.367
R1188 B.n405 B.n404 163.367
R1189 B.n404 B.n403 163.367
R1190 B.n403 B.n70 163.367
R1191 B.n399 B.n70 163.367
R1192 B.n399 B.n398 163.367
R1193 B.n398 B.n397 163.367
R1194 B.n397 B.n72 163.367
R1195 B.n393 B.n72 163.367
R1196 B.n393 B.n392 163.367
R1197 B.n392 B.n391 163.367
R1198 B.n391 B.n74 163.367
R1199 B.n387 B.n74 163.367
R1200 B.n387 B.n386 163.367
R1201 B.n386 B.n385 163.367
R1202 B.n385 B.n76 163.367
R1203 B.n381 B.n76 163.367
R1204 B.n381 B.n380 163.367
R1205 B.n380 B.n379 163.367
R1206 B.n379 B.n78 163.367
R1207 B.n375 B.n78 163.367
R1208 B.n375 B.n374 163.367
R1209 B.n374 B.n373 163.367
R1210 B.n373 B.n80 163.367
R1211 B.n369 B.n80 163.367
R1212 B.n369 B.n368 163.367
R1213 B.n368 B.n367 163.367
R1214 B.n367 B.n82 163.367
R1215 B.n363 B.n82 163.367
R1216 B.n363 B.n362 163.367
R1217 B.n362 B.n361 163.367
R1218 B.n361 B.n84 163.367
R1219 B.n357 B.n84 163.367
R1220 B.n357 B.n356 163.367
R1221 B.n356 B.n355 163.367
R1222 B.n355 B.n86 163.367
R1223 B.n351 B.n86 163.367
R1224 B.n351 B.n350 163.367
R1225 B.n350 B.n349 163.367
R1226 B.n349 B.n88 163.367
R1227 B.n345 B.n88 163.367
R1228 B.n345 B.n344 163.367
R1229 B.n344 B.n343 163.367
R1230 B.n343 B.n90 163.367
R1231 B.n339 B.n90 163.367
R1232 B.n339 B.n338 163.367
R1233 B.n338 B.n337 163.367
R1234 B.n337 B.n92 163.367
R1235 B.n333 B.n92 163.367
R1236 B.n333 B.n332 163.367
R1237 B.n332 B.n331 163.367
R1238 B.n331 B.n94 163.367
R1239 B.n327 B.n94 163.367
R1240 B.n327 B.n326 163.367
R1241 B.n326 B.n325 163.367
R1242 B.n325 B.n96 163.367
R1243 B.n542 B.n19 163.367
R1244 B.n538 B.n19 163.367
R1245 B.n538 B.n537 163.367
R1246 B.n537 B.n536 163.367
R1247 B.n536 B.n21 163.367
R1248 B.n532 B.n21 163.367
R1249 B.n532 B.n531 163.367
R1250 B.n531 B.n530 163.367
R1251 B.n530 B.n23 163.367
R1252 B.n526 B.n23 163.367
R1253 B.n526 B.n525 163.367
R1254 B.n525 B.n524 163.367
R1255 B.n524 B.n25 163.367
R1256 B.n520 B.n25 163.367
R1257 B.n520 B.n519 163.367
R1258 B.n519 B.n518 163.367
R1259 B.n518 B.n27 163.367
R1260 B.n514 B.n27 163.367
R1261 B.n514 B.n513 163.367
R1262 B.n513 B.n512 163.367
R1263 B.n512 B.n29 163.367
R1264 B.n508 B.n29 163.367
R1265 B.n508 B.n507 163.367
R1266 B.n507 B.n506 163.367
R1267 B.n506 B.n31 163.367
R1268 B.n502 B.n31 163.367
R1269 B.n502 B.n501 163.367
R1270 B.n501 B.n500 163.367
R1271 B.n500 B.n33 163.367
R1272 B.n496 B.n33 163.367
R1273 B.n496 B.n495 163.367
R1274 B.n495 B.n494 163.367
R1275 B.n494 B.n35 163.367
R1276 B.n489 B.n35 163.367
R1277 B.n489 B.n488 163.367
R1278 B.n488 B.n487 163.367
R1279 B.n487 B.n39 163.367
R1280 B.n483 B.n39 163.367
R1281 B.n483 B.n482 163.367
R1282 B.n482 B.n481 163.367
R1283 B.n481 B.n41 163.367
R1284 B.n477 B.n41 163.367
R1285 B.n477 B.n476 163.367
R1286 B.n476 B.n475 163.367
R1287 B.n475 B.n43 163.367
R1288 B.n471 B.n43 163.367
R1289 B.n471 B.n470 163.367
R1290 B.n470 B.n469 163.367
R1291 B.n469 B.n48 163.367
R1292 B.n465 B.n48 163.367
R1293 B.n465 B.n464 163.367
R1294 B.n464 B.n463 163.367
R1295 B.n463 B.n50 163.367
R1296 B.n459 B.n50 163.367
R1297 B.n459 B.n458 163.367
R1298 B.n458 B.n457 163.367
R1299 B.n457 B.n52 163.367
R1300 B.n453 B.n52 163.367
R1301 B.n453 B.n452 163.367
R1302 B.n452 B.n451 163.367
R1303 B.n451 B.n54 163.367
R1304 B.n447 B.n54 163.367
R1305 B.n447 B.n446 163.367
R1306 B.n446 B.n445 163.367
R1307 B.n445 B.n56 163.367
R1308 B.n441 B.n56 163.367
R1309 B.n441 B.n440 163.367
R1310 B.n440 B.n439 163.367
R1311 B.n439 B.n58 163.367
R1312 B.n435 B.n58 163.367
R1313 B.n435 B.n434 163.367
R1314 B.n434 B.n433 163.367
R1315 B.n433 B.n60 163.367
R1316 B.n429 B.n60 163.367
R1317 B.n429 B.n428 163.367
R1318 B.n428 B.n427 163.367
R1319 B.n427 B.n62 163.367
R1320 B.n544 B.n543 163.367
R1321 B.n544 B.n17 163.367
R1322 B.n548 B.n17 163.367
R1323 B.n549 B.n548 163.367
R1324 B.n550 B.n549 163.367
R1325 B.n550 B.n15 163.367
R1326 B.n554 B.n15 163.367
R1327 B.n555 B.n554 163.367
R1328 B.n556 B.n555 163.367
R1329 B.n556 B.n13 163.367
R1330 B.n560 B.n13 163.367
R1331 B.n561 B.n560 163.367
R1332 B.n562 B.n561 163.367
R1333 B.n562 B.n11 163.367
R1334 B.n566 B.n11 163.367
R1335 B.n567 B.n566 163.367
R1336 B.n568 B.n567 163.367
R1337 B.n568 B.n9 163.367
R1338 B.n572 B.n9 163.367
R1339 B.n573 B.n572 163.367
R1340 B.n574 B.n573 163.367
R1341 B.n574 B.n7 163.367
R1342 B.n578 B.n7 163.367
R1343 B.n579 B.n578 163.367
R1344 B.n580 B.n579 163.367
R1345 B.n580 B.n5 163.367
R1346 B.n584 B.n5 163.367
R1347 B.n585 B.n584 163.367
R1348 B.n586 B.n585 163.367
R1349 B.n586 B.n3 163.367
R1350 B.n590 B.n3 163.367
R1351 B.n591 B.n590 163.367
R1352 B.n154 B.n2 163.367
R1353 B.n155 B.n154 163.367
R1354 B.n155 B.n152 163.367
R1355 B.n159 B.n152 163.367
R1356 B.n160 B.n159 163.367
R1357 B.n161 B.n160 163.367
R1358 B.n161 B.n150 163.367
R1359 B.n165 B.n150 163.367
R1360 B.n166 B.n165 163.367
R1361 B.n167 B.n166 163.367
R1362 B.n167 B.n148 163.367
R1363 B.n171 B.n148 163.367
R1364 B.n172 B.n171 163.367
R1365 B.n173 B.n172 163.367
R1366 B.n173 B.n146 163.367
R1367 B.n177 B.n146 163.367
R1368 B.n178 B.n177 163.367
R1369 B.n179 B.n178 163.367
R1370 B.n179 B.n144 163.367
R1371 B.n183 B.n144 163.367
R1372 B.n184 B.n183 163.367
R1373 B.n185 B.n184 163.367
R1374 B.n185 B.n142 163.367
R1375 B.n189 B.n142 163.367
R1376 B.n190 B.n189 163.367
R1377 B.n191 B.n190 163.367
R1378 B.n191 B.n140 163.367
R1379 B.n195 B.n140 163.367
R1380 B.n196 B.n195 163.367
R1381 B.n197 B.n196 163.367
R1382 B.n197 B.n138 163.367
R1383 B.n201 B.n138 163.367
R1384 B.n253 B.n120 59.5399
R1385 B.n269 B.n268 59.5399
R1386 B.n46 B.n45 59.5399
R1387 B.n491 B.n37 59.5399
R1388 B.n541 B.n18 34.1859
R1389 B.n425 B.n424 34.1859
R1390 B.n323 B.n322 34.1859
R1391 B.n200 B.n137 34.1859
R1392 B.n120 B.n119 33.746
R1393 B.n268 B.n267 33.746
R1394 B.n45 B.n44 33.746
R1395 B.n37 B.n36 33.746
R1396 B B.n593 18.0485
R1397 B.n545 B.n18 10.6151
R1398 B.n546 B.n545 10.6151
R1399 B.n547 B.n546 10.6151
R1400 B.n547 B.n16 10.6151
R1401 B.n551 B.n16 10.6151
R1402 B.n552 B.n551 10.6151
R1403 B.n553 B.n552 10.6151
R1404 B.n553 B.n14 10.6151
R1405 B.n557 B.n14 10.6151
R1406 B.n558 B.n557 10.6151
R1407 B.n559 B.n558 10.6151
R1408 B.n559 B.n12 10.6151
R1409 B.n563 B.n12 10.6151
R1410 B.n564 B.n563 10.6151
R1411 B.n565 B.n564 10.6151
R1412 B.n565 B.n10 10.6151
R1413 B.n569 B.n10 10.6151
R1414 B.n570 B.n569 10.6151
R1415 B.n571 B.n570 10.6151
R1416 B.n571 B.n8 10.6151
R1417 B.n575 B.n8 10.6151
R1418 B.n576 B.n575 10.6151
R1419 B.n577 B.n576 10.6151
R1420 B.n577 B.n6 10.6151
R1421 B.n581 B.n6 10.6151
R1422 B.n582 B.n581 10.6151
R1423 B.n583 B.n582 10.6151
R1424 B.n583 B.n4 10.6151
R1425 B.n587 B.n4 10.6151
R1426 B.n588 B.n587 10.6151
R1427 B.n589 B.n588 10.6151
R1428 B.n589 B.n0 10.6151
R1429 B.n541 B.n540 10.6151
R1430 B.n540 B.n539 10.6151
R1431 B.n539 B.n20 10.6151
R1432 B.n535 B.n20 10.6151
R1433 B.n535 B.n534 10.6151
R1434 B.n534 B.n533 10.6151
R1435 B.n533 B.n22 10.6151
R1436 B.n529 B.n22 10.6151
R1437 B.n529 B.n528 10.6151
R1438 B.n528 B.n527 10.6151
R1439 B.n527 B.n24 10.6151
R1440 B.n523 B.n24 10.6151
R1441 B.n523 B.n522 10.6151
R1442 B.n522 B.n521 10.6151
R1443 B.n521 B.n26 10.6151
R1444 B.n517 B.n26 10.6151
R1445 B.n517 B.n516 10.6151
R1446 B.n516 B.n515 10.6151
R1447 B.n515 B.n28 10.6151
R1448 B.n511 B.n28 10.6151
R1449 B.n511 B.n510 10.6151
R1450 B.n510 B.n509 10.6151
R1451 B.n509 B.n30 10.6151
R1452 B.n505 B.n30 10.6151
R1453 B.n505 B.n504 10.6151
R1454 B.n504 B.n503 10.6151
R1455 B.n503 B.n32 10.6151
R1456 B.n499 B.n32 10.6151
R1457 B.n499 B.n498 10.6151
R1458 B.n498 B.n497 10.6151
R1459 B.n497 B.n34 10.6151
R1460 B.n493 B.n34 10.6151
R1461 B.n493 B.n492 10.6151
R1462 B.n490 B.n38 10.6151
R1463 B.n486 B.n38 10.6151
R1464 B.n486 B.n485 10.6151
R1465 B.n485 B.n484 10.6151
R1466 B.n484 B.n40 10.6151
R1467 B.n480 B.n40 10.6151
R1468 B.n480 B.n479 10.6151
R1469 B.n479 B.n478 10.6151
R1470 B.n478 B.n42 10.6151
R1471 B.n474 B.n473 10.6151
R1472 B.n473 B.n472 10.6151
R1473 B.n472 B.n47 10.6151
R1474 B.n468 B.n47 10.6151
R1475 B.n468 B.n467 10.6151
R1476 B.n467 B.n466 10.6151
R1477 B.n466 B.n49 10.6151
R1478 B.n462 B.n49 10.6151
R1479 B.n462 B.n461 10.6151
R1480 B.n461 B.n460 10.6151
R1481 B.n460 B.n51 10.6151
R1482 B.n456 B.n51 10.6151
R1483 B.n456 B.n455 10.6151
R1484 B.n455 B.n454 10.6151
R1485 B.n454 B.n53 10.6151
R1486 B.n450 B.n53 10.6151
R1487 B.n450 B.n449 10.6151
R1488 B.n449 B.n448 10.6151
R1489 B.n448 B.n55 10.6151
R1490 B.n444 B.n55 10.6151
R1491 B.n444 B.n443 10.6151
R1492 B.n443 B.n442 10.6151
R1493 B.n442 B.n57 10.6151
R1494 B.n438 B.n57 10.6151
R1495 B.n438 B.n437 10.6151
R1496 B.n437 B.n436 10.6151
R1497 B.n436 B.n59 10.6151
R1498 B.n432 B.n59 10.6151
R1499 B.n432 B.n431 10.6151
R1500 B.n431 B.n430 10.6151
R1501 B.n430 B.n61 10.6151
R1502 B.n426 B.n61 10.6151
R1503 B.n426 B.n425 10.6151
R1504 B.n424 B.n63 10.6151
R1505 B.n420 B.n63 10.6151
R1506 B.n420 B.n419 10.6151
R1507 B.n419 B.n418 10.6151
R1508 B.n418 B.n65 10.6151
R1509 B.n414 B.n65 10.6151
R1510 B.n414 B.n413 10.6151
R1511 B.n413 B.n412 10.6151
R1512 B.n412 B.n67 10.6151
R1513 B.n408 B.n67 10.6151
R1514 B.n408 B.n407 10.6151
R1515 B.n407 B.n406 10.6151
R1516 B.n406 B.n69 10.6151
R1517 B.n402 B.n69 10.6151
R1518 B.n402 B.n401 10.6151
R1519 B.n401 B.n400 10.6151
R1520 B.n400 B.n71 10.6151
R1521 B.n396 B.n71 10.6151
R1522 B.n396 B.n395 10.6151
R1523 B.n395 B.n394 10.6151
R1524 B.n394 B.n73 10.6151
R1525 B.n390 B.n73 10.6151
R1526 B.n390 B.n389 10.6151
R1527 B.n389 B.n388 10.6151
R1528 B.n388 B.n75 10.6151
R1529 B.n384 B.n75 10.6151
R1530 B.n384 B.n383 10.6151
R1531 B.n383 B.n382 10.6151
R1532 B.n382 B.n77 10.6151
R1533 B.n378 B.n77 10.6151
R1534 B.n378 B.n377 10.6151
R1535 B.n377 B.n376 10.6151
R1536 B.n376 B.n79 10.6151
R1537 B.n372 B.n79 10.6151
R1538 B.n372 B.n371 10.6151
R1539 B.n371 B.n370 10.6151
R1540 B.n370 B.n81 10.6151
R1541 B.n366 B.n81 10.6151
R1542 B.n366 B.n365 10.6151
R1543 B.n365 B.n364 10.6151
R1544 B.n364 B.n83 10.6151
R1545 B.n360 B.n83 10.6151
R1546 B.n360 B.n359 10.6151
R1547 B.n359 B.n358 10.6151
R1548 B.n358 B.n85 10.6151
R1549 B.n354 B.n85 10.6151
R1550 B.n354 B.n353 10.6151
R1551 B.n353 B.n352 10.6151
R1552 B.n352 B.n87 10.6151
R1553 B.n348 B.n87 10.6151
R1554 B.n348 B.n347 10.6151
R1555 B.n347 B.n346 10.6151
R1556 B.n346 B.n89 10.6151
R1557 B.n342 B.n89 10.6151
R1558 B.n342 B.n341 10.6151
R1559 B.n341 B.n340 10.6151
R1560 B.n340 B.n91 10.6151
R1561 B.n336 B.n91 10.6151
R1562 B.n336 B.n335 10.6151
R1563 B.n335 B.n334 10.6151
R1564 B.n334 B.n93 10.6151
R1565 B.n330 B.n93 10.6151
R1566 B.n330 B.n329 10.6151
R1567 B.n329 B.n328 10.6151
R1568 B.n328 B.n95 10.6151
R1569 B.n324 B.n95 10.6151
R1570 B.n324 B.n323 10.6151
R1571 B.n153 B.n1 10.6151
R1572 B.n156 B.n153 10.6151
R1573 B.n157 B.n156 10.6151
R1574 B.n158 B.n157 10.6151
R1575 B.n158 B.n151 10.6151
R1576 B.n162 B.n151 10.6151
R1577 B.n163 B.n162 10.6151
R1578 B.n164 B.n163 10.6151
R1579 B.n164 B.n149 10.6151
R1580 B.n168 B.n149 10.6151
R1581 B.n169 B.n168 10.6151
R1582 B.n170 B.n169 10.6151
R1583 B.n170 B.n147 10.6151
R1584 B.n174 B.n147 10.6151
R1585 B.n175 B.n174 10.6151
R1586 B.n176 B.n175 10.6151
R1587 B.n176 B.n145 10.6151
R1588 B.n180 B.n145 10.6151
R1589 B.n181 B.n180 10.6151
R1590 B.n182 B.n181 10.6151
R1591 B.n182 B.n143 10.6151
R1592 B.n186 B.n143 10.6151
R1593 B.n187 B.n186 10.6151
R1594 B.n188 B.n187 10.6151
R1595 B.n188 B.n141 10.6151
R1596 B.n192 B.n141 10.6151
R1597 B.n193 B.n192 10.6151
R1598 B.n194 B.n193 10.6151
R1599 B.n194 B.n139 10.6151
R1600 B.n198 B.n139 10.6151
R1601 B.n199 B.n198 10.6151
R1602 B.n200 B.n199 10.6151
R1603 B.n204 B.n137 10.6151
R1604 B.n205 B.n204 10.6151
R1605 B.n206 B.n205 10.6151
R1606 B.n206 B.n135 10.6151
R1607 B.n210 B.n135 10.6151
R1608 B.n211 B.n210 10.6151
R1609 B.n212 B.n211 10.6151
R1610 B.n212 B.n133 10.6151
R1611 B.n216 B.n133 10.6151
R1612 B.n217 B.n216 10.6151
R1613 B.n218 B.n217 10.6151
R1614 B.n218 B.n131 10.6151
R1615 B.n222 B.n131 10.6151
R1616 B.n223 B.n222 10.6151
R1617 B.n224 B.n223 10.6151
R1618 B.n224 B.n129 10.6151
R1619 B.n228 B.n129 10.6151
R1620 B.n229 B.n228 10.6151
R1621 B.n230 B.n229 10.6151
R1622 B.n230 B.n127 10.6151
R1623 B.n234 B.n127 10.6151
R1624 B.n235 B.n234 10.6151
R1625 B.n236 B.n235 10.6151
R1626 B.n236 B.n125 10.6151
R1627 B.n240 B.n125 10.6151
R1628 B.n241 B.n240 10.6151
R1629 B.n242 B.n241 10.6151
R1630 B.n242 B.n123 10.6151
R1631 B.n246 B.n123 10.6151
R1632 B.n247 B.n246 10.6151
R1633 B.n248 B.n247 10.6151
R1634 B.n248 B.n121 10.6151
R1635 B.n252 B.n121 10.6151
R1636 B.n255 B.n254 10.6151
R1637 B.n255 B.n117 10.6151
R1638 B.n259 B.n117 10.6151
R1639 B.n260 B.n259 10.6151
R1640 B.n261 B.n260 10.6151
R1641 B.n261 B.n115 10.6151
R1642 B.n265 B.n115 10.6151
R1643 B.n266 B.n265 10.6151
R1644 B.n270 B.n266 10.6151
R1645 B.n274 B.n113 10.6151
R1646 B.n275 B.n274 10.6151
R1647 B.n276 B.n275 10.6151
R1648 B.n276 B.n111 10.6151
R1649 B.n280 B.n111 10.6151
R1650 B.n281 B.n280 10.6151
R1651 B.n282 B.n281 10.6151
R1652 B.n282 B.n109 10.6151
R1653 B.n286 B.n109 10.6151
R1654 B.n287 B.n286 10.6151
R1655 B.n288 B.n287 10.6151
R1656 B.n288 B.n107 10.6151
R1657 B.n292 B.n107 10.6151
R1658 B.n293 B.n292 10.6151
R1659 B.n294 B.n293 10.6151
R1660 B.n294 B.n105 10.6151
R1661 B.n298 B.n105 10.6151
R1662 B.n299 B.n298 10.6151
R1663 B.n300 B.n299 10.6151
R1664 B.n300 B.n103 10.6151
R1665 B.n304 B.n103 10.6151
R1666 B.n305 B.n304 10.6151
R1667 B.n306 B.n305 10.6151
R1668 B.n306 B.n101 10.6151
R1669 B.n310 B.n101 10.6151
R1670 B.n311 B.n310 10.6151
R1671 B.n312 B.n311 10.6151
R1672 B.n312 B.n99 10.6151
R1673 B.n316 B.n99 10.6151
R1674 B.n317 B.n316 10.6151
R1675 B.n318 B.n317 10.6151
R1676 B.n318 B.n97 10.6151
R1677 B.n322 B.n97 10.6151
R1678 B.n492 B.n491 9.36635
R1679 B.n474 B.n46 9.36635
R1680 B.n253 B.n252 9.36635
R1681 B.n269 B.n113 9.36635
R1682 B.n593 B.n0 8.11757
R1683 B.n593 B.n1 8.11757
R1684 B.n491 B.n490 1.24928
R1685 B.n46 B.n42 1.24928
R1686 B.n254 B.n253 1.24928
R1687 B.n270 B.n269 1.24928
C0 B VDD2 1.27757f
C1 VP VDD2 0.393108f
C2 VN B 0.918389f
C3 B VTAIL 3.59357f
C4 VDD2 VDD1 1.18364f
C5 VN VP 5.74292f
C6 VTAIL VP 6.06918f
C7 VN VDD1 0.149642f
C8 VTAIL VDD1 7.37875f
C9 B w_n2710_n2862# 7.583601f
C10 VN VDD2 5.93258f
C11 VTAIL VDD2 7.42519f
C12 w_n2710_n2862# VP 5.4949f
C13 VN VTAIL 6.055069f
C14 w_n2710_n2862# VDD1 1.49437f
C15 w_n2710_n2862# VDD2 1.55912f
C16 B VP 1.49593f
C17 VN w_n2710_n2862# 5.1466f
C18 B VDD1 1.21889f
C19 w_n2710_n2862# VTAIL 3.55057f
C20 VP VDD1 6.17525f
C21 VDD2 VSUBS 1.370188f
C22 VDD1 VSUBS 1.811024f
C23 VTAIL VSUBS 0.98134f
C24 VN VSUBS 5.15306f
C25 VP VSUBS 2.259554f
C26 B VSUBS 3.461919f
C27 w_n2710_n2862# VSUBS 95.9015f
C28 B.n0 VSUBS 0.006943f
C29 B.n1 VSUBS 0.006943f
C30 B.n2 VSUBS 0.010269f
C31 B.n3 VSUBS 0.007869f
C32 B.n4 VSUBS 0.007869f
C33 B.n5 VSUBS 0.007869f
C34 B.n6 VSUBS 0.007869f
C35 B.n7 VSUBS 0.007869f
C36 B.n8 VSUBS 0.007869f
C37 B.n9 VSUBS 0.007869f
C38 B.n10 VSUBS 0.007869f
C39 B.n11 VSUBS 0.007869f
C40 B.n12 VSUBS 0.007869f
C41 B.n13 VSUBS 0.007869f
C42 B.n14 VSUBS 0.007869f
C43 B.n15 VSUBS 0.007869f
C44 B.n16 VSUBS 0.007869f
C45 B.n17 VSUBS 0.007869f
C46 B.n18 VSUBS 0.018383f
C47 B.n19 VSUBS 0.007869f
C48 B.n20 VSUBS 0.007869f
C49 B.n21 VSUBS 0.007869f
C50 B.n22 VSUBS 0.007869f
C51 B.n23 VSUBS 0.007869f
C52 B.n24 VSUBS 0.007869f
C53 B.n25 VSUBS 0.007869f
C54 B.n26 VSUBS 0.007869f
C55 B.n27 VSUBS 0.007869f
C56 B.n28 VSUBS 0.007869f
C57 B.n29 VSUBS 0.007869f
C58 B.n30 VSUBS 0.007869f
C59 B.n31 VSUBS 0.007869f
C60 B.n32 VSUBS 0.007869f
C61 B.n33 VSUBS 0.007869f
C62 B.n34 VSUBS 0.007869f
C63 B.n35 VSUBS 0.007869f
C64 B.t4 VSUBS 0.176063f
C65 B.t5 VSUBS 0.196892f
C66 B.t3 VSUBS 0.664247f
C67 B.n36 VSUBS 0.315725f
C68 B.n37 VSUBS 0.2359f
C69 B.n38 VSUBS 0.007869f
C70 B.n39 VSUBS 0.007869f
C71 B.n40 VSUBS 0.007869f
C72 B.n41 VSUBS 0.007869f
C73 B.n42 VSUBS 0.004398f
C74 B.n43 VSUBS 0.007869f
C75 B.t7 VSUBS 0.176066f
C76 B.t8 VSUBS 0.196895f
C77 B.t6 VSUBS 0.664247f
C78 B.n44 VSUBS 0.315723f
C79 B.n45 VSUBS 0.235897f
C80 B.n46 VSUBS 0.018232f
C81 B.n47 VSUBS 0.007869f
C82 B.n48 VSUBS 0.007869f
C83 B.n49 VSUBS 0.007869f
C84 B.n50 VSUBS 0.007869f
C85 B.n51 VSUBS 0.007869f
C86 B.n52 VSUBS 0.007869f
C87 B.n53 VSUBS 0.007869f
C88 B.n54 VSUBS 0.007869f
C89 B.n55 VSUBS 0.007869f
C90 B.n56 VSUBS 0.007869f
C91 B.n57 VSUBS 0.007869f
C92 B.n58 VSUBS 0.007869f
C93 B.n59 VSUBS 0.007869f
C94 B.n60 VSUBS 0.007869f
C95 B.n61 VSUBS 0.007869f
C96 B.n62 VSUBS 0.019575f
C97 B.n63 VSUBS 0.007869f
C98 B.n64 VSUBS 0.007869f
C99 B.n65 VSUBS 0.007869f
C100 B.n66 VSUBS 0.007869f
C101 B.n67 VSUBS 0.007869f
C102 B.n68 VSUBS 0.007869f
C103 B.n69 VSUBS 0.007869f
C104 B.n70 VSUBS 0.007869f
C105 B.n71 VSUBS 0.007869f
C106 B.n72 VSUBS 0.007869f
C107 B.n73 VSUBS 0.007869f
C108 B.n74 VSUBS 0.007869f
C109 B.n75 VSUBS 0.007869f
C110 B.n76 VSUBS 0.007869f
C111 B.n77 VSUBS 0.007869f
C112 B.n78 VSUBS 0.007869f
C113 B.n79 VSUBS 0.007869f
C114 B.n80 VSUBS 0.007869f
C115 B.n81 VSUBS 0.007869f
C116 B.n82 VSUBS 0.007869f
C117 B.n83 VSUBS 0.007869f
C118 B.n84 VSUBS 0.007869f
C119 B.n85 VSUBS 0.007869f
C120 B.n86 VSUBS 0.007869f
C121 B.n87 VSUBS 0.007869f
C122 B.n88 VSUBS 0.007869f
C123 B.n89 VSUBS 0.007869f
C124 B.n90 VSUBS 0.007869f
C125 B.n91 VSUBS 0.007869f
C126 B.n92 VSUBS 0.007869f
C127 B.n93 VSUBS 0.007869f
C128 B.n94 VSUBS 0.007869f
C129 B.n95 VSUBS 0.007869f
C130 B.n96 VSUBS 0.018383f
C131 B.n97 VSUBS 0.007869f
C132 B.n98 VSUBS 0.007869f
C133 B.n99 VSUBS 0.007869f
C134 B.n100 VSUBS 0.007869f
C135 B.n101 VSUBS 0.007869f
C136 B.n102 VSUBS 0.007869f
C137 B.n103 VSUBS 0.007869f
C138 B.n104 VSUBS 0.007869f
C139 B.n105 VSUBS 0.007869f
C140 B.n106 VSUBS 0.007869f
C141 B.n107 VSUBS 0.007869f
C142 B.n108 VSUBS 0.007869f
C143 B.n109 VSUBS 0.007869f
C144 B.n110 VSUBS 0.007869f
C145 B.n111 VSUBS 0.007869f
C146 B.n112 VSUBS 0.007869f
C147 B.n113 VSUBS 0.007406f
C148 B.n114 VSUBS 0.007869f
C149 B.n115 VSUBS 0.007869f
C150 B.n116 VSUBS 0.007869f
C151 B.n117 VSUBS 0.007869f
C152 B.n118 VSUBS 0.007869f
C153 B.t2 VSUBS 0.176063f
C154 B.t1 VSUBS 0.196892f
C155 B.t0 VSUBS 0.664247f
C156 B.n119 VSUBS 0.315725f
C157 B.n120 VSUBS 0.2359f
C158 B.n121 VSUBS 0.007869f
C159 B.n122 VSUBS 0.007869f
C160 B.n123 VSUBS 0.007869f
C161 B.n124 VSUBS 0.007869f
C162 B.n125 VSUBS 0.007869f
C163 B.n126 VSUBS 0.007869f
C164 B.n127 VSUBS 0.007869f
C165 B.n128 VSUBS 0.007869f
C166 B.n129 VSUBS 0.007869f
C167 B.n130 VSUBS 0.007869f
C168 B.n131 VSUBS 0.007869f
C169 B.n132 VSUBS 0.007869f
C170 B.n133 VSUBS 0.007869f
C171 B.n134 VSUBS 0.007869f
C172 B.n135 VSUBS 0.007869f
C173 B.n136 VSUBS 0.007869f
C174 B.n137 VSUBS 0.019575f
C175 B.n138 VSUBS 0.007869f
C176 B.n139 VSUBS 0.007869f
C177 B.n140 VSUBS 0.007869f
C178 B.n141 VSUBS 0.007869f
C179 B.n142 VSUBS 0.007869f
C180 B.n143 VSUBS 0.007869f
C181 B.n144 VSUBS 0.007869f
C182 B.n145 VSUBS 0.007869f
C183 B.n146 VSUBS 0.007869f
C184 B.n147 VSUBS 0.007869f
C185 B.n148 VSUBS 0.007869f
C186 B.n149 VSUBS 0.007869f
C187 B.n150 VSUBS 0.007869f
C188 B.n151 VSUBS 0.007869f
C189 B.n152 VSUBS 0.007869f
C190 B.n153 VSUBS 0.007869f
C191 B.n154 VSUBS 0.007869f
C192 B.n155 VSUBS 0.007869f
C193 B.n156 VSUBS 0.007869f
C194 B.n157 VSUBS 0.007869f
C195 B.n158 VSUBS 0.007869f
C196 B.n159 VSUBS 0.007869f
C197 B.n160 VSUBS 0.007869f
C198 B.n161 VSUBS 0.007869f
C199 B.n162 VSUBS 0.007869f
C200 B.n163 VSUBS 0.007869f
C201 B.n164 VSUBS 0.007869f
C202 B.n165 VSUBS 0.007869f
C203 B.n166 VSUBS 0.007869f
C204 B.n167 VSUBS 0.007869f
C205 B.n168 VSUBS 0.007869f
C206 B.n169 VSUBS 0.007869f
C207 B.n170 VSUBS 0.007869f
C208 B.n171 VSUBS 0.007869f
C209 B.n172 VSUBS 0.007869f
C210 B.n173 VSUBS 0.007869f
C211 B.n174 VSUBS 0.007869f
C212 B.n175 VSUBS 0.007869f
C213 B.n176 VSUBS 0.007869f
C214 B.n177 VSUBS 0.007869f
C215 B.n178 VSUBS 0.007869f
C216 B.n179 VSUBS 0.007869f
C217 B.n180 VSUBS 0.007869f
C218 B.n181 VSUBS 0.007869f
C219 B.n182 VSUBS 0.007869f
C220 B.n183 VSUBS 0.007869f
C221 B.n184 VSUBS 0.007869f
C222 B.n185 VSUBS 0.007869f
C223 B.n186 VSUBS 0.007869f
C224 B.n187 VSUBS 0.007869f
C225 B.n188 VSUBS 0.007869f
C226 B.n189 VSUBS 0.007869f
C227 B.n190 VSUBS 0.007869f
C228 B.n191 VSUBS 0.007869f
C229 B.n192 VSUBS 0.007869f
C230 B.n193 VSUBS 0.007869f
C231 B.n194 VSUBS 0.007869f
C232 B.n195 VSUBS 0.007869f
C233 B.n196 VSUBS 0.007869f
C234 B.n197 VSUBS 0.007869f
C235 B.n198 VSUBS 0.007869f
C236 B.n199 VSUBS 0.007869f
C237 B.n200 VSUBS 0.018383f
C238 B.n201 VSUBS 0.018383f
C239 B.n202 VSUBS 0.019575f
C240 B.n203 VSUBS 0.007869f
C241 B.n204 VSUBS 0.007869f
C242 B.n205 VSUBS 0.007869f
C243 B.n206 VSUBS 0.007869f
C244 B.n207 VSUBS 0.007869f
C245 B.n208 VSUBS 0.007869f
C246 B.n209 VSUBS 0.007869f
C247 B.n210 VSUBS 0.007869f
C248 B.n211 VSUBS 0.007869f
C249 B.n212 VSUBS 0.007869f
C250 B.n213 VSUBS 0.007869f
C251 B.n214 VSUBS 0.007869f
C252 B.n215 VSUBS 0.007869f
C253 B.n216 VSUBS 0.007869f
C254 B.n217 VSUBS 0.007869f
C255 B.n218 VSUBS 0.007869f
C256 B.n219 VSUBS 0.007869f
C257 B.n220 VSUBS 0.007869f
C258 B.n221 VSUBS 0.007869f
C259 B.n222 VSUBS 0.007869f
C260 B.n223 VSUBS 0.007869f
C261 B.n224 VSUBS 0.007869f
C262 B.n225 VSUBS 0.007869f
C263 B.n226 VSUBS 0.007869f
C264 B.n227 VSUBS 0.007869f
C265 B.n228 VSUBS 0.007869f
C266 B.n229 VSUBS 0.007869f
C267 B.n230 VSUBS 0.007869f
C268 B.n231 VSUBS 0.007869f
C269 B.n232 VSUBS 0.007869f
C270 B.n233 VSUBS 0.007869f
C271 B.n234 VSUBS 0.007869f
C272 B.n235 VSUBS 0.007869f
C273 B.n236 VSUBS 0.007869f
C274 B.n237 VSUBS 0.007869f
C275 B.n238 VSUBS 0.007869f
C276 B.n239 VSUBS 0.007869f
C277 B.n240 VSUBS 0.007869f
C278 B.n241 VSUBS 0.007869f
C279 B.n242 VSUBS 0.007869f
C280 B.n243 VSUBS 0.007869f
C281 B.n244 VSUBS 0.007869f
C282 B.n245 VSUBS 0.007869f
C283 B.n246 VSUBS 0.007869f
C284 B.n247 VSUBS 0.007869f
C285 B.n248 VSUBS 0.007869f
C286 B.n249 VSUBS 0.007869f
C287 B.n250 VSUBS 0.007869f
C288 B.n251 VSUBS 0.007869f
C289 B.n252 VSUBS 0.007406f
C290 B.n253 VSUBS 0.018232f
C291 B.n254 VSUBS 0.004398f
C292 B.n255 VSUBS 0.007869f
C293 B.n256 VSUBS 0.007869f
C294 B.n257 VSUBS 0.007869f
C295 B.n258 VSUBS 0.007869f
C296 B.n259 VSUBS 0.007869f
C297 B.n260 VSUBS 0.007869f
C298 B.n261 VSUBS 0.007869f
C299 B.n262 VSUBS 0.007869f
C300 B.n263 VSUBS 0.007869f
C301 B.n264 VSUBS 0.007869f
C302 B.n265 VSUBS 0.007869f
C303 B.n266 VSUBS 0.007869f
C304 B.t11 VSUBS 0.176066f
C305 B.t10 VSUBS 0.196895f
C306 B.t9 VSUBS 0.664247f
C307 B.n267 VSUBS 0.315723f
C308 B.n268 VSUBS 0.235897f
C309 B.n269 VSUBS 0.018232f
C310 B.n270 VSUBS 0.004398f
C311 B.n271 VSUBS 0.007869f
C312 B.n272 VSUBS 0.007869f
C313 B.n273 VSUBS 0.007869f
C314 B.n274 VSUBS 0.007869f
C315 B.n275 VSUBS 0.007869f
C316 B.n276 VSUBS 0.007869f
C317 B.n277 VSUBS 0.007869f
C318 B.n278 VSUBS 0.007869f
C319 B.n279 VSUBS 0.007869f
C320 B.n280 VSUBS 0.007869f
C321 B.n281 VSUBS 0.007869f
C322 B.n282 VSUBS 0.007869f
C323 B.n283 VSUBS 0.007869f
C324 B.n284 VSUBS 0.007869f
C325 B.n285 VSUBS 0.007869f
C326 B.n286 VSUBS 0.007869f
C327 B.n287 VSUBS 0.007869f
C328 B.n288 VSUBS 0.007869f
C329 B.n289 VSUBS 0.007869f
C330 B.n290 VSUBS 0.007869f
C331 B.n291 VSUBS 0.007869f
C332 B.n292 VSUBS 0.007869f
C333 B.n293 VSUBS 0.007869f
C334 B.n294 VSUBS 0.007869f
C335 B.n295 VSUBS 0.007869f
C336 B.n296 VSUBS 0.007869f
C337 B.n297 VSUBS 0.007869f
C338 B.n298 VSUBS 0.007869f
C339 B.n299 VSUBS 0.007869f
C340 B.n300 VSUBS 0.007869f
C341 B.n301 VSUBS 0.007869f
C342 B.n302 VSUBS 0.007869f
C343 B.n303 VSUBS 0.007869f
C344 B.n304 VSUBS 0.007869f
C345 B.n305 VSUBS 0.007869f
C346 B.n306 VSUBS 0.007869f
C347 B.n307 VSUBS 0.007869f
C348 B.n308 VSUBS 0.007869f
C349 B.n309 VSUBS 0.007869f
C350 B.n310 VSUBS 0.007869f
C351 B.n311 VSUBS 0.007869f
C352 B.n312 VSUBS 0.007869f
C353 B.n313 VSUBS 0.007869f
C354 B.n314 VSUBS 0.007869f
C355 B.n315 VSUBS 0.007869f
C356 B.n316 VSUBS 0.007869f
C357 B.n317 VSUBS 0.007869f
C358 B.n318 VSUBS 0.007869f
C359 B.n319 VSUBS 0.007869f
C360 B.n320 VSUBS 0.007869f
C361 B.n321 VSUBS 0.019575f
C362 B.n322 VSUBS 0.018686f
C363 B.n323 VSUBS 0.019271f
C364 B.n324 VSUBS 0.007869f
C365 B.n325 VSUBS 0.007869f
C366 B.n326 VSUBS 0.007869f
C367 B.n327 VSUBS 0.007869f
C368 B.n328 VSUBS 0.007869f
C369 B.n329 VSUBS 0.007869f
C370 B.n330 VSUBS 0.007869f
C371 B.n331 VSUBS 0.007869f
C372 B.n332 VSUBS 0.007869f
C373 B.n333 VSUBS 0.007869f
C374 B.n334 VSUBS 0.007869f
C375 B.n335 VSUBS 0.007869f
C376 B.n336 VSUBS 0.007869f
C377 B.n337 VSUBS 0.007869f
C378 B.n338 VSUBS 0.007869f
C379 B.n339 VSUBS 0.007869f
C380 B.n340 VSUBS 0.007869f
C381 B.n341 VSUBS 0.007869f
C382 B.n342 VSUBS 0.007869f
C383 B.n343 VSUBS 0.007869f
C384 B.n344 VSUBS 0.007869f
C385 B.n345 VSUBS 0.007869f
C386 B.n346 VSUBS 0.007869f
C387 B.n347 VSUBS 0.007869f
C388 B.n348 VSUBS 0.007869f
C389 B.n349 VSUBS 0.007869f
C390 B.n350 VSUBS 0.007869f
C391 B.n351 VSUBS 0.007869f
C392 B.n352 VSUBS 0.007869f
C393 B.n353 VSUBS 0.007869f
C394 B.n354 VSUBS 0.007869f
C395 B.n355 VSUBS 0.007869f
C396 B.n356 VSUBS 0.007869f
C397 B.n357 VSUBS 0.007869f
C398 B.n358 VSUBS 0.007869f
C399 B.n359 VSUBS 0.007869f
C400 B.n360 VSUBS 0.007869f
C401 B.n361 VSUBS 0.007869f
C402 B.n362 VSUBS 0.007869f
C403 B.n363 VSUBS 0.007869f
C404 B.n364 VSUBS 0.007869f
C405 B.n365 VSUBS 0.007869f
C406 B.n366 VSUBS 0.007869f
C407 B.n367 VSUBS 0.007869f
C408 B.n368 VSUBS 0.007869f
C409 B.n369 VSUBS 0.007869f
C410 B.n370 VSUBS 0.007869f
C411 B.n371 VSUBS 0.007869f
C412 B.n372 VSUBS 0.007869f
C413 B.n373 VSUBS 0.007869f
C414 B.n374 VSUBS 0.007869f
C415 B.n375 VSUBS 0.007869f
C416 B.n376 VSUBS 0.007869f
C417 B.n377 VSUBS 0.007869f
C418 B.n378 VSUBS 0.007869f
C419 B.n379 VSUBS 0.007869f
C420 B.n380 VSUBS 0.007869f
C421 B.n381 VSUBS 0.007869f
C422 B.n382 VSUBS 0.007869f
C423 B.n383 VSUBS 0.007869f
C424 B.n384 VSUBS 0.007869f
C425 B.n385 VSUBS 0.007869f
C426 B.n386 VSUBS 0.007869f
C427 B.n387 VSUBS 0.007869f
C428 B.n388 VSUBS 0.007869f
C429 B.n389 VSUBS 0.007869f
C430 B.n390 VSUBS 0.007869f
C431 B.n391 VSUBS 0.007869f
C432 B.n392 VSUBS 0.007869f
C433 B.n393 VSUBS 0.007869f
C434 B.n394 VSUBS 0.007869f
C435 B.n395 VSUBS 0.007869f
C436 B.n396 VSUBS 0.007869f
C437 B.n397 VSUBS 0.007869f
C438 B.n398 VSUBS 0.007869f
C439 B.n399 VSUBS 0.007869f
C440 B.n400 VSUBS 0.007869f
C441 B.n401 VSUBS 0.007869f
C442 B.n402 VSUBS 0.007869f
C443 B.n403 VSUBS 0.007869f
C444 B.n404 VSUBS 0.007869f
C445 B.n405 VSUBS 0.007869f
C446 B.n406 VSUBS 0.007869f
C447 B.n407 VSUBS 0.007869f
C448 B.n408 VSUBS 0.007869f
C449 B.n409 VSUBS 0.007869f
C450 B.n410 VSUBS 0.007869f
C451 B.n411 VSUBS 0.007869f
C452 B.n412 VSUBS 0.007869f
C453 B.n413 VSUBS 0.007869f
C454 B.n414 VSUBS 0.007869f
C455 B.n415 VSUBS 0.007869f
C456 B.n416 VSUBS 0.007869f
C457 B.n417 VSUBS 0.007869f
C458 B.n418 VSUBS 0.007869f
C459 B.n419 VSUBS 0.007869f
C460 B.n420 VSUBS 0.007869f
C461 B.n421 VSUBS 0.007869f
C462 B.n422 VSUBS 0.007869f
C463 B.n423 VSUBS 0.018383f
C464 B.n424 VSUBS 0.018383f
C465 B.n425 VSUBS 0.019575f
C466 B.n426 VSUBS 0.007869f
C467 B.n427 VSUBS 0.007869f
C468 B.n428 VSUBS 0.007869f
C469 B.n429 VSUBS 0.007869f
C470 B.n430 VSUBS 0.007869f
C471 B.n431 VSUBS 0.007869f
C472 B.n432 VSUBS 0.007869f
C473 B.n433 VSUBS 0.007869f
C474 B.n434 VSUBS 0.007869f
C475 B.n435 VSUBS 0.007869f
C476 B.n436 VSUBS 0.007869f
C477 B.n437 VSUBS 0.007869f
C478 B.n438 VSUBS 0.007869f
C479 B.n439 VSUBS 0.007869f
C480 B.n440 VSUBS 0.007869f
C481 B.n441 VSUBS 0.007869f
C482 B.n442 VSUBS 0.007869f
C483 B.n443 VSUBS 0.007869f
C484 B.n444 VSUBS 0.007869f
C485 B.n445 VSUBS 0.007869f
C486 B.n446 VSUBS 0.007869f
C487 B.n447 VSUBS 0.007869f
C488 B.n448 VSUBS 0.007869f
C489 B.n449 VSUBS 0.007869f
C490 B.n450 VSUBS 0.007869f
C491 B.n451 VSUBS 0.007869f
C492 B.n452 VSUBS 0.007869f
C493 B.n453 VSUBS 0.007869f
C494 B.n454 VSUBS 0.007869f
C495 B.n455 VSUBS 0.007869f
C496 B.n456 VSUBS 0.007869f
C497 B.n457 VSUBS 0.007869f
C498 B.n458 VSUBS 0.007869f
C499 B.n459 VSUBS 0.007869f
C500 B.n460 VSUBS 0.007869f
C501 B.n461 VSUBS 0.007869f
C502 B.n462 VSUBS 0.007869f
C503 B.n463 VSUBS 0.007869f
C504 B.n464 VSUBS 0.007869f
C505 B.n465 VSUBS 0.007869f
C506 B.n466 VSUBS 0.007869f
C507 B.n467 VSUBS 0.007869f
C508 B.n468 VSUBS 0.007869f
C509 B.n469 VSUBS 0.007869f
C510 B.n470 VSUBS 0.007869f
C511 B.n471 VSUBS 0.007869f
C512 B.n472 VSUBS 0.007869f
C513 B.n473 VSUBS 0.007869f
C514 B.n474 VSUBS 0.007406f
C515 B.n475 VSUBS 0.007869f
C516 B.n476 VSUBS 0.007869f
C517 B.n477 VSUBS 0.007869f
C518 B.n478 VSUBS 0.007869f
C519 B.n479 VSUBS 0.007869f
C520 B.n480 VSUBS 0.007869f
C521 B.n481 VSUBS 0.007869f
C522 B.n482 VSUBS 0.007869f
C523 B.n483 VSUBS 0.007869f
C524 B.n484 VSUBS 0.007869f
C525 B.n485 VSUBS 0.007869f
C526 B.n486 VSUBS 0.007869f
C527 B.n487 VSUBS 0.007869f
C528 B.n488 VSUBS 0.007869f
C529 B.n489 VSUBS 0.007869f
C530 B.n490 VSUBS 0.004398f
C531 B.n491 VSUBS 0.018232f
C532 B.n492 VSUBS 0.007406f
C533 B.n493 VSUBS 0.007869f
C534 B.n494 VSUBS 0.007869f
C535 B.n495 VSUBS 0.007869f
C536 B.n496 VSUBS 0.007869f
C537 B.n497 VSUBS 0.007869f
C538 B.n498 VSUBS 0.007869f
C539 B.n499 VSUBS 0.007869f
C540 B.n500 VSUBS 0.007869f
C541 B.n501 VSUBS 0.007869f
C542 B.n502 VSUBS 0.007869f
C543 B.n503 VSUBS 0.007869f
C544 B.n504 VSUBS 0.007869f
C545 B.n505 VSUBS 0.007869f
C546 B.n506 VSUBS 0.007869f
C547 B.n507 VSUBS 0.007869f
C548 B.n508 VSUBS 0.007869f
C549 B.n509 VSUBS 0.007869f
C550 B.n510 VSUBS 0.007869f
C551 B.n511 VSUBS 0.007869f
C552 B.n512 VSUBS 0.007869f
C553 B.n513 VSUBS 0.007869f
C554 B.n514 VSUBS 0.007869f
C555 B.n515 VSUBS 0.007869f
C556 B.n516 VSUBS 0.007869f
C557 B.n517 VSUBS 0.007869f
C558 B.n518 VSUBS 0.007869f
C559 B.n519 VSUBS 0.007869f
C560 B.n520 VSUBS 0.007869f
C561 B.n521 VSUBS 0.007869f
C562 B.n522 VSUBS 0.007869f
C563 B.n523 VSUBS 0.007869f
C564 B.n524 VSUBS 0.007869f
C565 B.n525 VSUBS 0.007869f
C566 B.n526 VSUBS 0.007869f
C567 B.n527 VSUBS 0.007869f
C568 B.n528 VSUBS 0.007869f
C569 B.n529 VSUBS 0.007869f
C570 B.n530 VSUBS 0.007869f
C571 B.n531 VSUBS 0.007869f
C572 B.n532 VSUBS 0.007869f
C573 B.n533 VSUBS 0.007869f
C574 B.n534 VSUBS 0.007869f
C575 B.n535 VSUBS 0.007869f
C576 B.n536 VSUBS 0.007869f
C577 B.n537 VSUBS 0.007869f
C578 B.n538 VSUBS 0.007869f
C579 B.n539 VSUBS 0.007869f
C580 B.n540 VSUBS 0.007869f
C581 B.n541 VSUBS 0.019575f
C582 B.n542 VSUBS 0.019575f
C583 B.n543 VSUBS 0.018383f
C584 B.n544 VSUBS 0.007869f
C585 B.n545 VSUBS 0.007869f
C586 B.n546 VSUBS 0.007869f
C587 B.n547 VSUBS 0.007869f
C588 B.n548 VSUBS 0.007869f
C589 B.n549 VSUBS 0.007869f
C590 B.n550 VSUBS 0.007869f
C591 B.n551 VSUBS 0.007869f
C592 B.n552 VSUBS 0.007869f
C593 B.n553 VSUBS 0.007869f
C594 B.n554 VSUBS 0.007869f
C595 B.n555 VSUBS 0.007869f
C596 B.n556 VSUBS 0.007869f
C597 B.n557 VSUBS 0.007869f
C598 B.n558 VSUBS 0.007869f
C599 B.n559 VSUBS 0.007869f
C600 B.n560 VSUBS 0.007869f
C601 B.n561 VSUBS 0.007869f
C602 B.n562 VSUBS 0.007869f
C603 B.n563 VSUBS 0.007869f
C604 B.n564 VSUBS 0.007869f
C605 B.n565 VSUBS 0.007869f
C606 B.n566 VSUBS 0.007869f
C607 B.n567 VSUBS 0.007869f
C608 B.n568 VSUBS 0.007869f
C609 B.n569 VSUBS 0.007869f
C610 B.n570 VSUBS 0.007869f
C611 B.n571 VSUBS 0.007869f
C612 B.n572 VSUBS 0.007869f
C613 B.n573 VSUBS 0.007869f
C614 B.n574 VSUBS 0.007869f
C615 B.n575 VSUBS 0.007869f
C616 B.n576 VSUBS 0.007869f
C617 B.n577 VSUBS 0.007869f
C618 B.n578 VSUBS 0.007869f
C619 B.n579 VSUBS 0.007869f
C620 B.n580 VSUBS 0.007869f
C621 B.n581 VSUBS 0.007869f
C622 B.n582 VSUBS 0.007869f
C623 B.n583 VSUBS 0.007869f
C624 B.n584 VSUBS 0.007869f
C625 B.n585 VSUBS 0.007869f
C626 B.n586 VSUBS 0.007869f
C627 B.n587 VSUBS 0.007869f
C628 B.n588 VSUBS 0.007869f
C629 B.n589 VSUBS 0.007869f
C630 B.n590 VSUBS 0.007869f
C631 B.n591 VSUBS 0.010269f
C632 B.n592 VSUBS 0.010939f
C633 B.n593 VSUBS 0.021753f
C634 VDD1.t6 VSUBS 0.189389f
C635 VDD1.t3 VSUBS 0.189389f
C636 VDD1.n0 VSUBS 1.43253f
C637 VDD1.t1 VSUBS 0.189389f
C638 VDD1.t0 VSUBS 0.189389f
C639 VDD1.n1 VSUBS 1.4316f
C640 VDD1.t5 VSUBS 0.189389f
C641 VDD1.t7 VSUBS 0.189389f
C642 VDD1.n2 VSUBS 1.4316f
C643 VDD1.n3 VSUBS 2.97664f
C644 VDD1.t4 VSUBS 0.189389f
C645 VDD1.t2 VSUBS 0.189389f
C646 VDD1.n4 VSUBS 1.42637f
C647 VDD1.n5 VSUBS 2.63149f
C648 VP.n0 VSUBS 0.043135f
C649 VP.t0 VSUBS 1.55733f
C650 VP.n1 VSUBS 0.061768f
C651 VP.n2 VSUBS 0.043135f
C652 VP.t2 VSUBS 1.55733f
C653 VP.n3 VSUBS 0.075411f
C654 VP.n4 VSUBS 0.043135f
C655 VP.n5 VSUBS 0.049435f
C656 VP.n6 VSUBS 0.043135f
C657 VP.t5 VSUBS 1.55733f
C658 VP.n7 VSUBS 0.061768f
C659 VP.n8 VSUBS 0.043135f
C660 VP.t3 VSUBS 1.55733f
C661 VP.n9 VSUBS 0.075411f
C662 VP.t1 VSUBS 1.67609f
C663 VP.t4 VSUBS 1.55733f
C664 VP.n10 VSUBS 0.663811f
C665 VP.n11 VSUBS 0.676986f
C666 VP.n12 VSUBS 0.266565f
C667 VP.n13 VSUBS 0.043135f
C668 VP.n14 VSUBS 0.034871f
C669 VP.n15 VSUBS 0.075411f
C670 VP.n16 VSUBS 0.577738f
C671 VP.n17 VSUBS 0.051022f
C672 VP.n18 VSUBS 0.043135f
C673 VP.n19 VSUBS 0.043135f
C674 VP.n20 VSUBS 0.043135f
C675 VP.n21 VSUBS 0.064172f
C676 VP.n22 VSUBS 0.049435f
C677 VP.n23 VSUBS 0.651046f
C678 VP.n24 VSUBS 1.87696f
C679 VP.t6 VSUBS 1.55733f
C680 VP.n25 VSUBS 0.651046f
C681 VP.n26 VSUBS 1.91282f
C682 VP.n27 VSUBS 0.043135f
C683 VP.n28 VSUBS 0.043135f
C684 VP.n29 VSUBS 0.064172f
C685 VP.n30 VSUBS 0.061768f
C686 VP.t7 VSUBS 1.55733f
C687 VP.n31 VSUBS 0.577738f
C688 VP.n32 VSUBS 0.051022f
C689 VP.n33 VSUBS 0.043135f
C690 VP.n34 VSUBS 0.043135f
C691 VP.n35 VSUBS 0.043135f
C692 VP.n36 VSUBS 0.034871f
C693 VP.n37 VSUBS 0.075411f
C694 VP.n38 VSUBS 0.577738f
C695 VP.n39 VSUBS 0.051022f
C696 VP.n40 VSUBS 0.043135f
C697 VP.n41 VSUBS 0.043135f
C698 VP.n42 VSUBS 0.043135f
C699 VP.n43 VSUBS 0.064172f
C700 VP.n44 VSUBS 0.049435f
C701 VP.n45 VSUBS 0.651046f
C702 VP.n46 VSUBS 0.042102f
C703 VTAIL.t14 VSUBS 0.189004f
C704 VTAIL.t10 VSUBS 0.189004f
C705 VTAIL.n0 VSUBS 1.3143f
C706 VTAIL.n1 VSUBS 0.640846f
C707 VTAIL.n2 VSUBS 0.028395f
C708 VTAIL.n3 VSUBS 0.025256f
C709 VTAIL.n4 VSUBS 0.013572f
C710 VTAIL.n5 VSUBS 0.032078f
C711 VTAIL.n6 VSUBS 0.013971f
C712 VTAIL.n7 VSUBS 0.025256f
C713 VTAIL.n8 VSUBS 0.01437f
C714 VTAIL.n9 VSUBS 0.032078f
C715 VTAIL.n10 VSUBS 0.01437f
C716 VTAIL.n11 VSUBS 0.025256f
C717 VTAIL.n12 VSUBS 0.013572f
C718 VTAIL.n13 VSUBS 0.032078f
C719 VTAIL.n14 VSUBS 0.01437f
C720 VTAIL.n15 VSUBS 0.960842f
C721 VTAIL.n16 VSUBS 0.013572f
C722 VTAIL.t15 VSUBS 0.068961f
C723 VTAIL.n17 VSUBS 0.170059f
C724 VTAIL.n18 VSUBS 0.024131f
C725 VTAIL.n19 VSUBS 0.024059f
C726 VTAIL.n20 VSUBS 0.032078f
C727 VTAIL.n21 VSUBS 0.01437f
C728 VTAIL.n22 VSUBS 0.013572f
C729 VTAIL.n23 VSUBS 0.025256f
C730 VTAIL.n24 VSUBS 0.025256f
C731 VTAIL.n25 VSUBS 0.013572f
C732 VTAIL.n26 VSUBS 0.01437f
C733 VTAIL.n27 VSUBS 0.032078f
C734 VTAIL.n28 VSUBS 0.032078f
C735 VTAIL.n29 VSUBS 0.01437f
C736 VTAIL.n30 VSUBS 0.013572f
C737 VTAIL.n31 VSUBS 0.025256f
C738 VTAIL.n32 VSUBS 0.025256f
C739 VTAIL.n33 VSUBS 0.013572f
C740 VTAIL.n34 VSUBS 0.013572f
C741 VTAIL.n35 VSUBS 0.01437f
C742 VTAIL.n36 VSUBS 0.032078f
C743 VTAIL.n37 VSUBS 0.032078f
C744 VTAIL.n38 VSUBS 0.032078f
C745 VTAIL.n39 VSUBS 0.013971f
C746 VTAIL.n40 VSUBS 0.013572f
C747 VTAIL.n41 VSUBS 0.025256f
C748 VTAIL.n42 VSUBS 0.025256f
C749 VTAIL.n43 VSUBS 0.013572f
C750 VTAIL.n44 VSUBS 0.01437f
C751 VTAIL.n45 VSUBS 0.032078f
C752 VTAIL.n46 VSUBS 0.079851f
C753 VTAIL.n47 VSUBS 0.01437f
C754 VTAIL.n48 VSUBS 0.013572f
C755 VTAIL.n49 VSUBS 0.066314f
C756 VTAIL.n50 VSUBS 0.040484f
C757 VTAIL.n51 VSUBS 0.18637f
C758 VTAIL.n52 VSUBS 0.028395f
C759 VTAIL.n53 VSUBS 0.025256f
C760 VTAIL.n54 VSUBS 0.013572f
C761 VTAIL.n55 VSUBS 0.032078f
C762 VTAIL.n56 VSUBS 0.013971f
C763 VTAIL.n57 VSUBS 0.025256f
C764 VTAIL.n58 VSUBS 0.01437f
C765 VTAIL.n59 VSUBS 0.032078f
C766 VTAIL.n60 VSUBS 0.01437f
C767 VTAIL.n61 VSUBS 0.025256f
C768 VTAIL.n62 VSUBS 0.013572f
C769 VTAIL.n63 VSUBS 0.032078f
C770 VTAIL.n64 VSUBS 0.01437f
C771 VTAIL.n65 VSUBS 0.960842f
C772 VTAIL.n66 VSUBS 0.013572f
C773 VTAIL.t2 VSUBS 0.068961f
C774 VTAIL.n67 VSUBS 0.170059f
C775 VTAIL.n68 VSUBS 0.024131f
C776 VTAIL.n69 VSUBS 0.024059f
C777 VTAIL.n70 VSUBS 0.032078f
C778 VTAIL.n71 VSUBS 0.01437f
C779 VTAIL.n72 VSUBS 0.013572f
C780 VTAIL.n73 VSUBS 0.025256f
C781 VTAIL.n74 VSUBS 0.025256f
C782 VTAIL.n75 VSUBS 0.013572f
C783 VTAIL.n76 VSUBS 0.01437f
C784 VTAIL.n77 VSUBS 0.032078f
C785 VTAIL.n78 VSUBS 0.032078f
C786 VTAIL.n79 VSUBS 0.01437f
C787 VTAIL.n80 VSUBS 0.013572f
C788 VTAIL.n81 VSUBS 0.025256f
C789 VTAIL.n82 VSUBS 0.025256f
C790 VTAIL.n83 VSUBS 0.013572f
C791 VTAIL.n84 VSUBS 0.013572f
C792 VTAIL.n85 VSUBS 0.01437f
C793 VTAIL.n86 VSUBS 0.032078f
C794 VTAIL.n87 VSUBS 0.032078f
C795 VTAIL.n88 VSUBS 0.032078f
C796 VTAIL.n89 VSUBS 0.013971f
C797 VTAIL.n90 VSUBS 0.013572f
C798 VTAIL.n91 VSUBS 0.025256f
C799 VTAIL.n92 VSUBS 0.025256f
C800 VTAIL.n93 VSUBS 0.013572f
C801 VTAIL.n94 VSUBS 0.01437f
C802 VTAIL.n95 VSUBS 0.032078f
C803 VTAIL.n96 VSUBS 0.079851f
C804 VTAIL.n97 VSUBS 0.01437f
C805 VTAIL.n98 VSUBS 0.013572f
C806 VTAIL.n99 VSUBS 0.066314f
C807 VTAIL.n100 VSUBS 0.040484f
C808 VTAIL.n101 VSUBS 0.18637f
C809 VTAIL.t0 VSUBS 0.189004f
C810 VTAIL.t4 VSUBS 0.189004f
C811 VTAIL.n102 VSUBS 1.3143f
C812 VTAIL.n103 VSUBS 0.758182f
C813 VTAIL.n104 VSUBS 0.028395f
C814 VTAIL.n105 VSUBS 0.025256f
C815 VTAIL.n106 VSUBS 0.013572f
C816 VTAIL.n107 VSUBS 0.032078f
C817 VTAIL.n108 VSUBS 0.013971f
C818 VTAIL.n109 VSUBS 0.025256f
C819 VTAIL.n110 VSUBS 0.01437f
C820 VTAIL.n111 VSUBS 0.032078f
C821 VTAIL.n112 VSUBS 0.01437f
C822 VTAIL.n113 VSUBS 0.025256f
C823 VTAIL.n114 VSUBS 0.013572f
C824 VTAIL.n115 VSUBS 0.032078f
C825 VTAIL.n116 VSUBS 0.01437f
C826 VTAIL.n117 VSUBS 0.960842f
C827 VTAIL.n118 VSUBS 0.013572f
C828 VTAIL.t7 VSUBS 0.068961f
C829 VTAIL.n119 VSUBS 0.170059f
C830 VTAIL.n120 VSUBS 0.024131f
C831 VTAIL.n121 VSUBS 0.024059f
C832 VTAIL.n122 VSUBS 0.032078f
C833 VTAIL.n123 VSUBS 0.01437f
C834 VTAIL.n124 VSUBS 0.013572f
C835 VTAIL.n125 VSUBS 0.025256f
C836 VTAIL.n126 VSUBS 0.025256f
C837 VTAIL.n127 VSUBS 0.013572f
C838 VTAIL.n128 VSUBS 0.01437f
C839 VTAIL.n129 VSUBS 0.032078f
C840 VTAIL.n130 VSUBS 0.032078f
C841 VTAIL.n131 VSUBS 0.01437f
C842 VTAIL.n132 VSUBS 0.013572f
C843 VTAIL.n133 VSUBS 0.025256f
C844 VTAIL.n134 VSUBS 0.025256f
C845 VTAIL.n135 VSUBS 0.013572f
C846 VTAIL.n136 VSUBS 0.013572f
C847 VTAIL.n137 VSUBS 0.01437f
C848 VTAIL.n138 VSUBS 0.032078f
C849 VTAIL.n139 VSUBS 0.032078f
C850 VTAIL.n140 VSUBS 0.032078f
C851 VTAIL.n141 VSUBS 0.013971f
C852 VTAIL.n142 VSUBS 0.013572f
C853 VTAIL.n143 VSUBS 0.025256f
C854 VTAIL.n144 VSUBS 0.025256f
C855 VTAIL.n145 VSUBS 0.013572f
C856 VTAIL.n146 VSUBS 0.01437f
C857 VTAIL.n147 VSUBS 0.032078f
C858 VTAIL.n148 VSUBS 0.079851f
C859 VTAIL.n149 VSUBS 0.01437f
C860 VTAIL.n150 VSUBS 0.013572f
C861 VTAIL.n151 VSUBS 0.066314f
C862 VTAIL.n152 VSUBS 0.040484f
C863 VTAIL.n153 VSUBS 1.27766f
C864 VTAIL.n154 VSUBS 0.028395f
C865 VTAIL.n155 VSUBS 0.025256f
C866 VTAIL.n156 VSUBS 0.013572f
C867 VTAIL.n157 VSUBS 0.032078f
C868 VTAIL.n158 VSUBS 0.013971f
C869 VTAIL.n159 VSUBS 0.025256f
C870 VTAIL.n160 VSUBS 0.013971f
C871 VTAIL.n161 VSUBS 0.013572f
C872 VTAIL.n162 VSUBS 0.032078f
C873 VTAIL.n163 VSUBS 0.032078f
C874 VTAIL.n164 VSUBS 0.01437f
C875 VTAIL.n165 VSUBS 0.025256f
C876 VTAIL.n166 VSUBS 0.013572f
C877 VTAIL.n167 VSUBS 0.032078f
C878 VTAIL.n168 VSUBS 0.01437f
C879 VTAIL.n169 VSUBS 0.960842f
C880 VTAIL.n170 VSUBS 0.013572f
C881 VTAIL.t13 VSUBS 0.068961f
C882 VTAIL.n171 VSUBS 0.170059f
C883 VTAIL.n172 VSUBS 0.024131f
C884 VTAIL.n173 VSUBS 0.024059f
C885 VTAIL.n174 VSUBS 0.032078f
C886 VTAIL.n175 VSUBS 0.01437f
C887 VTAIL.n176 VSUBS 0.013572f
C888 VTAIL.n177 VSUBS 0.025256f
C889 VTAIL.n178 VSUBS 0.025256f
C890 VTAIL.n179 VSUBS 0.013572f
C891 VTAIL.n180 VSUBS 0.01437f
C892 VTAIL.n181 VSUBS 0.032078f
C893 VTAIL.n182 VSUBS 0.032078f
C894 VTAIL.n183 VSUBS 0.01437f
C895 VTAIL.n184 VSUBS 0.013572f
C896 VTAIL.n185 VSUBS 0.025256f
C897 VTAIL.n186 VSUBS 0.025256f
C898 VTAIL.n187 VSUBS 0.013572f
C899 VTAIL.n188 VSUBS 0.01437f
C900 VTAIL.n189 VSUBS 0.032078f
C901 VTAIL.n190 VSUBS 0.032078f
C902 VTAIL.n191 VSUBS 0.01437f
C903 VTAIL.n192 VSUBS 0.013572f
C904 VTAIL.n193 VSUBS 0.025256f
C905 VTAIL.n194 VSUBS 0.025256f
C906 VTAIL.n195 VSUBS 0.013572f
C907 VTAIL.n196 VSUBS 0.01437f
C908 VTAIL.n197 VSUBS 0.032078f
C909 VTAIL.n198 VSUBS 0.079851f
C910 VTAIL.n199 VSUBS 0.01437f
C911 VTAIL.n200 VSUBS 0.013572f
C912 VTAIL.n201 VSUBS 0.066314f
C913 VTAIL.n202 VSUBS 0.040484f
C914 VTAIL.n203 VSUBS 1.27766f
C915 VTAIL.t11 VSUBS 0.189004f
C916 VTAIL.t9 VSUBS 0.189004f
C917 VTAIL.n204 VSUBS 1.31431f
C918 VTAIL.n205 VSUBS 0.758173f
C919 VTAIL.n206 VSUBS 0.028395f
C920 VTAIL.n207 VSUBS 0.025256f
C921 VTAIL.n208 VSUBS 0.013572f
C922 VTAIL.n209 VSUBS 0.032078f
C923 VTAIL.n210 VSUBS 0.013971f
C924 VTAIL.n211 VSUBS 0.025256f
C925 VTAIL.n212 VSUBS 0.013971f
C926 VTAIL.n213 VSUBS 0.013572f
C927 VTAIL.n214 VSUBS 0.032078f
C928 VTAIL.n215 VSUBS 0.032078f
C929 VTAIL.n216 VSUBS 0.01437f
C930 VTAIL.n217 VSUBS 0.025256f
C931 VTAIL.n218 VSUBS 0.013572f
C932 VTAIL.n219 VSUBS 0.032078f
C933 VTAIL.n220 VSUBS 0.01437f
C934 VTAIL.n221 VSUBS 0.960842f
C935 VTAIL.n222 VSUBS 0.013572f
C936 VTAIL.t12 VSUBS 0.068961f
C937 VTAIL.n223 VSUBS 0.170059f
C938 VTAIL.n224 VSUBS 0.024131f
C939 VTAIL.n225 VSUBS 0.024059f
C940 VTAIL.n226 VSUBS 0.032078f
C941 VTAIL.n227 VSUBS 0.01437f
C942 VTAIL.n228 VSUBS 0.013572f
C943 VTAIL.n229 VSUBS 0.025256f
C944 VTAIL.n230 VSUBS 0.025256f
C945 VTAIL.n231 VSUBS 0.013572f
C946 VTAIL.n232 VSUBS 0.01437f
C947 VTAIL.n233 VSUBS 0.032078f
C948 VTAIL.n234 VSUBS 0.032078f
C949 VTAIL.n235 VSUBS 0.01437f
C950 VTAIL.n236 VSUBS 0.013572f
C951 VTAIL.n237 VSUBS 0.025256f
C952 VTAIL.n238 VSUBS 0.025256f
C953 VTAIL.n239 VSUBS 0.013572f
C954 VTAIL.n240 VSUBS 0.01437f
C955 VTAIL.n241 VSUBS 0.032078f
C956 VTAIL.n242 VSUBS 0.032078f
C957 VTAIL.n243 VSUBS 0.01437f
C958 VTAIL.n244 VSUBS 0.013572f
C959 VTAIL.n245 VSUBS 0.025256f
C960 VTAIL.n246 VSUBS 0.025256f
C961 VTAIL.n247 VSUBS 0.013572f
C962 VTAIL.n248 VSUBS 0.01437f
C963 VTAIL.n249 VSUBS 0.032078f
C964 VTAIL.n250 VSUBS 0.079851f
C965 VTAIL.n251 VSUBS 0.01437f
C966 VTAIL.n252 VSUBS 0.013572f
C967 VTAIL.n253 VSUBS 0.066314f
C968 VTAIL.n254 VSUBS 0.040484f
C969 VTAIL.n255 VSUBS 0.18637f
C970 VTAIL.n256 VSUBS 0.028395f
C971 VTAIL.n257 VSUBS 0.025256f
C972 VTAIL.n258 VSUBS 0.013572f
C973 VTAIL.n259 VSUBS 0.032078f
C974 VTAIL.n260 VSUBS 0.013971f
C975 VTAIL.n261 VSUBS 0.025256f
C976 VTAIL.n262 VSUBS 0.013971f
C977 VTAIL.n263 VSUBS 0.013572f
C978 VTAIL.n264 VSUBS 0.032078f
C979 VTAIL.n265 VSUBS 0.032078f
C980 VTAIL.n266 VSUBS 0.01437f
C981 VTAIL.n267 VSUBS 0.025256f
C982 VTAIL.n268 VSUBS 0.013572f
C983 VTAIL.n269 VSUBS 0.032078f
C984 VTAIL.n270 VSUBS 0.01437f
C985 VTAIL.n271 VSUBS 0.960842f
C986 VTAIL.n272 VSUBS 0.013572f
C987 VTAIL.t1 VSUBS 0.068961f
C988 VTAIL.n273 VSUBS 0.170059f
C989 VTAIL.n274 VSUBS 0.024131f
C990 VTAIL.n275 VSUBS 0.024059f
C991 VTAIL.n276 VSUBS 0.032078f
C992 VTAIL.n277 VSUBS 0.01437f
C993 VTAIL.n278 VSUBS 0.013572f
C994 VTAIL.n279 VSUBS 0.025256f
C995 VTAIL.n280 VSUBS 0.025256f
C996 VTAIL.n281 VSUBS 0.013572f
C997 VTAIL.n282 VSUBS 0.01437f
C998 VTAIL.n283 VSUBS 0.032078f
C999 VTAIL.n284 VSUBS 0.032078f
C1000 VTAIL.n285 VSUBS 0.01437f
C1001 VTAIL.n286 VSUBS 0.013572f
C1002 VTAIL.n287 VSUBS 0.025256f
C1003 VTAIL.n288 VSUBS 0.025256f
C1004 VTAIL.n289 VSUBS 0.013572f
C1005 VTAIL.n290 VSUBS 0.01437f
C1006 VTAIL.n291 VSUBS 0.032078f
C1007 VTAIL.n292 VSUBS 0.032078f
C1008 VTAIL.n293 VSUBS 0.01437f
C1009 VTAIL.n294 VSUBS 0.013572f
C1010 VTAIL.n295 VSUBS 0.025256f
C1011 VTAIL.n296 VSUBS 0.025256f
C1012 VTAIL.n297 VSUBS 0.013572f
C1013 VTAIL.n298 VSUBS 0.01437f
C1014 VTAIL.n299 VSUBS 0.032078f
C1015 VTAIL.n300 VSUBS 0.079851f
C1016 VTAIL.n301 VSUBS 0.01437f
C1017 VTAIL.n302 VSUBS 0.013572f
C1018 VTAIL.n303 VSUBS 0.066314f
C1019 VTAIL.n304 VSUBS 0.040484f
C1020 VTAIL.n305 VSUBS 0.18637f
C1021 VTAIL.t3 VSUBS 0.189004f
C1022 VTAIL.t6 VSUBS 0.189004f
C1023 VTAIL.n306 VSUBS 1.31431f
C1024 VTAIL.n307 VSUBS 0.758173f
C1025 VTAIL.n308 VSUBS 0.028395f
C1026 VTAIL.n309 VSUBS 0.025256f
C1027 VTAIL.n310 VSUBS 0.013572f
C1028 VTAIL.n311 VSUBS 0.032078f
C1029 VTAIL.n312 VSUBS 0.013971f
C1030 VTAIL.n313 VSUBS 0.025256f
C1031 VTAIL.n314 VSUBS 0.013971f
C1032 VTAIL.n315 VSUBS 0.013572f
C1033 VTAIL.n316 VSUBS 0.032078f
C1034 VTAIL.n317 VSUBS 0.032078f
C1035 VTAIL.n318 VSUBS 0.01437f
C1036 VTAIL.n319 VSUBS 0.025256f
C1037 VTAIL.n320 VSUBS 0.013572f
C1038 VTAIL.n321 VSUBS 0.032078f
C1039 VTAIL.n322 VSUBS 0.01437f
C1040 VTAIL.n323 VSUBS 0.960842f
C1041 VTAIL.n324 VSUBS 0.013572f
C1042 VTAIL.t5 VSUBS 0.068961f
C1043 VTAIL.n325 VSUBS 0.170059f
C1044 VTAIL.n326 VSUBS 0.024131f
C1045 VTAIL.n327 VSUBS 0.024059f
C1046 VTAIL.n328 VSUBS 0.032078f
C1047 VTAIL.n329 VSUBS 0.01437f
C1048 VTAIL.n330 VSUBS 0.013572f
C1049 VTAIL.n331 VSUBS 0.025256f
C1050 VTAIL.n332 VSUBS 0.025256f
C1051 VTAIL.n333 VSUBS 0.013572f
C1052 VTAIL.n334 VSUBS 0.01437f
C1053 VTAIL.n335 VSUBS 0.032078f
C1054 VTAIL.n336 VSUBS 0.032078f
C1055 VTAIL.n337 VSUBS 0.01437f
C1056 VTAIL.n338 VSUBS 0.013572f
C1057 VTAIL.n339 VSUBS 0.025256f
C1058 VTAIL.n340 VSUBS 0.025256f
C1059 VTAIL.n341 VSUBS 0.013572f
C1060 VTAIL.n342 VSUBS 0.01437f
C1061 VTAIL.n343 VSUBS 0.032078f
C1062 VTAIL.n344 VSUBS 0.032078f
C1063 VTAIL.n345 VSUBS 0.01437f
C1064 VTAIL.n346 VSUBS 0.013572f
C1065 VTAIL.n347 VSUBS 0.025256f
C1066 VTAIL.n348 VSUBS 0.025256f
C1067 VTAIL.n349 VSUBS 0.013572f
C1068 VTAIL.n350 VSUBS 0.01437f
C1069 VTAIL.n351 VSUBS 0.032078f
C1070 VTAIL.n352 VSUBS 0.079851f
C1071 VTAIL.n353 VSUBS 0.01437f
C1072 VTAIL.n354 VSUBS 0.013572f
C1073 VTAIL.n355 VSUBS 0.066314f
C1074 VTAIL.n356 VSUBS 0.040484f
C1075 VTAIL.n357 VSUBS 1.27766f
C1076 VTAIL.n358 VSUBS 0.028395f
C1077 VTAIL.n359 VSUBS 0.025256f
C1078 VTAIL.n360 VSUBS 0.013572f
C1079 VTAIL.n361 VSUBS 0.032078f
C1080 VTAIL.n362 VSUBS 0.013971f
C1081 VTAIL.n363 VSUBS 0.025256f
C1082 VTAIL.n364 VSUBS 0.01437f
C1083 VTAIL.n365 VSUBS 0.032078f
C1084 VTAIL.n366 VSUBS 0.01437f
C1085 VTAIL.n367 VSUBS 0.025256f
C1086 VTAIL.n368 VSUBS 0.013572f
C1087 VTAIL.n369 VSUBS 0.032078f
C1088 VTAIL.n370 VSUBS 0.01437f
C1089 VTAIL.n371 VSUBS 0.960842f
C1090 VTAIL.n372 VSUBS 0.013572f
C1091 VTAIL.t8 VSUBS 0.068961f
C1092 VTAIL.n373 VSUBS 0.170059f
C1093 VTAIL.n374 VSUBS 0.024131f
C1094 VTAIL.n375 VSUBS 0.024059f
C1095 VTAIL.n376 VSUBS 0.032078f
C1096 VTAIL.n377 VSUBS 0.01437f
C1097 VTAIL.n378 VSUBS 0.013572f
C1098 VTAIL.n379 VSUBS 0.025256f
C1099 VTAIL.n380 VSUBS 0.025256f
C1100 VTAIL.n381 VSUBS 0.013572f
C1101 VTAIL.n382 VSUBS 0.01437f
C1102 VTAIL.n383 VSUBS 0.032078f
C1103 VTAIL.n384 VSUBS 0.032078f
C1104 VTAIL.n385 VSUBS 0.01437f
C1105 VTAIL.n386 VSUBS 0.013572f
C1106 VTAIL.n387 VSUBS 0.025256f
C1107 VTAIL.n388 VSUBS 0.025256f
C1108 VTAIL.n389 VSUBS 0.013572f
C1109 VTAIL.n390 VSUBS 0.013572f
C1110 VTAIL.n391 VSUBS 0.01437f
C1111 VTAIL.n392 VSUBS 0.032078f
C1112 VTAIL.n393 VSUBS 0.032078f
C1113 VTAIL.n394 VSUBS 0.032078f
C1114 VTAIL.n395 VSUBS 0.013971f
C1115 VTAIL.n396 VSUBS 0.013572f
C1116 VTAIL.n397 VSUBS 0.025256f
C1117 VTAIL.n398 VSUBS 0.025256f
C1118 VTAIL.n399 VSUBS 0.013572f
C1119 VTAIL.n400 VSUBS 0.01437f
C1120 VTAIL.n401 VSUBS 0.032078f
C1121 VTAIL.n402 VSUBS 0.079851f
C1122 VTAIL.n403 VSUBS 0.01437f
C1123 VTAIL.n404 VSUBS 0.013572f
C1124 VTAIL.n405 VSUBS 0.066314f
C1125 VTAIL.n406 VSUBS 0.040484f
C1126 VTAIL.n407 VSUBS 1.27292f
C1127 VDD2.t3 VSUBS 0.186493f
C1128 VDD2.t2 VSUBS 0.186493f
C1129 VDD2.n0 VSUBS 1.40971f
C1130 VDD2.t6 VSUBS 0.186493f
C1131 VDD2.t4 VSUBS 0.186493f
C1132 VDD2.n1 VSUBS 1.40971f
C1133 VDD2.n2 VSUBS 2.87837f
C1134 VDD2.t7 VSUBS 0.186493f
C1135 VDD2.t1 VSUBS 0.186493f
C1136 VDD2.n3 VSUBS 1.40457f
C1137 VDD2.n4 VSUBS 2.56131f
C1138 VDD2.t0 VSUBS 0.186493f
C1139 VDD2.t5 VSUBS 0.186493f
C1140 VDD2.n5 VSUBS 1.40968f
C1141 VN.n0 VSUBS 0.041743f
C1142 VN.t7 VSUBS 1.50705f
C1143 VN.n1 VSUBS 0.059774f
C1144 VN.n2 VSUBS 0.041743f
C1145 VN.t5 VSUBS 1.50705f
C1146 VN.n3 VSUBS 0.072977f
C1147 VN.t0 VSUBS 1.62197f
C1148 VN.t1 VSUBS 1.50705f
C1149 VN.n4 VSUBS 0.642381f
C1150 VN.n5 VSUBS 0.65513f
C1151 VN.n6 VSUBS 0.25796f
C1152 VN.n7 VSUBS 0.041743f
C1153 VN.n8 VSUBS 0.033745f
C1154 VN.n9 VSUBS 0.072977f
C1155 VN.n10 VSUBS 0.559086f
C1156 VN.n11 VSUBS 0.049375f
C1157 VN.n12 VSUBS 0.041743f
C1158 VN.n13 VSUBS 0.041743f
C1159 VN.n14 VSUBS 0.041743f
C1160 VN.n15 VSUBS 0.0621f
C1161 VN.n16 VSUBS 0.047839f
C1162 VN.n17 VSUBS 0.630027f
C1163 VN.n18 VSUBS 0.040742f
C1164 VN.n19 VSUBS 0.041743f
C1165 VN.t2 VSUBS 1.50705f
C1166 VN.n20 VSUBS 0.059774f
C1167 VN.n21 VSUBS 0.041743f
C1168 VN.t4 VSUBS 1.50705f
C1169 VN.n22 VSUBS 0.072977f
C1170 VN.t3 VSUBS 1.62197f
C1171 VN.t6 VSUBS 1.50705f
C1172 VN.n23 VSUBS 0.642381f
C1173 VN.n24 VSUBS 0.65513f
C1174 VN.n25 VSUBS 0.25796f
C1175 VN.n26 VSUBS 0.041743f
C1176 VN.n27 VSUBS 0.033745f
C1177 VN.n28 VSUBS 0.072977f
C1178 VN.n29 VSUBS 0.559086f
C1179 VN.n30 VSUBS 0.049375f
C1180 VN.n31 VSUBS 0.041743f
C1181 VN.n32 VSUBS 0.041743f
C1182 VN.n33 VSUBS 0.041743f
C1183 VN.n34 VSUBS 0.0621f
C1184 VN.n35 VSUBS 0.047839f
C1185 VN.n36 VSUBS 0.630027f
C1186 VN.n37 VSUBS 1.84372f
.ends

