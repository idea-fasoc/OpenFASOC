* NGSPICE file created from diff_pair_sample_0624.ext - technology: sky130A

.subckt diff_pair_sample_0624 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=0 ps=0 w=8.3 l=3.35
X1 VTAIL.t7 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=1.3695 ps=8.63 w=8.3 l=3.35
X2 VTAIL.t6 VP.t1 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=1.3695 ps=8.63 w=8.3 l=3.35
X3 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=0 ps=0 w=8.3 l=3.35
X4 VDD1.t0 VP.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3695 pd=8.63 as=3.237 ps=17.38 w=8.3 l=3.35
X5 VDD1.t1 VP.t3 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3695 pd=8.63 as=3.237 ps=17.38 w=8.3 l=3.35
X6 VDD2.t3 VN.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.3695 pd=8.63 as=3.237 ps=17.38 w=8.3 l=3.35
X7 VDD2.t2 VN.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.3695 pd=8.63 as=3.237 ps=17.38 w=8.3 l=3.35
X8 VTAIL.t1 VN.t2 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=1.3695 ps=8.63 w=8.3 l=3.35
X9 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=0 ps=0 w=8.3 l=3.35
X10 VTAIL.t0 VN.t3 VDD2.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=1.3695 ps=8.63 w=8.3 l=3.35
X11 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.237 pd=17.38 as=0 ps=0 w=8.3 l=3.35
R0 B.n691 B.n690 585
R1 B.n692 B.n691 585
R2 B.n255 B.n112 585
R3 B.n254 B.n253 585
R4 B.n252 B.n251 585
R5 B.n250 B.n249 585
R6 B.n248 B.n247 585
R7 B.n246 B.n245 585
R8 B.n244 B.n243 585
R9 B.n242 B.n241 585
R10 B.n240 B.n239 585
R11 B.n238 B.n237 585
R12 B.n236 B.n235 585
R13 B.n234 B.n233 585
R14 B.n232 B.n231 585
R15 B.n230 B.n229 585
R16 B.n228 B.n227 585
R17 B.n226 B.n225 585
R18 B.n224 B.n223 585
R19 B.n222 B.n221 585
R20 B.n220 B.n219 585
R21 B.n218 B.n217 585
R22 B.n216 B.n215 585
R23 B.n214 B.n213 585
R24 B.n212 B.n211 585
R25 B.n210 B.n209 585
R26 B.n208 B.n207 585
R27 B.n206 B.n205 585
R28 B.n204 B.n203 585
R29 B.n202 B.n201 585
R30 B.n200 B.n199 585
R31 B.n198 B.n197 585
R32 B.n196 B.n195 585
R33 B.n194 B.n193 585
R34 B.n192 B.n191 585
R35 B.n190 B.n189 585
R36 B.n188 B.n187 585
R37 B.n186 B.n185 585
R38 B.n184 B.n183 585
R39 B.n182 B.n181 585
R40 B.n180 B.n179 585
R41 B.n177 B.n176 585
R42 B.n175 B.n174 585
R43 B.n173 B.n172 585
R44 B.n171 B.n170 585
R45 B.n169 B.n168 585
R46 B.n167 B.n166 585
R47 B.n165 B.n164 585
R48 B.n163 B.n162 585
R49 B.n161 B.n160 585
R50 B.n159 B.n158 585
R51 B.n157 B.n156 585
R52 B.n155 B.n154 585
R53 B.n153 B.n152 585
R54 B.n151 B.n150 585
R55 B.n149 B.n148 585
R56 B.n147 B.n146 585
R57 B.n145 B.n144 585
R58 B.n143 B.n142 585
R59 B.n141 B.n140 585
R60 B.n139 B.n138 585
R61 B.n137 B.n136 585
R62 B.n135 B.n134 585
R63 B.n133 B.n132 585
R64 B.n131 B.n130 585
R65 B.n129 B.n128 585
R66 B.n127 B.n126 585
R67 B.n125 B.n124 585
R68 B.n123 B.n122 585
R69 B.n121 B.n120 585
R70 B.n119 B.n118 585
R71 B.n75 B.n74 585
R72 B.n689 B.n76 585
R73 B.n693 B.n76 585
R74 B.n688 B.n687 585
R75 B.n687 B.n72 585
R76 B.n686 B.n71 585
R77 B.n699 B.n71 585
R78 B.n685 B.n70 585
R79 B.n700 B.n70 585
R80 B.n684 B.n69 585
R81 B.n701 B.n69 585
R82 B.n683 B.n682 585
R83 B.n682 B.n65 585
R84 B.n681 B.n64 585
R85 B.n707 B.n64 585
R86 B.n680 B.n63 585
R87 B.n708 B.n63 585
R88 B.n679 B.n62 585
R89 B.n709 B.n62 585
R90 B.n678 B.n677 585
R91 B.n677 B.n58 585
R92 B.n676 B.n57 585
R93 B.n715 B.n57 585
R94 B.n675 B.n56 585
R95 B.n716 B.n56 585
R96 B.n674 B.n55 585
R97 B.n717 B.n55 585
R98 B.n673 B.n672 585
R99 B.n672 B.n51 585
R100 B.n671 B.n50 585
R101 B.n723 B.n50 585
R102 B.n670 B.n49 585
R103 B.n724 B.n49 585
R104 B.n669 B.n48 585
R105 B.n725 B.n48 585
R106 B.n668 B.n667 585
R107 B.n667 B.n44 585
R108 B.n666 B.n43 585
R109 B.n731 B.n43 585
R110 B.n665 B.n42 585
R111 B.n732 B.n42 585
R112 B.n664 B.n41 585
R113 B.n733 B.n41 585
R114 B.n663 B.n662 585
R115 B.n662 B.n37 585
R116 B.n661 B.n36 585
R117 B.n739 B.n36 585
R118 B.n660 B.n35 585
R119 B.n740 B.n35 585
R120 B.n659 B.n34 585
R121 B.n741 B.n34 585
R122 B.n658 B.n657 585
R123 B.n657 B.n30 585
R124 B.n656 B.n29 585
R125 B.n747 B.n29 585
R126 B.n655 B.n28 585
R127 B.n748 B.n28 585
R128 B.n654 B.n27 585
R129 B.n749 B.n27 585
R130 B.n653 B.n652 585
R131 B.n652 B.n23 585
R132 B.n651 B.n22 585
R133 B.n755 B.n22 585
R134 B.n650 B.n21 585
R135 B.n756 B.n21 585
R136 B.n649 B.n20 585
R137 B.n757 B.n20 585
R138 B.n648 B.n647 585
R139 B.n647 B.n19 585
R140 B.n646 B.n15 585
R141 B.n763 B.n15 585
R142 B.n645 B.n14 585
R143 B.n764 B.n14 585
R144 B.n644 B.n13 585
R145 B.n765 B.n13 585
R146 B.n643 B.n642 585
R147 B.n642 B.n12 585
R148 B.n641 B.n640 585
R149 B.n641 B.n8 585
R150 B.n639 B.n7 585
R151 B.n772 B.n7 585
R152 B.n638 B.n6 585
R153 B.n773 B.n6 585
R154 B.n637 B.n5 585
R155 B.n774 B.n5 585
R156 B.n636 B.n635 585
R157 B.n635 B.n4 585
R158 B.n634 B.n256 585
R159 B.n634 B.n633 585
R160 B.n624 B.n257 585
R161 B.n258 B.n257 585
R162 B.n626 B.n625 585
R163 B.n627 B.n626 585
R164 B.n623 B.n263 585
R165 B.n263 B.n262 585
R166 B.n622 B.n621 585
R167 B.n621 B.n620 585
R168 B.n265 B.n264 585
R169 B.n613 B.n265 585
R170 B.n612 B.n611 585
R171 B.n614 B.n612 585
R172 B.n610 B.n270 585
R173 B.n270 B.n269 585
R174 B.n609 B.n608 585
R175 B.n608 B.n607 585
R176 B.n272 B.n271 585
R177 B.n273 B.n272 585
R178 B.n600 B.n599 585
R179 B.n601 B.n600 585
R180 B.n598 B.n278 585
R181 B.n278 B.n277 585
R182 B.n597 B.n596 585
R183 B.n596 B.n595 585
R184 B.n280 B.n279 585
R185 B.n281 B.n280 585
R186 B.n588 B.n587 585
R187 B.n589 B.n588 585
R188 B.n586 B.n286 585
R189 B.n286 B.n285 585
R190 B.n585 B.n584 585
R191 B.n584 B.n583 585
R192 B.n288 B.n287 585
R193 B.n289 B.n288 585
R194 B.n576 B.n575 585
R195 B.n577 B.n576 585
R196 B.n574 B.n294 585
R197 B.n294 B.n293 585
R198 B.n573 B.n572 585
R199 B.n572 B.n571 585
R200 B.n296 B.n295 585
R201 B.n297 B.n296 585
R202 B.n564 B.n563 585
R203 B.n565 B.n564 585
R204 B.n562 B.n302 585
R205 B.n302 B.n301 585
R206 B.n561 B.n560 585
R207 B.n560 B.n559 585
R208 B.n304 B.n303 585
R209 B.n305 B.n304 585
R210 B.n552 B.n551 585
R211 B.n553 B.n552 585
R212 B.n550 B.n310 585
R213 B.n310 B.n309 585
R214 B.n549 B.n548 585
R215 B.n548 B.n547 585
R216 B.n312 B.n311 585
R217 B.n313 B.n312 585
R218 B.n540 B.n539 585
R219 B.n541 B.n540 585
R220 B.n538 B.n318 585
R221 B.n318 B.n317 585
R222 B.n537 B.n536 585
R223 B.n536 B.n535 585
R224 B.n320 B.n319 585
R225 B.n321 B.n320 585
R226 B.n528 B.n527 585
R227 B.n529 B.n528 585
R228 B.n526 B.n326 585
R229 B.n326 B.n325 585
R230 B.n525 B.n524 585
R231 B.n524 B.n523 585
R232 B.n328 B.n327 585
R233 B.n329 B.n328 585
R234 B.n516 B.n515 585
R235 B.n517 B.n516 585
R236 B.n332 B.n331 585
R237 B.n373 B.n372 585
R238 B.n374 B.n370 585
R239 B.n370 B.n333 585
R240 B.n376 B.n375 585
R241 B.n378 B.n369 585
R242 B.n381 B.n380 585
R243 B.n382 B.n368 585
R244 B.n384 B.n383 585
R245 B.n386 B.n367 585
R246 B.n389 B.n388 585
R247 B.n390 B.n366 585
R248 B.n392 B.n391 585
R249 B.n394 B.n365 585
R250 B.n397 B.n396 585
R251 B.n398 B.n364 585
R252 B.n400 B.n399 585
R253 B.n402 B.n363 585
R254 B.n405 B.n404 585
R255 B.n406 B.n362 585
R256 B.n408 B.n407 585
R257 B.n410 B.n361 585
R258 B.n413 B.n412 585
R259 B.n414 B.n360 585
R260 B.n416 B.n415 585
R261 B.n418 B.n359 585
R262 B.n421 B.n420 585
R263 B.n422 B.n358 585
R264 B.n424 B.n423 585
R265 B.n426 B.n357 585
R266 B.n429 B.n428 585
R267 B.n430 B.n354 585
R268 B.n433 B.n432 585
R269 B.n435 B.n353 585
R270 B.n438 B.n437 585
R271 B.n439 B.n352 585
R272 B.n441 B.n440 585
R273 B.n443 B.n351 585
R274 B.n446 B.n445 585
R275 B.n447 B.n350 585
R276 B.n452 B.n451 585
R277 B.n454 B.n349 585
R278 B.n457 B.n456 585
R279 B.n458 B.n348 585
R280 B.n460 B.n459 585
R281 B.n462 B.n347 585
R282 B.n465 B.n464 585
R283 B.n466 B.n346 585
R284 B.n468 B.n467 585
R285 B.n470 B.n345 585
R286 B.n473 B.n472 585
R287 B.n474 B.n344 585
R288 B.n476 B.n475 585
R289 B.n478 B.n343 585
R290 B.n481 B.n480 585
R291 B.n482 B.n342 585
R292 B.n484 B.n483 585
R293 B.n486 B.n341 585
R294 B.n489 B.n488 585
R295 B.n490 B.n340 585
R296 B.n492 B.n491 585
R297 B.n494 B.n339 585
R298 B.n497 B.n496 585
R299 B.n498 B.n338 585
R300 B.n500 B.n499 585
R301 B.n502 B.n337 585
R302 B.n505 B.n504 585
R303 B.n506 B.n336 585
R304 B.n508 B.n507 585
R305 B.n510 B.n335 585
R306 B.n513 B.n512 585
R307 B.n514 B.n334 585
R308 B.n519 B.n518 585
R309 B.n518 B.n517 585
R310 B.n520 B.n330 585
R311 B.n330 B.n329 585
R312 B.n522 B.n521 585
R313 B.n523 B.n522 585
R314 B.n324 B.n323 585
R315 B.n325 B.n324 585
R316 B.n531 B.n530 585
R317 B.n530 B.n529 585
R318 B.n532 B.n322 585
R319 B.n322 B.n321 585
R320 B.n534 B.n533 585
R321 B.n535 B.n534 585
R322 B.n316 B.n315 585
R323 B.n317 B.n316 585
R324 B.n543 B.n542 585
R325 B.n542 B.n541 585
R326 B.n544 B.n314 585
R327 B.n314 B.n313 585
R328 B.n546 B.n545 585
R329 B.n547 B.n546 585
R330 B.n308 B.n307 585
R331 B.n309 B.n308 585
R332 B.n555 B.n554 585
R333 B.n554 B.n553 585
R334 B.n556 B.n306 585
R335 B.n306 B.n305 585
R336 B.n558 B.n557 585
R337 B.n559 B.n558 585
R338 B.n300 B.n299 585
R339 B.n301 B.n300 585
R340 B.n567 B.n566 585
R341 B.n566 B.n565 585
R342 B.n568 B.n298 585
R343 B.n298 B.n297 585
R344 B.n570 B.n569 585
R345 B.n571 B.n570 585
R346 B.n292 B.n291 585
R347 B.n293 B.n292 585
R348 B.n579 B.n578 585
R349 B.n578 B.n577 585
R350 B.n580 B.n290 585
R351 B.n290 B.n289 585
R352 B.n582 B.n581 585
R353 B.n583 B.n582 585
R354 B.n284 B.n283 585
R355 B.n285 B.n284 585
R356 B.n591 B.n590 585
R357 B.n590 B.n589 585
R358 B.n592 B.n282 585
R359 B.n282 B.n281 585
R360 B.n594 B.n593 585
R361 B.n595 B.n594 585
R362 B.n276 B.n275 585
R363 B.n277 B.n276 585
R364 B.n603 B.n602 585
R365 B.n602 B.n601 585
R366 B.n604 B.n274 585
R367 B.n274 B.n273 585
R368 B.n606 B.n605 585
R369 B.n607 B.n606 585
R370 B.n268 B.n267 585
R371 B.n269 B.n268 585
R372 B.n616 B.n615 585
R373 B.n615 B.n614 585
R374 B.n617 B.n266 585
R375 B.n613 B.n266 585
R376 B.n619 B.n618 585
R377 B.n620 B.n619 585
R378 B.n261 B.n260 585
R379 B.n262 B.n261 585
R380 B.n629 B.n628 585
R381 B.n628 B.n627 585
R382 B.n630 B.n259 585
R383 B.n259 B.n258 585
R384 B.n632 B.n631 585
R385 B.n633 B.n632 585
R386 B.n3 B.n0 585
R387 B.n4 B.n3 585
R388 B.n771 B.n1 585
R389 B.n772 B.n771 585
R390 B.n770 B.n769 585
R391 B.n770 B.n8 585
R392 B.n768 B.n9 585
R393 B.n12 B.n9 585
R394 B.n767 B.n766 585
R395 B.n766 B.n765 585
R396 B.n11 B.n10 585
R397 B.n764 B.n11 585
R398 B.n762 B.n761 585
R399 B.n763 B.n762 585
R400 B.n760 B.n16 585
R401 B.n19 B.n16 585
R402 B.n759 B.n758 585
R403 B.n758 B.n757 585
R404 B.n18 B.n17 585
R405 B.n756 B.n18 585
R406 B.n754 B.n753 585
R407 B.n755 B.n754 585
R408 B.n752 B.n24 585
R409 B.n24 B.n23 585
R410 B.n751 B.n750 585
R411 B.n750 B.n749 585
R412 B.n26 B.n25 585
R413 B.n748 B.n26 585
R414 B.n746 B.n745 585
R415 B.n747 B.n746 585
R416 B.n744 B.n31 585
R417 B.n31 B.n30 585
R418 B.n743 B.n742 585
R419 B.n742 B.n741 585
R420 B.n33 B.n32 585
R421 B.n740 B.n33 585
R422 B.n738 B.n737 585
R423 B.n739 B.n738 585
R424 B.n736 B.n38 585
R425 B.n38 B.n37 585
R426 B.n735 B.n734 585
R427 B.n734 B.n733 585
R428 B.n40 B.n39 585
R429 B.n732 B.n40 585
R430 B.n730 B.n729 585
R431 B.n731 B.n730 585
R432 B.n728 B.n45 585
R433 B.n45 B.n44 585
R434 B.n727 B.n726 585
R435 B.n726 B.n725 585
R436 B.n47 B.n46 585
R437 B.n724 B.n47 585
R438 B.n722 B.n721 585
R439 B.n723 B.n722 585
R440 B.n720 B.n52 585
R441 B.n52 B.n51 585
R442 B.n719 B.n718 585
R443 B.n718 B.n717 585
R444 B.n54 B.n53 585
R445 B.n716 B.n54 585
R446 B.n714 B.n713 585
R447 B.n715 B.n714 585
R448 B.n712 B.n59 585
R449 B.n59 B.n58 585
R450 B.n711 B.n710 585
R451 B.n710 B.n709 585
R452 B.n61 B.n60 585
R453 B.n708 B.n61 585
R454 B.n706 B.n705 585
R455 B.n707 B.n706 585
R456 B.n704 B.n66 585
R457 B.n66 B.n65 585
R458 B.n703 B.n702 585
R459 B.n702 B.n701 585
R460 B.n68 B.n67 585
R461 B.n700 B.n68 585
R462 B.n698 B.n697 585
R463 B.n699 B.n698 585
R464 B.n696 B.n73 585
R465 B.n73 B.n72 585
R466 B.n695 B.n694 585
R467 B.n694 B.n693 585
R468 B.n775 B.n774 585
R469 B.n773 B.n2 585
R470 B.n694 B.n75 516.524
R471 B.n691 B.n76 516.524
R472 B.n516 B.n334 516.524
R473 B.n518 B.n332 516.524
R474 B.n116 B.t15 268.664
R475 B.n113 B.t11 268.664
R476 B.n448 B.t8 268.664
R477 B.n355 B.t4 268.664
R478 B.n692 B.n111 256.663
R479 B.n692 B.n110 256.663
R480 B.n692 B.n109 256.663
R481 B.n692 B.n108 256.663
R482 B.n692 B.n107 256.663
R483 B.n692 B.n106 256.663
R484 B.n692 B.n105 256.663
R485 B.n692 B.n104 256.663
R486 B.n692 B.n103 256.663
R487 B.n692 B.n102 256.663
R488 B.n692 B.n101 256.663
R489 B.n692 B.n100 256.663
R490 B.n692 B.n99 256.663
R491 B.n692 B.n98 256.663
R492 B.n692 B.n97 256.663
R493 B.n692 B.n96 256.663
R494 B.n692 B.n95 256.663
R495 B.n692 B.n94 256.663
R496 B.n692 B.n93 256.663
R497 B.n692 B.n92 256.663
R498 B.n692 B.n91 256.663
R499 B.n692 B.n90 256.663
R500 B.n692 B.n89 256.663
R501 B.n692 B.n88 256.663
R502 B.n692 B.n87 256.663
R503 B.n692 B.n86 256.663
R504 B.n692 B.n85 256.663
R505 B.n692 B.n84 256.663
R506 B.n692 B.n83 256.663
R507 B.n692 B.n82 256.663
R508 B.n692 B.n81 256.663
R509 B.n692 B.n80 256.663
R510 B.n692 B.n79 256.663
R511 B.n692 B.n78 256.663
R512 B.n692 B.n77 256.663
R513 B.n371 B.n333 256.663
R514 B.n377 B.n333 256.663
R515 B.n379 B.n333 256.663
R516 B.n385 B.n333 256.663
R517 B.n387 B.n333 256.663
R518 B.n393 B.n333 256.663
R519 B.n395 B.n333 256.663
R520 B.n401 B.n333 256.663
R521 B.n403 B.n333 256.663
R522 B.n409 B.n333 256.663
R523 B.n411 B.n333 256.663
R524 B.n417 B.n333 256.663
R525 B.n419 B.n333 256.663
R526 B.n425 B.n333 256.663
R527 B.n427 B.n333 256.663
R528 B.n434 B.n333 256.663
R529 B.n436 B.n333 256.663
R530 B.n442 B.n333 256.663
R531 B.n444 B.n333 256.663
R532 B.n453 B.n333 256.663
R533 B.n455 B.n333 256.663
R534 B.n461 B.n333 256.663
R535 B.n463 B.n333 256.663
R536 B.n469 B.n333 256.663
R537 B.n471 B.n333 256.663
R538 B.n477 B.n333 256.663
R539 B.n479 B.n333 256.663
R540 B.n485 B.n333 256.663
R541 B.n487 B.n333 256.663
R542 B.n493 B.n333 256.663
R543 B.n495 B.n333 256.663
R544 B.n501 B.n333 256.663
R545 B.n503 B.n333 256.663
R546 B.n509 B.n333 256.663
R547 B.n511 B.n333 256.663
R548 B.n777 B.n776 256.663
R549 B.n120 B.n119 163.367
R550 B.n124 B.n123 163.367
R551 B.n128 B.n127 163.367
R552 B.n132 B.n131 163.367
R553 B.n136 B.n135 163.367
R554 B.n140 B.n139 163.367
R555 B.n144 B.n143 163.367
R556 B.n148 B.n147 163.367
R557 B.n152 B.n151 163.367
R558 B.n156 B.n155 163.367
R559 B.n160 B.n159 163.367
R560 B.n164 B.n163 163.367
R561 B.n168 B.n167 163.367
R562 B.n172 B.n171 163.367
R563 B.n176 B.n175 163.367
R564 B.n181 B.n180 163.367
R565 B.n185 B.n184 163.367
R566 B.n189 B.n188 163.367
R567 B.n193 B.n192 163.367
R568 B.n197 B.n196 163.367
R569 B.n201 B.n200 163.367
R570 B.n205 B.n204 163.367
R571 B.n209 B.n208 163.367
R572 B.n213 B.n212 163.367
R573 B.n217 B.n216 163.367
R574 B.n221 B.n220 163.367
R575 B.n225 B.n224 163.367
R576 B.n229 B.n228 163.367
R577 B.n233 B.n232 163.367
R578 B.n237 B.n236 163.367
R579 B.n241 B.n240 163.367
R580 B.n245 B.n244 163.367
R581 B.n249 B.n248 163.367
R582 B.n253 B.n252 163.367
R583 B.n691 B.n112 163.367
R584 B.n516 B.n328 163.367
R585 B.n524 B.n328 163.367
R586 B.n524 B.n326 163.367
R587 B.n528 B.n326 163.367
R588 B.n528 B.n320 163.367
R589 B.n536 B.n320 163.367
R590 B.n536 B.n318 163.367
R591 B.n540 B.n318 163.367
R592 B.n540 B.n312 163.367
R593 B.n548 B.n312 163.367
R594 B.n548 B.n310 163.367
R595 B.n552 B.n310 163.367
R596 B.n552 B.n304 163.367
R597 B.n560 B.n304 163.367
R598 B.n560 B.n302 163.367
R599 B.n564 B.n302 163.367
R600 B.n564 B.n296 163.367
R601 B.n572 B.n296 163.367
R602 B.n572 B.n294 163.367
R603 B.n576 B.n294 163.367
R604 B.n576 B.n288 163.367
R605 B.n584 B.n288 163.367
R606 B.n584 B.n286 163.367
R607 B.n588 B.n286 163.367
R608 B.n588 B.n280 163.367
R609 B.n596 B.n280 163.367
R610 B.n596 B.n278 163.367
R611 B.n600 B.n278 163.367
R612 B.n600 B.n272 163.367
R613 B.n608 B.n272 163.367
R614 B.n608 B.n270 163.367
R615 B.n612 B.n270 163.367
R616 B.n612 B.n265 163.367
R617 B.n621 B.n265 163.367
R618 B.n621 B.n263 163.367
R619 B.n626 B.n263 163.367
R620 B.n626 B.n257 163.367
R621 B.n634 B.n257 163.367
R622 B.n635 B.n634 163.367
R623 B.n635 B.n5 163.367
R624 B.n6 B.n5 163.367
R625 B.n7 B.n6 163.367
R626 B.n641 B.n7 163.367
R627 B.n642 B.n641 163.367
R628 B.n642 B.n13 163.367
R629 B.n14 B.n13 163.367
R630 B.n15 B.n14 163.367
R631 B.n647 B.n15 163.367
R632 B.n647 B.n20 163.367
R633 B.n21 B.n20 163.367
R634 B.n22 B.n21 163.367
R635 B.n652 B.n22 163.367
R636 B.n652 B.n27 163.367
R637 B.n28 B.n27 163.367
R638 B.n29 B.n28 163.367
R639 B.n657 B.n29 163.367
R640 B.n657 B.n34 163.367
R641 B.n35 B.n34 163.367
R642 B.n36 B.n35 163.367
R643 B.n662 B.n36 163.367
R644 B.n662 B.n41 163.367
R645 B.n42 B.n41 163.367
R646 B.n43 B.n42 163.367
R647 B.n667 B.n43 163.367
R648 B.n667 B.n48 163.367
R649 B.n49 B.n48 163.367
R650 B.n50 B.n49 163.367
R651 B.n672 B.n50 163.367
R652 B.n672 B.n55 163.367
R653 B.n56 B.n55 163.367
R654 B.n57 B.n56 163.367
R655 B.n677 B.n57 163.367
R656 B.n677 B.n62 163.367
R657 B.n63 B.n62 163.367
R658 B.n64 B.n63 163.367
R659 B.n682 B.n64 163.367
R660 B.n682 B.n69 163.367
R661 B.n70 B.n69 163.367
R662 B.n71 B.n70 163.367
R663 B.n687 B.n71 163.367
R664 B.n687 B.n76 163.367
R665 B.n372 B.n370 163.367
R666 B.n376 B.n370 163.367
R667 B.n380 B.n378 163.367
R668 B.n384 B.n368 163.367
R669 B.n388 B.n386 163.367
R670 B.n392 B.n366 163.367
R671 B.n396 B.n394 163.367
R672 B.n400 B.n364 163.367
R673 B.n404 B.n402 163.367
R674 B.n408 B.n362 163.367
R675 B.n412 B.n410 163.367
R676 B.n416 B.n360 163.367
R677 B.n420 B.n418 163.367
R678 B.n424 B.n358 163.367
R679 B.n428 B.n426 163.367
R680 B.n433 B.n354 163.367
R681 B.n437 B.n435 163.367
R682 B.n441 B.n352 163.367
R683 B.n445 B.n443 163.367
R684 B.n452 B.n350 163.367
R685 B.n456 B.n454 163.367
R686 B.n460 B.n348 163.367
R687 B.n464 B.n462 163.367
R688 B.n468 B.n346 163.367
R689 B.n472 B.n470 163.367
R690 B.n476 B.n344 163.367
R691 B.n480 B.n478 163.367
R692 B.n484 B.n342 163.367
R693 B.n488 B.n486 163.367
R694 B.n492 B.n340 163.367
R695 B.n496 B.n494 163.367
R696 B.n500 B.n338 163.367
R697 B.n504 B.n502 163.367
R698 B.n508 B.n336 163.367
R699 B.n512 B.n510 163.367
R700 B.n518 B.n330 163.367
R701 B.n522 B.n330 163.367
R702 B.n522 B.n324 163.367
R703 B.n530 B.n324 163.367
R704 B.n530 B.n322 163.367
R705 B.n534 B.n322 163.367
R706 B.n534 B.n316 163.367
R707 B.n542 B.n316 163.367
R708 B.n542 B.n314 163.367
R709 B.n546 B.n314 163.367
R710 B.n546 B.n308 163.367
R711 B.n554 B.n308 163.367
R712 B.n554 B.n306 163.367
R713 B.n558 B.n306 163.367
R714 B.n558 B.n300 163.367
R715 B.n566 B.n300 163.367
R716 B.n566 B.n298 163.367
R717 B.n570 B.n298 163.367
R718 B.n570 B.n292 163.367
R719 B.n578 B.n292 163.367
R720 B.n578 B.n290 163.367
R721 B.n582 B.n290 163.367
R722 B.n582 B.n284 163.367
R723 B.n590 B.n284 163.367
R724 B.n590 B.n282 163.367
R725 B.n594 B.n282 163.367
R726 B.n594 B.n276 163.367
R727 B.n602 B.n276 163.367
R728 B.n602 B.n274 163.367
R729 B.n606 B.n274 163.367
R730 B.n606 B.n268 163.367
R731 B.n615 B.n268 163.367
R732 B.n615 B.n266 163.367
R733 B.n619 B.n266 163.367
R734 B.n619 B.n261 163.367
R735 B.n628 B.n261 163.367
R736 B.n628 B.n259 163.367
R737 B.n632 B.n259 163.367
R738 B.n632 B.n3 163.367
R739 B.n775 B.n3 163.367
R740 B.n771 B.n2 163.367
R741 B.n771 B.n770 163.367
R742 B.n770 B.n9 163.367
R743 B.n766 B.n9 163.367
R744 B.n766 B.n11 163.367
R745 B.n762 B.n11 163.367
R746 B.n762 B.n16 163.367
R747 B.n758 B.n16 163.367
R748 B.n758 B.n18 163.367
R749 B.n754 B.n18 163.367
R750 B.n754 B.n24 163.367
R751 B.n750 B.n24 163.367
R752 B.n750 B.n26 163.367
R753 B.n746 B.n26 163.367
R754 B.n746 B.n31 163.367
R755 B.n742 B.n31 163.367
R756 B.n742 B.n33 163.367
R757 B.n738 B.n33 163.367
R758 B.n738 B.n38 163.367
R759 B.n734 B.n38 163.367
R760 B.n734 B.n40 163.367
R761 B.n730 B.n40 163.367
R762 B.n730 B.n45 163.367
R763 B.n726 B.n45 163.367
R764 B.n726 B.n47 163.367
R765 B.n722 B.n47 163.367
R766 B.n722 B.n52 163.367
R767 B.n718 B.n52 163.367
R768 B.n718 B.n54 163.367
R769 B.n714 B.n54 163.367
R770 B.n714 B.n59 163.367
R771 B.n710 B.n59 163.367
R772 B.n710 B.n61 163.367
R773 B.n706 B.n61 163.367
R774 B.n706 B.n66 163.367
R775 B.n702 B.n66 163.367
R776 B.n702 B.n68 163.367
R777 B.n698 B.n68 163.367
R778 B.n698 B.n73 163.367
R779 B.n694 B.n73 163.367
R780 B.n113 B.t13 142.606
R781 B.n448 B.t10 142.606
R782 B.n116 B.t16 142.595
R783 B.n355 B.t7 142.595
R784 B.n517 B.n333 104.531
R785 B.n693 B.n692 104.531
R786 B.n77 B.n75 71.676
R787 B.n120 B.n78 71.676
R788 B.n124 B.n79 71.676
R789 B.n128 B.n80 71.676
R790 B.n132 B.n81 71.676
R791 B.n136 B.n82 71.676
R792 B.n140 B.n83 71.676
R793 B.n144 B.n84 71.676
R794 B.n148 B.n85 71.676
R795 B.n152 B.n86 71.676
R796 B.n156 B.n87 71.676
R797 B.n160 B.n88 71.676
R798 B.n164 B.n89 71.676
R799 B.n168 B.n90 71.676
R800 B.n172 B.n91 71.676
R801 B.n176 B.n92 71.676
R802 B.n181 B.n93 71.676
R803 B.n185 B.n94 71.676
R804 B.n189 B.n95 71.676
R805 B.n193 B.n96 71.676
R806 B.n197 B.n97 71.676
R807 B.n201 B.n98 71.676
R808 B.n205 B.n99 71.676
R809 B.n209 B.n100 71.676
R810 B.n213 B.n101 71.676
R811 B.n217 B.n102 71.676
R812 B.n221 B.n103 71.676
R813 B.n225 B.n104 71.676
R814 B.n229 B.n105 71.676
R815 B.n233 B.n106 71.676
R816 B.n237 B.n107 71.676
R817 B.n241 B.n108 71.676
R818 B.n245 B.n109 71.676
R819 B.n249 B.n110 71.676
R820 B.n253 B.n111 71.676
R821 B.n112 B.n111 71.676
R822 B.n252 B.n110 71.676
R823 B.n248 B.n109 71.676
R824 B.n244 B.n108 71.676
R825 B.n240 B.n107 71.676
R826 B.n236 B.n106 71.676
R827 B.n232 B.n105 71.676
R828 B.n228 B.n104 71.676
R829 B.n224 B.n103 71.676
R830 B.n220 B.n102 71.676
R831 B.n216 B.n101 71.676
R832 B.n212 B.n100 71.676
R833 B.n208 B.n99 71.676
R834 B.n204 B.n98 71.676
R835 B.n200 B.n97 71.676
R836 B.n196 B.n96 71.676
R837 B.n192 B.n95 71.676
R838 B.n188 B.n94 71.676
R839 B.n184 B.n93 71.676
R840 B.n180 B.n92 71.676
R841 B.n175 B.n91 71.676
R842 B.n171 B.n90 71.676
R843 B.n167 B.n89 71.676
R844 B.n163 B.n88 71.676
R845 B.n159 B.n87 71.676
R846 B.n155 B.n86 71.676
R847 B.n151 B.n85 71.676
R848 B.n147 B.n84 71.676
R849 B.n143 B.n83 71.676
R850 B.n139 B.n82 71.676
R851 B.n135 B.n81 71.676
R852 B.n131 B.n80 71.676
R853 B.n127 B.n79 71.676
R854 B.n123 B.n78 71.676
R855 B.n119 B.n77 71.676
R856 B.n371 B.n332 71.676
R857 B.n377 B.n376 71.676
R858 B.n380 B.n379 71.676
R859 B.n385 B.n384 71.676
R860 B.n388 B.n387 71.676
R861 B.n393 B.n392 71.676
R862 B.n396 B.n395 71.676
R863 B.n401 B.n400 71.676
R864 B.n404 B.n403 71.676
R865 B.n409 B.n408 71.676
R866 B.n412 B.n411 71.676
R867 B.n417 B.n416 71.676
R868 B.n420 B.n419 71.676
R869 B.n425 B.n424 71.676
R870 B.n428 B.n427 71.676
R871 B.n434 B.n433 71.676
R872 B.n437 B.n436 71.676
R873 B.n442 B.n441 71.676
R874 B.n445 B.n444 71.676
R875 B.n453 B.n452 71.676
R876 B.n456 B.n455 71.676
R877 B.n461 B.n460 71.676
R878 B.n464 B.n463 71.676
R879 B.n469 B.n468 71.676
R880 B.n472 B.n471 71.676
R881 B.n477 B.n476 71.676
R882 B.n480 B.n479 71.676
R883 B.n485 B.n484 71.676
R884 B.n488 B.n487 71.676
R885 B.n493 B.n492 71.676
R886 B.n496 B.n495 71.676
R887 B.n501 B.n500 71.676
R888 B.n504 B.n503 71.676
R889 B.n509 B.n508 71.676
R890 B.n512 B.n511 71.676
R891 B.n372 B.n371 71.676
R892 B.n378 B.n377 71.676
R893 B.n379 B.n368 71.676
R894 B.n386 B.n385 71.676
R895 B.n387 B.n366 71.676
R896 B.n394 B.n393 71.676
R897 B.n395 B.n364 71.676
R898 B.n402 B.n401 71.676
R899 B.n403 B.n362 71.676
R900 B.n410 B.n409 71.676
R901 B.n411 B.n360 71.676
R902 B.n418 B.n417 71.676
R903 B.n419 B.n358 71.676
R904 B.n426 B.n425 71.676
R905 B.n427 B.n354 71.676
R906 B.n435 B.n434 71.676
R907 B.n436 B.n352 71.676
R908 B.n443 B.n442 71.676
R909 B.n444 B.n350 71.676
R910 B.n454 B.n453 71.676
R911 B.n455 B.n348 71.676
R912 B.n462 B.n461 71.676
R913 B.n463 B.n346 71.676
R914 B.n470 B.n469 71.676
R915 B.n471 B.n344 71.676
R916 B.n478 B.n477 71.676
R917 B.n479 B.n342 71.676
R918 B.n486 B.n485 71.676
R919 B.n487 B.n340 71.676
R920 B.n494 B.n493 71.676
R921 B.n495 B.n338 71.676
R922 B.n502 B.n501 71.676
R923 B.n503 B.n336 71.676
R924 B.n510 B.n509 71.676
R925 B.n511 B.n334 71.676
R926 B.n776 B.n775 71.676
R927 B.n776 B.n2 71.676
R928 B.n117 B.n116 71.3702
R929 B.n114 B.n113 71.3702
R930 B.n449 B.n448 71.3702
R931 B.n356 B.n355 71.3702
R932 B.n114 B.t14 71.2356
R933 B.n449 B.t9 71.2356
R934 B.n117 B.t17 71.2258
R935 B.n356 B.t6 71.2258
R936 B.n178 B.n117 59.5399
R937 B.n115 B.n114 59.5399
R938 B.n450 B.n449 59.5399
R939 B.n431 B.n356 59.5399
R940 B.n517 B.n329 55.1018
R941 B.n523 B.n329 55.1018
R942 B.n523 B.n325 55.1018
R943 B.n529 B.n325 55.1018
R944 B.n529 B.n321 55.1018
R945 B.n535 B.n321 55.1018
R946 B.n535 B.n317 55.1018
R947 B.n541 B.n317 55.1018
R948 B.n547 B.n313 55.1018
R949 B.n547 B.n309 55.1018
R950 B.n553 B.n309 55.1018
R951 B.n553 B.n305 55.1018
R952 B.n559 B.n305 55.1018
R953 B.n559 B.n301 55.1018
R954 B.n565 B.n301 55.1018
R955 B.n565 B.n297 55.1018
R956 B.n571 B.n297 55.1018
R957 B.n571 B.n293 55.1018
R958 B.n577 B.n293 55.1018
R959 B.n577 B.n289 55.1018
R960 B.n583 B.n289 55.1018
R961 B.n589 B.n285 55.1018
R962 B.n589 B.n281 55.1018
R963 B.n595 B.n281 55.1018
R964 B.n595 B.n277 55.1018
R965 B.n601 B.n277 55.1018
R966 B.n601 B.n273 55.1018
R967 B.n607 B.n273 55.1018
R968 B.n607 B.n269 55.1018
R969 B.n614 B.n269 55.1018
R970 B.n614 B.n613 55.1018
R971 B.n620 B.n262 55.1018
R972 B.n627 B.n262 55.1018
R973 B.n627 B.n258 55.1018
R974 B.n633 B.n258 55.1018
R975 B.n633 B.n4 55.1018
R976 B.n774 B.n4 55.1018
R977 B.n774 B.n773 55.1018
R978 B.n773 B.n772 55.1018
R979 B.n772 B.n8 55.1018
R980 B.n12 B.n8 55.1018
R981 B.n765 B.n12 55.1018
R982 B.n765 B.n764 55.1018
R983 B.n764 B.n763 55.1018
R984 B.n757 B.n19 55.1018
R985 B.n757 B.n756 55.1018
R986 B.n756 B.n755 55.1018
R987 B.n755 B.n23 55.1018
R988 B.n749 B.n23 55.1018
R989 B.n749 B.n748 55.1018
R990 B.n748 B.n747 55.1018
R991 B.n747 B.n30 55.1018
R992 B.n741 B.n30 55.1018
R993 B.n741 B.n740 55.1018
R994 B.n739 B.n37 55.1018
R995 B.n733 B.n37 55.1018
R996 B.n733 B.n732 55.1018
R997 B.n732 B.n731 55.1018
R998 B.n731 B.n44 55.1018
R999 B.n725 B.n44 55.1018
R1000 B.n725 B.n724 55.1018
R1001 B.n724 B.n723 55.1018
R1002 B.n723 B.n51 55.1018
R1003 B.n717 B.n51 55.1018
R1004 B.n717 B.n716 55.1018
R1005 B.n716 B.n715 55.1018
R1006 B.n715 B.n58 55.1018
R1007 B.n709 B.n708 55.1018
R1008 B.n708 B.n707 55.1018
R1009 B.n707 B.n65 55.1018
R1010 B.n701 B.n65 55.1018
R1011 B.n701 B.n700 55.1018
R1012 B.n700 B.n699 55.1018
R1013 B.n699 B.n72 55.1018
R1014 B.n693 B.n72 55.1018
R1015 B.n583 B.t2 36.4646
R1016 B.t3 B.n739 36.4646
R1017 B.n541 B.t5 34.844
R1018 B.n709 B.t12 34.844
R1019 B.n519 B.n331 33.5615
R1020 B.n515 B.n514 33.5615
R1021 B.n690 B.n689 33.5615
R1022 B.n695 B.n74 33.5615
R1023 B.n620 B.t0 28.3615
R1024 B.n763 B.t1 28.3615
R1025 B.n613 B.t0 26.7408
R1026 B.n19 B.t1 26.7408
R1027 B.t5 B.n313 20.2583
R1028 B.t12 B.n58 20.2583
R1029 B.t2 B.n285 18.6377
R1030 B.n740 B.t3 18.6377
R1031 B B.n777 18.0485
R1032 B.n520 B.n519 10.6151
R1033 B.n521 B.n520 10.6151
R1034 B.n521 B.n323 10.6151
R1035 B.n531 B.n323 10.6151
R1036 B.n532 B.n531 10.6151
R1037 B.n533 B.n532 10.6151
R1038 B.n533 B.n315 10.6151
R1039 B.n543 B.n315 10.6151
R1040 B.n544 B.n543 10.6151
R1041 B.n545 B.n544 10.6151
R1042 B.n545 B.n307 10.6151
R1043 B.n555 B.n307 10.6151
R1044 B.n556 B.n555 10.6151
R1045 B.n557 B.n556 10.6151
R1046 B.n557 B.n299 10.6151
R1047 B.n567 B.n299 10.6151
R1048 B.n568 B.n567 10.6151
R1049 B.n569 B.n568 10.6151
R1050 B.n569 B.n291 10.6151
R1051 B.n579 B.n291 10.6151
R1052 B.n580 B.n579 10.6151
R1053 B.n581 B.n580 10.6151
R1054 B.n581 B.n283 10.6151
R1055 B.n591 B.n283 10.6151
R1056 B.n592 B.n591 10.6151
R1057 B.n593 B.n592 10.6151
R1058 B.n593 B.n275 10.6151
R1059 B.n603 B.n275 10.6151
R1060 B.n604 B.n603 10.6151
R1061 B.n605 B.n604 10.6151
R1062 B.n605 B.n267 10.6151
R1063 B.n616 B.n267 10.6151
R1064 B.n617 B.n616 10.6151
R1065 B.n618 B.n617 10.6151
R1066 B.n618 B.n260 10.6151
R1067 B.n629 B.n260 10.6151
R1068 B.n630 B.n629 10.6151
R1069 B.n631 B.n630 10.6151
R1070 B.n631 B.n0 10.6151
R1071 B.n373 B.n331 10.6151
R1072 B.n374 B.n373 10.6151
R1073 B.n375 B.n374 10.6151
R1074 B.n375 B.n369 10.6151
R1075 B.n381 B.n369 10.6151
R1076 B.n382 B.n381 10.6151
R1077 B.n383 B.n382 10.6151
R1078 B.n383 B.n367 10.6151
R1079 B.n389 B.n367 10.6151
R1080 B.n390 B.n389 10.6151
R1081 B.n391 B.n390 10.6151
R1082 B.n391 B.n365 10.6151
R1083 B.n397 B.n365 10.6151
R1084 B.n398 B.n397 10.6151
R1085 B.n399 B.n398 10.6151
R1086 B.n399 B.n363 10.6151
R1087 B.n405 B.n363 10.6151
R1088 B.n406 B.n405 10.6151
R1089 B.n407 B.n406 10.6151
R1090 B.n407 B.n361 10.6151
R1091 B.n413 B.n361 10.6151
R1092 B.n414 B.n413 10.6151
R1093 B.n415 B.n414 10.6151
R1094 B.n415 B.n359 10.6151
R1095 B.n421 B.n359 10.6151
R1096 B.n422 B.n421 10.6151
R1097 B.n423 B.n422 10.6151
R1098 B.n423 B.n357 10.6151
R1099 B.n429 B.n357 10.6151
R1100 B.n430 B.n429 10.6151
R1101 B.n432 B.n353 10.6151
R1102 B.n438 B.n353 10.6151
R1103 B.n439 B.n438 10.6151
R1104 B.n440 B.n439 10.6151
R1105 B.n440 B.n351 10.6151
R1106 B.n446 B.n351 10.6151
R1107 B.n447 B.n446 10.6151
R1108 B.n451 B.n447 10.6151
R1109 B.n457 B.n349 10.6151
R1110 B.n458 B.n457 10.6151
R1111 B.n459 B.n458 10.6151
R1112 B.n459 B.n347 10.6151
R1113 B.n465 B.n347 10.6151
R1114 B.n466 B.n465 10.6151
R1115 B.n467 B.n466 10.6151
R1116 B.n467 B.n345 10.6151
R1117 B.n473 B.n345 10.6151
R1118 B.n474 B.n473 10.6151
R1119 B.n475 B.n474 10.6151
R1120 B.n475 B.n343 10.6151
R1121 B.n481 B.n343 10.6151
R1122 B.n482 B.n481 10.6151
R1123 B.n483 B.n482 10.6151
R1124 B.n483 B.n341 10.6151
R1125 B.n489 B.n341 10.6151
R1126 B.n490 B.n489 10.6151
R1127 B.n491 B.n490 10.6151
R1128 B.n491 B.n339 10.6151
R1129 B.n497 B.n339 10.6151
R1130 B.n498 B.n497 10.6151
R1131 B.n499 B.n498 10.6151
R1132 B.n499 B.n337 10.6151
R1133 B.n505 B.n337 10.6151
R1134 B.n506 B.n505 10.6151
R1135 B.n507 B.n506 10.6151
R1136 B.n507 B.n335 10.6151
R1137 B.n513 B.n335 10.6151
R1138 B.n514 B.n513 10.6151
R1139 B.n515 B.n327 10.6151
R1140 B.n525 B.n327 10.6151
R1141 B.n526 B.n525 10.6151
R1142 B.n527 B.n526 10.6151
R1143 B.n527 B.n319 10.6151
R1144 B.n537 B.n319 10.6151
R1145 B.n538 B.n537 10.6151
R1146 B.n539 B.n538 10.6151
R1147 B.n539 B.n311 10.6151
R1148 B.n549 B.n311 10.6151
R1149 B.n550 B.n549 10.6151
R1150 B.n551 B.n550 10.6151
R1151 B.n551 B.n303 10.6151
R1152 B.n561 B.n303 10.6151
R1153 B.n562 B.n561 10.6151
R1154 B.n563 B.n562 10.6151
R1155 B.n563 B.n295 10.6151
R1156 B.n573 B.n295 10.6151
R1157 B.n574 B.n573 10.6151
R1158 B.n575 B.n574 10.6151
R1159 B.n575 B.n287 10.6151
R1160 B.n585 B.n287 10.6151
R1161 B.n586 B.n585 10.6151
R1162 B.n587 B.n586 10.6151
R1163 B.n587 B.n279 10.6151
R1164 B.n597 B.n279 10.6151
R1165 B.n598 B.n597 10.6151
R1166 B.n599 B.n598 10.6151
R1167 B.n599 B.n271 10.6151
R1168 B.n609 B.n271 10.6151
R1169 B.n610 B.n609 10.6151
R1170 B.n611 B.n610 10.6151
R1171 B.n611 B.n264 10.6151
R1172 B.n622 B.n264 10.6151
R1173 B.n623 B.n622 10.6151
R1174 B.n625 B.n623 10.6151
R1175 B.n625 B.n624 10.6151
R1176 B.n624 B.n256 10.6151
R1177 B.n636 B.n256 10.6151
R1178 B.n637 B.n636 10.6151
R1179 B.n638 B.n637 10.6151
R1180 B.n639 B.n638 10.6151
R1181 B.n640 B.n639 10.6151
R1182 B.n643 B.n640 10.6151
R1183 B.n644 B.n643 10.6151
R1184 B.n645 B.n644 10.6151
R1185 B.n646 B.n645 10.6151
R1186 B.n648 B.n646 10.6151
R1187 B.n649 B.n648 10.6151
R1188 B.n650 B.n649 10.6151
R1189 B.n651 B.n650 10.6151
R1190 B.n653 B.n651 10.6151
R1191 B.n654 B.n653 10.6151
R1192 B.n655 B.n654 10.6151
R1193 B.n656 B.n655 10.6151
R1194 B.n658 B.n656 10.6151
R1195 B.n659 B.n658 10.6151
R1196 B.n660 B.n659 10.6151
R1197 B.n661 B.n660 10.6151
R1198 B.n663 B.n661 10.6151
R1199 B.n664 B.n663 10.6151
R1200 B.n665 B.n664 10.6151
R1201 B.n666 B.n665 10.6151
R1202 B.n668 B.n666 10.6151
R1203 B.n669 B.n668 10.6151
R1204 B.n670 B.n669 10.6151
R1205 B.n671 B.n670 10.6151
R1206 B.n673 B.n671 10.6151
R1207 B.n674 B.n673 10.6151
R1208 B.n675 B.n674 10.6151
R1209 B.n676 B.n675 10.6151
R1210 B.n678 B.n676 10.6151
R1211 B.n679 B.n678 10.6151
R1212 B.n680 B.n679 10.6151
R1213 B.n681 B.n680 10.6151
R1214 B.n683 B.n681 10.6151
R1215 B.n684 B.n683 10.6151
R1216 B.n685 B.n684 10.6151
R1217 B.n686 B.n685 10.6151
R1218 B.n688 B.n686 10.6151
R1219 B.n689 B.n688 10.6151
R1220 B.n769 B.n1 10.6151
R1221 B.n769 B.n768 10.6151
R1222 B.n768 B.n767 10.6151
R1223 B.n767 B.n10 10.6151
R1224 B.n761 B.n10 10.6151
R1225 B.n761 B.n760 10.6151
R1226 B.n760 B.n759 10.6151
R1227 B.n759 B.n17 10.6151
R1228 B.n753 B.n17 10.6151
R1229 B.n753 B.n752 10.6151
R1230 B.n752 B.n751 10.6151
R1231 B.n751 B.n25 10.6151
R1232 B.n745 B.n25 10.6151
R1233 B.n745 B.n744 10.6151
R1234 B.n744 B.n743 10.6151
R1235 B.n743 B.n32 10.6151
R1236 B.n737 B.n32 10.6151
R1237 B.n737 B.n736 10.6151
R1238 B.n736 B.n735 10.6151
R1239 B.n735 B.n39 10.6151
R1240 B.n729 B.n39 10.6151
R1241 B.n729 B.n728 10.6151
R1242 B.n728 B.n727 10.6151
R1243 B.n727 B.n46 10.6151
R1244 B.n721 B.n46 10.6151
R1245 B.n721 B.n720 10.6151
R1246 B.n720 B.n719 10.6151
R1247 B.n719 B.n53 10.6151
R1248 B.n713 B.n53 10.6151
R1249 B.n713 B.n712 10.6151
R1250 B.n712 B.n711 10.6151
R1251 B.n711 B.n60 10.6151
R1252 B.n705 B.n60 10.6151
R1253 B.n705 B.n704 10.6151
R1254 B.n704 B.n703 10.6151
R1255 B.n703 B.n67 10.6151
R1256 B.n697 B.n67 10.6151
R1257 B.n697 B.n696 10.6151
R1258 B.n696 B.n695 10.6151
R1259 B.n118 B.n74 10.6151
R1260 B.n121 B.n118 10.6151
R1261 B.n122 B.n121 10.6151
R1262 B.n125 B.n122 10.6151
R1263 B.n126 B.n125 10.6151
R1264 B.n129 B.n126 10.6151
R1265 B.n130 B.n129 10.6151
R1266 B.n133 B.n130 10.6151
R1267 B.n134 B.n133 10.6151
R1268 B.n137 B.n134 10.6151
R1269 B.n138 B.n137 10.6151
R1270 B.n141 B.n138 10.6151
R1271 B.n142 B.n141 10.6151
R1272 B.n145 B.n142 10.6151
R1273 B.n146 B.n145 10.6151
R1274 B.n149 B.n146 10.6151
R1275 B.n150 B.n149 10.6151
R1276 B.n153 B.n150 10.6151
R1277 B.n154 B.n153 10.6151
R1278 B.n157 B.n154 10.6151
R1279 B.n158 B.n157 10.6151
R1280 B.n161 B.n158 10.6151
R1281 B.n162 B.n161 10.6151
R1282 B.n165 B.n162 10.6151
R1283 B.n166 B.n165 10.6151
R1284 B.n169 B.n166 10.6151
R1285 B.n170 B.n169 10.6151
R1286 B.n173 B.n170 10.6151
R1287 B.n174 B.n173 10.6151
R1288 B.n177 B.n174 10.6151
R1289 B.n182 B.n179 10.6151
R1290 B.n183 B.n182 10.6151
R1291 B.n186 B.n183 10.6151
R1292 B.n187 B.n186 10.6151
R1293 B.n190 B.n187 10.6151
R1294 B.n191 B.n190 10.6151
R1295 B.n194 B.n191 10.6151
R1296 B.n195 B.n194 10.6151
R1297 B.n199 B.n198 10.6151
R1298 B.n202 B.n199 10.6151
R1299 B.n203 B.n202 10.6151
R1300 B.n206 B.n203 10.6151
R1301 B.n207 B.n206 10.6151
R1302 B.n210 B.n207 10.6151
R1303 B.n211 B.n210 10.6151
R1304 B.n214 B.n211 10.6151
R1305 B.n215 B.n214 10.6151
R1306 B.n218 B.n215 10.6151
R1307 B.n219 B.n218 10.6151
R1308 B.n222 B.n219 10.6151
R1309 B.n223 B.n222 10.6151
R1310 B.n226 B.n223 10.6151
R1311 B.n227 B.n226 10.6151
R1312 B.n230 B.n227 10.6151
R1313 B.n231 B.n230 10.6151
R1314 B.n234 B.n231 10.6151
R1315 B.n235 B.n234 10.6151
R1316 B.n238 B.n235 10.6151
R1317 B.n239 B.n238 10.6151
R1318 B.n242 B.n239 10.6151
R1319 B.n243 B.n242 10.6151
R1320 B.n246 B.n243 10.6151
R1321 B.n247 B.n246 10.6151
R1322 B.n250 B.n247 10.6151
R1323 B.n251 B.n250 10.6151
R1324 B.n254 B.n251 10.6151
R1325 B.n255 B.n254 10.6151
R1326 B.n690 B.n255 10.6151
R1327 B.n777 B.n0 8.11757
R1328 B.n777 B.n1 8.11757
R1329 B.n432 B.n431 6.5566
R1330 B.n451 B.n450 6.5566
R1331 B.n179 B.n178 6.5566
R1332 B.n195 B.n115 6.5566
R1333 B.n431 B.n430 4.05904
R1334 B.n450 B.n349 4.05904
R1335 B.n178 B.n177 4.05904
R1336 B.n198 B.n115 4.05904
R1337 VP.n17 VP.n16 161.3
R1338 VP.n15 VP.n1 161.3
R1339 VP.n14 VP.n13 161.3
R1340 VP.n12 VP.n2 161.3
R1341 VP.n11 VP.n10 161.3
R1342 VP.n9 VP.n3 161.3
R1343 VP.n8 VP.n7 161.3
R1344 VP.n5 VP.t1 94.6782
R1345 VP.n5 VP.t3 93.5485
R1346 VP.n6 VP.n4 73.3375
R1347 VP.n18 VP.n0 73.3375
R1348 VP.n4 VP.t0 59.7109
R1349 VP.n0 VP.t2 59.7109
R1350 VP.n6 VP.n5 48.3428
R1351 VP.n10 VP.n2 40.4106
R1352 VP.n14 VP.n2 40.4106
R1353 VP.n9 VP.n8 24.3439
R1354 VP.n10 VP.n9 24.3439
R1355 VP.n15 VP.n14 24.3439
R1356 VP.n16 VP.n15 24.3439
R1357 VP.n8 VP.n4 16.554
R1358 VP.n16 VP.n0 16.554
R1359 VP.n7 VP.n6 0.355081
R1360 VP.n18 VP.n17 0.355081
R1361 VP VP.n18 0.26685
R1362 VP.n7 VP.n3 0.189894
R1363 VP.n11 VP.n3 0.189894
R1364 VP.n12 VP.n11 0.189894
R1365 VP.n13 VP.n12 0.189894
R1366 VP.n13 VP.n1 0.189894
R1367 VP.n17 VP.n1 0.189894
R1368 VDD1 VDD1.n1 107.323
R1369 VDD1 VDD1.n0 66.4689
R1370 VDD1.n0 VDD1.t2 2.38604
R1371 VDD1.n0 VDD1.t1 2.38604
R1372 VDD1.n1 VDD1.t3 2.38604
R1373 VDD1.n1 VDD1.t0 2.38604
R1374 VTAIL.n5 VTAIL.t6 52.1175
R1375 VTAIL.n4 VTAIL.t2 52.1175
R1376 VTAIL.n3 VTAIL.t0 52.1175
R1377 VTAIL.n6 VTAIL.t4 52.1175
R1378 VTAIL.n7 VTAIL.t3 52.1175
R1379 VTAIL.n0 VTAIL.t1 52.1175
R1380 VTAIL.n1 VTAIL.t5 52.1175
R1381 VTAIL.n2 VTAIL.t7 52.1175
R1382 VTAIL.n7 VTAIL.n6 22.6945
R1383 VTAIL.n3 VTAIL.n2 22.6945
R1384 VTAIL.n4 VTAIL.n3 3.17291
R1385 VTAIL.n6 VTAIL.n5 3.17291
R1386 VTAIL.n2 VTAIL.n1 3.17291
R1387 VTAIL VTAIL.n0 1.6449
R1388 VTAIL VTAIL.n7 1.52852
R1389 VTAIL.n5 VTAIL.n4 0.470328
R1390 VTAIL.n1 VTAIL.n0 0.470328
R1391 VN.n1 VN.t1 94.6784
R1392 VN.n0 VN.t2 94.6784
R1393 VN.n0 VN.t0 93.5485
R1394 VN.n1 VN.t3 93.5485
R1395 VN VN.n1 48.5083
R1396 VN VN.n0 2.42873
R1397 VDD2.n2 VDD2.n0 106.797
R1398 VDD2.n2 VDD2.n1 66.4107
R1399 VDD2.n1 VDD2.t0 2.38604
R1400 VDD2.n1 VDD2.t2 2.38604
R1401 VDD2.n0 VDD2.t1 2.38604
R1402 VDD2.n0 VDD2.t3 2.38604
R1403 VDD2 VDD2.n2 0.0586897
C0 VDD2 VN 3.52559f
C1 VTAIL VP 3.72933f
C2 VTAIL VDD1 4.78884f
C3 VDD2 VP 0.441542f
C4 VDD1 VDD2 1.20037f
C5 VTAIL VDD2 4.84807f
C6 VP VN 6.04959f
C7 VDD1 VN 0.14919f
C8 VDD1 VP 3.81702f
C9 VTAIL VN 3.71523f
C10 VDD2 B 3.913141f
C11 VDD1 B 8.00293f
C12 VTAIL B 8.253065f
C13 VN B 11.8735f
C14 VP B 10.289506f
C15 VDD2.t1 B 0.179653f
C16 VDD2.t3 B 0.179653f
C17 VDD2.n0 B 2.12808f
C18 VDD2.t0 B 0.179653f
C19 VDD2.t2 B 0.179653f
C20 VDD2.n1 B 1.56145f
C21 VDD2.n2 B 3.60596f
C22 VN.t0 B 1.99905f
C23 VN.t2 B 2.00811f
C24 VN.n0 B 1.18993f
C25 VN.t3 B 1.99905f
C26 VN.t1 B 2.00811f
C27 VN.n1 B 2.51414f
C28 VTAIL.t1 B 1.2704f
C29 VTAIL.n0 B 0.348575f
C30 VTAIL.t5 B 1.2704f
C31 VTAIL.n1 B 0.438854f
C32 VTAIL.t7 B 1.2704f
C33 VTAIL.n2 B 1.27035f
C34 VTAIL.t0 B 1.27041f
C35 VTAIL.n3 B 1.27034f
C36 VTAIL.t2 B 1.27041f
C37 VTAIL.n4 B 0.438845f
C38 VTAIL.t6 B 1.27041f
C39 VTAIL.n5 B 0.438845f
C40 VTAIL.t4 B 1.2704f
C41 VTAIL.n6 B 1.27035f
C42 VTAIL.t3 B 1.2704f
C43 VTAIL.n7 B 1.17319f
C44 VDD1.t2 B 0.183905f
C45 VDD1.t1 B 0.183905f
C46 VDD1.n0 B 1.59887f
C47 VDD1.t3 B 0.183905f
C48 VDD1.t0 B 0.183905f
C49 VDD1.n1 B 2.20437f
C50 VP.t2 B 1.75804f
C51 VP.n0 B 0.729724f
C52 VP.n1 B 0.023505f
C53 VP.n2 B 0.019021f
C54 VP.n3 B 0.023505f
C55 VP.t0 B 1.75804f
C56 VP.n4 B 0.729724f
C57 VP.t1 B 2.05877f
C58 VP.t3 B 2.04949f
C59 VP.n5 B 2.56791f
C60 VP.n6 B 1.27307f
C61 VP.n7 B 0.037943f
C62 VP.n8 B 0.037072f
C63 VP.n9 B 0.044028f
C64 VP.n10 B 0.046966f
C65 VP.n11 B 0.023505f
C66 VP.n12 B 0.023505f
C67 VP.n13 B 0.023505f
C68 VP.n14 B 0.046966f
C69 VP.n15 B 0.044028f
C70 VP.n16 B 0.037072f
C71 VP.n17 B 0.037943f
C72 VP.n18 B 0.055446f
.ends

