* NGSPICE file created from opamp_sample_0004.ext - technology: sky130A

.subckt opamp_sample_0004 GND VOUT VDD VN VP CS_BIAS DIFFPAIR_BIAS
X0 a_n18640_8567.t19 a_n7837_10186.t28 a_n5326_8245.t15 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X1 VDD.t157 a_n7837_10186.t29 a_n5326_8245.t12 VDD.t156 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X2 GND.t266 CS_BIAS.t32 VOUT.t10 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X3 GND.t154 GND.t151 GND.t153 GND.t152 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=0 ps=0 w=4.85 l=2.45
X4 CS_BIAS.t19 CS_BIAS.t18 GND.t265 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X5 a_n7837_10186.t8 VP.t6 a_n7336_n129.t20 GND.t3 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X6 VDD.t69 VDD.t67 VDD.t68 VDD.t10 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X7 GND.t150 GND.t148 VP.t5 GND.t149 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X8 a_n18640_8567.t2 VN.t6 a_n7336_n129.t2 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=3.9168 ps=12.32 w=5.44 l=5.27
X9 VOUT.t116 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X10 GND.t147 GND.t145 GND.t146 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X11 VDD.t66 VDD.t64 VDD.t65 VDD.t10 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X12 GND.t264 CS_BIAS.t33 VOUT.t51 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X13 a_n7336_n129.t8 DIFFPAIR_BIAS.t8 GND.t14 GND.t13 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
X14 VOUT.t50 CS_BIAS.t34 GND.t263 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X15 VOUT.t49 CS_BIAS.t35 GND.t262 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X16 VOUT.t48 CS_BIAS.t36 GND.t261 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X17 a_n7336_n129.t19 VP.t7 a_n7837_10186.t9 GND.t267 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X18 a_n7837_10186.t1 VP.t8 a_n7336_n129.t18 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X19 GND.t144 GND.t142 GND.t143 GND.t97 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=0 ps=0 w=5.44 l=5.27
X20 GND.t260 CS_BIAS.t37 VOUT.t47 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X21 CS_BIAS.t17 CS_BIAS.t16 GND.t259 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X22 GND.t141 GND.t139 GND.t140 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X23 GND.t258 CS_BIAS.t14 CS_BIAS.t15 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X24 GND.t257 CS_BIAS.t38 VOUT.t46 GND.t187 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X25 a_n7336_n129.t7 DIFFPAIR_BIAS.t9 GND.t12 GND.t11 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
X26 VOUT.t45 CS_BIAS.t39 GND.t256 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X27 a_8109_10383# a_8109_10383# a_8109_10383# VDD.t1 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=7.416 ps=23.48 w=5.15 l=3.71
X28 GND.t138 GND.t136 GND.t137 GND.t45 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X29 GND.t135 GND.t133 GND.t134 GND.t45 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X30 VDD.t63 VDD.t61 VDD.t62 VDD.t58 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X31 GND.t132 GND.t130 GND.t131 GND.t30 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X32 GND.t255 CS_BIAS.t40 VOUT.t44 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X33 a_n5326_8245.t11 a_n7837_10186.t30 VDD.t155 VDD.t154 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X34 VOUT.t43 CS_BIAS.t41 GND.t254 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X35 VDD.t153 a_n7837_10186.t31 a_n5326_8245.t3 VDD.t152 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X36 a_n7837_10186.t22 a_n7837_10186.t21 a_n7981_10383.t15 VDD.t143 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X37 GND.t129 GND.t127 VN.t5 GND.t128 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X38 GND.t126 GND.t124 VP.t4 GND.t125 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X39 GND.t123 GND.t121 GND.t122 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X40 a_n7981_10383.t7 a_n7837_10186.t32 VDD.t151 VDD.t150 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X41 VOUT.t115 a_n18640_8567.t20 VDD.t117 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X42 GND.t253 CS_BIAS.t42 VOUT.t42 GND.t187 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X43 VOUT.t114 a_n18640_8567.t21 VDD.t116 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X44 GND.t252 CS_BIAS.t43 VOUT.t41 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X45 a_n7336_n129.t4 VN.t7 a_n18640_8567.t4 GND.t7 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X46 VOUT.t40 CS_BIAS.t44 GND.t251 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X47 VDD.t60 VDD.t57 VDD.t59 VDD.t58 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X48 GND.t250 CS_BIAS.t45 VOUT.t39 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X49 VOUT.t37 CS_BIAS.t46 GND.t247 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X50 GND.t249 CS_BIAS.t47 VOUT.t38 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X51 GND.t248 CS_BIAS.t12 CS_BIAS.t13 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X52 GND.t246 CS_BIAS.t48 VOUT.t36 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X53 CS_BIAS.t11 CS_BIAS.t10 GND.t245 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X54 GND.t244 CS_BIAS.t49 VOUT.t35 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X55 GND.t235 CS_BIAS.t50 VOUT.t27 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X56 GND.t243 CS_BIAS.t51 VOUT.t34 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X57 GND.t120 GND.t118 GND.t119 GND.t30 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X58 VOUT.t33 CS_BIAS.t52 GND.t242 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X59 VOUT.t32 CS_BIAS.t53 GND.t241 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X60 VOUT.t31 CS_BIAS.t54 GND.t240 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X61 VDD.t56 VDD.t54 VDD.t55 VDD.t41 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X62 GND.t117 GND.t115 GND.t116 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X63 VDD.t53 VDD.t51 VDD.t52 VDD.t48 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X64 VDD.t149 a_n7837_10186.t33 a_n7981_10383.t6 VDD.t148 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X65 VOUT.t117 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X66 a_n5326_8245.t4 a_n7837_10186.t34 VDD.t147 VDD.t146 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X67 GND.t114 GND.t112 VN.t4 GND.t113 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X68 GND.t239 CS_BIAS.t55 VOUT.t30 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X69 GND.t238 CS_BIAS.t56 VOUT.t29 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X70 a_n7336_n129.t17 VP.t9 a_n7837_10186.t6 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X71 a_n7837_10186.t3 VP.t10 a_n7336_n129.t16 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X72 DIFFPAIR_BIAS.t7 DIFFPAIR_BIAS.t6 GND.t19 GND.t18 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
X73 VOUT.t113 a_n18640_8567.t22 VDD.t115 VDD.t99 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=3.4992 ps=11.16 w=4.86 l=5.24
X74 VOUT.t112 a_n18640_8567.t23 VDD.t114 VDD.t99 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=3.4992 ps=11.16 w=4.86 l=5.24
X75 a_n7981_10383.t14 a_n7837_10186.t11 a_n7837_10186.t12 VDD.t142 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X76 CS_BIAS.t9 CS_BIAS.t8 GND.t237 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X77 a_n18640_8567.t18 a_n7837_10186.t35 a_n5326_8245.t5 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X78 VOUT.t26 CS_BIAS.t57 GND.t234 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X79 GND.t236 CS_BIAS.t58 VOUT.t28 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X80 VDD.t113 a_n18640_8567.t24 VOUT.t111 VDD.t81 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=1.6038 ps=5.52 w=4.86 l=5.24
X81 VDD.t145 a_n7837_10186.t36 a_n7981_10383.t5 VDD.t144 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X82 CS_BIAS.t7 CS_BIAS.t6 GND.t233 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X83 VDD.t112 a_n18640_8567.t25 VOUT.t110 VDD.t81 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=1.6038 ps=5.52 w=4.86 l=5.24
X84 GND.t111 GND.t109 GND.t110 GND.t45 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X85 GND.t108 GND.t106 GND.t107 GND.t26 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=0 ps=0 w=5.44 l=5.27
X86 VDD.t50 VDD.t47 VDD.t49 VDD.t48 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X87 VOUT.t25 CS_BIAS.t59 GND.t232 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X88 a_n9139_10383# a_n9139_10383# a_n9139_10383# VDD.t0 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=7.416 ps=23.48 w=5.15 l=3.71
X89 GND.t105 GND.t103 VP.t3 GND.t104 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X90 VOUT.t24 CS_BIAS.t60 GND.t231 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X91 a_n7837_10186.t0 VP.t11 a_n7336_n129.t15 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=3.9168 ps=12.32 w=5.44 l=5.27
X92 a_n7336_n129.t14 VP.t12 a_n7837_10186.t27 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X93 VOUT.t23 CS_BIAS.t61 GND.t230 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X94 a_n5326_8245.t13 a_n7837_10186.t37 a_n18640_8567.t17 VDD.t143 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X95 VOUT.t109 a_n18640_8567.t26 VDD.t111 VDD.t110 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X96 GND.t102 GND.t100 GND.t101 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X97 VDD.t107 a_n18640_8567.t27 VOUT.t108 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X98 VOUT.t22 CS_BIAS.t62 GND.t229 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X99 VOUT.t21 CS_BIAS.t63 GND.t228 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X100 a_n18640_8567.t16 a_n7837_10186.t38 a_n5326_8245.t10 VDD.t142 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X101 VOUT.t107 a_n18640_8567.t28 VDD.t109 VDD.t85 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X102 a_n18640_8567.t7 VN.t8 a_n7336_n129.t21 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X103 VOUT.t118 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X104 VOUT.t20 CS_BIAS.t64 GND.t227 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X105 GND.t226 CS_BIAS.t65 VOUT.t19 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X106 a_n5326_8245.t6 a_n7837_10186.t39 a_n18640_8567.t15 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X107 GND.t92 GND.t90 VN.t3 GND.t91 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.39 ps=2.78 w=1 l=0.5
X108 GND.t95 GND.t93 GND.t94 GND.t30 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X109 a_n7837_10186.t4 VP.t13 a_n7336_n129.t13 GND.t4 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=3.9168 ps=12.32 w=5.44 l=5.27
X110 GND.t225 CS_BIAS.t66 VOUT.t18 GND.t187 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X111 GND.t224 CS_BIAS.t67 VOUT.t17 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X112 GND.t223 CS_BIAS.t68 VOUT.t16 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X113 VOUT.t15 CS_BIAS.t69 GND.t222 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X114 VDD.t108 a_n18640_8567.t29 VOUT.t106 VDD.t103 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X115 VDD.t106 a_n18640_8567.t30 VOUT.t105 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X116 a_n18640_8567.t11 VN.t9 a_n7336_n129.t25 GND.t9 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X117 VOUT.t14 CS_BIAS.t70 GND.t221 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X118 VDD.t105 a_n18640_8567.t31 VOUT.t104 VDD.t103 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X119 VDD.t98 a_n18640_8567.t32 VOUT.t103 VDD.t97 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X120 VDD.t104 a_n18640_8567.t33 VOUT.t102 VDD.t103 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X121 GND.t99 GND.t96 GND.t98 GND.t97 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=0 ps=0 w=5.44 l=5.27
X122 VN.t2 GND.t87 GND.t89 GND.t88 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X123 VOUT.t13 CS_BIAS.t71 GND.t220 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X124 VOUT.t9 CS_BIAS.t72 GND.t164 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X125 GND.t219 CS_BIAS.t73 VOUT.t12 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X126 VOUT.t101 a_n18640_8567.t34 VDD.t102 VDD.t83 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X127 a_n7336_n129.t22 VN.t10 a_n18640_8567.t8 GND.t17 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=1.7952 ps=6.1 w=5.44 l=5.27
X128 a_n5326_8245.t9 a_n7837_10186.t40 a_n18640_8567.t14 VDD.t136 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X129 GND.t218 CS_BIAS.t74 VOUT.t11 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X130 VDD.t141 a_n7837_10186.t41 a_n5326_8245.t2 VDD.t140 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X131 GND.t86 GND.t84 GND.t85 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X132 GND.t217 CS_BIAS.t75 VOUT.t61 GND.t187 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X133 VDD.t101 a_n18640_8567.t35 VOUT.t100 VDD.t70 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X134 VOUT.t56 CS_BIAS.t76 GND.t211 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X135 a_n7837_10186.t24 a_n7837_10186.t23 a_n7981_10383.t13 VDD.t127 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X136 GND.t216 CS_BIAS.t77 VOUT.t60 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X137 a_n7981_10383.t12 a_n7837_10186.t25 a_n7837_10186.t26 VDD.t139 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X138 VOUT.t59 CS_BIAS.t78 GND.t215 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X139 GND.t83 GND.t81 GND.t82 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X140 VOUT.t99 a_n18640_8567.t36 VDD.t100 VDD.t99 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=3.4992 ps=11.16 w=4.86 l=5.24
X141 DIFFPAIR_BIAS.t5 DIFFPAIR_BIAS.t4 GND.t2 GND.t1 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
X142 VDD.t138 a_n7837_10186.t42 a_n5326_8245.t1 VDD.t137 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X143 VOUT.t119 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X144 a_n7837_10186.t18 a_n7837_10186.t17 a_n7981_10383.t11 VDD.t136 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X145 a_n7981_10383.t4 a_n7837_10186.t43 VDD.t135 VDD.t134 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X146 GND.t214 CS_BIAS.t22 CS_BIAS.t23 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X147 GND.t213 CS_BIAS.t79 VOUT.t58 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X148 a_n7336_n129.t12 VP.t14 a_n7837_10186.t2 GND.t10 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=1.7952 ps=6.1 w=5.44 l=5.27
X149 VN.t1 GND.t78 GND.t80 GND.t79 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X150 VOUT.t120 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X151 VOUT.t57 CS_BIAS.t80 GND.t212 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X152 GND.t210 CS_BIAS.t20 CS_BIAS.t21 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X153 GND.t77 GND.t75 GND.t76 GND.t45 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X154 VDD.t46 VDD.t44 VDD.t45 VDD.t3 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X155 VOUT.t98 a_n18640_8567.t37 VDD.t96 VDD.t79 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X156 VOUT.t97 a_n18640_8567.t38 VDD.t95 VDD.t79 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X157 VOUT.t55 CS_BIAS.t81 GND.t209 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X158 GND.t74 GND.t72 GND.t73 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X159 VDD.t43 VDD.t40 VDD.t42 VDD.t41 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X160 a_n18640_8567.t1 VN.t11 a_n7336_n129.t1 GND.t3 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X161 VOUT.t121 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X162 a_n7336_n129.t27 DIFFPAIR_BIAS.t10 GND.t273 GND.t272 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
X163 VDD.t39 VDD.t37 VDD.t38 VDD.t22 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X164 VOUT.t54 CS_BIAS.t82 GND.t208 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X165 VDD.t36 VDD.t34 VDD.t35 VDD.t22 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X166 VOUT.t53 CS_BIAS.t83 GND.t207 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X167 a_n5326_8245.t14 a_n7837_10186.t44 VDD.t133 VDD.t132 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X168 VDD.t94 a_n18640_8567.t39 VOUT.t96 VDD.t91 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=1.6038 ps=5.52 w=4.86 l=5.24
X169 VP.t2 GND.t69 GND.t71 GND.t70 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X170 GND.t68 GND.t66 GND.t67 GND.t30 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X171 a_n18640_8567.t0 VN.t12 a_n7336_n129.t0 GND.t0 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X172 a_n7336_n129.t24 VN.t13 a_n18640_8567.t10 GND.t267 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X173 GND.t206 CS_BIAS.t84 VOUT.t52 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X174 VDD.t93 a_n18640_8567.t40 VOUT.t95 VDD.t91 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=1.6038 ps=5.52 w=4.86 l=5.24
X175 VOUT.t70 CS_BIAS.t85 GND.t205 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X176 VDD.t92 a_n18640_8567.t41 VOUT.t94 VDD.t91 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=1.6038 ps=5.52 w=4.86 l=5.24
X177 GND.t199 CS_BIAS.t86 VOUT.t66 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X178 VOUT.t69 CS_BIAS.t87 GND.t204 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X179 GND.t203 CS_BIAS.t88 VOUT.t68 GND.t187 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X180 CS_BIAS.t29 CS_BIAS.t28 GND.t202 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X181 CS_BIAS.t27 CS_BIAS.t26 GND.t201 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X182 GND.t200 CS_BIAS.t89 VOUT.t67 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X183 GND.t198 CS_BIAS.t90 VOUT.t65 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X184 GND.t197 CS_BIAS.t24 CS_BIAS.t25 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X185 GND.t196 CS_BIAS.t91 VOUT.t64 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X186 VOUT.t63 CS_BIAS.t92 GND.t195 GND.t194 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X187 VOUT.t93 a_n18640_8567.t42 VDD.t90 VDD.t77 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=3.4992 ps=11.16 w=4.86 l=5.24
X188 VOUT.t92 a_n18640_8567.t43 VDD.t89 VDD.t77 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=3.4992 ps=11.16 w=4.86 l=5.24
X189 GND.t65 GND.t63 GND.t64 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X190 VOUT.t91 a_n18640_8567.t44 VDD.t88 VDD.t85 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X191 VP.t1 GND.t60 GND.t62 GND.t61 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X192 VOUT.t62 CS_BIAS.t93 GND.t193 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X193 VOUT.t79 CS_BIAS.t94 GND.t192 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X194 GND.t191 CS_BIAS.t95 VOUT.t78 GND.t190 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X195 VOUT.t90 a_n18640_8567.t45 VDD.t87 VDD.t83 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X196 VOUT.t89 a_n18640_8567.t46 VDD.t86 VDD.t85 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X197 VOUT.t88 a_n18640_8567.t47 VDD.t84 VDD.t83 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X198 a_n7981_10383.t3 a_n7837_10186.t45 VDD.t131 VDD.t130 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X199 a_n5326_8245.t8 a_n7837_10186.t46 VDD.t129 VDD.t128 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X200 GND.t189 CS_BIAS.t96 VOUT.t77 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X201 GND.t188 CS_BIAS.t30 CS_BIAS.t31 GND.t187 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X202 VOUT.t76 CS_BIAS.t97 GND.t186 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X203 GND.t59 GND.t57 GND.t58 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X204 a_n18640_8567.t13 a_n7837_10186.t47 a_n5326_8245.t7 VDD.t120 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X205 a_n18640_8567.t5 VN.t14 a_n7336_n129.t5 GND.t6 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=3.9168 ps=12.32 w=5.44 l=5.27
X206 a_n7336_n129.t3 VN.t15 a_n18640_8567.t3 GND.t5 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X207 VOUT.t75 CS_BIAS.t98 GND.t185 GND.t163 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X208 GND.t56 GND.t54 GND.t55 GND.t45 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X209 GND.t184 CS_BIAS.t99 VOUT.t74 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X210 VOUT.t73 CS_BIAS.t100 GND.t183 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X211 a_n5326_8245.t16 a_n7837_10186.t48 a_n18640_8567.t12 VDD.t127 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X212 VDD.t33 VDD.t31 VDD.t32 VDD.t18 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X213 a_n7336_n129.t11 VP.t15 a_n7837_10186.t10 GND.t7 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X214 a_n7837_10186.t7 VP.t16 a_n7336_n129.t10 GND.t20 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X215 VDD.t126 a_n7837_10186.t49 a_n7981_10383.t2 VDD.t125 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X216 VDD.t82 a_n18640_8567.t48 VOUT.t87 VDD.t81 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=1.6038 ps=5.52 w=4.86 l=5.24
X217 VOUT.t86 a_n18640_8567.t49 VDD.t80 VDD.t79 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X218 a_n7837_10186.t14 a_n7837_10186.t13 a_n7981_10383.t10 VDD.t124 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X219 VOUT.t72 CS_BIAS.t101 GND.t182 GND.t181 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X220 GND.t180 CS_BIAS.t102 VOUT.t71 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X221 GND.t179 CS_BIAS.t2 CS_BIAS.t3 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X222 VN.t0 GND.t51 GND.t53 GND.t52 sky130_fd_pr__nfet_01v8 ad=0.165 pd=1.33 as=0.165 ps=1.33 w=1 l=0.5
X223 VDD.t30 VDD.t28 VDD.t29 VDD.t14 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X224 VDD.t27 VDD.t25 VDD.t26 VDD.t14 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X225 a_n7981_10383.t9 a_n7837_10186.t19 a_n7837_10186.t20 VDD.t123 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X226 VP.t0 GND.t48 GND.t50 GND.t49 sky130_fd_pr__nfet_01v8 ad=0.39 pd=2.78 as=0.165 ps=1.33 w=1 l=0.5
X227 a_n7336_n129.t9 VP.t17 a_n7837_10186.t5 GND.t17 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=1.7952 ps=6.1 w=5.44 l=5.27
X228 VDD.t24 VDD.t21 VDD.t23 VDD.t22 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X229 GND.t47 GND.t44 GND.t46 GND.t45 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X230 VDD.t20 VDD.t17 VDD.t19 VDD.t18 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=0 ps=0 w=5.15 l=3.71
X231 VDD.t122 a_n7837_10186.t50 a_n7981_10383.t1 VDD.t121 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=3.708 ps=11.74 w=5.15 l=3.71
X232 a_n7336_n129.t26 DIFFPAIR_BIAS.t11 GND.t271 GND.t270 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
X233 VDD.t16 VDD.t13 VDD.t15 VDD.t14 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X234 GND.t43 GND.t40 GND.t42 GND.t41 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=0 ps=0 w=4.85 l=2.45
X235 GND.t39 GND.t37 GND.t38 GND.t30 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X236 GND.t36 GND.t33 GND.t35 GND.t34 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X237 a_n7981_10383.t8 a_n7837_10186.t15 a_n7837_10186.t16 VDD.t120 sky130_fd_pr__pfet_01v8 ad=1.6995 pd=5.81 as=1.6995 ps=5.81 w=5.15 l=3.71
X238 a_n7336_n129.t6 VN.t16 a_n18640_8567.t6 GND.t8 sky130_fd_pr__nfet_01v8 ad=1.7952 pd=6.1 as=1.7952 ps=6.1 w=5.44 l=5.27
X239 GND.t178 CS_BIAS.t103 VOUT.t5 GND.t177 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X240 VOUT.t3 CS_BIAS.t104 GND.t174 GND.t173 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X241 GND.t176 CS_BIAS.t105 VOUT.t4 GND.t175 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X242 GND.t32 GND.t29 GND.t31 GND.t30 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X243 GND.t172 CS_BIAS.t0 CS_BIAS.t1 GND.t171 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0.9207 ps=3.45 w=2.79 l=5.03
X244 GND.t170 CS_BIAS.t106 VOUT.t2 GND.t169 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X245 VDD.t12 VDD.t9 VDD.t11 VDD.t10 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X246 a_n7336_n129.t23 VN.t17 a_n18640_8567.t9 GND.t10 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=1.7952 ps=6.1 w=5.44 l=5.27
X247 VOUT.t122 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X248 VOUT.t1 CS_BIAS.t107 GND.t168 GND.t167 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X249 GND.t28 GND.t25 GND.t27 GND.t26 sky130_fd_pr__nfet_01v8 ad=3.9168 pd=12.32 as=0 ps=0 w=5.44 l=5.27
X250 GND.t166 CS_BIAS.t108 VOUT.t0 GND.t165 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X251 GND.t162 CS_BIAS.t109 VOUT.t8 GND.t161 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X252 CS_BIAS.t5 CS_BIAS.t4 GND.t160 GND.t159 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X253 VOUT.t7 CS_BIAS.t110 GND.t158 GND.t157 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=2.0088 ps=7.02 w=2.79 l=5.03
X254 VOUT.t123 a_n5326_8245.t0 sky130_fd_pr__cap_mim_m3_1 l=14.74 w=14.15
X255 VOUT.t85 a_n18640_8567.t50 VDD.t78 VDD.t77 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=3.4992 ps=11.16 w=4.86 l=5.24
X256 VDD.t76 a_n18640_8567.t51 VOUT.t84 VDD.t73 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X257 VDD.t75 a_n18640_8567.t52 VOUT.t83 VDD.t73 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X258 DIFFPAIR_BIAS.t3 DIFFPAIR_BIAS.t2 GND.t16 GND.t15 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
X259 GND.t24 GND.t21 GND.t23 GND.t22 sky130_fd_pr__nfet_01v8 ad=2.0088 pd=7.02 as=0 ps=0 w=2.79 l=5.03
X260 a_n7981_10383.t0 a_n7837_10186.t51 VDD.t119 VDD.t118 sky130_fd_pr__pfet_01v8 ad=3.708 pd=11.74 as=1.6995 ps=5.81 w=5.15 l=3.71
X261 VDD.t8 VDD.t6 VDD.t7 VDD.t3 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X262 VDD.t74 a_n18640_8567.t53 VOUT.t82 VDD.t73 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X263 VDD.t72 a_n18640_8567.t54 VOUT.t81 VDD.t70 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X264 VDD.t5 VDD.t2 VDD.t4 VDD.t3 sky130_fd_pr__pfet_01v8 ad=3.4992 pd=11.16 as=0 ps=0 w=4.86 l=5.24
X265 VDD.t71 a_n18640_8567.t55 VOUT.t80 VDD.t70 sky130_fd_pr__pfet_01v8 ad=1.6038 pd=5.52 as=1.6038 ps=5.52 w=4.86 l=5.24
X266 VOUT.t6 CS_BIAS.t111 GND.t156 GND.t155 sky130_fd_pr__nfet_01v8 ad=0.9207 pd=3.45 as=0.9207 ps=3.45 w=2.79 l=5.03
X267 DIFFPAIR_BIAS.t1 DIFFPAIR_BIAS.t0 GND.t269 GND.t268 sky130_fd_pr__nfet_01v8 ad=3.492 pd=11.14 as=3.492 ps=11.14 w=4.85 l=2.45
R0 a_n7837_10186.n17 a_n7837_10186.t18 89.0675
R1 a_n7837_10186.t12 a_n7837_10186.n18 89.0675
R2 a_n7837_10186.n18 a_n7837_10186.t22 87.8118
R3 a_n7837_10186.n17 a_n7837_10186.t26 87.8106
R4 a_n7837_10186.n18 a_n7837_10186.n28 75.1885
R5 a_n7837_10186.n17 a_n7837_10186.n26 75.1885
R6 a_n7837_10186.n15 a_n7837_10186.n25 66.3231
R7 a_n7837_10186.n22 a_n7837_10186.n21 66.323
R8 a_n7837_10186.n22 a_n7837_10186.n19 66.323
R9 a_n7837_10186.n15 a_n7837_10186.n24 64.6191
R10 a_n7837_10186.n15 a_n7837_10186.n23 64.6191
R11 a_n7837_10186.n22 a_n7837_10186.n20 64.619
R12 a_n7837_10186.n15 a_n7837_10186.n22 37.3548
R13 a_n7837_10186.n8 a_n7837_10186.t51 65.9106
R14 a_n7837_10186.n13 a_n7837_10186.t33 67.0001
R15 a_n7837_10186.n13 a_n7837_10186.t45 64.1352
R16 a_n7837_10186.n8 a_n7837_10186.t36 65.9098
R17 a_n7837_10186.n8 a_n7837_10186.t43 65.9106
R18 a_n7837_10186.n10 a_n7837_10186.t49 64.1331
R19 a_n7837_10186.n10 a_n7837_10186.t32 67.0022
R20 a_n7837_10186.n8 a_n7837_10186.t50 65.9098
R21 a_n7837_10186.n8 a_n7837_10186.t34 65.9106
R22 a_n7837_10186.n12 a_n7837_10186.t29 66.6328
R23 a_n7837_10186.n12 a_n7837_10186.t44 64.3247
R24 a_n7837_10186.n8 a_n7837_10186.t31 65.9098
R25 a_n7837_10186.n8 a_n7837_10186.t46 65.9106
R26 a_n7837_10186.n9 a_n7837_10186.t41 64.0787
R27 a_n7837_10186.n9 a_n7837_10186.t30 67.107
R28 a_n7837_10186.n8 a_n7837_10186.t42 65.9098
R29 a_n7837_10186.n2 a_n7837_10186.t40 65.9106
R30 a_n7837_10186.n3 a_n7837_10186.t47 64.0569
R31 a_n7837_10186.n3 a_n7837_10186.t48 67.1572
R32 a_n7837_10186.n2 a_n7837_10186.t35 65.9098
R33 a_n7837_10186.n0 a_n7837_10186.t11 65.9107
R34 a_n7837_10186.n1 a_n7837_10186.t13 64.4727
R35 a_n7837_10186.n14 a_n7837_10186.t21 65.9106
R36 a_n7837_10186.n27 a_n7837_10186.t19 33.4547
R37 a_n7837_10186.n6 a_n7837_10186.t17 65.9106
R38 a_n7837_10186.n7 a_n7837_10186.t15 64.0569
R39 a_n7837_10186.n7 a_n7837_10186.t23 67.1572
R40 a_n7837_10186.n6 a_n7837_10186.t25 65.9098
R41 a_n7837_10186.n4 a_n7837_10186.t37 65.9106
R42 a_n7837_10186.n5 a_n7837_10186.t28 64.0569
R43 a_n7837_10186.n5 a_n7837_10186.t39 67.1572
R44 a_n7837_10186.n4 a_n7837_10186.t38 65.9098
R45 a_n7837_10186.n9 a_n7837_10186.n8 3.6043
R46 a_n7837_10186.n3 a_n7837_10186.n2 3.92555
R47 a_n7837_10186.n27 a_n7837_10186.n14 67.3006
R48 a_n7837_10186.n1 a_n7837_10186.n27 60.9891
R49 a_n7837_10186.n7 a_n7837_10186.n6 3.92555
R50 a_n7837_10186.n5 a_n7837_10186.n4 3.92555
R51 a_n7837_10186.n4 a_n7837_10186.n16 16.8579
R52 a_n7837_10186.n2 a_n7837_10186.n11 16.4336
R53 a_n7837_10186.n1 a_n7837_10186.n0 1.36255
R54 a_n7837_10186.n16 a_n7837_10186.n0 14.8011
R55 a_n7837_10186.n28 a_n7837_10186.t20 12.6238
R56 a_n7837_10186.n28 a_n7837_10186.t14 12.6238
R57 a_n7837_10186.n26 a_n7837_10186.t16 12.6238
R58 a_n7837_10186.n26 a_n7837_10186.t24 12.6238
R59 a_n7837_10186.n11 a_n7837_10186.n6 12.4223
R60 a_n7837_10186.n0 a_n7837_10186.n15 25.6229
R61 a_n7837_10186.n11 a_n7837_10186.n8 11.8295
R62 a_n7837_10186.n11 a_n7837_10186.n17 10.9708
R63 a_n7837_10186.n8 a_n7837_10186.n16 9.02643
R64 a_n7837_10186.n0 a_n7837_10186.n14 8.80874
R65 a_n7837_10186.n18 a_n7837_10186.n16 8.58024
R66 a_n7837_10186.n10 a_n7837_10186.n8 8.10362
R67 a_n7837_10186.n8 a_n7837_10186.n13 7.80594
R68 a_n7837_10186.n0 a_n7837_10186.n2 7.62812
R69 a_n7837_10186.n6 a_n7837_10186.n4 7.62812
R70 a_n7837_10186.n8 a_n7837_10186.n12 7.32566
R71 a_n7837_10186.n25 a_n7837_10186.t9 7.27991
R72 a_n7837_10186.n25 a_n7837_10186.t4 7.27991
R73 a_n7837_10186.n24 a_n7837_10186.t6 7.27991
R74 a_n7837_10186.n24 a_n7837_10186.t7 7.27991
R75 a_n7837_10186.n23 a_n7837_10186.t5 7.27991
R76 a_n7837_10186.n23 a_n7837_10186.t8 7.27991
R77 a_n7837_10186.n21 a_n7837_10186.t27 7.27991
R78 a_n7837_10186.n21 a_n7837_10186.t0 7.27991
R79 a_n7837_10186.n20 a_n7837_10186.t10 7.27991
R80 a_n7837_10186.n20 a_n7837_10186.t3 7.27991
R81 a_n7837_10186.n19 a_n7837_10186.t2 7.27991
R82 a_n7837_10186.n19 a_n7837_10186.t1 7.27991
R83 a_n5326_8245.n1 a_n5326_8245.t3 89.0675
R84 a_n5326_8245.n3 a_n5326_8245.t5 89.0675
R85 a_n5326_8245.n2 a_n5326_8245.t10 89.0664
R86 a_n5326_8245.n1 a_n5326_8245.t4 87.8118
R87 a_n5326_8245.n1 a_n5326_8245.t8 87.8118
R88 a_n5326_8245.n2 a_n5326_8245.t13 87.8118
R89 a_n5326_8245.n3 a_n5326_8245.t9 87.8118
R90 a_n5326_8245.t1 a_n5326_8245.n1 87.8118
R91 a_n5326_8245.n1 a_n5326_8245.n7 75.1885
R92 a_n5326_8245.n1 a_n5326_8245.n6 75.1885
R93 a_n5326_8245.n2 a_n5326_8245.n4 75.1885
R94 a_n5326_8245.n3 a_n5326_8245.n5 75.1885
R95 a_n5326_8245.n0 a_n5326_8245.n3 26.0066
R96 a_n5326_8245.n0 a_n5326_8245.t0 18.3772
R97 a_n5326_8245.n0 a_n5326_8245.n2 13.1351
R98 a_n5326_8245.n7 a_n5326_8245.t12 12.6238
R99 a_n5326_8245.n7 a_n5326_8245.t14 12.6238
R100 a_n5326_8245.n6 a_n5326_8245.t2 12.6238
R101 a_n5326_8245.n6 a_n5326_8245.t11 12.6238
R102 a_n5326_8245.n4 a_n5326_8245.t15 12.6238
R103 a_n5326_8245.n4 a_n5326_8245.t6 12.6238
R104 a_n5326_8245.n5 a_n5326_8245.t7 12.6238
R105 a_n5326_8245.n5 a_n5326_8245.t16 12.6238
R106 a_n5326_8245.n1 a_n5326_8245.n0 9.60179
R107 a_n18640_8567.n15 a_n18640_8567.n85 28.4611
R108 a_n18640_8567.n16 a_n18640_8567.n13 4.23161
R109 a_n18640_8567.n11 a_n18640_8567.n14 4.00359
R110 a_n18640_8567.n9 a_n18640_8567.n86 44.3987
R111 a_n18640_8567.n9 a_n18640_8567.n12 18.831
R112 a_n18640_8567.n6 a_n18640_8567.n10 6.43424
R113 a_n18640_8567.n6 a_n18640_8567.n87 161.3
R114 a_n18640_8567.n7 a_n18640_8567.n8 3.97245
R115 a_n18640_8567.n26 a_n18640_8567.n83 28.4611
R116 a_n18640_8567.n27 a_n18640_8567.n24 4.23161
R117 a_n18640_8567.n22 a_n18640_8567.n25 4.00359
R118 a_n18640_8567.n20 a_n18640_8567.n84 44.3987
R119 a_n18640_8567.n20 a_n18640_8567.n23 18.831
R120 a_n18640_8567.n17 a_n18640_8567.n21 6.43424
R121 a_n18640_8567.n17 a_n18640_8567.n88 161.3
R122 a_n18640_8567.n18 a_n18640_8567.n19 3.97245
R123 a_n18640_8567.n37 a_n18640_8567.n81 28.4611
R124 a_n18640_8567.n38 a_n18640_8567.n35 4.23161
R125 a_n18640_8567.n33 a_n18640_8567.n36 4.00359
R126 a_n18640_8567.n31 a_n18640_8567.n82 44.3987
R127 a_n18640_8567.n31 a_n18640_8567.n34 18.831
R128 a_n18640_8567.n28 a_n18640_8567.n32 6.43424
R129 a_n18640_8567.n28 a_n18640_8567.n89 161.3
R130 a_n18640_8567.n29 a_n18640_8567.n30 3.97245
R131 a_n18640_8567.n78 a_n18640_8567.n47 28.4611
R132 a_n18640_8567.n79 a_n18640_8567.n47 28.4611
R133 a_n18640_8567.n46 a_n18640_8567.n45 4.23161
R134 a_n18640_8567.n44 a_n18640_8567.n43 4.00359
R135 a_n18640_8567.n80 a_n18640_8567.n41 44.3987
R136 a_n18640_8567.n41 a_n18640_8567.n42 18.831
R137 a_n18640_8567.n39 a_n18640_8567.n40 6.43424
R138 a_n18640_8567.n75 a_n18640_8567.n56 28.4611
R139 a_n18640_8567.n76 a_n18640_8567.n56 28.4611
R140 a_n18640_8567.n55 a_n18640_8567.n54 4.23161
R141 a_n18640_8567.n53 a_n18640_8567.n52 4.00359
R142 a_n18640_8567.n77 a_n18640_8567.n50 44.3987
R143 a_n18640_8567.n50 a_n18640_8567.n51 18.831
R144 a_n18640_8567.n48 a_n18640_8567.n49 6.43424
R145 a_n18640_8567.n72 a_n18640_8567.n65 28.4611
R146 a_n18640_8567.n73 a_n18640_8567.n65 28.4611
R147 a_n18640_8567.n64 a_n18640_8567.n63 4.23161
R148 a_n18640_8567.n62 a_n18640_8567.n61 4.00359
R149 a_n18640_8567.n74 a_n18640_8567.n59 44.3987
R150 a_n18640_8567.n59 a_n18640_8567.n60 18.831
R151 a_n18640_8567.n57 a_n18640_8567.n58 6.43424
R152 a_n18640_8567.n92 a_n18640_8567.n90 96.0321
R153 a_n18640_8567.n140 a_n18640_8567.n139 96.0309
R154 a_n18640_8567.n92 a_n18640_8567.n91 94.7763
R155 a_n18640_8567.n141 a_n18640_8567.n140 94.7763
R156 a_n18640_8567.n66 a_n18640_8567.n67 20.4673
R157 a_n18640_8567.n68 a_n18640_8567.n69 20.4673
R158 a_n18640_8567.n70 a_n18640_8567.n71 20.4673
R159 a_n18640_8567.n0 a_n18640_8567.n1 2.07196
R160 a_n18640_8567.n2 a_n18640_8567.n3 2.07196
R161 a_n18640_8567.n4 a_n18640_8567.n5 2.07196
R162 a_n18640_8567.n101 a_n18640_8567.n93 66.3231
R163 a_n18640_8567.n98 a_n18640_8567.n97 66.323
R164 a_n18640_8567.n98 a_n18640_8567.n95 66.323
R165 a_n18640_8567.n100 a_n18640_8567.n99 64.6191
R166 a_n18640_8567.n101 a_n18640_8567.n94 64.6191
R167 a_n18640_8567.n98 a_n18640_8567.n96 64.619
R168 a_n18640_8567.n134 a_n18640_8567.n133 59.0433
R169 a_n18640_8567.n128 a_n18640_8567.n127 59.0433
R170 a_n18640_8567.n123 a_n18640_8567.n122 59.0433
R171 a_n18640_8567.n115 a_n18640_8567.n114 59.0433
R172 a_n18640_8567.n109 a_n18640_8567.n108 59.0433
R173 a_n18640_8567.n104 a_n18640_8567.n103 59.0433
R174 a_n18640_8567.n115 a_n18640_8567.t41 56.3025
R175 a_n18640_8567.n109 a_n18640_8567.t39 56.3025
R176 a_n18640_8567.n104 a_n18640_8567.t40 56.3025
R177 a_n18640_8567.n134 a_n18640_8567.t36 56.3024
R178 a_n18640_8567.n128 a_n18640_8567.t23 56.3024
R179 a_n18640_8567.n123 a_n18640_8567.t22 56.3024
R180 a_n18640_8567.n100 a_n18640_8567.n98 38.3131
R181 a_n18640_8567.n140 a_n18640_8567.n138 33.9236
R182 a_n18640_8567.n1 a_n18640_8567.n78 113.552
R183 a_n18640_8567.n3 a_n18640_8567.n75 113.552
R184 a_n18640_8567.n5 a_n18640_8567.n72 113.552
R185 a_n18640_8567.n8 a_n18640_8567.n67 109.871
R186 a_n18640_8567.n87 a_n18640_8567.n8 73.501
R187 a_n18640_8567.n12 a_n18640_8567.n10 125.445
R188 a_n18640_8567.n12 a_n18640_8567.n131 38.2112
R189 a_n18640_8567.n14 a_n18640_8567.n86 101.389
R190 a_n18640_8567.n132 a_n18640_8567.n14 70.8162
R191 a_n18640_8567.n132 a_n18640_8567.n16 50.5784
R192 a_n18640_8567.n16 a_n18640_8567.n85 117.103
R193 a_n18640_8567.n85 a_n18640_8567.n133 46.6587
R194 a_n18640_8567.n19 a_n18640_8567.n69 109.871
R195 a_n18640_8567.n88 a_n18640_8567.n19 73.501
R196 a_n18640_8567.n23 a_n18640_8567.n21 125.445
R197 a_n18640_8567.n23 a_n18640_8567.n125 38.2112
R198 a_n18640_8567.n25 a_n18640_8567.n84 101.389
R199 a_n18640_8567.n126 a_n18640_8567.n25 70.8162
R200 a_n18640_8567.n126 a_n18640_8567.n27 50.5784
R201 a_n18640_8567.n27 a_n18640_8567.n83 117.103
R202 a_n18640_8567.n83 a_n18640_8567.n127 46.6587
R203 a_n18640_8567.n30 a_n18640_8567.n71 109.871
R204 a_n18640_8567.n89 a_n18640_8567.n30 73.501
R205 a_n18640_8567.n34 a_n18640_8567.n32 125.445
R206 a_n18640_8567.n34 a_n18640_8567.n120 38.2112
R207 a_n18640_8567.n36 a_n18640_8567.n82 101.389
R208 a_n18640_8567.n121 a_n18640_8567.n36 70.8162
R209 a_n18640_8567.n121 a_n18640_8567.n38 50.5784
R210 a_n18640_8567.n38 a_n18640_8567.n81 117.103
R211 a_n18640_8567.n81 a_n18640_8567.n122 46.6587
R212 a_n18640_8567.n40 a_n18640_8567.n42 125.445
R213 a_n18640_8567.n113 a_n18640_8567.n42 38.2112
R214 a_n18640_8567.n44 a_n18640_8567.n80 101.389
R215 a_n18640_8567.n116 a_n18640_8567.n44 70.8162
R216 a_n18640_8567.n46 a_n18640_8567.n116 50.5784
R217 a_n18640_8567.n79 a_n18640_8567.n46 117.103
R218 a_n18640_8567.n117 a_n18640_8567.n79 46.6587
R219 a_n18640_8567.n78 a_n18640_8567.n117 36.8219
R220 a_n18640_8567.n49 a_n18640_8567.n51 125.445
R221 a_n18640_8567.n107 a_n18640_8567.n51 38.2112
R222 a_n18640_8567.n53 a_n18640_8567.n77 101.389
R223 a_n18640_8567.n110 a_n18640_8567.n53 70.8162
R224 a_n18640_8567.n55 a_n18640_8567.n110 50.5784
R225 a_n18640_8567.n76 a_n18640_8567.n55 117.103
R226 a_n18640_8567.n111 a_n18640_8567.n76 46.6587
R227 a_n18640_8567.n75 a_n18640_8567.n111 36.8219
R228 a_n18640_8567.n58 a_n18640_8567.n60 125.445
R229 a_n18640_8567.n102 a_n18640_8567.n60 38.2112
R230 a_n18640_8567.n62 a_n18640_8567.n74 101.389
R231 a_n18640_8567.n105 a_n18640_8567.n62 70.8162
R232 a_n18640_8567.n64 a_n18640_8567.n105 50.5784
R233 a_n18640_8567.n73 a_n18640_8567.n64 117.103
R234 a_n18640_8567.n106 a_n18640_8567.n73 46.6587
R235 a_n18640_8567.n72 a_n18640_8567.n106 36.8219
R236 a_n18640_8567.n67 a_n18640_8567.t48 37.8581
R237 a_n18640_8567.n130 a_n18640_8567.t49 22.3528
R238 a_n18640_8567.n131 a_n18640_8567.t33 22.3528
R239 a_n18640_8567.n132 a_n18640_8567.t34 22.3528
R240 a_n18640_8567.n133 a_n18640_8567.t35 22.3528
R241 a_n18640_8567.n69 a_n18640_8567.t24 37.8581
R242 a_n18640_8567.n124 a_n18640_8567.t37 22.3528
R243 a_n18640_8567.n125 a_n18640_8567.t29 22.3528
R244 a_n18640_8567.n126 a_n18640_8567.t47 22.3528
R245 a_n18640_8567.n127 a_n18640_8567.t55 22.3528
R246 a_n18640_8567.n71 a_n18640_8567.t25 37.8581
R247 a_n18640_8567.n119 a_n18640_8567.t38 22.3528
R248 a_n18640_8567.n120 a_n18640_8567.t31 22.3528
R249 a_n18640_8567.n121 a_n18640_8567.t45 22.3528
R250 a_n18640_8567.n122 a_n18640_8567.t54 22.3528
R251 a_n18640_8567.n114 a_n18640_8567.t28 22.3528
R252 a_n18640_8567.n113 a_n18640_8567.t27 22.3528
R253 a_n18640_8567.n116 a_n18640_8567.t26 22.3528
R254 a_n18640_8567.n117 a_n18640_8567.t53 22.3528
R255 a_n18640_8567.n1 a_n18640_8567.t50 53.1633
R256 a_n18640_8567.n108 a_n18640_8567.t44 22.3528
R257 a_n18640_8567.n107 a_n18640_8567.t30 22.3528
R258 a_n18640_8567.n110 a_n18640_8567.t20 22.3528
R259 a_n18640_8567.n111 a_n18640_8567.t52 22.3528
R260 a_n18640_8567.n3 a_n18640_8567.t43 53.1633
R261 a_n18640_8567.n103 a_n18640_8567.t46 22.3528
R262 a_n18640_8567.n102 a_n18640_8567.t32 22.3528
R263 a_n18640_8567.n105 a_n18640_8567.t21 22.3528
R264 a_n18640_8567.n106 a_n18640_8567.t51 22.3528
R265 a_n18640_8567.n5 a_n18640_8567.t42 53.1633
R266 a_n18640_8567.n86 a_n18640_8567.n131 43.4724
R267 a_n18640_8567.n84 a_n18640_8567.n125 43.4724
R268 a_n18640_8567.n82 a_n18640_8567.n120 43.4724
R269 a_n18640_8567.n80 a_n18640_8567.n113 43.4724
R270 a_n18640_8567.n77 a_n18640_8567.n107 43.4724
R271 a_n18640_8567.n74 a_n18640_8567.n102 43.4724
R272 a_n18640_8567.n138 a_n18640_8567.n92 20.1226
R273 a_n18640_8567.n10 a_n18640_8567.n130 63.5531
R274 a_n18640_8567.n21 a_n18640_8567.n124 63.5531
R275 a_n18640_8567.n32 a_n18640_8567.n119 63.5531
R276 a_n18640_8567.n114 a_n18640_8567.n40 63.5531
R277 a_n18640_8567.n108 a_n18640_8567.n49 63.5531
R278 a_n18640_8567.n103 a_n18640_8567.n58 63.5531
R279 a_n18640_8567.n139 a_n18640_8567.t15 12.6238
R280 a_n18640_8567.n139 a_n18640_8567.t16 12.6238
R281 a_n18640_8567.n91 a_n18640_8567.t12 12.6238
R282 a_n18640_8567.n91 a_n18640_8567.t18 12.6238
R283 a_n18640_8567.n90 a_n18640_8567.t14 12.6238
R284 a_n18640_8567.n90 a_n18640_8567.t13 12.6238
R285 a_n18640_8567.n141 a_n18640_8567.t17 12.6238
R286 a_n18640_8567.t19 a_n18640_8567.n141 12.6238
R287 a_n18640_8567.n137 a_n18640_8567.n101 12.3618
R288 a_n18640_8567.n138 a_n18640_8567.n137 11.4887
R289 a_n18640_8567.n129 a_n18640_8567.n70 8.51486
R290 a_n18640_8567.n112 a_n18640_8567.n4 8.51486
R291 a_n18640_8567.n136 a_n18640_8567.n118 8.1057
R292 a_n18640_8567.n130 a_n18640_8567.n87 7.37805
R293 a_n18640_8567.n124 a_n18640_8567.n88 7.37805
R294 a_n18640_8567.n119 a_n18640_8567.n89 7.37805
R295 a_n18640_8567.n99 a_n18640_8567.t3 7.27991
R296 a_n18640_8567.n99 a_n18640_8567.t5 7.27991
R297 a_n18640_8567.n94 a_n18640_8567.t4 7.27991
R298 a_n18640_8567.n94 a_n18640_8567.t0 7.27991
R299 a_n18640_8567.n93 a_n18640_8567.t9 7.27991
R300 a_n18640_8567.n93 a_n18640_8567.t11 7.27991
R301 a_n18640_8567.n97 a_n18640_8567.t10 7.27991
R302 a_n18640_8567.n97 a_n18640_8567.t2 7.27991
R303 a_n18640_8567.n96 a_n18640_8567.t6 7.27991
R304 a_n18640_8567.n96 a_n18640_8567.t7 7.27991
R305 a_n18640_8567.n95 a_n18640_8567.t8 7.27991
R306 a_n18640_8567.n95 a_n18640_8567.t1 7.27991
R307 a_n18640_8567.n136 a_n18640_8567.n135 6.94637
R308 a_n18640_8567.n135 a_n18640_8567.n66 5.41448
R309 a_n18640_8567.n129 a_n18640_8567.n68 5.41448
R310 a_n18640_8567.n118 a_n18640_8567.n0 5.41448
R311 a_n18640_8567.n112 a_n18640_8567.n2 5.41448
R312 a_n18640_8567.n137 a_n18640_8567.n136 3.4105
R313 a_n18640_8567.n135 a_n18640_8567.n129 3.10088
R314 a_n18640_8567.n118 a_n18640_8567.n112 3.10088
R315 a_n18640_8567.n4 a_n18640_8567.n65 2.35976
R316 a_n18640_8567.n2 a_n18640_8567.n56 2.35976
R317 a_n18640_8567.n0 a_n18640_8567.n47 2.35976
R318 a_n18640_8567.n70 a_n18640_8567.n29 1.98097
R319 a_n18640_8567.n68 a_n18640_8567.n18 1.98097
R320 a_n18640_8567.n66 a_n18640_8567.n7 1.98097
R321 a_n18640_8567.n57 a_n18640_8567.n104 1.71922
R322 a_n18640_8567.n48 a_n18640_8567.n109 1.71922
R323 a_n18640_8567.n39 a_n18640_8567.n115 1.71922
R324 a_n18640_8567.n101 a_n18640_8567.n100 1.70452
R325 a_n18640_8567.n65 a_n18640_8567.n63 1.51565
R326 a_n18640_8567.n63 a_n18640_8567.n61 1.51565
R327 a_n18640_8567.n61 a_n18640_8567.n59 1.51565
R328 a_n18640_8567.n59 a_n18640_8567.n57 1.51565
R329 a_n18640_8567.n56 a_n18640_8567.n54 1.51565
R330 a_n18640_8567.n54 a_n18640_8567.n52 1.51565
R331 a_n18640_8567.n52 a_n18640_8567.n50 1.51565
R332 a_n18640_8567.n50 a_n18640_8567.n48 1.51565
R333 a_n18640_8567.n47 a_n18640_8567.n45 1.51565
R334 a_n18640_8567.n45 a_n18640_8567.n43 1.51565
R335 a_n18640_8567.n43 a_n18640_8567.n41 1.51565
R336 a_n18640_8567.n41 a_n18640_8567.n39 1.51565
R337 a_n18640_8567.n33 a_n18640_8567.n35 1.51565
R338 a_n18640_8567.n31 a_n18640_8567.n33 1.51565
R339 a_n18640_8567.n28 a_n18640_8567.n31 1.51565
R340 a_n18640_8567.n29 a_n18640_8567.n28 1.51565
R341 a_n18640_8567.n22 a_n18640_8567.n24 1.51565
R342 a_n18640_8567.n20 a_n18640_8567.n22 1.51565
R343 a_n18640_8567.n17 a_n18640_8567.n20 1.51565
R344 a_n18640_8567.n18 a_n18640_8567.n17 1.51565
R345 a_n18640_8567.n11 a_n18640_8567.n13 1.51565
R346 a_n18640_8567.n9 a_n18640_8567.n11 1.51565
R347 a_n18640_8567.n6 a_n18640_8567.n9 1.51565
R348 a_n18640_8567.n7 a_n18640_8567.n6 1.51565
R349 a_n18640_8567.n13 a_n18640_8567.n15 1.13686
R350 a_n18640_8567.n24 a_n18640_8567.n26 1.13686
R351 a_n18640_8567.n35 a_n18640_8567.n37 1.13686
R352 a_n18640_8567.n15 a_n18640_8567.n134 0.961639
R353 a_n18640_8567.n26 a_n18640_8567.n128 0.961639
R354 a_n18640_8567.n37 a_n18640_8567.n123 0.961639
R355 VDD.n4221 VDD.n3999 458.05
R356 VDD.n4078 VDD.n4001 458.05
R357 VDD.n3680 VDD.n286 458.05
R358 VDD.n3686 VDD.n288 458.05
R359 VDD.n2196 VDD.n1074 458.05
R360 VDD.n1194 VDD.n1076 458.05
R361 VDD.n1675 VDD.n1497 458.05
R362 VDD.n1671 VDD.n1495 458.05
R363 VDD.n3172 VDD.n621 291.221
R364 VDD.n3522 VDD.n341 291.221
R365 VDD.n3478 VDD.n338 291.221
R366 VDD.n3125 VDD.n3124 291.221
R367 VDD.n2783 VDD.n654 291.221
R368 VDD.n2735 VDD.n2734 291.221
R369 VDD.n2224 VDD.n931 291.221
R370 VDD.n2405 VDD.n933 291.221
R371 VDD.n3457 VDD.n339 291.221
R372 VDD.n3525 VDD.n3524 291.221
R373 VDD.n2893 VDD.n2807 291.221
R374 VDD.n3176 VDD.n625 291.221
R375 VDD.n2720 VDD.n2719 291.221
R376 VDD.n2668 VDD.n641 291.221
R377 VDD.n2398 VDD.n932 291.221
R378 VDD.n2407 VDD.n930 291.221
R379 VDD.n1170 VDD.t54 242.726
R380 VDD.n675 VDD.t31 242.726
R381 VDD.n1047 VDD.t40 242.726
R382 VDD.n657 VDD.t17 242.726
R383 VDD.n2845 VDD.t47 242.726
R384 VDD.n356 VDD.t61 242.726
R385 VDD.n2810 VDD.t51 242.726
R386 VDD.n328 VDD.t57 242.726
R387 VDD.n1500 VDD.t13 232.528
R388 VDD.n1574 VDD.t25 232.528
R389 VDD.n1546 VDD.t28 232.528
R390 VDD.n1195 VDD.t44 232.528
R391 VDD.n1129 VDD.t6 232.528
R392 VDD.n1111 VDD.t2 232.528
R393 VDD.n4080 VDD.t21 232.528
R394 VDD.n4059 VDD.t37 232.528
R395 VDD.n4041 VDD.t34 232.528
R396 VDD.n3592 VDD.t64 232.528
R397 VDD.n3632 VDD.t67 232.528
R398 VDD.n3549 VDD.t9 232.528
R399 VDD.n1500 VDD.t16 197.928
R400 VDD.n1574 VDD.t27 197.928
R401 VDD.n1546 VDD.t30 197.928
R402 VDD.n1195 VDD.t45 197.928
R403 VDD.n1129 VDD.t7 197.928
R404 VDD.n1111 VDD.t4 197.928
R405 VDD.n4080 VDD.t23 197.928
R406 VDD.n4059 VDD.t38 197.928
R407 VDD.n4041 VDD.t35 197.928
R408 VDD.n3592 VDD.t66 197.928
R409 VDD.n3632 VDD.t69 197.928
R410 VDD.n3549 VDD.t12 197.928
R411 VDD.n1074 VDD.n1070 189.749
R412 VDD.n3686 VDD.n291 189.749
R413 VDD.n3680 VDD.n3679 188.06
R414 VDD.n1200 VDD.n1194 188.06
R415 VDD.n2194 VDD.t1 187.629
R416 VDD.n3688 VDD.t0 187.629
R417 VDD.n3459 VDD.n339 185
R418 VDD.n3523 VDD.n339 185
R419 VDD.n3461 VDD.n3460 185
R420 VDD.n3460 VDD.n337 185
R421 VDD.n3462 VDD.n366 185
R422 VDD.n3472 VDD.n366 185
R423 VDD.n3463 VDD.n374 185
R424 VDD.n374 VDD.n364 185
R425 VDD.n3465 VDD.n3464 185
R426 VDD.n3466 VDD.n3465 185
R427 VDD.n3430 VDD.n373 185
R428 VDD.n373 VDD.n370 185
R429 VDD.n3429 VDD.n3428 185
R430 VDD.n3428 VDD.n3427 185
R431 VDD.n376 VDD.n375 185
R432 VDD.n377 VDD.n376 185
R433 VDD.n3420 VDD.n3419 185
R434 VDD.n3421 VDD.n3420 185
R435 VDD.n3418 VDD.n385 185
R436 VDD.n391 VDD.n385 185
R437 VDD.n3417 VDD.n3416 185
R438 VDD.n3416 VDD.n3415 185
R439 VDD.n387 VDD.n386 185
R440 VDD.n388 VDD.n387 185
R441 VDD.n3408 VDD.n3407 185
R442 VDD.n3409 VDD.n3408 185
R443 VDD.n3406 VDD.n398 185
R444 VDD.n398 VDD.n395 185
R445 VDD.n3405 VDD.n3404 185
R446 VDD.n3404 VDD.n3403 185
R447 VDD.n400 VDD.n399 185
R448 VDD.n401 VDD.n400 185
R449 VDD.n3396 VDD.n3395 185
R450 VDD.n3397 VDD.n3396 185
R451 VDD.n3394 VDD.n410 185
R452 VDD.n410 VDD.n407 185
R453 VDD.n3393 VDD.n3392 185
R454 VDD.n3392 VDD.n3391 185
R455 VDD.n412 VDD.n411 185
R456 VDD.n413 VDD.n412 185
R457 VDD.n3384 VDD.n3383 185
R458 VDD.n3385 VDD.n3384 185
R459 VDD.n3382 VDD.n422 185
R460 VDD.n422 VDD.n419 185
R461 VDD.n3381 VDD.n3380 185
R462 VDD.n3380 VDD.n3379 185
R463 VDD.n424 VDD.n423 185
R464 VDD.n425 VDD.n424 185
R465 VDD.n3372 VDD.n3371 185
R466 VDD.n3373 VDD.n3372 185
R467 VDD.n3370 VDD.n433 185
R468 VDD.n3026 VDD.n433 185
R469 VDD.n3369 VDD.n3368 185
R470 VDD.n3368 VDD.n3367 185
R471 VDD.n435 VDD.n434 185
R472 VDD.n436 VDD.n435 185
R473 VDD.n3360 VDD.n3359 185
R474 VDD.n3361 VDD.n3360 185
R475 VDD.n3358 VDD.n445 185
R476 VDD.n445 VDD.n442 185
R477 VDD.n3357 VDD.n3356 185
R478 VDD.n3356 VDD.n3355 185
R479 VDD.n447 VDD.n446 185
R480 VDD.n448 VDD.n447 185
R481 VDD.n3348 VDD.n3347 185
R482 VDD.n3349 VDD.n3348 185
R483 VDD.n3346 VDD.n457 185
R484 VDD.n457 VDD.n454 185
R485 VDD.n3345 VDD.n3344 185
R486 VDD.n3344 VDD.n3343 185
R487 VDD.n459 VDD.n458 185
R488 VDD.n460 VDD.n459 185
R489 VDD.n3336 VDD.n3335 185
R490 VDD.n3337 VDD.n3336 185
R491 VDD.n3334 VDD.n469 185
R492 VDD.n469 VDD.n466 185
R493 VDD.n3333 VDD.n3332 185
R494 VDD.n3332 VDD.n3331 185
R495 VDD.n471 VDD.n470 185
R496 VDD.n480 VDD.n471 185
R497 VDD.n3324 VDD.n3323 185
R498 VDD.n3325 VDD.n3324 185
R499 VDD.n3322 VDD.n481 185
R500 VDD.n481 VDD.n477 185
R501 VDD.n3321 VDD.n3320 185
R502 VDD.n3320 VDD.n3319 185
R503 VDD.n483 VDD.n482 185
R504 VDD.n484 VDD.n483 185
R505 VDD.n3312 VDD.n3311 185
R506 VDD.n3313 VDD.n3312 185
R507 VDD.n3310 VDD.n493 185
R508 VDD.n493 VDD.n490 185
R509 VDD.n3309 VDD.n3308 185
R510 VDD.n3308 VDD.n3307 185
R511 VDD.n495 VDD.n494 185
R512 VDD.n496 VDD.n495 185
R513 VDD.n3300 VDD.n3299 185
R514 VDD.n3301 VDD.n3300 185
R515 VDD.n3298 VDD.n505 185
R516 VDD.n505 VDD.n502 185
R517 VDD.n3297 VDD.n3296 185
R518 VDD.n3296 VDD.n3295 185
R519 VDD.n507 VDD.n506 185
R520 VDD.n516 VDD.n507 185
R521 VDD.n3288 VDD.n3287 185
R522 VDD.n3289 VDD.n3288 185
R523 VDD.n3286 VDD.n517 185
R524 VDD.n517 VDD.n513 185
R525 VDD.n3285 VDD.n3284 185
R526 VDD.n3284 VDD.n3283 185
R527 VDD.n519 VDD.n518 185
R528 VDD.n520 VDD.n519 185
R529 VDD.n3276 VDD.n3275 185
R530 VDD.n3277 VDD.n3276 185
R531 VDD.n3274 VDD.n528 185
R532 VDD.n534 VDD.n528 185
R533 VDD.n3273 VDD.n3272 185
R534 VDD.n3272 VDD.n3271 185
R535 VDD.n530 VDD.n529 185
R536 VDD.n531 VDD.n530 185
R537 VDD.n3264 VDD.n3263 185
R538 VDD.n3265 VDD.n3264 185
R539 VDD.n3262 VDD.n541 185
R540 VDD.n541 VDD.n538 185
R541 VDD.n3261 VDD.n3260 185
R542 VDD.n3260 VDD.n3259 185
R543 VDD.n543 VDD.n542 185
R544 VDD.n544 VDD.n543 185
R545 VDD.n3252 VDD.n3251 185
R546 VDD.n3253 VDD.n3252 185
R547 VDD.n3250 VDD.n553 185
R548 VDD.n553 VDD.n550 185
R549 VDD.n3249 VDD.n3248 185
R550 VDD.n3248 VDD.n3247 185
R551 VDD.n555 VDD.n554 185
R552 VDD.n556 VDD.n555 185
R553 VDD.n3240 VDD.n3239 185
R554 VDD.n3241 VDD.n3240 185
R555 VDD.n3238 VDD.n565 185
R556 VDD.n565 VDD.n562 185
R557 VDD.n3237 VDD.n3236 185
R558 VDD.n3236 VDD.n3235 185
R559 VDD.n567 VDD.n566 185
R560 VDD.n568 VDD.n567 185
R561 VDD.n3228 VDD.n3227 185
R562 VDD.n3229 VDD.n3228 185
R563 VDD.n3226 VDD.n577 185
R564 VDD.n577 VDD.n574 185
R565 VDD.n3225 VDD.n3224 185
R566 VDD.n3224 VDD.n3223 185
R567 VDD.n579 VDD.n578 185
R568 VDD.n580 VDD.n579 185
R569 VDD.n3216 VDD.n3215 185
R570 VDD.n3217 VDD.n3216 185
R571 VDD.n3214 VDD.n589 185
R572 VDD.n589 VDD.n586 185
R573 VDD.n3213 VDD.n3212 185
R574 VDD.n3212 VDD.n3211 185
R575 VDD.n591 VDD.n590 185
R576 VDD.n592 VDD.n591 185
R577 VDD.n3204 VDD.n3203 185
R578 VDD.n3205 VDD.n3204 185
R579 VDD.n3202 VDD.n600 185
R580 VDD.n605 VDD.n600 185
R581 VDD.n3201 VDD.n3200 185
R582 VDD.n3200 VDD.n3199 185
R583 VDD.n602 VDD.n601 185
R584 VDD.n612 VDD.n602 185
R585 VDD.n3192 VDD.n3191 185
R586 VDD.n3193 VDD.n3192 185
R587 VDD.n3190 VDD.n613 185
R588 VDD.n613 VDD.n609 185
R589 VDD.n3189 VDD.n3188 185
R590 VDD.n3188 VDD.n3187 185
R591 VDD.n615 VDD.n614 185
R592 VDD.n616 VDD.n615 185
R593 VDD.n3180 VDD.n3179 185
R594 VDD.n3181 VDD.n3180 185
R595 VDD.n3178 VDD.n625 185
R596 VDD.n625 VDD.n622 185
R597 VDD.n3177 VDD.n3176 185
R598 VDD.n627 VDD.n626 185
R599 VDD.n2848 VDD.n2847 185
R600 VDD.n2850 VDD.n2849 185
R601 VDD.n2852 VDD.n2851 185
R602 VDD.n2854 VDD.n2853 185
R603 VDD.n2856 VDD.n2855 185
R604 VDD.n2858 VDD.n2857 185
R605 VDD.n2860 VDD.n2859 185
R606 VDD.n2862 VDD.n2861 185
R607 VDD.n2864 VDD.n2863 185
R608 VDD.n2866 VDD.n2865 185
R609 VDD.n2868 VDD.n2867 185
R610 VDD.n2870 VDD.n2869 185
R611 VDD.n2872 VDD.n2871 185
R612 VDD.n2874 VDD.n2873 185
R613 VDD.n2876 VDD.n2875 185
R614 VDD.n2878 VDD.n2877 185
R615 VDD.n2880 VDD.n2879 185
R616 VDD.n2882 VDD.n2881 185
R617 VDD.n2884 VDD.n2883 185
R618 VDD.n2887 VDD.n2886 185
R619 VDD.n2889 VDD.n2888 185
R620 VDD.n2891 VDD.n2890 185
R621 VDD.n2892 VDD.n2807 185
R622 VDD.n3174 VDD.n2807 185
R623 VDD.n3526 VDD.n3525 185
R624 VDD.n3527 VDD.n333 185
R625 VDD.n3529 VDD.n3528 185
R626 VDD.n3531 VDD.n332 185
R627 VDD.n3533 VDD.n3532 185
R628 VDD.n3534 VDD.n327 185
R629 VDD.n3536 VDD.n3535 185
R630 VDD.n3538 VDD.n325 185
R631 VDD.n3540 VDD.n3539 185
R632 VDD.n3541 VDD.n324 185
R633 VDD.n3543 VDD.n3542 185
R634 VDD.n3545 VDD.n321 185
R635 VDD.n3547 VDD.n3546 185
R636 VDD.n3438 VDD.n320 185
R637 VDD.n3440 VDD.n3439 185
R638 VDD.n3442 VDD.n3436 185
R639 VDD.n3444 VDD.n3443 185
R640 VDD.n3445 VDD.n3435 185
R641 VDD.n3447 VDD.n3446 185
R642 VDD.n3449 VDD.n3433 185
R643 VDD.n3451 VDD.n3450 185
R644 VDD.n3452 VDD.n3432 185
R645 VDD.n3454 VDD.n3453 185
R646 VDD.n3456 VDD.n3431 185
R647 VDD.n3458 VDD.n3457 185
R648 VDD.n3457 VDD.n323 185
R649 VDD.n3524 VDD.n334 185
R650 VDD.n3524 VDD.n3523 185
R651 VDD.n2989 VDD.n336 185
R652 VDD.n337 VDD.n336 185
R653 VDD.n2990 VDD.n365 185
R654 VDD.n3472 VDD.n365 185
R655 VDD.n2992 VDD.n2991 185
R656 VDD.n2991 VDD.n364 185
R657 VDD.n2993 VDD.n372 185
R658 VDD.n3466 VDD.n372 185
R659 VDD.n2995 VDD.n2994 185
R660 VDD.n2994 VDD.n370 185
R661 VDD.n2996 VDD.n379 185
R662 VDD.n3427 VDD.n379 185
R663 VDD.n2998 VDD.n2997 185
R664 VDD.n2997 VDD.n377 185
R665 VDD.n2999 VDD.n384 185
R666 VDD.n3421 VDD.n384 185
R667 VDD.n3001 VDD.n3000 185
R668 VDD.n3000 VDD.n391 185
R669 VDD.n3002 VDD.n390 185
R670 VDD.n3415 VDD.n390 185
R671 VDD.n3004 VDD.n3003 185
R672 VDD.n3003 VDD.n388 185
R673 VDD.n3005 VDD.n397 185
R674 VDD.n3409 VDD.n397 185
R675 VDD.n3007 VDD.n3006 185
R676 VDD.n3006 VDD.n395 185
R677 VDD.n3008 VDD.n403 185
R678 VDD.n3403 VDD.n403 185
R679 VDD.n3010 VDD.n3009 185
R680 VDD.n3009 VDD.n401 185
R681 VDD.n3011 VDD.n409 185
R682 VDD.n3397 VDD.n409 185
R683 VDD.n3013 VDD.n3012 185
R684 VDD.n3012 VDD.n407 185
R685 VDD.n3014 VDD.n415 185
R686 VDD.n3391 VDD.n415 185
R687 VDD.n3016 VDD.n3015 185
R688 VDD.n3015 VDD.n413 185
R689 VDD.n3017 VDD.n421 185
R690 VDD.n3385 VDD.n421 185
R691 VDD.n3019 VDD.n3018 185
R692 VDD.n3018 VDD.n419 185
R693 VDD.n3020 VDD.n427 185
R694 VDD.n3379 VDD.n427 185
R695 VDD.n3022 VDD.n3021 185
R696 VDD.n3021 VDD.n425 185
R697 VDD.n3023 VDD.n432 185
R698 VDD.n3373 VDD.n432 185
R699 VDD.n3025 VDD.n3024 185
R700 VDD.n3026 VDD.n3025 185
R701 VDD.n2988 VDD.n438 185
R702 VDD.n3367 VDD.n438 185
R703 VDD.n2987 VDD.n2986 185
R704 VDD.n2986 VDD.n436 185
R705 VDD.n2985 VDD.n444 185
R706 VDD.n3361 VDD.n444 185
R707 VDD.n2984 VDD.n2983 185
R708 VDD.n2983 VDD.n442 185
R709 VDD.n2982 VDD.n450 185
R710 VDD.n3355 VDD.n450 185
R711 VDD.n2981 VDD.n2980 185
R712 VDD.n2980 VDD.n448 185
R713 VDD.n2979 VDD.n456 185
R714 VDD.n3349 VDD.n456 185
R715 VDD.n2978 VDD.n2977 185
R716 VDD.n2977 VDD.n454 185
R717 VDD.n2976 VDD.n462 185
R718 VDD.n3343 VDD.n462 185
R719 VDD.n2975 VDD.n2974 185
R720 VDD.n2974 VDD.n460 185
R721 VDD.n2973 VDD.n468 185
R722 VDD.n3337 VDD.n468 185
R723 VDD.n2972 VDD.n2971 185
R724 VDD.n2971 VDD.n466 185
R725 VDD.n2970 VDD.n473 185
R726 VDD.n3331 VDD.n473 185
R727 VDD.n2969 VDD.n2968 185
R728 VDD.n2968 VDD.n480 185
R729 VDD.n2967 VDD.n479 185
R730 VDD.n3325 VDD.n479 185
R731 VDD.n2966 VDD.n2965 185
R732 VDD.n2965 VDD.n477 185
R733 VDD.n2964 VDD.n486 185
R734 VDD.n3319 VDD.n486 185
R735 VDD.n2963 VDD.n2962 185
R736 VDD.n2962 VDD.n484 185
R737 VDD.n2961 VDD.n492 185
R738 VDD.n3313 VDD.n492 185
R739 VDD.n2960 VDD.n2959 185
R740 VDD.n2959 VDD.n490 185
R741 VDD.n2958 VDD.n498 185
R742 VDD.n3307 VDD.n498 185
R743 VDD.n2957 VDD.n2956 185
R744 VDD.n2956 VDD.n496 185
R745 VDD.n2955 VDD.n504 185
R746 VDD.n3301 VDD.n504 185
R747 VDD.n2954 VDD.n2953 185
R748 VDD.n2953 VDD.n502 185
R749 VDD.n2952 VDD.n509 185
R750 VDD.n3295 VDD.n509 185
R751 VDD.n2951 VDD.n2950 185
R752 VDD.n2950 VDD.n516 185
R753 VDD.n2949 VDD.n515 185
R754 VDD.n3289 VDD.n515 185
R755 VDD.n2948 VDD.n2947 185
R756 VDD.n2947 VDD.n513 185
R757 VDD.n2946 VDD.n522 185
R758 VDD.n3283 VDD.n522 185
R759 VDD.n2945 VDD.n2944 185
R760 VDD.n2944 VDD.n520 185
R761 VDD.n2943 VDD.n527 185
R762 VDD.n3277 VDD.n527 185
R763 VDD.n2942 VDD.n2941 185
R764 VDD.n2941 VDD.n534 185
R765 VDD.n2940 VDD.n533 185
R766 VDD.n3271 VDD.n533 185
R767 VDD.n2939 VDD.n2938 185
R768 VDD.n2938 VDD.n531 185
R769 VDD.n2937 VDD.n540 185
R770 VDD.n3265 VDD.n540 185
R771 VDD.n2936 VDD.n2935 185
R772 VDD.n2935 VDD.n538 185
R773 VDD.n2934 VDD.n546 185
R774 VDD.n3259 VDD.n546 185
R775 VDD.n2933 VDD.n2932 185
R776 VDD.n2932 VDD.n544 185
R777 VDD.n2931 VDD.n552 185
R778 VDD.n3253 VDD.n552 185
R779 VDD.n2930 VDD.n2929 185
R780 VDD.n2929 VDD.n550 185
R781 VDD.n2928 VDD.n558 185
R782 VDD.n3247 VDD.n558 185
R783 VDD.n2927 VDD.n2926 185
R784 VDD.n2926 VDD.n556 185
R785 VDD.n2925 VDD.n564 185
R786 VDD.n3241 VDD.n564 185
R787 VDD.n2924 VDD.n2923 185
R788 VDD.n2923 VDD.n562 185
R789 VDD.n2922 VDD.n570 185
R790 VDD.n3235 VDD.n570 185
R791 VDD.n2921 VDD.n2920 185
R792 VDD.n2920 VDD.n568 185
R793 VDD.n2919 VDD.n576 185
R794 VDD.n3229 VDD.n576 185
R795 VDD.n2918 VDD.n2917 185
R796 VDD.n2917 VDD.n574 185
R797 VDD.n2916 VDD.n582 185
R798 VDD.n3223 VDD.n582 185
R799 VDD.n2915 VDD.n2914 185
R800 VDD.n2914 VDD.n580 185
R801 VDD.n2913 VDD.n588 185
R802 VDD.n3217 VDD.n588 185
R803 VDD.n2912 VDD.n2911 185
R804 VDD.n2911 VDD.n586 185
R805 VDD.n2910 VDD.n594 185
R806 VDD.n3211 VDD.n594 185
R807 VDD.n2909 VDD.n2908 185
R808 VDD.n2908 VDD.n592 185
R809 VDD.n2907 VDD.n599 185
R810 VDD.n3205 VDD.n599 185
R811 VDD.n2906 VDD.n2905 185
R812 VDD.n2905 VDD.n605 185
R813 VDD.n2904 VDD.n604 185
R814 VDD.n3199 VDD.n604 185
R815 VDD.n2903 VDD.n2902 185
R816 VDD.n2902 VDD.n612 185
R817 VDD.n2901 VDD.n611 185
R818 VDD.n3193 VDD.n611 185
R819 VDD.n2900 VDD.n2899 185
R820 VDD.n2899 VDD.n609 185
R821 VDD.n2898 VDD.n618 185
R822 VDD.n3187 VDD.n618 185
R823 VDD.n2897 VDD.n2896 185
R824 VDD.n2896 VDD.n616 185
R825 VDD.n2895 VDD.n624 185
R826 VDD.n3181 VDD.n624 185
R827 VDD.n2894 VDD.n2893 185
R828 VDD.n2893 VDD.n622 185
R829 VDD.n2197 VDD.n2196 185
R830 VDD.n2196 VDD.n2195 185
R831 VDD.n1073 VDD.n1072 185
R832 VDD.n1075 VDD.n1073 185
R833 VDD.n2095 VDD.n2094 185
R834 VDD.n2096 VDD.n2095 185
R835 VDD.n1206 VDD.n1205 185
R836 VDD.n1205 VDD.n1204 185
R837 VDD.n2090 VDD.n2089 185
R838 VDD.n2089 VDD.n2088 185
R839 VDD.n1209 VDD.n1208 185
R840 VDD.n1210 VDD.n1209 185
R841 VDD.n2077 VDD.n2076 185
R842 VDD.n2078 VDD.n2077 185
R843 VDD.n1218 VDD.n1217 185
R844 VDD.n2069 VDD.n1217 185
R845 VDD.n2072 VDD.n2071 185
R846 VDD.n2071 VDD.n2070 185
R847 VDD.n1221 VDD.n1220 185
R848 VDD.n1222 VDD.n1221 185
R849 VDD.n2060 VDD.n2059 185
R850 VDD.n2061 VDD.n2060 185
R851 VDD.n1230 VDD.n1229 185
R852 VDD.n1229 VDD.n1228 185
R853 VDD.n2055 VDD.n2054 185
R854 VDD.n2054 VDD.n2053 185
R855 VDD.n1233 VDD.n1232 185
R856 VDD.n1234 VDD.n1233 185
R857 VDD.n2044 VDD.n2043 185
R858 VDD.n2045 VDD.n2044 185
R859 VDD.n1242 VDD.n1241 185
R860 VDD.n1241 VDD.n1240 185
R861 VDD.n2039 VDD.n2038 185
R862 VDD.n2038 VDD.n2037 185
R863 VDD.n1245 VDD.n1244 185
R864 VDD.n1246 VDD.n1245 185
R865 VDD.n2028 VDD.n2027 185
R866 VDD.n2029 VDD.n2028 185
R867 VDD.n1254 VDD.n1253 185
R868 VDD.n1253 VDD.n1252 185
R869 VDD.n2023 VDD.n2022 185
R870 VDD.n2022 VDD.n2021 185
R871 VDD.n1257 VDD.n1256 185
R872 VDD.t77 VDD.n1257 185
R873 VDD.n2012 VDD.n2011 185
R874 VDD.n2013 VDD.n2012 185
R875 VDD.n1265 VDD.n1264 185
R876 VDD.n1264 VDD.n1263 185
R877 VDD.n2007 VDD.n2006 185
R878 VDD.n2006 VDD.n2005 185
R879 VDD.n1268 VDD.n1267 185
R880 VDD.n1269 VDD.n1268 185
R881 VDD.n1996 VDD.n1995 185
R882 VDD.n1997 VDD.n1996 185
R883 VDD.n1277 VDD.n1276 185
R884 VDD.n1276 VDD.n1275 185
R885 VDD.n1991 VDD.n1990 185
R886 VDD.n1990 VDD.n1989 185
R887 VDD.n1280 VDD.n1279 185
R888 VDD.n1281 VDD.n1280 185
R889 VDD.n1980 VDD.n1979 185
R890 VDD.n1981 VDD.n1980 185
R891 VDD.n1289 VDD.n1288 185
R892 VDD.n1288 VDD.n1287 185
R893 VDD.n1975 VDD.n1974 185
R894 VDD.n1974 VDD.n1973 185
R895 VDD.n1292 VDD.n1291 185
R896 VDD.n1299 VDD.n1292 185
R897 VDD.n1964 VDD.n1963 185
R898 VDD.n1965 VDD.n1964 185
R899 VDD.n1301 VDD.n1300 185
R900 VDD.n1300 VDD.n1298 185
R901 VDD.n1959 VDD.n1958 185
R902 VDD.n1958 VDD.n1957 185
R903 VDD.n1304 VDD.n1303 185
R904 VDD.n1305 VDD.n1304 185
R905 VDD.n1948 VDD.n1947 185
R906 VDD.n1949 VDD.n1948 185
R907 VDD.n1313 VDD.n1312 185
R908 VDD.n1312 VDD.n1311 185
R909 VDD.n1943 VDD.n1942 185
R910 VDD.n1942 VDD.n1941 185
R911 VDD.n1316 VDD.n1315 185
R912 VDD.n1317 VDD.n1316 185
R913 VDD.n1932 VDD.n1931 185
R914 VDD.n1933 VDD.n1932 185
R915 VDD.n1325 VDD.n1324 185
R916 VDD.n1324 VDD.n1323 185
R917 VDD.n1927 VDD.n1926 185
R918 VDD.n1926 VDD.n1925 185
R919 VDD.n1328 VDD.n1327 185
R920 VDD.n1335 VDD.n1328 185
R921 VDD.n1916 VDD.n1915 185
R922 VDD.n1917 VDD.n1916 185
R923 VDD.n1337 VDD.n1336 185
R924 VDD.n1336 VDD.n1334 185
R925 VDD.n1911 VDD.n1910 185
R926 VDD.n1910 VDD.n1909 185
R927 VDD.n1340 VDD.n1339 185
R928 VDD.n1341 VDD.n1340 185
R929 VDD.n1900 VDD.n1899 185
R930 VDD.n1901 VDD.n1900 185
R931 VDD.n1349 VDD.n1348 185
R932 VDD.n1348 VDD.n1347 185
R933 VDD.n1876 VDD.n1875 185
R934 VDD.n1875 VDD.n1874 185
R935 VDD.n1352 VDD.n1351 185
R936 VDD.n1353 VDD.n1352 185
R937 VDD.n1865 VDD.n1864 185
R938 VDD.n1866 VDD.n1865 185
R939 VDD.n1361 VDD.n1360 185
R940 VDD.n1360 VDD.n1359 185
R941 VDD.n1860 VDD.n1859 185
R942 VDD.n1859 VDD.n1858 185
R943 VDD.n1364 VDD.n1363 185
R944 VDD.n1371 VDD.n1364 185
R945 VDD.n1849 VDD.n1848 185
R946 VDD.n1850 VDD.n1849 185
R947 VDD.n1373 VDD.n1372 185
R948 VDD.n1372 VDD.n1370 185
R949 VDD.n1844 VDD.n1843 185
R950 VDD.n1843 VDD.n1842 185
R951 VDD.n1376 VDD.n1375 185
R952 VDD.n1377 VDD.n1376 185
R953 VDD.n1833 VDD.n1832 185
R954 VDD.n1834 VDD.n1833 185
R955 VDD.n1385 VDD.n1384 185
R956 VDD.n1384 VDD.n1383 185
R957 VDD.n1828 VDD.n1827 185
R958 VDD.n1827 VDD.n1826 185
R959 VDD.n1388 VDD.n1387 185
R960 VDD.n1389 VDD.n1388 185
R961 VDD.n1817 VDD.n1816 185
R962 VDD.n1818 VDD.n1817 185
R963 VDD.n1397 VDD.n1396 185
R964 VDD.n1396 VDD.n1395 185
R965 VDD.n1812 VDD.n1811 185
R966 VDD.n1811 VDD.n1810 185
R967 VDD.n1400 VDD.n1399 185
R968 VDD.n1407 VDD.n1400 185
R969 VDD.n1801 VDD.n1800 185
R970 VDD.n1802 VDD.n1801 185
R971 VDD.n1409 VDD.n1408 185
R972 VDD.n1408 VDD.n1406 185
R973 VDD.n1796 VDD.n1795 185
R974 VDD.n1795 VDD.n1794 185
R975 VDD.n1412 VDD.n1411 185
R976 VDD.n1413 VDD.n1412 185
R977 VDD.n1785 VDD.n1784 185
R978 VDD.n1786 VDD.n1785 185
R979 VDD.n1421 VDD.n1420 185
R980 VDD.n1420 VDD.n1419 185
R981 VDD.n1780 VDD.n1779 185
R982 VDD.n1779 VDD.n1778 185
R983 VDD.n1424 VDD.n1423 185
R984 VDD.n1425 VDD.n1424 185
R985 VDD.n1769 VDD.n1768 185
R986 VDD.n1770 VDD.n1769 185
R987 VDD.n1433 VDD.n1432 185
R988 VDD.n1432 VDD.n1431 185
R989 VDD.n1764 VDD.n1763 185
R990 VDD.n1763 VDD.t91 185
R991 VDD.n1436 VDD.n1435 185
R992 VDD.n1437 VDD.n1436 185
R993 VDD.n1754 VDD.n1753 185
R994 VDD.n1755 VDD.n1754 185
R995 VDD.n1445 VDD.n1444 185
R996 VDD.n1444 VDD.n1443 185
R997 VDD.n1749 VDD.n1748 185
R998 VDD.n1748 VDD.n1747 185
R999 VDD.n1448 VDD.n1447 185
R1000 VDD.n1449 VDD.n1448 185
R1001 VDD.n1738 VDD.n1737 185
R1002 VDD.n1739 VDD.n1738 185
R1003 VDD.n1457 VDD.n1456 185
R1004 VDD.n1456 VDD.n1455 185
R1005 VDD.n1733 VDD.n1732 185
R1006 VDD.n1732 VDD.n1731 185
R1007 VDD.n1460 VDD.n1459 185
R1008 VDD.n1461 VDD.n1460 185
R1009 VDD.n1722 VDD.n1721 185
R1010 VDD.n1723 VDD.n1722 185
R1011 VDD.n1469 VDD.n1468 185
R1012 VDD.n1468 VDD.n1467 185
R1013 VDD.n1717 VDD.n1716 185
R1014 VDD.n1716 VDD.n1715 185
R1015 VDD.n1472 VDD.n1471 185
R1016 VDD.n1473 VDD.n1472 185
R1017 VDD.n1706 VDD.n1705 185
R1018 VDD.n1707 VDD.n1706 185
R1019 VDD.n1480 VDD.n1479 185
R1020 VDD.n1698 VDD.n1479 185
R1021 VDD.n1701 VDD.n1700 185
R1022 VDD.n1700 VDD.n1699 185
R1023 VDD.n1483 VDD.n1482 185
R1024 VDD.n1484 VDD.n1483 185
R1025 VDD.n1689 VDD.n1688 185
R1026 VDD.n1690 VDD.n1689 185
R1027 VDD.n1492 VDD.n1491 185
R1028 VDD.n1491 VDD.n1490 185
R1029 VDD.n1684 VDD.n1683 185
R1030 VDD.n1683 VDD.n1682 185
R1031 VDD.n1495 VDD.n1494 185
R1032 VDD.n1496 VDD.n1495 185
R1033 VDD.n1671 VDD.n1670 185
R1034 VDD.n1669 VDD.n1527 185
R1035 VDD.n1529 VDD.n1526 185
R1036 VDD.n1673 VDD.n1526 185
R1037 VDD.n1665 VDD.n1531 185
R1038 VDD.n1664 VDD.n1532 185
R1039 VDD.n1663 VDD.n1533 185
R1040 VDD.n1536 VDD.n1534 185
R1041 VDD.n1659 VDD.n1537 185
R1042 VDD.n1658 VDD.n1538 185
R1043 VDD.n1657 VDD.n1539 185
R1044 VDD.n1542 VDD.n1540 185
R1045 VDD.n1653 VDD.n1543 185
R1046 VDD.n1652 VDD.n1544 185
R1047 VDD.n1651 VDD.n1545 185
R1048 VDD.n1550 VDD.n1548 185
R1049 VDD.n1647 VDD.n1551 185
R1050 VDD.n1646 VDD.n1552 185
R1051 VDD.n1645 VDD.n1553 185
R1052 VDD.n1556 VDD.n1554 185
R1053 VDD.n1641 VDD.n1557 185
R1054 VDD.n1640 VDD.n1558 185
R1055 VDD.n1639 VDD.n1559 185
R1056 VDD.n1562 VDD.n1560 185
R1057 VDD.n1635 VDD.n1563 185
R1058 VDD.n1634 VDD.n1564 185
R1059 VDD.n1633 VDD.n1565 185
R1060 VDD.n1568 VDD.n1566 185
R1061 VDD.n1629 VDD.n1569 185
R1062 VDD.n1628 VDD.n1570 185
R1063 VDD.n1627 VDD.n1571 185
R1064 VDD.n1577 VDD.n1572 185
R1065 VDD.n1623 VDD.n1578 185
R1066 VDD.n1622 VDD.n1579 185
R1067 VDD.n1621 VDD.n1580 185
R1068 VDD.n1583 VDD.n1581 185
R1069 VDD.n1617 VDD.n1584 185
R1070 VDD.n1616 VDD.n1585 185
R1071 VDD.n1615 VDD.n1586 185
R1072 VDD.n1589 VDD.n1587 185
R1073 VDD.n1611 VDD.n1590 185
R1074 VDD.n1610 VDD.n1591 185
R1075 VDD.n1609 VDD.n1592 185
R1076 VDD.n1595 VDD.n1593 185
R1077 VDD.n1605 VDD.n1596 185
R1078 VDD.n1604 VDD.n1597 185
R1079 VDD.n1603 VDD.n1598 185
R1080 VDD.n1600 VDD.n1599 185
R1081 VDD.n1503 VDD.n1502 185
R1082 VDD.n1676 VDD.n1675 185
R1083 VDD.n1199 VDD.n1198 185
R1084 VDD.n1197 VDD.n1146 185
R1085 VDD.n2105 VDD.n2104 185
R1086 VDD.n2107 VDD.n2106 185
R1087 VDD.n2109 VDD.n2108 185
R1088 VDD.n2111 VDD.n2110 185
R1089 VDD.n2113 VDD.n2112 185
R1090 VDD.n2115 VDD.n2114 185
R1091 VDD.n2117 VDD.n2116 185
R1092 VDD.n2119 VDD.n2118 185
R1093 VDD.n2121 VDD.n2120 185
R1094 VDD.n2123 VDD.n2122 185
R1095 VDD.n2125 VDD.n2124 185
R1096 VDD.n2127 VDD.n2126 185
R1097 VDD.n2129 VDD.n2128 185
R1098 VDD.n2131 VDD.n2130 185
R1099 VDD.n2133 VDD.n2132 185
R1100 VDD.n2135 VDD.n2134 185
R1101 VDD.n2137 VDD.n2136 185
R1102 VDD.n2139 VDD.n2138 185
R1103 VDD.n2141 VDD.n2140 185
R1104 VDD.n2143 VDD.n2142 185
R1105 VDD.n2145 VDD.n2144 185
R1106 VDD.n2147 VDD.n2146 185
R1107 VDD.n2149 VDD.n2148 185
R1108 VDD.n2151 VDD.n2150 185
R1109 VDD.n2153 VDD.n2152 185
R1110 VDD.n2155 VDD.n2154 185
R1111 VDD.n2157 VDD.n2156 185
R1112 VDD.n2159 VDD.n2158 185
R1113 VDD.n2161 VDD.n2160 185
R1114 VDD.n2163 VDD.n2162 185
R1115 VDD.n1113 VDD.n1110 185
R1116 VDD.n2167 VDD.n1114 185
R1117 VDD.n2169 VDD.n2168 185
R1118 VDD.n2171 VDD.n2170 185
R1119 VDD.n2173 VDD.n2172 185
R1120 VDD.n2175 VDD.n2174 185
R1121 VDD.n2177 VDD.n2176 185
R1122 VDD.n2179 VDD.n2178 185
R1123 VDD.n2181 VDD.n2180 185
R1124 VDD.n2183 VDD.n2182 185
R1125 VDD.n2185 VDD.n2184 185
R1126 VDD.n2187 VDD.n2186 185
R1127 VDD.n2189 VDD.n2188 185
R1128 VDD.n2192 VDD.n2191 185
R1129 VDD.n2190 VDD.n1100 185
R1130 VDD.n2194 VDD.n1074 185
R1131 VDD.n2100 VDD.n1076 185
R1132 VDD.n2195 VDD.n1076 185
R1133 VDD.n2099 VDD.n2098 185
R1134 VDD.n2098 VDD.n1075 185
R1135 VDD.n2097 VDD.n1202 185
R1136 VDD.n2097 VDD.n2096 185
R1137 VDD.n1213 VDD.n1203 185
R1138 VDD.n1204 VDD.n1203 185
R1139 VDD.n2087 VDD.n2086 185
R1140 VDD.n2088 VDD.n2087 185
R1141 VDD.n1212 VDD.n1211 185
R1142 VDD.n1211 VDD.n1210 185
R1143 VDD.n2080 VDD.n2079 185
R1144 VDD.n2079 VDD.n2078 185
R1145 VDD.n1216 VDD.n1215 185
R1146 VDD.n2069 VDD.n1216 185
R1147 VDD.n2068 VDD.n2067 185
R1148 VDD.n2070 VDD.n2068 185
R1149 VDD.n1224 VDD.n1223 185
R1150 VDD.n1223 VDD.n1222 185
R1151 VDD.n2063 VDD.n2062 185
R1152 VDD.n2062 VDD.n2061 185
R1153 VDD.n1227 VDD.n1226 185
R1154 VDD.n1228 VDD.n1227 185
R1155 VDD.n2052 VDD.n2051 185
R1156 VDD.n2053 VDD.n2052 185
R1157 VDD.n1236 VDD.n1235 185
R1158 VDD.n1235 VDD.n1234 185
R1159 VDD.n2047 VDD.n2046 185
R1160 VDD.n2046 VDD.n2045 185
R1161 VDD.n1239 VDD.n1238 185
R1162 VDD.n1240 VDD.n1239 185
R1163 VDD.n2036 VDD.n2035 185
R1164 VDD.n2037 VDD.n2036 185
R1165 VDD.n1248 VDD.n1247 185
R1166 VDD.n1247 VDD.n1246 185
R1167 VDD.n2031 VDD.n2030 185
R1168 VDD.n2030 VDD.n2029 185
R1169 VDD.n1251 VDD.n1250 185
R1170 VDD.n1252 VDD.n1251 185
R1171 VDD.n2020 VDD.n2019 185
R1172 VDD.n2021 VDD.n2020 185
R1173 VDD.n1259 VDD.n1258 185
R1174 VDD.n1258 VDD.t77 185
R1175 VDD.n2015 VDD.n2014 185
R1176 VDD.n2014 VDD.n2013 185
R1177 VDD.n1262 VDD.n1261 185
R1178 VDD.n1263 VDD.n1262 185
R1179 VDD.n2004 VDD.n2003 185
R1180 VDD.n2005 VDD.n2004 185
R1181 VDD.n1271 VDD.n1270 185
R1182 VDD.n1270 VDD.n1269 185
R1183 VDD.n1999 VDD.n1998 185
R1184 VDD.n1998 VDD.n1997 185
R1185 VDD.n1274 VDD.n1273 185
R1186 VDD.n1275 VDD.n1274 185
R1187 VDD.n1988 VDD.n1987 185
R1188 VDD.n1989 VDD.n1988 185
R1189 VDD.n1283 VDD.n1282 185
R1190 VDD.n1282 VDD.n1281 185
R1191 VDD.n1983 VDD.n1982 185
R1192 VDD.n1982 VDD.n1981 185
R1193 VDD.n1286 VDD.n1285 185
R1194 VDD.n1287 VDD.n1286 185
R1195 VDD.n1972 VDD.n1971 185
R1196 VDD.n1973 VDD.n1972 185
R1197 VDD.n1294 VDD.n1293 185
R1198 VDD.n1299 VDD.n1293 185
R1199 VDD.n1967 VDD.n1966 185
R1200 VDD.n1966 VDD.n1965 185
R1201 VDD.n1297 VDD.n1296 185
R1202 VDD.n1298 VDD.n1297 185
R1203 VDD.n1956 VDD.n1955 185
R1204 VDD.n1957 VDD.n1956 185
R1205 VDD.n1307 VDD.n1306 185
R1206 VDD.n1306 VDD.n1305 185
R1207 VDD.n1951 VDD.n1950 185
R1208 VDD.n1950 VDD.n1949 185
R1209 VDD.n1310 VDD.n1309 185
R1210 VDD.n1311 VDD.n1310 185
R1211 VDD.n1940 VDD.n1939 185
R1212 VDD.n1941 VDD.n1940 185
R1213 VDD.n1319 VDD.n1318 185
R1214 VDD.n1318 VDD.n1317 185
R1215 VDD.n1935 VDD.n1934 185
R1216 VDD.n1934 VDD.n1933 185
R1217 VDD.n1322 VDD.n1321 185
R1218 VDD.n1323 VDD.n1322 185
R1219 VDD.n1924 VDD.n1923 185
R1220 VDD.n1925 VDD.n1924 185
R1221 VDD.n1330 VDD.n1329 185
R1222 VDD.n1335 VDD.n1329 185
R1223 VDD.n1919 VDD.n1918 185
R1224 VDD.n1918 VDD.n1917 185
R1225 VDD.n1333 VDD.n1332 185
R1226 VDD.n1334 VDD.n1333 185
R1227 VDD.n1908 VDD.n1907 185
R1228 VDD.n1909 VDD.n1908 185
R1229 VDD.n1343 VDD.n1342 185
R1230 VDD.n1342 VDD.n1341 185
R1231 VDD.n1903 VDD.n1902 185
R1232 VDD.n1902 VDD.n1901 185
R1233 VDD.n1346 VDD.n1345 185
R1234 VDD.n1347 VDD.n1346 185
R1235 VDD.n1873 VDD.n1872 185
R1236 VDD.n1874 VDD.n1873 185
R1237 VDD.n1355 VDD.n1354 185
R1238 VDD.n1354 VDD.n1353 185
R1239 VDD.n1868 VDD.n1867 185
R1240 VDD.n1867 VDD.n1866 185
R1241 VDD.n1358 VDD.n1357 185
R1242 VDD.n1359 VDD.n1358 185
R1243 VDD.n1857 VDD.n1856 185
R1244 VDD.n1858 VDD.n1857 185
R1245 VDD.n1366 VDD.n1365 185
R1246 VDD.n1371 VDD.n1365 185
R1247 VDD.n1852 VDD.n1851 185
R1248 VDD.n1851 VDD.n1850 185
R1249 VDD.n1369 VDD.n1368 185
R1250 VDD.n1370 VDD.n1369 185
R1251 VDD.n1841 VDD.n1840 185
R1252 VDD.n1842 VDD.n1841 185
R1253 VDD.n1379 VDD.n1378 185
R1254 VDD.n1378 VDD.n1377 185
R1255 VDD.n1836 VDD.n1835 185
R1256 VDD.n1835 VDD.n1834 185
R1257 VDD.n1382 VDD.n1381 185
R1258 VDD.n1383 VDD.n1382 185
R1259 VDD.n1825 VDD.n1824 185
R1260 VDD.n1826 VDD.n1825 185
R1261 VDD.n1391 VDD.n1390 185
R1262 VDD.n1390 VDD.n1389 185
R1263 VDD.n1820 VDD.n1819 185
R1264 VDD.n1819 VDD.n1818 185
R1265 VDD.n1394 VDD.n1393 185
R1266 VDD.n1395 VDD.n1394 185
R1267 VDD.n1809 VDD.n1808 185
R1268 VDD.n1810 VDD.n1809 185
R1269 VDD.n1402 VDD.n1401 185
R1270 VDD.n1407 VDD.n1401 185
R1271 VDD.n1804 VDD.n1803 185
R1272 VDD.n1803 VDD.n1802 185
R1273 VDD.n1405 VDD.n1404 185
R1274 VDD.n1406 VDD.n1405 185
R1275 VDD.n1793 VDD.n1792 185
R1276 VDD.n1794 VDD.n1793 185
R1277 VDD.n1415 VDD.n1414 185
R1278 VDD.n1414 VDD.n1413 185
R1279 VDD.n1788 VDD.n1787 185
R1280 VDD.n1787 VDD.n1786 185
R1281 VDD.n1418 VDD.n1417 185
R1282 VDD.n1419 VDD.n1418 185
R1283 VDD.n1777 VDD.n1776 185
R1284 VDD.n1778 VDD.n1777 185
R1285 VDD.n1427 VDD.n1426 185
R1286 VDD.n1426 VDD.n1425 185
R1287 VDD.n1772 VDD.n1771 185
R1288 VDD.n1771 VDD.n1770 185
R1289 VDD.n1430 VDD.n1429 185
R1290 VDD.n1431 VDD.n1430 185
R1291 VDD.n1762 VDD.n1761 185
R1292 VDD.t91 VDD.n1762 185
R1293 VDD.n1439 VDD.n1438 185
R1294 VDD.n1438 VDD.n1437 185
R1295 VDD.n1757 VDD.n1756 185
R1296 VDD.n1756 VDD.n1755 185
R1297 VDD.n1442 VDD.n1441 185
R1298 VDD.n1443 VDD.n1442 185
R1299 VDD.n1746 VDD.n1745 185
R1300 VDD.n1747 VDD.n1746 185
R1301 VDD.n1451 VDD.n1450 185
R1302 VDD.n1450 VDD.n1449 185
R1303 VDD.n1741 VDD.n1740 185
R1304 VDD.n1740 VDD.n1739 185
R1305 VDD.n1454 VDD.n1453 185
R1306 VDD.n1455 VDD.n1454 185
R1307 VDD.n1730 VDD.n1729 185
R1308 VDD.n1731 VDD.n1730 185
R1309 VDD.n1463 VDD.n1462 185
R1310 VDD.n1462 VDD.n1461 185
R1311 VDD.n1725 VDD.n1724 185
R1312 VDD.n1724 VDD.n1723 185
R1313 VDD.n1466 VDD.n1465 185
R1314 VDD.n1467 VDD.n1466 185
R1315 VDD.n1714 VDD.n1713 185
R1316 VDD.n1715 VDD.n1714 185
R1317 VDD.n1475 VDD.n1474 185
R1318 VDD.n1474 VDD.n1473 185
R1319 VDD.n1709 VDD.n1708 185
R1320 VDD.n1708 VDD.n1707 185
R1321 VDD.n1478 VDD.n1477 185
R1322 VDD.n1698 VDD.n1478 185
R1323 VDD.n1697 VDD.n1696 185
R1324 VDD.n1699 VDD.n1697 185
R1325 VDD.n1486 VDD.n1485 185
R1326 VDD.n1485 VDD.n1484 185
R1327 VDD.n1692 VDD.n1691 185
R1328 VDD.n1691 VDD.n1690 185
R1329 VDD.n1489 VDD.n1488 185
R1330 VDD.n1490 VDD.n1489 185
R1331 VDD.n1681 VDD.n1680 185
R1332 VDD.n1682 VDD.n1681 185
R1333 VDD.n1498 VDD.n1497 185
R1334 VDD.n1497 VDD.n1496 185
R1335 VDD.n656 VDD.n654 185
R1336 VDD.n654 VDD.n628 185
R1337 VDD.n2731 VDD.n2730 185
R1338 VDD.n2732 VDD.n2731 185
R1339 VDD.n2729 VDD.n666 185
R1340 VDD.n666 VDD.n663 185
R1341 VDD.n2728 VDD.n2727 185
R1342 VDD.n2727 VDD.n2726 185
R1343 VDD.n668 VDD.n667 185
R1344 VDD.n669 VDD.n668 185
R1345 VDD.n2659 VDD.n2658 185
R1346 VDD.n2660 VDD.n2659 185
R1347 VDD.n2657 VDD.n682 185
R1348 VDD.n682 VDD.n679 185
R1349 VDD.n2656 VDD.n2655 185
R1350 VDD.n2655 VDD.n2654 185
R1351 VDD.n684 VDD.n683 185
R1352 VDD.n685 VDD.n684 185
R1353 VDD.n2645 VDD.n2644 185
R1354 VDD.n2646 VDD.n2645 185
R1355 VDD.n2643 VDD.n695 185
R1356 VDD.n695 VDD.n692 185
R1357 VDD.n2642 VDD.n2641 185
R1358 VDD.n2641 VDD.n2640 185
R1359 VDD.n697 VDD.n696 185
R1360 VDD.n698 VDD.n697 185
R1361 VDD.n2633 VDD.n2632 185
R1362 VDD.n2634 VDD.n2633 185
R1363 VDD.n2631 VDD.n707 185
R1364 VDD.n707 VDD.n704 185
R1365 VDD.n2630 VDD.n2629 185
R1366 VDD.n2629 VDD.n2628 185
R1367 VDD.n709 VDD.n708 185
R1368 VDD.n710 VDD.n709 185
R1369 VDD.n2621 VDD.n2620 185
R1370 VDD.n2622 VDD.n2621 185
R1371 VDD.n2619 VDD.n719 185
R1372 VDD.n719 VDD.n716 185
R1373 VDD.n2618 VDD.n2617 185
R1374 VDD.n2617 VDD.n2616 185
R1375 VDD.n721 VDD.n720 185
R1376 VDD.n730 VDD.n721 185
R1377 VDD.n2609 VDD.n2608 185
R1378 VDD.n2610 VDD.n2609 185
R1379 VDD.n2607 VDD.n731 185
R1380 VDD.n731 VDD.n727 185
R1381 VDD.n2606 VDD.n2605 185
R1382 VDD.n2605 VDD.n2604 185
R1383 VDD.n733 VDD.n732 185
R1384 VDD.n734 VDD.n733 185
R1385 VDD.n2597 VDD.n2596 185
R1386 VDD.n2598 VDD.n2597 185
R1387 VDD.n2595 VDD.n742 185
R1388 VDD.n748 VDD.n742 185
R1389 VDD.n2594 VDD.n2593 185
R1390 VDD.n2593 VDD.n2592 185
R1391 VDD.n744 VDD.n743 185
R1392 VDD.n745 VDD.n744 185
R1393 VDD.n2585 VDD.n2584 185
R1394 VDD.n2586 VDD.n2585 185
R1395 VDD.n2583 VDD.n755 185
R1396 VDD.n755 VDD.n752 185
R1397 VDD.n2582 VDD.n2581 185
R1398 VDD.n2581 VDD.n2580 185
R1399 VDD.n757 VDD.n756 185
R1400 VDD.n758 VDD.n757 185
R1401 VDD.n2573 VDD.n2572 185
R1402 VDD.n2574 VDD.n2573 185
R1403 VDD.n2571 VDD.n767 185
R1404 VDD.n767 VDD.n764 185
R1405 VDD.n2570 VDD.n2569 185
R1406 VDD.n2569 VDD.n2568 185
R1407 VDD.n769 VDD.n768 185
R1408 VDD.n770 VDD.n769 185
R1409 VDD.n2561 VDD.n2560 185
R1410 VDD.n2562 VDD.n2561 185
R1411 VDD.n2559 VDD.n779 185
R1412 VDD.n779 VDD.n776 185
R1413 VDD.n2558 VDD.n2557 185
R1414 VDD.n2557 VDD.n2556 185
R1415 VDD.n781 VDD.n780 185
R1416 VDD.n782 VDD.n781 185
R1417 VDD.n2549 VDD.n2548 185
R1418 VDD.n2550 VDD.n2549 185
R1419 VDD.n2547 VDD.n791 185
R1420 VDD.n791 VDD.n788 185
R1421 VDD.n2546 VDD.n2545 185
R1422 VDD.n2545 VDD.n2544 185
R1423 VDD.n793 VDD.n792 185
R1424 VDD.n794 VDD.n793 185
R1425 VDD.n2537 VDD.n2536 185
R1426 VDD.n2538 VDD.n2537 185
R1427 VDD.n2535 VDD.n802 185
R1428 VDD.n808 VDD.n802 185
R1429 VDD.n2534 VDD.n2533 185
R1430 VDD.n2533 VDD.n2532 185
R1431 VDD.n804 VDD.n803 185
R1432 VDD.n805 VDD.n804 185
R1433 VDD.n2525 VDD.n2524 185
R1434 VDD.n2526 VDD.n2525 185
R1435 VDD.n2523 VDD.n815 185
R1436 VDD.n815 VDD.n812 185
R1437 VDD.n2522 VDD.n2521 185
R1438 VDD.n2521 VDD.n2520 185
R1439 VDD.n817 VDD.n816 185
R1440 VDD.n818 VDD.n817 185
R1441 VDD.n2513 VDD.n2512 185
R1442 VDD.n2514 VDD.n2513 185
R1443 VDD.n2511 VDD.n827 185
R1444 VDD.n827 VDD.n824 185
R1445 VDD.n2510 VDD.n2509 185
R1446 VDD.n2509 VDD.n2508 185
R1447 VDD.n829 VDD.n828 185
R1448 VDD.n830 VDD.n829 185
R1449 VDD.n2501 VDD.n2500 185
R1450 VDD.n2502 VDD.n2501 185
R1451 VDD.n2499 VDD.n839 185
R1452 VDD.n839 VDD.n836 185
R1453 VDD.n2498 VDD.n2497 185
R1454 VDD.n2497 VDD.n2496 185
R1455 VDD.n841 VDD.n840 185
R1456 VDD.n842 VDD.n841 185
R1457 VDD.n2489 VDD.n2488 185
R1458 VDD.n2490 VDD.n2489 185
R1459 VDD.n2487 VDD.n851 185
R1460 VDD.n851 VDD.n848 185
R1461 VDD.n2486 VDD.n2485 185
R1462 VDD.n2485 VDD.n2484 185
R1463 VDD.n853 VDD.n852 185
R1464 VDD.n2357 VDD.n853 185
R1465 VDD.n2477 VDD.n2476 185
R1466 VDD.n2478 VDD.n2477 185
R1467 VDD.n2475 VDD.n862 185
R1468 VDD.n862 VDD.n859 185
R1469 VDD.n2474 VDD.n2473 185
R1470 VDD.n2473 VDD.n2472 185
R1471 VDD.n864 VDD.n863 185
R1472 VDD.n865 VDD.n864 185
R1473 VDD.n2465 VDD.n2464 185
R1474 VDD.n2466 VDD.n2465 185
R1475 VDD.n2463 VDD.n874 185
R1476 VDD.n874 VDD.n871 185
R1477 VDD.n2462 VDD.n2461 185
R1478 VDD.n2461 VDD.n2460 185
R1479 VDD.n876 VDD.n875 185
R1480 VDD.n877 VDD.n876 185
R1481 VDD.n2453 VDD.n2452 185
R1482 VDD.n2454 VDD.n2453 185
R1483 VDD.n2451 VDD.n886 185
R1484 VDD.n886 VDD.n883 185
R1485 VDD.n2450 VDD.n2449 185
R1486 VDD.n2449 VDD.n2448 185
R1487 VDD.n888 VDD.n887 185
R1488 VDD.n889 VDD.n888 185
R1489 VDD.n2441 VDD.n2440 185
R1490 VDD.n2442 VDD.n2441 185
R1491 VDD.n2439 VDD.n897 185
R1492 VDD.n903 VDD.n897 185
R1493 VDD.n2438 VDD.n2437 185
R1494 VDD.n2437 VDD.n2436 185
R1495 VDD.n899 VDD.n898 185
R1496 VDD.n900 VDD.n899 185
R1497 VDD.n2429 VDD.n2428 185
R1498 VDD.n2430 VDD.n2429 185
R1499 VDD.n2427 VDD.n910 185
R1500 VDD.n910 VDD.n907 185
R1501 VDD.n2426 VDD.n2425 185
R1502 VDD.n2425 VDD.n2424 185
R1503 VDD.n912 VDD.n911 185
R1504 VDD.n913 VDD.n912 185
R1505 VDD.n2417 VDD.n2416 185
R1506 VDD.n2418 VDD.n2417 185
R1507 VDD.n2415 VDD.n922 185
R1508 VDD.n922 VDD.n919 185
R1509 VDD.n2414 VDD.n2413 185
R1510 VDD.n2413 VDD.n2412 185
R1511 VDD.n924 VDD.n923 185
R1512 VDD.n925 VDD.n924 185
R1513 VDD.n2405 VDD.n2404 185
R1514 VDD.n2406 VDD.n2405 185
R1515 VDD.n2403 VDD.n933 185
R1516 VDD.n2402 VDD.n2401 185
R1517 VDD.n935 VDD.n934 185
R1518 VDD.n2399 VDD.n935 185
R1519 VDD.n1051 VDD.n1050 185
R1520 VDD.n1053 VDD.n1052 185
R1521 VDD.n1055 VDD.n1054 185
R1522 VDD.n1057 VDD.n1056 185
R1523 VDD.n1059 VDD.n1058 185
R1524 VDD.n1061 VDD.n1060 185
R1525 VDD.n1063 VDD.n1062 185
R1526 VDD.n1065 VDD.n1064 185
R1527 VDD.n1067 VDD.n1066 185
R1528 VDD.n2201 VDD.n2200 185
R1529 VDD.n2203 VDD.n2202 185
R1530 VDD.n2205 VDD.n2204 185
R1531 VDD.n2207 VDD.n2206 185
R1532 VDD.n2209 VDD.n2208 185
R1533 VDD.n2211 VDD.n2210 185
R1534 VDD.n2213 VDD.n2212 185
R1535 VDD.n2215 VDD.n2214 185
R1536 VDD.n2217 VDD.n2216 185
R1537 VDD.n2219 VDD.n2218 185
R1538 VDD.n2221 VDD.n2220 185
R1539 VDD.n2223 VDD.n2222 185
R1540 VDD.n2225 VDD.n2224 185
R1541 VDD.n2736 VDD.n2735 185
R1542 VDD.n2738 VDD.n2737 185
R1543 VDD.n2740 VDD.n2739 185
R1544 VDD.n2742 VDD.n2741 185
R1545 VDD.n2744 VDD.n2743 185
R1546 VDD.n2746 VDD.n2745 185
R1547 VDD.n2748 VDD.n2747 185
R1548 VDD.n2750 VDD.n2749 185
R1549 VDD.n2752 VDD.n2751 185
R1550 VDD.n2754 VDD.n2753 185
R1551 VDD.n2756 VDD.n2755 185
R1552 VDD.n2758 VDD.n2757 185
R1553 VDD.n2760 VDD.n2759 185
R1554 VDD.n2762 VDD.n2761 185
R1555 VDD.n2764 VDD.n2763 185
R1556 VDD.n2766 VDD.n2765 185
R1557 VDD.n2768 VDD.n2767 185
R1558 VDD.n2770 VDD.n2769 185
R1559 VDD.n2772 VDD.n2771 185
R1560 VDD.n2774 VDD.n2773 185
R1561 VDD.n2776 VDD.n2775 185
R1562 VDD.n2778 VDD.n2777 185
R1563 VDD.n2780 VDD.n2779 185
R1564 VDD.n2781 VDD.n655 185
R1565 VDD.n2783 VDD.n2782 185
R1566 VDD.n2784 VDD.n2783 185
R1567 VDD.n2734 VDD.n660 185
R1568 VDD.n2734 VDD.n628 185
R1569 VDD.n2733 VDD.n662 185
R1570 VDD.n2733 VDD.n2732 185
R1571 VDD.n2263 VDD.n661 185
R1572 VDD.n663 VDD.n661 185
R1573 VDD.n2264 VDD.n670 185
R1574 VDD.n2726 VDD.n670 185
R1575 VDD.n2266 VDD.n2265 185
R1576 VDD.n2265 VDD.n669 185
R1577 VDD.n2267 VDD.n680 185
R1578 VDD.n2660 VDD.n680 185
R1579 VDD.n2269 VDD.n2268 185
R1580 VDD.n2268 VDD.n679 185
R1581 VDD.n2270 VDD.n686 185
R1582 VDD.n2654 VDD.n686 185
R1583 VDD.n2272 VDD.n2271 185
R1584 VDD.n2271 VDD.n685 185
R1585 VDD.n2273 VDD.n693 185
R1586 VDD.n2646 VDD.n693 185
R1587 VDD.n2275 VDD.n2274 185
R1588 VDD.n2274 VDD.n692 185
R1589 VDD.n2276 VDD.n699 185
R1590 VDD.n2640 VDD.n699 185
R1591 VDD.n2278 VDD.n2277 185
R1592 VDD.n2277 VDD.n698 185
R1593 VDD.n2279 VDD.n705 185
R1594 VDD.n2634 VDD.n705 185
R1595 VDD.n2281 VDD.n2280 185
R1596 VDD.n2280 VDD.n704 185
R1597 VDD.n2282 VDD.n711 185
R1598 VDD.n2628 VDD.n711 185
R1599 VDD.n2284 VDD.n2283 185
R1600 VDD.n2283 VDD.n710 185
R1601 VDD.n2285 VDD.n717 185
R1602 VDD.n2622 VDD.n717 185
R1603 VDD.n2287 VDD.n2286 185
R1604 VDD.n2286 VDD.n716 185
R1605 VDD.n2288 VDD.n722 185
R1606 VDD.n2616 VDD.n722 185
R1607 VDD.n2290 VDD.n2289 185
R1608 VDD.n2289 VDD.n730 185
R1609 VDD.n2291 VDD.n728 185
R1610 VDD.n2610 VDD.n728 185
R1611 VDD.n2293 VDD.n2292 185
R1612 VDD.n2292 VDD.n727 185
R1613 VDD.n2294 VDD.n735 185
R1614 VDD.n2604 VDD.n735 185
R1615 VDD.n2296 VDD.n2295 185
R1616 VDD.n2295 VDD.n734 185
R1617 VDD.n2297 VDD.n740 185
R1618 VDD.n2598 VDD.n740 185
R1619 VDD.n2299 VDD.n2298 185
R1620 VDD.n2298 VDD.n748 185
R1621 VDD.n2300 VDD.n746 185
R1622 VDD.n2592 VDD.n746 185
R1623 VDD.n2302 VDD.n2301 185
R1624 VDD.n2301 VDD.n745 185
R1625 VDD.n2303 VDD.n753 185
R1626 VDD.n2586 VDD.n753 185
R1627 VDD.n2305 VDD.n2304 185
R1628 VDD.n2304 VDD.n752 185
R1629 VDD.n2306 VDD.n759 185
R1630 VDD.n2580 VDD.n759 185
R1631 VDD.n2308 VDD.n2307 185
R1632 VDD.n2307 VDD.n758 185
R1633 VDD.n2309 VDD.n765 185
R1634 VDD.n2574 VDD.n765 185
R1635 VDD.n2311 VDD.n2310 185
R1636 VDD.n2310 VDD.n764 185
R1637 VDD.n2312 VDD.n771 185
R1638 VDD.n2568 VDD.n771 185
R1639 VDD.n2314 VDD.n2313 185
R1640 VDD.n2313 VDD.n770 185
R1641 VDD.n2315 VDD.n777 185
R1642 VDD.n2562 VDD.n777 185
R1643 VDD.n2317 VDD.n2316 185
R1644 VDD.n2316 VDD.n776 185
R1645 VDD.n2318 VDD.n783 185
R1646 VDD.n2556 VDD.n783 185
R1647 VDD.n2320 VDD.n2319 185
R1648 VDD.n2319 VDD.n782 185
R1649 VDD.n2321 VDD.n789 185
R1650 VDD.n2550 VDD.n789 185
R1651 VDD.n2323 VDD.n2322 185
R1652 VDD.n2322 VDD.n788 185
R1653 VDD.n2324 VDD.n795 185
R1654 VDD.n2544 VDD.n795 185
R1655 VDD.n2326 VDD.n2325 185
R1656 VDD.n2325 VDD.n794 185
R1657 VDD.n2327 VDD.n800 185
R1658 VDD.n2538 VDD.n800 185
R1659 VDD.n2329 VDD.n2328 185
R1660 VDD.n2328 VDD.n808 185
R1661 VDD.n2330 VDD.n806 185
R1662 VDD.n2532 VDD.n806 185
R1663 VDD.n2332 VDD.n2331 185
R1664 VDD.n2331 VDD.n805 185
R1665 VDD.n2333 VDD.n813 185
R1666 VDD.n2526 VDD.n813 185
R1667 VDD.n2335 VDD.n2334 185
R1668 VDD.n2334 VDD.n812 185
R1669 VDD.n2336 VDD.n819 185
R1670 VDD.n2520 VDD.n819 185
R1671 VDD.n2338 VDD.n2337 185
R1672 VDD.n2337 VDD.n818 185
R1673 VDD.n2339 VDD.n825 185
R1674 VDD.n2514 VDD.n825 185
R1675 VDD.n2341 VDD.n2340 185
R1676 VDD.n2340 VDD.n824 185
R1677 VDD.n2342 VDD.n831 185
R1678 VDD.n2508 VDD.n831 185
R1679 VDD.n2344 VDD.n2343 185
R1680 VDD.n2343 VDD.n830 185
R1681 VDD.n2345 VDD.n837 185
R1682 VDD.n2502 VDD.n837 185
R1683 VDD.n2347 VDD.n2346 185
R1684 VDD.n2346 VDD.n836 185
R1685 VDD.n2348 VDD.n843 185
R1686 VDD.n2496 VDD.n843 185
R1687 VDD.n2350 VDD.n2349 185
R1688 VDD.n2349 VDD.n842 185
R1689 VDD.n2351 VDD.n849 185
R1690 VDD.n2490 VDD.n849 185
R1691 VDD.n2353 VDD.n2352 185
R1692 VDD.n2352 VDD.n848 185
R1693 VDD.n2354 VDD.n854 185
R1694 VDD.n2484 VDD.n854 185
R1695 VDD.n2356 VDD.n2355 185
R1696 VDD.n2357 VDD.n2356 185
R1697 VDD.n2262 VDD.n860 185
R1698 VDD.n2478 VDD.n860 185
R1699 VDD.n2261 VDD.n2260 185
R1700 VDD.n2260 VDD.n859 185
R1701 VDD.n2259 VDD.n866 185
R1702 VDD.n2472 VDD.n866 185
R1703 VDD.n2258 VDD.n2257 185
R1704 VDD.n2257 VDD.n865 185
R1705 VDD.n2256 VDD.n872 185
R1706 VDD.n2466 VDD.n872 185
R1707 VDD.n2255 VDD.n2254 185
R1708 VDD.n2254 VDD.n871 185
R1709 VDD.n2253 VDD.n878 185
R1710 VDD.n2460 VDD.n878 185
R1711 VDD.n2252 VDD.n2251 185
R1712 VDD.n2251 VDD.n877 185
R1713 VDD.n2250 VDD.n884 185
R1714 VDD.n2454 VDD.n884 185
R1715 VDD.n2249 VDD.n2248 185
R1716 VDD.n2248 VDD.n883 185
R1717 VDD.n2247 VDD.n890 185
R1718 VDD.n2448 VDD.n890 185
R1719 VDD.n2246 VDD.n2245 185
R1720 VDD.n2245 VDD.n889 185
R1721 VDD.n2244 VDD.n895 185
R1722 VDD.n2442 VDD.n895 185
R1723 VDD.n2243 VDD.n2242 185
R1724 VDD.n2242 VDD.n903 185
R1725 VDD.n2241 VDD.n901 185
R1726 VDD.n2436 VDD.n901 185
R1727 VDD.n2240 VDD.n2239 185
R1728 VDD.n2239 VDD.n900 185
R1729 VDD.n2238 VDD.n908 185
R1730 VDD.n2430 VDD.n908 185
R1731 VDD.n2237 VDD.n2236 185
R1732 VDD.n2236 VDD.n907 185
R1733 VDD.n2235 VDD.n914 185
R1734 VDD.n2424 VDD.n914 185
R1735 VDD.n2234 VDD.n2233 185
R1736 VDD.n2233 VDD.n913 185
R1737 VDD.n2232 VDD.n920 185
R1738 VDD.n2418 VDD.n920 185
R1739 VDD.n2231 VDD.n2230 185
R1740 VDD.n2230 VDD.n919 185
R1741 VDD.n2229 VDD.n926 185
R1742 VDD.n2412 VDD.n926 185
R1743 VDD.n2228 VDD.n2227 185
R1744 VDD.n2227 VDD.n925 185
R1745 VDD.n2226 VDD.n931 185
R1746 VDD.n2406 VDD.n931 185
R1747 VDD.n3999 VDD.n3998 185
R1748 VDD.n4223 VDD.n3999 185
R1749 VDD.n4226 VDD.n4225 185
R1750 VDD.n4225 VDD.n4224 185
R1751 VDD.n4227 VDD.n3993 185
R1752 VDD.n3993 VDD.n3992 185
R1753 VDD.n4229 VDD.n4228 185
R1754 VDD.n4230 VDD.n4229 185
R1755 VDD.n3987 VDD.n3986 185
R1756 VDD.n4231 VDD.n3987 185
R1757 VDD.n4234 VDD.n4233 185
R1758 VDD.n4233 VDD.n4232 185
R1759 VDD.n4235 VDD.n3981 185
R1760 VDD.n3988 VDD.n3981 185
R1761 VDD.n4237 VDD.n4236 185
R1762 VDD.n4238 VDD.n4237 185
R1763 VDD.n3977 VDD.n3976 185
R1764 VDD.n4239 VDD.n3977 185
R1765 VDD.n4242 VDD.n4241 185
R1766 VDD.n4241 VDD.n4240 185
R1767 VDD.n4243 VDD.n3971 185
R1768 VDD.n3971 VDD.n3970 185
R1769 VDD.n4245 VDD.n4244 185
R1770 VDD.n4246 VDD.n4245 185
R1771 VDD.n3966 VDD.n3965 185
R1772 VDD.n4247 VDD.n3966 185
R1773 VDD.n4250 VDD.n4249 185
R1774 VDD.n4249 VDD.n4248 185
R1775 VDD.n4251 VDD.n3960 185
R1776 VDD.n3960 VDD.n3959 185
R1777 VDD.n4253 VDD.n4252 185
R1778 VDD.n4254 VDD.n4253 185
R1779 VDD.n3955 VDD.n3954 185
R1780 VDD.n4255 VDD.n3955 185
R1781 VDD.n4258 VDD.n4257 185
R1782 VDD.n4257 VDD.n4256 185
R1783 VDD.n4259 VDD.n3949 185
R1784 VDD.n3949 VDD.n3948 185
R1785 VDD.n4261 VDD.n4260 185
R1786 VDD.n4262 VDD.n4261 185
R1787 VDD.n116 VDD.n115 185
R1788 VDD.n117 VDD.n116 185
R1789 VDD.n4269 VDD.n4268 185
R1790 VDD.n4268 VDD.t99 185
R1791 VDD.n4270 VDD.n110 185
R1792 VDD.n110 VDD.n109 185
R1793 VDD.n4272 VDD.n4271 185
R1794 VDD.n4273 VDD.n4272 185
R1795 VDD.n105 VDD.n104 185
R1796 VDD.n4274 VDD.n105 185
R1797 VDD.n4277 VDD.n4276 185
R1798 VDD.n4276 VDD.n4275 185
R1799 VDD.n4278 VDD.n99 185
R1800 VDD.n99 VDD.n98 185
R1801 VDD.n4280 VDD.n4279 185
R1802 VDD.n4281 VDD.n4280 185
R1803 VDD.n94 VDD.n93 185
R1804 VDD.n4282 VDD.n94 185
R1805 VDD.n4285 VDD.n4284 185
R1806 VDD.n4284 VDD.n4283 185
R1807 VDD.n4286 VDD.n88 185
R1808 VDD.n88 VDD.n87 185
R1809 VDD.n4288 VDD.n4287 185
R1810 VDD.n4289 VDD.n4288 185
R1811 VDD.n83 VDD.n82 185
R1812 VDD.n4290 VDD.n83 185
R1813 VDD.n4293 VDD.n4292 185
R1814 VDD.n4292 VDD.n4291 185
R1815 VDD.n4294 VDD.n77 185
R1816 VDD.n77 VDD.n76 185
R1817 VDD.n4296 VDD.n4295 185
R1818 VDD.n4297 VDD.n4296 185
R1819 VDD.n72 VDD.n71 185
R1820 VDD.n4298 VDD.n72 185
R1821 VDD.n4301 VDD.n4300 185
R1822 VDD.n4300 VDD.n4299 185
R1823 VDD.n4302 VDD.n66 185
R1824 VDD.n66 VDD.n65 185
R1825 VDD.n4304 VDD.n4303 185
R1826 VDD.n4305 VDD.n4304 185
R1827 VDD.n61 VDD.n60 185
R1828 VDD.n4306 VDD.n61 185
R1829 VDD.n4309 VDD.n4308 185
R1830 VDD.n4308 VDD.n4307 185
R1831 VDD.n4310 VDD.n55 185
R1832 VDD.n55 VDD.n54 185
R1833 VDD.n4312 VDD.n4311 185
R1834 VDD.n4313 VDD.n4312 185
R1835 VDD.n50 VDD.n49 185
R1836 VDD.n4314 VDD.n50 185
R1837 VDD.n4317 VDD.n4316 185
R1838 VDD.n4316 VDD.n4315 185
R1839 VDD.n4318 VDD.n44 185
R1840 VDD.n44 VDD.n43 185
R1841 VDD.n4320 VDD.n4319 185
R1842 VDD.n4321 VDD.n4320 185
R1843 VDD.n38 VDD.n37 185
R1844 VDD.n4322 VDD.n38 185
R1845 VDD.n4325 VDD.n4324 185
R1846 VDD.n4324 VDD.n4323 185
R1847 VDD.n4326 VDD.n36 185
R1848 VDD.n39 VDD.n36 185
R1849 VDD.n3895 VDD.n35 185
R1850 VDD.n3896 VDD.n3895 185
R1851 VDD.n3894 VDD.n3893 185
R1852 VDD.n3894 VDD.n145 185
R1853 VDD.n147 VDD.n146 185
R1854 VDD.n3886 VDD.n146 185
R1855 VDD.n3889 VDD.n3888 185
R1856 VDD.n3888 VDD.n3887 185
R1857 VDD.n150 VDD.n149 185
R1858 VDD.n151 VDD.n150 185
R1859 VDD.n3876 VDD.n3875 185
R1860 VDD.n3877 VDD.n3876 185
R1861 VDD.n158 VDD.n157 185
R1862 VDD.n3868 VDD.n157 185
R1863 VDD.n3871 VDD.n3870 185
R1864 VDD.n3870 VDD.n3869 185
R1865 VDD.n161 VDD.n160 185
R1866 VDD.n162 VDD.n161 185
R1867 VDD.n3857 VDD.n3856 185
R1868 VDD.n3858 VDD.n3857 185
R1869 VDD.n170 VDD.n169 185
R1870 VDD.n169 VDD.n168 185
R1871 VDD.n3852 VDD.n3851 185
R1872 VDD.n3851 VDD.n3850 185
R1873 VDD.n173 VDD.n172 185
R1874 VDD.n174 VDD.n173 185
R1875 VDD.n3841 VDD.n3840 185
R1876 VDD.n3842 VDD.n3841 185
R1877 VDD.n182 VDD.n181 185
R1878 VDD.n181 VDD.n180 185
R1879 VDD.n3836 VDD.n3835 185
R1880 VDD.n3835 VDD.n3834 185
R1881 VDD.n185 VDD.n184 185
R1882 VDD.n186 VDD.n185 185
R1883 VDD.n3825 VDD.n3824 185
R1884 VDD.n3826 VDD.n3825 185
R1885 VDD.n193 VDD.n192 185
R1886 VDD.n3817 VDD.n192 185
R1887 VDD.n3820 VDD.n3819 185
R1888 VDD.n3819 VDD.n3818 185
R1889 VDD.n196 VDD.n195 185
R1890 VDD.n197 VDD.n196 185
R1891 VDD.n3808 VDD.n3807 185
R1892 VDD.n3809 VDD.n3808 185
R1893 VDD.n205 VDD.n204 185
R1894 VDD.n204 VDD.n203 185
R1895 VDD.n3803 VDD.n3802 185
R1896 VDD.n3802 VDD.n3801 185
R1897 VDD.n208 VDD.n207 185
R1898 VDD.n209 VDD.n208 185
R1899 VDD.n3792 VDD.n3791 185
R1900 VDD.n3793 VDD.n3792 185
R1901 VDD.n217 VDD.n216 185
R1902 VDD.n216 VDD.n215 185
R1903 VDD.n3787 VDD.n3786 185
R1904 VDD.n3786 VDD.n3785 185
R1905 VDD.n220 VDD.n219 185
R1906 VDD.n221 VDD.n220 185
R1907 VDD.n3777 VDD.n3776 185
R1908 VDD.t81 VDD.n3777 185
R1909 VDD.n229 VDD.n228 185
R1910 VDD.n228 VDD.n227 185
R1911 VDD.n3772 VDD.n3771 185
R1912 VDD.n3771 VDD.n3770 185
R1913 VDD.n232 VDD.n231 185
R1914 VDD.n233 VDD.n232 185
R1915 VDD.n3761 VDD.n3760 185
R1916 VDD.n3762 VDD.n3761 185
R1917 VDD.n241 VDD.n240 185
R1918 VDD.n240 VDD.n239 185
R1919 VDD.n3756 VDD.n3755 185
R1920 VDD.n3755 VDD.n3754 185
R1921 VDD.n244 VDD.n243 185
R1922 VDD.n245 VDD.n244 185
R1923 VDD.n3745 VDD.n3744 185
R1924 VDD.n3746 VDD.n3745 185
R1925 VDD.n253 VDD.n252 185
R1926 VDD.n252 VDD.n251 185
R1927 VDD.n3740 VDD.n3739 185
R1928 VDD.n3739 VDD.n3738 185
R1929 VDD.n256 VDD.n255 185
R1930 VDD.n257 VDD.n256 185
R1931 VDD.n3729 VDD.n3728 185
R1932 VDD.n3730 VDD.n3729 185
R1933 VDD.n265 VDD.n264 185
R1934 VDD.n264 VDD.n263 185
R1935 VDD.n3724 VDD.n3723 185
R1936 VDD.n3723 VDD.n3722 185
R1937 VDD.n268 VDD.n267 185
R1938 VDD.n275 VDD.n268 185
R1939 VDD.n3713 VDD.n3712 185
R1940 VDD.n3714 VDD.n3713 185
R1941 VDD.n277 VDD.n276 185
R1942 VDD.n276 VDD.n274 185
R1943 VDD.n3708 VDD.n3707 185
R1944 VDD.n3707 VDD.n3706 185
R1945 VDD.n280 VDD.n279 185
R1946 VDD.n281 VDD.n280 185
R1947 VDD.n3697 VDD.n3696 185
R1948 VDD.n3698 VDD.n3697 185
R1949 VDD.n289 VDD.n288 185
R1950 VDD.n288 VDD.n287 185
R1951 VDD.n3685 VDD.n3684 185
R1952 VDD.n3683 VDD.n3682 185
R1953 VDD.n3688 VDD.n3682 185
R1954 VDD.n297 VDD.n294 185
R1955 VDD.n3691 VDD.n3690 185
R1956 VDD.n296 VDD.n295 185
R1957 VDD.n3572 VDD.n3571 185
R1958 VDD.n3570 VDD.n3569 185
R1959 VDD.n3577 VDD.n3576 185
R1960 VDD.n3579 VDD.n3578 185
R1961 VDD.n3582 VDD.n3581 185
R1962 VDD.n3580 VDD.n3567 185
R1963 VDD.n3587 VDD.n3586 185
R1964 VDD.n3589 VDD.n3588 185
R1965 VDD.n3594 VDD.n3591 185
R1966 VDD.n3590 VDD.n3565 185
R1967 VDD.n3599 VDD.n3598 185
R1968 VDD.n3601 VDD.n3600 185
R1969 VDD.n3604 VDD.n3603 185
R1970 VDD.n3602 VDD.n3563 185
R1971 VDD.n3609 VDD.n3608 185
R1972 VDD.n3611 VDD.n3610 185
R1973 VDD.n3614 VDD.n3613 185
R1974 VDD.n3612 VDD.n3561 185
R1975 VDD.n3619 VDD.n3618 185
R1976 VDD.n3621 VDD.n3620 185
R1977 VDD.n3624 VDD.n3623 185
R1978 VDD.n3622 VDD.n3559 185
R1979 VDD.n3629 VDD.n3628 185
R1980 VDD.n3631 VDD.n3630 185
R1981 VDD.n3637 VDD.n3636 185
R1982 VDD.n3635 VDD.n3557 185
R1983 VDD.n3642 VDD.n3641 185
R1984 VDD.n3644 VDD.n3643 185
R1985 VDD.n3647 VDD.n3646 185
R1986 VDD.n3645 VDD.n3555 185
R1987 VDD.n3652 VDD.n3651 185
R1988 VDD.n3654 VDD.n3653 185
R1989 VDD.n3657 VDD.n3656 185
R1990 VDD.n3655 VDD.n3553 185
R1991 VDD.n3662 VDD.n3661 185
R1992 VDD.n3664 VDD.n3663 185
R1993 VDD.n3667 VDD.n3666 185
R1994 VDD.n3665 VDD.n3551 185
R1995 VDD.n3672 VDD.n3671 185
R1996 VDD.n3674 VDD.n3673 185
R1997 VDD.n3677 VDD.n3676 185
R1998 VDD.n3678 VDD.n319 185
R1999 VDD.n4079 VDD.n4078 185
R2000 VDD.n4126 VDD.n4125 185
R2001 VDD.n4128 VDD.n4127 185
R2002 VDD.n4130 VDD.n4129 185
R2003 VDD.n4132 VDD.n4131 185
R2004 VDD.n4134 VDD.n4133 185
R2005 VDD.n4136 VDD.n4135 185
R2006 VDD.n4138 VDD.n4137 185
R2007 VDD.n4140 VDD.n4139 185
R2008 VDD.n4142 VDD.n4141 185
R2009 VDD.n4144 VDD.n4143 185
R2010 VDD.n4146 VDD.n4145 185
R2011 VDD.n4148 VDD.n4147 185
R2012 VDD.n4150 VDD.n4149 185
R2013 VDD.n4152 VDD.n4151 185
R2014 VDD.n4154 VDD.n4153 185
R2015 VDD.n4156 VDD.n4155 185
R2016 VDD.n4158 VDD.n4157 185
R2017 VDD.n4160 VDD.n4159 185
R2018 VDD.n4162 VDD.n4161 185
R2019 VDD.n4164 VDD.n4163 185
R2020 VDD.n4166 VDD.n4165 185
R2021 VDD.n4168 VDD.n4167 185
R2022 VDD.n4170 VDD.n4169 185
R2023 VDD.n4172 VDD.n4171 185
R2024 VDD.n4174 VDD.n4173 185
R2025 VDD.n4176 VDD.n4175 185
R2026 VDD.n4178 VDD.n4177 185
R2027 VDD.n4180 VDD.n4179 185
R2028 VDD.n4182 VDD.n4181 185
R2029 VDD.n4184 VDD.n4183 185
R2030 VDD.n4186 VDD.n4185 185
R2031 VDD.n4188 VDD.n4187 185
R2032 VDD.n4043 VDD.n4040 185
R2033 VDD.n4192 VDD.n4044 185
R2034 VDD.n4194 VDD.n4193 185
R2035 VDD.n4196 VDD.n4195 185
R2036 VDD.n4198 VDD.n4197 185
R2037 VDD.n4200 VDD.n4199 185
R2038 VDD.n4202 VDD.n4201 185
R2039 VDD.n4204 VDD.n4203 185
R2040 VDD.n4206 VDD.n4205 185
R2041 VDD.n4208 VDD.n4207 185
R2042 VDD.n4210 VDD.n4209 185
R2043 VDD.n4212 VDD.n4211 185
R2044 VDD.n4215 VDD.n4214 185
R2045 VDD.n4213 VDD.n4029 185
R2046 VDD.n4219 VDD.n4026 185
R2047 VDD.n4221 VDD.n4220 185
R2048 VDD.n4222 VDD.n4221 185
R2049 VDD.n4121 VDD.n4001 185
R2050 VDD.n4223 VDD.n4001 185
R2051 VDD.n4120 VDD.n4000 185
R2052 VDD.n4224 VDD.n4000 185
R2053 VDD.n4119 VDD.n4118 185
R2054 VDD.n4118 VDD.n3992 185
R2055 VDD.n4083 VDD.n3991 185
R2056 VDD.n4230 VDD.n3991 185
R2057 VDD.n4114 VDD.n3990 185
R2058 VDD.n4231 VDD.n3990 185
R2059 VDD.n4113 VDD.n3989 185
R2060 VDD.n4232 VDD.n3989 185
R2061 VDD.n4112 VDD.n4111 185
R2062 VDD.n4111 VDD.n3988 185
R2063 VDD.n4085 VDD.n3980 185
R2064 VDD.n4238 VDD.n3980 185
R2065 VDD.n4107 VDD.n3979 185
R2066 VDD.n4239 VDD.n3979 185
R2067 VDD.n4106 VDD.n3978 185
R2068 VDD.n4240 VDD.n3978 185
R2069 VDD.n4105 VDD.n4104 185
R2070 VDD.n4104 VDD.n3970 185
R2071 VDD.n4087 VDD.n3969 185
R2072 VDD.n4246 VDD.n3969 185
R2073 VDD.n4100 VDD.n3968 185
R2074 VDD.n4247 VDD.n3968 185
R2075 VDD.n4099 VDD.n3967 185
R2076 VDD.n4248 VDD.n3967 185
R2077 VDD.n4098 VDD.n4097 185
R2078 VDD.n4097 VDD.n3959 185
R2079 VDD.n4089 VDD.n3958 185
R2080 VDD.n4254 VDD.n3958 185
R2081 VDD.n4093 VDD.n3957 185
R2082 VDD.n4255 VDD.n3957 185
R2083 VDD.n4092 VDD.n3956 185
R2084 VDD.n4256 VDD.n3956 185
R2085 VDD.n3947 VDD.n3946 185
R2086 VDD.n3948 VDD.n3947 185
R2087 VDD.n4264 VDD.n4263 185
R2088 VDD.n4263 VDD.n4262 185
R2089 VDD.n4265 VDD.n119 185
R2090 VDD.n119 VDD.n117 185
R2091 VDD.n4267 VDD.n4266 185
R2092 VDD.t99 VDD.n4267 185
R2093 VDD.n120 VDD.n118 185
R2094 VDD.n118 VDD.n109 185
R2095 VDD.n3940 VDD.n108 185
R2096 VDD.n4273 VDD.n108 185
R2097 VDD.n3939 VDD.n107 185
R2098 VDD.n4274 VDD.n107 185
R2099 VDD.n3938 VDD.n106 185
R2100 VDD.n4275 VDD.n106 185
R2101 VDD.n123 VDD.n122 185
R2102 VDD.n122 VDD.n98 185
R2103 VDD.n3934 VDD.n97 185
R2104 VDD.n4281 VDD.n97 185
R2105 VDD.n3933 VDD.n96 185
R2106 VDD.n4282 VDD.n96 185
R2107 VDD.n3932 VDD.n95 185
R2108 VDD.n4283 VDD.n95 185
R2109 VDD.n126 VDD.n125 185
R2110 VDD.n125 VDD.n87 185
R2111 VDD.n3928 VDD.n86 185
R2112 VDD.n4289 VDD.n86 185
R2113 VDD.n3927 VDD.n85 185
R2114 VDD.n4290 VDD.n85 185
R2115 VDD.n3926 VDD.n84 185
R2116 VDD.n4291 VDD.n84 185
R2117 VDD.n129 VDD.n128 185
R2118 VDD.n128 VDD.n76 185
R2119 VDD.n3922 VDD.n75 185
R2120 VDD.n4297 VDD.n75 185
R2121 VDD.n3921 VDD.n74 185
R2122 VDD.n4298 VDD.n74 185
R2123 VDD.n3920 VDD.n73 185
R2124 VDD.n4299 VDD.n73 185
R2125 VDD.n132 VDD.n131 185
R2126 VDD.n131 VDD.n65 185
R2127 VDD.n3916 VDD.n64 185
R2128 VDD.n4305 VDD.n64 185
R2129 VDD.n3915 VDD.n63 185
R2130 VDD.n4306 VDD.n63 185
R2131 VDD.n3914 VDD.n62 185
R2132 VDD.n4307 VDD.n62 185
R2133 VDD.n135 VDD.n134 185
R2134 VDD.n134 VDD.n54 185
R2135 VDD.n3910 VDD.n53 185
R2136 VDD.n4313 VDD.n53 185
R2137 VDD.n3909 VDD.n52 185
R2138 VDD.n4314 VDD.n52 185
R2139 VDD.n3908 VDD.n51 185
R2140 VDD.n4315 VDD.n51 185
R2141 VDD.n138 VDD.n137 185
R2142 VDD.n137 VDD.n43 185
R2143 VDD.n3904 VDD.n42 185
R2144 VDD.n4321 VDD.n42 185
R2145 VDD.n3903 VDD.n41 185
R2146 VDD.n4322 VDD.n41 185
R2147 VDD.n3902 VDD.n40 185
R2148 VDD.n4323 VDD.n40 185
R2149 VDD.n144 VDD.n140 185
R2150 VDD.n144 VDD.n39 185
R2151 VDD.n3898 VDD.n3897 185
R2152 VDD.n3897 VDD.n3896 185
R2153 VDD.n143 VDD.n142 185
R2154 VDD.n145 VDD.n143 185
R2155 VDD.n3885 VDD.n3884 185
R2156 VDD.n3886 VDD.n3885 185
R2157 VDD.n153 VDD.n152 185
R2158 VDD.n3887 VDD.n152 185
R2159 VDD.n3880 VDD.n3879 185
R2160 VDD.n3879 VDD.n151 185
R2161 VDD.n3878 VDD.n155 185
R2162 VDD.n3878 VDD.n3877 185
R2163 VDD.n3865 VDD.n156 185
R2164 VDD.n3868 VDD.n156 185
R2165 VDD.n3867 VDD.n3866 185
R2166 VDD.n3869 VDD.n3867 185
R2167 VDD.n164 VDD.n163 185
R2168 VDD.n163 VDD.n162 185
R2169 VDD.n3860 VDD.n3859 185
R2170 VDD.n3859 VDD.n3858 185
R2171 VDD.n167 VDD.n166 185
R2172 VDD.n168 VDD.n167 185
R2173 VDD.n3849 VDD.n3848 185
R2174 VDD.n3850 VDD.n3849 185
R2175 VDD.n176 VDD.n175 185
R2176 VDD.n175 VDD.n174 185
R2177 VDD.n3844 VDD.n3843 185
R2178 VDD.n3843 VDD.n3842 185
R2179 VDD.n179 VDD.n178 185
R2180 VDD.n180 VDD.n179 185
R2181 VDD.n3833 VDD.n3832 185
R2182 VDD.n3834 VDD.n3833 185
R2183 VDD.n188 VDD.n187 185
R2184 VDD.n187 VDD.n186 185
R2185 VDD.n3828 VDD.n3827 185
R2186 VDD.n3827 VDD.n3826 185
R2187 VDD.n191 VDD.n190 185
R2188 VDD.n3817 VDD.n191 185
R2189 VDD.n3816 VDD.n3815 185
R2190 VDD.n3818 VDD.n3816 185
R2191 VDD.n199 VDD.n198 185
R2192 VDD.n198 VDD.n197 185
R2193 VDD.n3811 VDD.n3810 185
R2194 VDD.n3810 VDD.n3809 185
R2195 VDD.n202 VDD.n201 185
R2196 VDD.n203 VDD.n202 185
R2197 VDD.n3800 VDD.n3799 185
R2198 VDD.n3801 VDD.n3800 185
R2199 VDD.n211 VDD.n210 185
R2200 VDD.n210 VDD.n209 185
R2201 VDD.n3795 VDD.n3794 185
R2202 VDD.n3794 VDD.n3793 185
R2203 VDD.n214 VDD.n213 185
R2204 VDD.n215 VDD.n214 185
R2205 VDD.n3784 VDD.n3783 185
R2206 VDD.n3785 VDD.n3784 185
R2207 VDD.n223 VDD.n222 185
R2208 VDD.n222 VDD.n221 185
R2209 VDD.n3779 VDD.n3778 185
R2210 VDD.n3778 VDD.t81 185
R2211 VDD.n226 VDD.n225 185
R2212 VDD.n227 VDD.n226 185
R2213 VDD.n3769 VDD.n3768 185
R2214 VDD.n3770 VDD.n3769 185
R2215 VDD.n235 VDD.n234 185
R2216 VDD.n234 VDD.n233 185
R2217 VDD.n3764 VDD.n3763 185
R2218 VDD.n3763 VDD.n3762 185
R2219 VDD.n238 VDD.n237 185
R2220 VDD.n239 VDD.n238 185
R2221 VDD.n3753 VDD.n3752 185
R2222 VDD.n3754 VDD.n3753 185
R2223 VDD.n247 VDD.n246 185
R2224 VDD.n246 VDD.n245 185
R2225 VDD.n3748 VDD.n3747 185
R2226 VDD.n3747 VDD.n3746 185
R2227 VDD.n250 VDD.n249 185
R2228 VDD.n251 VDD.n250 185
R2229 VDD.n3737 VDD.n3736 185
R2230 VDD.n3738 VDD.n3737 185
R2231 VDD.n259 VDD.n258 185
R2232 VDD.n258 VDD.n257 185
R2233 VDD.n3732 VDD.n3731 185
R2234 VDD.n3731 VDD.n3730 185
R2235 VDD.n262 VDD.n261 185
R2236 VDD.n263 VDD.n262 185
R2237 VDD.n3721 VDD.n3720 185
R2238 VDD.n3722 VDD.n3721 185
R2239 VDD.n270 VDD.n269 185
R2240 VDD.n275 VDD.n269 185
R2241 VDD.n3716 VDD.n3715 185
R2242 VDD.n3715 VDD.n3714 185
R2243 VDD.n273 VDD.n272 185
R2244 VDD.n274 VDD.n273 185
R2245 VDD.n3705 VDD.n3704 185
R2246 VDD.n3706 VDD.n3705 185
R2247 VDD.n283 VDD.n282 185
R2248 VDD.n282 VDD.n281 185
R2249 VDD.n3700 VDD.n3699 185
R2250 VDD.n3699 VDD.n3698 185
R2251 VDD.n286 VDD.n285 185
R2252 VDD.n287 VDD.n286 185
R2253 VDD.n3172 VDD.n3171 185
R2254 VDD.n3170 VDD.n2809 185
R2255 VDD.n3169 VDD.n2808 185
R2256 VDD.n3174 VDD.n2808 185
R2257 VDD.n3168 VDD.n3167 185
R2258 VDD.n3166 VDD.n3165 185
R2259 VDD.n3164 VDD.n3163 185
R2260 VDD.n3162 VDD.n3161 185
R2261 VDD.n3160 VDD.n3159 185
R2262 VDD.n3158 VDD.n3157 185
R2263 VDD.n3156 VDD.n3155 185
R2264 VDD.n3154 VDD.n3153 185
R2265 VDD.n3152 VDD.n3151 185
R2266 VDD.n3150 VDD.n3149 185
R2267 VDD.n3148 VDD.n3147 185
R2268 VDD.n3146 VDD.n3145 185
R2269 VDD.n3144 VDD.n3143 185
R2270 VDD.n3142 VDD.n3141 185
R2271 VDD.n3140 VDD.n3139 185
R2272 VDD.n3138 VDD.n3137 185
R2273 VDD.n3136 VDD.n3135 185
R2274 VDD.n3134 VDD.n3133 185
R2275 VDD.n3132 VDD.n3131 185
R2276 VDD.n3130 VDD.n3129 185
R2277 VDD.n3128 VDD.n3127 185
R2278 VDD.n3126 VDD.n3125 185
R2279 VDD.n3479 VDD.n3478 185
R2280 VDD.n3480 VDD.n361 185
R2281 VDD.n3482 VDD.n3481 185
R2282 VDD.n3484 VDD.n360 185
R2283 VDD.n3486 VDD.n3485 185
R2284 VDD.n3487 VDD.n355 185
R2285 VDD.n3489 VDD.n3488 185
R2286 VDD.n3491 VDD.n353 185
R2287 VDD.n3493 VDD.n3492 185
R2288 VDD.n3494 VDD.n352 185
R2289 VDD.n3496 VDD.n3495 185
R2290 VDD.n3498 VDD.n351 185
R2291 VDD.n3499 VDD.n290 185
R2292 VDD.n3501 VDD.n349 185
R2293 VDD.n3503 VDD.n3502 185
R2294 VDD.n3504 VDD.n348 185
R2295 VDD.n3506 VDD.n3505 185
R2296 VDD.n3508 VDD.n346 185
R2297 VDD.n3510 VDD.n3509 185
R2298 VDD.n3511 VDD.n345 185
R2299 VDD.n3513 VDD.n3512 185
R2300 VDD.n3515 VDD.n344 185
R2301 VDD.n3516 VDD.n343 185
R2302 VDD.n3519 VDD.n3518 185
R2303 VDD.n3520 VDD.n341 185
R2304 VDD.n341 VDD.n323 185
R2305 VDD.n3476 VDD.n338 185
R2306 VDD.n3523 VDD.n338 185
R2307 VDD.n3475 VDD.n3474 185
R2308 VDD.n3474 VDD.n337 185
R2309 VDD.n3473 VDD.n362 185
R2310 VDD.n3473 VDD.n3472 185
R2311 VDD.n2813 VDD.n363 185
R2312 VDD.n364 VDD.n363 185
R2313 VDD.n2814 VDD.n371 185
R2314 VDD.n3466 VDD.n371 185
R2315 VDD.n2816 VDD.n2815 185
R2316 VDD.n2815 VDD.n370 185
R2317 VDD.n2817 VDD.n378 185
R2318 VDD.n3427 VDD.n378 185
R2319 VDD.n2819 VDD.n2818 185
R2320 VDD.n2818 VDD.n377 185
R2321 VDD.n2820 VDD.n383 185
R2322 VDD.n3421 VDD.n383 185
R2323 VDD.n2822 VDD.n2821 185
R2324 VDD.n2821 VDD.n391 185
R2325 VDD.n2823 VDD.n389 185
R2326 VDD.n3415 VDD.n389 185
R2327 VDD.n2825 VDD.n2824 185
R2328 VDD.n2824 VDD.n388 185
R2329 VDD.n2826 VDD.n396 185
R2330 VDD.n3409 VDD.n396 185
R2331 VDD.n2828 VDD.n2827 185
R2332 VDD.n2827 VDD.n395 185
R2333 VDD.n2829 VDD.n402 185
R2334 VDD.n3403 VDD.n402 185
R2335 VDD.n2831 VDD.n2830 185
R2336 VDD.n2830 VDD.n401 185
R2337 VDD.n2832 VDD.n408 185
R2338 VDD.n3397 VDD.n408 185
R2339 VDD.n2834 VDD.n2833 185
R2340 VDD.n2833 VDD.n407 185
R2341 VDD.n2835 VDD.n414 185
R2342 VDD.n3391 VDD.n414 185
R2343 VDD.n2837 VDD.n2836 185
R2344 VDD.n2836 VDD.n413 185
R2345 VDD.n2838 VDD.n420 185
R2346 VDD.n3385 VDD.n420 185
R2347 VDD.n2840 VDD.n2839 185
R2348 VDD.n2839 VDD.n419 185
R2349 VDD.n2841 VDD.n426 185
R2350 VDD.n3379 VDD.n426 185
R2351 VDD.n2843 VDD.n2842 185
R2352 VDD.n2842 VDD.n425 185
R2353 VDD.n2844 VDD.n431 185
R2354 VDD.n3373 VDD.n431 185
R2355 VDD.n3028 VDD.n3027 185
R2356 VDD.n3027 VDD.n3026 185
R2357 VDD.n3029 VDD.n437 185
R2358 VDD.n3367 VDD.n437 185
R2359 VDD.n3031 VDD.n3030 185
R2360 VDD.n3030 VDD.n436 185
R2361 VDD.n3032 VDD.n443 185
R2362 VDD.n3361 VDD.n443 185
R2363 VDD.n3034 VDD.n3033 185
R2364 VDD.n3033 VDD.n442 185
R2365 VDD.n3035 VDD.n449 185
R2366 VDD.n3355 VDD.n449 185
R2367 VDD.n3037 VDD.n3036 185
R2368 VDD.n3036 VDD.n448 185
R2369 VDD.n3038 VDD.n455 185
R2370 VDD.n3349 VDD.n455 185
R2371 VDD.n3040 VDD.n3039 185
R2372 VDD.n3039 VDD.n454 185
R2373 VDD.n3041 VDD.n461 185
R2374 VDD.n3343 VDD.n461 185
R2375 VDD.n3043 VDD.n3042 185
R2376 VDD.n3042 VDD.n460 185
R2377 VDD.n3044 VDD.n467 185
R2378 VDD.n3337 VDD.n467 185
R2379 VDD.n3046 VDD.n3045 185
R2380 VDD.n3045 VDD.n466 185
R2381 VDD.n3047 VDD.n472 185
R2382 VDD.n3331 VDD.n472 185
R2383 VDD.n3049 VDD.n3048 185
R2384 VDD.n3048 VDD.n480 185
R2385 VDD.n3050 VDD.n478 185
R2386 VDD.n3325 VDD.n478 185
R2387 VDD.n3052 VDD.n3051 185
R2388 VDD.n3051 VDD.n477 185
R2389 VDD.n3053 VDD.n485 185
R2390 VDD.n3319 VDD.n485 185
R2391 VDD.n3055 VDD.n3054 185
R2392 VDD.n3054 VDD.n484 185
R2393 VDD.n3056 VDD.n491 185
R2394 VDD.n3313 VDD.n491 185
R2395 VDD.n3058 VDD.n3057 185
R2396 VDD.n3057 VDD.n490 185
R2397 VDD.n3059 VDD.n497 185
R2398 VDD.n3307 VDD.n497 185
R2399 VDD.n3061 VDD.n3060 185
R2400 VDD.n3060 VDD.n496 185
R2401 VDD.n3062 VDD.n503 185
R2402 VDD.n3301 VDD.n503 185
R2403 VDD.n3064 VDD.n3063 185
R2404 VDD.n3063 VDD.n502 185
R2405 VDD.n3065 VDD.n508 185
R2406 VDD.n3295 VDD.n508 185
R2407 VDD.n3067 VDD.n3066 185
R2408 VDD.n3066 VDD.n516 185
R2409 VDD.n3068 VDD.n514 185
R2410 VDD.n3289 VDD.n514 185
R2411 VDD.n3070 VDD.n3069 185
R2412 VDD.n3069 VDD.n513 185
R2413 VDD.n3071 VDD.n521 185
R2414 VDD.n3283 VDD.n521 185
R2415 VDD.n3073 VDD.n3072 185
R2416 VDD.n3072 VDD.n520 185
R2417 VDD.n3074 VDD.n526 185
R2418 VDD.n3277 VDD.n526 185
R2419 VDD.n3076 VDD.n3075 185
R2420 VDD.n3075 VDD.n534 185
R2421 VDD.n3077 VDD.n532 185
R2422 VDD.n3271 VDD.n532 185
R2423 VDD.n3079 VDD.n3078 185
R2424 VDD.n3078 VDD.n531 185
R2425 VDD.n3080 VDD.n539 185
R2426 VDD.n3265 VDD.n539 185
R2427 VDD.n3082 VDD.n3081 185
R2428 VDD.n3081 VDD.n538 185
R2429 VDD.n3083 VDD.n545 185
R2430 VDD.n3259 VDD.n545 185
R2431 VDD.n3085 VDD.n3084 185
R2432 VDD.n3084 VDD.n544 185
R2433 VDD.n3086 VDD.n551 185
R2434 VDD.n3253 VDD.n551 185
R2435 VDD.n3088 VDD.n3087 185
R2436 VDD.n3087 VDD.n550 185
R2437 VDD.n3089 VDD.n557 185
R2438 VDD.n3247 VDD.n557 185
R2439 VDD.n3091 VDD.n3090 185
R2440 VDD.n3090 VDD.n556 185
R2441 VDD.n3092 VDD.n563 185
R2442 VDD.n3241 VDD.n563 185
R2443 VDD.n3094 VDD.n3093 185
R2444 VDD.n3093 VDD.n562 185
R2445 VDD.n3095 VDD.n569 185
R2446 VDD.n3235 VDD.n569 185
R2447 VDD.n3097 VDD.n3096 185
R2448 VDD.n3096 VDD.n568 185
R2449 VDD.n3098 VDD.n575 185
R2450 VDD.n3229 VDD.n575 185
R2451 VDD.n3100 VDD.n3099 185
R2452 VDD.n3099 VDD.n574 185
R2453 VDD.n3101 VDD.n581 185
R2454 VDD.n3223 VDD.n581 185
R2455 VDD.n3103 VDD.n3102 185
R2456 VDD.n3102 VDD.n580 185
R2457 VDD.n3104 VDD.n587 185
R2458 VDD.n3217 VDD.n587 185
R2459 VDD.n3106 VDD.n3105 185
R2460 VDD.n3105 VDD.n586 185
R2461 VDD.n3107 VDD.n593 185
R2462 VDD.n3211 VDD.n593 185
R2463 VDD.n3109 VDD.n3108 185
R2464 VDD.n3108 VDD.n592 185
R2465 VDD.n3110 VDD.n598 185
R2466 VDD.n3205 VDD.n598 185
R2467 VDD.n3112 VDD.n3111 185
R2468 VDD.n3111 VDD.n605 185
R2469 VDD.n3113 VDD.n603 185
R2470 VDD.n3199 VDD.n603 185
R2471 VDD.n3115 VDD.n3114 185
R2472 VDD.n3114 VDD.n612 185
R2473 VDD.n3116 VDD.n610 185
R2474 VDD.n3193 VDD.n610 185
R2475 VDD.n3118 VDD.n3117 185
R2476 VDD.n3117 VDD.n609 185
R2477 VDD.n3119 VDD.n617 185
R2478 VDD.n3187 VDD.n617 185
R2479 VDD.n3121 VDD.n3120 185
R2480 VDD.n3120 VDD.n616 185
R2481 VDD.n3122 VDD.n623 185
R2482 VDD.n3181 VDD.n623 185
R2483 VDD.n3124 VDD.n3123 185
R2484 VDD.n3124 VDD.n622 185
R2485 VDD.n621 VDD.n620 185
R2486 VDD.n622 VDD.n621 185
R2487 VDD.n3183 VDD.n3182 185
R2488 VDD.n3182 VDD.n3181 185
R2489 VDD.n3184 VDD.n619 185
R2490 VDD.n619 VDD.n616 185
R2491 VDD.n3186 VDD.n3185 185
R2492 VDD.n3187 VDD.n3186 185
R2493 VDD.n608 VDD.n607 185
R2494 VDD.n609 VDD.n608 185
R2495 VDD.n3195 VDD.n3194 185
R2496 VDD.n3194 VDD.n3193 185
R2497 VDD.n3196 VDD.n606 185
R2498 VDD.n612 VDD.n606 185
R2499 VDD.n3198 VDD.n3197 185
R2500 VDD.n3199 VDD.n3198 185
R2501 VDD.n597 VDD.n596 185
R2502 VDD.n605 VDD.n597 185
R2503 VDD.n3207 VDD.n3206 185
R2504 VDD.n3206 VDD.n3205 185
R2505 VDD.n3208 VDD.n595 185
R2506 VDD.n595 VDD.n592 185
R2507 VDD.n3210 VDD.n3209 185
R2508 VDD.n3211 VDD.n3210 185
R2509 VDD.n585 VDD.n584 185
R2510 VDD.n586 VDD.n585 185
R2511 VDD.n3219 VDD.n3218 185
R2512 VDD.n3218 VDD.n3217 185
R2513 VDD.n3220 VDD.n583 185
R2514 VDD.n583 VDD.n580 185
R2515 VDD.n3222 VDD.n3221 185
R2516 VDD.n3223 VDD.n3222 185
R2517 VDD.n573 VDD.n572 185
R2518 VDD.n574 VDD.n573 185
R2519 VDD.n3231 VDD.n3230 185
R2520 VDD.n3230 VDD.n3229 185
R2521 VDD.n3232 VDD.n571 185
R2522 VDD.n571 VDD.n568 185
R2523 VDD.n3234 VDD.n3233 185
R2524 VDD.n3235 VDD.n3234 185
R2525 VDD.n561 VDD.n560 185
R2526 VDD.n562 VDD.n561 185
R2527 VDD.n3243 VDD.n3242 185
R2528 VDD.n3242 VDD.n3241 185
R2529 VDD.n3244 VDD.n559 185
R2530 VDD.n559 VDD.n556 185
R2531 VDD.n3246 VDD.n3245 185
R2532 VDD.n3247 VDD.n3246 185
R2533 VDD.n549 VDD.n548 185
R2534 VDD.n550 VDD.n549 185
R2535 VDD.n3255 VDD.n3254 185
R2536 VDD.n3254 VDD.n3253 185
R2537 VDD.n3256 VDD.n547 185
R2538 VDD.n547 VDD.n544 185
R2539 VDD.n3258 VDD.n3257 185
R2540 VDD.n3259 VDD.n3258 185
R2541 VDD.n537 VDD.n536 185
R2542 VDD.n538 VDD.n537 185
R2543 VDD.n3267 VDD.n3266 185
R2544 VDD.n3266 VDD.n3265 185
R2545 VDD.n3268 VDD.n535 185
R2546 VDD.n535 VDD.n531 185
R2547 VDD.n3270 VDD.n3269 185
R2548 VDD.n3271 VDD.n3270 185
R2549 VDD.n525 VDD.n524 185
R2550 VDD.n534 VDD.n525 185
R2551 VDD.n3279 VDD.n3278 185
R2552 VDD.n3278 VDD.n3277 185
R2553 VDD.n3280 VDD.n523 185
R2554 VDD.n523 VDD.n520 185
R2555 VDD.n3282 VDD.n3281 185
R2556 VDD.n3283 VDD.n3282 185
R2557 VDD.n512 VDD.n511 185
R2558 VDD.n513 VDD.n512 185
R2559 VDD.n3291 VDD.n3290 185
R2560 VDD.n3290 VDD.n3289 185
R2561 VDD.n3292 VDD.n510 185
R2562 VDD.n516 VDD.n510 185
R2563 VDD.n3294 VDD.n3293 185
R2564 VDD.n3295 VDD.n3294 185
R2565 VDD.n501 VDD.n500 185
R2566 VDD.n502 VDD.n501 185
R2567 VDD.n3303 VDD.n3302 185
R2568 VDD.n3302 VDD.n3301 185
R2569 VDD.n3304 VDD.n499 185
R2570 VDD.n499 VDD.n496 185
R2571 VDD.n3306 VDD.n3305 185
R2572 VDD.n3307 VDD.n3306 185
R2573 VDD.n489 VDD.n488 185
R2574 VDD.n490 VDD.n489 185
R2575 VDD.n3315 VDD.n3314 185
R2576 VDD.n3314 VDD.n3313 185
R2577 VDD.n3316 VDD.n487 185
R2578 VDD.n487 VDD.n484 185
R2579 VDD.n3318 VDD.n3317 185
R2580 VDD.n3319 VDD.n3318 185
R2581 VDD.n476 VDD.n475 185
R2582 VDD.n477 VDD.n476 185
R2583 VDD.n3327 VDD.n3326 185
R2584 VDD.n3326 VDD.n3325 185
R2585 VDD.n3328 VDD.n474 185
R2586 VDD.n480 VDD.n474 185
R2587 VDD.n3330 VDD.n3329 185
R2588 VDD.n3331 VDD.n3330 185
R2589 VDD.n465 VDD.n464 185
R2590 VDD.n466 VDD.n465 185
R2591 VDD.n3339 VDD.n3338 185
R2592 VDD.n3338 VDD.n3337 185
R2593 VDD.n3340 VDD.n463 185
R2594 VDD.n463 VDD.n460 185
R2595 VDD.n3342 VDD.n3341 185
R2596 VDD.n3343 VDD.n3342 185
R2597 VDD.n453 VDD.n452 185
R2598 VDD.n454 VDD.n453 185
R2599 VDD.n3351 VDD.n3350 185
R2600 VDD.n3350 VDD.n3349 185
R2601 VDD.n3352 VDD.n451 185
R2602 VDD.n451 VDD.n448 185
R2603 VDD.n3354 VDD.n3353 185
R2604 VDD.n3355 VDD.n3354 185
R2605 VDD.n441 VDD.n440 185
R2606 VDD.n442 VDD.n441 185
R2607 VDD.n3363 VDD.n3362 185
R2608 VDD.n3362 VDD.n3361 185
R2609 VDD.n3364 VDD.n439 185
R2610 VDD.n439 VDD.n436 185
R2611 VDD.n3366 VDD.n3365 185
R2612 VDD.n3367 VDD.n3366 185
R2613 VDD.n430 VDD.n429 185
R2614 VDD.n3026 VDD.n430 185
R2615 VDD.n3375 VDD.n3374 185
R2616 VDD.n3374 VDD.n3373 185
R2617 VDD.n3376 VDD.n428 185
R2618 VDD.n428 VDD.n425 185
R2619 VDD.n3378 VDD.n3377 185
R2620 VDD.n3379 VDD.n3378 185
R2621 VDD.n418 VDD.n417 185
R2622 VDD.n419 VDD.n418 185
R2623 VDD.n3387 VDD.n3386 185
R2624 VDD.n3386 VDD.n3385 185
R2625 VDD.n3388 VDD.n416 185
R2626 VDD.n416 VDD.n413 185
R2627 VDD.n3390 VDD.n3389 185
R2628 VDD.n3391 VDD.n3390 185
R2629 VDD.n406 VDD.n405 185
R2630 VDD.n407 VDD.n406 185
R2631 VDD.n3399 VDD.n3398 185
R2632 VDD.n3398 VDD.n3397 185
R2633 VDD.n3400 VDD.n404 185
R2634 VDD.n404 VDD.n401 185
R2635 VDD.n3402 VDD.n3401 185
R2636 VDD.n3403 VDD.n3402 185
R2637 VDD.n394 VDD.n393 185
R2638 VDD.n395 VDD.n394 185
R2639 VDD.n3411 VDD.n3410 185
R2640 VDD.n3410 VDD.n3409 185
R2641 VDD.n3412 VDD.n392 185
R2642 VDD.n392 VDD.n388 185
R2643 VDD.n3414 VDD.n3413 185
R2644 VDD.n3415 VDD.n3414 185
R2645 VDD.n382 VDD.n381 185
R2646 VDD.n391 VDD.n382 185
R2647 VDD.n3423 VDD.n3422 185
R2648 VDD.n3422 VDD.n3421 185
R2649 VDD.n3424 VDD.n380 185
R2650 VDD.n380 VDD.n377 185
R2651 VDD.n3426 VDD.n3425 185
R2652 VDD.n3427 VDD.n3426 185
R2653 VDD.n369 VDD.n368 185
R2654 VDD.n370 VDD.n369 185
R2655 VDD.n3468 VDD.n3467 185
R2656 VDD.n3467 VDD.n3466 185
R2657 VDD.n3469 VDD.n367 185
R2658 VDD.n367 VDD.n364 185
R2659 VDD.n3471 VDD.n3470 185
R2660 VDD.n3472 VDD.n3471 185
R2661 VDD.n342 VDD.n340 185
R2662 VDD.n340 VDD.n337 185
R2663 VDD.n3522 VDD.n3521 185
R2664 VDD.n3523 VDD.n3522 185
R2665 VDD.n2721 VDD.n2720 185
R2666 VDD.n2720 VDD.n628 185
R2667 VDD.n2722 VDD.n665 185
R2668 VDD.n2732 VDD.n665 185
R2669 VDD.n2723 VDD.n673 185
R2670 VDD.n673 VDD.n663 185
R2671 VDD.n2725 VDD.n2724 185
R2672 VDD.n2726 VDD.n2725 185
R2673 VDD.n674 VDD.n672 185
R2674 VDD.n672 VDD.n669 185
R2675 VDD.n2650 VDD.n681 185
R2676 VDD.n2660 VDD.n681 185
R2677 VDD.n2651 VDD.n689 185
R2678 VDD.n689 VDD.n679 185
R2679 VDD.n2653 VDD.n2652 185
R2680 VDD.n2654 VDD.n2653 185
R2681 VDD.n2649 VDD.n688 185
R2682 VDD.n688 VDD.n685 185
R2683 VDD.n2648 VDD.n2647 185
R2684 VDD.n2647 VDD.n2646 185
R2685 VDD.n691 VDD.n690 185
R2686 VDD.n692 VDD.n691 185
R2687 VDD.n2639 VDD.n2638 185
R2688 VDD.n2640 VDD.n2639 185
R2689 VDD.n2637 VDD.n701 185
R2690 VDD.n701 VDD.n698 185
R2691 VDD.n2636 VDD.n2635 185
R2692 VDD.n2635 VDD.n2634 185
R2693 VDD.n703 VDD.n702 185
R2694 VDD.n704 VDD.n703 185
R2695 VDD.n2627 VDD.n2626 185
R2696 VDD.n2628 VDD.n2627 185
R2697 VDD.n2625 VDD.n713 185
R2698 VDD.n713 VDD.n710 185
R2699 VDD.n2624 VDD.n2623 185
R2700 VDD.n2623 VDD.n2622 185
R2701 VDD.n715 VDD.n714 185
R2702 VDD.n716 VDD.n715 185
R2703 VDD.n2615 VDD.n2614 185
R2704 VDD.n2616 VDD.n2615 185
R2705 VDD.n2613 VDD.n724 185
R2706 VDD.n730 VDD.n724 185
R2707 VDD.n2612 VDD.n2611 185
R2708 VDD.n2611 VDD.n2610 185
R2709 VDD.n726 VDD.n725 185
R2710 VDD.n727 VDD.n726 185
R2711 VDD.n2603 VDD.n2602 185
R2712 VDD.n2604 VDD.n2603 185
R2713 VDD.n2601 VDD.n737 185
R2714 VDD.n737 VDD.n734 185
R2715 VDD.n2600 VDD.n2599 185
R2716 VDD.n2599 VDD.n2598 185
R2717 VDD.n739 VDD.n738 185
R2718 VDD.n748 VDD.n739 185
R2719 VDD.n2591 VDD.n2590 185
R2720 VDD.n2592 VDD.n2591 185
R2721 VDD.n2589 VDD.n749 185
R2722 VDD.n749 VDD.n745 185
R2723 VDD.n2588 VDD.n2587 185
R2724 VDD.n2587 VDD.n2586 185
R2725 VDD.n751 VDD.n750 185
R2726 VDD.n752 VDD.n751 185
R2727 VDD.n2579 VDD.n2578 185
R2728 VDD.n2580 VDD.n2579 185
R2729 VDD.n2577 VDD.n761 185
R2730 VDD.n761 VDD.n758 185
R2731 VDD.n2576 VDD.n2575 185
R2732 VDD.n2575 VDD.n2574 185
R2733 VDD.n763 VDD.n762 185
R2734 VDD.n764 VDD.n763 185
R2735 VDD.n2567 VDD.n2566 185
R2736 VDD.n2568 VDD.n2567 185
R2737 VDD.n2565 VDD.n773 185
R2738 VDD.n773 VDD.n770 185
R2739 VDD.n2564 VDD.n2563 185
R2740 VDD.n2563 VDD.n2562 185
R2741 VDD.n775 VDD.n774 185
R2742 VDD.n776 VDD.n775 185
R2743 VDD.n2555 VDD.n2554 185
R2744 VDD.n2556 VDD.n2555 185
R2745 VDD.n2553 VDD.n785 185
R2746 VDD.n785 VDD.n782 185
R2747 VDD.n2552 VDD.n2551 185
R2748 VDD.n2551 VDD.n2550 185
R2749 VDD.n787 VDD.n786 185
R2750 VDD.n788 VDD.n787 185
R2751 VDD.n2543 VDD.n2542 185
R2752 VDD.n2544 VDD.n2543 185
R2753 VDD.n2541 VDD.n797 185
R2754 VDD.n797 VDD.n794 185
R2755 VDD.n2540 VDD.n2539 185
R2756 VDD.n2539 VDD.n2538 185
R2757 VDD.n799 VDD.n798 185
R2758 VDD.n808 VDD.n799 185
R2759 VDD.n2531 VDD.n2530 185
R2760 VDD.n2532 VDD.n2531 185
R2761 VDD.n2529 VDD.n809 185
R2762 VDD.n809 VDD.n805 185
R2763 VDD.n2528 VDD.n2527 185
R2764 VDD.n2527 VDD.n2526 185
R2765 VDD.n811 VDD.n810 185
R2766 VDD.n812 VDD.n811 185
R2767 VDD.n2519 VDD.n2518 185
R2768 VDD.n2520 VDD.n2519 185
R2769 VDD.n2517 VDD.n821 185
R2770 VDD.n821 VDD.n818 185
R2771 VDD.n2516 VDD.n2515 185
R2772 VDD.n2515 VDD.n2514 185
R2773 VDD.n823 VDD.n822 185
R2774 VDD.n824 VDD.n823 185
R2775 VDD.n2507 VDD.n2506 185
R2776 VDD.n2508 VDD.n2507 185
R2777 VDD.n2505 VDD.n833 185
R2778 VDD.n833 VDD.n830 185
R2779 VDD.n2504 VDD.n2503 185
R2780 VDD.n2503 VDD.n2502 185
R2781 VDD.n835 VDD.n834 185
R2782 VDD.n836 VDD.n835 185
R2783 VDD.n2495 VDD.n2494 185
R2784 VDD.n2496 VDD.n2495 185
R2785 VDD.n2493 VDD.n845 185
R2786 VDD.n845 VDD.n842 185
R2787 VDD.n2492 VDD.n2491 185
R2788 VDD.n2491 VDD.n2490 185
R2789 VDD.n847 VDD.n846 185
R2790 VDD.n848 VDD.n847 185
R2791 VDD.n2483 VDD.n2482 185
R2792 VDD.n2484 VDD.n2483 185
R2793 VDD.n2481 VDD.n856 185
R2794 VDD.n2357 VDD.n856 185
R2795 VDD.n2480 VDD.n2479 185
R2796 VDD.n2479 VDD.n2478 185
R2797 VDD.n858 VDD.n857 185
R2798 VDD.n859 VDD.n858 185
R2799 VDD.n2471 VDD.n2470 185
R2800 VDD.n2472 VDD.n2471 185
R2801 VDD.n2469 VDD.n868 185
R2802 VDD.n868 VDD.n865 185
R2803 VDD.n2468 VDD.n2467 185
R2804 VDD.n2467 VDD.n2466 185
R2805 VDD.n870 VDD.n869 185
R2806 VDD.n871 VDD.n870 185
R2807 VDD.n2459 VDD.n2458 185
R2808 VDD.n2460 VDD.n2459 185
R2809 VDD.n2457 VDD.n880 185
R2810 VDD.n880 VDD.n877 185
R2811 VDD.n2456 VDD.n2455 185
R2812 VDD.n2455 VDD.n2454 185
R2813 VDD.n882 VDD.n881 185
R2814 VDD.n883 VDD.n882 185
R2815 VDD.n2447 VDD.n2446 185
R2816 VDD.n2448 VDD.n2447 185
R2817 VDD.n2445 VDD.n892 185
R2818 VDD.n892 VDD.n889 185
R2819 VDD.n2444 VDD.n2443 185
R2820 VDD.n2443 VDD.n2442 185
R2821 VDD.n894 VDD.n893 185
R2822 VDD.n903 VDD.n894 185
R2823 VDD.n2435 VDD.n2434 185
R2824 VDD.n2436 VDD.n2435 185
R2825 VDD.n2433 VDD.n904 185
R2826 VDD.n904 VDD.n900 185
R2827 VDD.n2432 VDD.n2431 185
R2828 VDD.n2431 VDD.n2430 185
R2829 VDD.n906 VDD.n905 185
R2830 VDD.n907 VDD.n906 185
R2831 VDD.n2423 VDD.n2422 185
R2832 VDD.n2424 VDD.n2423 185
R2833 VDD.n2421 VDD.n916 185
R2834 VDD.n916 VDD.n913 185
R2835 VDD.n2420 VDD.n2419 185
R2836 VDD.n2419 VDD.n2418 185
R2837 VDD.n918 VDD.n917 185
R2838 VDD.n919 VDD.n918 185
R2839 VDD.n2411 VDD.n2410 185
R2840 VDD.n2412 VDD.n2411 185
R2841 VDD.n2409 VDD.n928 185
R2842 VDD.n928 VDD.n925 185
R2843 VDD.n2408 VDD.n2407 185
R2844 VDD.n2407 VDD.n2406 185
R2845 VDD.n2670 VDD.n641 185
R2846 VDD.n2784 VDD.n641 185
R2847 VDD.n2672 VDD.n2671 185
R2848 VDD.n2674 VDD.n2673 185
R2849 VDD.n2676 VDD.n2675 185
R2850 VDD.n2679 VDD.n2678 185
R2851 VDD.n2681 VDD.n2680 185
R2852 VDD.n2683 VDD.n2682 185
R2853 VDD.n2685 VDD.n2684 185
R2854 VDD.n2687 VDD.n2686 185
R2855 VDD.n2689 VDD.n2688 185
R2856 VDD.n2691 VDD.n2690 185
R2857 VDD.n2693 VDD.n2692 185
R2858 VDD.n2695 VDD.n2694 185
R2859 VDD.n2697 VDD.n2696 185
R2860 VDD.n2699 VDD.n2698 185
R2861 VDD.n2701 VDD.n2700 185
R2862 VDD.n2703 VDD.n2702 185
R2863 VDD.n2705 VDD.n2704 185
R2864 VDD.n2707 VDD.n2706 185
R2865 VDD.n2709 VDD.n2708 185
R2866 VDD.n2711 VDD.n2710 185
R2867 VDD.n2713 VDD.n2712 185
R2868 VDD.n2715 VDD.n2714 185
R2869 VDD.n2717 VDD.n2716 185
R2870 VDD.n2719 VDD.n2718 185
R2871 VDD.n2669 VDD.n2668 185
R2872 VDD.n2668 VDD.n628 185
R2873 VDD.n2667 VDD.n664 185
R2874 VDD.n2732 VDD.n664 185
R2875 VDD.n2666 VDD.n2665 185
R2876 VDD.n2665 VDD.n663 185
R2877 VDD.n2664 VDD.n671 185
R2878 VDD.n2726 VDD.n671 185
R2879 VDD.n2663 VDD.n2662 185
R2880 VDD.n2662 VDD.n669 185
R2881 VDD.n2661 VDD.n677 185
R2882 VDD.n2661 VDD.n2660 185
R2883 VDD.n961 VDD.n678 185
R2884 VDD.n679 VDD.n678 185
R2885 VDD.n962 VDD.n687 185
R2886 VDD.n2654 VDD.n687 185
R2887 VDD.n964 VDD.n963 185
R2888 VDD.n963 VDD.n685 185
R2889 VDD.n965 VDD.n694 185
R2890 VDD.n2646 VDD.n694 185
R2891 VDD.n967 VDD.n966 185
R2892 VDD.n966 VDD.n692 185
R2893 VDD.n968 VDD.n700 185
R2894 VDD.n2640 VDD.n700 185
R2895 VDD.n970 VDD.n969 185
R2896 VDD.n969 VDD.n698 185
R2897 VDD.n971 VDD.n706 185
R2898 VDD.n2634 VDD.n706 185
R2899 VDD.n973 VDD.n972 185
R2900 VDD.n972 VDD.n704 185
R2901 VDD.n974 VDD.n712 185
R2902 VDD.n2628 VDD.n712 185
R2903 VDD.n976 VDD.n975 185
R2904 VDD.n975 VDD.n710 185
R2905 VDD.n977 VDD.n718 185
R2906 VDD.n2622 VDD.n718 185
R2907 VDD.n979 VDD.n978 185
R2908 VDD.n978 VDD.n716 185
R2909 VDD.n980 VDD.n723 185
R2910 VDD.n2616 VDD.n723 185
R2911 VDD.n982 VDD.n981 185
R2912 VDD.n981 VDD.n730 185
R2913 VDD.n983 VDD.n729 185
R2914 VDD.n2610 VDD.n729 185
R2915 VDD.n985 VDD.n984 185
R2916 VDD.n984 VDD.n727 185
R2917 VDD.n986 VDD.n736 185
R2918 VDD.n2604 VDD.n736 185
R2919 VDD.n988 VDD.n987 185
R2920 VDD.n987 VDD.n734 185
R2921 VDD.n989 VDD.n741 185
R2922 VDD.n2598 VDD.n741 185
R2923 VDD.n991 VDD.n990 185
R2924 VDD.n990 VDD.n748 185
R2925 VDD.n992 VDD.n747 185
R2926 VDD.n2592 VDD.n747 185
R2927 VDD.n994 VDD.n993 185
R2928 VDD.n993 VDD.n745 185
R2929 VDD.n995 VDD.n754 185
R2930 VDD.n2586 VDD.n754 185
R2931 VDD.n997 VDD.n996 185
R2932 VDD.n996 VDD.n752 185
R2933 VDD.n998 VDD.n760 185
R2934 VDD.n2580 VDD.n760 185
R2935 VDD.n1000 VDD.n999 185
R2936 VDD.n999 VDD.n758 185
R2937 VDD.n1001 VDD.n766 185
R2938 VDD.n2574 VDD.n766 185
R2939 VDD.n1003 VDD.n1002 185
R2940 VDD.n1002 VDD.n764 185
R2941 VDD.n1004 VDD.n772 185
R2942 VDD.n2568 VDD.n772 185
R2943 VDD.n1006 VDD.n1005 185
R2944 VDD.n1005 VDD.n770 185
R2945 VDD.n1007 VDD.n778 185
R2946 VDD.n2562 VDD.n778 185
R2947 VDD.n1009 VDD.n1008 185
R2948 VDD.n1008 VDD.n776 185
R2949 VDD.n1010 VDD.n784 185
R2950 VDD.n2556 VDD.n784 185
R2951 VDD.n1012 VDD.n1011 185
R2952 VDD.n1011 VDD.n782 185
R2953 VDD.n1013 VDD.n790 185
R2954 VDD.n2550 VDD.n790 185
R2955 VDD.n1015 VDD.n1014 185
R2956 VDD.n1014 VDD.n788 185
R2957 VDD.n1016 VDD.n796 185
R2958 VDD.n2544 VDD.n796 185
R2959 VDD.n1018 VDD.n1017 185
R2960 VDD.n1017 VDD.n794 185
R2961 VDD.n1019 VDD.n801 185
R2962 VDD.n2538 VDD.n801 185
R2963 VDD.n1021 VDD.n1020 185
R2964 VDD.n1020 VDD.n808 185
R2965 VDD.n1022 VDD.n807 185
R2966 VDD.n2532 VDD.n807 185
R2967 VDD.n1024 VDD.n1023 185
R2968 VDD.n1023 VDD.n805 185
R2969 VDD.n1025 VDD.n814 185
R2970 VDD.n2526 VDD.n814 185
R2971 VDD.n1027 VDD.n1026 185
R2972 VDD.n1026 VDD.n812 185
R2973 VDD.n1028 VDD.n820 185
R2974 VDD.n2520 VDD.n820 185
R2975 VDD.n1030 VDD.n1029 185
R2976 VDD.n1029 VDD.n818 185
R2977 VDD.n1031 VDD.n826 185
R2978 VDD.n2514 VDD.n826 185
R2979 VDD.n1033 VDD.n1032 185
R2980 VDD.n1032 VDD.n824 185
R2981 VDD.n1034 VDD.n832 185
R2982 VDD.n2508 VDD.n832 185
R2983 VDD.n1036 VDD.n1035 185
R2984 VDD.n1035 VDD.n830 185
R2985 VDD.n1037 VDD.n838 185
R2986 VDD.n2502 VDD.n838 185
R2987 VDD.n1039 VDD.n1038 185
R2988 VDD.n1038 VDD.n836 185
R2989 VDD.n1040 VDD.n844 185
R2990 VDD.n2496 VDD.n844 185
R2991 VDD.n1042 VDD.n1041 185
R2992 VDD.n1041 VDD.n842 185
R2993 VDD.n1043 VDD.n850 185
R2994 VDD.n2490 VDD.n850 185
R2995 VDD.n1045 VDD.n1044 185
R2996 VDD.n1044 VDD.n848 185
R2997 VDD.n1046 VDD.n855 185
R2998 VDD.n2484 VDD.n855 185
R2999 VDD.n2359 VDD.n2358 185
R3000 VDD.n2358 VDD.n2357 185
R3001 VDD.n2360 VDD.n861 185
R3002 VDD.n2478 VDD.n861 185
R3003 VDD.n2362 VDD.n2361 185
R3004 VDD.n2361 VDD.n859 185
R3005 VDD.n2363 VDD.n867 185
R3006 VDD.n2472 VDD.n867 185
R3007 VDD.n2365 VDD.n2364 185
R3008 VDD.n2364 VDD.n865 185
R3009 VDD.n2366 VDD.n873 185
R3010 VDD.n2466 VDD.n873 185
R3011 VDD.n2368 VDD.n2367 185
R3012 VDD.n2367 VDD.n871 185
R3013 VDD.n2369 VDD.n879 185
R3014 VDD.n2460 VDD.n879 185
R3015 VDD.n2371 VDD.n2370 185
R3016 VDD.n2370 VDD.n877 185
R3017 VDD.n2372 VDD.n885 185
R3018 VDD.n2454 VDD.n885 185
R3019 VDD.n2374 VDD.n2373 185
R3020 VDD.n2373 VDD.n883 185
R3021 VDD.n2375 VDD.n891 185
R3022 VDD.n2448 VDD.n891 185
R3023 VDD.n2377 VDD.n2376 185
R3024 VDD.n2376 VDD.n889 185
R3025 VDD.n2378 VDD.n896 185
R3026 VDD.n2442 VDD.n896 185
R3027 VDD.n2380 VDD.n2379 185
R3028 VDD.n2379 VDD.n903 185
R3029 VDD.n2381 VDD.n902 185
R3030 VDD.n2436 VDD.n902 185
R3031 VDD.n2383 VDD.n2382 185
R3032 VDD.n2382 VDD.n900 185
R3033 VDD.n2384 VDD.n909 185
R3034 VDD.n2430 VDD.n909 185
R3035 VDD.n2386 VDD.n2385 185
R3036 VDD.n2385 VDD.n907 185
R3037 VDD.n2387 VDD.n915 185
R3038 VDD.n2424 VDD.n915 185
R3039 VDD.n2389 VDD.n2388 185
R3040 VDD.n2388 VDD.n913 185
R3041 VDD.n2390 VDD.n921 185
R3042 VDD.n2418 VDD.n921 185
R3043 VDD.n2392 VDD.n2391 185
R3044 VDD.n2391 VDD.n919 185
R3045 VDD.n2393 VDD.n927 185
R3046 VDD.n2412 VDD.n927 185
R3047 VDD.n2395 VDD.n2394 185
R3048 VDD.n2394 VDD.n925 185
R3049 VDD.n2396 VDD.n932 185
R3050 VDD.n2406 VDD.n932 185
R3051 VDD.n930 VDD.n929 185
R3052 VDD.n1148 VDD.n1147 185
R3053 VDD.n1150 VDD.n1149 185
R3054 VDD.n1152 VDD.n1151 185
R3055 VDD.n1154 VDD.n1153 185
R3056 VDD.n1156 VDD.n1155 185
R3057 VDD.n1158 VDD.n1157 185
R3058 VDD.n1160 VDD.n1159 185
R3059 VDD.n1162 VDD.n1161 185
R3060 VDD.n1164 VDD.n1163 185
R3061 VDD.n1166 VDD.n1165 185
R3062 VDD.n1168 VDD.n1167 185
R3063 VDD.n1193 VDD.n1169 185
R3064 VDD.n1192 VDD.n1191 185
R3065 VDD.n1190 VDD.n1189 185
R3066 VDD.n1188 VDD.n1187 185
R3067 VDD.n1186 VDD.n1185 185
R3068 VDD.n1184 VDD.n1183 185
R3069 VDD.n1182 VDD.n1181 185
R3070 VDD.n1180 VDD.n1179 185
R3071 VDD.n1178 VDD.n1177 185
R3072 VDD.n1175 VDD.n1174 185
R3073 VDD.n1173 VDD.n1172 185
R3074 VDD.n960 VDD.n959 185
R3075 VDD.n2398 VDD.n2397 185
R3076 VDD.n2399 VDD.n2398 185
R3077 VDD.t1 VDD.t128 165.478
R3078 VDD.t144 VDD.t0 165.478
R3079 VDD.n1170 VDD.t56 165.321
R3080 VDD.n675 VDD.t32 165.321
R3081 VDD.n1047 VDD.t43 165.321
R3082 VDD.n657 VDD.t19 165.321
R3083 VDD.n2845 VDD.t50 165.321
R3084 VDD.n356 VDD.t62 165.321
R3085 VDD.n2810 VDD.t53 165.321
R3086 VDD.n328 VDD.t59 165.321
R3087 VDD.n4221 VDD.n4026 146.341
R3088 VDD.n4214 VDD.n4213 146.341
R3089 VDD.n4211 VDD.n4210 146.341
R3090 VDD.n4207 VDD.n4206 146.341
R3091 VDD.n4203 VDD.n4202 146.341
R3092 VDD.n4199 VDD.n4198 146.341
R3093 VDD.n4195 VDD.n4194 146.341
R3094 VDD.n4044 VDD.n4043 146.341
R3095 VDD.n4187 VDD.n4186 146.341
R3096 VDD.n4183 VDD.n4182 146.341
R3097 VDD.n4179 VDD.n4178 146.341
R3098 VDD.n4175 VDD.n4174 146.341
R3099 VDD.n4171 VDD.n4170 146.341
R3100 VDD.n4167 VDD.n4166 146.341
R3101 VDD.n4163 VDD.n4162 146.341
R3102 VDD.n4159 VDD.n4158 146.341
R3103 VDD.n4155 VDD.n4154 146.341
R3104 VDD.n4151 VDD.n4150 146.341
R3105 VDD.n4147 VDD.n4146 146.341
R3106 VDD.n4143 VDD.n4142 146.341
R3107 VDD.n4139 VDD.n4138 146.341
R3108 VDD.n4135 VDD.n4134 146.341
R3109 VDD.n4131 VDD.n4130 146.341
R3110 VDD.n4127 VDD.n4126 146.341
R3111 VDD.n3699 VDD.n286 146.341
R3112 VDD.n3699 VDD.n282 146.341
R3113 VDD.n3705 VDD.n282 146.341
R3114 VDD.n3705 VDD.n273 146.341
R3115 VDD.n3715 VDD.n273 146.341
R3116 VDD.n3715 VDD.n269 146.341
R3117 VDD.n3721 VDD.n269 146.341
R3118 VDD.n3721 VDD.n262 146.341
R3119 VDD.n3731 VDD.n262 146.341
R3120 VDD.n3731 VDD.n258 146.341
R3121 VDD.n3737 VDD.n258 146.341
R3122 VDD.n3737 VDD.n250 146.341
R3123 VDD.n3747 VDD.n250 146.341
R3124 VDD.n3747 VDD.n246 146.341
R3125 VDD.n3753 VDD.n246 146.341
R3126 VDD.n3753 VDD.n238 146.341
R3127 VDD.n3763 VDD.n238 146.341
R3128 VDD.n3763 VDD.n234 146.341
R3129 VDD.n3769 VDD.n234 146.341
R3130 VDD.n3769 VDD.n226 146.341
R3131 VDD.n3778 VDD.n226 146.341
R3132 VDD.n3778 VDD.n222 146.341
R3133 VDD.n3784 VDD.n222 146.341
R3134 VDD.n3784 VDD.n214 146.341
R3135 VDD.n3794 VDD.n214 146.341
R3136 VDD.n3794 VDD.n210 146.341
R3137 VDD.n3800 VDD.n210 146.341
R3138 VDD.n3800 VDD.n202 146.341
R3139 VDD.n3810 VDD.n202 146.341
R3140 VDD.n3810 VDD.n198 146.341
R3141 VDD.n3816 VDD.n198 146.341
R3142 VDD.n3816 VDD.n191 146.341
R3143 VDD.n3827 VDD.n191 146.341
R3144 VDD.n3827 VDD.n187 146.341
R3145 VDD.n3833 VDD.n187 146.341
R3146 VDD.n3833 VDD.n179 146.341
R3147 VDD.n3843 VDD.n179 146.341
R3148 VDD.n3843 VDD.n175 146.341
R3149 VDD.n3849 VDD.n175 146.341
R3150 VDD.n3849 VDD.n167 146.341
R3151 VDD.n3859 VDD.n167 146.341
R3152 VDD.n3859 VDD.n163 146.341
R3153 VDD.n3867 VDD.n163 146.341
R3154 VDD.n3867 VDD.n156 146.341
R3155 VDD.n3878 VDD.n156 146.341
R3156 VDD.n3879 VDD.n3878 146.341
R3157 VDD.n3879 VDD.n152 146.341
R3158 VDD.n3885 VDD.n152 146.341
R3159 VDD.n3885 VDD.n143 146.341
R3160 VDD.n3897 VDD.n143 146.341
R3161 VDD.n3897 VDD.n144 146.341
R3162 VDD.n144 VDD.n40 146.341
R3163 VDD.n41 VDD.n40 146.341
R3164 VDD.n42 VDD.n41 146.341
R3165 VDD.n137 VDD.n42 146.341
R3166 VDD.n137 VDD.n51 146.341
R3167 VDD.n52 VDD.n51 146.341
R3168 VDD.n53 VDD.n52 146.341
R3169 VDD.n134 VDD.n53 146.341
R3170 VDD.n134 VDD.n62 146.341
R3171 VDD.n63 VDD.n62 146.341
R3172 VDD.n64 VDD.n63 146.341
R3173 VDD.n131 VDD.n64 146.341
R3174 VDD.n131 VDD.n73 146.341
R3175 VDD.n74 VDD.n73 146.341
R3176 VDD.n75 VDD.n74 146.341
R3177 VDD.n128 VDD.n75 146.341
R3178 VDD.n128 VDD.n84 146.341
R3179 VDD.n85 VDD.n84 146.341
R3180 VDD.n86 VDD.n85 146.341
R3181 VDD.n125 VDD.n86 146.341
R3182 VDD.n125 VDD.n95 146.341
R3183 VDD.n96 VDD.n95 146.341
R3184 VDD.n97 VDD.n96 146.341
R3185 VDD.n122 VDD.n97 146.341
R3186 VDD.n122 VDD.n106 146.341
R3187 VDD.n107 VDD.n106 146.341
R3188 VDD.n108 VDD.n107 146.341
R3189 VDD.n118 VDD.n108 146.341
R3190 VDD.n4267 VDD.n118 146.341
R3191 VDD.n4267 VDD.n119 146.341
R3192 VDD.n4263 VDD.n119 146.341
R3193 VDD.n4263 VDD.n3947 146.341
R3194 VDD.n3956 VDD.n3947 146.341
R3195 VDD.n3957 VDD.n3956 146.341
R3196 VDD.n3958 VDD.n3957 146.341
R3197 VDD.n4097 VDD.n3958 146.341
R3198 VDD.n4097 VDD.n3967 146.341
R3199 VDD.n3968 VDD.n3967 146.341
R3200 VDD.n3969 VDD.n3968 146.341
R3201 VDD.n4104 VDD.n3969 146.341
R3202 VDD.n4104 VDD.n3978 146.341
R3203 VDD.n3979 VDD.n3978 146.341
R3204 VDD.n3980 VDD.n3979 146.341
R3205 VDD.n4111 VDD.n3980 146.341
R3206 VDD.n4111 VDD.n3989 146.341
R3207 VDD.n3990 VDD.n3989 146.341
R3208 VDD.n3991 VDD.n3990 146.341
R3209 VDD.n4118 VDD.n3991 146.341
R3210 VDD.n4118 VDD.n4000 146.341
R3211 VDD.n4001 VDD.n4000 146.341
R3212 VDD.n3685 VDD.n3682 146.341
R3213 VDD.n3682 VDD.n297 146.341
R3214 VDD.n3690 VDD.n296 146.341
R3215 VDD.n3571 VDD.n3570 146.341
R3216 VDD.n3578 VDD.n3577 146.341
R3217 VDD.n3581 VDD.n3580 146.341
R3218 VDD.n3588 VDD.n3587 146.341
R3219 VDD.n3591 VDD.n3590 146.341
R3220 VDD.n3600 VDD.n3599 146.341
R3221 VDD.n3603 VDD.n3602 146.341
R3222 VDD.n3610 VDD.n3609 146.341
R3223 VDD.n3613 VDD.n3612 146.341
R3224 VDD.n3620 VDD.n3619 146.341
R3225 VDD.n3623 VDD.n3622 146.341
R3226 VDD.n3630 VDD.n3629 146.341
R3227 VDD.n3636 VDD.n3635 146.341
R3228 VDD.n3643 VDD.n3642 146.341
R3229 VDD.n3646 VDD.n3645 146.341
R3230 VDD.n3653 VDD.n3652 146.341
R3231 VDD.n3656 VDD.n3655 146.341
R3232 VDD.n3663 VDD.n3662 146.341
R3233 VDD.n3666 VDD.n3665 146.341
R3234 VDD.n3673 VDD.n3672 146.341
R3235 VDD.n3676 VDD.n319 146.341
R3236 VDD.n3697 VDD.n288 146.341
R3237 VDD.n3697 VDD.n280 146.341
R3238 VDD.n3707 VDD.n280 146.341
R3239 VDD.n3707 VDD.n276 146.341
R3240 VDD.n3713 VDD.n276 146.341
R3241 VDD.n3713 VDD.n268 146.341
R3242 VDD.n3723 VDD.n268 146.341
R3243 VDD.n3723 VDD.n264 146.341
R3244 VDD.n3729 VDD.n264 146.341
R3245 VDD.n3729 VDD.n256 146.341
R3246 VDD.n3739 VDD.n256 146.341
R3247 VDD.n3739 VDD.n252 146.341
R3248 VDD.n3745 VDD.n252 146.341
R3249 VDD.n3745 VDD.n244 146.341
R3250 VDD.n3755 VDD.n244 146.341
R3251 VDD.n3755 VDD.n240 146.341
R3252 VDD.n3761 VDD.n240 146.341
R3253 VDD.n3761 VDD.n232 146.341
R3254 VDD.n3771 VDD.n232 146.341
R3255 VDD.n3771 VDD.n228 146.341
R3256 VDD.n3777 VDD.n228 146.341
R3257 VDD.n3777 VDD.n220 146.341
R3258 VDD.n3786 VDD.n220 146.341
R3259 VDD.n3786 VDD.n216 146.341
R3260 VDD.n3792 VDD.n216 146.341
R3261 VDD.n3792 VDD.n208 146.341
R3262 VDD.n3802 VDD.n208 146.341
R3263 VDD.n3802 VDD.n204 146.341
R3264 VDD.n3808 VDD.n204 146.341
R3265 VDD.n3808 VDD.n196 146.341
R3266 VDD.n3819 VDD.n196 146.341
R3267 VDD.n3819 VDD.n192 146.341
R3268 VDD.n3825 VDD.n192 146.341
R3269 VDD.n3825 VDD.n185 146.341
R3270 VDD.n3835 VDD.n185 146.341
R3271 VDD.n3835 VDD.n181 146.341
R3272 VDD.n3841 VDD.n181 146.341
R3273 VDD.n3841 VDD.n173 146.341
R3274 VDD.n3851 VDD.n173 146.341
R3275 VDD.n3851 VDD.n169 146.341
R3276 VDD.n3857 VDD.n169 146.341
R3277 VDD.n3857 VDD.n161 146.341
R3278 VDD.n3870 VDD.n161 146.341
R3279 VDD.n3870 VDD.n157 146.341
R3280 VDD.n3876 VDD.n157 146.341
R3281 VDD.n3876 VDD.n150 146.341
R3282 VDD.n3888 VDD.n150 146.341
R3283 VDD.n3888 VDD.n146 146.341
R3284 VDD.n3894 VDD.n146 146.341
R3285 VDD.n3895 VDD.n3894 146.341
R3286 VDD.n3895 VDD.n36 146.341
R3287 VDD.n4324 VDD.n36 146.341
R3288 VDD.n4324 VDD.n38 146.341
R3289 VDD.n4320 VDD.n38 146.341
R3290 VDD.n4320 VDD.n44 146.341
R3291 VDD.n4316 VDD.n44 146.341
R3292 VDD.n4316 VDD.n50 146.341
R3293 VDD.n4312 VDD.n50 146.341
R3294 VDD.n4312 VDD.n55 146.341
R3295 VDD.n4308 VDD.n55 146.341
R3296 VDD.n4308 VDD.n61 146.341
R3297 VDD.n4304 VDD.n61 146.341
R3298 VDD.n4304 VDD.n66 146.341
R3299 VDD.n4300 VDD.n66 146.341
R3300 VDD.n4300 VDD.n72 146.341
R3301 VDD.n4296 VDD.n72 146.341
R3302 VDD.n4296 VDD.n77 146.341
R3303 VDD.n4292 VDD.n77 146.341
R3304 VDD.n4292 VDD.n83 146.341
R3305 VDD.n4288 VDD.n83 146.341
R3306 VDD.n4288 VDD.n88 146.341
R3307 VDD.n4284 VDD.n88 146.341
R3308 VDD.n4284 VDD.n94 146.341
R3309 VDD.n4280 VDD.n94 146.341
R3310 VDD.n4280 VDD.n99 146.341
R3311 VDD.n4276 VDD.n99 146.341
R3312 VDD.n4276 VDD.n105 146.341
R3313 VDD.n4272 VDD.n105 146.341
R3314 VDD.n4272 VDD.n110 146.341
R3315 VDD.n4268 VDD.n110 146.341
R3316 VDD.n4268 VDD.n116 146.341
R3317 VDD.n4261 VDD.n116 146.341
R3318 VDD.n4261 VDD.n3949 146.341
R3319 VDD.n4257 VDD.n3949 146.341
R3320 VDD.n4257 VDD.n3955 146.341
R3321 VDD.n4253 VDD.n3955 146.341
R3322 VDD.n4253 VDD.n3960 146.341
R3323 VDD.n4249 VDD.n3960 146.341
R3324 VDD.n4249 VDD.n3966 146.341
R3325 VDD.n4245 VDD.n3966 146.341
R3326 VDD.n4245 VDD.n3971 146.341
R3327 VDD.n4241 VDD.n3971 146.341
R3328 VDD.n4241 VDD.n3977 146.341
R3329 VDD.n4237 VDD.n3977 146.341
R3330 VDD.n4237 VDD.n3981 146.341
R3331 VDD.n4233 VDD.n3981 146.341
R3332 VDD.n4233 VDD.n3987 146.341
R3333 VDD.n4229 VDD.n3987 146.341
R3334 VDD.n4229 VDD.n3993 146.341
R3335 VDD.n4225 VDD.n3993 146.341
R3336 VDD.n4225 VDD.n3999 146.341
R3337 VDD.n1100 VDD.n1074 146.341
R3338 VDD.n2192 VDD.n2189 146.341
R3339 VDD.n2186 VDD.n2185 146.341
R3340 VDD.n2182 VDD.n2181 146.341
R3341 VDD.n2178 VDD.n2177 146.341
R3342 VDD.n2174 VDD.n2173 146.341
R3343 VDD.n2170 VDD.n2169 146.341
R3344 VDD.n1114 VDD.n1113 146.341
R3345 VDD.n2162 VDD.n2161 146.341
R3346 VDD.n2158 VDD.n2157 146.341
R3347 VDD.n2154 VDD.n2153 146.341
R3348 VDD.n2150 VDD.n2149 146.341
R3349 VDD.n2146 VDD.n2145 146.341
R3350 VDD.n2142 VDD.n2141 146.341
R3351 VDD.n2138 VDD.n2137 146.341
R3352 VDD.n2134 VDD.n2133 146.341
R3353 VDD.n2130 VDD.n2129 146.341
R3354 VDD.n2126 VDD.n2125 146.341
R3355 VDD.n2122 VDD.n2121 146.341
R3356 VDD.n2118 VDD.n2117 146.341
R3357 VDD.n2114 VDD.n2113 146.341
R3358 VDD.n2110 VDD.n2109 146.341
R3359 VDD.n2106 VDD.n2105 146.341
R3360 VDD.n1198 VDD.n1197 146.341
R3361 VDD.n1681 VDD.n1497 146.341
R3362 VDD.n1681 VDD.n1489 146.341
R3363 VDD.n1691 VDD.n1489 146.341
R3364 VDD.n1691 VDD.n1485 146.341
R3365 VDD.n1697 VDD.n1485 146.341
R3366 VDD.n1697 VDD.n1478 146.341
R3367 VDD.n1708 VDD.n1478 146.341
R3368 VDD.n1708 VDD.n1474 146.341
R3369 VDD.n1714 VDD.n1474 146.341
R3370 VDD.n1714 VDD.n1466 146.341
R3371 VDD.n1724 VDD.n1466 146.341
R3372 VDD.n1724 VDD.n1462 146.341
R3373 VDD.n1730 VDD.n1462 146.341
R3374 VDD.n1730 VDD.n1454 146.341
R3375 VDD.n1740 VDD.n1454 146.341
R3376 VDD.n1740 VDD.n1450 146.341
R3377 VDD.n1746 VDD.n1450 146.341
R3378 VDD.n1746 VDD.n1442 146.341
R3379 VDD.n1756 VDD.n1442 146.341
R3380 VDD.n1756 VDD.n1438 146.341
R3381 VDD.n1762 VDD.n1438 146.341
R3382 VDD.n1762 VDD.n1430 146.341
R3383 VDD.n1771 VDD.n1430 146.341
R3384 VDD.n1771 VDD.n1426 146.341
R3385 VDD.n1777 VDD.n1426 146.341
R3386 VDD.n1777 VDD.n1418 146.341
R3387 VDD.n1787 VDD.n1418 146.341
R3388 VDD.n1787 VDD.n1414 146.341
R3389 VDD.n1793 VDD.n1414 146.341
R3390 VDD.n1793 VDD.n1405 146.341
R3391 VDD.n1803 VDD.n1405 146.341
R3392 VDD.n1803 VDD.n1401 146.341
R3393 VDD.n1809 VDD.n1401 146.341
R3394 VDD.n1809 VDD.n1394 146.341
R3395 VDD.n1819 VDD.n1394 146.341
R3396 VDD.n1819 VDD.n1390 146.341
R3397 VDD.n1825 VDD.n1390 146.341
R3398 VDD.n1825 VDD.n1382 146.341
R3399 VDD.n1835 VDD.n1382 146.341
R3400 VDD.n1835 VDD.n1378 146.341
R3401 VDD.n1841 VDD.n1378 146.341
R3402 VDD.n1841 VDD.n1369 146.341
R3403 VDD.n1851 VDD.n1369 146.341
R3404 VDD.n1851 VDD.n1365 146.341
R3405 VDD.n1857 VDD.n1365 146.341
R3406 VDD.n1857 VDD.n1358 146.341
R3407 VDD.n1867 VDD.n1358 146.341
R3408 VDD.n1867 VDD.n1354 146.341
R3409 VDD.n1873 VDD.n1354 146.341
R3410 VDD.n1873 VDD.n1346 146.341
R3411 VDD.n1902 VDD.n1346 146.341
R3412 VDD.n1902 VDD.n1342 146.341
R3413 VDD.n1908 VDD.n1342 146.341
R3414 VDD.n1908 VDD.n1333 146.341
R3415 VDD.n1918 VDD.n1333 146.341
R3416 VDD.n1918 VDD.n1329 146.341
R3417 VDD.n1924 VDD.n1329 146.341
R3418 VDD.n1924 VDD.n1322 146.341
R3419 VDD.n1934 VDD.n1322 146.341
R3420 VDD.n1934 VDD.n1318 146.341
R3421 VDD.n1940 VDD.n1318 146.341
R3422 VDD.n1940 VDD.n1310 146.341
R3423 VDD.n1950 VDD.n1310 146.341
R3424 VDD.n1950 VDD.n1306 146.341
R3425 VDD.n1956 VDD.n1306 146.341
R3426 VDD.n1956 VDD.n1297 146.341
R3427 VDD.n1966 VDD.n1297 146.341
R3428 VDD.n1966 VDD.n1293 146.341
R3429 VDD.n1972 VDD.n1293 146.341
R3430 VDD.n1972 VDD.n1286 146.341
R3431 VDD.n1982 VDD.n1286 146.341
R3432 VDD.n1982 VDD.n1282 146.341
R3433 VDD.n1988 VDD.n1282 146.341
R3434 VDD.n1988 VDD.n1274 146.341
R3435 VDD.n1998 VDD.n1274 146.341
R3436 VDD.n1998 VDD.n1270 146.341
R3437 VDD.n2004 VDD.n1270 146.341
R3438 VDD.n2004 VDD.n1262 146.341
R3439 VDD.n2014 VDD.n1262 146.341
R3440 VDD.n2014 VDD.n1258 146.341
R3441 VDD.n2020 VDD.n1258 146.341
R3442 VDD.n2020 VDD.n1251 146.341
R3443 VDD.n2030 VDD.n1251 146.341
R3444 VDD.n2030 VDD.n1247 146.341
R3445 VDD.n2036 VDD.n1247 146.341
R3446 VDD.n2036 VDD.n1239 146.341
R3447 VDD.n2046 VDD.n1239 146.341
R3448 VDD.n2046 VDD.n1235 146.341
R3449 VDD.n2052 VDD.n1235 146.341
R3450 VDD.n2052 VDD.n1227 146.341
R3451 VDD.n2062 VDD.n1227 146.341
R3452 VDD.n2062 VDD.n1223 146.341
R3453 VDD.n2068 VDD.n1223 146.341
R3454 VDD.n2068 VDD.n1216 146.341
R3455 VDD.n2079 VDD.n1216 146.341
R3456 VDD.n2079 VDD.n1211 146.341
R3457 VDD.n2087 VDD.n1211 146.341
R3458 VDD.n2087 VDD.n1203 146.341
R3459 VDD.n2097 VDD.n1203 146.341
R3460 VDD.n2098 VDD.n2097 146.341
R3461 VDD.n2098 VDD.n1076 146.341
R3462 VDD.n1527 VDD.n1526 146.341
R3463 VDD.n1531 VDD.n1526 146.341
R3464 VDD.n1533 VDD.n1532 146.341
R3465 VDD.n1537 VDD.n1536 146.341
R3466 VDD.n1539 VDD.n1538 146.341
R3467 VDD.n1543 VDD.n1542 146.341
R3468 VDD.n1545 VDD.n1544 146.341
R3469 VDD.n1551 VDD.n1550 146.341
R3470 VDD.n1553 VDD.n1552 146.341
R3471 VDD.n1557 VDD.n1556 146.341
R3472 VDD.n1559 VDD.n1558 146.341
R3473 VDD.n1563 VDD.n1562 146.341
R3474 VDD.n1565 VDD.n1564 146.341
R3475 VDD.n1569 VDD.n1568 146.341
R3476 VDD.n1571 VDD.n1570 146.341
R3477 VDD.n1578 VDD.n1577 146.341
R3478 VDD.n1580 VDD.n1579 146.341
R3479 VDD.n1584 VDD.n1583 146.341
R3480 VDD.n1586 VDD.n1585 146.341
R3481 VDD.n1590 VDD.n1589 146.341
R3482 VDD.n1592 VDD.n1591 146.341
R3483 VDD.n1596 VDD.n1595 146.341
R3484 VDD.n1598 VDD.n1597 146.341
R3485 VDD.n1599 VDD.n1503 146.341
R3486 VDD.n1683 VDD.n1495 146.341
R3487 VDD.n1683 VDD.n1491 146.341
R3488 VDD.n1689 VDD.n1491 146.341
R3489 VDD.n1689 VDD.n1483 146.341
R3490 VDD.n1700 VDD.n1483 146.341
R3491 VDD.n1700 VDD.n1479 146.341
R3492 VDD.n1706 VDD.n1479 146.341
R3493 VDD.n1706 VDD.n1472 146.341
R3494 VDD.n1716 VDD.n1472 146.341
R3495 VDD.n1716 VDD.n1468 146.341
R3496 VDD.n1722 VDD.n1468 146.341
R3497 VDD.n1722 VDD.n1460 146.341
R3498 VDD.n1732 VDD.n1460 146.341
R3499 VDD.n1732 VDD.n1456 146.341
R3500 VDD.n1738 VDD.n1456 146.341
R3501 VDD.n1738 VDD.n1448 146.341
R3502 VDD.n1748 VDD.n1448 146.341
R3503 VDD.n1748 VDD.n1444 146.341
R3504 VDD.n1754 VDD.n1444 146.341
R3505 VDD.n1754 VDD.n1436 146.341
R3506 VDD.n1763 VDD.n1436 146.341
R3507 VDD.n1763 VDD.n1432 146.341
R3508 VDD.n1769 VDD.n1432 146.341
R3509 VDD.n1769 VDD.n1424 146.341
R3510 VDD.n1779 VDD.n1424 146.341
R3511 VDD.n1779 VDD.n1420 146.341
R3512 VDD.n1785 VDD.n1420 146.341
R3513 VDD.n1785 VDD.n1412 146.341
R3514 VDD.n1795 VDD.n1412 146.341
R3515 VDD.n1795 VDD.n1408 146.341
R3516 VDD.n1801 VDD.n1408 146.341
R3517 VDD.n1801 VDD.n1400 146.341
R3518 VDD.n1811 VDD.n1400 146.341
R3519 VDD.n1811 VDD.n1396 146.341
R3520 VDD.n1817 VDD.n1396 146.341
R3521 VDD.n1817 VDD.n1388 146.341
R3522 VDD.n1827 VDD.n1388 146.341
R3523 VDD.n1827 VDD.n1384 146.341
R3524 VDD.n1833 VDD.n1384 146.341
R3525 VDD.n1833 VDD.n1376 146.341
R3526 VDD.n1843 VDD.n1376 146.341
R3527 VDD.n1843 VDD.n1372 146.341
R3528 VDD.n1849 VDD.n1372 146.341
R3529 VDD.n1849 VDD.n1364 146.341
R3530 VDD.n1859 VDD.n1364 146.341
R3531 VDD.n1859 VDD.n1360 146.341
R3532 VDD.n1865 VDD.n1360 146.341
R3533 VDD.n1865 VDD.n1352 146.341
R3534 VDD.n1875 VDD.n1352 146.341
R3535 VDD.n1875 VDD.n1348 146.341
R3536 VDD.n1900 VDD.n1348 146.341
R3537 VDD.n1900 VDD.n1340 146.341
R3538 VDD.n1910 VDD.n1340 146.341
R3539 VDD.n1910 VDD.n1336 146.341
R3540 VDD.n1916 VDD.n1336 146.341
R3541 VDD.n1916 VDD.n1328 146.341
R3542 VDD.n1926 VDD.n1328 146.341
R3543 VDD.n1926 VDD.n1324 146.341
R3544 VDD.n1932 VDD.n1324 146.341
R3545 VDD.n1932 VDD.n1316 146.341
R3546 VDD.n1942 VDD.n1316 146.341
R3547 VDD.n1942 VDD.n1312 146.341
R3548 VDD.n1948 VDD.n1312 146.341
R3549 VDD.n1948 VDD.n1304 146.341
R3550 VDD.n1958 VDD.n1304 146.341
R3551 VDD.n1958 VDD.n1300 146.341
R3552 VDD.n1964 VDD.n1300 146.341
R3553 VDD.n1964 VDD.n1292 146.341
R3554 VDD.n1974 VDD.n1292 146.341
R3555 VDD.n1974 VDD.n1288 146.341
R3556 VDD.n1980 VDD.n1288 146.341
R3557 VDD.n1980 VDD.n1280 146.341
R3558 VDD.n1990 VDD.n1280 146.341
R3559 VDD.n1990 VDD.n1276 146.341
R3560 VDD.n1996 VDD.n1276 146.341
R3561 VDD.n1996 VDD.n1268 146.341
R3562 VDD.n2006 VDD.n1268 146.341
R3563 VDD.n2006 VDD.n1264 146.341
R3564 VDD.n2012 VDD.n1264 146.341
R3565 VDD.n2012 VDD.n1257 146.341
R3566 VDD.n2022 VDD.n1257 146.341
R3567 VDD.n2022 VDD.n1253 146.341
R3568 VDD.n2028 VDD.n1253 146.341
R3569 VDD.n2028 VDD.n1245 146.341
R3570 VDD.n2038 VDD.n1245 146.341
R3571 VDD.n2038 VDD.n1241 146.341
R3572 VDD.n2044 VDD.n1241 146.341
R3573 VDD.n2044 VDD.n1233 146.341
R3574 VDD.n2054 VDD.n1233 146.341
R3575 VDD.n2054 VDD.n1229 146.341
R3576 VDD.n2060 VDD.n1229 146.341
R3577 VDD.n2060 VDD.n1221 146.341
R3578 VDD.n2071 VDD.n1221 146.341
R3579 VDD.n2071 VDD.n1217 146.341
R3580 VDD.n2077 VDD.n1217 146.341
R3581 VDD.n2077 VDD.n1209 146.341
R3582 VDD.n2089 VDD.n1209 146.341
R3583 VDD.n2089 VDD.n1205 146.341
R3584 VDD.n2095 VDD.n1205 146.341
R3585 VDD.n2095 VDD.n1073 146.341
R3586 VDD.n2196 VDD.n1073 146.341
R3587 VDD.n2399 VDD.t128 118.465
R3588 VDD.n323 VDD.t144 118.465
R3589 VDD.n3174 VDD.n2784 103.746
R3590 VDD.n1501 VDD.n1500 101.624
R3591 VDD.n1575 VDD.n1574 101.624
R3592 VDD.n1547 VDD.n1546 101.624
R3593 VDD.n1196 VDD.n1195 101.624
R3594 VDD.n1130 VDD.n1129 101.624
R3595 VDD.n1112 VDD.n1111 101.624
R3596 VDD.n4081 VDD.n4080 101.624
R3597 VDD.n4060 VDD.n4059 101.624
R3598 VDD.n4042 VDD.n4041 101.624
R3599 VDD.n3593 VDD.n3592 101.624
R3600 VDD.n3633 VDD.n3632 101.624
R3601 VDD.n3550 VDD.n3549 101.624
R3602 VDD.n3182 VDD.n621 99.5127
R3603 VDD.n3182 VDD.n619 99.5127
R3604 VDD.n3186 VDD.n619 99.5127
R3605 VDD.n3186 VDD.n608 99.5127
R3606 VDD.n3194 VDD.n608 99.5127
R3607 VDD.n3194 VDD.n606 99.5127
R3608 VDD.n3198 VDD.n606 99.5127
R3609 VDD.n3198 VDD.n597 99.5127
R3610 VDD.n3206 VDD.n597 99.5127
R3611 VDD.n3206 VDD.n595 99.5127
R3612 VDD.n3210 VDD.n595 99.5127
R3613 VDD.n3210 VDD.n585 99.5127
R3614 VDD.n3218 VDD.n585 99.5127
R3615 VDD.n3218 VDD.n583 99.5127
R3616 VDD.n3222 VDD.n583 99.5127
R3617 VDD.n3222 VDD.n573 99.5127
R3618 VDD.n3230 VDD.n573 99.5127
R3619 VDD.n3230 VDD.n571 99.5127
R3620 VDD.n3234 VDD.n571 99.5127
R3621 VDD.n3234 VDD.n561 99.5127
R3622 VDD.n3242 VDD.n561 99.5127
R3623 VDD.n3242 VDD.n559 99.5127
R3624 VDD.n3246 VDD.n559 99.5127
R3625 VDD.n3246 VDD.n549 99.5127
R3626 VDD.n3254 VDD.n549 99.5127
R3627 VDD.n3254 VDD.n547 99.5127
R3628 VDD.n3258 VDD.n547 99.5127
R3629 VDD.n3258 VDD.n537 99.5127
R3630 VDD.n3266 VDD.n537 99.5127
R3631 VDD.n3266 VDD.n535 99.5127
R3632 VDD.n3270 VDD.n535 99.5127
R3633 VDD.n3270 VDD.n525 99.5127
R3634 VDD.n3278 VDD.n525 99.5127
R3635 VDD.n3278 VDD.n523 99.5127
R3636 VDD.n3282 VDD.n523 99.5127
R3637 VDD.n3282 VDD.n512 99.5127
R3638 VDD.n3290 VDD.n512 99.5127
R3639 VDD.n3290 VDD.n510 99.5127
R3640 VDD.n3294 VDD.n510 99.5127
R3641 VDD.n3294 VDD.n501 99.5127
R3642 VDD.n3302 VDD.n501 99.5127
R3643 VDD.n3302 VDD.n499 99.5127
R3644 VDD.n3306 VDD.n499 99.5127
R3645 VDD.n3306 VDD.n489 99.5127
R3646 VDD.n3314 VDD.n489 99.5127
R3647 VDD.n3314 VDD.n487 99.5127
R3648 VDD.n3318 VDD.n487 99.5127
R3649 VDD.n3318 VDD.n476 99.5127
R3650 VDD.n3326 VDD.n476 99.5127
R3651 VDD.n3326 VDD.n474 99.5127
R3652 VDD.n3330 VDD.n474 99.5127
R3653 VDD.n3330 VDD.n465 99.5127
R3654 VDD.n3338 VDD.n465 99.5127
R3655 VDD.n3338 VDD.n463 99.5127
R3656 VDD.n3342 VDD.n463 99.5127
R3657 VDD.n3342 VDD.n453 99.5127
R3658 VDD.n3350 VDD.n453 99.5127
R3659 VDD.n3350 VDD.n451 99.5127
R3660 VDD.n3354 VDD.n451 99.5127
R3661 VDD.n3354 VDD.n441 99.5127
R3662 VDD.n3362 VDD.n441 99.5127
R3663 VDD.n3362 VDD.n439 99.5127
R3664 VDD.n3366 VDD.n439 99.5127
R3665 VDD.n3366 VDD.n430 99.5127
R3666 VDD.n3374 VDD.n430 99.5127
R3667 VDD.n3374 VDD.n428 99.5127
R3668 VDD.n3378 VDD.n428 99.5127
R3669 VDD.n3378 VDD.n418 99.5127
R3670 VDD.n3386 VDD.n418 99.5127
R3671 VDD.n3386 VDD.n416 99.5127
R3672 VDD.n3390 VDD.n416 99.5127
R3673 VDD.n3390 VDD.n406 99.5127
R3674 VDD.n3398 VDD.n406 99.5127
R3675 VDD.n3398 VDD.n404 99.5127
R3676 VDD.n3402 VDD.n404 99.5127
R3677 VDD.n3402 VDD.n394 99.5127
R3678 VDD.n3410 VDD.n394 99.5127
R3679 VDD.n3410 VDD.n392 99.5127
R3680 VDD.n3414 VDD.n392 99.5127
R3681 VDD.n3414 VDD.n382 99.5127
R3682 VDD.n3422 VDD.n382 99.5127
R3683 VDD.n3422 VDD.n380 99.5127
R3684 VDD.n3426 VDD.n380 99.5127
R3685 VDD.n3426 VDD.n369 99.5127
R3686 VDD.n3467 VDD.n369 99.5127
R3687 VDD.n3467 VDD.n367 99.5127
R3688 VDD.n3471 VDD.n367 99.5127
R3689 VDD.n3471 VDD.n340 99.5127
R3690 VDD.n3522 VDD.n340 99.5127
R3691 VDD.n3518 VDD.n341 99.5127
R3692 VDD.n3516 VDD.n3515 99.5127
R3693 VDD.n3513 VDD.n345 99.5127
R3694 VDD.n3509 VDD.n3508 99.5127
R3695 VDD.n3506 VDD.n348 99.5127
R3696 VDD.n3502 VDD.n3501 99.5127
R3697 VDD.n3499 VDD.n3498 99.5127
R3698 VDD.n3496 VDD.n352 99.5127
R3699 VDD.n3492 VDD.n3491 99.5127
R3700 VDD.n3489 VDD.n355 99.5127
R3701 VDD.n3485 VDD.n3484 99.5127
R3702 VDD.n3482 VDD.n361 99.5127
R3703 VDD.n3124 VDD.n623 99.5127
R3704 VDD.n3120 VDD.n623 99.5127
R3705 VDD.n3120 VDD.n617 99.5127
R3706 VDD.n3117 VDD.n617 99.5127
R3707 VDD.n3117 VDD.n610 99.5127
R3708 VDD.n3114 VDD.n610 99.5127
R3709 VDD.n3114 VDD.n603 99.5127
R3710 VDD.n3111 VDD.n603 99.5127
R3711 VDD.n3111 VDD.n598 99.5127
R3712 VDD.n3108 VDD.n598 99.5127
R3713 VDD.n3108 VDD.n593 99.5127
R3714 VDD.n3105 VDD.n593 99.5127
R3715 VDD.n3105 VDD.n587 99.5127
R3716 VDD.n3102 VDD.n587 99.5127
R3717 VDD.n3102 VDD.n581 99.5127
R3718 VDD.n3099 VDD.n581 99.5127
R3719 VDD.n3099 VDD.n575 99.5127
R3720 VDD.n3096 VDD.n575 99.5127
R3721 VDD.n3096 VDD.n569 99.5127
R3722 VDD.n3093 VDD.n569 99.5127
R3723 VDD.n3093 VDD.n563 99.5127
R3724 VDD.n3090 VDD.n563 99.5127
R3725 VDD.n3090 VDD.n557 99.5127
R3726 VDD.n3087 VDD.n557 99.5127
R3727 VDD.n3087 VDD.n551 99.5127
R3728 VDD.n3084 VDD.n551 99.5127
R3729 VDD.n3084 VDD.n545 99.5127
R3730 VDD.n3081 VDD.n545 99.5127
R3731 VDD.n3081 VDD.n539 99.5127
R3732 VDD.n3078 VDD.n539 99.5127
R3733 VDD.n3078 VDD.n532 99.5127
R3734 VDD.n3075 VDD.n532 99.5127
R3735 VDD.n3075 VDD.n526 99.5127
R3736 VDD.n3072 VDD.n526 99.5127
R3737 VDD.n3072 VDD.n521 99.5127
R3738 VDD.n3069 VDD.n521 99.5127
R3739 VDD.n3069 VDD.n514 99.5127
R3740 VDD.n3066 VDD.n514 99.5127
R3741 VDD.n3066 VDD.n508 99.5127
R3742 VDD.n3063 VDD.n508 99.5127
R3743 VDD.n3063 VDD.n503 99.5127
R3744 VDD.n3060 VDD.n503 99.5127
R3745 VDD.n3060 VDD.n497 99.5127
R3746 VDD.n3057 VDD.n497 99.5127
R3747 VDD.n3057 VDD.n491 99.5127
R3748 VDD.n3054 VDD.n491 99.5127
R3749 VDD.n3054 VDD.n485 99.5127
R3750 VDD.n3051 VDD.n485 99.5127
R3751 VDD.n3051 VDD.n478 99.5127
R3752 VDD.n3048 VDD.n478 99.5127
R3753 VDD.n3048 VDD.n472 99.5127
R3754 VDD.n3045 VDD.n472 99.5127
R3755 VDD.n3045 VDD.n467 99.5127
R3756 VDD.n3042 VDD.n467 99.5127
R3757 VDD.n3042 VDD.n461 99.5127
R3758 VDD.n3039 VDD.n461 99.5127
R3759 VDD.n3039 VDD.n455 99.5127
R3760 VDD.n3036 VDD.n455 99.5127
R3761 VDD.n3036 VDD.n449 99.5127
R3762 VDD.n3033 VDD.n449 99.5127
R3763 VDD.n3033 VDD.n443 99.5127
R3764 VDD.n3030 VDD.n443 99.5127
R3765 VDD.n3030 VDD.n437 99.5127
R3766 VDD.n3027 VDD.n437 99.5127
R3767 VDD.n3027 VDD.n431 99.5127
R3768 VDD.n2842 VDD.n431 99.5127
R3769 VDD.n2842 VDD.n426 99.5127
R3770 VDD.n2839 VDD.n426 99.5127
R3771 VDD.n2839 VDD.n420 99.5127
R3772 VDD.n2836 VDD.n420 99.5127
R3773 VDD.n2836 VDD.n414 99.5127
R3774 VDD.n2833 VDD.n414 99.5127
R3775 VDD.n2833 VDD.n408 99.5127
R3776 VDD.n2830 VDD.n408 99.5127
R3777 VDD.n2830 VDD.n402 99.5127
R3778 VDD.n2827 VDD.n402 99.5127
R3779 VDD.n2827 VDD.n396 99.5127
R3780 VDD.n2824 VDD.n396 99.5127
R3781 VDD.n2824 VDD.n389 99.5127
R3782 VDD.n2821 VDD.n389 99.5127
R3783 VDD.n2821 VDD.n383 99.5127
R3784 VDD.n2818 VDD.n383 99.5127
R3785 VDD.n2818 VDD.n378 99.5127
R3786 VDD.n2815 VDD.n378 99.5127
R3787 VDD.n2815 VDD.n371 99.5127
R3788 VDD.n371 VDD.n363 99.5127
R3789 VDD.n3473 VDD.n363 99.5127
R3790 VDD.n3474 VDD.n3473 99.5127
R3791 VDD.n3474 VDD.n338 99.5127
R3792 VDD.n2809 VDD.n2808 99.5127
R3793 VDD.n3167 VDD.n2808 99.5127
R3794 VDD.n3165 VDD.n3164 99.5127
R3795 VDD.n3161 VDD.n3160 99.5127
R3796 VDD.n3157 VDD.n3156 99.5127
R3797 VDD.n3153 VDD.n3152 99.5127
R3798 VDD.n3149 VDD.n3148 99.5127
R3799 VDD.n3145 VDD.n3144 99.5127
R3800 VDD.n3141 VDD.n3140 99.5127
R3801 VDD.n3137 VDD.n3136 99.5127
R3802 VDD.n3133 VDD.n3132 99.5127
R3803 VDD.n3129 VDD.n3128 99.5127
R3804 VDD.n2783 VDD.n655 99.5127
R3805 VDD.n2779 VDD.n2778 99.5127
R3806 VDD.n2775 VDD.n2774 99.5127
R3807 VDD.n2771 VDD.n2770 99.5127
R3808 VDD.n2767 VDD.n2766 99.5127
R3809 VDD.n2763 VDD.n2762 99.5127
R3810 VDD.n2759 VDD.n2758 99.5127
R3811 VDD.n2755 VDD.n2754 99.5127
R3812 VDD.n2751 VDD.n2750 99.5127
R3813 VDD.n2747 VDD.n2746 99.5127
R3814 VDD.n2743 VDD.n2742 99.5127
R3815 VDD.n2739 VDD.n2738 99.5127
R3816 VDD.n2227 VDD.n931 99.5127
R3817 VDD.n2227 VDD.n926 99.5127
R3818 VDD.n2230 VDD.n926 99.5127
R3819 VDD.n2230 VDD.n920 99.5127
R3820 VDD.n2233 VDD.n920 99.5127
R3821 VDD.n2233 VDD.n914 99.5127
R3822 VDD.n2236 VDD.n914 99.5127
R3823 VDD.n2236 VDD.n908 99.5127
R3824 VDD.n2239 VDD.n908 99.5127
R3825 VDD.n2239 VDD.n901 99.5127
R3826 VDD.n2242 VDD.n901 99.5127
R3827 VDD.n2242 VDD.n895 99.5127
R3828 VDD.n2245 VDD.n895 99.5127
R3829 VDD.n2245 VDD.n890 99.5127
R3830 VDD.n2248 VDD.n890 99.5127
R3831 VDD.n2248 VDD.n884 99.5127
R3832 VDD.n2251 VDD.n884 99.5127
R3833 VDD.n2251 VDD.n878 99.5127
R3834 VDD.n2254 VDD.n878 99.5127
R3835 VDD.n2254 VDD.n872 99.5127
R3836 VDD.n2257 VDD.n872 99.5127
R3837 VDD.n2257 VDD.n866 99.5127
R3838 VDD.n2260 VDD.n866 99.5127
R3839 VDD.n2260 VDD.n860 99.5127
R3840 VDD.n2356 VDD.n860 99.5127
R3841 VDD.n2356 VDD.n854 99.5127
R3842 VDD.n2352 VDD.n854 99.5127
R3843 VDD.n2352 VDD.n849 99.5127
R3844 VDD.n2349 VDD.n849 99.5127
R3845 VDD.n2349 VDD.n843 99.5127
R3846 VDD.n2346 VDD.n843 99.5127
R3847 VDD.n2346 VDD.n837 99.5127
R3848 VDD.n2343 VDD.n837 99.5127
R3849 VDD.n2343 VDD.n831 99.5127
R3850 VDD.n2340 VDD.n831 99.5127
R3851 VDD.n2340 VDD.n825 99.5127
R3852 VDD.n2337 VDD.n825 99.5127
R3853 VDD.n2337 VDD.n819 99.5127
R3854 VDD.n2334 VDD.n819 99.5127
R3855 VDD.n2334 VDD.n813 99.5127
R3856 VDD.n2331 VDD.n813 99.5127
R3857 VDD.n2331 VDD.n806 99.5127
R3858 VDD.n2328 VDD.n806 99.5127
R3859 VDD.n2328 VDD.n800 99.5127
R3860 VDD.n2325 VDD.n800 99.5127
R3861 VDD.n2325 VDD.n795 99.5127
R3862 VDD.n2322 VDD.n795 99.5127
R3863 VDD.n2322 VDD.n789 99.5127
R3864 VDD.n2319 VDD.n789 99.5127
R3865 VDD.n2319 VDD.n783 99.5127
R3866 VDD.n2316 VDD.n783 99.5127
R3867 VDD.n2316 VDD.n777 99.5127
R3868 VDD.n2313 VDD.n777 99.5127
R3869 VDD.n2313 VDD.n771 99.5127
R3870 VDD.n2310 VDD.n771 99.5127
R3871 VDD.n2310 VDD.n765 99.5127
R3872 VDD.n2307 VDD.n765 99.5127
R3873 VDD.n2307 VDD.n759 99.5127
R3874 VDD.n2304 VDD.n759 99.5127
R3875 VDD.n2304 VDD.n753 99.5127
R3876 VDD.n2301 VDD.n753 99.5127
R3877 VDD.n2301 VDD.n746 99.5127
R3878 VDD.n2298 VDD.n746 99.5127
R3879 VDD.n2298 VDD.n740 99.5127
R3880 VDD.n2295 VDD.n740 99.5127
R3881 VDD.n2295 VDD.n735 99.5127
R3882 VDD.n2292 VDD.n735 99.5127
R3883 VDD.n2292 VDD.n728 99.5127
R3884 VDD.n2289 VDD.n728 99.5127
R3885 VDD.n2289 VDD.n722 99.5127
R3886 VDD.n2286 VDD.n722 99.5127
R3887 VDD.n2286 VDD.n717 99.5127
R3888 VDD.n2283 VDD.n717 99.5127
R3889 VDD.n2283 VDD.n711 99.5127
R3890 VDD.n2280 VDD.n711 99.5127
R3891 VDD.n2280 VDD.n705 99.5127
R3892 VDD.n2277 VDD.n705 99.5127
R3893 VDD.n2277 VDD.n699 99.5127
R3894 VDD.n2274 VDD.n699 99.5127
R3895 VDD.n2274 VDD.n693 99.5127
R3896 VDD.n2271 VDD.n693 99.5127
R3897 VDD.n2271 VDD.n686 99.5127
R3898 VDD.n2268 VDD.n686 99.5127
R3899 VDD.n2268 VDD.n680 99.5127
R3900 VDD.n2265 VDD.n680 99.5127
R3901 VDD.n2265 VDD.n670 99.5127
R3902 VDD.n670 VDD.n661 99.5127
R3903 VDD.n2733 VDD.n661 99.5127
R3904 VDD.n2734 VDD.n2733 99.5127
R3905 VDD.n2401 VDD.n935 99.5127
R3906 VDD.n1050 VDD.n935 99.5127
R3907 VDD.n1054 VDD.n1053 99.5127
R3908 VDD.n1058 VDD.n1057 99.5127
R3909 VDD.n1062 VDD.n1061 99.5127
R3910 VDD.n1066 VDD.n1065 99.5127
R3911 VDD.n2202 VDD.n2201 99.5127
R3912 VDD.n2206 VDD.n2205 99.5127
R3913 VDD.n2210 VDD.n2209 99.5127
R3914 VDD.n2214 VDD.n2213 99.5127
R3915 VDD.n2218 VDD.n2217 99.5127
R3916 VDD.n2222 VDD.n2221 99.5127
R3917 VDD.n2405 VDD.n924 99.5127
R3918 VDD.n2413 VDD.n924 99.5127
R3919 VDD.n2413 VDD.n922 99.5127
R3920 VDD.n2417 VDD.n922 99.5127
R3921 VDD.n2417 VDD.n912 99.5127
R3922 VDD.n2425 VDD.n912 99.5127
R3923 VDD.n2425 VDD.n910 99.5127
R3924 VDD.n2429 VDD.n910 99.5127
R3925 VDD.n2429 VDD.n899 99.5127
R3926 VDD.n2437 VDD.n899 99.5127
R3927 VDD.n2437 VDD.n897 99.5127
R3928 VDD.n2441 VDD.n897 99.5127
R3929 VDD.n2441 VDD.n888 99.5127
R3930 VDD.n2449 VDD.n888 99.5127
R3931 VDD.n2449 VDD.n886 99.5127
R3932 VDD.n2453 VDD.n886 99.5127
R3933 VDD.n2453 VDD.n876 99.5127
R3934 VDD.n2461 VDD.n876 99.5127
R3935 VDD.n2461 VDD.n874 99.5127
R3936 VDD.n2465 VDD.n874 99.5127
R3937 VDD.n2465 VDD.n864 99.5127
R3938 VDD.n2473 VDD.n864 99.5127
R3939 VDD.n2473 VDD.n862 99.5127
R3940 VDD.n2477 VDD.n862 99.5127
R3941 VDD.n2477 VDD.n853 99.5127
R3942 VDD.n2485 VDD.n853 99.5127
R3943 VDD.n2485 VDD.n851 99.5127
R3944 VDD.n2489 VDD.n851 99.5127
R3945 VDD.n2489 VDD.n841 99.5127
R3946 VDD.n2497 VDD.n841 99.5127
R3947 VDD.n2497 VDD.n839 99.5127
R3948 VDD.n2501 VDD.n839 99.5127
R3949 VDD.n2501 VDD.n829 99.5127
R3950 VDD.n2509 VDD.n829 99.5127
R3951 VDD.n2509 VDD.n827 99.5127
R3952 VDD.n2513 VDD.n827 99.5127
R3953 VDD.n2513 VDD.n817 99.5127
R3954 VDD.n2521 VDD.n817 99.5127
R3955 VDD.n2521 VDD.n815 99.5127
R3956 VDD.n2525 VDD.n815 99.5127
R3957 VDD.n2525 VDD.n804 99.5127
R3958 VDD.n2533 VDD.n804 99.5127
R3959 VDD.n2533 VDD.n802 99.5127
R3960 VDD.n2537 VDD.n802 99.5127
R3961 VDD.n2537 VDD.n793 99.5127
R3962 VDD.n2545 VDD.n793 99.5127
R3963 VDD.n2545 VDD.n791 99.5127
R3964 VDD.n2549 VDD.n791 99.5127
R3965 VDD.n2549 VDD.n781 99.5127
R3966 VDD.n2557 VDD.n781 99.5127
R3967 VDD.n2557 VDD.n779 99.5127
R3968 VDD.n2561 VDD.n779 99.5127
R3969 VDD.n2561 VDD.n769 99.5127
R3970 VDD.n2569 VDD.n769 99.5127
R3971 VDD.n2569 VDD.n767 99.5127
R3972 VDD.n2573 VDD.n767 99.5127
R3973 VDD.n2573 VDD.n757 99.5127
R3974 VDD.n2581 VDD.n757 99.5127
R3975 VDD.n2581 VDD.n755 99.5127
R3976 VDD.n2585 VDD.n755 99.5127
R3977 VDD.n2585 VDD.n744 99.5127
R3978 VDD.n2593 VDD.n744 99.5127
R3979 VDD.n2593 VDD.n742 99.5127
R3980 VDD.n2597 VDD.n742 99.5127
R3981 VDD.n2597 VDD.n733 99.5127
R3982 VDD.n2605 VDD.n733 99.5127
R3983 VDD.n2605 VDD.n731 99.5127
R3984 VDD.n2609 VDD.n731 99.5127
R3985 VDD.n2609 VDD.n721 99.5127
R3986 VDD.n2617 VDD.n721 99.5127
R3987 VDD.n2617 VDD.n719 99.5127
R3988 VDD.n2621 VDD.n719 99.5127
R3989 VDD.n2621 VDD.n709 99.5127
R3990 VDD.n2629 VDD.n709 99.5127
R3991 VDD.n2629 VDD.n707 99.5127
R3992 VDD.n2633 VDD.n707 99.5127
R3993 VDD.n2633 VDD.n697 99.5127
R3994 VDD.n2641 VDD.n697 99.5127
R3995 VDD.n2641 VDD.n695 99.5127
R3996 VDD.n2645 VDD.n695 99.5127
R3997 VDD.n2645 VDD.n684 99.5127
R3998 VDD.n2655 VDD.n684 99.5127
R3999 VDD.n2655 VDD.n682 99.5127
R4000 VDD.n2659 VDD.n682 99.5127
R4001 VDD.n2659 VDD.n668 99.5127
R4002 VDD.n2727 VDD.n668 99.5127
R4003 VDD.n2727 VDD.n666 99.5127
R4004 VDD.n2731 VDD.n666 99.5127
R4005 VDD.n2731 VDD.n654 99.5127
R4006 VDD.n3457 VDD.n3456 99.5127
R4007 VDD.n3454 VDD.n3432 99.5127
R4008 VDD.n3450 VDD.n3449 99.5127
R4009 VDD.n3447 VDD.n3435 99.5127
R4010 VDD.n3443 VDD.n3442 99.5127
R4011 VDD.n3440 VDD.n3438 99.5127
R4012 VDD.n3546 VDD.n3545 99.5127
R4013 VDD.n3543 VDD.n324 99.5127
R4014 VDD.n3539 VDD.n3538 99.5127
R4015 VDD.n3536 VDD.n327 99.5127
R4016 VDD.n3532 VDD.n3531 99.5127
R4017 VDD.n3529 VDD.n333 99.5127
R4018 VDD.n2893 VDD.n624 99.5127
R4019 VDD.n2896 VDD.n624 99.5127
R4020 VDD.n2896 VDD.n618 99.5127
R4021 VDD.n2899 VDD.n618 99.5127
R4022 VDD.n2899 VDD.n611 99.5127
R4023 VDD.n2902 VDD.n611 99.5127
R4024 VDD.n2902 VDD.n604 99.5127
R4025 VDD.n2905 VDD.n604 99.5127
R4026 VDD.n2905 VDD.n599 99.5127
R4027 VDD.n2908 VDD.n599 99.5127
R4028 VDD.n2908 VDD.n594 99.5127
R4029 VDD.n2911 VDD.n594 99.5127
R4030 VDD.n2911 VDD.n588 99.5127
R4031 VDD.n2914 VDD.n588 99.5127
R4032 VDD.n2914 VDD.n582 99.5127
R4033 VDD.n2917 VDD.n582 99.5127
R4034 VDD.n2917 VDD.n576 99.5127
R4035 VDD.n2920 VDD.n576 99.5127
R4036 VDD.n2920 VDD.n570 99.5127
R4037 VDD.n2923 VDD.n570 99.5127
R4038 VDD.n2923 VDD.n564 99.5127
R4039 VDD.n2926 VDD.n564 99.5127
R4040 VDD.n2926 VDD.n558 99.5127
R4041 VDD.n2929 VDD.n558 99.5127
R4042 VDD.n2929 VDD.n552 99.5127
R4043 VDD.n2932 VDD.n552 99.5127
R4044 VDD.n2932 VDD.n546 99.5127
R4045 VDD.n2935 VDD.n546 99.5127
R4046 VDD.n2935 VDD.n540 99.5127
R4047 VDD.n2938 VDD.n540 99.5127
R4048 VDD.n2938 VDD.n533 99.5127
R4049 VDD.n2941 VDD.n533 99.5127
R4050 VDD.n2941 VDD.n527 99.5127
R4051 VDD.n2944 VDD.n527 99.5127
R4052 VDD.n2944 VDD.n522 99.5127
R4053 VDD.n2947 VDD.n522 99.5127
R4054 VDD.n2947 VDD.n515 99.5127
R4055 VDD.n2950 VDD.n515 99.5127
R4056 VDD.n2950 VDD.n509 99.5127
R4057 VDD.n2953 VDD.n509 99.5127
R4058 VDD.n2953 VDD.n504 99.5127
R4059 VDD.n2956 VDD.n504 99.5127
R4060 VDD.n2956 VDD.n498 99.5127
R4061 VDD.n2959 VDD.n498 99.5127
R4062 VDD.n2959 VDD.n492 99.5127
R4063 VDD.n2962 VDD.n492 99.5127
R4064 VDD.n2962 VDD.n486 99.5127
R4065 VDD.n2965 VDD.n486 99.5127
R4066 VDD.n2965 VDD.n479 99.5127
R4067 VDD.n2968 VDD.n479 99.5127
R4068 VDD.n2968 VDD.n473 99.5127
R4069 VDD.n2971 VDD.n473 99.5127
R4070 VDD.n2971 VDD.n468 99.5127
R4071 VDD.n2974 VDD.n468 99.5127
R4072 VDD.n2974 VDD.n462 99.5127
R4073 VDD.n2977 VDD.n462 99.5127
R4074 VDD.n2977 VDD.n456 99.5127
R4075 VDD.n2980 VDD.n456 99.5127
R4076 VDD.n2980 VDD.n450 99.5127
R4077 VDD.n2983 VDD.n450 99.5127
R4078 VDD.n2983 VDD.n444 99.5127
R4079 VDD.n2986 VDD.n444 99.5127
R4080 VDD.n2986 VDD.n438 99.5127
R4081 VDD.n3025 VDD.n438 99.5127
R4082 VDD.n3025 VDD.n432 99.5127
R4083 VDD.n3021 VDD.n432 99.5127
R4084 VDD.n3021 VDD.n427 99.5127
R4085 VDD.n3018 VDD.n427 99.5127
R4086 VDD.n3018 VDD.n421 99.5127
R4087 VDD.n3015 VDD.n421 99.5127
R4088 VDD.n3015 VDD.n415 99.5127
R4089 VDD.n3012 VDD.n415 99.5127
R4090 VDD.n3012 VDD.n409 99.5127
R4091 VDD.n3009 VDD.n409 99.5127
R4092 VDD.n3009 VDD.n403 99.5127
R4093 VDD.n3006 VDD.n403 99.5127
R4094 VDD.n3006 VDD.n397 99.5127
R4095 VDD.n3003 VDD.n397 99.5127
R4096 VDD.n3003 VDD.n390 99.5127
R4097 VDD.n3000 VDD.n390 99.5127
R4098 VDD.n3000 VDD.n384 99.5127
R4099 VDD.n2997 VDD.n384 99.5127
R4100 VDD.n2997 VDD.n379 99.5127
R4101 VDD.n2994 VDD.n379 99.5127
R4102 VDD.n2994 VDD.n372 99.5127
R4103 VDD.n2991 VDD.n372 99.5127
R4104 VDD.n2991 VDD.n365 99.5127
R4105 VDD.n365 VDD.n336 99.5127
R4106 VDD.n3524 VDD.n336 99.5127
R4107 VDD.n2847 VDD.n627 99.5127
R4108 VDD.n2851 VDD.n2850 99.5127
R4109 VDD.n2855 VDD.n2854 99.5127
R4110 VDD.n2859 VDD.n2858 99.5127
R4111 VDD.n2863 VDD.n2862 99.5127
R4112 VDD.n2867 VDD.n2866 99.5127
R4113 VDD.n2871 VDD.n2870 99.5127
R4114 VDD.n2875 VDD.n2874 99.5127
R4115 VDD.n2879 VDD.n2878 99.5127
R4116 VDD.n2883 VDD.n2882 99.5127
R4117 VDD.n2888 VDD.n2887 99.5127
R4118 VDD.n2890 VDD.n2807 99.5127
R4119 VDD.n3180 VDD.n625 99.5127
R4120 VDD.n3180 VDD.n615 99.5127
R4121 VDD.n3188 VDD.n615 99.5127
R4122 VDD.n3188 VDD.n613 99.5127
R4123 VDD.n3192 VDD.n613 99.5127
R4124 VDD.n3192 VDD.n602 99.5127
R4125 VDD.n3200 VDD.n602 99.5127
R4126 VDD.n3200 VDD.n600 99.5127
R4127 VDD.n3204 VDD.n600 99.5127
R4128 VDD.n3204 VDD.n591 99.5127
R4129 VDD.n3212 VDD.n591 99.5127
R4130 VDD.n3212 VDD.n589 99.5127
R4131 VDD.n3216 VDD.n589 99.5127
R4132 VDD.n3216 VDD.n579 99.5127
R4133 VDD.n3224 VDD.n579 99.5127
R4134 VDD.n3224 VDD.n577 99.5127
R4135 VDD.n3228 VDD.n577 99.5127
R4136 VDD.n3228 VDD.n567 99.5127
R4137 VDD.n3236 VDD.n567 99.5127
R4138 VDD.n3236 VDD.n565 99.5127
R4139 VDD.n3240 VDD.n565 99.5127
R4140 VDD.n3240 VDD.n555 99.5127
R4141 VDD.n3248 VDD.n555 99.5127
R4142 VDD.n3248 VDD.n553 99.5127
R4143 VDD.n3252 VDD.n553 99.5127
R4144 VDD.n3252 VDD.n543 99.5127
R4145 VDD.n3260 VDD.n543 99.5127
R4146 VDD.n3260 VDD.n541 99.5127
R4147 VDD.n3264 VDD.n541 99.5127
R4148 VDD.n3264 VDD.n530 99.5127
R4149 VDD.n3272 VDD.n530 99.5127
R4150 VDD.n3272 VDD.n528 99.5127
R4151 VDD.n3276 VDD.n528 99.5127
R4152 VDD.n3276 VDD.n519 99.5127
R4153 VDD.n3284 VDD.n519 99.5127
R4154 VDD.n3284 VDD.n517 99.5127
R4155 VDD.n3288 VDD.n517 99.5127
R4156 VDD.n3288 VDD.n507 99.5127
R4157 VDD.n3296 VDD.n507 99.5127
R4158 VDD.n3296 VDD.n505 99.5127
R4159 VDD.n3300 VDD.n505 99.5127
R4160 VDD.n3300 VDD.n495 99.5127
R4161 VDD.n3308 VDD.n495 99.5127
R4162 VDD.n3308 VDD.n493 99.5127
R4163 VDD.n3312 VDD.n493 99.5127
R4164 VDD.n3312 VDD.n483 99.5127
R4165 VDD.n3320 VDD.n483 99.5127
R4166 VDD.n3320 VDD.n481 99.5127
R4167 VDD.n3324 VDD.n481 99.5127
R4168 VDD.n3324 VDD.n471 99.5127
R4169 VDD.n3332 VDD.n471 99.5127
R4170 VDD.n3332 VDD.n469 99.5127
R4171 VDD.n3336 VDD.n469 99.5127
R4172 VDD.n3336 VDD.n459 99.5127
R4173 VDD.n3344 VDD.n459 99.5127
R4174 VDD.n3344 VDD.n457 99.5127
R4175 VDD.n3348 VDD.n457 99.5127
R4176 VDD.n3348 VDD.n447 99.5127
R4177 VDD.n3356 VDD.n447 99.5127
R4178 VDD.n3356 VDD.n445 99.5127
R4179 VDD.n3360 VDD.n445 99.5127
R4180 VDD.n3360 VDD.n435 99.5127
R4181 VDD.n3368 VDD.n435 99.5127
R4182 VDD.n3368 VDD.n433 99.5127
R4183 VDD.n3372 VDD.n433 99.5127
R4184 VDD.n3372 VDD.n424 99.5127
R4185 VDD.n3380 VDD.n424 99.5127
R4186 VDD.n3380 VDD.n422 99.5127
R4187 VDD.n3384 VDD.n422 99.5127
R4188 VDD.n3384 VDD.n412 99.5127
R4189 VDD.n3392 VDD.n412 99.5127
R4190 VDD.n3392 VDD.n410 99.5127
R4191 VDD.n3396 VDD.n410 99.5127
R4192 VDD.n3396 VDD.n400 99.5127
R4193 VDD.n3404 VDD.n400 99.5127
R4194 VDD.n3404 VDD.n398 99.5127
R4195 VDD.n3408 VDD.n398 99.5127
R4196 VDD.n3408 VDD.n387 99.5127
R4197 VDD.n3416 VDD.n387 99.5127
R4198 VDD.n3416 VDD.n385 99.5127
R4199 VDD.n3420 VDD.n385 99.5127
R4200 VDD.n3420 VDD.n376 99.5127
R4201 VDD.n3428 VDD.n376 99.5127
R4202 VDD.n3428 VDD.n373 99.5127
R4203 VDD.n3465 VDD.n373 99.5127
R4204 VDD.n3465 VDD.n374 99.5127
R4205 VDD.n374 VDD.n366 99.5127
R4206 VDD.n3460 VDD.n366 99.5127
R4207 VDD.n3460 VDD.n339 99.5127
R4208 VDD.n2716 VDD.n2715 99.5127
R4209 VDD.n2712 VDD.n2711 99.5127
R4210 VDD.n2708 VDD.n2707 99.5127
R4211 VDD.n2704 VDD.n2703 99.5127
R4212 VDD.n2700 VDD.n2699 99.5127
R4213 VDD.n2696 VDD.n2695 99.5127
R4214 VDD.n2692 VDD.n2691 99.5127
R4215 VDD.n2688 VDD.n2687 99.5127
R4216 VDD.n2684 VDD.n2683 99.5127
R4217 VDD.n2680 VDD.n2679 99.5127
R4218 VDD.n2675 VDD.n2674 99.5127
R4219 VDD.n2671 VDD.n641 99.5127
R4220 VDD.n2394 VDD.n932 99.5127
R4221 VDD.n2394 VDD.n927 99.5127
R4222 VDD.n2391 VDD.n927 99.5127
R4223 VDD.n2391 VDD.n921 99.5127
R4224 VDD.n2388 VDD.n921 99.5127
R4225 VDD.n2388 VDD.n915 99.5127
R4226 VDD.n2385 VDD.n915 99.5127
R4227 VDD.n2385 VDD.n909 99.5127
R4228 VDD.n2382 VDD.n909 99.5127
R4229 VDD.n2382 VDD.n902 99.5127
R4230 VDD.n2379 VDD.n902 99.5127
R4231 VDD.n2379 VDD.n896 99.5127
R4232 VDD.n2376 VDD.n896 99.5127
R4233 VDD.n2376 VDD.n891 99.5127
R4234 VDD.n2373 VDD.n891 99.5127
R4235 VDD.n2373 VDD.n885 99.5127
R4236 VDD.n2370 VDD.n885 99.5127
R4237 VDD.n2370 VDD.n879 99.5127
R4238 VDD.n2367 VDD.n879 99.5127
R4239 VDD.n2367 VDD.n873 99.5127
R4240 VDD.n2364 VDD.n873 99.5127
R4241 VDD.n2364 VDD.n867 99.5127
R4242 VDD.n2361 VDD.n867 99.5127
R4243 VDD.n2361 VDD.n861 99.5127
R4244 VDD.n2358 VDD.n861 99.5127
R4245 VDD.n2358 VDD.n855 99.5127
R4246 VDD.n1044 VDD.n855 99.5127
R4247 VDD.n1044 VDD.n850 99.5127
R4248 VDD.n1041 VDD.n850 99.5127
R4249 VDD.n1041 VDD.n844 99.5127
R4250 VDD.n1038 VDD.n844 99.5127
R4251 VDD.n1038 VDD.n838 99.5127
R4252 VDD.n1035 VDD.n838 99.5127
R4253 VDD.n1035 VDD.n832 99.5127
R4254 VDD.n1032 VDD.n832 99.5127
R4255 VDD.n1032 VDD.n826 99.5127
R4256 VDD.n1029 VDD.n826 99.5127
R4257 VDD.n1029 VDD.n820 99.5127
R4258 VDD.n1026 VDD.n820 99.5127
R4259 VDD.n1026 VDD.n814 99.5127
R4260 VDD.n1023 VDD.n814 99.5127
R4261 VDD.n1023 VDD.n807 99.5127
R4262 VDD.n1020 VDD.n807 99.5127
R4263 VDD.n1020 VDD.n801 99.5127
R4264 VDD.n1017 VDD.n801 99.5127
R4265 VDD.n1017 VDD.n796 99.5127
R4266 VDD.n1014 VDD.n796 99.5127
R4267 VDD.n1014 VDD.n790 99.5127
R4268 VDD.n1011 VDD.n790 99.5127
R4269 VDD.n1011 VDD.n784 99.5127
R4270 VDD.n1008 VDD.n784 99.5127
R4271 VDD.n1008 VDD.n778 99.5127
R4272 VDD.n1005 VDD.n778 99.5127
R4273 VDD.n1005 VDD.n772 99.5127
R4274 VDD.n1002 VDD.n772 99.5127
R4275 VDD.n1002 VDD.n766 99.5127
R4276 VDD.n999 VDD.n766 99.5127
R4277 VDD.n999 VDD.n760 99.5127
R4278 VDD.n996 VDD.n760 99.5127
R4279 VDD.n996 VDD.n754 99.5127
R4280 VDD.n993 VDD.n754 99.5127
R4281 VDD.n993 VDD.n747 99.5127
R4282 VDD.n990 VDD.n747 99.5127
R4283 VDD.n990 VDD.n741 99.5127
R4284 VDD.n987 VDD.n741 99.5127
R4285 VDD.n987 VDD.n736 99.5127
R4286 VDD.n984 VDD.n736 99.5127
R4287 VDD.n984 VDD.n729 99.5127
R4288 VDD.n981 VDD.n729 99.5127
R4289 VDD.n981 VDD.n723 99.5127
R4290 VDD.n978 VDD.n723 99.5127
R4291 VDD.n978 VDD.n718 99.5127
R4292 VDD.n975 VDD.n718 99.5127
R4293 VDD.n975 VDD.n712 99.5127
R4294 VDD.n972 VDD.n712 99.5127
R4295 VDD.n972 VDD.n706 99.5127
R4296 VDD.n969 VDD.n706 99.5127
R4297 VDD.n969 VDD.n700 99.5127
R4298 VDD.n966 VDD.n700 99.5127
R4299 VDD.n966 VDD.n694 99.5127
R4300 VDD.n963 VDD.n694 99.5127
R4301 VDD.n963 VDD.n687 99.5127
R4302 VDD.n687 VDD.n678 99.5127
R4303 VDD.n2661 VDD.n678 99.5127
R4304 VDD.n2662 VDD.n2661 99.5127
R4305 VDD.n2662 VDD.n671 99.5127
R4306 VDD.n2665 VDD.n671 99.5127
R4307 VDD.n2665 VDD.n664 99.5127
R4308 VDD.n2668 VDD.n664 99.5127
R4309 VDD.n1149 VDD.n1148 99.5127
R4310 VDD.n1153 VDD.n1152 99.5127
R4311 VDD.n1157 VDD.n1156 99.5127
R4312 VDD.n1161 VDD.n1160 99.5127
R4313 VDD.n1165 VDD.n1164 99.5127
R4314 VDD.n1169 VDD.n1168 99.5127
R4315 VDD.n1191 VDD.n1190 99.5127
R4316 VDD.n1187 VDD.n1186 99.5127
R4317 VDD.n1183 VDD.n1182 99.5127
R4318 VDD.n1179 VDD.n1178 99.5127
R4319 VDD.n1174 VDD.n1173 99.5127
R4320 VDD.n2398 VDD.n959 99.5127
R4321 VDD.n2407 VDD.n928 99.5127
R4322 VDD.n2411 VDD.n928 99.5127
R4323 VDD.n2411 VDD.n918 99.5127
R4324 VDD.n2419 VDD.n918 99.5127
R4325 VDD.n2419 VDD.n916 99.5127
R4326 VDD.n2423 VDD.n916 99.5127
R4327 VDD.n2423 VDD.n906 99.5127
R4328 VDD.n2431 VDD.n906 99.5127
R4329 VDD.n2431 VDD.n904 99.5127
R4330 VDD.n2435 VDD.n904 99.5127
R4331 VDD.n2435 VDD.n894 99.5127
R4332 VDD.n2443 VDD.n894 99.5127
R4333 VDD.n2443 VDD.n892 99.5127
R4334 VDD.n2447 VDD.n892 99.5127
R4335 VDD.n2447 VDD.n882 99.5127
R4336 VDD.n2455 VDD.n882 99.5127
R4337 VDD.n2455 VDD.n880 99.5127
R4338 VDD.n2459 VDD.n880 99.5127
R4339 VDD.n2459 VDD.n870 99.5127
R4340 VDD.n2467 VDD.n870 99.5127
R4341 VDD.n2467 VDD.n868 99.5127
R4342 VDD.n2471 VDD.n868 99.5127
R4343 VDD.n2471 VDD.n858 99.5127
R4344 VDD.n2479 VDD.n858 99.5127
R4345 VDD.n2479 VDD.n856 99.5127
R4346 VDD.n2483 VDD.n856 99.5127
R4347 VDD.n2483 VDD.n847 99.5127
R4348 VDD.n2491 VDD.n847 99.5127
R4349 VDD.n2491 VDD.n845 99.5127
R4350 VDD.n2495 VDD.n845 99.5127
R4351 VDD.n2495 VDD.n835 99.5127
R4352 VDD.n2503 VDD.n835 99.5127
R4353 VDD.n2503 VDD.n833 99.5127
R4354 VDD.n2507 VDD.n833 99.5127
R4355 VDD.n2507 VDD.n823 99.5127
R4356 VDD.n2515 VDD.n823 99.5127
R4357 VDD.n2515 VDD.n821 99.5127
R4358 VDD.n2519 VDD.n821 99.5127
R4359 VDD.n2519 VDD.n811 99.5127
R4360 VDD.n2527 VDD.n811 99.5127
R4361 VDD.n2527 VDD.n809 99.5127
R4362 VDD.n2531 VDD.n809 99.5127
R4363 VDD.n2531 VDD.n799 99.5127
R4364 VDD.n2539 VDD.n799 99.5127
R4365 VDD.n2539 VDD.n797 99.5127
R4366 VDD.n2543 VDD.n797 99.5127
R4367 VDD.n2543 VDD.n787 99.5127
R4368 VDD.n2551 VDD.n787 99.5127
R4369 VDD.n2551 VDD.n785 99.5127
R4370 VDD.n2555 VDD.n785 99.5127
R4371 VDD.n2555 VDD.n775 99.5127
R4372 VDD.n2563 VDD.n775 99.5127
R4373 VDD.n2563 VDD.n773 99.5127
R4374 VDD.n2567 VDD.n773 99.5127
R4375 VDD.n2567 VDD.n763 99.5127
R4376 VDD.n2575 VDD.n763 99.5127
R4377 VDD.n2575 VDD.n761 99.5127
R4378 VDD.n2579 VDD.n761 99.5127
R4379 VDD.n2579 VDD.n751 99.5127
R4380 VDD.n2587 VDD.n751 99.5127
R4381 VDD.n2587 VDD.n749 99.5127
R4382 VDD.n2591 VDD.n749 99.5127
R4383 VDD.n2591 VDD.n739 99.5127
R4384 VDD.n2599 VDD.n739 99.5127
R4385 VDD.n2599 VDD.n737 99.5127
R4386 VDD.n2603 VDD.n737 99.5127
R4387 VDD.n2603 VDD.n726 99.5127
R4388 VDD.n2611 VDD.n726 99.5127
R4389 VDD.n2611 VDD.n724 99.5127
R4390 VDD.n2615 VDD.n724 99.5127
R4391 VDD.n2615 VDD.n715 99.5127
R4392 VDD.n2623 VDD.n715 99.5127
R4393 VDD.n2623 VDD.n713 99.5127
R4394 VDD.n2627 VDD.n713 99.5127
R4395 VDD.n2627 VDD.n703 99.5127
R4396 VDD.n2635 VDD.n703 99.5127
R4397 VDD.n2635 VDD.n701 99.5127
R4398 VDD.n2639 VDD.n701 99.5127
R4399 VDD.n2639 VDD.n691 99.5127
R4400 VDD.n2647 VDD.n691 99.5127
R4401 VDD.n2647 VDD.n688 99.5127
R4402 VDD.n2653 VDD.n688 99.5127
R4403 VDD.n2653 VDD.n689 99.5127
R4404 VDD.n689 VDD.n681 99.5127
R4405 VDD.n681 VDD.n672 99.5127
R4406 VDD.n2725 VDD.n672 99.5127
R4407 VDD.n2725 VDD.n673 99.5127
R4408 VDD.n673 VDD.n665 99.5127
R4409 VDD.n2720 VDD.n665 99.5127
R4410 VDD.n1501 VDD.t15 96.3032
R4411 VDD.n1575 VDD.t26 96.3032
R4412 VDD.n1547 VDD.t29 96.3032
R4413 VDD.n1196 VDD.t46 96.3032
R4414 VDD.n1130 VDD.t8 96.3032
R4415 VDD.n1112 VDD.t5 96.3032
R4416 VDD.n4081 VDD.t24 96.3032
R4417 VDD.n4060 VDD.t39 96.3032
R4418 VDD.n4042 VDD.t36 96.3032
R4419 VDD.n3593 VDD.t65 96.3032
R4420 VDD.n3633 VDD.t68 96.3032
R4421 VDD.n3550 VDD.t11 96.3032
R4422 VDD.n9 VDD.n7 96.0321
R4423 VDD.n2 VDD.n0 96.0321
R4424 VDD.n9 VDD.n8 94.7763
R4425 VDD.n11 VDD.n10 94.7763
R4426 VDD.n13 VDD.n12 94.7763
R4427 VDD.n6 VDD.n5 94.7763
R4428 VDD.n4 VDD.n3 94.7763
R4429 VDD.n2 VDD.n1 94.7763
R4430 VDD.n1171 VDD.t55 93.369
R4431 VDD.n676 VDD.t33 93.369
R4432 VDD.n1048 VDD.t42 93.369
R4433 VDD.n658 VDD.t20 93.369
R4434 VDD.n2846 VDD.t49 93.369
R4435 VDD.n357 VDD.t63 93.369
R4436 VDD.n2811 VDD.t52 93.369
R4437 VDD.n329 VDD.t60 93.369
R4438 VDD.n28 VDD.t112 91.1447
R4439 VDD.n22 VDD.t113 91.1447
R4440 VDD.n17 VDD.t82 91.1447
R4441 VDD.n1891 VDD.t90 91.1447
R4442 VDD.n1885 VDD.t89 91.1447
R4443 VDD.n1880 VDD.t78 91.1447
R4444 VDD.n31 VDD.t115 89.4493
R4445 VDD.n25 VDD.t114 89.4493
R4446 VDD.n20 VDD.t100 89.4493
R4447 VDD.n1894 VDD.t93 89.4493
R4448 VDD.n1888 VDD.t94 89.4493
R4449 VDD.n1883 VDD.t92 89.4493
R4450 VDD.n30 VDD.n29 76.0728
R4451 VDD.n28 VDD.n27 76.0728
R4452 VDD.n24 VDD.n23 76.0728
R4453 VDD.n22 VDD.n21 76.0728
R4454 VDD.n19 VDD.n18 76.0728
R4455 VDD.n17 VDD.n16 76.0728
R4456 VDD.n1891 VDD.n1890 76.0728
R4457 VDD.n1893 VDD.n1892 76.0728
R4458 VDD.n1885 VDD.n1884 76.0728
R4459 VDD.n1887 VDD.n1886 76.0728
R4460 VDD.n1880 VDD.n1879 76.0728
R4461 VDD.n1882 VDD.n1881 76.0728
R4462 VDD.n3175 VDD.n3174 72.8958
R4463 VDD.n3174 VDD.n2796 72.8958
R4464 VDD.n3174 VDD.n2797 72.8958
R4465 VDD.n3174 VDD.n2798 72.8958
R4466 VDD.n3174 VDD.n2799 72.8958
R4467 VDD.n3174 VDD.n2800 72.8958
R4468 VDD.n3174 VDD.n2801 72.8958
R4469 VDD.n3174 VDD.n2802 72.8958
R4470 VDD.n3174 VDD.n2803 72.8958
R4471 VDD.n3174 VDD.n2804 72.8958
R4472 VDD.n3174 VDD.n2805 72.8958
R4473 VDD.n3174 VDD.n2806 72.8958
R4474 VDD.n335 VDD.n323 72.8958
R4475 VDD.n3530 VDD.n323 72.8958
R4476 VDD.n331 VDD.n323 72.8958
R4477 VDD.n3537 VDD.n323 72.8958
R4478 VDD.n326 VDD.n323 72.8958
R4479 VDD.n3544 VDD.n323 72.8958
R4480 VDD.n323 VDD.n322 72.8958
R4481 VDD.n3441 VDD.n323 72.8958
R4482 VDD.n3437 VDD.n323 72.8958
R4483 VDD.n3448 VDD.n323 72.8958
R4484 VDD.n3434 VDD.n323 72.8958
R4485 VDD.n3455 VDD.n323 72.8958
R4486 VDD.n2400 VDD.n2399 72.8958
R4487 VDD.n2399 VDD.n936 72.8958
R4488 VDD.n2399 VDD.n937 72.8958
R4489 VDD.n2399 VDD.n938 72.8958
R4490 VDD.n2399 VDD.n939 72.8958
R4491 VDD.n2399 VDD.n940 72.8958
R4492 VDD.n2399 VDD.n941 72.8958
R4493 VDD.n2399 VDD.n942 72.8958
R4494 VDD.n2399 VDD.n943 72.8958
R4495 VDD.n2399 VDD.n944 72.8958
R4496 VDD.n2399 VDD.n945 72.8958
R4497 VDD.n2399 VDD.n946 72.8958
R4498 VDD.n2784 VDD.n642 72.8958
R4499 VDD.n2784 VDD.n643 72.8958
R4500 VDD.n2784 VDD.n644 72.8958
R4501 VDD.n2784 VDD.n645 72.8958
R4502 VDD.n2784 VDD.n646 72.8958
R4503 VDD.n2784 VDD.n647 72.8958
R4504 VDD.n2784 VDD.n648 72.8958
R4505 VDD.n2784 VDD.n649 72.8958
R4506 VDD.n2784 VDD.n650 72.8958
R4507 VDD.n2784 VDD.n651 72.8958
R4508 VDD.n2784 VDD.n652 72.8958
R4509 VDD.n2784 VDD.n653 72.8958
R4510 VDD.n3174 VDD.n3173 72.8958
R4511 VDD.n3174 VDD.n2785 72.8958
R4512 VDD.n3174 VDD.n2786 72.8958
R4513 VDD.n3174 VDD.n2787 72.8958
R4514 VDD.n3174 VDD.n2788 72.8958
R4515 VDD.n3174 VDD.n2789 72.8958
R4516 VDD.n3174 VDD.n2790 72.8958
R4517 VDD.n3174 VDD.n2791 72.8958
R4518 VDD.n3174 VDD.n2792 72.8958
R4519 VDD.n3174 VDD.n2793 72.8958
R4520 VDD.n3174 VDD.n2794 72.8958
R4521 VDD.n3174 VDD.n2795 72.8958
R4522 VDD.n3477 VDD.n323 72.8958
R4523 VDD.n3483 VDD.n323 72.8958
R4524 VDD.n359 VDD.n323 72.8958
R4525 VDD.n3490 VDD.n323 72.8958
R4526 VDD.n354 VDD.n323 72.8958
R4527 VDD.n3497 VDD.n323 72.8958
R4528 VDD.n3500 VDD.n323 72.8958
R4529 VDD.n350 VDD.n323 72.8958
R4530 VDD.n3507 VDD.n323 72.8958
R4531 VDD.n347 VDD.n323 72.8958
R4532 VDD.n3514 VDD.n323 72.8958
R4533 VDD.n3517 VDD.n323 72.8958
R4534 VDD.n2784 VDD.n640 72.8958
R4535 VDD.n2784 VDD.n639 72.8958
R4536 VDD.n2784 VDD.n638 72.8958
R4537 VDD.n2784 VDD.n637 72.8958
R4538 VDD.n2784 VDD.n636 72.8958
R4539 VDD.n2784 VDD.n635 72.8958
R4540 VDD.n2784 VDD.n634 72.8958
R4541 VDD.n2784 VDD.n633 72.8958
R4542 VDD.n2784 VDD.n632 72.8958
R4543 VDD.n2784 VDD.n631 72.8958
R4544 VDD.n2784 VDD.n630 72.8958
R4545 VDD.n2784 VDD.n629 72.8958
R4546 VDD.n2399 VDD.n947 72.8958
R4547 VDD.n2399 VDD.n948 72.8958
R4548 VDD.n2399 VDD.n949 72.8958
R4549 VDD.n2399 VDD.n950 72.8958
R4550 VDD.n2399 VDD.n951 72.8958
R4551 VDD.n2399 VDD.n952 72.8958
R4552 VDD.n2399 VDD.n953 72.8958
R4553 VDD.n2399 VDD.n954 72.8958
R4554 VDD.n2399 VDD.n955 72.8958
R4555 VDD.n2399 VDD.n956 72.8958
R4556 VDD.n2399 VDD.n957 72.8958
R4557 VDD.n2399 VDD.n958 72.8958
R4558 VDD.n1171 VDD.n1170 71.952
R4559 VDD.n676 VDD.n675 71.952
R4560 VDD.n1048 VDD.n1047 71.952
R4561 VDD.n658 VDD.n657 71.952
R4562 VDD.n2846 VDD.n2845 71.952
R4563 VDD.n357 VDD.n356 71.952
R4564 VDD.n2811 VDD.n2810 71.952
R4565 VDD.n329 VDD.n328 71.952
R4566 VDD.n1673 VDD.n1672 66.2847
R4567 VDD.n1673 VDD.n1504 66.2847
R4568 VDD.n1673 VDD.n1505 66.2847
R4569 VDD.n1673 VDD.n1506 66.2847
R4570 VDD.n1673 VDD.n1507 66.2847
R4571 VDD.n1673 VDD.n1508 66.2847
R4572 VDD.n1673 VDD.n1509 66.2847
R4573 VDD.n1673 VDD.n1510 66.2847
R4574 VDD.n1673 VDD.n1511 66.2847
R4575 VDD.n1673 VDD.n1512 66.2847
R4576 VDD.n1673 VDD.n1513 66.2847
R4577 VDD.n1673 VDD.n1514 66.2847
R4578 VDD.n1673 VDD.n1515 66.2847
R4579 VDD.n1673 VDD.n1516 66.2847
R4580 VDD.n1673 VDD.n1517 66.2847
R4581 VDD.n1673 VDD.n1518 66.2847
R4582 VDD.n1673 VDD.n1519 66.2847
R4583 VDD.n1673 VDD.n1520 66.2847
R4584 VDD.n1673 VDD.n1521 66.2847
R4585 VDD.n1673 VDD.n1522 66.2847
R4586 VDD.n1673 VDD.n1523 66.2847
R4587 VDD.n1673 VDD.n1524 66.2847
R4588 VDD.n1673 VDD.n1525 66.2847
R4589 VDD.n1674 VDD.n1673 66.2847
R4590 VDD.n2194 VDD.n1077 66.2847
R4591 VDD.n2194 VDD.n1078 66.2847
R4592 VDD.n2194 VDD.n1079 66.2847
R4593 VDD.n2194 VDD.n1080 66.2847
R4594 VDD.n2194 VDD.n1081 66.2847
R4595 VDD.n2194 VDD.n1082 66.2847
R4596 VDD.n2194 VDD.n1083 66.2847
R4597 VDD.n2194 VDD.n1084 66.2847
R4598 VDD.n2194 VDD.n1085 66.2847
R4599 VDD.n2194 VDD.n1086 66.2847
R4600 VDD.n2194 VDD.n1087 66.2847
R4601 VDD.n2194 VDD.n1088 66.2847
R4602 VDD.n2194 VDD.n1089 66.2847
R4603 VDD.n2194 VDD.n1090 66.2847
R4604 VDD.n2194 VDD.n1091 66.2847
R4605 VDD.n2194 VDD.n1092 66.2847
R4606 VDD.n2194 VDD.n1093 66.2847
R4607 VDD.n2194 VDD.n1094 66.2847
R4608 VDD.n2194 VDD.n1095 66.2847
R4609 VDD.n2194 VDD.n1096 66.2847
R4610 VDD.n2194 VDD.n1097 66.2847
R4611 VDD.n2194 VDD.n1098 66.2847
R4612 VDD.n2194 VDD.n1099 66.2847
R4613 VDD.n2194 VDD.n2193 66.2847
R4614 VDD.n3688 VDD.n3687 66.2847
R4615 VDD.n3689 VDD.n3688 66.2847
R4616 VDD.n3688 VDD.n298 66.2847
R4617 VDD.n3688 VDD.n299 66.2847
R4618 VDD.n3688 VDD.n300 66.2847
R4619 VDD.n3688 VDD.n301 66.2847
R4620 VDD.n3688 VDD.n302 66.2847
R4621 VDD.n3688 VDD.n303 66.2847
R4622 VDD.n3688 VDD.n304 66.2847
R4623 VDD.n3688 VDD.n305 66.2847
R4624 VDD.n3688 VDD.n306 66.2847
R4625 VDD.n3688 VDD.n307 66.2847
R4626 VDD.n3688 VDD.n308 66.2847
R4627 VDD.n3688 VDD.n309 66.2847
R4628 VDD.n3688 VDD.n310 66.2847
R4629 VDD.n3688 VDD.n311 66.2847
R4630 VDD.n3688 VDD.n312 66.2847
R4631 VDD.n3688 VDD.n313 66.2847
R4632 VDD.n3688 VDD.n314 66.2847
R4633 VDD.n3688 VDD.n315 66.2847
R4634 VDD.n3688 VDD.n316 66.2847
R4635 VDD.n3688 VDD.n317 66.2847
R4636 VDD.n3688 VDD.n318 66.2847
R4637 VDD.n3688 VDD.n3681 66.2847
R4638 VDD.n4222 VDD.n4002 66.2847
R4639 VDD.n4222 VDD.n4003 66.2847
R4640 VDD.n4222 VDD.n4004 66.2847
R4641 VDD.n4222 VDD.n4005 66.2847
R4642 VDD.n4222 VDD.n4006 66.2847
R4643 VDD.n4222 VDD.n4007 66.2847
R4644 VDD.n4222 VDD.n4008 66.2847
R4645 VDD.n4222 VDD.n4009 66.2847
R4646 VDD.n4222 VDD.n4010 66.2847
R4647 VDD.n4222 VDD.n4011 66.2847
R4648 VDD.n4222 VDD.n4012 66.2847
R4649 VDD.n4222 VDD.n4013 66.2847
R4650 VDD.n4222 VDD.n4014 66.2847
R4651 VDD.n4222 VDD.n4015 66.2847
R4652 VDD.n4222 VDD.n4016 66.2847
R4653 VDD.n4222 VDD.n4017 66.2847
R4654 VDD.n4222 VDD.n4018 66.2847
R4655 VDD.n4222 VDD.n4019 66.2847
R4656 VDD.n4222 VDD.n4020 66.2847
R4657 VDD.n4222 VDD.n4021 66.2847
R4658 VDD.n4222 VDD.n4022 66.2847
R4659 VDD.n4222 VDD.n4023 66.2847
R4660 VDD.n4222 VDD.n4024 66.2847
R4661 VDD.n4222 VDD.n4025 66.2847
R4662 VDD.n4213 VDD.n4025 52.4337
R4663 VDD.n4211 VDD.n4024 52.4337
R4664 VDD.n4207 VDD.n4023 52.4337
R4665 VDD.n4203 VDD.n4022 52.4337
R4666 VDD.n4199 VDD.n4021 52.4337
R4667 VDD.n4195 VDD.n4020 52.4337
R4668 VDD.n4044 VDD.n4019 52.4337
R4669 VDD.n4187 VDD.n4018 52.4337
R4670 VDD.n4183 VDD.n4017 52.4337
R4671 VDD.n4179 VDD.n4016 52.4337
R4672 VDD.n4175 VDD.n4015 52.4337
R4673 VDD.n4171 VDD.n4014 52.4337
R4674 VDD.n4167 VDD.n4013 52.4337
R4675 VDD.n4163 VDD.n4012 52.4337
R4676 VDD.n4159 VDD.n4011 52.4337
R4677 VDD.n4155 VDD.n4010 52.4337
R4678 VDD.n4151 VDD.n4009 52.4337
R4679 VDD.n4147 VDD.n4008 52.4337
R4680 VDD.n4143 VDD.n4007 52.4337
R4681 VDD.n4139 VDD.n4006 52.4337
R4682 VDD.n4135 VDD.n4005 52.4337
R4683 VDD.n4131 VDD.n4004 52.4337
R4684 VDD.n4127 VDD.n4003 52.4337
R4685 VDD.n4078 VDD.n4002 52.4337
R4686 VDD.n3687 VDD.n3686 52.4337
R4687 VDD.n3689 VDD.n297 52.4337
R4688 VDD.n298 VDD.n296 52.4337
R4689 VDD.n3570 VDD.n299 52.4337
R4690 VDD.n3578 VDD.n300 52.4337
R4691 VDD.n3580 VDD.n301 52.4337
R4692 VDD.n3588 VDD.n302 52.4337
R4693 VDD.n3590 VDD.n303 52.4337
R4694 VDD.n3600 VDD.n304 52.4337
R4695 VDD.n3602 VDD.n305 52.4337
R4696 VDD.n3610 VDD.n306 52.4337
R4697 VDD.n3612 VDD.n307 52.4337
R4698 VDD.n3620 VDD.n308 52.4337
R4699 VDD.n3622 VDD.n309 52.4337
R4700 VDD.n3630 VDD.n310 52.4337
R4701 VDD.n3635 VDD.n311 52.4337
R4702 VDD.n3643 VDD.n312 52.4337
R4703 VDD.n3645 VDD.n313 52.4337
R4704 VDD.n3653 VDD.n314 52.4337
R4705 VDD.n3655 VDD.n315 52.4337
R4706 VDD.n3663 VDD.n316 52.4337
R4707 VDD.n3665 VDD.n317 52.4337
R4708 VDD.n3673 VDD.n318 52.4337
R4709 VDD.n3681 VDD.n319 52.4337
R4710 VDD.n2193 VDD.n2192 52.4337
R4711 VDD.n2186 VDD.n1099 52.4337
R4712 VDD.n2182 VDD.n1098 52.4337
R4713 VDD.n2178 VDD.n1097 52.4337
R4714 VDD.n2174 VDD.n1096 52.4337
R4715 VDD.n2170 VDD.n1095 52.4337
R4716 VDD.n1114 VDD.n1094 52.4337
R4717 VDD.n2162 VDD.n1093 52.4337
R4718 VDD.n2158 VDD.n1092 52.4337
R4719 VDD.n2154 VDD.n1091 52.4337
R4720 VDD.n2150 VDD.n1090 52.4337
R4721 VDD.n2146 VDD.n1089 52.4337
R4722 VDD.n2142 VDD.n1088 52.4337
R4723 VDD.n2138 VDD.n1087 52.4337
R4724 VDD.n2134 VDD.n1086 52.4337
R4725 VDD.n2130 VDD.n1085 52.4337
R4726 VDD.n2126 VDD.n1084 52.4337
R4727 VDD.n2122 VDD.n1083 52.4337
R4728 VDD.n2118 VDD.n1082 52.4337
R4729 VDD.n2114 VDD.n1081 52.4337
R4730 VDD.n2110 VDD.n1080 52.4337
R4731 VDD.n2106 VDD.n1079 52.4337
R4732 VDD.n1197 VDD.n1078 52.4337
R4733 VDD.n1194 VDD.n1077 52.4337
R4734 VDD.n1672 VDD.n1671 52.4337
R4735 VDD.n1531 VDD.n1504 52.4337
R4736 VDD.n1533 VDD.n1505 52.4337
R4737 VDD.n1537 VDD.n1506 52.4337
R4738 VDD.n1539 VDD.n1507 52.4337
R4739 VDD.n1543 VDD.n1508 52.4337
R4740 VDD.n1545 VDD.n1509 52.4337
R4741 VDD.n1551 VDD.n1510 52.4337
R4742 VDD.n1553 VDD.n1511 52.4337
R4743 VDD.n1557 VDD.n1512 52.4337
R4744 VDD.n1559 VDD.n1513 52.4337
R4745 VDD.n1563 VDD.n1514 52.4337
R4746 VDD.n1565 VDD.n1515 52.4337
R4747 VDD.n1569 VDD.n1516 52.4337
R4748 VDD.n1571 VDD.n1517 52.4337
R4749 VDD.n1578 VDD.n1518 52.4337
R4750 VDD.n1580 VDD.n1519 52.4337
R4751 VDD.n1584 VDD.n1520 52.4337
R4752 VDD.n1586 VDD.n1521 52.4337
R4753 VDD.n1590 VDD.n1522 52.4337
R4754 VDD.n1592 VDD.n1523 52.4337
R4755 VDD.n1596 VDD.n1524 52.4337
R4756 VDD.n1598 VDD.n1525 52.4337
R4757 VDD.n1674 VDD.n1503 52.4337
R4758 VDD.n1672 VDD.n1527 52.4337
R4759 VDD.n1532 VDD.n1504 52.4337
R4760 VDD.n1536 VDD.n1505 52.4337
R4761 VDD.n1538 VDD.n1506 52.4337
R4762 VDD.n1542 VDD.n1507 52.4337
R4763 VDD.n1544 VDD.n1508 52.4337
R4764 VDD.n1550 VDD.n1509 52.4337
R4765 VDD.n1552 VDD.n1510 52.4337
R4766 VDD.n1556 VDD.n1511 52.4337
R4767 VDD.n1558 VDD.n1512 52.4337
R4768 VDD.n1562 VDD.n1513 52.4337
R4769 VDD.n1564 VDD.n1514 52.4337
R4770 VDD.n1568 VDD.n1515 52.4337
R4771 VDD.n1570 VDD.n1516 52.4337
R4772 VDD.n1577 VDD.n1517 52.4337
R4773 VDD.n1579 VDD.n1518 52.4337
R4774 VDD.n1583 VDD.n1519 52.4337
R4775 VDD.n1585 VDD.n1520 52.4337
R4776 VDD.n1589 VDD.n1521 52.4337
R4777 VDD.n1591 VDD.n1522 52.4337
R4778 VDD.n1595 VDD.n1523 52.4337
R4779 VDD.n1597 VDD.n1524 52.4337
R4780 VDD.n1599 VDD.n1525 52.4337
R4781 VDD.n1675 VDD.n1674 52.4337
R4782 VDD.n1198 VDD.n1077 52.4337
R4783 VDD.n2105 VDD.n1078 52.4337
R4784 VDD.n2109 VDD.n1079 52.4337
R4785 VDD.n2113 VDD.n1080 52.4337
R4786 VDD.n2117 VDD.n1081 52.4337
R4787 VDD.n2121 VDD.n1082 52.4337
R4788 VDD.n2125 VDD.n1083 52.4337
R4789 VDD.n2129 VDD.n1084 52.4337
R4790 VDD.n2133 VDD.n1085 52.4337
R4791 VDD.n2137 VDD.n1086 52.4337
R4792 VDD.n2141 VDD.n1087 52.4337
R4793 VDD.n2145 VDD.n1088 52.4337
R4794 VDD.n2149 VDD.n1089 52.4337
R4795 VDD.n2153 VDD.n1090 52.4337
R4796 VDD.n2157 VDD.n1091 52.4337
R4797 VDD.n2161 VDD.n1092 52.4337
R4798 VDD.n1113 VDD.n1093 52.4337
R4799 VDD.n2169 VDD.n1094 52.4337
R4800 VDD.n2173 VDD.n1095 52.4337
R4801 VDD.n2177 VDD.n1096 52.4337
R4802 VDD.n2181 VDD.n1097 52.4337
R4803 VDD.n2185 VDD.n1098 52.4337
R4804 VDD.n2189 VDD.n1099 52.4337
R4805 VDD.n2193 VDD.n1100 52.4337
R4806 VDD.n3687 VDD.n3685 52.4337
R4807 VDD.n3690 VDD.n3689 52.4337
R4808 VDD.n3571 VDD.n298 52.4337
R4809 VDD.n3577 VDD.n299 52.4337
R4810 VDD.n3581 VDD.n300 52.4337
R4811 VDD.n3587 VDD.n301 52.4337
R4812 VDD.n3591 VDD.n302 52.4337
R4813 VDD.n3599 VDD.n303 52.4337
R4814 VDD.n3603 VDD.n304 52.4337
R4815 VDD.n3609 VDD.n305 52.4337
R4816 VDD.n3613 VDD.n306 52.4337
R4817 VDD.n3619 VDD.n307 52.4337
R4818 VDD.n3623 VDD.n308 52.4337
R4819 VDD.n3629 VDD.n309 52.4337
R4820 VDD.n3636 VDD.n310 52.4337
R4821 VDD.n3642 VDD.n311 52.4337
R4822 VDD.n3646 VDD.n312 52.4337
R4823 VDD.n3652 VDD.n313 52.4337
R4824 VDD.n3656 VDD.n314 52.4337
R4825 VDD.n3662 VDD.n315 52.4337
R4826 VDD.n3666 VDD.n316 52.4337
R4827 VDD.n3672 VDD.n317 52.4337
R4828 VDD.n3676 VDD.n318 52.4337
R4829 VDD.n3681 VDD.n3680 52.4337
R4830 VDD.n4126 VDD.n4002 52.4337
R4831 VDD.n4130 VDD.n4003 52.4337
R4832 VDD.n4134 VDD.n4004 52.4337
R4833 VDD.n4138 VDD.n4005 52.4337
R4834 VDD.n4142 VDD.n4006 52.4337
R4835 VDD.n4146 VDD.n4007 52.4337
R4836 VDD.n4150 VDD.n4008 52.4337
R4837 VDD.n4154 VDD.n4009 52.4337
R4838 VDD.n4158 VDD.n4010 52.4337
R4839 VDD.n4162 VDD.n4011 52.4337
R4840 VDD.n4166 VDD.n4012 52.4337
R4841 VDD.n4170 VDD.n4013 52.4337
R4842 VDD.n4174 VDD.n4014 52.4337
R4843 VDD.n4178 VDD.n4015 52.4337
R4844 VDD.n4182 VDD.n4016 52.4337
R4845 VDD.n4186 VDD.n4017 52.4337
R4846 VDD.n4043 VDD.n4018 52.4337
R4847 VDD.n4194 VDD.n4019 52.4337
R4848 VDD.n4198 VDD.n4020 52.4337
R4849 VDD.n4202 VDD.n4021 52.4337
R4850 VDD.n4206 VDD.n4022 52.4337
R4851 VDD.n4210 VDD.n4023 52.4337
R4852 VDD.n4214 VDD.n4024 52.4337
R4853 VDD.n4026 VDD.n4025 52.4337
R4854 VDD.n3517 VDD.n3516 39.2114
R4855 VDD.n3514 VDD.n3513 39.2114
R4856 VDD.n3509 VDD.n347 39.2114
R4857 VDD.n3507 VDD.n3506 39.2114
R4858 VDD.n3502 VDD.n350 39.2114
R4859 VDD.n3500 VDD.n3499 39.2114
R4860 VDD.n3497 VDD.n3496 39.2114
R4861 VDD.n3492 VDD.n354 39.2114
R4862 VDD.n3490 VDD.n3489 39.2114
R4863 VDD.n3485 VDD.n359 39.2114
R4864 VDD.n3483 VDD.n3482 39.2114
R4865 VDD.n3478 VDD.n3477 39.2114
R4866 VDD.n3173 VDD.n3172 39.2114
R4867 VDD.n3167 VDD.n2785 39.2114
R4868 VDD.n3164 VDD.n2786 39.2114
R4869 VDD.n3160 VDD.n2787 39.2114
R4870 VDD.n3156 VDD.n2788 39.2114
R4871 VDD.n3152 VDD.n2789 39.2114
R4872 VDD.n3148 VDD.n2790 39.2114
R4873 VDD.n3144 VDD.n2791 39.2114
R4874 VDD.n3140 VDD.n2792 39.2114
R4875 VDD.n3136 VDD.n2793 39.2114
R4876 VDD.n3132 VDD.n2794 39.2114
R4877 VDD.n3128 VDD.n2795 39.2114
R4878 VDD.n2779 VDD.n653 39.2114
R4879 VDD.n2775 VDD.n652 39.2114
R4880 VDD.n2771 VDD.n651 39.2114
R4881 VDD.n2767 VDD.n650 39.2114
R4882 VDD.n2763 VDD.n649 39.2114
R4883 VDD.n2759 VDD.n648 39.2114
R4884 VDD.n2755 VDD.n647 39.2114
R4885 VDD.n2751 VDD.n646 39.2114
R4886 VDD.n2747 VDD.n645 39.2114
R4887 VDD.n2743 VDD.n644 39.2114
R4888 VDD.n2739 VDD.n643 39.2114
R4889 VDD.n2735 VDD.n642 39.2114
R4890 VDD.n2400 VDD.n933 39.2114
R4891 VDD.n1050 VDD.n936 39.2114
R4892 VDD.n1054 VDD.n937 39.2114
R4893 VDD.n1058 VDD.n938 39.2114
R4894 VDD.n1062 VDD.n939 39.2114
R4895 VDD.n1066 VDD.n940 39.2114
R4896 VDD.n2202 VDD.n941 39.2114
R4897 VDD.n2206 VDD.n942 39.2114
R4898 VDD.n2210 VDD.n943 39.2114
R4899 VDD.n2214 VDD.n944 39.2114
R4900 VDD.n2218 VDD.n945 39.2114
R4901 VDD.n2222 VDD.n946 39.2114
R4902 VDD.n3455 VDD.n3454 39.2114
R4903 VDD.n3450 VDD.n3434 39.2114
R4904 VDD.n3448 VDD.n3447 39.2114
R4905 VDD.n3443 VDD.n3437 39.2114
R4906 VDD.n3441 VDD.n3440 39.2114
R4907 VDD.n3546 VDD.n322 39.2114
R4908 VDD.n3544 VDD.n3543 39.2114
R4909 VDD.n3539 VDD.n326 39.2114
R4910 VDD.n3537 VDD.n3536 39.2114
R4911 VDD.n3532 VDD.n331 39.2114
R4912 VDD.n3530 VDD.n3529 39.2114
R4913 VDD.n3525 VDD.n335 39.2114
R4914 VDD.n3176 VDD.n3175 39.2114
R4915 VDD.n2847 VDD.n2796 39.2114
R4916 VDD.n2851 VDD.n2797 39.2114
R4917 VDD.n2855 VDD.n2798 39.2114
R4918 VDD.n2859 VDD.n2799 39.2114
R4919 VDD.n2863 VDD.n2800 39.2114
R4920 VDD.n2867 VDD.n2801 39.2114
R4921 VDD.n2871 VDD.n2802 39.2114
R4922 VDD.n2875 VDD.n2803 39.2114
R4923 VDD.n2879 VDD.n2804 39.2114
R4924 VDD.n2883 VDD.n2805 39.2114
R4925 VDD.n2888 VDD.n2806 39.2114
R4926 VDD.n3175 VDD.n627 39.2114
R4927 VDD.n2850 VDD.n2796 39.2114
R4928 VDD.n2854 VDD.n2797 39.2114
R4929 VDD.n2858 VDD.n2798 39.2114
R4930 VDD.n2862 VDD.n2799 39.2114
R4931 VDD.n2866 VDD.n2800 39.2114
R4932 VDD.n2870 VDD.n2801 39.2114
R4933 VDD.n2874 VDD.n2802 39.2114
R4934 VDD.n2878 VDD.n2803 39.2114
R4935 VDD.n2882 VDD.n2804 39.2114
R4936 VDD.n2887 VDD.n2805 39.2114
R4937 VDD.n2890 VDD.n2806 39.2114
R4938 VDD.n335 VDD.n333 39.2114
R4939 VDD.n3531 VDD.n3530 39.2114
R4940 VDD.n331 VDD.n327 39.2114
R4941 VDD.n3538 VDD.n3537 39.2114
R4942 VDD.n326 VDD.n324 39.2114
R4943 VDD.n3545 VDD.n3544 39.2114
R4944 VDD.n3438 VDD.n322 39.2114
R4945 VDD.n3442 VDD.n3441 39.2114
R4946 VDD.n3437 VDD.n3435 39.2114
R4947 VDD.n3449 VDD.n3448 39.2114
R4948 VDD.n3434 VDD.n3432 39.2114
R4949 VDD.n3456 VDD.n3455 39.2114
R4950 VDD.n2401 VDD.n2400 39.2114
R4951 VDD.n1053 VDD.n936 39.2114
R4952 VDD.n1057 VDD.n937 39.2114
R4953 VDD.n1061 VDD.n938 39.2114
R4954 VDD.n1065 VDD.n939 39.2114
R4955 VDD.n2201 VDD.n940 39.2114
R4956 VDD.n2205 VDD.n941 39.2114
R4957 VDD.n2209 VDD.n942 39.2114
R4958 VDD.n2213 VDD.n943 39.2114
R4959 VDD.n2217 VDD.n944 39.2114
R4960 VDD.n2221 VDD.n945 39.2114
R4961 VDD.n2224 VDD.n946 39.2114
R4962 VDD.n2738 VDD.n642 39.2114
R4963 VDD.n2742 VDD.n643 39.2114
R4964 VDD.n2746 VDD.n644 39.2114
R4965 VDD.n2750 VDD.n645 39.2114
R4966 VDD.n2754 VDD.n646 39.2114
R4967 VDD.n2758 VDD.n647 39.2114
R4968 VDD.n2762 VDD.n648 39.2114
R4969 VDD.n2766 VDD.n649 39.2114
R4970 VDD.n2770 VDD.n650 39.2114
R4971 VDD.n2774 VDD.n651 39.2114
R4972 VDD.n2778 VDD.n652 39.2114
R4973 VDD.n655 VDD.n653 39.2114
R4974 VDD.n3173 VDD.n2809 39.2114
R4975 VDD.n3165 VDD.n2785 39.2114
R4976 VDD.n3161 VDD.n2786 39.2114
R4977 VDD.n3157 VDD.n2787 39.2114
R4978 VDD.n3153 VDD.n2788 39.2114
R4979 VDD.n3149 VDD.n2789 39.2114
R4980 VDD.n3145 VDD.n2790 39.2114
R4981 VDD.n3141 VDD.n2791 39.2114
R4982 VDD.n3137 VDD.n2792 39.2114
R4983 VDD.n3133 VDD.n2793 39.2114
R4984 VDD.n3129 VDD.n2794 39.2114
R4985 VDD.n3125 VDD.n2795 39.2114
R4986 VDD.n3477 VDD.n361 39.2114
R4987 VDD.n3484 VDD.n3483 39.2114
R4988 VDD.n359 VDD.n355 39.2114
R4989 VDD.n3491 VDD.n3490 39.2114
R4990 VDD.n354 VDD.n352 39.2114
R4991 VDD.n3498 VDD.n3497 39.2114
R4992 VDD.n3501 VDD.n3500 39.2114
R4993 VDD.n350 VDD.n348 39.2114
R4994 VDD.n3508 VDD.n3507 39.2114
R4995 VDD.n347 VDD.n345 39.2114
R4996 VDD.n3515 VDD.n3514 39.2114
R4997 VDD.n3518 VDD.n3517 39.2114
R4998 VDD.n2719 VDD.n629 39.2114
R4999 VDD.n2715 VDD.n630 39.2114
R5000 VDD.n2711 VDD.n631 39.2114
R5001 VDD.n2707 VDD.n632 39.2114
R5002 VDD.n2703 VDD.n633 39.2114
R5003 VDD.n2699 VDD.n634 39.2114
R5004 VDD.n2695 VDD.n635 39.2114
R5005 VDD.n2691 VDD.n636 39.2114
R5006 VDD.n2687 VDD.n637 39.2114
R5007 VDD.n2683 VDD.n638 39.2114
R5008 VDD.n2679 VDD.n639 39.2114
R5009 VDD.n2674 VDD.n640 39.2114
R5010 VDD.n947 VDD.n930 39.2114
R5011 VDD.n1149 VDD.n948 39.2114
R5012 VDD.n1153 VDD.n949 39.2114
R5013 VDD.n1157 VDD.n950 39.2114
R5014 VDD.n1161 VDD.n951 39.2114
R5015 VDD.n1165 VDD.n952 39.2114
R5016 VDD.n1169 VDD.n953 39.2114
R5017 VDD.n1190 VDD.n954 39.2114
R5018 VDD.n1186 VDD.n955 39.2114
R5019 VDD.n1182 VDD.n956 39.2114
R5020 VDD.n1178 VDD.n957 39.2114
R5021 VDD.n1173 VDD.n958 39.2114
R5022 VDD.n2671 VDD.n640 39.2114
R5023 VDD.n2675 VDD.n639 39.2114
R5024 VDD.n2680 VDD.n638 39.2114
R5025 VDD.n2684 VDD.n637 39.2114
R5026 VDD.n2688 VDD.n636 39.2114
R5027 VDD.n2692 VDD.n635 39.2114
R5028 VDD.n2696 VDD.n634 39.2114
R5029 VDD.n2700 VDD.n633 39.2114
R5030 VDD.n2704 VDD.n632 39.2114
R5031 VDD.n2708 VDD.n631 39.2114
R5032 VDD.n2712 VDD.n630 39.2114
R5033 VDD.n2716 VDD.n629 39.2114
R5034 VDD.n1148 VDD.n947 39.2114
R5035 VDD.n1152 VDD.n948 39.2114
R5036 VDD.n1156 VDD.n949 39.2114
R5037 VDD.n1160 VDD.n950 39.2114
R5038 VDD.n1164 VDD.n951 39.2114
R5039 VDD.n1168 VDD.n952 39.2114
R5040 VDD.n1191 VDD.n953 39.2114
R5041 VDD.n1187 VDD.n954 39.2114
R5042 VDD.n1183 VDD.n955 39.2114
R5043 VDD.n1179 VDD.n956 39.2114
R5044 VDD.n1174 VDD.n957 39.2114
R5045 VDD.n959 VDD.n958 39.2114
R5046 VDD.n2404 VDD.n2403 31.0639
R5047 VDD.n2782 VDD.n656 31.0639
R5048 VDD.n2736 VDD.n660 31.0639
R5049 VDD.n2226 VDD.n2225 31.0639
R5050 VDD.n3126 VDD.n3123 31.0639
R5051 VDD.n3479 VDD.n3476 31.0639
R5052 VDD.n3171 VDD.n620 31.0639
R5053 VDD.n3521 VDD.n3520 31.0639
R5054 VDD.n3459 VDD.n3458 31.0639
R5055 VDD.n3526 VDD.n334 31.0639
R5056 VDD.n2894 VDD.n2892 31.0639
R5057 VDD.n3178 VDD.n3177 31.0639
R5058 VDD.n2408 VDD.n929 31.0639
R5059 VDD.n2721 VDD.n2718 31.0639
R5060 VDD.n2670 VDD.n2669 31.0639
R5061 VDD.n2397 VDD.n2396 31.0639
R5062 VDD.n1502 VDD.n1501 30.8369
R5063 VDD.n1576 VDD.n1575 30.8369
R5064 VDD.n1548 VDD.n1547 30.8369
R5065 VDD.n1199 VDD.n1196 30.8369
R5066 VDD.n1131 VDD.n1130 30.8369
R5067 VDD.n2167 VDD.n1112 30.8369
R5068 VDD.n4125 VDD.n4081 30.8369
R5069 VDD.n4061 VDD.n4060 30.8369
R5070 VDD.n4192 VDD.n4042 30.8369
R5071 VDD.n3594 VDD.n3593 30.8369
R5072 VDD.n3634 VDD.n3633 30.8369
R5073 VDD.n3678 VDD.n3550 30.8369
R5074 VDD.n1673 VDD.n1496 25.5796
R5075 VDD.n2195 VDD.n2194 25.5796
R5076 VDD.n3688 VDD.n287 25.5796
R5077 VDD.n4223 VDD.n4222 25.5796
R5078 VDD.n1176 VDD.n1171 24.049
R5079 VDD.n2677 VDD.n676 24.049
R5080 VDD.n1049 VDD.n1048 24.049
R5081 VDD.n659 VDD.n658 24.049
R5082 VDD.n2885 VDD.n2846 24.049
R5083 VDD.n358 VDD.n357 24.049
R5084 VDD.n2812 VDD.n2811 24.049
R5085 VDD.n330 VDD.n329 24.049
R5086 VDD.n1680 VDD.n1498 19.3944
R5087 VDD.n1680 VDD.n1488 19.3944
R5088 VDD.n1692 VDD.n1488 19.3944
R5089 VDD.n1692 VDD.n1486 19.3944
R5090 VDD.n1696 VDD.n1486 19.3944
R5091 VDD.n1696 VDD.n1477 19.3944
R5092 VDD.n1709 VDD.n1477 19.3944
R5093 VDD.n1709 VDD.n1475 19.3944
R5094 VDD.n1713 VDD.n1475 19.3944
R5095 VDD.n1713 VDD.n1465 19.3944
R5096 VDD.n1725 VDD.n1465 19.3944
R5097 VDD.n1725 VDD.n1463 19.3944
R5098 VDD.n1729 VDD.n1463 19.3944
R5099 VDD.n1729 VDD.n1453 19.3944
R5100 VDD.n1741 VDD.n1453 19.3944
R5101 VDD.n1741 VDD.n1451 19.3944
R5102 VDD.n1745 VDD.n1451 19.3944
R5103 VDD.n1745 VDD.n1441 19.3944
R5104 VDD.n1757 VDD.n1441 19.3944
R5105 VDD.n1757 VDD.n1439 19.3944
R5106 VDD.n1761 VDD.n1439 19.3944
R5107 VDD.n1761 VDD.n1429 19.3944
R5108 VDD.n1772 VDD.n1429 19.3944
R5109 VDD.n1772 VDD.n1427 19.3944
R5110 VDD.n1776 VDD.n1427 19.3944
R5111 VDD.n1776 VDD.n1417 19.3944
R5112 VDD.n1788 VDD.n1417 19.3944
R5113 VDD.n1788 VDD.n1415 19.3944
R5114 VDD.n1792 VDD.n1415 19.3944
R5115 VDD.n1792 VDD.n1404 19.3944
R5116 VDD.n1804 VDD.n1404 19.3944
R5117 VDD.n1804 VDD.n1402 19.3944
R5118 VDD.n1808 VDD.n1402 19.3944
R5119 VDD.n1808 VDD.n1393 19.3944
R5120 VDD.n1820 VDD.n1393 19.3944
R5121 VDD.n1820 VDD.n1391 19.3944
R5122 VDD.n1824 VDD.n1391 19.3944
R5123 VDD.n1824 VDD.n1381 19.3944
R5124 VDD.n1836 VDD.n1381 19.3944
R5125 VDD.n1836 VDD.n1379 19.3944
R5126 VDD.n1840 VDD.n1379 19.3944
R5127 VDD.n1840 VDD.n1368 19.3944
R5128 VDD.n1852 VDD.n1368 19.3944
R5129 VDD.n1852 VDD.n1366 19.3944
R5130 VDD.n1856 VDD.n1366 19.3944
R5131 VDD.n1856 VDD.n1357 19.3944
R5132 VDD.n1868 VDD.n1357 19.3944
R5133 VDD.n1868 VDD.n1355 19.3944
R5134 VDD.n1872 VDD.n1355 19.3944
R5135 VDD.n1872 VDD.n1345 19.3944
R5136 VDD.n1903 VDD.n1345 19.3944
R5137 VDD.n1903 VDD.n1343 19.3944
R5138 VDD.n1907 VDD.n1343 19.3944
R5139 VDD.n1907 VDD.n1332 19.3944
R5140 VDD.n1919 VDD.n1332 19.3944
R5141 VDD.n1919 VDD.n1330 19.3944
R5142 VDD.n1923 VDD.n1330 19.3944
R5143 VDD.n1923 VDD.n1321 19.3944
R5144 VDD.n1935 VDD.n1321 19.3944
R5145 VDD.n1935 VDD.n1319 19.3944
R5146 VDD.n1939 VDD.n1319 19.3944
R5147 VDD.n1939 VDD.n1309 19.3944
R5148 VDD.n1951 VDD.n1309 19.3944
R5149 VDD.n1951 VDD.n1307 19.3944
R5150 VDD.n1955 VDD.n1307 19.3944
R5151 VDD.n1955 VDD.n1296 19.3944
R5152 VDD.n1967 VDD.n1296 19.3944
R5153 VDD.n1967 VDD.n1294 19.3944
R5154 VDD.n1971 VDD.n1294 19.3944
R5155 VDD.n1971 VDD.n1285 19.3944
R5156 VDD.n1983 VDD.n1285 19.3944
R5157 VDD.n1983 VDD.n1283 19.3944
R5158 VDD.n1987 VDD.n1283 19.3944
R5159 VDD.n1987 VDD.n1273 19.3944
R5160 VDD.n1999 VDD.n1273 19.3944
R5161 VDD.n1999 VDD.n1271 19.3944
R5162 VDD.n2003 VDD.n1271 19.3944
R5163 VDD.n2003 VDD.n1261 19.3944
R5164 VDD.n2015 VDD.n1261 19.3944
R5165 VDD.n2015 VDD.n1259 19.3944
R5166 VDD.n2019 VDD.n1259 19.3944
R5167 VDD.n2019 VDD.n1250 19.3944
R5168 VDD.n2031 VDD.n1250 19.3944
R5169 VDD.n2031 VDD.n1248 19.3944
R5170 VDD.n2035 VDD.n1248 19.3944
R5171 VDD.n2035 VDD.n1238 19.3944
R5172 VDD.n2047 VDD.n1238 19.3944
R5173 VDD.n2047 VDD.n1236 19.3944
R5174 VDD.n2051 VDD.n1236 19.3944
R5175 VDD.n2051 VDD.n1226 19.3944
R5176 VDD.n2063 VDD.n1226 19.3944
R5177 VDD.n2063 VDD.n1224 19.3944
R5178 VDD.n2067 VDD.n1224 19.3944
R5179 VDD.n2067 VDD.n1215 19.3944
R5180 VDD.n2080 VDD.n1215 19.3944
R5181 VDD.n2080 VDD.n1212 19.3944
R5182 VDD.n2086 VDD.n1212 19.3944
R5183 VDD.n2086 VDD.n1213 19.3944
R5184 VDD.n1213 VDD.n1202 19.3944
R5185 VDD.n2099 VDD.n1202 19.3944
R5186 VDD.n2100 VDD.n2099 19.3944
R5187 VDD.n1623 VDD.n1622 19.3944
R5188 VDD.n1622 VDD.n1621 19.3944
R5189 VDD.n1621 VDD.n1581 19.3944
R5190 VDD.n1617 VDD.n1581 19.3944
R5191 VDD.n1617 VDD.n1616 19.3944
R5192 VDD.n1616 VDD.n1615 19.3944
R5193 VDD.n1615 VDD.n1587 19.3944
R5194 VDD.n1611 VDD.n1587 19.3944
R5195 VDD.n1611 VDD.n1610 19.3944
R5196 VDD.n1610 VDD.n1609 19.3944
R5197 VDD.n1609 VDD.n1593 19.3944
R5198 VDD.n1605 VDD.n1593 19.3944
R5199 VDD.n1605 VDD.n1604 19.3944
R5200 VDD.n1604 VDD.n1603 19.3944
R5201 VDD.n1603 VDD.n1600 19.3944
R5202 VDD.n1647 VDD.n1646 19.3944
R5203 VDD.n1646 VDD.n1645 19.3944
R5204 VDD.n1645 VDD.n1554 19.3944
R5205 VDD.n1641 VDD.n1554 19.3944
R5206 VDD.n1641 VDD.n1640 19.3944
R5207 VDD.n1640 VDD.n1639 19.3944
R5208 VDD.n1639 VDD.n1560 19.3944
R5209 VDD.n1635 VDD.n1560 19.3944
R5210 VDD.n1635 VDD.n1634 19.3944
R5211 VDD.n1634 VDD.n1633 19.3944
R5212 VDD.n1633 VDD.n1566 19.3944
R5213 VDD.n1629 VDD.n1566 19.3944
R5214 VDD.n1629 VDD.n1628 19.3944
R5215 VDD.n1628 VDD.n1627 19.3944
R5216 VDD.n1627 VDD.n1572 19.3944
R5217 VDD.n1670 VDD.n1669 19.3944
R5218 VDD.n1669 VDD.n1529 19.3944
R5219 VDD.n1665 VDD.n1529 19.3944
R5220 VDD.n1665 VDD.n1664 19.3944
R5221 VDD.n1664 VDD.n1663 19.3944
R5222 VDD.n1663 VDD.n1534 19.3944
R5223 VDD.n1659 VDD.n1534 19.3944
R5224 VDD.n1659 VDD.n1658 19.3944
R5225 VDD.n1658 VDD.n1657 19.3944
R5226 VDD.n1657 VDD.n1540 19.3944
R5227 VDD.n1653 VDD.n1540 19.3944
R5228 VDD.n1653 VDD.n1652 19.3944
R5229 VDD.n1652 VDD.n1651 19.3944
R5230 VDD.n2132 VDD.n2131 19.3944
R5231 VDD.n2131 VDD.n2128 19.3944
R5232 VDD.n2128 VDD.n2127 19.3944
R5233 VDD.n2127 VDD.n2124 19.3944
R5234 VDD.n2124 VDD.n2123 19.3944
R5235 VDD.n2123 VDD.n2120 19.3944
R5236 VDD.n2120 VDD.n2119 19.3944
R5237 VDD.n2119 VDD.n2116 19.3944
R5238 VDD.n2116 VDD.n2115 19.3944
R5239 VDD.n2115 VDD.n2112 19.3944
R5240 VDD.n2112 VDD.n2111 19.3944
R5241 VDD.n2111 VDD.n2108 19.3944
R5242 VDD.n2108 VDD.n2107 19.3944
R5243 VDD.n2107 VDD.n2104 19.3944
R5244 VDD.n2163 VDD.n1110 19.3944
R5245 VDD.n2163 VDD.n2160 19.3944
R5246 VDD.n2160 VDD.n2159 19.3944
R5247 VDD.n2159 VDD.n2156 19.3944
R5248 VDD.n2156 VDD.n2155 19.3944
R5249 VDD.n2155 VDD.n2152 19.3944
R5250 VDD.n2152 VDD.n2151 19.3944
R5251 VDD.n2151 VDD.n2148 19.3944
R5252 VDD.n2148 VDD.n2147 19.3944
R5253 VDD.n2147 VDD.n2144 19.3944
R5254 VDD.n2144 VDD.n2143 19.3944
R5255 VDD.n2143 VDD.n2140 19.3944
R5256 VDD.n2140 VDD.n2139 19.3944
R5257 VDD.n2139 VDD.n2136 19.3944
R5258 VDD.n2136 VDD.n2135 19.3944
R5259 VDD.n2191 VDD.n2190 19.3944
R5260 VDD.n2188 VDD.n2187 19.3944
R5261 VDD.n2187 VDD.n2184 19.3944
R5262 VDD.n2184 VDD.n2183 19.3944
R5263 VDD.n2183 VDD.n2180 19.3944
R5264 VDD.n2180 VDD.n2179 19.3944
R5265 VDD.n2179 VDD.n2176 19.3944
R5266 VDD.n2176 VDD.n2175 19.3944
R5267 VDD.n2175 VDD.n2172 19.3944
R5268 VDD.n2172 VDD.n2171 19.3944
R5269 VDD.n2171 VDD.n2168 19.3944
R5270 VDD.n1684 VDD.n1494 19.3944
R5271 VDD.n1684 VDD.n1492 19.3944
R5272 VDD.n1688 VDD.n1492 19.3944
R5273 VDD.n1688 VDD.n1482 19.3944
R5274 VDD.n1701 VDD.n1482 19.3944
R5275 VDD.n1701 VDD.n1480 19.3944
R5276 VDD.n1705 VDD.n1480 19.3944
R5277 VDD.n1705 VDD.n1471 19.3944
R5278 VDD.n1717 VDD.n1471 19.3944
R5279 VDD.n1717 VDD.n1469 19.3944
R5280 VDD.n1721 VDD.n1469 19.3944
R5281 VDD.n1721 VDD.n1459 19.3944
R5282 VDD.n1733 VDD.n1459 19.3944
R5283 VDD.n1733 VDD.n1457 19.3944
R5284 VDD.n1737 VDD.n1457 19.3944
R5285 VDD.n1737 VDD.n1447 19.3944
R5286 VDD.n1749 VDD.n1447 19.3944
R5287 VDD.n1749 VDD.n1445 19.3944
R5288 VDD.n1753 VDD.n1445 19.3944
R5289 VDD.n1753 VDD.n1435 19.3944
R5290 VDD.n1764 VDD.n1435 19.3944
R5291 VDD.n1764 VDD.n1433 19.3944
R5292 VDD.n1768 VDD.n1433 19.3944
R5293 VDD.n1768 VDD.n1423 19.3944
R5294 VDD.n1780 VDD.n1423 19.3944
R5295 VDD.n1780 VDD.n1421 19.3944
R5296 VDD.n1784 VDD.n1421 19.3944
R5297 VDD.n1784 VDD.n1411 19.3944
R5298 VDD.n1796 VDD.n1411 19.3944
R5299 VDD.n1796 VDD.n1409 19.3944
R5300 VDD.n1800 VDD.n1409 19.3944
R5301 VDD.n1800 VDD.n1399 19.3944
R5302 VDD.n1812 VDD.n1399 19.3944
R5303 VDD.n1812 VDD.n1397 19.3944
R5304 VDD.n1816 VDD.n1397 19.3944
R5305 VDD.n1816 VDD.n1387 19.3944
R5306 VDD.n1828 VDD.n1387 19.3944
R5307 VDD.n1828 VDD.n1385 19.3944
R5308 VDD.n1832 VDD.n1385 19.3944
R5309 VDD.n1832 VDD.n1375 19.3944
R5310 VDD.n1844 VDD.n1375 19.3944
R5311 VDD.n1844 VDD.n1373 19.3944
R5312 VDD.n1848 VDD.n1373 19.3944
R5313 VDD.n1848 VDD.n1363 19.3944
R5314 VDD.n1860 VDD.n1363 19.3944
R5315 VDD.n1860 VDD.n1361 19.3944
R5316 VDD.n1864 VDD.n1361 19.3944
R5317 VDD.n1864 VDD.n1351 19.3944
R5318 VDD.n1876 VDD.n1351 19.3944
R5319 VDD.n1876 VDD.n1349 19.3944
R5320 VDD.n1899 VDD.n1349 19.3944
R5321 VDD.n1899 VDD.n1339 19.3944
R5322 VDD.n1911 VDD.n1339 19.3944
R5323 VDD.n1911 VDD.n1337 19.3944
R5324 VDD.n1915 VDD.n1337 19.3944
R5325 VDD.n1915 VDD.n1327 19.3944
R5326 VDD.n1927 VDD.n1327 19.3944
R5327 VDD.n1927 VDD.n1325 19.3944
R5328 VDD.n1931 VDD.n1325 19.3944
R5329 VDD.n1931 VDD.n1315 19.3944
R5330 VDD.n1943 VDD.n1315 19.3944
R5331 VDD.n1943 VDD.n1313 19.3944
R5332 VDD.n1947 VDD.n1313 19.3944
R5333 VDD.n1947 VDD.n1303 19.3944
R5334 VDD.n1959 VDD.n1303 19.3944
R5335 VDD.n1959 VDD.n1301 19.3944
R5336 VDD.n1963 VDD.n1301 19.3944
R5337 VDD.n1963 VDD.n1291 19.3944
R5338 VDD.n1975 VDD.n1291 19.3944
R5339 VDD.n1975 VDD.n1289 19.3944
R5340 VDD.n1979 VDD.n1289 19.3944
R5341 VDD.n1979 VDD.n1279 19.3944
R5342 VDD.n1991 VDD.n1279 19.3944
R5343 VDD.n1991 VDD.n1277 19.3944
R5344 VDD.n1995 VDD.n1277 19.3944
R5345 VDD.n1995 VDD.n1267 19.3944
R5346 VDD.n2007 VDD.n1267 19.3944
R5347 VDD.n2007 VDD.n1265 19.3944
R5348 VDD.n2011 VDD.n1265 19.3944
R5349 VDD.n2011 VDD.n1256 19.3944
R5350 VDD.n2023 VDD.n1256 19.3944
R5351 VDD.n2023 VDD.n1254 19.3944
R5352 VDD.n2027 VDD.n1254 19.3944
R5353 VDD.n2027 VDD.n1244 19.3944
R5354 VDD.n2039 VDD.n1244 19.3944
R5355 VDD.n2039 VDD.n1242 19.3944
R5356 VDD.n2043 VDD.n1242 19.3944
R5357 VDD.n2043 VDD.n1232 19.3944
R5358 VDD.n2055 VDD.n1232 19.3944
R5359 VDD.n2055 VDD.n1230 19.3944
R5360 VDD.n2059 VDD.n1230 19.3944
R5361 VDD.n2059 VDD.n1220 19.3944
R5362 VDD.n2072 VDD.n1220 19.3944
R5363 VDD.n2072 VDD.n1218 19.3944
R5364 VDD.n2076 VDD.n1218 19.3944
R5365 VDD.n2076 VDD.n1208 19.3944
R5366 VDD.n2090 VDD.n1208 19.3944
R5367 VDD.n2090 VDD.n1206 19.3944
R5368 VDD.n2094 VDD.n1206 19.3944
R5369 VDD.n2094 VDD.n1072 19.3944
R5370 VDD.n2197 VDD.n1072 19.3944
R5371 VDD.n3696 VDD.n289 19.3944
R5372 VDD.n3696 VDD.n279 19.3944
R5373 VDD.n3708 VDD.n279 19.3944
R5374 VDD.n3708 VDD.n277 19.3944
R5375 VDD.n3712 VDD.n277 19.3944
R5376 VDD.n3712 VDD.n267 19.3944
R5377 VDD.n3724 VDD.n267 19.3944
R5378 VDD.n3724 VDD.n265 19.3944
R5379 VDD.n3728 VDD.n265 19.3944
R5380 VDD.n3728 VDD.n255 19.3944
R5381 VDD.n3740 VDD.n255 19.3944
R5382 VDD.n3740 VDD.n253 19.3944
R5383 VDD.n3744 VDD.n253 19.3944
R5384 VDD.n3744 VDD.n243 19.3944
R5385 VDD.n3756 VDD.n243 19.3944
R5386 VDD.n3756 VDD.n241 19.3944
R5387 VDD.n3760 VDD.n241 19.3944
R5388 VDD.n3760 VDD.n231 19.3944
R5389 VDD.n3772 VDD.n231 19.3944
R5390 VDD.n3772 VDD.n229 19.3944
R5391 VDD.n3776 VDD.n229 19.3944
R5392 VDD.n3776 VDD.n219 19.3944
R5393 VDD.n3787 VDD.n219 19.3944
R5394 VDD.n3787 VDD.n217 19.3944
R5395 VDD.n3791 VDD.n217 19.3944
R5396 VDD.n3791 VDD.n207 19.3944
R5397 VDD.n3803 VDD.n207 19.3944
R5398 VDD.n3803 VDD.n205 19.3944
R5399 VDD.n3807 VDD.n205 19.3944
R5400 VDD.n3807 VDD.n195 19.3944
R5401 VDD.n3820 VDD.n195 19.3944
R5402 VDD.n3820 VDD.n193 19.3944
R5403 VDD.n3824 VDD.n193 19.3944
R5404 VDD.n3824 VDD.n184 19.3944
R5405 VDD.n3836 VDD.n184 19.3944
R5406 VDD.n3836 VDD.n182 19.3944
R5407 VDD.n3840 VDD.n182 19.3944
R5408 VDD.n3840 VDD.n172 19.3944
R5409 VDD.n3852 VDD.n172 19.3944
R5410 VDD.n3852 VDD.n170 19.3944
R5411 VDD.n3856 VDD.n170 19.3944
R5412 VDD.n3856 VDD.n160 19.3944
R5413 VDD.n3871 VDD.n160 19.3944
R5414 VDD.n3871 VDD.n158 19.3944
R5415 VDD.n3875 VDD.n158 19.3944
R5416 VDD.n3875 VDD.n149 19.3944
R5417 VDD.n3889 VDD.n149 19.3944
R5418 VDD.n3889 VDD.n147 19.3944
R5419 VDD.n3893 VDD.n147 19.3944
R5420 VDD.n3893 VDD.n35 19.3944
R5421 VDD.n4326 VDD.n35 19.3944
R5422 VDD.n4326 VDD.n4325 19.3944
R5423 VDD.n4325 VDD.n37 19.3944
R5424 VDD.n4319 VDD.n37 19.3944
R5425 VDD.n4319 VDD.n4318 19.3944
R5426 VDD.n4318 VDD.n4317 19.3944
R5427 VDD.n4317 VDD.n49 19.3944
R5428 VDD.n4311 VDD.n49 19.3944
R5429 VDD.n4311 VDD.n4310 19.3944
R5430 VDD.n4310 VDD.n4309 19.3944
R5431 VDD.n4309 VDD.n60 19.3944
R5432 VDD.n4303 VDD.n60 19.3944
R5433 VDD.n4303 VDD.n4302 19.3944
R5434 VDD.n4302 VDD.n4301 19.3944
R5435 VDD.n4301 VDD.n71 19.3944
R5436 VDD.n4295 VDD.n71 19.3944
R5437 VDD.n4295 VDD.n4294 19.3944
R5438 VDD.n4294 VDD.n4293 19.3944
R5439 VDD.n4293 VDD.n82 19.3944
R5440 VDD.n4287 VDD.n82 19.3944
R5441 VDD.n4287 VDD.n4286 19.3944
R5442 VDD.n4286 VDD.n4285 19.3944
R5443 VDD.n4285 VDD.n93 19.3944
R5444 VDD.n4279 VDD.n93 19.3944
R5445 VDD.n4279 VDD.n4278 19.3944
R5446 VDD.n4278 VDD.n4277 19.3944
R5447 VDD.n4277 VDD.n104 19.3944
R5448 VDD.n4271 VDD.n104 19.3944
R5449 VDD.n4271 VDD.n4270 19.3944
R5450 VDD.n4270 VDD.n4269 19.3944
R5451 VDD.n4269 VDD.n115 19.3944
R5452 VDD.n4260 VDD.n115 19.3944
R5453 VDD.n4260 VDD.n4259 19.3944
R5454 VDD.n4259 VDD.n4258 19.3944
R5455 VDD.n4258 VDD.n3954 19.3944
R5456 VDD.n4252 VDD.n3954 19.3944
R5457 VDD.n4252 VDD.n4251 19.3944
R5458 VDD.n4251 VDD.n4250 19.3944
R5459 VDD.n4250 VDD.n3965 19.3944
R5460 VDD.n4244 VDD.n3965 19.3944
R5461 VDD.n4244 VDD.n4243 19.3944
R5462 VDD.n4243 VDD.n4242 19.3944
R5463 VDD.n4242 VDD.n3976 19.3944
R5464 VDD.n4236 VDD.n3976 19.3944
R5465 VDD.n4236 VDD.n4235 19.3944
R5466 VDD.n4235 VDD.n4234 19.3944
R5467 VDD.n4234 VDD.n3986 19.3944
R5468 VDD.n4228 VDD.n3986 19.3944
R5469 VDD.n4228 VDD.n4227 19.3944
R5470 VDD.n4227 VDD.n4226 19.3944
R5471 VDD.n4226 VDD.n3998 19.3944
R5472 VDD.n4157 VDD.n4156 19.3944
R5473 VDD.n4156 VDD.n4153 19.3944
R5474 VDD.n4153 VDD.n4152 19.3944
R5475 VDD.n4152 VDD.n4149 19.3944
R5476 VDD.n4149 VDD.n4148 19.3944
R5477 VDD.n4148 VDD.n4145 19.3944
R5478 VDD.n4145 VDD.n4144 19.3944
R5479 VDD.n4144 VDD.n4141 19.3944
R5480 VDD.n4141 VDD.n4140 19.3944
R5481 VDD.n4140 VDD.n4137 19.3944
R5482 VDD.n4137 VDD.n4136 19.3944
R5483 VDD.n4136 VDD.n4133 19.3944
R5484 VDD.n4133 VDD.n4132 19.3944
R5485 VDD.n4132 VDD.n4129 19.3944
R5486 VDD.n4129 VDD.n4128 19.3944
R5487 VDD.n4188 VDD.n4040 19.3944
R5488 VDD.n4188 VDD.n4185 19.3944
R5489 VDD.n4185 VDD.n4184 19.3944
R5490 VDD.n4184 VDD.n4181 19.3944
R5491 VDD.n4181 VDD.n4180 19.3944
R5492 VDD.n4180 VDD.n4177 19.3944
R5493 VDD.n4177 VDD.n4176 19.3944
R5494 VDD.n4176 VDD.n4173 19.3944
R5495 VDD.n4173 VDD.n4172 19.3944
R5496 VDD.n4172 VDD.n4169 19.3944
R5497 VDD.n4169 VDD.n4168 19.3944
R5498 VDD.n4168 VDD.n4165 19.3944
R5499 VDD.n4165 VDD.n4164 19.3944
R5500 VDD.n4164 VDD.n4161 19.3944
R5501 VDD.n4161 VDD.n4160 19.3944
R5502 VDD.n4220 VDD.n4219 19.3944
R5503 VDD.n4219 VDD.n4029 19.3944
R5504 VDD.n4215 VDD.n4029 19.3944
R5505 VDD.n4215 VDD.n4212 19.3944
R5506 VDD.n4212 VDD.n4209 19.3944
R5507 VDD.n4209 VDD.n4208 19.3944
R5508 VDD.n4208 VDD.n4205 19.3944
R5509 VDD.n4205 VDD.n4204 19.3944
R5510 VDD.n4204 VDD.n4201 19.3944
R5511 VDD.n4201 VDD.n4200 19.3944
R5512 VDD.n4200 VDD.n4197 19.3944
R5513 VDD.n4197 VDD.n4196 19.3944
R5514 VDD.n4196 VDD.n4193 19.3944
R5515 VDD.n3700 VDD.n285 19.3944
R5516 VDD.n3700 VDD.n283 19.3944
R5517 VDD.n3704 VDD.n283 19.3944
R5518 VDD.n3704 VDD.n272 19.3944
R5519 VDD.n3716 VDD.n272 19.3944
R5520 VDD.n3716 VDD.n270 19.3944
R5521 VDD.n3720 VDD.n270 19.3944
R5522 VDD.n3720 VDD.n261 19.3944
R5523 VDD.n3732 VDD.n261 19.3944
R5524 VDD.n3732 VDD.n259 19.3944
R5525 VDD.n3736 VDD.n259 19.3944
R5526 VDD.n3736 VDD.n249 19.3944
R5527 VDD.n3748 VDD.n249 19.3944
R5528 VDD.n3748 VDD.n247 19.3944
R5529 VDD.n3752 VDD.n247 19.3944
R5530 VDD.n3752 VDD.n237 19.3944
R5531 VDD.n3764 VDD.n237 19.3944
R5532 VDD.n3764 VDD.n235 19.3944
R5533 VDD.n3768 VDD.n235 19.3944
R5534 VDD.n3768 VDD.n225 19.3944
R5535 VDD.n3779 VDD.n225 19.3944
R5536 VDD.n3779 VDD.n223 19.3944
R5537 VDD.n3783 VDD.n223 19.3944
R5538 VDD.n3783 VDD.n213 19.3944
R5539 VDD.n3795 VDD.n213 19.3944
R5540 VDD.n3795 VDD.n211 19.3944
R5541 VDD.n3799 VDD.n211 19.3944
R5542 VDD.n3799 VDD.n201 19.3944
R5543 VDD.n3811 VDD.n201 19.3944
R5544 VDD.n3811 VDD.n199 19.3944
R5545 VDD.n3815 VDD.n199 19.3944
R5546 VDD.n3815 VDD.n190 19.3944
R5547 VDD.n3828 VDD.n190 19.3944
R5548 VDD.n3828 VDD.n188 19.3944
R5549 VDD.n3832 VDD.n188 19.3944
R5550 VDD.n3832 VDD.n178 19.3944
R5551 VDD.n3844 VDD.n178 19.3944
R5552 VDD.n3844 VDD.n176 19.3944
R5553 VDD.n3848 VDD.n176 19.3944
R5554 VDD.n3848 VDD.n166 19.3944
R5555 VDD.n3860 VDD.n166 19.3944
R5556 VDD.n3860 VDD.n164 19.3944
R5557 VDD.n3866 VDD.n164 19.3944
R5558 VDD.n3866 VDD.n3865 19.3944
R5559 VDD.n3865 VDD.n155 19.3944
R5560 VDD.n3880 VDD.n155 19.3944
R5561 VDD.n3880 VDD.n153 19.3944
R5562 VDD.n3884 VDD.n153 19.3944
R5563 VDD.n3884 VDD.n142 19.3944
R5564 VDD.n3898 VDD.n142 19.3944
R5565 VDD.n3898 VDD.n140 19.3944
R5566 VDD.n3902 VDD.n140 19.3944
R5567 VDD.n3903 VDD.n3902 19.3944
R5568 VDD.n3904 VDD.n3903 19.3944
R5569 VDD.n3904 VDD.n138 19.3944
R5570 VDD.n3908 VDD.n138 19.3944
R5571 VDD.n3909 VDD.n3908 19.3944
R5572 VDD.n3910 VDD.n3909 19.3944
R5573 VDD.n3910 VDD.n135 19.3944
R5574 VDD.n3914 VDD.n135 19.3944
R5575 VDD.n3915 VDD.n3914 19.3944
R5576 VDD.n3916 VDD.n3915 19.3944
R5577 VDD.n3916 VDD.n132 19.3944
R5578 VDD.n3920 VDD.n132 19.3944
R5579 VDD.n3921 VDD.n3920 19.3944
R5580 VDD.n3922 VDD.n3921 19.3944
R5581 VDD.n3922 VDD.n129 19.3944
R5582 VDD.n3926 VDD.n129 19.3944
R5583 VDD.n3927 VDD.n3926 19.3944
R5584 VDD.n3928 VDD.n3927 19.3944
R5585 VDD.n3928 VDD.n126 19.3944
R5586 VDD.n3932 VDD.n126 19.3944
R5587 VDD.n3933 VDD.n3932 19.3944
R5588 VDD.n3934 VDD.n3933 19.3944
R5589 VDD.n3934 VDD.n123 19.3944
R5590 VDD.n3938 VDD.n123 19.3944
R5591 VDD.n3939 VDD.n3938 19.3944
R5592 VDD.n3940 VDD.n3939 19.3944
R5593 VDD.n3940 VDD.n120 19.3944
R5594 VDD.n4266 VDD.n120 19.3944
R5595 VDD.n4266 VDD.n4265 19.3944
R5596 VDD.n4265 VDD.n4264 19.3944
R5597 VDD.n4264 VDD.n3946 19.3944
R5598 VDD.n4092 VDD.n3946 19.3944
R5599 VDD.n4093 VDD.n4092 19.3944
R5600 VDD.n4093 VDD.n4089 19.3944
R5601 VDD.n4098 VDD.n4089 19.3944
R5602 VDD.n4099 VDD.n4098 19.3944
R5603 VDD.n4100 VDD.n4099 19.3944
R5604 VDD.n4100 VDD.n4087 19.3944
R5605 VDD.n4105 VDD.n4087 19.3944
R5606 VDD.n4106 VDD.n4105 19.3944
R5607 VDD.n4107 VDD.n4106 19.3944
R5608 VDD.n4107 VDD.n4085 19.3944
R5609 VDD.n4112 VDD.n4085 19.3944
R5610 VDD.n4113 VDD.n4112 19.3944
R5611 VDD.n4114 VDD.n4113 19.3944
R5612 VDD.n4114 VDD.n4083 19.3944
R5613 VDD.n4119 VDD.n4083 19.3944
R5614 VDD.n4120 VDD.n4119 19.3944
R5615 VDD.n4121 VDD.n4120 19.3944
R5616 VDD.n3684 VDD.n3683 19.3944
R5617 VDD.n3691 VDD.n294 19.3944
R5618 VDD.n3691 VDD.n295 19.3944
R5619 VDD.n3572 VDD.n295 19.3944
R5620 VDD.n3572 VDD.n3569 19.3944
R5621 VDD.n3576 VDD.n3569 19.3944
R5622 VDD.n3579 VDD.n3576 19.3944
R5623 VDD.n3582 VDD.n3579 19.3944
R5624 VDD.n3582 VDD.n3567 19.3944
R5625 VDD.n3586 VDD.n3567 19.3944
R5626 VDD.n3589 VDD.n3586 19.3944
R5627 VDD.n3598 VDD.n3565 19.3944
R5628 VDD.n3601 VDD.n3598 19.3944
R5629 VDD.n3604 VDD.n3601 19.3944
R5630 VDD.n3604 VDD.n3563 19.3944
R5631 VDD.n3608 VDD.n3563 19.3944
R5632 VDD.n3611 VDD.n3608 19.3944
R5633 VDD.n3614 VDD.n3611 19.3944
R5634 VDD.n3614 VDD.n3561 19.3944
R5635 VDD.n3618 VDD.n3561 19.3944
R5636 VDD.n3621 VDD.n3618 19.3944
R5637 VDD.n3624 VDD.n3621 19.3944
R5638 VDD.n3624 VDD.n3559 19.3944
R5639 VDD.n3628 VDD.n3559 19.3944
R5640 VDD.n3631 VDD.n3628 19.3944
R5641 VDD.n3637 VDD.n3631 19.3944
R5642 VDD.n3641 VDD.n3557 19.3944
R5643 VDD.n3644 VDD.n3641 19.3944
R5644 VDD.n3647 VDD.n3644 19.3944
R5645 VDD.n3647 VDD.n3555 19.3944
R5646 VDD.n3651 VDD.n3555 19.3944
R5647 VDD.n3654 VDD.n3651 19.3944
R5648 VDD.n3657 VDD.n3654 19.3944
R5649 VDD.n3657 VDD.n3553 19.3944
R5650 VDD.n3661 VDD.n3553 19.3944
R5651 VDD.n3664 VDD.n3661 19.3944
R5652 VDD.n3667 VDD.n3664 19.3944
R5653 VDD.n3667 VDD.n3551 19.3944
R5654 VDD.n3671 VDD.n3551 19.3944
R5655 VDD.n3674 VDD.n3671 19.3944
R5656 VDD.n1600 VDD.n1502 16.8732
R5657 VDD.n1199 VDD.n1146 16.8732
R5658 VDD.n4128 VDD.n4125 16.8732
R5659 VDD.n3678 VDD.n3677 16.8732
R5660 VDD.n2784 VDD.n628 15.8624
R5661 VDD.n3174 VDD.n622 15.8624
R5662 VDD.n1682 VDD.n1496 14.2905
R5663 VDD.n1682 VDD.n1490 14.2905
R5664 VDD.n1690 VDD.n1490 14.2905
R5665 VDD.n1690 VDD.n1484 14.2905
R5666 VDD.n1699 VDD.n1484 14.2905
R5667 VDD.n1699 VDD.n1698 14.2905
R5668 VDD.n1707 VDD.n1473 14.2905
R5669 VDD.n1715 VDD.n1473 14.2905
R5670 VDD.n1715 VDD.n1467 14.2905
R5671 VDD.n1723 VDD.n1467 14.2905
R5672 VDD.n1723 VDD.n1461 14.2905
R5673 VDD.n1731 VDD.n1461 14.2905
R5674 VDD.n1731 VDD.n1455 14.2905
R5675 VDD.n1739 VDD.n1455 14.2905
R5676 VDD.n1739 VDD.n1449 14.2905
R5677 VDD.n1747 VDD.n1449 14.2905
R5678 VDD.n1747 VDD.n1443 14.2905
R5679 VDD.n1755 VDD.n1443 14.2905
R5680 VDD.n1755 VDD.n1437 14.2905
R5681 VDD.t91 VDD.n1437 14.2905
R5682 VDD.t91 VDD.n1431 14.2905
R5683 VDD.n1770 VDD.n1431 14.2905
R5684 VDD.n1770 VDD.n1425 14.2905
R5685 VDD.n1778 VDD.n1425 14.2905
R5686 VDD.n1778 VDD.n1419 14.2905
R5687 VDD.n1786 VDD.n1419 14.2905
R5688 VDD.n1786 VDD.n1413 14.2905
R5689 VDD.n1794 VDD.n1413 14.2905
R5690 VDD.n1794 VDD.n1406 14.2905
R5691 VDD.n1802 VDD.n1406 14.2905
R5692 VDD.n1802 VDD.n1407 14.2905
R5693 VDD.n1810 VDD.n1395 14.2905
R5694 VDD.n1818 VDD.n1395 14.2905
R5695 VDD.n1818 VDD.n1389 14.2905
R5696 VDD.n1826 VDD.n1389 14.2905
R5697 VDD.n1826 VDD.n1383 14.2905
R5698 VDD.n1834 VDD.n1383 14.2905
R5699 VDD.n1834 VDD.n1377 14.2905
R5700 VDD.n1842 VDD.n1377 14.2905
R5701 VDD.n1842 VDD.n1370 14.2905
R5702 VDD.n1850 VDD.n1370 14.2905
R5703 VDD.n1850 VDD.n1371 14.2905
R5704 VDD.n1858 VDD.n1359 14.2905
R5705 VDD.n1866 VDD.n1359 14.2905
R5706 VDD.n1866 VDD.n1353 14.2905
R5707 VDD.n1874 VDD.n1353 14.2905
R5708 VDD.n1874 VDD.n1347 14.2905
R5709 VDD.n1901 VDD.n1347 14.2905
R5710 VDD.n1901 VDD.n1341 14.2905
R5711 VDD.n1909 VDD.n1341 14.2905
R5712 VDD.n1909 VDD.n1334 14.2905
R5713 VDD.n1917 VDD.n1334 14.2905
R5714 VDD.n1917 VDD.n1335 14.2905
R5715 VDD.n1925 VDD.n1323 14.2905
R5716 VDD.n1933 VDD.n1323 14.2905
R5717 VDD.n1933 VDD.n1317 14.2905
R5718 VDD.n1941 VDD.n1317 14.2905
R5719 VDD.n1941 VDD.n1311 14.2905
R5720 VDD.n1949 VDD.n1311 14.2905
R5721 VDD.n1949 VDD.n1305 14.2905
R5722 VDD.n1957 VDD.n1305 14.2905
R5723 VDD.n1957 VDD.n1298 14.2905
R5724 VDD.n1965 VDD.n1298 14.2905
R5725 VDD.n1965 VDD.n1299 14.2905
R5726 VDD.n1973 VDD.n1287 14.2905
R5727 VDD.n1981 VDD.n1287 14.2905
R5728 VDD.n1981 VDD.n1281 14.2905
R5729 VDD.n1989 VDD.n1281 14.2905
R5730 VDD.n1989 VDD.n1275 14.2905
R5731 VDD.n1997 VDD.n1275 14.2905
R5732 VDD.n1997 VDD.n1269 14.2905
R5733 VDD.n2005 VDD.n1269 14.2905
R5734 VDD.n2005 VDD.n1263 14.2905
R5735 VDD.n2013 VDD.n1263 14.2905
R5736 VDD.n2013 VDD.t77 14.2905
R5737 VDD.n2021 VDD.t77 14.2905
R5738 VDD.n2021 VDD.n1252 14.2905
R5739 VDD.n2029 VDD.n1252 14.2905
R5740 VDD.n2029 VDD.n1246 14.2905
R5741 VDD.n2037 VDD.n1246 14.2905
R5742 VDD.n2037 VDD.n1240 14.2905
R5743 VDD.n2045 VDD.n1240 14.2905
R5744 VDD.n2045 VDD.n1234 14.2905
R5745 VDD.n2053 VDD.n1234 14.2905
R5746 VDD.n2053 VDD.n1228 14.2905
R5747 VDD.n2061 VDD.n1228 14.2905
R5748 VDD.n2061 VDD.n1222 14.2905
R5749 VDD.n2070 VDD.n1222 14.2905
R5750 VDD.n2070 VDD.n2069 14.2905
R5751 VDD.n2078 VDD.n1210 14.2905
R5752 VDD.n2088 VDD.n1210 14.2905
R5753 VDD.n2088 VDD.n1204 14.2905
R5754 VDD.n2096 VDD.n1204 14.2905
R5755 VDD.n2096 VDD.n1075 14.2905
R5756 VDD.n2195 VDD.n1075 14.2905
R5757 VDD.n3698 VDD.n287 14.2905
R5758 VDD.n3698 VDD.n281 14.2905
R5759 VDD.n3706 VDD.n281 14.2905
R5760 VDD.n3706 VDD.n274 14.2905
R5761 VDD.n3714 VDD.n274 14.2905
R5762 VDD.n3714 VDD.n275 14.2905
R5763 VDD.n3722 VDD.n263 14.2905
R5764 VDD.n3730 VDD.n263 14.2905
R5765 VDD.n3730 VDD.n257 14.2905
R5766 VDD.n3738 VDD.n257 14.2905
R5767 VDD.n3738 VDD.n251 14.2905
R5768 VDD.n3746 VDD.n251 14.2905
R5769 VDD.n3746 VDD.n245 14.2905
R5770 VDD.n3754 VDD.n245 14.2905
R5771 VDD.n3754 VDD.n239 14.2905
R5772 VDD.n3762 VDD.n239 14.2905
R5773 VDD.n3762 VDD.n233 14.2905
R5774 VDD.n3770 VDD.n233 14.2905
R5775 VDD.n3770 VDD.n227 14.2905
R5776 VDD.t81 VDD.n227 14.2905
R5777 VDD.t81 VDD.n221 14.2905
R5778 VDD.n3785 VDD.n221 14.2905
R5779 VDD.n3785 VDD.n215 14.2905
R5780 VDD.n3793 VDD.n215 14.2905
R5781 VDD.n3793 VDD.n209 14.2905
R5782 VDD.n3801 VDD.n209 14.2905
R5783 VDD.n3801 VDD.n203 14.2905
R5784 VDD.n3809 VDD.n203 14.2905
R5785 VDD.n3809 VDD.n197 14.2905
R5786 VDD.n3818 VDD.n197 14.2905
R5787 VDD.n3818 VDD.n3817 14.2905
R5788 VDD.n3826 VDD.n186 14.2905
R5789 VDD.n3834 VDD.n186 14.2905
R5790 VDD.n3834 VDD.n180 14.2905
R5791 VDD.n3842 VDD.n180 14.2905
R5792 VDD.n3842 VDD.n174 14.2905
R5793 VDD.n3850 VDD.n174 14.2905
R5794 VDD.n3850 VDD.n168 14.2905
R5795 VDD.n3858 VDD.n168 14.2905
R5796 VDD.n3858 VDD.n162 14.2905
R5797 VDD.n3869 VDD.n162 14.2905
R5798 VDD.n3869 VDD.n3868 14.2905
R5799 VDD.n3877 VDD.n151 14.2905
R5800 VDD.n3887 VDD.n151 14.2905
R5801 VDD.n3887 VDD.n3886 14.2905
R5802 VDD.n3886 VDD.n145 14.2905
R5803 VDD.n3896 VDD.n145 14.2905
R5804 VDD.n3896 VDD.n39 14.2905
R5805 VDD.n4323 VDD.n39 14.2905
R5806 VDD.n4323 VDD.n4322 14.2905
R5807 VDD.n4322 VDD.n4321 14.2905
R5808 VDD.n4321 VDD.n43 14.2905
R5809 VDD.n4315 VDD.n43 14.2905
R5810 VDD.n4314 VDD.n4313 14.2905
R5811 VDD.n4313 VDD.n54 14.2905
R5812 VDD.n4307 VDD.n54 14.2905
R5813 VDD.n4307 VDD.n4306 14.2905
R5814 VDD.n4306 VDD.n4305 14.2905
R5815 VDD.n4305 VDD.n65 14.2905
R5816 VDD.n4299 VDD.n65 14.2905
R5817 VDD.n4299 VDD.n4298 14.2905
R5818 VDD.n4298 VDD.n4297 14.2905
R5819 VDD.n4297 VDD.n76 14.2905
R5820 VDD.n4291 VDD.n76 14.2905
R5821 VDD.n4290 VDD.n4289 14.2905
R5822 VDD.n4289 VDD.n87 14.2905
R5823 VDD.n4283 VDD.n87 14.2905
R5824 VDD.n4283 VDD.n4282 14.2905
R5825 VDD.n4282 VDD.n4281 14.2905
R5826 VDD.n4281 VDD.n98 14.2905
R5827 VDD.n4275 VDD.n98 14.2905
R5828 VDD.n4275 VDD.n4274 14.2905
R5829 VDD.n4274 VDD.n4273 14.2905
R5830 VDD.n4273 VDD.n109 14.2905
R5831 VDD.t99 VDD.n109 14.2905
R5832 VDD.t99 VDD.n117 14.2905
R5833 VDD.n4262 VDD.n117 14.2905
R5834 VDD.n4262 VDD.n3948 14.2905
R5835 VDD.n4256 VDD.n3948 14.2905
R5836 VDD.n4256 VDD.n4255 14.2905
R5837 VDD.n4255 VDD.n4254 14.2905
R5838 VDD.n4254 VDD.n3959 14.2905
R5839 VDD.n4248 VDD.n3959 14.2905
R5840 VDD.n4248 VDD.n4247 14.2905
R5841 VDD.n4247 VDD.n4246 14.2905
R5842 VDD.n4246 VDD.n3970 14.2905
R5843 VDD.n4240 VDD.n3970 14.2905
R5844 VDD.n4240 VDD.n4239 14.2905
R5845 VDD.n4239 VDD.n4238 14.2905
R5846 VDD.n4232 VDD.n3988 14.2905
R5847 VDD.n4232 VDD.n4231 14.2905
R5848 VDD.n4231 VDD.n4230 14.2905
R5849 VDD.n4230 VDD.n3992 14.2905
R5850 VDD.n4224 VDD.n3992 14.2905
R5851 VDD.n4224 VDD.n4223 14.2905
R5852 VDD.n1651 VDD.n1548 14.1581
R5853 VDD.n2168 VDD.n2167 14.1581
R5854 VDD.n4193 VDD.n4192 14.1581
R5855 VDD.n3594 VDD.n3589 14.1581
R5856 VDD.n29 VDD.t87 13.377
R5857 VDD.n29 VDD.t72 13.377
R5858 VDD.n27 VDD.t95 13.377
R5859 VDD.n27 VDD.t105 13.377
R5860 VDD.n23 VDD.t84 13.377
R5861 VDD.n23 VDD.t71 13.377
R5862 VDD.n21 VDD.t96 13.377
R5863 VDD.n21 VDD.t108 13.377
R5864 VDD.n18 VDD.t102 13.377
R5865 VDD.n18 VDD.t101 13.377
R5866 VDD.n16 VDD.t80 13.377
R5867 VDD.n16 VDD.t104 13.377
R5868 VDD.n1890 VDD.t116 13.377
R5869 VDD.n1890 VDD.t76 13.377
R5870 VDD.n1892 VDD.t86 13.377
R5871 VDD.n1892 VDD.t98 13.377
R5872 VDD.n1884 VDD.t117 13.377
R5873 VDD.n1884 VDD.t75 13.377
R5874 VDD.n1886 VDD.t88 13.377
R5875 VDD.n1886 VDD.t106 13.377
R5876 VDD.n1879 VDD.t111 13.377
R5877 VDD.n1879 VDD.t74 13.377
R5878 VDD.n1881 VDD.t109 13.377
R5879 VDD.n1881 VDD.t107 13.377
R5880 VDD.n7 VDD.t131 12.6238
R5881 VDD.n7 VDD.t145 12.6238
R5882 VDD.n8 VDD.t119 12.6238
R5883 VDD.n8 VDD.t149 12.6238
R5884 VDD.n10 VDD.t151 12.6238
R5885 VDD.n10 VDD.t122 12.6238
R5886 VDD.n12 VDD.t135 12.6238
R5887 VDD.n12 VDD.t126 12.6238
R5888 VDD.n5 VDD.t133 12.6238
R5889 VDD.n5 VDD.t153 12.6238
R5890 VDD.n3 VDD.t147 12.6238
R5891 VDD.n3 VDD.t157 12.6238
R5892 VDD.n1 VDD.t155 12.6238
R5893 VDD.n1 VDD.t138 12.6238
R5894 VDD.n0 VDD.t129 12.6238
R5895 VDD.n0 VDD.t141 12.6238
R5896 VDD.n1647 VDD.n1548 11.8308
R5897 VDD.n2167 VDD.n1110 11.8308
R5898 VDD.n4192 VDD.n4040 11.8308
R5899 VDD.n3594 VDD.n3565 11.8308
R5900 VDD.n1407 VDD.t85 11.4325
R5901 VDD.n1973 VDD.t73 11.4325
R5902 VDD.n3817 VDD.t79 11.4325
R5903 VDD.t70 VDD.n4290 11.4325
R5904 VDD.n2404 VDD.n923 10.6151
R5905 VDD.n2414 VDD.n923 10.6151
R5906 VDD.n2415 VDD.n2414 10.6151
R5907 VDD.n2416 VDD.n2415 10.6151
R5908 VDD.n2416 VDD.n911 10.6151
R5909 VDD.n2426 VDD.n911 10.6151
R5910 VDD.n2427 VDD.n2426 10.6151
R5911 VDD.n2428 VDD.n2427 10.6151
R5912 VDD.n2428 VDD.n898 10.6151
R5913 VDD.n2438 VDD.n898 10.6151
R5914 VDD.n2439 VDD.n2438 10.6151
R5915 VDD.n2440 VDD.n2439 10.6151
R5916 VDD.n2440 VDD.n887 10.6151
R5917 VDD.n2450 VDD.n887 10.6151
R5918 VDD.n2451 VDD.n2450 10.6151
R5919 VDD.n2452 VDD.n2451 10.6151
R5920 VDD.n2452 VDD.n875 10.6151
R5921 VDD.n2462 VDD.n875 10.6151
R5922 VDD.n2463 VDD.n2462 10.6151
R5923 VDD.n2464 VDD.n2463 10.6151
R5924 VDD.n2464 VDD.n863 10.6151
R5925 VDD.n2474 VDD.n863 10.6151
R5926 VDD.n2475 VDD.n2474 10.6151
R5927 VDD.n2476 VDD.n2475 10.6151
R5928 VDD.n2476 VDD.n852 10.6151
R5929 VDD.n2486 VDD.n852 10.6151
R5930 VDD.n2487 VDD.n2486 10.6151
R5931 VDD.n2488 VDD.n2487 10.6151
R5932 VDD.n2488 VDD.n840 10.6151
R5933 VDD.n2498 VDD.n840 10.6151
R5934 VDD.n2499 VDD.n2498 10.6151
R5935 VDD.n2500 VDD.n2499 10.6151
R5936 VDD.n2500 VDD.n828 10.6151
R5937 VDD.n2510 VDD.n828 10.6151
R5938 VDD.n2511 VDD.n2510 10.6151
R5939 VDD.n2512 VDD.n2511 10.6151
R5940 VDD.n2512 VDD.n816 10.6151
R5941 VDD.n2522 VDD.n816 10.6151
R5942 VDD.n2523 VDD.n2522 10.6151
R5943 VDD.n2524 VDD.n2523 10.6151
R5944 VDD.n2524 VDD.n803 10.6151
R5945 VDD.n2534 VDD.n803 10.6151
R5946 VDD.n2535 VDD.n2534 10.6151
R5947 VDD.n2536 VDD.n2535 10.6151
R5948 VDD.n2536 VDD.n792 10.6151
R5949 VDD.n2546 VDD.n792 10.6151
R5950 VDD.n2547 VDD.n2546 10.6151
R5951 VDD.n2548 VDD.n2547 10.6151
R5952 VDD.n2548 VDD.n780 10.6151
R5953 VDD.n2558 VDD.n780 10.6151
R5954 VDD.n2559 VDD.n2558 10.6151
R5955 VDD.n2560 VDD.n2559 10.6151
R5956 VDD.n2560 VDD.n768 10.6151
R5957 VDD.n2570 VDD.n768 10.6151
R5958 VDD.n2571 VDD.n2570 10.6151
R5959 VDD.n2572 VDD.n2571 10.6151
R5960 VDD.n2572 VDD.n756 10.6151
R5961 VDD.n2582 VDD.n756 10.6151
R5962 VDD.n2583 VDD.n2582 10.6151
R5963 VDD.n2584 VDD.n2583 10.6151
R5964 VDD.n2584 VDD.n743 10.6151
R5965 VDD.n2594 VDD.n743 10.6151
R5966 VDD.n2595 VDD.n2594 10.6151
R5967 VDD.n2596 VDD.n2595 10.6151
R5968 VDD.n2596 VDD.n732 10.6151
R5969 VDD.n2606 VDD.n732 10.6151
R5970 VDD.n2607 VDD.n2606 10.6151
R5971 VDD.n2608 VDD.n2607 10.6151
R5972 VDD.n2608 VDD.n720 10.6151
R5973 VDD.n2618 VDD.n720 10.6151
R5974 VDD.n2619 VDD.n2618 10.6151
R5975 VDD.n2620 VDD.n2619 10.6151
R5976 VDD.n2620 VDD.n708 10.6151
R5977 VDD.n2630 VDD.n708 10.6151
R5978 VDD.n2631 VDD.n2630 10.6151
R5979 VDD.n2632 VDD.n2631 10.6151
R5980 VDD.n2632 VDD.n696 10.6151
R5981 VDD.n2642 VDD.n696 10.6151
R5982 VDD.n2643 VDD.n2642 10.6151
R5983 VDD.n2644 VDD.n2643 10.6151
R5984 VDD.n2644 VDD.n683 10.6151
R5985 VDD.n2656 VDD.n683 10.6151
R5986 VDD.n2657 VDD.n2656 10.6151
R5987 VDD.n2658 VDD.n2657 10.6151
R5988 VDD.n2658 VDD.n667 10.6151
R5989 VDD.n2728 VDD.n667 10.6151
R5990 VDD.n2729 VDD.n2728 10.6151
R5991 VDD.n2730 VDD.n2729 10.6151
R5992 VDD.n2730 VDD.n656 10.6151
R5993 VDD.n2782 VDD.n2781 10.6151
R5994 VDD.n2781 VDD.n2780 10.6151
R5995 VDD.n2780 VDD.n2777 10.6151
R5996 VDD.n2777 VDD.n2776 10.6151
R5997 VDD.n2776 VDD.n2773 10.6151
R5998 VDD.n2773 VDD.n2772 10.6151
R5999 VDD.n2772 VDD.n2769 10.6151
R6000 VDD.n2769 VDD.n2768 10.6151
R6001 VDD.n2768 VDD.n2765 10.6151
R6002 VDD.n2765 VDD.n2764 10.6151
R6003 VDD.n2764 VDD.n2761 10.6151
R6004 VDD.n2761 VDD.n2760 10.6151
R6005 VDD.n2760 VDD.n2757 10.6151
R6006 VDD.n2757 VDD.n2756 10.6151
R6007 VDD.n2756 VDD.n2753 10.6151
R6008 VDD.n2753 VDD.n2752 10.6151
R6009 VDD.n2752 VDD.n2749 10.6151
R6010 VDD.n2749 VDD.n2748 10.6151
R6011 VDD.n2748 VDD.n2745 10.6151
R6012 VDD.n2745 VDD.n2744 10.6151
R6013 VDD.n2741 VDD.n2740 10.6151
R6014 VDD.n2740 VDD.n2737 10.6151
R6015 VDD.n2737 VDD.n2736 10.6151
R6016 VDD.n2228 VDD.n2226 10.6151
R6017 VDD.n2229 VDD.n2228 10.6151
R6018 VDD.n2231 VDD.n2229 10.6151
R6019 VDD.n2232 VDD.n2231 10.6151
R6020 VDD.n2234 VDD.n2232 10.6151
R6021 VDD.n2235 VDD.n2234 10.6151
R6022 VDD.n2237 VDD.n2235 10.6151
R6023 VDD.n2238 VDD.n2237 10.6151
R6024 VDD.n2240 VDD.n2238 10.6151
R6025 VDD.n2241 VDD.n2240 10.6151
R6026 VDD.n2243 VDD.n2241 10.6151
R6027 VDD.n2244 VDD.n2243 10.6151
R6028 VDD.n2246 VDD.n2244 10.6151
R6029 VDD.n2247 VDD.n2246 10.6151
R6030 VDD.n2249 VDD.n2247 10.6151
R6031 VDD.n2250 VDD.n2249 10.6151
R6032 VDD.n2252 VDD.n2250 10.6151
R6033 VDD.n2253 VDD.n2252 10.6151
R6034 VDD.n2255 VDD.n2253 10.6151
R6035 VDD.n2256 VDD.n2255 10.6151
R6036 VDD.n2258 VDD.n2256 10.6151
R6037 VDD.n2259 VDD.n2258 10.6151
R6038 VDD.n2261 VDD.n2259 10.6151
R6039 VDD.n2262 VDD.n2261 10.6151
R6040 VDD.n2355 VDD.n2262 10.6151
R6041 VDD.n2355 VDD.n2354 10.6151
R6042 VDD.n2354 VDD.n2353 10.6151
R6043 VDD.n2353 VDD.n2351 10.6151
R6044 VDD.n2351 VDD.n2350 10.6151
R6045 VDD.n2350 VDD.n2348 10.6151
R6046 VDD.n2348 VDD.n2347 10.6151
R6047 VDD.n2347 VDD.n2345 10.6151
R6048 VDD.n2345 VDD.n2344 10.6151
R6049 VDD.n2344 VDD.n2342 10.6151
R6050 VDD.n2342 VDD.n2341 10.6151
R6051 VDD.n2341 VDD.n2339 10.6151
R6052 VDD.n2339 VDD.n2338 10.6151
R6053 VDD.n2338 VDD.n2336 10.6151
R6054 VDD.n2336 VDD.n2335 10.6151
R6055 VDD.n2335 VDD.n2333 10.6151
R6056 VDD.n2333 VDD.n2332 10.6151
R6057 VDD.n2332 VDD.n2330 10.6151
R6058 VDD.n2330 VDD.n2329 10.6151
R6059 VDD.n2329 VDD.n2327 10.6151
R6060 VDD.n2327 VDD.n2326 10.6151
R6061 VDD.n2326 VDD.n2324 10.6151
R6062 VDD.n2324 VDD.n2323 10.6151
R6063 VDD.n2323 VDD.n2321 10.6151
R6064 VDD.n2321 VDD.n2320 10.6151
R6065 VDD.n2320 VDD.n2318 10.6151
R6066 VDD.n2318 VDD.n2317 10.6151
R6067 VDD.n2317 VDD.n2315 10.6151
R6068 VDD.n2315 VDD.n2314 10.6151
R6069 VDD.n2314 VDD.n2312 10.6151
R6070 VDD.n2312 VDD.n2311 10.6151
R6071 VDD.n2311 VDD.n2309 10.6151
R6072 VDD.n2309 VDD.n2308 10.6151
R6073 VDD.n2308 VDD.n2306 10.6151
R6074 VDD.n2306 VDD.n2305 10.6151
R6075 VDD.n2305 VDD.n2303 10.6151
R6076 VDD.n2303 VDD.n2302 10.6151
R6077 VDD.n2302 VDD.n2300 10.6151
R6078 VDD.n2300 VDD.n2299 10.6151
R6079 VDD.n2299 VDD.n2297 10.6151
R6080 VDD.n2297 VDD.n2296 10.6151
R6081 VDD.n2296 VDD.n2294 10.6151
R6082 VDD.n2294 VDD.n2293 10.6151
R6083 VDD.n2293 VDD.n2291 10.6151
R6084 VDD.n2291 VDD.n2290 10.6151
R6085 VDD.n2290 VDD.n2288 10.6151
R6086 VDD.n2288 VDD.n2287 10.6151
R6087 VDD.n2287 VDD.n2285 10.6151
R6088 VDD.n2285 VDD.n2284 10.6151
R6089 VDD.n2284 VDD.n2282 10.6151
R6090 VDD.n2282 VDD.n2281 10.6151
R6091 VDD.n2281 VDD.n2279 10.6151
R6092 VDD.n2279 VDD.n2278 10.6151
R6093 VDD.n2278 VDD.n2276 10.6151
R6094 VDD.n2276 VDD.n2275 10.6151
R6095 VDD.n2275 VDD.n2273 10.6151
R6096 VDD.n2273 VDD.n2272 10.6151
R6097 VDD.n2272 VDD.n2270 10.6151
R6098 VDD.n2270 VDD.n2269 10.6151
R6099 VDD.n2269 VDD.n2267 10.6151
R6100 VDD.n2267 VDD.n2266 10.6151
R6101 VDD.n2266 VDD.n2264 10.6151
R6102 VDD.n2264 VDD.n2263 10.6151
R6103 VDD.n2263 VDD.n662 10.6151
R6104 VDD.n662 VDD.n660 10.6151
R6105 VDD.n2403 VDD.n2402 10.6151
R6106 VDD.n2402 VDD.n934 10.6151
R6107 VDD.n1051 VDD.n934 10.6151
R6108 VDD.n1052 VDD.n1051 10.6151
R6109 VDD.n1055 VDD.n1052 10.6151
R6110 VDD.n1056 VDD.n1055 10.6151
R6111 VDD.n1059 VDD.n1056 10.6151
R6112 VDD.n1060 VDD.n1059 10.6151
R6113 VDD.n1063 VDD.n1060 10.6151
R6114 VDD.n1064 VDD.n1063 10.6151
R6115 VDD.n1067 VDD.n1064 10.6151
R6116 VDD.n2200 VDD.n1067 10.6151
R6117 VDD.n2203 VDD.n2200 10.6151
R6118 VDD.n2204 VDD.n2203 10.6151
R6119 VDD.n2207 VDD.n2204 10.6151
R6120 VDD.n2208 VDD.n2207 10.6151
R6121 VDD.n2211 VDD.n2208 10.6151
R6122 VDD.n2212 VDD.n2211 10.6151
R6123 VDD.n2215 VDD.n2212 10.6151
R6124 VDD.n2216 VDD.n2215 10.6151
R6125 VDD.n2220 VDD.n2219 10.6151
R6126 VDD.n2223 VDD.n2220 10.6151
R6127 VDD.n2225 VDD.n2223 10.6151
R6128 VDD.n3123 VDD.n3122 10.6151
R6129 VDD.n3122 VDD.n3121 10.6151
R6130 VDD.n3121 VDD.n3119 10.6151
R6131 VDD.n3119 VDD.n3118 10.6151
R6132 VDD.n3118 VDD.n3116 10.6151
R6133 VDD.n3116 VDD.n3115 10.6151
R6134 VDD.n3115 VDD.n3113 10.6151
R6135 VDD.n3113 VDD.n3112 10.6151
R6136 VDD.n3112 VDD.n3110 10.6151
R6137 VDD.n3110 VDD.n3109 10.6151
R6138 VDD.n3109 VDD.n3107 10.6151
R6139 VDD.n3107 VDD.n3106 10.6151
R6140 VDD.n3106 VDD.n3104 10.6151
R6141 VDD.n3104 VDD.n3103 10.6151
R6142 VDD.n3103 VDD.n3101 10.6151
R6143 VDD.n3101 VDD.n3100 10.6151
R6144 VDD.n3100 VDD.n3098 10.6151
R6145 VDD.n3098 VDD.n3097 10.6151
R6146 VDD.n3097 VDD.n3095 10.6151
R6147 VDD.n3095 VDD.n3094 10.6151
R6148 VDD.n3094 VDD.n3092 10.6151
R6149 VDD.n3092 VDD.n3091 10.6151
R6150 VDD.n3091 VDD.n3089 10.6151
R6151 VDD.n3089 VDD.n3088 10.6151
R6152 VDD.n3088 VDD.n3086 10.6151
R6153 VDD.n3086 VDD.n3085 10.6151
R6154 VDD.n3085 VDD.n3083 10.6151
R6155 VDD.n3083 VDD.n3082 10.6151
R6156 VDD.n3082 VDD.n3080 10.6151
R6157 VDD.n3080 VDD.n3079 10.6151
R6158 VDD.n3079 VDD.n3077 10.6151
R6159 VDD.n3077 VDD.n3076 10.6151
R6160 VDD.n3076 VDD.n3074 10.6151
R6161 VDD.n3074 VDD.n3073 10.6151
R6162 VDD.n3073 VDD.n3071 10.6151
R6163 VDD.n3071 VDD.n3070 10.6151
R6164 VDD.n3070 VDD.n3068 10.6151
R6165 VDD.n3068 VDD.n3067 10.6151
R6166 VDD.n3067 VDD.n3065 10.6151
R6167 VDD.n3065 VDD.n3064 10.6151
R6168 VDD.n3064 VDD.n3062 10.6151
R6169 VDD.n3062 VDD.n3061 10.6151
R6170 VDD.n3061 VDD.n3059 10.6151
R6171 VDD.n3059 VDD.n3058 10.6151
R6172 VDD.n3058 VDD.n3056 10.6151
R6173 VDD.n3056 VDD.n3055 10.6151
R6174 VDD.n3055 VDD.n3053 10.6151
R6175 VDD.n3053 VDD.n3052 10.6151
R6176 VDD.n3052 VDD.n3050 10.6151
R6177 VDD.n3050 VDD.n3049 10.6151
R6178 VDD.n3049 VDD.n3047 10.6151
R6179 VDD.n3047 VDD.n3046 10.6151
R6180 VDD.n3046 VDD.n3044 10.6151
R6181 VDD.n3044 VDD.n3043 10.6151
R6182 VDD.n3043 VDD.n3041 10.6151
R6183 VDD.n3041 VDD.n3040 10.6151
R6184 VDD.n3040 VDD.n3038 10.6151
R6185 VDD.n3038 VDD.n3037 10.6151
R6186 VDD.n3037 VDD.n3035 10.6151
R6187 VDD.n3035 VDD.n3034 10.6151
R6188 VDD.n3034 VDD.n3032 10.6151
R6189 VDD.n3032 VDD.n3031 10.6151
R6190 VDD.n3031 VDD.n3029 10.6151
R6191 VDD.n3029 VDD.n3028 10.6151
R6192 VDD.n3028 VDD.n2844 10.6151
R6193 VDD.n2844 VDD.n2843 10.6151
R6194 VDD.n2843 VDD.n2841 10.6151
R6195 VDD.n2841 VDD.n2840 10.6151
R6196 VDD.n2840 VDD.n2838 10.6151
R6197 VDD.n2838 VDD.n2837 10.6151
R6198 VDD.n2837 VDD.n2835 10.6151
R6199 VDD.n2835 VDD.n2834 10.6151
R6200 VDD.n2834 VDD.n2832 10.6151
R6201 VDD.n2832 VDD.n2831 10.6151
R6202 VDD.n2831 VDD.n2829 10.6151
R6203 VDD.n2829 VDD.n2828 10.6151
R6204 VDD.n2828 VDD.n2826 10.6151
R6205 VDD.n2826 VDD.n2825 10.6151
R6206 VDD.n2825 VDD.n2823 10.6151
R6207 VDD.n2823 VDD.n2822 10.6151
R6208 VDD.n2822 VDD.n2820 10.6151
R6209 VDD.n2820 VDD.n2819 10.6151
R6210 VDD.n2819 VDD.n2817 10.6151
R6211 VDD.n2817 VDD.n2816 10.6151
R6212 VDD.n2816 VDD.n2814 10.6151
R6213 VDD.n2814 VDD.n2813 10.6151
R6214 VDD.n2813 VDD.n362 10.6151
R6215 VDD.n3475 VDD.n362 10.6151
R6216 VDD.n3476 VDD.n3475 10.6151
R6217 VDD.n3171 VDD.n3170 10.6151
R6218 VDD.n3170 VDD.n3169 10.6151
R6219 VDD.n3169 VDD.n3168 10.6151
R6220 VDD.n3168 VDD.n3166 10.6151
R6221 VDD.n3166 VDD.n3163 10.6151
R6222 VDD.n3163 VDD.n3162 10.6151
R6223 VDD.n3162 VDD.n3159 10.6151
R6224 VDD.n3159 VDD.n3158 10.6151
R6225 VDD.n3158 VDD.n3155 10.6151
R6226 VDD.n3155 VDD.n3154 10.6151
R6227 VDD.n3154 VDD.n3151 10.6151
R6228 VDD.n3151 VDD.n3150 10.6151
R6229 VDD.n3150 VDD.n3147 10.6151
R6230 VDD.n3147 VDD.n3146 10.6151
R6231 VDD.n3146 VDD.n3143 10.6151
R6232 VDD.n3143 VDD.n3142 10.6151
R6233 VDD.n3142 VDD.n3139 10.6151
R6234 VDD.n3139 VDD.n3138 10.6151
R6235 VDD.n3138 VDD.n3135 10.6151
R6236 VDD.n3135 VDD.n3134 10.6151
R6237 VDD.n3131 VDD.n3130 10.6151
R6238 VDD.n3130 VDD.n3127 10.6151
R6239 VDD.n3127 VDD.n3126 10.6151
R6240 VDD.n3183 VDD.n620 10.6151
R6241 VDD.n3184 VDD.n3183 10.6151
R6242 VDD.n3185 VDD.n3184 10.6151
R6243 VDD.n3185 VDD.n607 10.6151
R6244 VDD.n3195 VDD.n607 10.6151
R6245 VDD.n3196 VDD.n3195 10.6151
R6246 VDD.n3197 VDD.n3196 10.6151
R6247 VDD.n3197 VDD.n596 10.6151
R6248 VDD.n3207 VDD.n596 10.6151
R6249 VDD.n3208 VDD.n3207 10.6151
R6250 VDD.n3209 VDD.n3208 10.6151
R6251 VDD.n3209 VDD.n584 10.6151
R6252 VDD.n3219 VDD.n584 10.6151
R6253 VDD.n3220 VDD.n3219 10.6151
R6254 VDD.n3221 VDD.n3220 10.6151
R6255 VDD.n3221 VDD.n572 10.6151
R6256 VDD.n3231 VDD.n572 10.6151
R6257 VDD.n3232 VDD.n3231 10.6151
R6258 VDD.n3233 VDD.n3232 10.6151
R6259 VDD.n3233 VDD.n560 10.6151
R6260 VDD.n3243 VDD.n560 10.6151
R6261 VDD.n3244 VDD.n3243 10.6151
R6262 VDD.n3245 VDD.n3244 10.6151
R6263 VDD.n3245 VDD.n548 10.6151
R6264 VDD.n3255 VDD.n548 10.6151
R6265 VDD.n3256 VDD.n3255 10.6151
R6266 VDD.n3257 VDD.n3256 10.6151
R6267 VDD.n3257 VDD.n536 10.6151
R6268 VDD.n3267 VDD.n536 10.6151
R6269 VDD.n3268 VDD.n3267 10.6151
R6270 VDD.n3269 VDD.n3268 10.6151
R6271 VDD.n3269 VDD.n524 10.6151
R6272 VDD.n3279 VDD.n524 10.6151
R6273 VDD.n3280 VDD.n3279 10.6151
R6274 VDD.n3281 VDD.n3280 10.6151
R6275 VDD.n3281 VDD.n511 10.6151
R6276 VDD.n3291 VDD.n511 10.6151
R6277 VDD.n3292 VDD.n3291 10.6151
R6278 VDD.n3293 VDD.n3292 10.6151
R6279 VDD.n3293 VDD.n500 10.6151
R6280 VDD.n3303 VDD.n500 10.6151
R6281 VDD.n3304 VDD.n3303 10.6151
R6282 VDD.n3305 VDD.n3304 10.6151
R6283 VDD.n3305 VDD.n488 10.6151
R6284 VDD.n3315 VDD.n488 10.6151
R6285 VDD.n3316 VDD.n3315 10.6151
R6286 VDD.n3317 VDD.n3316 10.6151
R6287 VDD.n3317 VDD.n475 10.6151
R6288 VDD.n3327 VDD.n475 10.6151
R6289 VDD.n3328 VDD.n3327 10.6151
R6290 VDD.n3329 VDD.n3328 10.6151
R6291 VDD.n3329 VDD.n464 10.6151
R6292 VDD.n3339 VDD.n464 10.6151
R6293 VDD.n3340 VDD.n3339 10.6151
R6294 VDD.n3341 VDD.n3340 10.6151
R6295 VDD.n3341 VDD.n452 10.6151
R6296 VDD.n3351 VDD.n452 10.6151
R6297 VDD.n3352 VDD.n3351 10.6151
R6298 VDD.n3353 VDD.n3352 10.6151
R6299 VDD.n3353 VDD.n440 10.6151
R6300 VDD.n3363 VDD.n440 10.6151
R6301 VDD.n3364 VDD.n3363 10.6151
R6302 VDD.n3365 VDD.n3364 10.6151
R6303 VDD.n3365 VDD.n429 10.6151
R6304 VDD.n3375 VDD.n429 10.6151
R6305 VDD.n3376 VDD.n3375 10.6151
R6306 VDD.n3377 VDD.n3376 10.6151
R6307 VDD.n3377 VDD.n417 10.6151
R6308 VDD.n3387 VDD.n417 10.6151
R6309 VDD.n3388 VDD.n3387 10.6151
R6310 VDD.n3389 VDD.n3388 10.6151
R6311 VDD.n3389 VDD.n405 10.6151
R6312 VDD.n3399 VDD.n405 10.6151
R6313 VDD.n3400 VDD.n3399 10.6151
R6314 VDD.n3401 VDD.n3400 10.6151
R6315 VDD.n3401 VDD.n393 10.6151
R6316 VDD.n3411 VDD.n393 10.6151
R6317 VDD.n3412 VDD.n3411 10.6151
R6318 VDD.n3413 VDD.n3412 10.6151
R6319 VDD.n3413 VDD.n381 10.6151
R6320 VDD.n3423 VDD.n381 10.6151
R6321 VDD.n3424 VDD.n3423 10.6151
R6322 VDD.n3425 VDD.n3424 10.6151
R6323 VDD.n3425 VDD.n368 10.6151
R6324 VDD.n3468 VDD.n368 10.6151
R6325 VDD.n3469 VDD.n3468 10.6151
R6326 VDD.n3470 VDD.n3469 10.6151
R6327 VDD.n3470 VDD.n342 10.6151
R6328 VDD.n3521 VDD.n342 10.6151
R6329 VDD.n3520 VDD.n3519 10.6151
R6330 VDD.n3519 VDD.n343 10.6151
R6331 VDD.n344 VDD.n343 10.6151
R6332 VDD.n3512 VDD.n344 10.6151
R6333 VDD.n3512 VDD.n3511 10.6151
R6334 VDD.n3511 VDD.n3510 10.6151
R6335 VDD.n3510 VDD.n346 10.6151
R6336 VDD.n3505 VDD.n346 10.6151
R6337 VDD.n3505 VDD.n3504 10.6151
R6338 VDD.n3504 VDD.n3503 10.6151
R6339 VDD.n3503 VDD.n349 10.6151
R6340 VDD.n349 VDD.n290 10.6151
R6341 VDD.n351 VDD.n290 10.6151
R6342 VDD.n3495 VDD.n351 10.6151
R6343 VDD.n3495 VDD.n3494 10.6151
R6344 VDD.n3494 VDD.n3493 10.6151
R6345 VDD.n3493 VDD.n353 10.6151
R6346 VDD.n3488 VDD.n353 10.6151
R6347 VDD.n3488 VDD.n3487 10.6151
R6348 VDD.n3487 VDD.n3486 10.6151
R6349 VDD.n3481 VDD.n360 10.6151
R6350 VDD.n3481 VDD.n3480 10.6151
R6351 VDD.n3480 VDD.n3479 10.6151
R6352 VDD.n3458 VDD.n3431 10.6151
R6353 VDD.n3453 VDD.n3431 10.6151
R6354 VDD.n3453 VDD.n3452 10.6151
R6355 VDD.n3452 VDD.n3451 10.6151
R6356 VDD.n3451 VDD.n3433 10.6151
R6357 VDD.n3446 VDD.n3433 10.6151
R6358 VDD.n3446 VDD.n3445 10.6151
R6359 VDD.n3445 VDD.n3444 10.6151
R6360 VDD.n3444 VDD.n3436 10.6151
R6361 VDD.n3439 VDD.n3436 10.6151
R6362 VDD.n3439 VDD.n320 10.6151
R6363 VDD.n3547 VDD.n320 10.6151
R6364 VDD.n3547 VDD.n321 10.6151
R6365 VDD.n3542 VDD.n321 10.6151
R6366 VDD.n3542 VDD.n3541 10.6151
R6367 VDD.n3541 VDD.n3540 10.6151
R6368 VDD.n3540 VDD.n325 10.6151
R6369 VDD.n3535 VDD.n325 10.6151
R6370 VDD.n3535 VDD.n3534 10.6151
R6371 VDD.n3534 VDD.n3533 10.6151
R6372 VDD.n3528 VDD.n332 10.6151
R6373 VDD.n3528 VDD.n3527 10.6151
R6374 VDD.n3527 VDD.n3526 10.6151
R6375 VDD.n2895 VDD.n2894 10.6151
R6376 VDD.n2897 VDD.n2895 10.6151
R6377 VDD.n2898 VDD.n2897 10.6151
R6378 VDD.n2900 VDD.n2898 10.6151
R6379 VDD.n2901 VDD.n2900 10.6151
R6380 VDD.n2903 VDD.n2901 10.6151
R6381 VDD.n2904 VDD.n2903 10.6151
R6382 VDD.n2906 VDD.n2904 10.6151
R6383 VDD.n2907 VDD.n2906 10.6151
R6384 VDD.n2909 VDD.n2907 10.6151
R6385 VDD.n2910 VDD.n2909 10.6151
R6386 VDD.n2912 VDD.n2910 10.6151
R6387 VDD.n2913 VDD.n2912 10.6151
R6388 VDD.n2915 VDD.n2913 10.6151
R6389 VDD.n2916 VDD.n2915 10.6151
R6390 VDD.n2918 VDD.n2916 10.6151
R6391 VDD.n2919 VDD.n2918 10.6151
R6392 VDD.n2921 VDD.n2919 10.6151
R6393 VDD.n2922 VDD.n2921 10.6151
R6394 VDD.n2924 VDD.n2922 10.6151
R6395 VDD.n2925 VDD.n2924 10.6151
R6396 VDD.n2927 VDD.n2925 10.6151
R6397 VDD.n2928 VDD.n2927 10.6151
R6398 VDD.n2930 VDD.n2928 10.6151
R6399 VDD.n2931 VDD.n2930 10.6151
R6400 VDD.n2933 VDD.n2931 10.6151
R6401 VDD.n2934 VDD.n2933 10.6151
R6402 VDD.n2936 VDD.n2934 10.6151
R6403 VDD.n2937 VDD.n2936 10.6151
R6404 VDD.n2939 VDD.n2937 10.6151
R6405 VDD.n2940 VDD.n2939 10.6151
R6406 VDD.n2942 VDD.n2940 10.6151
R6407 VDD.n2943 VDD.n2942 10.6151
R6408 VDD.n2945 VDD.n2943 10.6151
R6409 VDD.n2946 VDD.n2945 10.6151
R6410 VDD.n2948 VDD.n2946 10.6151
R6411 VDD.n2949 VDD.n2948 10.6151
R6412 VDD.n2951 VDD.n2949 10.6151
R6413 VDD.n2952 VDD.n2951 10.6151
R6414 VDD.n2954 VDD.n2952 10.6151
R6415 VDD.n2955 VDD.n2954 10.6151
R6416 VDD.n2957 VDD.n2955 10.6151
R6417 VDD.n2958 VDD.n2957 10.6151
R6418 VDD.n2960 VDD.n2958 10.6151
R6419 VDD.n2961 VDD.n2960 10.6151
R6420 VDD.n2963 VDD.n2961 10.6151
R6421 VDD.n2964 VDD.n2963 10.6151
R6422 VDD.n2966 VDD.n2964 10.6151
R6423 VDD.n2967 VDD.n2966 10.6151
R6424 VDD.n2969 VDD.n2967 10.6151
R6425 VDD.n2970 VDD.n2969 10.6151
R6426 VDD.n2972 VDD.n2970 10.6151
R6427 VDD.n2973 VDD.n2972 10.6151
R6428 VDD.n2975 VDD.n2973 10.6151
R6429 VDD.n2976 VDD.n2975 10.6151
R6430 VDD.n2978 VDD.n2976 10.6151
R6431 VDD.n2979 VDD.n2978 10.6151
R6432 VDD.n2981 VDD.n2979 10.6151
R6433 VDD.n2982 VDD.n2981 10.6151
R6434 VDD.n2984 VDD.n2982 10.6151
R6435 VDD.n2985 VDD.n2984 10.6151
R6436 VDD.n2987 VDD.n2985 10.6151
R6437 VDD.n2988 VDD.n2987 10.6151
R6438 VDD.n3024 VDD.n2988 10.6151
R6439 VDD.n3024 VDD.n3023 10.6151
R6440 VDD.n3023 VDD.n3022 10.6151
R6441 VDD.n3022 VDD.n3020 10.6151
R6442 VDD.n3020 VDD.n3019 10.6151
R6443 VDD.n3019 VDD.n3017 10.6151
R6444 VDD.n3017 VDD.n3016 10.6151
R6445 VDD.n3016 VDD.n3014 10.6151
R6446 VDD.n3014 VDD.n3013 10.6151
R6447 VDD.n3013 VDD.n3011 10.6151
R6448 VDD.n3011 VDD.n3010 10.6151
R6449 VDD.n3010 VDD.n3008 10.6151
R6450 VDD.n3008 VDD.n3007 10.6151
R6451 VDD.n3007 VDD.n3005 10.6151
R6452 VDD.n3005 VDD.n3004 10.6151
R6453 VDD.n3004 VDD.n3002 10.6151
R6454 VDD.n3002 VDD.n3001 10.6151
R6455 VDD.n3001 VDD.n2999 10.6151
R6456 VDD.n2999 VDD.n2998 10.6151
R6457 VDD.n2998 VDD.n2996 10.6151
R6458 VDD.n2996 VDD.n2995 10.6151
R6459 VDD.n2995 VDD.n2993 10.6151
R6460 VDD.n2993 VDD.n2992 10.6151
R6461 VDD.n2992 VDD.n2990 10.6151
R6462 VDD.n2990 VDD.n2989 10.6151
R6463 VDD.n2989 VDD.n334 10.6151
R6464 VDD.n3177 VDD.n626 10.6151
R6465 VDD.n2848 VDD.n626 10.6151
R6466 VDD.n2849 VDD.n2848 10.6151
R6467 VDD.n2852 VDD.n2849 10.6151
R6468 VDD.n2853 VDD.n2852 10.6151
R6469 VDD.n2856 VDD.n2853 10.6151
R6470 VDD.n2857 VDD.n2856 10.6151
R6471 VDD.n2860 VDD.n2857 10.6151
R6472 VDD.n2861 VDD.n2860 10.6151
R6473 VDD.n2864 VDD.n2861 10.6151
R6474 VDD.n2865 VDD.n2864 10.6151
R6475 VDD.n2868 VDD.n2865 10.6151
R6476 VDD.n2869 VDD.n2868 10.6151
R6477 VDD.n2872 VDD.n2869 10.6151
R6478 VDD.n2873 VDD.n2872 10.6151
R6479 VDD.n2876 VDD.n2873 10.6151
R6480 VDD.n2877 VDD.n2876 10.6151
R6481 VDD.n2880 VDD.n2877 10.6151
R6482 VDD.n2881 VDD.n2880 10.6151
R6483 VDD.n2884 VDD.n2881 10.6151
R6484 VDD.n2889 VDD.n2886 10.6151
R6485 VDD.n2891 VDD.n2889 10.6151
R6486 VDD.n2892 VDD.n2891 10.6151
R6487 VDD.n3179 VDD.n3178 10.6151
R6488 VDD.n3179 VDD.n614 10.6151
R6489 VDD.n3189 VDD.n614 10.6151
R6490 VDD.n3190 VDD.n3189 10.6151
R6491 VDD.n3191 VDD.n3190 10.6151
R6492 VDD.n3191 VDD.n601 10.6151
R6493 VDD.n3201 VDD.n601 10.6151
R6494 VDD.n3202 VDD.n3201 10.6151
R6495 VDD.n3203 VDD.n3202 10.6151
R6496 VDD.n3203 VDD.n590 10.6151
R6497 VDD.n3213 VDD.n590 10.6151
R6498 VDD.n3214 VDD.n3213 10.6151
R6499 VDD.n3215 VDD.n3214 10.6151
R6500 VDD.n3215 VDD.n578 10.6151
R6501 VDD.n3225 VDD.n578 10.6151
R6502 VDD.n3226 VDD.n3225 10.6151
R6503 VDD.n3227 VDD.n3226 10.6151
R6504 VDD.n3227 VDD.n566 10.6151
R6505 VDD.n3237 VDD.n566 10.6151
R6506 VDD.n3238 VDD.n3237 10.6151
R6507 VDD.n3239 VDD.n3238 10.6151
R6508 VDD.n3239 VDD.n554 10.6151
R6509 VDD.n3249 VDD.n554 10.6151
R6510 VDD.n3250 VDD.n3249 10.6151
R6511 VDD.n3251 VDD.n3250 10.6151
R6512 VDD.n3251 VDD.n542 10.6151
R6513 VDD.n3261 VDD.n542 10.6151
R6514 VDD.n3262 VDD.n3261 10.6151
R6515 VDD.n3263 VDD.n3262 10.6151
R6516 VDD.n3263 VDD.n529 10.6151
R6517 VDD.n3273 VDD.n529 10.6151
R6518 VDD.n3274 VDD.n3273 10.6151
R6519 VDD.n3275 VDD.n3274 10.6151
R6520 VDD.n3275 VDD.n518 10.6151
R6521 VDD.n3285 VDD.n518 10.6151
R6522 VDD.n3286 VDD.n3285 10.6151
R6523 VDD.n3287 VDD.n3286 10.6151
R6524 VDD.n3287 VDD.n506 10.6151
R6525 VDD.n3297 VDD.n506 10.6151
R6526 VDD.n3298 VDD.n3297 10.6151
R6527 VDD.n3299 VDD.n3298 10.6151
R6528 VDD.n3299 VDD.n494 10.6151
R6529 VDD.n3309 VDD.n494 10.6151
R6530 VDD.n3310 VDD.n3309 10.6151
R6531 VDD.n3311 VDD.n3310 10.6151
R6532 VDD.n3311 VDD.n482 10.6151
R6533 VDD.n3321 VDD.n482 10.6151
R6534 VDD.n3322 VDD.n3321 10.6151
R6535 VDD.n3323 VDD.n3322 10.6151
R6536 VDD.n3323 VDD.n470 10.6151
R6537 VDD.n3333 VDD.n470 10.6151
R6538 VDD.n3334 VDD.n3333 10.6151
R6539 VDD.n3335 VDD.n3334 10.6151
R6540 VDD.n3335 VDD.n458 10.6151
R6541 VDD.n3345 VDD.n458 10.6151
R6542 VDD.n3346 VDD.n3345 10.6151
R6543 VDD.n3347 VDD.n3346 10.6151
R6544 VDD.n3347 VDD.n446 10.6151
R6545 VDD.n3357 VDD.n446 10.6151
R6546 VDD.n3358 VDD.n3357 10.6151
R6547 VDD.n3359 VDD.n3358 10.6151
R6548 VDD.n3359 VDD.n434 10.6151
R6549 VDD.n3369 VDD.n434 10.6151
R6550 VDD.n3370 VDD.n3369 10.6151
R6551 VDD.n3371 VDD.n3370 10.6151
R6552 VDD.n3371 VDD.n423 10.6151
R6553 VDD.n3381 VDD.n423 10.6151
R6554 VDD.n3382 VDD.n3381 10.6151
R6555 VDD.n3383 VDD.n3382 10.6151
R6556 VDD.n3383 VDD.n411 10.6151
R6557 VDD.n3393 VDD.n411 10.6151
R6558 VDD.n3394 VDD.n3393 10.6151
R6559 VDD.n3395 VDD.n3394 10.6151
R6560 VDD.n3395 VDD.n399 10.6151
R6561 VDD.n3405 VDD.n399 10.6151
R6562 VDD.n3406 VDD.n3405 10.6151
R6563 VDD.n3407 VDD.n3406 10.6151
R6564 VDD.n3407 VDD.n386 10.6151
R6565 VDD.n3417 VDD.n386 10.6151
R6566 VDD.n3418 VDD.n3417 10.6151
R6567 VDD.n3419 VDD.n3418 10.6151
R6568 VDD.n3419 VDD.n375 10.6151
R6569 VDD.n3429 VDD.n375 10.6151
R6570 VDD.n3430 VDD.n3429 10.6151
R6571 VDD.n3464 VDD.n3430 10.6151
R6572 VDD.n3464 VDD.n3463 10.6151
R6573 VDD.n3463 VDD.n3462 10.6151
R6574 VDD.n3462 VDD.n3461 10.6151
R6575 VDD.n3461 VDD.n3459 10.6151
R6576 VDD.n2409 VDD.n2408 10.6151
R6577 VDD.n2410 VDD.n2409 10.6151
R6578 VDD.n2410 VDD.n917 10.6151
R6579 VDD.n2420 VDD.n917 10.6151
R6580 VDD.n2421 VDD.n2420 10.6151
R6581 VDD.n2422 VDD.n2421 10.6151
R6582 VDD.n2422 VDD.n905 10.6151
R6583 VDD.n2432 VDD.n905 10.6151
R6584 VDD.n2433 VDD.n2432 10.6151
R6585 VDD.n2434 VDD.n2433 10.6151
R6586 VDD.n2434 VDD.n893 10.6151
R6587 VDD.n2444 VDD.n893 10.6151
R6588 VDD.n2445 VDD.n2444 10.6151
R6589 VDD.n2446 VDD.n2445 10.6151
R6590 VDD.n2446 VDD.n881 10.6151
R6591 VDD.n2456 VDD.n881 10.6151
R6592 VDD.n2457 VDD.n2456 10.6151
R6593 VDD.n2458 VDD.n2457 10.6151
R6594 VDD.n2458 VDD.n869 10.6151
R6595 VDD.n2468 VDD.n869 10.6151
R6596 VDD.n2469 VDD.n2468 10.6151
R6597 VDD.n2470 VDD.n2469 10.6151
R6598 VDD.n2470 VDD.n857 10.6151
R6599 VDD.n2480 VDD.n857 10.6151
R6600 VDD.n2481 VDD.n2480 10.6151
R6601 VDD.n2482 VDD.n2481 10.6151
R6602 VDD.n2482 VDD.n846 10.6151
R6603 VDD.n2492 VDD.n846 10.6151
R6604 VDD.n2493 VDD.n2492 10.6151
R6605 VDD.n2494 VDD.n2493 10.6151
R6606 VDD.n2494 VDD.n834 10.6151
R6607 VDD.n2504 VDD.n834 10.6151
R6608 VDD.n2505 VDD.n2504 10.6151
R6609 VDD.n2506 VDD.n2505 10.6151
R6610 VDD.n2506 VDD.n822 10.6151
R6611 VDD.n2516 VDD.n822 10.6151
R6612 VDD.n2517 VDD.n2516 10.6151
R6613 VDD.n2518 VDD.n2517 10.6151
R6614 VDD.n2518 VDD.n810 10.6151
R6615 VDD.n2528 VDD.n810 10.6151
R6616 VDD.n2529 VDD.n2528 10.6151
R6617 VDD.n2530 VDD.n2529 10.6151
R6618 VDD.n2530 VDD.n798 10.6151
R6619 VDD.n2540 VDD.n798 10.6151
R6620 VDD.n2541 VDD.n2540 10.6151
R6621 VDD.n2542 VDD.n2541 10.6151
R6622 VDD.n2542 VDD.n786 10.6151
R6623 VDD.n2552 VDD.n786 10.6151
R6624 VDD.n2553 VDD.n2552 10.6151
R6625 VDD.n2554 VDD.n2553 10.6151
R6626 VDD.n2554 VDD.n774 10.6151
R6627 VDD.n2564 VDD.n774 10.6151
R6628 VDD.n2565 VDD.n2564 10.6151
R6629 VDD.n2566 VDD.n2565 10.6151
R6630 VDD.n2566 VDD.n762 10.6151
R6631 VDD.n2576 VDD.n762 10.6151
R6632 VDD.n2577 VDD.n2576 10.6151
R6633 VDD.n2578 VDD.n2577 10.6151
R6634 VDD.n2578 VDD.n750 10.6151
R6635 VDD.n2588 VDD.n750 10.6151
R6636 VDD.n2589 VDD.n2588 10.6151
R6637 VDD.n2590 VDD.n2589 10.6151
R6638 VDD.n2590 VDD.n738 10.6151
R6639 VDD.n2600 VDD.n738 10.6151
R6640 VDD.n2601 VDD.n2600 10.6151
R6641 VDD.n2602 VDD.n2601 10.6151
R6642 VDD.n2602 VDD.n725 10.6151
R6643 VDD.n2612 VDD.n725 10.6151
R6644 VDD.n2613 VDD.n2612 10.6151
R6645 VDD.n2614 VDD.n2613 10.6151
R6646 VDD.n2614 VDD.n714 10.6151
R6647 VDD.n2624 VDD.n714 10.6151
R6648 VDD.n2625 VDD.n2624 10.6151
R6649 VDD.n2626 VDD.n2625 10.6151
R6650 VDD.n2626 VDD.n702 10.6151
R6651 VDD.n2636 VDD.n702 10.6151
R6652 VDD.n2637 VDD.n2636 10.6151
R6653 VDD.n2638 VDD.n2637 10.6151
R6654 VDD.n2638 VDD.n690 10.6151
R6655 VDD.n2648 VDD.n690 10.6151
R6656 VDD.n2649 VDD.n2648 10.6151
R6657 VDD.n2652 VDD.n2649 10.6151
R6658 VDD.n2652 VDD.n2651 10.6151
R6659 VDD.n2651 VDD.n2650 10.6151
R6660 VDD.n2650 VDD.n674 10.6151
R6661 VDD.n2724 VDD.n674 10.6151
R6662 VDD.n2724 VDD.n2723 10.6151
R6663 VDD.n2723 VDD.n2722 10.6151
R6664 VDD.n2722 VDD.n2721 10.6151
R6665 VDD.n2718 VDD.n2717 10.6151
R6666 VDD.n2717 VDD.n2714 10.6151
R6667 VDD.n2714 VDD.n2713 10.6151
R6668 VDD.n2713 VDD.n2710 10.6151
R6669 VDD.n2710 VDD.n2709 10.6151
R6670 VDD.n2709 VDD.n2706 10.6151
R6671 VDD.n2706 VDD.n2705 10.6151
R6672 VDD.n2705 VDD.n2702 10.6151
R6673 VDD.n2702 VDD.n2701 10.6151
R6674 VDD.n2701 VDD.n2698 10.6151
R6675 VDD.n2698 VDD.n2697 10.6151
R6676 VDD.n2697 VDD.n2694 10.6151
R6677 VDD.n2694 VDD.n2693 10.6151
R6678 VDD.n2693 VDD.n2690 10.6151
R6679 VDD.n2690 VDD.n2689 10.6151
R6680 VDD.n2689 VDD.n2686 10.6151
R6681 VDD.n2686 VDD.n2685 10.6151
R6682 VDD.n2685 VDD.n2682 10.6151
R6683 VDD.n2682 VDD.n2681 10.6151
R6684 VDD.n2681 VDD.n2678 10.6151
R6685 VDD.n2676 VDD.n2673 10.6151
R6686 VDD.n2673 VDD.n2672 10.6151
R6687 VDD.n2672 VDD.n2670 10.6151
R6688 VDD.n2396 VDD.n2395 10.6151
R6689 VDD.n2395 VDD.n2393 10.6151
R6690 VDD.n2393 VDD.n2392 10.6151
R6691 VDD.n2392 VDD.n2390 10.6151
R6692 VDD.n2390 VDD.n2389 10.6151
R6693 VDD.n2389 VDD.n2387 10.6151
R6694 VDD.n2387 VDD.n2386 10.6151
R6695 VDD.n2386 VDD.n2384 10.6151
R6696 VDD.n2384 VDD.n2383 10.6151
R6697 VDD.n2383 VDD.n2381 10.6151
R6698 VDD.n2381 VDD.n2380 10.6151
R6699 VDD.n2380 VDD.n2378 10.6151
R6700 VDD.n2378 VDD.n2377 10.6151
R6701 VDD.n2377 VDD.n2375 10.6151
R6702 VDD.n2375 VDD.n2374 10.6151
R6703 VDD.n2374 VDD.n2372 10.6151
R6704 VDD.n2372 VDD.n2371 10.6151
R6705 VDD.n2371 VDD.n2369 10.6151
R6706 VDD.n2369 VDD.n2368 10.6151
R6707 VDD.n2368 VDD.n2366 10.6151
R6708 VDD.n2366 VDD.n2365 10.6151
R6709 VDD.n2365 VDD.n2363 10.6151
R6710 VDD.n2363 VDD.n2362 10.6151
R6711 VDD.n2362 VDD.n2360 10.6151
R6712 VDD.n2360 VDD.n2359 10.6151
R6713 VDD.n2359 VDD.n1046 10.6151
R6714 VDD.n1046 VDD.n1045 10.6151
R6715 VDD.n1045 VDD.n1043 10.6151
R6716 VDD.n1043 VDD.n1042 10.6151
R6717 VDD.n1042 VDD.n1040 10.6151
R6718 VDD.n1040 VDD.n1039 10.6151
R6719 VDD.n1039 VDD.n1037 10.6151
R6720 VDD.n1037 VDD.n1036 10.6151
R6721 VDD.n1036 VDD.n1034 10.6151
R6722 VDD.n1034 VDD.n1033 10.6151
R6723 VDD.n1033 VDD.n1031 10.6151
R6724 VDD.n1031 VDD.n1030 10.6151
R6725 VDD.n1030 VDD.n1028 10.6151
R6726 VDD.n1028 VDD.n1027 10.6151
R6727 VDD.n1027 VDD.n1025 10.6151
R6728 VDD.n1025 VDD.n1024 10.6151
R6729 VDD.n1024 VDD.n1022 10.6151
R6730 VDD.n1022 VDD.n1021 10.6151
R6731 VDD.n1021 VDD.n1019 10.6151
R6732 VDD.n1019 VDD.n1018 10.6151
R6733 VDD.n1018 VDD.n1016 10.6151
R6734 VDD.n1016 VDD.n1015 10.6151
R6735 VDD.n1015 VDD.n1013 10.6151
R6736 VDD.n1013 VDD.n1012 10.6151
R6737 VDD.n1012 VDD.n1010 10.6151
R6738 VDD.n1010 VDD.n1009 10.6151
R6739 VDD.n1009 VDD.n1007 10.6151
R6740 VDD.n1007 VDD.n1006 10.6151
R6741 VDD.n1006 VDD.n1004 10.6151
R6742 VDD.n1004 VDD.n1003 10.6151
R6743 VDD.n1003 VDD.n1001 10.6151
R6744 VDD.n1001 VDD.n1000 10.6151
R6745 VDD.n1000 VDD.n998 10.6151
R6746 VDD.n998 VDD.n997 10.6151
R6747 VDD.n997 VDD.n995 10.6151
R6748 VDD.n995 VDD.n994 10.6151
R6749 VDD.n994 VDD.n992 10.6151
R6750 VDD.n992 VDD.n991 10.6151
R6751 VDD.n991 VDD.n989 10.6151
R6752 VDD.n989 VDD.n988 10.6151
R6753 VDD.n988 VDD.n986 10.6151
R6754 VDD.n986 VDD.n985 10.6151
R6755 VDD.n985 VDD.n983 10.6151
R6756 VDD.n983 VDD.n982 10.6151
R6757 VDD.n982 VDD.n980 10.6151
R6758 VDD.n980 VDD.n979 10.6151
R6759 VDD.n979 VDD.n977 10.6151
R6760 VDD.n977 VDD.n976 10.6151
R6761 VDD.n976 VDD.n974 10.6151
R6762 VDD.n974 VDD.n973 10.6151
R6763 VDD.n973 VDD.n971 10.6151
R6764 VDD.n971 VDD.n970 10.6151
R6765 VDD.n970 VDD.n968 10.6151
R6766 VDD.n968 VDD.n967 10.6151
R6767 VDD.n967 VDD.n965 10.6151
R6768 VDD.n965 VDD.n964 10.6151
R6769 VDD.n964 VDD.n962 10.6151
R6770 VDD.n962 VDD.n961 10.6151
R6771 VDD.n961 VDD.n677 10.6151
R6772 VDD.n2663 VDD.n677 10.6151
R6773 VDD.n2664 VDD.n2663 10.6151
R6774 VDD.n2666 VDD.n2664 10.6151
R6775 VDD.n2667 VDD.n2666 10.6151
R6776 VDD.n2669 VDD.n2667 10.6151
R6777 VDD.n1147 VDD.n929 10.6151
R6778 VDD.n1150 VDD.n1147 10.6151
R6779 VDD.n1151 VDD.n1150 10.6151
R6780 VDD.n1154 VDD.n1151 10.6151
R6781 VDD.n1155 VDD.n1154 10.6151
R6782 VDD.n1158 VDD.n1155 10.6151
R6783 VDD.n1159 VDD.n1158 10.6151
R6784 VDD.n1162 VDD.n1159 10.6151
R6785 VDD.n1163 VDD.n1162 10.6151
R6786 VDD.n1166 VDD.n1163 10.6151
R6787 VDD.n1167 VDD.n1166 10.6151
R6788 VDD.n1193 VDD.n1167 10.6151
R6789 VDD.n1193 VDD.n1192 10.6151
R6790 VDD.n1192 VDD.n1189 10.6151
R6791 VDD.n1189 VDD.n1188 10.6151
R6792 VDD.n1188 VDD.n1185 10.6151
R6793 VDD.n1185 VDD.n1184 10.6151
R6794 VDD.n1184 VDD.n1181 10.6151
R6795 VDD.n1181 VDD.n1180 10.6151
R6796 VDD.n1180 VDD.n1177 10.6151
R6797 VDD.n1175 VDD.n1172 10.6151
R6798 VDD.n1172 VDD.n960 10.6151
R6799 VDD.n2397 VDD.n960 10.6151
R6800 VDD.n2200 VDD.n2199 10.3189
R6801 VDD.n3693 VDD.n290 10.3189
R6802 VDD.n3548 VDD.n3547 10.3189
R6803 VDD.n2102 VDD.n1193 10.3189
R6804 VDD.n2406 VDD.n925 9.71771
R6805 VDD.n2412 VDD.n925 9.71771
R6806 VDD.n2412 VDD.n919 9.71771
R6807 VDD.n2418 VDD.n919 9.71771
R6808 VDD.n2418 VDD.n913 9.71771
R6809 VDD.n2424 VDD.n913 9.71771
R6810 VDD.n2424 VDD.n907 9.71771
R6811 VDD.n2430 VDD.n907 9.71771
R6812 VDD.n2436 VDD.n900 9.71771
R6813 VDD.n2436 VDD.n903 9.71771
R6814 VDD.n2442 VDD.n889 9.71771
R6815 VDD.n2448 VDD.n889 9.71771
R6816 VDD.n2448 VDD.n883 9.71771
R6817 VDD.n2454 VDD.n883 9.71771
R6818 VDD.n2454 VDD.n877 9.71771
R6819 VDD.n2460 VDD.n877 9.71771
R6820 VDD.n2460 VDD.n871 9.71771
R6821 VDD.n2466 VDD.n871 9.71771
R6822 VDD.n2466 VDD.n865 9.71771
R6823 VDD.n2472 VDD.n865 9.71771
R6824 VDD.n2472 VDD.n859 9.71771
R6825 VDD.n2478 VDD.n859 9.71771
R6826 VDD.n2484 VDD.n848 9.71771
R6827 VDD.n2490 VDD.n848 9.71771
R6828 VDD.n2490 VDD.n842 9.71771
R6829 VDD.n2496 VDD.n842 9.71771
R6830 VDD.n2496 VDD.n836 9.71771
R6831 VDD.n2502 VDD.n836 9.71771
R6832 VDD.n2502 VDD.n830 9.71771
R6833 VDD.n2508 VDD.n830 9.71771
R6834 VDD.n2508 VDD.n824 9.71771
R6835 VDD.n2514 VDD.n824 9.71771
R6836 VDD.n2514 VDD.n818 9.71771
R6837 VDD.n2520 VDD.n818 9.71771
R6838 VDD.n2526 VDD.n812 9.71771
R6839 VDD.n2526 VDD.n805 9.71771
R6840 VDD.n2532 VDD.n805 9.71771
R6841 VDD.n2532 VDD.n808 9.71771
R6842 VDD.n2538 VDD.n794 9.71771
R6843 VDD.n2544 VDD.n794 9.71771
R6844 VDD.n2544 VDD.n788 9.71771
R6845 VDD.n2550 VDD.n788 9.71771
R6846 VDD.n2550 VDD.n782 9.71771
R6847 VDD.n2556 VDD.n782 9.71771
R6848 VDD.n2562 VDD.n776 9.71771
R6849 VDD.n2562 VDD.n770 9.71771
R6850 VDD.n2568 VDD.n770 9.71771
R6851 VDD.n2568 VDD.n764 9.71771
R6852 VDD.n2574 VDD.n764 9.71771
R6853 VDD.n2580 VDD.n758 9.71771
R6854 VDD.n2580 VDD.n752 9.71771
R6855 VDD.n2586 VDD.n752 9.71771
R6856 VDD.n2586 VDD.n745 9.71771
R6857 VDD.n2592 VDD.n745 9.71771
R6858 VDD.n2592 VDD.n748 9.71771
R6859 VDD.n2598 VDD.n734 9.71771
R6860 VDD.n2604 VDD.n734 9.71771
R6861 VDD.n2604 VDD.n727 9.71771
R6862 VDD.n2610 VDD.n727 9.71771
R6863 VDD.n2610 VDD.n730 9.71771
R6864 VDD.n2616 VDD.n716 9.71771
R6865 VDD.n2622 VDD.n716 9.71771
R6866 VDD.n2622 VDD.n710 9.71771
R6867 VDD.n2628 VDD.n710 9.71771
R6868 VDD.n2628 VDD.n704 9.71771
R6869 VDD.n2634 VDD.n704 9.71771
R6870 VDD.n2634 VDD.n698 9.71771
R6871 VDD.n2640 VDD.n698 9.71771
R6872 VDD.n2640 VDD.n692 9.71771
R6873 VDD.n2646 VDD.n692 9.71771
R6874 VDD.n2654 VDD.n685 9.71771
R6875 VDD.n2660 VDD.n679 9.71771
R6876 VDD.n2660 VDD.n669 9.71771
R6877 VDD.n2726 VDD.n669 9.71771
R6878 VDD.n2726 VDD.n663 9.71771
R6879 VDD.n2732 VDD.n663 9.71771
R6880 VDD.n2732 VDD.n628 9.71771
R6881 VDD.n3181 VDD.n622 9.71771
R6882 VDD.n3181 VDD.n616 9.71771
R6883 VDD.n3187 VDD.n616 9.71771
R6884 VDD.n3187 VDD.n609 9.71771
R6885 VDD.n3193 VDD.n609 9.71771
R6886 VDD.n3193 VDD.n612 9.71771
R6887 VDD.n3199 VDD.n605 9.71771
R6888 VDD.n3205 VDD.n592 9.71771
R6889 VDD.n3211 VDD.n592 9.71771
R6890 VDD.n3211 VDD.n586 9.71771
R6891 VDD.n3217 VDD.n586 9.71771
R6892 VDD.n3217 VDD.n580 9.71771
R6893 VDD.n3223 VDD.n580 9.71771
R6894 VDD.n3223 VDD.n574 9.71771
R6895 VDD.n3229 VDD.n574 9.71771
R6896 VDD.n3229 VDD.n568 9.71771
R6897 VDD.n3235 VDD.n568 9.71771
R6898 VDD.n3241 VDD.n562 9.71771
R6899 VDD.n3241 VDD.n556 9.71771
R6900 VDD.n3247 VDD.n556 9.71771
R6901 VDD.n3247 VDD.n550 9.71771
R6902 VDD.n3253 VDD.n550 9.71771
R6903 VDD.n3259 VDD.n544 9.71771
R6904 VDD.n3259 VDD.n538 9.71771
R6905 VDD.n3265 VDD.n538 9.71771
R6906 VDD.n3265 VDD.n531 9.71771
R6907 VDD.n3271 VDD.n531 9.71771
R6908 VDD.n3271 VDD.n534 9.71771
R6909 VDD.n3277 VDD.n520 9.71771
R6910 VDD.n3283 VDD.n520 9.71771
R6911 VDD.n3283 VDD.n513 9.71771
R6912 VDD.n3289 VDD.n513 9.71771
R6913 VDD.n3289 VDD.n516 9.71771
R6914 VDD.n3295 VDD.n502 9.71771
R6915 VDD.n3301 VDD.n502 9.71771
R6916 VDD.n3301 VDD.n496 9.71771
R6917 VDD.n3307 VDD.n496 9.71771
R6918 VDD.n3307 VDD.n490 9.71771
R6919 VDD.n3313 VDD.n490 9.71771
R6920 VDD.n3319 VDD.n484 9.71771
R6921 VDD.n3319 VDD.n477 9.71771
R6922 VDD.n3325 VDD.n477 9.71771
R6923 VDD.n3325 VDD.n480 9.71771
R6924 VDD.n3331 VDD.n466 9.71771
R6925 VDD.n3337 VDD.n466 9.71771
R6926 VDD.n3337 VDD.n460 9.71771
R6927 VDD.n3343 VDD.n460 9.71771
R6928 VDD.n3343 VDD.n454 9.71771
R6929 VDD.n3349 VDD.n454 9.71771
R6930 VDD.n3349 VDD.n448 9.71771
R6931 VDD.n3355 VDD.n448 9.71771
R6932 VDD.n3355 VDD.n442 9.71771
R6933 VDD.n3361 VDD.n442 9.71771
R6934 VDD.n3361 VDD.n436 9.71771
R6935 VDD.n3367 VDD.n436 9.71771
R6936 VDD.n3373 VDD.n425 9.71771
R6937 VDD.n3379 VDD.n425 9.71771
R6938 VDD.n3379 VDD.n419 9.71771
R6939 VDD.n3385 VDD.n419 9.71771
R6940 VDD.n3385 VDD.n413 9.71771
R6941 VDD.n3391 VDD.n413 9.71771
R6942 VDD.n3391 VDD.n407 9.71771
R6943 VDD.n3397 VDD.n407 9.71771
R6944 VDD.n3397 VDD.n401 9.71771
R6945 VDD.n3403 VDD.n401 9.71771
R6946 VDD.n3403 VDD.n395 9.71771
R6947 VDD.n3409 VDD.n395 9.71771
R6948 VDD.n3415 VDD.n388 9.71771
R6949 VDD.n3415 VDD.n391 9.71771
R6950 VDD.n3421 VDD.n377 9.71771
R6951 VDD.n3427 VDD.n377 9.71771
R6952 VDD.n3427 VDD.n370 9.71771
R6953 VDD.n3466 VDD.n370 9.71771
R6954 VDD.n3466 VDD.n364 9.71771
R6955 VDD.n3472 VDD.n364 9.71771
R6956 VDD.n3472 VDD.n337 9.71771
R6957 VDD.n3523 VDD.n337 9.71771
R6958 VDD.n2406 VDD.t140 9.43191
R6959 VDD.n3523 VDD.t130 9.43191
R6960 VDD.n2165 VDD.n1110 9.3005
R6961 VDD.n2164 VDD.n2163 9.3005
R6962 VDD.n2160 VDD.n1115 9.3005
R6963 VDD.n2159 VDD.n1116 9.3005
R6964 VDD.n2156 VDD.n1117 9.3005
R6965 VDD.n2155 VDD.n1118 9.3005
R6966 VDD.n2152 VDD.n1119 9.3005
R6967 VDD.n2151 VDD.n1120 9.3005
R6968 VDD.n2148 VDD.n1121 9.3005
R6969 VDD.n2147 VDD.n1122 9.3005
R6970 VDD.n2144 VDD.n1123 9.3005
R6971 VDD.n2143 VDD.n1124 9.3005
R6972 VDD.n2140 VDD.n1125 9.3005
R6973 VDD.n2139 VDD.n1126 9.3005
R6974 VDD.n2136 VDD.n1127 9.3005
R6975 VDD.n2135 VDD.n1128 9.3005
R6976 VDD.n2132 VDD.n1132 9.3005
R6977 VDD.n2131 VDD.n1133 9.3005
R6978 VDD.n2128 VDD.n1134 9.3005
R6979 VDD.n2127 VDD.n1135 9.3005
R6980 VDD.n2124 VDD.n1136 9.3005
R6981 VDD.n2123 VDD.n1137 9.3005
R6982 VDD.n2120 VDD.n1138 9.3005
R6983 VDD.n2119 VDD.n1139 9.3005
R6984 VDD.n2116 VDD.n1140 9.3005
R6985 VDD.n2115 VDD.n1141 9.3005
R6986 VDD.n2112 VDD.n1142 9.3005
R6987 VDD.n2111 VDD.n1143 9.3005
R6988 VDD.n2108 VDD.n1144 9.3005
R6989 VDD.n2107 VDD.n1145 9.3005
R6990 VDD.n2167 VDD.n2166 9.3005
R6991 VDD.n2187 VDD.n1068 9.3005
R6992 VDD.n2184 VDD.n1101 9.3005
R6993 VDD.n2183 VDD.n1102 9.3005
R6994 VDD.n2180 VDD.n1103 9.3005
R6995 VDD.n2179 VDD.n1104 9.3005
R6996 VDD.n2176 VDD.n1105 9.3005
R6997 VDD.n2175 VDD.n1106 9.3005
R6998 VDD.n2172 VDD.n1107 9.3005
R6999 VDD.n2171 VDD.n1108 9.3005
R7000 VDD.n2168 VDD.n1109 9.3005
R7001 VDD.n1899 VDD.n1898 9.3005
R7002 VDD.n1339 VDD.n1338 9.3005
R7003 VDD.n1912 VDD.n1911 9.3005
R7004 VDD.n1913 VDD.n1337 9.3005
R7005 VDD.n1915 VDD.n1914 9.3005
R7006 VDD.n1327 VDD.n1326 9.3005
R7007 VDD.n1928 VDD.n1927 9.3005
R7008 VDD.n1929 VDD.n1325 9.3005
R7009 VDD.n1931 VDD.n1930 9.3005
R7010 VDD.n1315 VDD.n1314 9.3005
R7011 VDD.n1944 VDD.n1943 9.3005
R7012 VDD.n1945 VDD.n1313 9.3005
R7013 VDD.n1947 VDD.n1946 9.3005
R7014 VDD.n1303 VDD.n1302 9.3005
R7015 VDD.n1960 VDD.n1959 9.3005
R7016 VDD.n1961 VDD.n1301 9.3005
R7017 VDD.n1963 VDD.n1962 9.3005
R7018 VDD.n1291 VDD.n1290 9.3005
R7019 VDD.n1976 VDD.n1975 9.3005
R7020 VDD.n1977 VDD.n1289 9.3005
R7021 VDD.n1979 VDD.n1978 9.3005
R7022 VDD.n1279 VDD.n1278 9.3005
R7023 VDD.n1992 VDD.n1991 9.3005
R7024 VDD.n1993 VDD.n1277 9.3005
R7025 VDD.n1995 VDD.n1994 9.3005
R7026 VDD.n1267 VDD.n1266 9.3005
R7027 VDD.n2008 VDD.n2007 9.3005
R7028 VDD.n2009 VDD.n1265 9.3005
R7029 VDD.n2011 VDD.n2010 9.3005
R7030 VDD.n1256 VDD.n1255 9.3005
R7031 VDD.n2024 VDD.n2023 9.3005
R7032 VDD.n2025 VDD.n1254 9.3005
R7033 VDD.n2027 VDD.n2026 9.3005
R7034 VDD.n1244 VDD.n1243 9.3005
R7035 VDD.n2040 VDD.n2039 9.3005
R7036 VDD.n2041 VDD.n1242 9.3005
R7037 VDD.n2043 VDD.n2042 9.3005
R7038 VDD.n1232 VDD.n1231 9.3005
R7039 VDD.n2056 VDD.n2055 9.3005
R7040 VDD.n2057 VDD.n1230 9.3005
R7041 VDD.n2059 VDD.n2058 9.3005
R7042 VDD.n1220 VDD.n1219 9.3005
R7043 VDD.n2073 VDD.n2072 9.3005
R7044 VDD.n2074 VDD.n1218 9.3005
R7045 VDD.n2076 VDD.n2075 9.3005
R7046 VDD.n1208 VDD.n1207 9.3005
R7047 VDD.n2091 VDD.n2090 9.3005
R7048 VDD.n2092 VDD.n1206 9.3005
R7049 VDD.n2094 VDD.n2093 9.3005
R7050 VDD.n1072 VDD.n1071 9.3005
R7051 VDD.n2198 VDD.n2197 9.3005
R7052 VDD.n3701 VDD.n3700 9.3005
R7053 VDD.n3702 VDD.n283 9.3005
R7054 VDD.n3704 VDD.n3703 9.3005
R7055 VDD.n272 VDD.n271 9.3005
R7056 VDD.n3717 VDD.n3716 9.3005
R7057 VDD.n3718 VDD.n270 9.3005
R7058 VDD.n3720 VDD.n3719 9.3005
R7059 VDD.n261 VDD.n260 9.3005
R7060 VDD.n3733 VDD.n3732 9.3005
R7061 VDD.n3734 VDD.n259 9.3005
R7062 VDD.n3736 VDD.n3735 9.3005
R7063 VDD.n249 VDD.n248 9.3005
R7064 VDD.n3749 VDD.n3748 9.3005
R7065 VDD.n3750 VDD.n247 9.3005
R7066 VDD.n3752 VDD.n3751 9.3005
R7067 VDD.n237 VDD.n236 9.3005
R7068 VDD.n3765 VDD.n3764 9.3005
R7069 VDD.n3766 VDD.n235 9.3005
R7070 VDD.n3768 VDD.n3767 9.3005
R7071 VDD.n225 VDD.n224 9.3005
R7072 VDD.n3780 VDD.n3779 9.3005
R7073 VDD.n3781 VDD.n223 9.3005
R7074 VDD.n3783 VDD.n3782 9.3005
R7075 VDD.n213 VDD.n212 9.3005
R7076 VDD.n3796 VDD.n3795 9.3005
R7077 VDD.n3797 VDD.n211 9.3005
R7078 VDD.n3799 VDD.n3798 9.3005
R7079 VDD.n201 VDD.n200 9.3005
R7080 VDD.n3812 VDD.n3811 9.3005
R7081 VDD.n3813 VDD.n199 9.3005
R7082 VDD.n3815 VDD.n3814 9.3005
R7083 VDD.n190 VDD.n189 9.3005
R7084 VDD.n3829 VDD.n3828 9.3005
R7085 VDD.n3830 VDD.n188 9.3005
R7086 VDD.n3832 VDD.n3831 9.3005
R7087 VDD.n178 VDD.n177 9.3005
R7088 VDD.n3845 VDD.n3844 9.3005
R7089 VDD.n3846 VDD.n176 9.3005
R7090 VDD.n3848 VDD.n3847 9.3005
R7091 VDD.n166 VDD.n165 9.3005
R7092 VDD.n3861 VDD.n3860 9.3005
R7093 VDD.n3862 VDD.n164 9.3005
R7094 VDD.n3866 VDD.n3863 9.3005
R7095 VDD.n3865 VDD.n3864 9.3005
R7096 VDD.n155 VDD.n154 9.3005
R7097 VDD.n3881 VDD.n3880 9.3005
R7098 VDD.n3882 VDD.n153 9.3005
R7099 VDD.n3884 VDD.n3883 9.3005
R7100 VDD.n142 VDD.n141 9.3005
R7101 VDD.n3899 VDD.n3898 9.3005
R7102 VDD.n3900 VDD.n140 9.3005
R7103 VDD.n3902 VDD.n3901 9.3005
R7104 VDD.n3903 VDD.n139 9.3005
R7105 VDD.n3905 VDD.n3904 9.3005
R7106 VDD.n3906 VDD.n138 9.3005
R7107 VDD.n3908 VDD.n3907 9.3005
R7108 VDD.n3909 VDD.n136 9.3005
R7109 VDD.n3911 VDD.n3910 9.3005
R7110 VDD.n3912 VDD.n135 9.3005
R7111 VDD.n3914 VDD.n3913 9.3005
R7112 VDD.n3915 VDD.n133 9.3005
R7113 VDD.n3917 VDD.n3916 9.3005
R7114 VDD.n3918 VDD.n132 9.3005
R7115 VDD.n3920 VDD.n3919 9.3005
R7116 VDD.n3921 VDD.n130 9.3005
R7117 VDD.n3923 VDD.n3922 9.3005
R7118 VDD.n3924 VDD.n129 9.3005
R7119 VDD.n3926 VDD.n3925 9.3005
R7120 VDD.n3927 VDD.n127 9.3005
R7121 VDD.n3929 VDD.n3928 9.3005
R7122 VDD.n3930 VDD.n126 9.3005
R7123 VDD.n3932 VDD.n3931 9.3005
R7124 VDD.n3933 VDD.n124 9.3005
R7125 VDD.n3935 VDD.n3934 9.3005
R7126 VDD.n3936 VDD.n123 9.3005
R7127 VDD.n3938 VDD.n3937 9.3005
R7128 VDD.n3939 VDD.n121 9.3005
R7129 VDD.n3941 VDD.n3940 9.3005
R7130 VDD.n3942 VDD.n120 9.3005
R7131 VDD.n4266 VDD.n3943 9.3005
R7132 VDD.n4265 VDD.n3944 9.3005
R7133 VDD.n4264 VDD.n3945 9.3005
R7134 VDD.n4090 VDD.n3946 9.3005
R7135 VDD.n4092 VDD.n4091 9.3005
R7136 VDD.n4094 VDD.n4093 9.3005
R7137 VDD.n4095 VDD.n4089 9.3005
R7138 VDD.n4098 VDD.n4096 9.3005
R7139 VDD.n4099 VDD.n4088 9.3005
R7140 VDD.n4101 VDD.n4100 9.3005
R7141 VDD.n4102 VDD.n4087 9.3005
R7142 VDD.n4105 VDD.n4103 9.3005
R7143 VDD.n4106 VDD.n4086 9.3005
R7144 VDD.n4108 VDD.n4107 9.3005
R7145 VDD.n4109 VDD.n4085 9.3005
R7146 VDD.n4112 VDD.n4110 9.3005
R7147 VDD.n4113 VDD.n4084 9.3005
R7148 VDD.n4115 VDD.n4114 9.3005
R7149 VDD.n4116 VDD.n4083 9.3005
R7150 VDD.n4119 VDD.n4117 9.3005
R7151 VDD.n4120 VDD.n4082 9.3005
R7152 VDD.n4122 VDD.n4121 9.3005
R7153 VDD.n285 VDD.n284 9.3005
R7154 VDD.n4219 VDD.n4218 9.3005
R7155 VDD.n4217 VDD.n4029 9.3005
R7156 VDD.n4216 VDD.n4215 9.3005
R7157 VDD.n4212 VDD.n4030 9.3005
R7158 VDD.n4209 VDD.n4031 9.3005
R7159 VDD.n4208 VDD.n4032 9.3005
R7160 VDD.n4205 VDD.n4033 9.3005
R7161 VDD.n4204 VDD.n4034 9.3005
R7162 VDD.n4201 VDD.n4035 9.3005
R7163 VDD.n4200 VDD.n4036 9.3005
R7164 VDD.n4197 VDD.n4037 9.3005
R7165 VDD.n4196 VDD.n4038 9.3005
R7166 VDD.n4193 VDD.n4039 9.3005
R7167 VDD.n4192 VDD.n4191 9.3005
R7168 VDD.n4190 VDD.n4040 9.3005
R7169 VDD.n4189 VDD.n4188 9.3005
R7170 VDD.n4185 VDD.n4045 9.3005
R7171 VDD.n4184 VDD.n4046 9.3005
R7172 VDD.n4181 VDD.n4047 9.3005
R7173 VDD.n4180 VDD.n4048 9.3005
R7174 VDD.n4177 VDD.n4049 9.3005
R7175 VDD.n4176 VDD.n4050 9.3005
R7176 VDD.n4173 VDD.n4051 9.3005
R7177 VDD.n4172 VDD.n4052 9.3005
R7178 VDD.n4169 VDD.n4053 9.3005
R7179 VDD.n4168 VDD.n4054 9.3005
R7180 VDD.n4165 VDD.n4055 9.3005
R7181 VDD.n4164 VDD.n4056 9.3005
R7182 VDD.n4161 VDD.n4057 9.3005
R7183 VDD.n4160 VDD.n4058 9.3005
R7184 VDD.n4157 VDD.n4062 9.3005
R7185 VDD.n4156 VDD.n4063 9.3005
R7186 VDD.n4153 VDD.n4064 9.3005
R7187 VDD.n4152 VDD.n4065 9.3005
R7188 VDD.n4149 VDD.n4066 9.3005
R7189 VDD.n4148 VDD.n4067 9.3005
R7190 VDD.n4145 VDD.n4068 9.3005
R7191 VDD.n4144 VDD.n4069 9.3005
R7192 VDD.n4141 VDD.n4070 9.3005
R7193 VDD.n4140 VDD.n4071 9.3005
R7194 VDD.n4137 VDD.n4072 9.3005
R7195 VDD.n4136 VDD.n4073 9.3005
R7196 VDD.n4133 VDD.n4074 9.3005
R7197 VDD.n4132 VDD.n4075 9.3005
R7198 VDD.n4129 VDD.n4076 9.3005
R7199 VDD.n4128 VDD.n4077 9.3005
R7200 VDD.n4125 VDD.n4124 9.3005
R7201 VDD.n4123 VDD.n4079 9.3005
R7202 VDD.n4220 VDD.n4028 9.3005
R7203 VDD.n4327 VDD.n4326 9.3005
R7204 VDD.n4325 VDD.n34 9.3005
R7205 VDD.n45 VDD.n37 9.3005
R7206 VDD.n4319 VDD.n46 9.3005
R7207 VDD.n4318 VDD.n47 9.3005
R7208 VDD.n4317 VDD.n48 9.3005
R7209 VDD.n56 VDD.n49 9.3005
R7210 VDD.n4311 VDD.n57 9.3005
R7211 VDD.n4310 VDD.n58 9.3005
R7212 VDD.n4309 VDD.n59 9.3005
R7213 VDD.n67 VDD.n60 9.3005
R7214 VDD.n4303 VDD.n68 9.3005
R7215 VDD.n4302 VDD.n69 9.3005
R7216 VDD.n4301 VDD.n70 9.3005
R7217 VDD.n78 VDD.n71 9.3005
R7218 VDD.n4295 VDD.n79 9.3005
R7219 VDD.n4294 VDD.n80 9.3005
R7220 VDD.n4293 VDD.n81 9.3005
R7221 VDD.n89 VDD.n82 9.3005
R7222 VDD.n4287 VDD.n90 9.3005
R7223 VDD.n4286 VDD.n91 9.3005
R7224 VDD.n4285 VDD.n92 9.3005
R7225 VDD.n100 VDD.n93 9.3005
R7226 VDD.n4279 VDD.n101 9.3005
R7227 VDD.n4278 VDD.n102 9.3005
R7228 VDD.n4277 VDD.n103 9.3005
R7229 VDD.n111 VDD.n104 9.3005
R7230 VDD.n4271 VDD.n112 9.3005
R7231 VDD.n4270 VDD.n113 9.3005
R7232 VDD.n4269 VDD.n114 9.3005
R7233 VDD.n3950 VDD.n115 9.3005
R7234 VDD.n4260 VDD.n3951 9.3005
R7235 VDD.n4259 VDD.n3952 9.3005
R7236 VDD.n4258 VDD.n3953 9.3005
R7237 VDD.n3961 VDD.n3954 9.3005
R7238 VDD.n4252 VDD.n3962 9.3005
R7239 VDD.n4251 VDD.n3963 9.3005
R7240 VDD.n4250 VDD.n3964 9.3005
R7241 VDD.n3972 VDD.n3965 9.3005
R7242 VDD.n4244 VDD.n3973 9.3005
R7243 VDD.n4243 VDD.n3974 9.3005
R7244 VDD.n4242 VDD.n3975 9.3005
R7245 VDD.n3982 VDD.n3976 9.3005
R7246 VDD.n4236 VDD.n3983 9.3005
R7247 VDD.n4235 VDD.n3984 9.3005
R7248 VDD.n4234 VDD.n3985 9.3005
R7249 VDD.n3994 VDD.n3986 9.3005
R7250 VDD.n4228 VDD.n3995 9.3005
R7251 VDD.n4227 VDD.n3996 9.3005
R7252 VDD.n4226 VDD.n3997 9.3005
R7253 VDD.n4027 VDD.n3998 9.3005
R7254 VDD.n3696 VDD.n3695 9.3005
R7255 VDD.n279 VDD.n278 9.3005
R7256 VDD.n3709 VDD.n3708 9.3005
R7257 VDD.n3710 VDD.n277 9.3005
R7258 VDD.n3712 VDD.n3711 9.3005
R7259 VDD.n267 VDD.n266 9.3005
R7260 VDD.n3725 VDD.n3724 9.3005
R7261 VDD.n3726 VDD.n265 9.3005
R7262 VDD.n3728 VDD.n3727 9.3005
R7263 VDD.n255 VDD.n254 9.3005
R7264 VDD.n3741 VDD.n3740 9.3005
R7265 VDD.n3742 VDD.n253 9.3005
R7266 VDD.n3744 VDD.n3743 9.3005
R7267 VDD.n243 VDD.n242 9.3005
R7268 VDD.n3757 VDD.n3756 9.3005
R7269 VDD.n3758 VDD.n241 9.3005
R7270 VDD.n3760 VDD.n3759 9.3005
R7271 VDD.n231 VDD.n230 9.3005
R7272 VDD.n3773 VDD.n3772 9.3005
R7273 VDD.n3774 VDD.n229 9.3005
R7274 VDD.n3776 VDD.n3775 9.3005
R7275 VDD.n219 VDD.n218 9.3005
R7276 VDD.n3788 VDD.n3787 9.3005
R7277 VDD.n3789 VDD.n217 9.3005
R7278 VDD.n3791 VDD.n3790 9.3005
R7279 VDD.n207 VDD.n206 9.3005
R7280 VDD.n3804 VDD.n3803 9.3005
R7281 VDD.n3805 VDD.n205 9.3005
R7282 VDD.n3807 VDD.n3806 9.3005
R7283 VDD.n195 VDD.n194 9.3005
R7284 VDD.n3821 VDD.n3820 9.3005
R7285 VDD.n3822 VDD.n193 9.3005
R7286 VDD.n3824 VDD.n3823 9.3005
R7287 VDD.n184 VDD.n183 9.3005
R7288 VDD.n3837 VDD.n3836 9.3005
R7289 VDD.n3838 VDD.n182 9.3005
R7290 VDD.n3840 VDD.n3839 9.3005
R7291 VDD.n172 VDD.n171 9.3005
R7292 VDD.n3853 VDD.n3852 9.3005
R7293 VDD.n3854 VDD.n170 9.3005
R7294 VDD.n3856 VDD.n3855 9.3005
R7295 VDD.n160 VDD.n159 9.3005
R7296 VDD.n3872 VDD.n3871 9.3005
R7297 VDD.n3873 VDD.n158 9.3005
R7298 VDD.n3875 VDD.n3874 9.3005
R7299 VDD.n149 VDD.n148 9.3005
R7300 VDD.n3890 VDD.n3889 9.3005
R7301 VDD.n3891 VDD.n147 9.3005
R7302 VDD.n3893 VDD.n3892 9.3005
R7303 VDD.n35 VDD.n33 9.3005
R7304 VDD.n3694 VDD.n289 9.3005
R7305 VDD.n3589 VDD.n3566 9.3005
R7306 VDD.n3586 VDD.n3585 9.3005
R7307 VDD.n3584 VDD.n3567 9.3005
R7308 VDD.n3583 VDD.n3582 9.3005
R7309 VDD.n3579 VDD.n3568 9.3005
R7310 VDD.n3576 VDD.n3575 9.3005
R7311 VDD.n3574 VDD.n3569 9.3005
R7312 VDD.n3573 VDD.n3572 9.3005
R7313 VDD.n295 VDD.n293 9.3005
R7314 VDD.n3692 VDD.n3691 9.3005
R7315 VDD.n3595 VDD.n3594 9.3005
R7316 VDD.n3638 VDD.n3637 9.3005
R7317 VDD.n3631 VDD.n3558 9.3005
R7318 VDD.n3628 VDD.n3627 9.3005
R7319 VDD.n3626 VDD.n3559 9.3005
R7320 VDD.n3625 VDD.n3624 9.3005
R7321 VDD.n3621 VDD.n3560 9.3005
R7322 VDD.n3618 VDD.n3617 9.3005
R7323 VDD.n3616 VDD.n3561 9.3005
R7324 VDD.n3615 VDD.n3614 9.3005
R7325 VDD.n3611 VDD.n3562 9.3005
R7326 VDD.n3608 VDD.n3607 9.3005
R7327 VDD.n3606 VDD.n3563 9.3005
R7328 VDD.n3605 VDD.n3604 9.3005
R7329 VDD.n3601 VDD.n3564 9.3005
R7330 VDD.n3598 VDD.n3597 9.3005
R7331 VDD.n3596 VDD.n3565 9.3005
R7332 VDD.n3671 VDD.n3670 9.3005
R7333 VDD.n3669 VDD.n3551 9.3005
R7334 VDD.n3668 VDD.n3667 9.3005
R7335 VDD.n3664 VDD.n3552 9.3005
R7336 VDD.n3661 VDD.n3660 9.3005
R7337 VDD.n3659 VDD.n3553 9.3005
R7338 VDD.n3658 VDD.n3657 9.3005
R7339 VDD.n3654 VDD.n3554 9.3005
R7340 VDD.n3651 VDD.n3650 9.3005
R7341 VDD.n3649 VDD.n3555 9.3005
R7342 VDD.n3648 VDD.n3647 9.3005
R7343 VDD.n3644 VDD.n3556 9.3005
R7344 VDD.n3641 VDD.n3640 9.3005
R7345 VDD.n3639 VDD.n3557 9.3005
R7346 VDD.n1680 VDD.n1679 9.3005
R7347 VDD.n1488 VDD.n1487 9.3005
R7348 VDD.n1693 VDD.n1692 9.3005
R7349 VDD.n1694 VDD.n1486 9.3005
R7350 VDD.n1696 VDD.n1695 9.3005
R7351 VDD.n1477 VDD.n1476 9.3005
R7352 VDD.n1710 VDD.n1709 9.3005
R7353 VDD.n1711 VDD.n1475 9.3005
R7354 VDD.n1713 VDD.n1712 9.3005
R7355 VDD.n1465 VDD.n1464 9.3005
R7356 VDD.n1726 VDD.n1725 9.3005
R7357 VDD.n1727 VDD.n1463 9.3005
R7358 VDD.n1729 VDD.n1728 9.3005
R7359 VDD.n1453 VDD.n1452 9.3005
R7360 VDD.n1742 VDD.n1741 9.3005
R7361 VDD.n1743 VDD.n1451 9.3005
R7362 VDD.n1745 VDD.n1744 9.3005
R7363 VDD.n1441 VDD.n1440 9.3005
R7364 VDD.n1758 VDD.n1757 9.3005
R7365 VDD.n1759 VDD.n1439 9.3005
R7366 VDD.n1761 VDD.n1760 9.3005
R7367 VDD.n1429 VDD.n1428 9.3005
R7368 VDD.n1773 VDD.n1772 9.3005
R7369 VDD.n1774 VDD.n1427 9.3005
R7370 VDD.n1776 VDD.n1775 9.3005
R7371 VDD.n1417 VDD.n1416 9.3005
R7372 VDD.n1789 VDD.n1788 9.3005
R7373 VDD.n1790 VDD.n1415 9.3005
R7374 VDD.n1792 VDD.n1791 9.3005
R7375 VDD.n1404 VDD.n1403 9.3005
R7376 VDD.n1805 VDD.n1804 9.3005
R7377 VDD.n1806 VDD.n1402 9.3005
R7378 VDD.n1808 VDD.n1807 9.3005
R7379 VDD.n1393 VDD.n1392 9.3005
R7380 VDD.n1821 VDD.n1820 9.3005
R7381 VDD.n1822 VDD.n1391 9.3005
R7382 VDD.n1824 VDD.n1823 9.3005
R7383 VDD.n1381 VDD.n1380 9.3005
R7384 VDD.n1837 VDD.n1836 9.3005
R7385 VDD.n1838 VDD.n1379 9.3005
R7386 VDD.n1840 VDD.n1839 9.3005
R7387 VDD.n1368 VDD.n1367 9.3005
R7388 VDD.n1853 VDD.n1852 9.3005
R7389 VDD.n1854 VDD.n1366 9.3005
R7390 VDD.n1856 VDD.n1855 9.3005
R7391 VDD.n1357 VDD.n1356 9.3005
R7392 VDD.n1869 VDD.n1868 9.3005
R7393 VDD.n1870 VDD.n1355 9.3005
R7394 VDD.n1872 VDD.n1871 9.3005
R7395 VDD.n1345 VDD.n1344 9.3005
R7396 VDD.n1904 VDD.n1903 9.3005
R7397 VDD.n1905 VDD.n1343 9.3005
R7398 VDD.n1907 VDD.n1906 9.3005
R7399 VDD.n1332 VDD.n1331 9.3005
R7400 VDD.n1920 VDD.n1919 9.3005
R7401 VDD.n1921 VDD.n1330 9.3005
R7402 VDD.n1923 VDD.n1922 9.3005
R7403 VDD.n1321 VDD.n1320 9.3005
R7404 VDD.n1936 VDD.n1935 9.3005
R7405 VDD.n1937 VDD.n1319 9.3005
R7406 VDD.n1939 VDD.n1938 9.3005
R7407 VDD.n1309 VDD.n1308 9.3005
R7408 VDD.n1952 VDD.n1951 9.3005
R7409 VDD.n1953 VDD.n1307 9.3005
R7410 VDD.n1955 VDD.n1954 9.3005
R7411 VDD.n1296 VDD.n1295 9.3005
R7412 VDD.n1968 VDD.n1967 9.3005
R7413 VDD.n1969 VDD.n1294 9.3005
R7414 VDD.n1971 VDD.n1970 9.3005
R7415 VDD.n1285 VDD.n1284 9.3005
R7416 VDD.n1984 VDD.n1983 9.3005
R7417 VDD.n1985 VDD.n1283 9.3005
R7418 VDD.n1987 VDD.n1986 9.3005
R7419 VDD.n1273 VDD.n1272 9.3005
R7420 VDD.n2000 VDD.n1999 9.3005
R7421 VDD.n2001 VDD.n1271 9.3005
R7422 VDD.n2003 VDD.n2002 9.3005
R7423 VDD.n1261 VDD.n1260 9.3005
R7424 VDD.n2016 VDD.n2015 9.3005
R7425 VDD.n2017 VDD.n1259 9.3005
R7426 VDD.n2019 VDD.n2018 9.3005
R7427 VDD.n1250 VDD.n1249 9.3005
R7428 VDD.n2032 VDD.n2031 9.3005
R7429 VDD.n2033 VDD.n1248 9.3005
R7430 VDD.n2035 VDD.n2034 9.3005
R7431 VDD.n1238 VDD.n1237 9.3005
R7432 VDD.n2048 VDD.n2047 9.3005
R7433 VDD.n2049 VDD.n1236 9.3005
R7434 VDD.n2051 VDD.n2050 9.3005
R7435 VDD.n1226 VDD.n1225 9.3005
R7436 VDD.n2064 VDD.n2063 9.3005
R7437 VDD.n2065 VDD.n1224 9.3005
R7438 VDD.n2067 VDD.n2066 9.3005
R7439 VDD.n1215 VDD.n1214 9.3005
R7440 VDD.n2081 VDD.n2080 9.3005
R7441 VDD.n2082 VDD.n1212 9.3005
R7442 VDD.n2086 VDD.n2085 9.3005
R7443 VDD.n2084 VDD.n1213 9.3005
R7444 VDD.n2083 VDD.n1202 9.3005
R7445 VDD.n2099 VDD.n1201 9.3005
R7446 VDD.n2101 VDD.n2100 9.3005
R7447 VDD.n1678 VDD.n1498 9.3005
R7448 VDD.n1601 VDD.n1600 9.3005
R7449 VDD.n1603 VDD.n1602 9.3005
R7450 VDD.n1604 VDD.n1594 9.3005
R7451 VDD.n1606 VDD.n1605 9.3005
R7452 VDD.n1607 VDD.n1593 9.3005
R7453 VDD.n1609 VDD.n1608 9.3005
R7454 VDD.n1610 VDD.n1588 9.3005
R7455 VDD.n1612 VDD.n1611 9.3005
R7456 VDD.n1613 VDD.n1587 9.3005
R7457 VDD.n1615 VDD.n1614 9.3005
R7458 VDD.n1616 VDD.n1582 9.3005
R7459 VDD.n1618 VDD.n1617 9.3005
R7460 VDD.n1619 VDD.n1581 9.3005
R7461 VDD.n1621 VDD.n1620 9.3005
R7462 VDD.n1622 VDD.n1573 9.3005
R7463 VDD.n1624 VDD.n1623 9.3005
R7464 VDD.n1625 VDD.n1572 9.3005
R7465 VDD.n1627 VDD.n1626 9.3005
R7466 VDD.n1628 VDD.n1567 9.3005
R7467 VDD.n1630 VDD.n1629 9.3005
R7468 VDD.n1631 VDD.n1566 9.3005
R7469 VDD.n1633 VDD.n1632 9.3005
R7470 VDD.n1634 VDD.n1561 9.3005
R7471 VDD.n1636 VDD.n1635 9.3005
R7472 VDD.n1637 VDD.n1560 9.3005
R7473 VDD.n1639 VDD.n1638 9.3005
R7474 VDD.n1640 VDD.n1555 9.3005
R7475 VDD.n1642 VDD.n1641 9.3005
R7476 VDD.n1643 VDD.n1554 9.3005
R7477 VDD.n1645 VDD.n1644 9.3005
R7478 VDD.n1646 VDD.n1549 9.3005
R7479 VDD.n1648 VDD.n1647 9.3005
R7480 VDD.n1651 VDD.n1650 9.3005
R7481 VDD.n1652 VDD.n1541 9.3005
R7482 VDD.n1654 VDD.n1653 9.3005
R7483 VDD.n1655 VDD.n1540 9.3005
R7484 VDD.n1657 VDD.n1656 9.3005
R7485 VDD.n1658 VDD.n1535 9.3005
R7486 VDD.n1660 VDD.n1659 9.3005
R7487 VDD.n1661 VDD.n1534 9.3005
R7488 VDD.n1663 VDD.n1662 9.3005
R7489 VDD.n1664 VDD.n1530 9.3005
R7490 VDD.n1666 VDD.n1665 9.3005
R7491 VDD.n1667 VDD.n1529 9.3005
R7492 VDD.n1669 VDD.n1668 9.3005
R7493 VDD.n1670 VDD.n1528 9.3005
R7494 VDD.n1649 VDD.n1548 9.3005
R7495 VDD.n1502 VDD.n1499 9.3005
R7496 VDD.n1677 VDD.n1676 9.3005
R7497 VDD.n1685 VDD.n1684 9.3005
R7498 VDD.n1686 VDD.n1492 9.3005
R7499 VDD.n1688 VDD.n1687 9.3005
R7500 VDD.n1482 VDD.n1481 9.3005
R7501 VDD.n1702 VDD.n1701 9.3005
R7502 VDD.n1703 VDD.n1480 9.3005
R7503 VDD.n1705 VDD.n1704 9.3005
R7504 VDD.n1471 VDD.n1470 9.3005
R7505 VDD.n1718 VDD.n1717 9.3005
R7506 VDD.n1719 VDD.n1469 9.3005
R7507 VDD.n1721 VDD.n1720 9.3005
R7508 VDD.n1459 VDD.n1458 9.3005
R7509 VDD.n1734 VDD.n1733 9.3005
R7510 VDD.n1735 VDD.n1457 9.3005
R7511 VDD.n1737 VDD.n1736 9.3005
R7512 VDD.n1447 VDD.n1446 9.3005
R7513 VDD.n1750 VDD.n1749 9.3005
R7514 VDD.n1751 VDD.n1445 9.3005
R7515 VDD.n1753 VDD.n1752 9.3005
R7516 VDD.n1435 VDD.n1434 9.3005
R7517 VDD.n1765 VDD.n1764 9.3005
R7518 VDD.n1766 VDD.n1433 9.3005
R7519 VDD.n1768 VDD.n1767 9.3005
R7520 VDD.n1423 VDD.n1422 9.3005
R7521 VDD.n1781 VDD.n1780 9.3005
R7522 VDD.n1782 VDD.n1421 9.3005
R7523 VDD.n1784 VDD.n1783 9.3005
R7524 VDD.n1411 VDD.n1410 9.3005
R7525 VDD.n1797 VDD.n1796 9.3005
R7526 VDD.n1798 VDD.n1409 9.3005
R7527 VDD.n1800 VDD.n1799 9.3005
R7528 VDD.n1399 VDD.n1398 9.3005
R7529 VDD.n1813 VDD.n1812 9.3005
R7530 VDD.n1814 VDD.n1397 9.3005
R7531 VDD.n1816 VDD.n1815 9.3005
R7532 VDD.n1387 VDD.n1386 9.3005
R7533 VDD.n1829 VDD.n1828 9.3005
R7534 VDD.n1830 VDD.n1385 9.3005
R7535 VDD.n1832 VDD.n1831 9.3005
R7536 VDD.n1375 VDD.n1374 9.3005
R7537 VDD.n1845 VDD.n1844 9.3005
R7538 VDD.n1846 VDD.n1373 9.3005
R7539 VDD.n1848 VDD.n1847 9.3005
R7540 VDD.n1363 VDD.n1362 9.3005
R7541 VDD.n1861 VDD.n1860 9.3005
R7542 VDD.n1862 VDD.n1361 9.3005
R7543 VDD.n1864 VDD.n1863 9.3005
R7544 VDD.n1351 VDD.n1350 9.3005
R7545 VDD.n1877 VDD.n1876 9.3005
R7546 VDD.n1878 VDD.n1349 9.3005
R7547 VDD.n1494 VDD.n1493 9.3005
R7548 VDD.n1707 VDD.t14 9.14611
R7549 VDD.n2069 VDD.t3 9.14611
R7550 VDD.n3722 VDD.t10 9.14611
R7551 VDD.n4238 VDD.t22 9.14611
R7552 VDD.n1676 VDD.n1502 9.11565
R7553 VDD.n4125 VDD.n4079 9.11565
R7554 VDD.t123 VDD.n812 9.00321
R7555 VDD.n2556 VDD.t124 9.00321
R7556 VDD.n3295 VDD.t120 9.00321
R7557 VDD.n480 VDD.t127 9.00321
R7558 VDD.n1371 VDD.t97 8.57451
R7559 VDD.n1925 VDD.t110 8.57451
R7560 VDD.n903 VDD.t154 8.57451
R7561 VDD.t148 VDD.n388 8.57451
R7562 VDD.n3868 VDD.t103 8.57451
R7563 VDD.t83 VDD.n4314 8.57451
R7564 VDD.n2744 VDD.n659 8.42977
R7565 VDD.n2216 VDD.n1049 8.42977
R7566 VDD.n3134 VDD.n2812 8.42977
R7567 VDD.n3486 VDD.n358 8.42977
R7568 VDD.n3533 VDD.n330 8.42977
R7569 VDD.n2885 VDD.n2884 8.42977
R7570 VDD.n2678 VDD.n2677 8.42977
R7571 VDD.n1177 VDD.n1176 8.42977
R7572 VDD.n15 VDD.n14 8.34259
R7573 VDD.n4329 VDD.n4328 8.15
R7574 VDD.n1897 VDD.n1896 8.15
R7575 VDD.t41 VDD.n900 7.86001
R7576 VDD.n2646 VDD.t18 7.86001
R7577 VDD.n3205 VDD.t48 7.86001
R7578 VDD.n391 VDD.t58 7.86001
R7579 VDD.n2484 VDD.t143 7.57421
R7580 VDD.n748 VDD.t142 7.57421
R7581 VDD.t136 VDD.n544 7.57421
R7582 VDD.n3367 VDD.t139 7.57421
R7583 VDD.t152 VDD.n679 7.28841
R7584 VDD.n612 VDD.t134 7.28841
R7585 VDD.n2478 VDD.t137 7.14551
R7586 VDD.n3373 VDD.t118 7.14551
R7587 VDD.n808 VDD.t146 6.71681
R7588 VDD.t121 VDD.n484 6.71681
R7589 VDD.n2399 VDD.t140 6.43101
R7590 VDD.t130 VDD.n323 6.43101
R7591 VDD.n2616 VDD.t132 5.8594
R7592 VDD.n3235 VDD.t125 5.8594
R7593 VDD.n26 VDD.n20 5.8288
R7594 VDD.n1889 VDD.n1883 5.8288
R7595 VDD.n1576 VDD.n1572 5.81868
R7596 VDD.n2135 VDD.n1131 5.81868
R7597 VDD.n4160 VDD.n4061 5.81868
R7598 VDD.n3637 VDD.n3634 5.81868
R7599 VDD.n1858 VDD.t97 5.7165
R7600 VDD.n1335 VDD.t110 5.7165
R7601 VDD.n3877 VDD.t103 5.7165
R7602 VDD.n4315 VDD.t83 5.7165
R7603 VDD.n2574 VDD.t156 5.2878
R7604 VDD.n3277 VDD.t150 5.2878
R7605 VDD.n1698 VDD.t14 5.1449
R7606 VDD.n2078 VDD.t3 5.1449
R7607 VDD.n275 VDD.t10 5.1449
R7608 VDD.n3988 VDD.t22 5.1449
R7609 VDD.n4329 VDD.n32 5.06146
R7610 VDD.n1896 VDD.n1895 5.06146
R7611 VDD.n2104 VDD.n2103 4.74817
R7612 VDD.n2190 VDD.n1070 4.74817
R7613 VDD.n2191 VDD.n1069 4.74817
R7614 VDD.n2188 VDD.n1069 4.74817
R7615 VDD.n294 VDD.n292 4.74817
R7616 VDD.n3683 VDD.n292 4.74817
R7617 VDD.n3684 VDD.n291 4.74817
R7618 VDD.n3677 VDD.n3675 4.74817
R7619 VDD.n3675 VDD.n3674 4.74817
R7620 VDD.n2103 VDD.n1146 4.74817
R7621 VDD.n32 VDD.n31 4.63843
R7622 VDD.n26 VDD.n25 4.63843
R7623 VDD.n1895 VDD.n1894 4.63843
R7624 VDD.n1889 VDD.n1888 4.63843
R7625 VDD.t156 VDD.n758 4.4304
R7626 VDD.n534 VDD.t150 4.4304
R7627 VDD.n730 VDD.t132 3.8588
R7628 VDD.t125 VDD.n562 3.8588
R7629 VDD.n3679 VDD.n3548 3.12168
R7630 VDD.n2102 VDD.n1200 3.12168
R7631 VDD.n1200 VDD.n1199 3.05965
R7632 VDD.n3679 VDD.n3678 3.05965
R7633 VDD.n2538 VDD.t146 3.0014
R7634 VDD.n3313 VDD.t121 3.0014
R7635 VDD.n1810 VDD.t85 2.8585
R7636 VDD.n1299 VDD.t73 2.8585
R7637 VDD.n3826 VDD.t79 2.8585
R7638 VDD.n4291 VDD.t70 2.8585
R7639 VDD.n2357 VDD.t137 2.5727
R7640 VDD.n3026 VDD.t118 2.5727
R7641 VDD.n2654 VDD.t152 2.4298
R7642 VDD.n3199 VDD.t134 2.4298
R7643 VDD.n1896 VDD.n15 2.33734
R7644 VDD VDD.n4329 2.32951
R7645 VDD.n2199 VDD.n1070 2.27742
R7646 VDD.n2199 VDD.n1069 2.27742
R7647 VDD.n3693 VDD.n292 2.27742
R7648 VDD.n3693 VDD.n291 2.27742
R7649 VDD.n3675 VDD.n3548 2.27742
R7650 VDD.n2103 VDD.n2102 2.27742
R7651 VDD.n2741 VDD.n659 2.18587
R7652 VDD.n2219 VDD.n1049 2.18587
R7653 VDD.n3131 VDD.n2812 2.18587
R7654 VDD.n360 VDD.n358 2.18587
R7655 VDD.n332 VDD.n330 2.18587
R7656 VDD.n2886 VDD.n2885 2.18587
R7657 VDD.n2677 VDD.n2676 2.18587
R7658 VDD.n1176 VDD.n1175 2.18587
R7659 VDD.n2357 VDD.t143 2.144
R7660 VDD.n2598 VDD.t142 2.144
R7661 VDD.n3253 VDD.t136 2.144
R7662 VDD.n3026 VDD.t139 2.144
R7663 VDD.n2430 VDD.t41 1.8582
R7664 VDD.t18 VDD.n685 1.8582
R7665 VDD.n605 VDD.t48 1.8582
R7666 VDD.n3421 VDD.t58 1.8582
R7667 VDD.n30 VDD.n28 1.6959
R7668 VDD.n31 VDD.n30 1.6959
R7669 VDD.n24 VDD.n22 1.6959
R7670 VDD.n25 VDD.n24 1.6959
R7671 VDD.n19 VDD.n17 1.6959
R7672 VDD.n20 VDD.n19 1.6959
R7673 VDD.n1894 VDD.n1893 1.6959
R7674 VDD.n1893 VDD.n1891 1.6959
R7675 VDD.n1888 VDD.n1887 1.6959
R7676 VDD.n1887 VDD.n1885 1.6959
R7677 VDD.n1883 VDD.n1882 1.6959
R7678 VDD.n1882 VDD.n1880 1.6959
R7679 VDD.n4 VDD.n2 1.55438
R7680 VDD.n11 VDD.n9 1.55438
R7681 VDD.n6 VDD.n4 1.25625
R7682 VDD.n13 VDD.n11 1.25625
R7683 VDD.n32 VDD.n26 1.19087
R7684 VDD.n1895 VDD.n1889 1.19087
R7685 VDD.n2442 VDD.t154 1.1437
R7686 VDD.n3409 VDD.t148 1.1437
R7687 VDD.n14 VDD.n6 0.984695
R7688 VDD.n14 VDD.n13 0.984695
R7689 VDD.n1623 VDD.n1576 0.776258
R7690 VDD.n2132 VDD.n1131 0.776258
R7691 VDD.n4157 VDD.n4061 0.776258
R7692 VDD.n3634 VDD.n3557 0.776258
R7693 VDD.n2520 VDD.t123 0.715001
R7694 VDD.t124 VDD.n776 0.715001
R7695 VDD.n516 VDD.t120 0.715001
R7696 VDD.n3331 VDD.t127 0.715001
R7697 VDD.n4123 VDD.n4122 0.477634
R7698 VDD.n4028 VDD.n4027 0.477634
R7699 VDD.n1678 VDD.n1677 0.477634
R7700 VDD.n1528 VDD.n1493 0.477634
R7701 VDD.n2199 VDD.n2198 0.416658
R7702 VDD.n3548 VDD.n284 0.416658
R7703 VDD.n3694 VDD.n3693 0.416658
R7704 VDD.n2102 VDD.n2101 0.416658
R7705 VDD.n1101 VDD.n1068 0.152939
R7706 VDD.n1102 VDD.n1101 0.152939
R7707 VDD.n1103 VDD.n1102 0.152939
R7708 VDD.n1104 VDD.n1103 0.152939
R7709 VDD.n1105 VDD.n1104 0.152939
R7710 VDD.n1106 VDD.n1105 0.152939
R7711 VDD.n1107 VDD.n1106 0.152939
R7712 VDD.n1108 VDD.n1107 0.152939
R7713 VDD.n1109 VDD.n1108 0.152939
R7714 VDD.n2166 VDD.n1109 0.152939
R7715 VDD.n2166 VDD.n2165 0.152939
R7716 VDD.n2165 VDD.n2164 0.152939
R7717 VDD.n2164 VDD.n1115 0.152939
R7718 VDD.n1116 VDD.n1115 0.152939
R7719 VDD.n1117 VDD.n1116 0.152939
R7720 VDD.n1118 VDD.n1117 0.152939
R7721 VDD.n1119 VDD.n1118 0.152939
R7722 VDD.n1120 VDD.n1119 0.152939
R7723 VDD.n1121 VDD.n1120 0.152939
R7724 VDD.n1122 VDD.n1121 0.152939
R7725 VDD.n1123 VDD.n1122 0.152939
R7726 VDD.n1124 VDD.n1123 0.152939
R7727 VDD.n1125 VDD.n1124 0.152939
R7728 VDD.n1126 VDD.n1125 0.152939
R7729 VDD.n1127 VDD.n1126 0.152939
R7730 VDD.n1128 VDD.n1127 0.152939
R7731 VDD.n1132 VDD.n1128 0.152939
R7732 VDD.n1133 VDD.n1132 0.152939
R7733 VDD.n1134 VDD.n1133 0.152939
R7734 VDD.n1135 VDD.n1134 0.152939
R7735 VDD.n1136 VDD.n1135 0.152939
R7736 VDD.n1137 VDD.n1136 0.152939
R7737 VDD.n1138 VDD.n1137 0.152939
R7738 VDD.n1139 VDD.n1138 0.152939
R7739 VDD.n1140 VDD.n1139 0.152939
R7740 VDD.n1141 VDD.n1140 0.152939
R7741 VDD.n1142 VDD.n1141 0.152939
R7742 VDD.n1143 VDD.n1142 0.152939
R7743 VDD.n1144 VDD.n1143 0.152939
R7744 VDD.n1145 VDD.n1144 0.152939
R7745 VDD.n1898 VDD.n1338 0.152939
R7746 VDD.n1912 VDD.n1338 0.152939
R7747 VDD.n1913 VDD.n1912 0.152939
R7748 VDD.n1914 VDD.n1913 0.152939
R7749 VDD.n1914 VDD.n1326 0.152939
R7750 VDD.n1928 VDD.n1326 0.152939
R7751 VDD.n1929 VDD.n1928 0.152939
R7752 VDD.n1930 VDD.n1929 0.152939
R7753 VDD.n1930 VDD.n1314 0.152939
R7754 VDD.n1944 VDD.n1314 0.152939
R7755 VDD.n1945 VDD.n1944 0.152939
R7756 VDD.n1946 VDD.n1945 0.152939
R7757 VDD.n1946 VDD.n1302 0.152939
R7758 VDD.n1960 VDD.n1302 0.152939
R7759 VDD.n1961 VDD.n1960 0.152939
R7760 VDD.n1962 VDD.n1961 0.152939
R7761 VDD.n1962 VDD.n1290 0.152939
R7762 VDD.n1976 VDD.n1290 0.152939
R7763 VDD.n1977 VDD.n1976 0.152939
R7764 VDD.n1978 VDD.n1977 0.152939
R7765 VDD.n1978 VDD.n1278 0.152939
R7766 VDD.n1992 VDD.n1278 0.152939
R7767 VDD.n1993 VDD.n1992 0.152939
R7768 VDD.n1994 VDD.n1993 0.152939
R7769 VDD.n1994 VDD.n1266 0.152939
R7770 VDD.n2008 VDD.n1266 0.152939
R7771 VDD.n2009 VDD.n2008 0.152939
R7772 VDD.n2010 VDD.n2009 0.152939
R7773 VDD.n2010 VDD.n1255 0.152939
R7774 VDD.n2024 VDD.n1255 0.152939
R7775 VDD.n2025 VDD.n2024 0.152939
R7776 VDD.n2026 VDD.n2025 0.152939
R7777 VDD.n2026 VDD.n1243 0.152939
R7778 VDD.n2040 VDD.n1243 0.152939
R7779 VDD.n2041 VDD.n2040 0.152939
R7780 VDD.n2042 VDD.n2041 0.152939
R7781 VDD.n2042 VDD.n1231 0.152939
R7782 VDD.n2056 VDD.n1231 0.152939
R7783 VDD.n2057 VDD.n2056 0.152939
R7784 VDD.n2058 VDD.n2057 0.152939
R7785 VDD.n2058 VDD.n1219 0.152939
R7786 VDD.n2073 VDD.n1219 0.152939
R7787 VDD.n2074 VDD.n2073 0.152939
R7788 VDD.n2075 VDD.n2074 0.152939
R7789 VDD.n2075 VDD.n1207 0.152939
R7790 VDD.n2091 VDD.n1207 0.152939
R7791 VDD.n2092 VDD.n2091 0.152939
R7792 VDD.n2093 VDD.n2092 0.152939
R7793 VDD.n2093 VDD.n1071 0.152939
R7794 VDD.n2198 VDD.n1071 0.152939
R7795 VDD.n3701 VDD.n284 0.152939
R7796 VDD.n3702 VDD.n3701 0.152939
R7797 VDD.n3703 VDD.n3702 0.152939
R7798 VDD.n3703 VDD.n271 0.152939
R7799 VDD.n3717 VDD.n271 0.152939
R7800 VDD.n3718 VDD.n3717 0.152939
R7801 VDD.n3719 VDD.n3718 0.152939
R7802 VDD.n3719 VDD.n260 0.152939
R7803 VDD.n3733 VDD.n260 0.152939
R7804 VDD.n3734 VDD.n3733 0.152939
R7805 VDD.n3735 VDD.n3734 0.152939
R7806 VDD.n3735 VDD.n248 0.152939
R7807 VDD.n3749 VDD.n248 0.152939
R7808 VDD.n3750 VDD.n3749 0.152939
R7809 VDD.n3751 VDD.n3750 0.152939
R7810 VDD.n3751 VDD.n236 0.152939
R7811 VDD.n3765 VDD.n236 0.152939
R7812 VDD.n3766 VDD.n3765 0.152939
R7813 VDD.n3767 VDD.n3766 0.152939
R7814 VDD.n3767 VDD.n224 0.152939
R7815 VDD.n3780 VDD.n224 0.152939
R7816 VDD.n3781 VDD.n3780 0.152939
R7817 VDD.n3782 VDD.n3781 0.152939
R7818 VDD.n3782 VDD.n212 0.152939
R7819 VDD.n3796 VDD.n212 0.152939
R7820 VDD.n3797 VDD.n3796 0.152939
R7821 VDD.n3798 VDD.n3797 0.152939
R7822 VDD.n3798 VDD.n200 0.152939
R7823 VDD.n3812 VDD.n200 0.152939
R7824 VDD.n3813 VDD.n3812 0.152939
R7825 VDD.n3814 VDD.n3813 0.152939
R7826 VDD.n3814 VDD.n189 0.152939
R7827 VDD.n3829 VDD.n189 0.152939
R7828 VDD.n3830 VDD.n3829 0.152939
R7829 VDD.n3831 VDD.n3830 0.152939
R7830 VDD.n3831 VDD.n177 0.152939
R7831 VDD.n3845 VDD.n177 0.152939
R7832 VDD.n3846 VDD.n3845 0.152939
R7833 VDD.n3847 VDD.n3846 0.152939
R7834 VDD.n3847 VDD.n165 0.152939
R7835 VDD.n3861 VDD.n165 0.152939
R7836 VDD.n3862 VDD.n3861 0.152939
R7837 VDD.n3863 VDD.n3862 0.152939
R7838 VDD.n3864 VDD.n3863 0.152939
R7839 VDD.n3864 VDD.n154 0.152939
R7840 VDD.n3881 VDD.n154 0.152939
R7841 VDD.n3882 VDD.n3881 0.152939
R7842 VDD.n3883 VDD.n3882 0.152939
R7843 VDD.n3883 VDD.n141 0.152939
R7844 VDD.n3899 VDD.n141 0.152939
R7845 VDD.n3900 VDD.n3899 0.152939
R7846 VDD.n3901 VDD.n3900 0.152939
R7847 VDD.n3901 VDD.n139 0.152939
R7848 VDD.n3905 VDD.n139 0.152939
R7849 VDD.n3906 VDD.n3905 0.152939
R7850 VDD.n3907 VDD.n3906 0.152939
R7851 VDD.n3907 VDD.n136 0.152939
R7852 VDD.n3911 VDD.n136 0.152939
R7853 VDD.n3912 VDD.n3911 0.152939
R7854 VDD.n3913 VDD.n3912 0.152939
R7855 VDD.n3913 VDD.n133 0.152939
R7856 VDD.n3917 VDD.n133 0.152939
R7857 VDD.n3918 VDD.n3917 0.152939
R7858 VDD.n3919 VDD.n3918 0.152939
R7859 VDD.n3919 VDD.n130 0.152939
R7860 VDD.n3923 VDD.n130 0.152939
R7861 VDD.n3924 VDD.n3923 0.152939
R7862 VDD.n3925 VDD.n3924 0.152939
R7863 VDD.n3925 VDD.n127 0.152939
R7864 VDD.n3929 VDD.n127 0.152939
R7865 VDD.n3930 VDD.n3929 0.152939
R7866 VDD.n3931 VDD.n3930 0.152939
R7867 VDD.n3931 VDD.n124 0.152939
R7868 VDD.n3935 VDD.n124 0.152939
R7869 VDD.n3936 VDD.n3935 0.152939
R7870 VDD.n3937 VDD.n3936 0.152939
R7871 VDD.n3937 VDD.n121 0.152939
R7872 VDD.n3941 VDD.n121 0.152939
R7873 VDD.n3942 VDD.n3941 0.152939
R7874 VDD.n3943 VDD.n3942 0.152939
R7875 VDD.n3944 VDD.n3943 0.152939
R7876 VDD.n3945 VDD.n3944 0.152939
R7877 VDD.n4090 VDD.n3945 0.152939
R7878 VDD.n4091 VDD.n4090 0.152939
R7879 VDD.n4094 VDD.n4091 0.152939
R7880 VDD.n4095 VDD.n4094 0.152939
R7881 VDD.n4096 VDD.n4095 0.152939
R7882 VDD.n4096 VDD.n4088 0.152939
R7883 VDD.n4101 VDD.n4088 0.152939
R7884 VDD.n4102 VDD.n4101 0.152939
R7885 VDD.n4103 VDD.n4102 0.152939
R7886 VDD.n4103 VDD.n4086 0.152939
R7887 VDD.n4108 VDD.n4086 0.152939
R7888 VDD.n4109 VDD.n4108 0.152939
R7889 VDD.n4110 VDD.n4109 0.152939
R7890 VDD.n4110 VDD.n4084 0.152939
R7891 VDD.n4115 VDD.n4084 0.152939
R7892 VDD.n4116 VDD.n4115 0.152939
R7893 VDD.n4117 VDD.n4116 0.152939
R7894 VDD.n4117 VDD.n4082 0.152939
R7895 VDD.n4122 VDD.n4082 0.152939
R7896 VDD.n4218 VDD.n4028 0.152939
R7897 VDD.n4218 VDD.n4217 0.152939
R7898 VDD.n4217 VDD.n4216 0.152939
R7899 VDD.n4216 VDD.n4030 0.152939
R7900 VDD.n4031 VDD.n4030 0.152939
R7901 VDD.n4032 VDD.n4031 0.152939
R7902 VDD.n4033 VDD.n4032 0.152939
R7903 VDD.n4034 VDD.n4033 0.152939
R7904 VDD.n4035 VDD.n4034 0.152939
R7905 VDD.n4036 VDD.n4035 0.152939
R7906 VDD.n4037 VDD.n4036 0.152939
R7907 VDD.n4038 VDD.n4037 0.152939
R7908 VDD.n4039 VDD.n4038 0.152939
R7909 VDD.n4191 VDD.n4039 0.152939
R7910 VDD.n4191 VDD.n4190 0.152939
R7911 VDD.n4190 VDD.n4189 0.152939
R7912 VDD.n4189 VDD.n4045 0.152939
R7913 VDD.n4046 VDD.n4045 0.152939
R7914 VDD.n4047 VDD.n4046 0.152939
R7915 VDD.n4048 VDD.n4047 0.152939
R7916 VDD.n4049 VDD.n4048 0.152939
R7917 VDD.n4050 VDD.n4049 0.152939
R7918 VDD.n4051 VDD.n4050 0.152939
R7919 VDD.n4052 VDD.n4051 0.152939
R7920 VDD.n4053 VDD.n4052 0.152939
R7921 VDD.n4054 VDD.n4053 0.152939
R7922 VDD.n4055 VDD.n4054 0.152939
R7923 VDD.n4056 VDD.n4055 0.152939
R7924 VDD.n4057 VDD.n4056 0.152939
R7925 VDD.n4058 VDD.n4057 0.152939
R7926 VDD.n4062 VDD.n4058 0.152939
R7927 VDD.n4063 VDD.n4062 0.152939
R7928 VDD.n4064 VDD.n4063 0.152939
R7929 VDD.n4065 VDD.n4064 0.152939
R7930 VDD.n4066 VDD.n4065 0.152939
R7931 VDD.n4067 VDD.n4066 0.152939
R7932 VDD.n4068 VDD.n4067 0.152939
R7933 VDD.n4069 VDD.n4068 0.152939
R7934 VDD.n4070 VDD.n4069 0.152939
R7935 VDD.n4071 VDD.n4070 0.152939
R7936 VDD.n4072 VDD.n4071 0.152939
R7937 VDD.n4073 VDD.n4072 0.152939
R7938 VDD.n4074 VDD.n4073 0.152939
R7939 VDD.n4075 VDD.n4074 0.152939
R7940 VDD.n4076 VDD.n4075 0.152939
R7941 VDD.n4077 VDD.n4076 0.152939
R7942 VDD.n4124 VDD.n4077 0.152939
R7943 VDD.n4124 VDD.n4123 0.152939
R7944 VDD.n4327 VDD.n34 0.152939
R7945 VDD.n45 VDD.n34 0.152939
R7946 VDD.n46 VDD.n45 0.152939
R7947 VDD.n47 VDD.n46 0.152939
R7948 VDD.n48 VDD.n47 0.152939
R7949 VDD.n56 VDD.n48 0.152939
R7950 VDD.n57 VDD.n56 0.152939
R7951 VDD.n58 VDD.n57 0.152939
R7952 VDD.n59 VDD.n58 0.152939
R7953 VDD.n67 VDD.n59 0.152939
R7954 VDD.n68 VDD.n67 0.152939
R7955 VDD.n69 VDD.n68 0.152939
R7956 VDD.n70 VDD.n69 0.152939
R7957 VDD.n78 VDD.n70 0.152939
R7958 VDD.n79 VDD.n78 0.152939
R7959 VDD.n80 VDD.n79 0.152939
R7960 VDD.n81 VDD.n80 0.152939
R7961 VDD.n89 VDD.n81 0.152939
R7962 VDD.n90 VDD.n89 0.152939
R7963 VDD.n91 VDD.n90 0.152939
R7964 VDD.n92 VDD.n91 0.152939
R7965 VDD.n100 VDD.n92 0.152939
R7966 VDD.n101 VDD.n100 0.152939
R7967 VDD.n102 VDD.n101 0.152939
R7968 VDD.n103 VDD.n102 0.152939
R7969 VDD.n111 VDD.n103 0.152939
R7970 VDD.n112 VDD.n111 0.152939
R7971 VDD.n113 VDD.n112 0.152939
R7972 VDD.n114 VDD.n113 0.152939
R7973 VDD.n3950 VDD.n114 0.152939
R7974 VDD.n3951 VDD.n3950 0.152939
R7975 VDD.n3952 VDD.n3951 0.152939
R7976 VDD.n3953 VDD.n3952 0.152939
R7977 VDD.n3961 VDD.n3953 0.152939
R7978 VDD.n3962 VDD.n3961 0.152939
R7979 VDD.n3963 VDD.n3962 0.152939
R7980 VDD.n3964 VDD.n3963 0.152939
R7981 VDD.n3972 VDD.n3964 0.152939
R7982 VDD.n3973 VDD.n3972 0.152939
R7983 VDD.n3974 VDD.n3973 0.152939
R7984 VDD.n3975 VDD.n3974 0.152939
R7985 VDD.n3982 VDD.n3975 0.152939
R7986 VDD.n3983 VDD.n3982 0.152939
R7987 VDD.n3984 VDD.n3983 0.152939
R7988 VDD.n3985 VDD.n3984 0.152939
R7989 VDD.n3994 VDD.n3985 0.152939
R7990 VDD.n3995 VDD.n3994 0.152939
R7991 VDD.n3996 VDD.n3995 0.152939
R7992 VDD.n3997 VDD.n3996 0.152939
R7993 VDD.n4027 VDD.n3997 0.152939
R7994 VDD.n3695 VDD.n3694 0.152939
R7995 VDD.n3695 VDD.n278 0.152939
R7996 VDD.n3709 VDD.n278 0.152939
R7997 VDD.n3710 VDD.n3709 0.152939
R7998 VDD.n3711 VDD.n3710 0.152939
R7999 VDD.n3711 VDD.n266 0.152939
R8000 VDD.n3725 VDD.n266 0.152939
R8001 VDD.n3726 VDD.n3725 0.152939
R8002 VDD.n3727 VDD.n3726 0.152939
R8003 VDD.n3727 VDD.n254 0.152939
R8004 VDD.n3741 VDD.n254 0.152939
R8005 VDD.n3742 VDD.n3741 0.152939
R8006 VDD.n3743 VDD.n3742 0.152939
R8007 VDD.n3743 VDD.n242 0.152939
R8008 VDD.n3757 VDD.n242 0.152939
R8009 VDD.n3758 VDD.n3757 0.152939
R8010 VDD.n3759 VDD.n3758 0.152939
R8011 VDD.n3759 VDD.n230 0.152939
R8012 VDD.n3773 VDD.n230 0.152939
R8013 VDD.n3774 VDD.n3773 0.152939
R8014 VDD.n3775 VDD.n3774 0.152939
R8015 VDD.n3775 VDD.n218 0.152939
R8016 VDD.n3788 VDD.n218 0.152939
R8017 VDD.n3789 VDD.n3788 0.152939
R8018 VDD.n3790 VDD.n3789 0.152939
R8019 VDD.n3790 VDD.n206 0.152939
R8020 VDD.n3804 VDD.n206 0.152939
R8021 VDD.n3805 VDD.n3804 0.152939
R8022 VDD.n3806 VDD.n3805 0.152939
R8023 VDD.n3806 VDD.n194 0.152939
R8024 VDD.n3821 VDD.n194 0.152939
R8025 VDD.n3822 VDD.n3821 0.152939
R8026 VDD.n3823 VDD.n3822 0.152939
R8027 VDD.n3823 VDD.n183 0.152939
R8028 VDD.n3837 VDD.n183 0.152939
R8029 VDD.n3838 VDD.n3837 0.152939
R8030 VDD.n3839 VDD.n3838 0.152939
R8031 VDD.n3839 VDD.n171 0.152939
R8032 VDD.n3853 VDD.n171 0.152939
R8033 VDD.n3854 VDD.n3853 0.152939
R8034 VDD.n3855 VDD.n3854 0.152939
R8035 VDD.n3855 VDD.n159 0.152939
R8036 VDD.n3872 VDD.n159 0.152939
R8037 VDD.n3873 VDD.n3872 0.152939
R8038 VDD.n3874 VDD.n3873 0.152939
R8039 VDD.n3874 VDD.n148 0.152939
R8040 VDD.n3890 VDD.n148 0.152939
R8041 VDD.n3891 VDD.n3890 0.152939
R8042 VDD.n3892 VDD.n3891 0.152939
R8043 VDD.n3892 VDD.n33 0.152939
R8044 VDD.n3692 VDD.n293 0.152939
R8045 VDD.n3573 VDD.n293 0.152939
R8046 VDD.n3574 VDD.n3573 0.152939
R8047 VDD.n3575 VDD.n3574 0.152939
R8048 VDD.n3575 VDD.n3568 0.152939
R8049 VDD.n3583 VDD.n3568 0.152939
R8050 VDD.n3584 VDD.n3583 0.152939
R8051 VDD.n3585 VDD.n3584 0.152939
R8052 VDD.n3585 VDD.n3566 0.152939
R8053 VDD.n3595 VDD.n3566 0.152939
R8054 VDD.n3596 VDD.n3595 0.152939
R8055 VDD.n3597 VDD.n3596 0.152939
R8056 VDD.n3597 VDD.n3564 0.152939
R8057 VDD.n3605 VDD.n3564 0.152939
R8058 VDD.n3606 VDD.n3605 0.152939
R8059 VDD.n3607 VDD.n3606 0.152939
R8060 VDD.n3607 VDD.n3562 0.152939
R8061 VDD.n3615 VDD.n3562 0.152939
R8062 VDD.n3616 VDD.n3615 0.152939
R8063 VDD.n3617 VDD.n3616 0.152939
R8064 VDD.n3617 VDD.n3560 0.152939
R8065 VDD.n3625 VDD.n3560 0.152939
R8066 VDD.n3626 VDD.n3625 0.152939
R8067 VDD.n3627 VDD.n3626 0.152939
R8068 VDD.n3627 VDD.n3558 0.152939
R8069 VDD.n3638 VDD.n3558 0.152939
R8070 VDD.n3639 VDD.n3638 0.152939
R8071 VDD.n3640 VDD.n3639 0.152939
R8072 VDD.n3640 VDD.n3556 0.152939
R8073 VDD.n3648 VDD.n3556 0.152939
R8074 VDD.n3649 VDD.n3648 0.152939
R8075 VDD.n3650 VDD.n3649 0.152939
R8076 VDD.n3650 VDD.n3554 0.152939
R8077 VDD.n3658 VDD.n3554 0.152939
R8078 VDD.n3659 VDD.n3658 0.152939
R8079 VDD.n3660 VDD.n3659 0.152939
R8080 VDD.n3660 VDD.n3552 0.152939
R8081 VDD.n3668 VDD.n3552 0.152939
R8082 VDD.n3669 VDD.n3668 0.152939
R8083 VDD.n3670 VDD.n3669 0.152939
R8084 VDD.n1679 VDD.n1678 0.152939
R8085 VDD.n1679 VDD.n1487 0.152939
R8086 VDD.n1693 VDD.n1487 0.152939
R8087 VDD.n1694 VDD.n1693 0.152939
R8088 VDD.n1695 VDD.n1694 0.152939
R8089 VDD.n1695 VDD.n1476 0.152939
R8090 VDD.n1710 VDD.n1476 0.152939
R8091 VDD.n1711 VDD.n1710 0.152939
R8092 VDD.n1712 VDD.n1711 0.152939
R8093 VDD.n1712 VDD.n1464 0.152939
R8094 VDD.n1726 VDD.n1464 0.152939
R8095 VDD.n1727 VDD.n1726 0.152939
R8096 VDD.n1728 VDD.n1727 0.152939
R8097 VDD.n1728 VDD.n1452 0.152939
R8098 VDD.n1742 VDD.n1452 0.152939
R8099 VDD.n1743 VDD.n1742 0.152939
R8100 VDD.n1744 VDD.n1743 0.152939
R8101 VDD.n1744 VDD.n1440 0.152939
R8102 VDD.n1758 VDD.n1440 0.152939
R8103 VDD.n1759 VDD.n1758 0.152939
R8104 VDD.n1760 VDD.n1759 0.152939
R8105 VDD.n1760 VDD.n1428 0.152939
R8106 VDD.n1773 VDD.n1428 0.152939
R8107 VDD.n1774 VDD.n1773 0.152939
R8108 VDD.n1775 VDD.n1774 0.152939
R8109 VDD.n1775 VDD.n1416 0.152939
R8110 VDD.n1789 VDD.n1416 0.152939
R8111 VDD.n1790 VDD.n1789 0.152939
R8112 VDD.n1791 VDD.n1790 0.152939
R8113 VDD.n1791 VDD.n1403 0.152939
R8114 VDD.n1805 VDD.n1403 0.152939
R8115 VDD.n1806 VDD.n1805 0.152939
R8116 VDD.n1807 VDD.n1806 0.152939
R8117 VDD.n1807 VDD.n1392 0.152939
R8118 VDD.n1821 VDD.n1392 0.152939
R8119 VDD.n1822 VDD.n1821 0.152939
R8120 VDD.n1823 VDD.n1822 0.152939
R8121 VDD.n1823 VDD.n1380 0.152939
R8122 VDD.n1837 VDD.n1380 0.152939
R8123 VDD.n1838 VDD.n1837 0.152939
R8124 VDD.n1839 VDD.n1838 0.152939
R8125 VDD.n1839 VDD.n1367 0.152939
R8126 VDD.n1853 VDD.n1367 0.152939
R8127 VDD.n1854 VDD.n1853 0.152939
R8128 VDD.n1855 VDD.n1854 0.152939
R8129 VDD.n1855 VDD.n1356 0.152939
R8130 VDD.n1869 VDD.n1356 0.152939
R8131 VDD.n1870 VDD.n1869 0.152939
R8132 VDD.n1871 VDD.n1870 0.152939
R8133 VDD.n1871 VDD.n1344 0.152939
R8134 VDD.n1904 VDD.n1344 0.152939
R8135 VDD.n1905 VDD.n1904 0.152939
R8136 VDD.n1906 VDD.n1905 0.152939
R8137 VDD.n1906 VDD.n1331 0.152939
R8138 VDD.n1920 VDD.n1331 0.152939
R8139 VDD.n1921 VDD.n1920 0.152939
R8140 VDD.n1922 VDD.n1921 0.152939
R8141 VDD.n1922 VDD.n1320 0.152939
R8142 VDD.n1936 VDD.n1320 0.152939
R8143 VDD.n1937 VDD.n1936 0.152939
R8144 VDD.n1938 VDD.n1937 0.152939
R8145 VDD.n1938 VDD.n1308 0.152939
R8146 VDD.n1952 VDD.n1308 0.152939
R8147 VDD.n1953 VDD.n1952 0.152939
R8148 VDD.n1954 VDD.n1953 0.152939
R8149 VDD.n1954 VDD.n1295 0.152939
R8150 VDD.n1968 VDD.n1295 0.152939
R8151 VDD.n1969 VDD.n1968 0.152939
R8152 VDD.n1970 VDD.n1969 0.152939
R8153 VDD.n1970 VDD.n1284 0.152939
R8154 VDD.n1984 VDD.n1284 0.152939
R8155 VDD.n1985 VDD.n1984 0.152939
R8156 VDD.n1986 VDD.n1985 0.152939
R8157 VDD.n1986 VDD.n1272 0.152939
R8158 VDD.n2000 VDD.n1272 0.152939
R8159 VDD.n2001 VDD.n2000 0.152939
R8160 VDD.n2002 VDD.n2001 0.152939
R8161 VDD.n2002 VDD.n1260 0.152939
R8162 VDD.n2016 VDD.n1260 0.152939
R8163 VDD.n2017 VDD.n2016 0.152939
R8164 VDD.n2018 VDD.n2017 0.152939
R8165 VDD.n2018 VDD.n1249 0.152939
R8166 VDD.n2032 VDD.n1249 0.152939
R8167 VDD.n2033 VDD.n2032 0.152939
R8168 VDD.n2034 VDD.n2033 0.152939
R8169 VDD.n2034 VDD.n1237 0.152939
R8170 VDD.n2048 VDD.n1237 0.152939
R8171 VDD.n2049 VDD.n2048 0.152939
R8172 VDD.n2050 VDD.n2049 0.152939
R8173 VDD.n2050 VDD.n1225 0.152939
R8174 VDD.n2064 VDD.n1225 0.152939
R8175 VDD.n2065 VDD.n2064 0.152939
R8176 VDD.n2066 VDD.n2065 0.152939
R8177 VDD.n2066 VDD.n1214 0.152939
R8178 VDD.n2081 VDD.n1214 0.152939
R8179 VDD.n2082 VDD.n2081 0.152939
R8180 VDD.n2085 VDD.n2082 0.152939
R8181 VDD.n2085 VDD.n2084 0.152939
R8182 VDD.n2084 VDD.n2083 0.152939
R8183 VDD.n2083 VDD.n1201 0.152939
R8184 VDD.n2101 VDD.n1201 0.152939
R8185 VDD.n1668 VDD.n1528 0.152939
R8186 VDD.n1668 VDD.n1667 0.152939
R8187 VDD.n1667 VDD.n1666 0.152939
R8188 VDD.n1666 VDD.n1530 0.152939
R8189 VDD.n1662 VDD.n1530 0.152939
R8190 VDD.n1662 VDD.n1661 0.152939
R8191 VDD.n1661 VDD.n1660 0.152939
R8192 VDD.n1660 VDD.n1535 0.152939
R8193 VDD.n1656 VDD.n1535 0.152939
R8194 VDD.n1656 VDD.n1655 0.152939
R8195 VDD.n1655 VDD.n1654 0.152939
R8196 VDD.n1654 VDD.n1541 0.152939
R8197 VDD.n1650 VDD.n1541 0.152939
R8198 VDD.n1650 VDD.n1649 0.152939
R8199 VDD.n1649 VDD.n1648 0.152939
R8200 VDD.n1648 VDD.n1549 0.152939
R8201 VDD.n1644 VDD.n1549 0.152939
R8202 VDD.n1644 VDD.n1643 0.152939
R8203 VDD.n1643 VDD.n1642 0.152939
R8204 VDD.n1642 VDD.n1555 0.152939
R8205 VDD.n1638 VDD.n1555 0.152939
R8206 VDD.n1638 VDD.n1637 0.152939
R8207 VDD.n1637 VDD.n1636 0.152939
R8208 VDD.n1636 VDD.n1561 0.152939
R8209 VDD.n1632 VDD.n1561 0.152939
R8210 VDD.n1632 VDD.n1631 0.152939
R8211 VDD.n1631 VDD.n1630 0.152939
R8212 VDD.n1630 VDD.n1567 0.152939
R8213 VDD.n1626 VDD.n1567 0.152939
R8214 VDD.n1626 VDD.n1625 0.152939
R8215 VDD.n1625 VDD.n1624 0.152939
R8216 VDD.n1624 VDD.n1573 0.152939
R8217 VDD.n1620 VDD.n1573 0.152939
R8218 VDD.n1620 VDD.n1619 0.152939
R8219 VDD.n1619 VDD.n1618 0.152939
R8220 VDD.n1618 VDD.n1582 0.152939
R8221 VDD.n1614 VDD.n1582 0.152939
R8222 VDD.n1614 VDD.n1613 0.152939
R8223 VDD.n1613 VDD.n1612 0.152939
R8224 VDD.n1612 VDD.n1588 0.152939
R8225 VDD.n1608 VDD.n1588 0.152939
R8226 VDD.n1608 VDD.n1607 0.152939
R8227 VDD.n1607 VDD.n1606 0.152939
R8228 VDD.n1606 VDD.n1594 0.152939
R8229 VDD.n1602 VDD.n1594 0.152939
R8230 VDD.n1602 VDD.n1601 0.152939
R8231 VDD.n1601 VDD.n1499 0.152939
R8232 VDD.n1677 VDD.n1499 0.152939
R8233 VDD.n1685 VDD.n1493 0.152939
R8234 VDD.n1686 VDD.n1685 0.152939
R8235 VDD.n1687 VDD.n1686 0.152939
R8236 VDD.n1687 VDD.n1481 0.152939
R8237 VDD.n1702 VDD.n1481 0.152939
R8238 VDD.n1703 VDD.n1702 0.152939
R8239 VDD.n1704 VDD.n1703 0.152939
R8240 VDD.n1704 VDD.n1470 0.152939
R8241 VDD.n1718 VDD.n1470 0.152939
R8242 VDD.n1719 VDD.n1718 0.152939
R8243 VDD.n1720 VDD.n1719 0.152939
R8244 VDD.n1720 VDD.n1458 0.152939
R8245 VDD.n1734 VDD.n1458 0.152939
R8246 VDD.n1735 VDD.n1734 0.152939
R8247 VDD.n1736 VDD.n1735 0.152939
R8248 VDD.n1736 VDD.n1446 0.152939
R8249 VDD.n1750 VDD.n1446 0.152939
R8250 VDD.n1751 VDD.n1750 0.152939
R8251 VDD.n1752 VDD.n1751 0.152939
R8252 VDD.n1752 VDD.n1434 0.152939
R8253 VDD.n1765 VDD.n1434 0.152939
R8254 VDD.n1766 VDD.n1765 0.152939
R8255 VDD.n1767 VDD.n1766 0.152939
R8256 VDD.n1767 VDD.n1422 0.152939
R8257 VDD.n1781 VDD.n1422 0.152939
R8258 VDD.n1782 VDD.n1781 0.152939
R8259 VDD.n1783 VDD.n1782 0.152939
R8260 VDD.n1783 VDD.n1410 0.152939
R8261 VDD.n1797 VDD.n1410 0.152939
R8262 VDD.n1798 VDD.n1797 0.152939
R8263 VDD.n1799 VDD.n1798 0.152939
R8264 VDD.n1799 VDD.n1398 0.152939
R8265 VDD.n1813 VDD.n1398 0.152939
R8266 VDD.n1814 VDD.n1813 0.152939
R8267 VDD.n1815 VDD.n1814 0.152939
R8268 VDD.n1815 VDD.n1386 0.152939
R8269 VDD.n1829 VDD.n1386 0.152939
R8270 VDD.n1830 VDD.n1829 0.152939
R8271 VDD.n1831 VDD.n1830 0.152939
R8272 VDD.n1831 VDD.n1374 0.152939
R8273 VDD.n1845 VDD.n1374 0.152939
R8274 VDD.n1846 VDD.n1845 0.152939
R8275 VDD.n1847 VDD.n1846 0.152939
R8276 VDD.n1847 VDD.n1362 0.152939
R8277 VDD.n1861 VDD.n1362 0.152939
R8278 VDD.n1862 VDD.n1861 0.152939
R8279 VDD.n1863 VDD.n1862 0.152939
R8280 VDD.n1863 VDD.n1350 0.152939
R8281 VDD.n1877 VDD.n1350 0.152939
R8282 VDD.n1878 VDD.n1877 0.152939
R8283 VDD.n1898 VDD.n1897 0.0695946
R8284 VDD.n4328 VDD.n4327 0.0695946
R8285 VDD.n4328 VDD.n33 0.0695946
R8286 VDD.n1897 VDD.n1878 0.0695946
R8287 VDD.n2199 VDD.n1068 0.0614756
R8288 VDD.n2102 VDD.n1145 0.0614756
R8289 VDD.n3693 VDD.n3692 0.0614756
R8290 VDD.n3670 VDD.n3548 0.0614756
R8291 VDD VDD.n15 0.00833333
R8292 CS_BIAS.n879 CS_BIAS.n878 161.3
R8293 CS_BIAS.n877 CS_BIAS.n737 161.3
R8294 CS_BIAS.n876 CS_BIAS.n875 161.3
R8295 CS_BIAS.n874 CS_BIAS.n738 161.3
R8296 CS_BIAS.n873 CS_BIAS.n872 161.3
R8297 CS_BIAS.n871 CS_BIAS.n739 161.3
R8298 CS_BIAS.n870 CS_BIAS.n869 161.3
R8299 CS_BIAS.n868 CS_BIAS.n740 161.3
R8300 CS_BIAS.n867 CS_BIAS.n866 161.3
R8301 CS_BIAS.n865 CS_BIAS.n741 161.3
R8302 CS_BIAS.n864 CS_BIAS.n863 161.3
R8303 CS_BIAS.n862 CS_BIAS.n861 161.3
R8304 CS_BIAS.n860 CS_BIAS.n743 161.3
R8305 CS_BIAS.n859 CS_BIAS.n858 161.3
R8306 CS_BIAS.n857 CS_BIAS.n744 161.3
R8307 CS_BIAS.n856 CS_BIAS.n855 161.3
R8308 CS_BIAS.n854 CS_BIAS.n745 161.3
R8309 CS_BIAS.n853 CS_BIAS.n852 161.3
R8310 CS_BIAS.n851 CS_BIAS.n746 161.3
R8311 CS_BIAS.n850 CS_BIAS.n849 161.3
R8312 CS_BIAS.n848 CS_BIAS.n747 161.3
R8313 CS_BIAS.n847 CS_BIAS.n846 161.3
R8314 CS_BIAS.n845 CS_BIAS.n844 161.3
R8315 CS_BIAS.n843 CS_BIAS.n749 161.3
R8316 CS_BIAS.n842 CS_BIAS.n841 161.3
R8317 CS_BIAS.n840 CS_BIAS.n750 161.3
R8318 CS_BIAS.n839 CS_BIAS.n838 161.3
R8319 CS_BIAS.n837 CS_BIAS.n751 161.3
R8320 CS_BIAS.n836 CS_BIAS.n835 161.3
R8321 CS_BIAS.n834 CS_BIAS.n752 161.3
R8322 CS_BIAS.n833 CS_BIAS.n832 161.3
R8323 CS_BIAS.n831 CS_BIAS.n753 161.3
R8324 CS_BIAS.n830 CS_BIAS.n829 161.3
R8325 CS_BIAS.n828 CS_BIAS.n754 161.3
R8326 CS_BIAS.n827 CS_BIAS.n826 161.3
R8327 CS_BIAS.n825 CS_BIAS.n755 161.3
R8328 CS_BIAS.n824 CS_BIAS.n823 161.3
R8329 CS_BIAS.n822 CS_BIAS.n757 161.3
R8330 CS_BIAS.n821 CS_BIAS.n820 161.3
R8331 CS_BIAS.n819 CS_BIAS.n758 161.3
R8332 CS_BIAS.n818 CS_BIAS.n817 161.3
R8333 CS_BIAS.n816 CS_BIAS.n759 161.3
R8334 CS_BIAS.n815 CS_BIAS.n814 161.3
R8335 CS_BIAS.n813 CS_BIAS.n760 161.3
R8336 CS_BIAS.n812 CS_BIAS.n811 161.3
R8337 CS_BIAS.n810 CS_BIAS.n809 161.3
R8338 CS_BIAS.n808 CS_BIAS.n762 161.3
R8339 CS_BIAS.n807 CS_BIAS.n806 161.3
R8340 CS_BIAS.n805 CS_BIAS.n763 161.3
R8341 CS_BIAS.n804 CS_BIAS.n803 161.3
R8342 CS_BIAS.n802 CS_BIAS.n764 161.3
R8343 CS_BIAS.n801 CS_BIAS.n800 161.3
R8344 CS_BIAS.n799 CS_BIAS.n765 161.3
R8345 CS_BIAS.n798 CS_BIAS.n797 161.3
R8346 CS_BIAS.n796 CS_BIAS.n766 161.3
R8347 CS_BIAS.n795 CS_BIAS.n794 161.3
R8348 CS_BIAS.n793 CS_BIAS.n767 161.3
R8349 CS_BIAS.n792 CS_BIAS.n791 161.3
R8350 CS_BIAS.n790 CS_BIAS.n768 161.3
R8351 CS_BIAS.n789 CS_BIAS.n788 161.3
R8352 CS_BIAS.n787 CS_BIAS.n770 161.3
R8353 CS_BIAS.n786 CS_BIAS.n785 161.3
R8354 CS_BIAS.n784 CS_BIAS.n771 161.3
R8355 CS_BIAS.n783 CS_BIAS.n782 161.3
R8356 CS_BIAS.n781 CS_BIAS.n772 161.3
R8357 CS_BIAS.n780 CS_BIAS.n779 161.3
R8358 CS_BIAS.n778 CS_BIAS.n773 161.3
R8359 CS_BIAS.n777 CS_BIAS.n776 161.3
R8360 CS_BIAS.n631 CS_BIAS.n630 161.3
R8361 CS_BIAS.n632 CS_BIAS.n627 161.3
R8362 CS_BIAS.n634 CS_BIAS.n633 161.3
R8363 CS_BIAS.n635 CS_BIAS.n626 161.3
R8364 CS_BIAS.n637 CS_BIAS.n636 161.3
R8365 CS_BIAS.n638 CS_BIAS.n625 161.3
R8366 CS_BIAS.n640 CS_BIAS.n639 161.3
R8367 CS_BIAS.n641 CS_BIAS.n624 161.3
R8368 CS_BIAS.n643 CS_BIAS.n642 161.3
R8369 CS_BIAS.n644 CS_BIAS.n622 161.3
R8370 CS_BIAS.n646 CS_BIAS.n645 161.3
R8371 CS_BIAS.n647 CS_BIAS.n621 161.3
R8372 CS_BIAS.n649 CS_BIAS.n648 161.3
R8373 CS_BIAS.n650 CS_BIAS.n620 161.3
R8374 CS_BIAS.n652 CS_BIAS.n651 161.3
R8375 CS_BIAS.n653 CS_BIAS.n619 161.3
R8376 CS_BIAS.n655 CS_BIAS.n654 161.3
R8377 CS_BIAS.n656 CS_BIAS.n618 161.3
R8378 CS_BIAS.n658 CS_BIAS.n657 161.3
R8379 CS_BIAS.n659 CS_BIAS.n617 161.3
R8380 CS_BIAS.n661 CS_BIAS.n660 161.3
R8381 CS_BIAS.n662 CS_BIAS.n616 161.3
R8382 CS_BIAS.n664 CS_BIAS.n663 161.3
R8383 CS_BIAS.n666 CS_BIAS.n665 161.3
R8384 CS_BIAS.n667 CS_BIAS.n614 161.3
R8385 CS_BIAS.n669 CS_BIAS.n668 161.3
R8386 CS_BIAS.n670 CS_BIAS.n613 161.3
R8387 CS_BIAS.n672 CS_BIAS.n671 161.3
R8388 CS_BIAS.n673 CS_BIAS.n612 161.3
R8389 CS_BIAS.n675 CS_BIAS.n674 161.3
R8390 CS_BIAS.n676 CS_BIAS.n611 161.3
R8391 CS_BIAS.n678 CS_BIAS.n677 161.3
R8392 CS_BIAS.n679 CS_BIAS.n609 161.3
R8393 CS_BIAS.n681 CS_BIAS.n680 161.3
R8394 CS_BIAS.n682 CS_BIAS.n608 161.3
R8395 CS_BIAS.n684 CS_BIAS.n683 161.3
R8396 CS_BIAS.n685 CS_BIAS.n607 161.3
R8397 CS_BIAS.n687 CS_BIAS.n686 161.3
R8398 CS_BIAS.n688 CS_BIAS.n606 161.3
R8399 CS_BIAS.n690 CS_BIAS.n689 161.3
R8400 CS_BIAS.n691 CS_BIAS.n605 161.3
R8401 CS_BIAS.n693 CS_BIAS.n692 161.3
R8402 CS_BIAS.n694 CS_BIAS.n604 161.3
R8403 CS_BIAS.n696 CS_BIAS.n695 161.3
R8404 CS_BIAS.n697 CS_BIAS.n603 161.3
R8405 CS_BIAS.n699 CS_BIAS.n698 161.3
R8406 CS_BIAS.n701 CS_BIAS.n700 161.3
R8407 CS_BIAS.n702 CS_BIAS.n601 161.3
R8408 CS_BIAS.n704 CS_BIAS.n703 161.3
R8409 CS_BIAS.n705 CS_BIAS.n600 161.3
R8410 CS_BIAS.n707 CS_BIAS.n706 161.3
R8411 CS_BIAS.n708 CS_BIAS.n599 161.3
R8412 CS_BIAS.n710 CS_BIAS.n709 161.3
R8413 CS_BIAS.n711 CS_BIAS.n598 161.3
R8414 CS_BIAS.n713 CS_BIAS.n712 161.3
R8415 CS_BIAS.n714 CS_BIAS.n597 161.3
R8416 CS_BIAS.n716 CS_BIAS.n715 161.3
R8417 CS_BIAS.n718 CS_BIAS.n717 161.3
R8418 CS_BIAS.n719 CS_BIAS.n595 161.3
R8419 CS_BIAS.n721 CS_BIAS.n720 161.3
R8420 CS_BIAS.n722 CS_BIAS.n594 161.3
R8421 CS_BIAS.n724 CS_BIAS.n723 161.3
R8422 CS_BIAS.n725 CS_BIAS.n593 161.3
R8423 CS_BIAS.n727 CS_BIAS.n726 161.3
R8424 CS_BIAS.n728 CS_BIAS.n592 161.3
R8425 CS_BIAS.n730 CS_BIAS.n729 161.3
R8426 CS_BIAS.n731 CS_BIAS.n591 161.3
R8427 CS_BIAS.n733 CS_BIAS.n732 161.3
R8428 CS_BIAS.n485 CS_BIAS.n484 161.3
R8429 CS_BIAS.n486 CS_BIAS.n481 161.3
R8430 CS_BIAS.n488 CS_BIAS.n487 161.3
R8431 CS_BIAS.n489 CS_BIAS.n480 161.3
R8432 CS_BIAS.n491 CS_BIAS.n490 161.3
R8433 CS_BIAS.n492 CS_BIAS.n479 161.3
R8434 CS_BIAS.n494 CS_BIAS.n493 161.3
R8435 CS_BIAS.n495 CS_BIAS.n478 161.3
R8436 CS_BIAS.n497 CS_BIAS.n496 161.3
R8437 CS_BIAS.n498 CS_BIAS.n476 161.3
R8438 CS_BIAS.n500 CS_BIAS.n499 161.3
R8439 CS_BIAS.n501 CS_BIAS.n475 161.3
R8440 CS_BIAS.n503 CS_BIAS.n502 161.3
R8441 CS_BIAS.n504 CS_BIAS.n474 161.3
R8442 CS_BIAS.n506 CS_BIAS.n505 161.3
R8443 CS_BIAS.n507 CS_BIAS.n473 161.3
R8444 CS_BIAS.n509 CS_BIAS.n508 161.3
R8445 CS_BIAS.n510 CS_BIAS.n472 161.3
R8446 CS_BIAS.n512 CS_BIAS.n511 161.3
R8447 CS_BIAS.n513 CS_BIAS.n471 161.3
R8448 CS_BIAS.n515 CS_BIAS.n514 161.3
R8449 CS_BIAS.n516 CS_BIAS.n470 161.3
R8450 CS_BIAS.n518 CS_BIAS.n517 161.3
R8451 CS_BIAS.n520 CS_BIAS.n519 161.3
R8452 CS_BIAS.n521 CS_BIAS.n468 161.3
R8453 CS_BIAS.n523 CS_BIAS.n522 161.3
R8454 CS_BIAS.n524 CS_BIAS.n467 161.3
R8455 CS_BIAS.n526 CS_BIAS.n525 161.3
R8456 CS_BIAS.n527 CS_BIAS.n466 161.3
R8457 CS_BIAS.n529 CS_BIAS.n528 161.3
R8458 CS_BIAS.n530 CS_BIAS.n465 161.3
R8459 CS_BIAS.n532 CS_BIAS.n531 161.3
R8460 CS_BIAS.n533 CS_BIAS.n463 161.3
R8461 CS_BIAS.n535 CS_BIAS.n534 161.3
R8462 CS_BIAS.n536 CS_BIAS.n462 161.3
R8463 CS_BIAS.n538 CS_BIAS.n537 161.3
R8464 CS_BIAS.n539 CS_BIAS.n461 161.3
R8465 CS_BIAS.n541 CS_BIAS.n540 161.3
R8466 CS_BIAS.n542 CS_BIAS.n460 161.3
R8467 CS_BIAS.n544 CS_BIAS.n543 161.3
R8468 CS_BIAS.n545 CS_BIAS.n459 161.3
R8469 CS_BIAS.n547 CS_BIAS.n546 161.3
R8470 CS_BIAS.n548 CS_BIAS.n458 161.3
R8471 CS_BIAS.n550 CS_BIAS.n549 161.3
R8472 CS_BIAS.n551 CS_BIAS.n457 161.3
R8473 CS_BIAS.n553 CS_BIAS.n552 161.3
R8474 CS_BIAS.n555 CS_BIAS.n554 161.3
R8475 CS_BIAS.n556 CS_BIAS.n455 161.3
R8476 CS_BIAS.n558 CS_BIAS.n557 161.3
R8477 CS_BIAS.n559 CS_BIAS.n454 161.3
R8478 CS_BIAS.n561 CS_BIAS.n560 161.3
R8479 CS_BIAS.n562 CS_BIAS.n453 161.3
R8480 CS_BIAS.n564 CS_BIAS.n563 161.3
R8481 CS_BIAS.n565 CS_BIAS.n452 161.3
R8482 CS_BIAS.n567 CS_BIAS.n566 161.3
R8483 CS_BIAS.n568 CS_BIAS.n451 161.3
R8484 CS_BIAS.n570 CS_BIAS.n569 161.3
R8485 CS_BIAS.n572 CS_BIAS.n571 161.3
R8486 CS_BIAS.n573 CS_BIAS.n449 161.3
R8487 CS_BIAS.n575 CS_BIAS.n574 161.3
R8488 CS_BIAS.n576 CS_BIAS.n448 161.3
R8489 CS_BIAS.n578 CS_BIAS.n577 161.3
R8490 CS_BIAS.n579 CS_BIAS.n447 161.3
R8491 CS_BIAS.n581 CS_BIAS.n580 161.3
R8492 CS_BIAS.n582 CS_BIAS.n446 161.3
R8493 CS_BIAS.n584 CS_BIAS.n583 161.3
R8494 CS_BIAS.n585 CS_BIAS.n445 161.3
R8495 CS_BIAS.n587 CS_BIAS.n586 161.3
R8496 CS_BIAS.n339 CS_BIAS.n338 161.3
R8497 CS_BIAS.n340 CS_BIAS.n335 161.3
R8498 CS_BIAS.n342 CS_BIAS.n341 161.3
R8499 CS_BIAS.n343 CS_BIAS.n334 161.3
R8500 CS_BIAS.n345 CS_BIAS.n344 161.3
R8501 CS_BIAS.n346 CS_BIAS.n333 161.3
R8502 CS_BIAS.n348 CS_BIAS.n347 161.3
R8503 CS_BIAS.n349 CS_BIAS.n332 161.3
R8504 CS_BIAS.n351 CS_BIAS.n350 161.3
R8505 CS_BIAS.n352 CS_BIAS.n330 161.3
R8506 CS_BIAS.n354 CS_BIAS.n353 161.3
R8507 CS_BIAS.n355 CS_BIAS.n329 161.3
R8508 CS_BIAS.n357 CS_BIAS.n356 161.3
R8509 CS_BIAS.n358 CS_BIAS.n328 161.3
R8510 CS_BIAS.n360 CS_BIAS.n359 161.3
R8511 CS_BIAS.n361 CS_BIAS.n327 161.3
R8512 CS_BIAS.n363 CS_BIAS.n362 161.3
R8513 CS_BIAS.n364 CS_BIAS.n326 161.3
R8514 CS_BIAS.n366 CS_BIAS.n365 161.3
R8515 CS_BIAS.n367 CS_BIAS.n325 161.3
R8516 CS_BIAS.n369 CS_BIAS.n368 161.3
R8517 CS_BIAS.n370 CS_BIAS.n324 161.3
R8518 CS_BIAS.n372 CS_BIAS.n371 161.3
R8519 CS_BIAS.n374 CS_BIAS.n373 161.3
R8520 CS_BIAS.n375 CS_BIAS.n322 161.3
R8521 CS_BIAS.n377 CS_BIAS.n376 161.3
R8522 CS_BIAS.n378 CS_BIAS.n321 161.3
R8523 CS_BIAS.n380 CS_BIAS.n379 161.3
R8524 CS_BIAS.n381 CS_BIAS.n320 161.3
R8525 CS_BIAS.n383 CS_BIAS.n382 161.3
R8526 CS_BIAS.n384 CS_BIAS.n319 161.3
R8527 CS_BIAS.n386 CS_BIAS.n385 161.3
R8528 CS_BIAS.n387 CS_BIAS.n317 161.3
R8529 CS_BIAS.n389 CS_BIAS.n388 161.3
R8530 CS_BIAS.n390 CS_BIAS.n316 161.3
R8531 CS_BIAS.n392 CS_BIAS.n391 161.3
R8532 CS_BIAS.n393 CS_BIAS.n315 161.3
R8533 CS_BIAS.n395 CS_BIAS.n394 161.3
R8534 CS_BIAS.n396 CS_BIAS.n314 161.3
R8535 CS_BIAS.n398 CS_BIAS.n397 161.3
R8536 CS_BIAS.n399 CS_BIAS.n313 161.3
R8537 CS_BIAS.n401 CS_BIAS.n400 161.3
R8538 CS_BIAS.n402 CS_BIAS.n312 161.3
R8539 CS_BIAS.n404 CS_BIAS.n403 161.3
R8540 CS_BIAS.n405 CS_BIAS.n311 161.3
R8541 CS_BIAS.n407 CS_BIAS.n406 161.3
R8542 CS_BIAS.n409 CS_BIAS.n408 161.3
R8543 CS_BIAS.n410 CS_BIAS.n309 161.3
R8544 CS_BIAS.n412 CS_BIAS.n411 161.3
R8545 CS_BIAS.n413 CS_BIAS.n308 161.3
R8546 CS_BIAS.n415 CS_BIAS.n414 161.3
R8547 CS_BIAS.n416 CS_BIAS.n307 161.3
R8548 CS_BIAS.n418 CS_BIAS.n417 161.3
R8549 CS_BIAS.n419 CS_BIAS.n306 161.3
R8550 CS_BIAS.n421 CS_BIAS.n420 161.3
R8551 CS_BIAS.n422 CS_BIAS.n305 161.3
R8552 CS_BIAS.n424 CS_BIAS.n423 161.3
R8553 CS_BIAS.n426 CS_BIAS.n425 161.3
R8554 CS_BIAS.n427 CS_BIAS.n303 161.3
R8555 CS_BIAS.n429 CS_BIAS.n428 161.3
R8556 CS_BIAS.n430 CS_BIAS.n302 161.3
R8557 CS_BIAS.n432 CS_BIAS.n431 161.3
R8558 CS_BIAS.n433 CS_BIAS.n301 161.3
R8559 CS_BIAS.n435 CS_BIAS.n434 161.3
R8560 CS_BIAS.n436 CS_BIAS.n300 161.3
R8561 CS_BIAS.n438 CS_BIAS.n437 161.3
R8562 CS_BIAS.n439 CS_BIAS.n299 161.3
R8563 CS_BIAS.n441 CS_BIAS.n440 161.3
R8564 CS_BIAS.n63 CS_BIAS.n62 161.3
R8565 CS_BIAS.n64 CS_BIAS.n59 161.3
R8566 CS_BIAS.n66 CS_BIAS.n65 161.3
R8567 CS_BIAS.n67 CS_BIAS.n58 161.3
R8568 CS_BIAS.n69 CS_BIAS.n68 161.3
R8569 CS_BIAS.n70 CS_BIAS.n57 161.3
R8570 CS_BIAS.n72 CS_BIAS.n71 161.3
R8571 CS_BIAS.n73 CS_BIAS.n56 161.3
R8572 CS_BIAS.n75 CS_BIAS.n74 161.3
R8573 CS_BIAS.n76 CS_BIAS.n54 161.3
R8574 CS_BIAS.n78 CS_BIAS.n77 161.3
R8575 CS_BIAS.n79 CS_BIAS.n53 161.3
R8576 CS_BIAS.n81 CS_BIAS.n80 161.3
R8577 CS_BIAS.n82 CS_BIAS.n52 161.3
R8578 CS_BIAS.n84 CS_BIAS.n83 161.3
R8579 CS_BIAS.n85 CS_BIAS.n51 161.3
R8580 CS_BIAS.n87 CS_BIAS.n86 161.3
R8581 CS_BIAS.n88 CS_BIAS.n50 161.3
R8582 CS_BIAS.n90 CS_BIAS.n89 161.3
R8583 CS_BIAS.n91 CS_BIAS.n49 161.3
R8584 CS_BIAS.n93 CS_BIAS.n92 161.3
R8585 CS_BIAS.n94 CS_BIAS.n48 161.3
R8586 CS_BIAS.n96 CS_BIAS.n95 161.3
R8587 CS_BIAS.n98 CS_BIAS.n97 161.3
R8588 CS_BIAS.n99 CS_BIAS.n46 161.3
R8589 CS_BIAS.n101 CS_BIAS.n100 161.3
R8590 CS_BIAS.n102 CS_BIAS.n45 161.3
R8591 CS_BIAS.n104 CS_BIAS.n103 161.3
R8592 CS_BIAS.n105 CS_BIAS.n44 161.3
R8593 CS_BIAS.n107 CS_BIAS.n106 161.3
R8594 CS_BIAS.n108 CS_BIAS.n43 161.3
R8595 CS_BIAS.n110 CS_BIAS.n109 161.3
R8596 CS_BIAS.n111 CS_BIAS.n41 161.3
R8597 CS_BIAS.n113 CS_BIAS.n112 161.3
R8598 CS_BIAS.n114 CS_BIAS.n40 161.3
R8599 CS_BIAS.n116 CS_BIAS.n115 161.3
R8600 CS_BIAS.n117 CS_BIAS.n39 161.3
R8601 CS_BIAS.n119 CS_BIAS.n118 161.3
R8602 CS_BIAS.n120 CS_BIAS.n38 161.3
R8603 CS_BIAS.n122 CS_BIAS.n121 161.3
R8604 CS_BIAS.n123 CS_BIAS.n37 161.3
R8605 CS_BIAS.n125 CS_BIAS.n124 161.3
R8606 CS_BIAS.n126 CS_BIAS.n36 161.3
R8607 CS_BIAS.n128 CS_BIAS.n127 161.3
R8608 CS_BIAS.n129 CS_BIAS.n35 161.3
R8609 CS_BIAS.n131 CS_BIAS.n130 161.3
R8610 CS_BIAS.n133 CS_BIAS.n132 161.3
R8611 CS_BIAS.n134 CS_BIAS.n33 161.3
R8612 CS_BIAS.n136 CS_BIAS.n135 161.3
R8613 CS_BIAS.n137 CS_BIAS.n32 161.3
R8614 CS_BIAS.n139 CS_BIAS.n138 161.3
R8615 CS_BIAS.n140 CS_BIAS.n31 161.3
R8616 CS_BIAS.n142 CS_BIAS.n141 161.3
R8617 CS_BIAS.n143 CS_BIAS.n30 161.3
R8618 CS_BIAS.n145 CS_BIAS.n144 161.3
R8619 CS_BIAS.n146 CS_BIAS.n29 161.3
R8620 CS_BIAS.n148 CS_BIAS.n147 161.3
R8621 CS_BIAS.n150 CS_BIAS.n149 161.3
R8622 CS_BIAS.n151 CS_BIAS.n27 161.3
R8623 CS_BIAS.n153 CS_BIAS.n152 161.3
R8624 CS_BIAS.n154 CS_BIAS.n26 161.3
R8625 CS_BIAS.n156 CS_BIAS.n155 161.3
R8626 CS_BIAS.n157 CS_BIAS.n25 161.3
R8627 CS_BIAS.n159 CS_BIAS.n158 161.3
R8628 CS_BIAS.n160 CS_BIAS.n24 161.3
R8629 CS_BIAS.n162 CS_BIAS.n161 161.3
R8630 CS_BIAS.n163 CS_BIAS.n23 161.3
R8631 CS_BIAS.n165 CS_BIAS.n164 161.3
R8632 CS_BIAS.n194 CS_BIAS.n193 161.3
R8633 CS_BIAS.n195 CS_BIAS.n190 161.3
R8634 CS_BIAS.n197 CS_BIAS.n196 161.3
R8635 CS_BIAS.n198 CS_BIAS.n189 161.3
R8636 CS_BIAS.n200 CS_BIAS.n199 161.3
R8637 CS_BIAS.n201 CS_BIAS.n188 161.3
R8638 CS_BIAS.n203 CS_BIAS.n202 161.3
R8639 CS_BIAS.n204 CS_BIAS.n187 161.3
R8640 CS_BIAS.n206 CS_BIAS.n205 161.3
R8641 CS_BIAS.n207 CS_BIAS.n185 161.3
R8642 CS_BIAS.n209 CS_BIAS.n208 161.3
R8643 CS_BIAS.n210 CS_BIAS.n184 161.3
R8644 CS_BIAS.n212 CS_BIAS.n211 161.3
R8645 CS_BIAS.n213 CS_BIAS.n183 161.3
R8646 CS_BIAS.n215 CS_BIAS.n214 161.3
R8647 CS_BIAS.n216 CS_BIAS.n182 161.3
R8648 CS_BIAS.n218 CS_BIAS.n217 161.3
R8649 CS_BIAS.n219 CS_BIAS.n181 161.3
R8650 CS_BIAS.n221 CS_BIAS.n220 161.3
R8651 CS_BIAS.n222 CS_BIAS.n180 161.3
R8652 CS_BIAS.n224 CS_BIAS.n223 161.3
R8653 CS_BIAS.n225 CS_BIAS.n179 161.3
R8654 CS_BIAS.n227 CS_BIAS.n226 161.3
R8655 CS_BIAS.n229 CS_BIAS.n228 161.3
R8656 CS_BIAS.n230 CS_BIAS.n177 161.3
R8657 CS_BIAS.n232 CS_BIAS.n231 161.3
R8658 CS_BIAS.n233 CS_BIAS.n176 161.3
R8659 CS_BIAS.n235 CS_BIAS.n234 161.3
R8660 CS_BIAS.n236 CS_BIAS.n175 161.3
R8661 CS_BIAS.n238 CS_BIAS.n237 161.3
R8662 CS_BIAS.n239 CS_BIAS.n21 161.3
R8663 CS_BIAS.n241 CS_BIAS.n240 161.3
R8664 CS_BIAS.n242 CS_BIAS.n19 161.3
R8665 CS_BIAS.n244 CS_BIAS.n243 161.3
R8666 CS_BIAS.n245 CS_BIAS.n18 161.3
R8667 CS_BIAS.n247 CS_BIAS.n246 161.3
R8668 CS_BIAS.n248 CS_BIAS.n17 161.3
R8669 CS_BIAS.n250 CS_BIAS.n249 161.3
R8670 CS_BIAS.n251 CS_BIAS.n16 161.3
R8671 CS_BIAS.n253 CS_BIAS.n252 161.3
R8672 CS_BIAS.n254 CS_BIAS.n15 161.3
R8673 CS_BIAS.n256 CS_BIAS.n255 161.3
R8674 CS_BIAS.n257 CS_BIAS.n14 161.3
R8675 CS_BIAS.n259 CS_BIAS.n258 161.3
R8676 CS_BIAS.n260 CS_BIAS.n13 161.3
R8677 CS_BIAS.n262 CS_BIAS.n261 161.3
R8678 CS_BIAS.n264 CS_BIAS.n263 161.3
R8679 CS_BIAS.n265 CS_BIAS.n11 161.3
R8680 CS_BIAS.n267 CS_BIAS.n266 161.3
R8681 CS_BIAS.n268 CS_BIAS.n10 161.3
R8682 CS_BIAS.n270 CS_BIAS.n269 161.3
R8683 CS_BIAS.n271 CS_BIAS.n9 161.3
R8684 CS_BIAS.n273 CS_BIAS.n272 161.3
R8685 CS_BIAS.n274 CS_BIAS.n8 161.3
R8686 CS_BIAS.n276 CS_BIAS.n275 161.3
R8687 CS_BIAS.n277 CS_BIAS.n7 161.3
R8688 CS_BIAS.n279 CS_BIAS.n278 161.3
R8689 CS_BIAS.n281 CS_BIAS.n280 161.3
R8690 CS_BIAS.n282 CS_BIAS.n5 161.3
R8691 CS_BIAS.n284 CS_BIAS.n283 161.3
R8692 CS_BIAS.n285 CS_BIAS.n4 161.3
R8693 CS_BIAS.n287 CS_BIAS.n286 161.3
R8694 CS_BIAS.n288 CS_BIAS.n3 161.3
R8695 CS_BIAS.n290 CS_BIAS.n289 161.3
R8696 CS_BIAS.n291 CS_BIAS.n2 161.3
R8697 CS_BIAS.n293 CS_BIAS.n292 161.3
R8698 CS_BIAS.n294 CS_BIAS.n1 161.3
R8699 CS_BIAS.n296 CS_BIAS.n295 161.3
R8700 CS_BIAS.n1761 CS_BIAS.n1760 161.3
R8701 CS_BIAS.n1759 CS_BIAS.n1619 161.3
R8702 CS_BIAS.n1758 CS_BIAS.n1757 161.3
R8703 CS_BIAS.n1756 CS_BIAS.n1620 161.3
R8704 CS_BIAS.n1755 CS_BIAS.n1754 161.3
R8705 CS_BIAS.n1753 CS_BIAS.n1621 161.3
R8706 CS_BIAS.n1752 CS_BIAS.n1751 161.3
R8707 CS_BIAS.n1750 CS_BIAS.n1622 161.3
R8708 CS_BIAS.n1749 CS_BIAS.n1748 161.3
R8709 CS_BIAS.n1747 CS_BIAS.n1623 161.3
R8710 CS_BIAS.n1746 CS_BIAS.n1745 161.3
R8711 CS_BIAS.n1744 CS_BIAS.n1743 161.3
R8712 CS_BIAS.n1742 CS_BIAS.n1625 161.3
R8713 CS_BIAS.n1741 CS_BIAS.n1740 161.3
R8714 CS_BIAS.n1739 CS_BIAS.n1626 161.3
R8715 CS_BIAS.n1738 CS_BIAS.n1737 161.3
R8716 CS_BIAS.n1736 CS_BIAS.n1627 161.3
R8717 CS_BIAS.n1735 CS_BIAS.n1734 161.3
R8718 CS_BIAS.n1733 CS_BIAS.n1628 161.3
R8719 CS_BIAS.n1732 CS_BIAS.n1731 161.3
R8720 CS_BIAS.n1730 CS_BIAS.n1629 161.3
R8721 CS_BIAS.n1729 CS_BIAS.n1728 161.3
R8722 CS_BIAS.n1727 CS_BIAS.n1726 161.3
R8723 CS_BIAS.n1725 CS_BIAS.n1631 161.3
R8724 CS_BIAS.n1724 CS_BIAS.n1723 161.3
R8725 CS_BIAS.n1722 CS_BIAS.n1632 161.3
R8726 CS_BIAS.n1721 CS_BIAS.n1720 161.3
R8727 CS_BIAS.n1719 CS_BIAS.n1633 161.3
R8728 CS_BIAS.n1718 CS_BIAS.n1717 161.3
R8729 CS_BIAS.n1716 CS_BIAS.n1634 161.3
R8730 CS_BIAS.n1715 CS_BIAS.n1714 161.3
R8731 CS_BIAS.n1713 CS_BIAS.n1635 161.3
R8732 CS_BIAS.n1712 CS_BIAS.n1711 161.3
R8733 CS_BIAS.n1710 CS_BIAS.n1636 161.3
R8734 CS_BIAS.n1709 CS_BIAS.n1708 161.3
R8735 CS_BIAS.n1706 CS_BIAS.n1637 161.3
R8736 CS_BIAS.n1705 CS_BIAS.n1704 161.3
R8737 CS_BIAS.n1703 CS_BIAS.n1638 161.3
R8738 CS_BIAS.n1702 CS_BIAS.n1701 161.3
R8739 CS_BIAS.n1700 CS_BIAS.n1639 161.3
R8740 CS_BIAS.n1699 CS_BIAS.n1698 161.3
R8741 CS_BIAS.n1697 CS_BIAS.n1640 161.3
R8742 CS_BIAS.n1696 CS_BIAS.n1695 161.3
R8743 CS_BIAS.n1694 CS_BIAS.n1641 161.3
R8744 CS_BIAS.n1693 CS_BIAS.n1692 161.3
R8745 CS_BIAS.n1691 CS_BIAS.n1690 161.3
R8746 CS_BIAS.n1689 CS_BIAS.n1643 161.3
R8747 CS_BIAS.n1688 CS_BIAS.n1687 161.3
R8748 CS_BIAS.n1686 CS_BIAS.n1644 161.3
R8749 CS_BIAS.n1685 CS_BIAS.n1684 161.3
R8750 CS_BIAS.n1683 CS_BIAS.n1645 161.3
R8751 CS_BIAS.n1682 CS_BIAS.n1681 161.3
R8752 CS_BIAS.n1680 CS_BIAS.n1646 161.3
R8753 CS_BIAS.n1679 CS_BIAS.n1678 161.3
R8754 CS_BIAS.n1677 CS_BIAS.n1647 161.3
R8755 CS_BIAS.n1676 CS_BIAS.n1675 161.3
R8756 CS_BIAS.n1674 CS_BIAS.n1648 161.3
R8757 CS_BIAS.n1673 CS_BIAS.n1672 161.3
R8758 CS_BIAS.n1670 CS_BIAS.n1649 161.3
R8759 CS_BIAS.n1669 CS_BIAS.n1668 161.3
R8760 CS_BIAS.n1667 CS_BIAS.n1650 161.3
R8761 CS_BIAS.n1666 CS_BIAS.n1665 161.3
R8762 CS_BIAS.n1664 CS_BIAS.n1651 161.3
R8763 CS_BIAS.n1663 CS_BIAS.n1662 161.3
R8764 CS_BIAS.n1661 CS_BIAS.n1652 161.3
R8765 CS_BIAS.n1660 CS_BIAS.n1659 161.3
R8766 CS_BIAS.n1658 CS_BIAS.n1653 161.3
R8767 CS_BIAS.n1657 CS_BIAS.n1656 161.3
R8768 CS_BIAS.n1615 CS_BIAS.n1614 161.3
R8769 CS_BIAS.n1613 CS_BIAS.n1473 161.3
R8770 CS_BIAS.n1612 CS_BIAS.n1611 161.3
R8771 CS_BIAS.n1610 CS_BIAS.n1474 161.3
R8772 CS_BIAS.n1609 CS_BIAS.n1608 161.3
R8773 CS_BIAS.n1607 CS_BIAS.n1475 161.3
R8774 CS_BIAS.n1606 CS_BIAS.n1605 161.3
R8775 CS_BIAS.n1604 CS_BIAS.n1476 161.3
R8776 CS_BIAS.n1603 CS_BIAS.n1602 161.3
R8777 CS_BIAS.n1601 CS_BIAS.n1477 161.3
R8778 CS_BIAS.n1600 CS_BIAS.n1599 161.3
R8779 CS_BIAS.n1598 CS_BIAS.n1597 161.3
R8780 CS_BIAS.n1596 CS_BIAS.n1479 161.3
R8781 CS_BIAS.n1595 CS_BIAS.n1594 161.3
R8782 CS_BIAS.n1593 CS_BIAS.n1480 161.3
R8783 CS_BIAS.n1592 CS_BIAS.n1591 161.3
R8784 CS_BIAS.n1590 CS_BIAS.n1481 161.3
R8785 CS_BIAS.n1589 CS_BIAS.n1588 161.3
R8786 CS_BIAS.n1587 CS_BIAS.n1482 161.3
R8787 CS_BIAS.n1586 CS_BIAS.n1585 161.3
R8788 CS_BIAS.n1584 CS_BIAS.n1483 161.3
R8789 CS_BIAS.n1583 CS_BIAS.n1582 161.3
R8790 CS_BIAS.n1581 CS_BIAS.n1580 161.3
R8791 CS_BIAS.n1579 CS_BIAS.n1485 161.3
R8792 CS_BIAS.n1578 CS_BIAS.n1577 161.3
R8793 CS_BIAS.n1576 CS_BIAS.n1486 161.3
R8794 CS_BIAS.n1575 CS_BIAS.n1574 161.3
R8795 CS_BIAS.n1573 CS_BIAS.n1487 161.3
R8796 CS_BIAS.n1572 CS_BIAS.n1571 161.3
R8797 CS_BIAS.n1570 CS_BIAS.n1488 161.3
R8798 CS_BIAS.n1569 CS_BIAS.n1568 161.3
R8799 CS_BIAS.n1567 CS_BIAS.n1489 161.3
R8800 CS_BIAS.n1566 CS_BIAS.n1565 161.3
R8801 CS_BIAS.n1564 CS_BIAS.n1490 161.3
R8802 CS_BIAS.n1563 CS_BIAS.n1562 161.3
R8803 CS_BIAS.n1560 CS_BIAS.n1491 161.3
R8804 CS_BIAS.n1559 CS_BIAS.n1558 161.3
R8805 CS_BIAS.n1557 CS_BIAS.n1492 161.3
R8806 CS_BIAS.n1556 CS_BIAS.n1555 161.3
R8807 CS_BIAS.n1554 CS_BIAS.n1493 161.3
R8808 CS_BIAS.n1553 CS_BIAS.n1552 161.3
R8809 CS_BIAS.n1551 CS_BIAS.n1494 161.3
R8810 CS_BIAS.n1550 CS_BIAS.n1549 161.3
R8811 CS_BIAS.n1548 CS_BIAS.n1495 161.3
R8812 CS_BIAS.n1547 CS_BIAS.n1546 161.3
R8813 CS_BIAS.n1545 CS_BIAS.n1544 161.3
R8814 CS_BIAS.n1543 CS_BIAS.n1497 161.3
R8815 CS_BIAS.n1542 CS_BIAS.n1541 161.3
R8816 CS_BIAS.n1540 CS_BIAS.n1498 161.3
R8817 CS_BIAS.n1539 CS_BIAS.n1538 161.3
R8818 CS_BIAS.n1537 CS_BIAS.n1499 161.3
R8819 CS_BIAS.n1536 CS_BIAS.n1535 161.3
R8820 CS_BIAS.n1534 CS_BIAS.n1500 161.3
R8821 CS_BIAS.n1533 CS_BIAS.n1532 161.3
R8822 CS_BIAS.n1531 CS_BIAS.n1501 161.3
R8823 CS_BIAS.n1530 CS_BIAS.n1529 161.3
R8824 CS_BIAS.n1528 CS_BIAS.n1502 161.3
R8825 CS_BIAS.n1527 CS_BIAS.n1526 161.3
R8826 CS_BIAS.n1524 CS_BIAS.n1503 161.3
R8827 CS_BIAS.n1523 CS_BIAS.n1522 161.3
R8828 CS_BIAS.n1521 CS_BIAS.n1504 161.3
R8829 CS_BIAS.n1520 CS_BIAS.n1519 161.3
R8830 CS_BIAS.n1518 CS_BIAS.n1505 161.3
R8831 CS_BIAS.n1517 CS_BIAS.n1516 161.3
R8832 CS_BIAS.n1515 CS_BIAS.n1506 161.3
R8833 CS_BIAS.n1514 CS_BIAS.n1513 161.3
R8834 CS_BIAS.n1512 CS_BIAS.n1507 161.3
R8835 CS_BIAS.n1511 CS_BIAS.n1510 161.3
R8836 CS_BIAS.n1469 CS_BIAS.n1468 161.3
R8837 CS_BIAS.n1467 CS_BIAS.n1327 161.3
R8838 CS_BIAS.n1466 CS_BIAS.n1465 161.3
R8839 CS_BIAS.n1464 CS_BIAS.n1328 161.3
R8840 CS_BIAS.n1463 CS_BIAS.n1462 161.3
R8841 CS_BIAS.n1461 CS_BIAS.n1329 161.3
R8842 CS_BIAS.n1460 CS_BIAS.n1459 161.3
R8843 CS_BIAS.n1458 CS_BIAS.n1330 161.3
R8844 CS_BIAS.n1457 CS_BIAS.n1456 161.3
R8845 CS_BIAS.n1455 CS_BIAS.n1331 161.3
R8846 CS_BIAS.n1454 CS_BIAS.n1453 161.3
R8847 CS_BIAS.n1452 CS_BIAS.n1451 161.3
R8848 CS_BIAS.n1450 CS_BIAS.n1333 161.3
R8849 CS_BIAS.n1449 CS_BIAS.n1448 161.3
R8850 CS_BIAS.n1447 CS_BIAS.n1334 161.3
R8851 CS_BIAS.n1446 CS_BIAS.n1445 161.3
R8852 CS_BIAS.n1444 CS_BIAS.n1335 161.3
R8853 CS_BIAS.n1443 CS_BIAS.n1442 161.3
R8854 CS_BIAS.n1441 CS_BIAS.n1336 161.3
R8855 CS_BIAS.n1440 CS_BIAS.n1439 161.3
R8856 CS_BIAS.n1438 CS_BIAS.n1337 161.3
R8857 CS_BIAS.n1437 CS_BIAS.n1436 161.3
R8858 CS_BIAS.n1435 CS_BIAS.n1434 161.3
R8859 CS_BIAS.n1433 CS_BIAS.n1339 161.3
R8860 CS_BIAS.n1432 CS_BIAS.n1431 161.3
R8861 CS_BIAS.n1430 CS_BIAS.n1340 161.3
R8862 CS_BIAS.n1429 CS_BIAS.n1428 161.3
R8863 CS_BIAS.n1427 CS_BIAS.n1341 161.3
R8864 CS_BIAS.n1426 CS_BIAS.n1425 161.3
R8865 CS_BIAS.n1424 CS_BIAS.n1342 161.3
R8866 CS_BIAS.n1423 CS_BIAS.n1422 161.3
R8867 CS_BIAS.n1421 CS_BIAS.n1343 161.3
R8868 CS_BIAS.n1420 CS_BIAS.n1419 161.3
R8869 CS_BIAS.n1418 CS_BIAS.n1344 161.3
R8870 CS_BIAS.n1417 CS_BIAS.n1416 161.3
R8871 CS_BIAS.n1414 CS_BIAS.n1345 161.3
R8872 CS_BIAS.n1413 CS_BIAS.n1412 161.3
R8873 CS_BIAS.n1411 CS_BIAS.n1346 161.3
R8874 CS_BIAS.n1410 CS_BIAS.n1409 161.3
R8875 CS_BIAS.n1408 CS_BIAS.n1347 161.3
R8876 CS_BIAS.n1407 CS_BIAS.n1406 161.3
R8877 CS_BIAS.n1405 CS_BIAS.n1348 161.3
R8878 CS_BIAS.n1404 CS_BIAS.n1403 161.3
R8879 CS_BIAS.n1402 CS_BIAS.n1349 161.3
R8880 CS_BIAS.n1401 CS_BIAS.n1400 161.3
R8881 CS_BIAS.n1399 CS_BIAS.n1398 161.3
R8882 CS_BIAS.n1397 CS_BIAS.n1351 161.3
R8883 CS_BIAS.n1396 CS_BIAS.n1395 161.3
R8884 CS_BIAS.n1394 CS_BIAS.n1352 161.3
R8885 CS_BIAS.n1393 CS_BIAS.n1392 161.3
R8886 CS_BIAS.n1391 CS_BIAS.n1353 161.3
R8887 CS_BIAS.n1390 CS_BIAS.n1389 161.3
R8888 CS_BIAS.n1388 CS_BIAS.n1354 161.3
R8889 CS_BIAS.n1387 CS_BIAS.n1386 161.3
R8890 CS_BIAS.n1385 CS_BIAS.n1355 161.3
R8891 CS_BIAS.n1384 CS_BIAS.n1383 161.3
R8892 CS_BIAS.n1382 CS_BIAS.n1356 161.3
R8893 CS_BIAS.n1381 CS_BIAS.n1380 161.3
R8894 CS_BIAS.n1378 CS_BIAS.n1357 161.3
R8895 CS_BIAS.n1377 CS_BIAS.n1376 161.3
R8896 CS_BIAS.n1375 CS_BIAS.n1358 161.3
R8897 CS_BIAS.n1374 CS_BIAS.n1373 161.3
R8898 CS_BIAS.n1372 CS_BIAS.n1359 161.3
R8899 CS_BIAS.n1371 CS_BIAS.n1370 161.3
R8900 CS_BIAS.n1369 CS_BIAS.n1360 161.3
R8901 CS_BIAS.n1368 CS_BIAS.n1367 161.3
R8902 CS_BIAS.n1366 CS_BIAS.n1361 161.3
R8903 CS_BIAS.n1365 CS_BIAS.n1364 161.3
R8904 CS_BIAS.n1323 CS_BIAS.n1322 161.3
R8905 CS_BIAS.n1321 CS_BIAS.n1181 161.3
R8906 CS_BIAS.n1320 CS_BIAS.n1319 161.3
R8907 CS_BIAS.n1318 CS_BIAS.n1182 161.3
R8908 CS_BIAS.n1317 CS_BIAS.n1316 161.3
R8909 CS_BIAS.n1315 CS_BIAS.n1183 161.3
R8910 CS_BIAS.n1314 CS_BIAS.n1313 161.3
R8911 CS_BIAS.n1312 CS_BIAS.n1184 161.3
R8912 CS_BIAS.n1311 CS_BIAS.n1310 161.3
R8913 CS_BIAS.n1309 CS_BIAS.n1185 161.3
R8914 CS_BIAS.n1308 CS_BIAS.n1307 161.3
R8915 CS_BIAS.n1306 CS_BIAS.n1305 161.3
R8916 CS_BIAS.n1304 CS_BIAS.n1187 161.3
R8917 CS_BIAS.n1303 CS_BIAS.n1302 161.3
R8918 CS_BIAS.n1301 CS_BIAS.n1188 161.3
R8919 CS_BIAS.n1300 CS_BIAS.n1299 161.3
R8920 CS_BIAS.n1298 CS_BIAS.n1189 161.3
R8921 CS_BIAS.n1297 CS_BIAS.n1296 161.3
R8922 CS_BIAS.n1295 CS_BIAS.n1190 161.3
R8923 CS_BIAS.n1294 CS_BIAS.n1293 161.3
R8924 CS_BIAS.n1292 CS_BIAS.n1191 161.3
R8925 CS_BIAS.n1291 CS_BIAS.n1290 161.3
R8926 CS_BIAS.n1289 CS_BIAS.n1288 161.3
R8927 CS_BIAS.n1287 CS_BIAS.n1193 161.3
R8928 CS_BIAS.n1286 CS_BIAS.n1285 161.3
R8929 CS_BIAS.n1284 CS_BIAS.n1194 161.3
R8930 CS_BIAS.n1283 CS_BIAS.n1282 161.3
R8931 CS_BIAS.n1281 CS_BIAS.n1195 161.3
R8932 CS_BIAS.n1280 CS_BIAS.n1279 161.3
R8933 CS_BIAS.n1278 CS_BIAS.n1196 161.3
R8934 CS_BIAS.n1277 CS_BIAS.n1276 161.3
R8935 CS_BIAS.n1275 CS_BIAS.n1197 161.3
R8936 CS_BIAS.n1274 CS_BIAS.n1273 161.3
R8937 CS_BIAS.n1272 CS_BIAS.n1198 161.3
R8938 CS_BIAS.n1271 CS_BIAS.n1270 161.3
R8939 CS_BIAS.n1268 CS_BIAS.n1199 161.3
R8940 CS_BIAS.n1267 CS_BIAS.n1266 161.3
R8941 CS_BIAS.n1265 CS_BIAS.n1200 161.3
R8942 CS_BIAS.n1264 CS_BIAS.n1263 161.3
R8943 CS_BIAS.n1262 CS_BIAS.n1201 161.3
R8944 CS_BIAS.n1261 CS_BIAS.n1260 161.3
R8945 CS_BIAS.n1259 CS_BIAS.n1202 161.3
R8946 CS_BIAS.n1258 CS_BIAS.n1257 161.3
R8947 CS_BIAS.n1256 CS_BIAS.n1203 161.3
R8948 CS_BIAS.n1255 CS_BIAS.n1254 161.3
R8949 CS_BIAS.n1253 CS_BIAS.n1252 161.3
R8950 CS_BIAS.n1251 CS_BIAS.n1205 161.3
R8951 CS_BIAS.n1250 CS_BIAS.n1249 161.3
R8952 CS_BIAS.n1248 CS_BIAS.n1206 161.3
R8953 CS_BIAS.n1247 CS_BIAS.n1246 161.3
R8954 CS_BIAS.n1245 CS_BIAS.n1207 161.3
R8955 CS_BIAS.n1244 CS_BIAS.n1243 161.3
R8956 CS_BIAS.n1242 CS_BIAS.n1208 161.3
R8957 CS_BIAS.n1241 CS_BIAS.n1240 161.3
R8958 CS_BIAS.n1239 CS_BIAS.n1209 161.3
R8959 CS_BIAS.n1238 CS_BIAS.n1237 161.3
R8960 CS_BIAS.n1236 CS_BIAS.n1210 161.3
R8961 CS_BIAS.n1235 CS_BIAS.n1234 161.3
R8962 CS_BIAS.n1232 CS_BIAS.n1211 161.3
R8963 CS_BIAS.n1231 CS_BIAS.n1230 161.3
R8964 CS_BIAS.n1229 CS_BIAS.n1212 161.3
R8965 CS_BIAS.n1228 CS_BIAS.n1227 161.3
R8966 CS_BIAS.n1226 CS_BIAS.n1213 161.3
R8967 CS_BIAS.n1225 CS_BIAS.n1224 161.3
R8968 CS_BIAS.n1223 CS_BIAS.n1214 161.3
R8969 CS_BIAS.n1222 CS_BIAS.n1221 161.3
R8970 CS_BIAS.n1220 CS_BIAS.n1215 161.3
R8971 CS_BIAS.n1219 CS_BIAS.n1218 161.3
R8972 CS_BIAS.n1049 CS_BIAS.n1048 161.3
R8973 CS_BIAS.n1047 CS_BIAS.n907 161.3
R8974 CS_BIAS.n1046 CS_BIAS.n1045 161.3
R8975 CS_BIAS.n1044 CS_BIAS.n908 161.3
R8976 CS_BIAS.n1043 CS_BIAS.n1042 161.3
R8977 CS_BIAS.n1041 CS_BIAS.n909 161.3
R8978 CS_BIAS.n1040 CS_BIAS.n1039 161.3
R8979 CS_BIAS.n1038 CS_BIAS.n910 161.3
R8980 CS_BIAS.n1037 CS_BIAS.n1036 161.3
R8981 CS_BIAS.n1035 CS_BIAS.n911 161.3
R8982 CS_BIAS.n1034 CS_BIAS.n1033 161.3
R8983 CS_BIAS.n1032 CS_BIAS.n1031 161.3
R8984 CS_BIAS.n1030 CS_BIAS.n913 161.3
R8985 CS_BIAS.n1029 CS_BIAS.n1028 161.3
R8986 CS_BIAS.n1027 CS_BIAS.n914 161.3
R8987 CS_BIAS.n1026 CS_BIAS.n1025 161.3
R8988 CS_BIAS.n1024 CS_BIAS.n915 161.3
R8989 CS_BIAS.n1023 CS_BIAS.n1022 161.3
R8990 CS_BIAS.n1021 CS_BIAS.n916 161.3
R8991 CS_BIAS.n1020 CS_BIAS.n1019 161.3
R8992 CS_BIAS.n1018 CS_BIAS.n917 161.3
R8993 CS_BIAS.n1017 CS_BIAS.n1016 161.3
R8994 CS_BIAS.n1015 CS_BIAS.n1014 161.3
R8995 CS_BIAS.n1013 CS_BIAS.n919 161.3
R8996 CS_BIAS.n1012 CS_BIAS.n1011 161.3
R8997 CS_BIAS.n1010 CS_BIAS.n920 161.3
R8998 CS_BIAS.n1009 CS_BIAS.n1008 161.3
R8999 CS_BIAS.n1007 CS_BIAS.n921 161.3
R9000 CS_BIAS.n1006 CS_BIAS.n1005 161.3
R9001 CS_BIAS.n1004 CS_BIAS.n922 161.3
R9002 CS_BIAS.n1003 CS_BIAS.n1002 161.3
R9003 CS_BIAS.n1001 CS_BIAS.n923 161.3
R9004 CS_BIAS.n1000 CS_BIAS.n999 161.3
R9005 CS_BIAS.n998 CS_BIAS.n924 161.3
R9006 CS_BIAS.n997 CS_BIAS.n996 161.3
R9007 CS_BIAS.n994 CS_BIAS.n925 161.3
R9008 CS_BIAS.n993 CS_BIAS.n992 161.3
R9009 CS_BIAS.n991 CS_BIAS.n926 161.3
R9010 CS_BIAS.n990 CS_BIAS.n989 161.3
R9011 CS_BIAS.n988 CS_BIAS.n927 161.3
R9012 CS_BIAS.n987 CS_BIAS.n986 161.3
R9013 CS_BIAS.n985 CS_BIAS.n928 161.3
R9014 CS_BIAS.n984 CS_BIAS.n983 161.3
R9015 CS_BIAS.n982 CS_BIAS.n929 161.3
R9016 CS_BIAS.n981 CS_BIAS.n980 161.3
R9017 CS_BIAS.n979 CS_BIAS.n978 161.3
R9018 CS_BIAS.n977 CS_BIAS.n931 161.3
R9019 CS_BIAS.n976 CS_BIAS.n975 161.3
R9020 CS_BIAS.n974 CS_BIAS.n932 161.3
R9021 CS_BIAS.n973 CS_BIAS.n972 161.3
R9022 CS_BIAS.n971 CS_BIAS.n933 161.3
R9023 CS_BIAS.n970 CS_BIAS.n969 161.3
R9024 CS_BIAS.n968 CS_BIAS.n934 161.3
R9025 CS_BIAS.n967 CS_BIAS.n966 161.3
R9026 CS_BIAS.n965 CS_BIAS.n935 161.3
R9027 CS_BIAS.n964 CS_BIAS.n963 161.3
R9028 CS_BIAS.n962 CS_BIAS.n936 161.3
R9029 CS_BIAS.n961 CS_BIAS.n960 161.3
R9030 CS_BIAS.n958 CS_BIAS.n937 161.3
R9031 CS_BIAS.n957 CS_BIAS.n956 161.3
R9032 CS_BIAS.n955 CS_BIAS.n938 161.3
R9033 CS_BIAS.n954 CS_BIAS.n953 161.3
R9034 CS_BIAS.n952 CS_BIAS.n939 161.3
R9035 CS_BIAS.n951 CS_BIAS.n950 161.3
R9036 CS_BIAS.n949 CS_BIAS.n940 161.3
R9037 CS_BIAS.n948 CS_BIAS.n947 161.3
R9038 CS_BIAS.n946 CS_BIAS.n941 161.3
R9039 CS_BIAS.n945 CS_BIAS.n944 161.3
R9040 CS_BIAS.n1116 CS_BIAS.n1115 161.3
R9041 CS_BIAS.n1114 CS_BIAS.n1057 161.3
R9042 CS_BIAS.n1113 CS_BIAS.n1112 161.3
R9043 CS_BIAS.n1111 CS_BIAS.n1058 161.3
R9044 CS_BIAS.n1110 CS_BIAS.n1109 161.3
R9045 CS_BIAS.n1108 CS_BIAS.n1107 161.3
R9046 CS_BIAS.n1106 CS_BIAS.n1060 161.3
R9047 CS_BIAS.n1105 CS_BIAS.n1104 161.3
R9048 CS_BIAS.n1103 CS_BIAS.n1061 161.3
R9049 CS_BIAS.n1102 CS_BIAS.n1101 161.3
R9050 CS_BIAS.n1100 CS_BIAS.n1062 161.3
R9051 CS_BIAS.n1099 CS_BIAS.n1098 161.3
R9052 CS_BIAS.n1097 CS_BIAS.n1063 161.3
R9053 CS_BIAS.n1096 CS_BIAS.n1095 161.3
R9054 CS_BIAS.n1094 CS_BIAS.n1064 161.3
R9055 CS_BIAS.n1093 CS_BIAS.n1092 161.3
R9056 CS_BIAS.n1091 CS_BIAS.n1065 161.3
R9057 CS_BIAS.n1090 CS_BIAS.n1089 161.3
R9058 CS_BIAS.n1087 CS_BIAS.n1066 161.3
R9059 CS_BIAS.n1086 CS_BIAS.n1085 161.3
R9060 CS_BIAS.n1084 CS_BIAS.n1067 161.3
R9061 CS_BIAS.n1083 CS_BIAS.n1082 161.3
R9062 CS_BIAS.n1081 CS_BIAS.n1068 161.3
R9063 CS_BIAS.n1080 CS_BIAS.n1079 161.3
R9064 CS_BIAS.n1078 CS_BIAS.n1069 161.3
R9065 CS_BIAS.n1077 CS_BIAS.n1076 161.3
R9066 CS_BIAS.n1075 CS_BIAS.n1070 161.3
R9067 CS_BIAS.n1074 CS_BIAS.n1073 161.3
R9068 CS_BIAS.n1117 CS_BIAS.n1056 161.3
R9069 CS_BIAS.n1178 CS_BIAS.n1177 161.3
R9070 CS_BIAS.n1176 CS_BIAS.n883 161.3
R9071 CS_BIAS.n1175 CS_BIAS.n1174 161.3
R9072 CS_BIAS.n1173 CS_BIAS.n884 161.3
R9073 CS_BIAS.n1172 CS_BIAS.n1171 161.3
R9074 CS_BIAS.n1170 CS_BIAS.n885 161.3
R9075 CS_BIAS.n1169 CS_BIAS.n1168 161.3
R9076 CS_BIAS.n1167 CS_BIAS.n886 161.3
R9077 CS_BIAS.n1166 CS_BIAS.n1165 161.3
R9078 CS_BIAS.n1164 CS_BIAS.n887 161.3
R9079 CS_BIAS.n1163 CS_BIAS.n1162 161.3
R9080 CS_BIAS.n1161 CS_BIAS.n1160 161.3
R9081 CS_BIAS.n1159 CS_BIAS.n889 161.3
R9082 CS_BIAS.n1158 CS_BIAS.n1157 161.3
R9083 CS_BIAS.n1156 CS_BIAS.n890 161.3
R9084 CS_BIAS.n1155 CS_BIAS.n1154 161.3
R9085 CS_BIAS.n1153 CS_BIAS.n891 161.3
R9086 CS_BIAS.n1152 CS_BIAS.n1151 161.3
R9087 CS_BIAS.n1150 CS_BIAS.n892 161.3
R9088 CS_BIAS.n1149 CS_BIAS.n1148 161.3
R9089 CS_BIAS.n1147 CS_BIAS.n893 161.3
R9090 CS_BIAS.n1146 CS_BIAS.n1145 161.3
R9091 CS_BIAS.n1144 CS_BIAS.n1143 161.3
R9092 CS_BIAS.n1142 CS_BIAS.n895 161.3
R9093 CS_BIAS.n1141 CS_BIAS.n1140 161.3
R9094 CS_BIAS.n1139 CS_BIAS.n896 161.3
R9095 CS_BIAS.n1138 CS_BIAS.n1137 161.3
R9096 CS_BIAS.n1136 CS_BIAS.n897 161.3
R9097 CS_BIAS.n1135 CS_BIAS.n1134 161.3
R9098 CS_BIAS.n1133 CS_BIAS.n898 161.3
R9099 CS_BIAS.n1132 CS_BIAS.n1131 161.3
R9100 CS_BIAS.n1130 CS_BIAS.n899 161.3
R9101 CS_BIAS.n1129 CS_BIAS.n1128 161.3
R9102 CS_BIAS.n1127 CS_BIAS.n900 161.3
R9103 CS_BIAS.n1126 CS_BIAS.n1125 161.3
R9104 CS_BIAS.n1123 CS_BIAS.n901 161.3
R9105 CS_BIAS.n1122 CS_BIAS.n1121 161.3
R9106 CS_BIAS.n1120 CS_BIAS.n902 161.3
R9107 CS_BIAS.n1119 CS_BIAS.n1118 161.3
R9108 CS_BIAS.n173 CS_BIAS.n171 78.5929
R9109 CS_BIAS.n905 CS_BIAS.n903 78.5929
R9110 CS_BIAS.n173 CS_BIAS.n172 76.9579
R9111 CS_BIAS.n170 CS_BIAS.n169 76.9579
R9112 CS_BIAS.n168 CS_BIAS.n167 76.9579
R9113 CS_BIAS.n1052 CS_BIAS.n1051 76.9579
R9114 CS_BIAS.n1054 CS_BIAS.n1053 76.9579
R9115 CS_BIAS.n905 CS_BIAS.n904 76.9579
R9116 CS_BIAS.n802 CS_BIAS.n801 73.0308
R9117 CS_BIAS.n837 CS_BIAS.n836 73.0308
R9118 CS_BIAS.n691 CS_BIAS.n690 73.0308
R9119 CS_BIAS.n656 CS_BIAS.n655 73.0308
R9120 CS_BIAS.n545 CS_BIAS.n544 73.0308
R9121 CS_BIAS.n510 CS_BIAS.n509 73.0308
R9122 CS_BIAS.n399 CS_BIAS.n398 73.0308
R9123 CS_BIAS.n364 CS_BIAS.n363 73.0308
R9124 CS_BIAS.n123 CS_BIAS.n122 73.0308
R9125 CS_BIAS.n88 CS_BIAS.n87 73.0308
R9126 CS_BIAS.n254 CS_BIAS.n253 73.0308
R9127 CS_BIAS.n219 CS_BIAS.n218 73.0308
R9128 CS_BIAS.n1683 CS_BIAS.n1682 73.0308
R9129 CS_BIAS.n1719 CS_BIAS.n1718 73.0308
R9130 CS_BIAS.n1537 CS_BIAS.n1536 73.0308
R9131 CS_BIAS.n1573 CS_BIAS.n1572 73.0308
R9132 CS_BIAS.n1391 CS_BIAS.n1390 73.0308
R9133 CS_BIAS.n1427 CS_BIAS.n1426 73.0308
R9134 CS_BIAS.n1245 CS_BIAS.n1244 73.0308
R9135 CS_BIAS.n1281 CS_BIAS.n1280 73.0308
R9136 CS_BIAS.n971 CS_BIAS.n970 73.0308
R9137 CS_BIAS.n1007 CS_BIAS.n1006 73.0308
R9138 CS_BIAS.n1136 CS_BIAS.n1135 73.0308
R9139 CS_BIAS.n1100 CS_BIAS.n1099 73.0308
R9140 CS_BIAS.n785 CS_BIAS.n784 68.1745
R9141 CS_BIAS.n854 CS_BIAS.n853 68.1745
R9142 CS_BIAS.n708 CS_BIAS.n707 68.1745
R9143 CS_BIAS.n639 CS_BIAS.n638 68.1745
R9144 CS_BIAS.n562 CS_BIAS.n561 68.1745
R9145 CS_BIAS.n493 CS_BIAS.n492 68.1745
R9146 CS_BIAS.n416 CS_BIAS.n415 68.1745
R9147 CS_BIAS.n347 CS_BIAS.n346 68.1745
R9148 CS_BIAS.n140 CS_BIAS.n139 68.1745
R9149 CS_BIAS.n71 CS_BIAS.n70 68.1745
R9150 CS_BIAS.n271 CS_BIAS.n270 68.1745
R9151 CS_BIAS.n202 CS_BIAS.n201 68.1745
R9152 CS_BIAS.n1665 CS_BIAS.n1664 68.1745
R9153 CS_BIAS.n1736 CS_BIAS.n1735 68.1745
R9154 CS_BIAS.n1519 CS_BIAS.n1518 68.1745
R9155 CS_BIAS.n1590 CS_BIAS.n1589 68.1745
R9156 CS_BIAS.n1373 CS_BIAS.n1372 68.1745
R9157 CS_BIAS.n1444 CS_BIAS.n1443 68.1745
R9158 CS_BIAS.n1227 CS_BIAS.n1226 68.1745
R9159 CS_BIAS.n1298 CS_BIAS.n1297 68.1745
R9160 CS_BIAS.n953 CS_BIAS.n952 68.1745
R9161 CS_BIAS.n1024 CS_BIAS.n1023 68.1745
R9162 CS_BIAS.n1153 CS_BIAS.n1152 68.1745
R9163 CS_BIAS.n1082 CS_BIAS.n1081 68.1745
R9164 CS_BIAS.n629 CS_BIAS.n628 65.1383
R9165 CS_BIAS.n483 CS_BIAS.n482 65.1383
R9166 CS_BIAS.n337 CS_BIAS.n336 65.1383
R9167 CS_BIAS.n61 CS_BIAS.n60 65.1383
R9168 CS_BIAS.n192 CS_BIAS.n191 65.1383
R9169 CS_BIAS.n775 CS_BIAS.n774 65.1383
R9170 CS_BIAS.n1655 CS_BIAS.n1654 65.1383
R9171 CS_BIAS.n1509 CS_BIAS.n1508 65.1383
R9172 CS_BIAS.n1363 CS_BIAS.n1362 65.1383
R9173 CS_BIAS.n1217 CS_BIAS.n1216 65.1383
R9174 CS_BIAS.n943 CS_BIAS.n942 65.1383
R9175 CS_BIAS.n1072 CS_BIAS.n1071 65.1383
R9176 CS_BIAS.n872 CS_BIAS.n871 63.3181
R9177 CS_BIAS.n726 CS_BIAS.n725 63.3181
R9178 CS_BIAS.n580 CS_BIAS.n579 63.3181
R9179 CS_BIAS.n434 CS_BIAS.n433 63.3181
R9180 CS_BIAS.n158 CS_BIAS.n157 63.3181
R9181 CS_BIAS.n289 CS_BIAS.n288 63.3181
R9182 CS_BIAS.n1754 CS_BIAS.n1753 63.3181
R9183 CS_BIAS.n1608 CS_BIAS.n1607 63.3181
R9184 CS_BIAS.n1462 CS_BIAS.n1461 63.3181
R9185 CS_BIAS.n1316 CS_BIAS.n1315 63.3181
R9186 CS_BIAS.n1042 CS_BIAS.n1041 63.3181
R9187 CS_BIAS.n1171 CS_BIAS.n1170 63.3181
R9188 CS_BIAS.n880 CS_BIAS.n736 58.5103
R9189 CS_BIAS.n734 CS_BIAS.n590 58.5103
R9190 CS_BIAS.n588 CS_BIAS.n444 58.5103
R9191 CS_BIAS.n442 CS_BIAS.n298 58.5103
R9192 CS_BIAS.n166 CS_BIAS.n22 58.5103
R9193 CS_BIAS.n297 CS_BIAS.n0 58.5103
R9194 CS_BIAS.n1762 CS_BIAS.n1618 58.5103
R9195 CS_BIAS.n1616 CS_BIAS.n1472 58.5103
R9196 CS_BIAS.n1470 CS_BIAS.n1326 58.5103
R9197 CS_BIAS.n1324 CS_BIAS.n1180 58.5103
R9198 CS_BIAS.n1050 CS_BIAS.n906 58.5103
R9199 CS_BIAS.n1179 CS_BIAS.n882 58.5103
R9200 CS_BIAS.n819 CS_BIAS.n818 56.5193
R9201 CS_BIAS.n820 CS_BIAS.n819 56.5193
R9202 CS_BIAS.n674 CS_BIAS.n673 56.5193
R9203 CS_BIAS.n673 CS_BIAS.n672 56.5193
R9204 CS_BIAS.n528 CS_BIAS.n527 56.5193
R9205 CS_BIAS.n527 CS_BIAS.n526 56.5193
R9206 CS_BIAS.n382 CS_BIAS.n381 56.5193
R9207 CS_BIAS.n381 CS_BIAS.n380 56.5193
R9208 CS_BIAS.n106 CS_BIAS.n105 56.5193
R9209 CS_BIAS.n105 CS_BIAS.n104 56.5193
R9210 CS_BIAS.n237 CS_BIAS.n236 56.5193
R9211 CS_BIAS.n236 CS_BIAS.n235 56.5193
R9212 CS_BIAS.n1700 CS_BIAS.n1699 56.5193
R9213 CS_BIAS.n1701 CS_BIAS.n1700 56.5193
R9214 CS_BIAS.n1554 CS_BIAS.n1553 56.5193
R9215 CS_BIAS.n1555 CS_BIAS.n1554 56.5193
R9216 CS_BIAS.n1408 CS_BIAS.n1407 56.5193
R9217 CS_BIAS.n1409 CS_BIAS.n1408 56.5193
R9218 CS_BIAS.n1262 CS_BIAS.n1261 56.5193
R9219 CS_BIAS.n1263 CS_BIAS.n1262 56.5193
R9220 CS_BIAS.n988 CS_BIAS.n987 56.5193
R9221 CS_BIAS.n989 CS_BIAS.n988 56.5193
R9222 CS_BIAS.n1118 CS_BIAS.n1117 56.5193
R9223 CS_BIAS.n1117 CS_BIAS.n1116 56.5193
R9224 CS_BIAS.n871 CS_BIAS.n870 49.7204
R9225 CS_BIAS.n725 CS_BIAS.n724 49.7204
R9226 CS_BIAS.n579 CS_BIAS.n578 49.7204
R9227 CS_BIAS.n433 CS_BIAS.n432 49.7204
R9228 CS_BIAS.n157 CS_BIAS.n156 49.7204
R9229 CS_BIAS.n288 CS_BIAS.n287 49.7204
R9230 CS_BIAS.n1753 CS_BIAS.n1752 49.7204
R9231 CS_BIAS.n1607 CS_BIAS.n1606 49.7204
R9232 CS_BIAS.n1461 CS_BIAS.n1460 49.7204
R9233 CS_BIAS.n1315 CS_BIAS.n1314 49.7204
R9234 CS_BIAS.n1041 CS_BIAS.n1040 49.7204
R9235 CS_BIAS.n1170 CS_BIAS.n1169 49.7204
R9236 CS_BIAS.n775 CS_BIAS.t101 46.6798
R9237 CS_BIAS.n1655 CS_BIAS.t42 46.6798
R9238 CS_BIAS.n1509 CS_BIAS.t88 46.6798
R9239 CS_BIAS.n1363 CS_BIAS.t75 46.6798
R9240 CS_BIAS.n1217 CS_BIAS.t66 46.6798
R9241 CS_BIAS.n943 CS_BIAS.t30 46.6798
R9242 CS_BIAS.n1072 CS_BIAS.t38 46.6798
R9243 CS_BIAS.n629 CS_BIAS.t60 46.6796
R9244 CS_BIAS.n483 CS_BIAS.t71 46.6796
R9245 CS_BIAS.n337 CS_BIAS.t39 46.6796
R9246 CS_BIAS.n61 CS_BIAS.t18 46.6796
R9247 CS_BIAS.n192 CS_BIAS.t61 46.6796
R9248 CS_BIAS.n784 CS_BIAS.n783 44.8641
R9249 CS_BIAS.n855 CS_BIAS.n854 44.8641
R9250 CS_BIAS.n709 CS_BIAS.n708 44.8641
R9251 CS_BIAS.n638 CS_BIAS.n637 44.8641
R9252 CS_BIAS.n563 CS_BIAS.n562 44.8641
R9253 CS_BIAS.n492 CS_BIAS.n491 44.8641
R9254 CS_BIAS.n417 CS_BIAS.n416 44.8641
R9255 CS_BIAS.n346 CS_BIAS.n345 44.8641
R9256 CS_BIAS.n141 CS_BIAS.n140 44.8641
R9257 CS_BIAS.n70 CS_BIAS.n69 44.8641
R9258 CS_BIAS.n272 CS_BIAS.n271 44.8641
R9259 CS_BIAS.n201 CS_BIAS.n200 44.8641
R9260 CS_BIAS.n1664 CS_BIAS.n1663 44.8641
R9261 CS_BIAS.n1737 CS_BIAS.n1736 44.8641
R9262 CS_BIAS.n1518 CS_BIAS.n1517 44.8641
R9263 CS_BIAS.n1591 CS_BIAS.n1590 44.8641
R9264 CS_BIAS.n1372 CS_BIAS.n1371 44.8641
R9265 CS_BIAS.n1445 CS_BIAS.n1444 44.8641
R9266 CS_BIAS.n1226 CS_BIAS.n1225 44.8641
R9267 CS_BIAS.n1299 CS_BIAS.n1298 44.8641
R9268 CS_BIAS.n952 CS_BIAS.n951 44.8641
R9269 CS_BIAS.n1025 CS_BIAS.n1024 44.8641
R9270 CS_BIAS.n1154 CS_BIAS.n1153 44.8641
R9271 CS_BIAS.n1081 CS_BIAS.n1080 44.8641
R9272 CS_BIAS.n803 CS_BIAS.n802 38.0652
R9273 CS_BIAS.n836 CS_BIAS.n752 38.0652
R9274 CS_BIAS.n690 CS_BIAS.n606 38.0652
R9275 CS_BIAS.n657 CS_BIAS.n656 38.0652
R9276 CS_BIAS.n544 CS_BIAS.n460 38.0652
R9277 CS_BIAS.n511 CS_BIAS.n510 38.0652
R9278 CS_BIAS.n398 CS_BIAS.n314 38.0652
R9279 CS_BIAS.n365 CS_BIAS.n364 38.0652
R9280 CS_BIAS.n122 CS_BIAS.n38 38.0652
R9281 CS_BIAS.n89 CS_BIAS.n88 38.0652
R9282 CS_BIAS.n253 CS_BIAS.n16 38.0652
R9283 CS_BIAS.n220 CS_BIAS.n219 38.0652
R9284 CS_BIAS.n1684 CS_BIAS.n1683 38.0652
R9285 CS_BIAS.n1718 CS_BIAS.n1634 38.0652
R9286 CS_BIAS.n1538 CS_BIAS.n1537 38.0652
R9287 CS_BIAS.n1572 CS_BIAS.n1488 38.0652
R9288 CS_BIAS.n1392 CS_BIAS.n1391 38.0652
R9289 CS_BIAS.n1426 CS_BIAS.n1342 38.0652
R9290 CS_BIAS.n1246 CS_BIAS.n1245 38.0652
R9291 CS_BIAS.n1280 CS_BIAS.n1196 38.0652
R9292 CS_BIAS.n972 CS_BIAS.n971 38.0652
R9293 CS_BIAS.n1006 CS_BIAS.n922 38.0652
R9294 CS_BIAS.n1135 CS_BIAS.n898 38.0652
R9295 CS_BIAS.n1101 CS_BIAS.n1100 38.0652
R9296 CS_BIAS.n801 CS_BIAS.n765 26.41
R9297 CS_BIAS.n838 CS_BIAS.n837 26.41
R9298 CS_BIAS.n692 CS_BIAS.n691 26.41
R9299 CS_BIAS.n655 CS_BIAS.n619 26.41
R9300 CS_BIAS.n546 CS_BIAS.n545 26.41
R9301 CS_BIAS.n509 CS_BIAS.n473 26.41
R9302 CS_BIAS.n400 CS_BIAS.n399 26.41
R9303 CS_BIAS.n363 CS_BIAS.n327 26.41
R9304 CS_BIAS.n124 CS_BIAS.n123 26.41
R9305 CS_BIAS.n87 CS_BIAS.n51 26.41
R9306 CS_BIAS.n255 CS_BIAS.n254 26.41
R9307 CS_BIAS.n218 CS_BIAS.n182 26.41
R9308 CS_BIAS.n1682 CS_BIAS.n1646 26.41
R9309 CS_BIAS.n1720 CS_BIAS.n1719 26.41
R9310 CS_BIAS.n1536 CS_BIAS.n1500 26.41
R9311 CS_BIAS.n1574 CS_BIAS.n1573 26.41
R9312 CS_BIAS.n1390 CS_BIAS.n1354 26.41
R9313 CS_BIAS.n1428 CS_BIAS.n1427 26.41
R9314 CS_BIAS.n1244 CS_BIAS.n1208 26.41
R9315 CS_BIAS.n1282 CS_BIAS.n1281 26.41
R9316 CS_BIAS.n970 CS_BIAS.n934 26.41
R9317 CS_BIAS.n1008 CS_BIAS.n1007 26.41
R9318 CS_BIAS.n1137 CS_BIAS.n1136 26.41
R9319 CS_BIAS.n1099 CS_BIAS.n1063 26.41
R9320 CS_BIAS.n783 CS_BIAS.n772 24.4675
R9321 CS_BIAS.n779 CS_BIAS.n772 24.4675
R9322 CS_BIAS.n779 CS_BIAS.n778 24.4675
R9323 CS_BIAS.n778 CS_BIAS.n777 24.4675
R9324 CS_BIAS.n797 CS_BIAS.n765 24.4675
R9325 CS_BIAS.n797 CS_BIAS.n796 24.4675
R9326 CS_BIAS.n796 CS_BIAS.n795 24.4675
R9327 CS_BIAS.n795 CS_BIAS.n767 24.4675
R9328 CS_BIAS.n791 CS_BIAS.n790 24.4675
R9329 CS_BIAS.n790 CS_BIAS.n789 24.4675
R9330 CS_BIAS.n789 CS_BIAS.n770 24.4675
R9331 CS_BIAS.n785 CS_BIAS.n770 24.4675
R9332 CS_BIAS.n818 CS_BIAS.n759 24.4675
R9333 CS_BIAS.n814 CS_BIAS.n759 24.4675
R9334 CS_BIAS.n814 CS_BIAS.n813 24.4675
R9335 CS_BIAS.n813 CS_BIAS.n812 24.4675
R9336 CS_BIAS.n809 CS_BIAS.n808 24.4675
R9337 CS_BIAS.n808 CS_BIAS.n807 24.4675
R9338 CS_BIAS.n807 CS_BIAS.n763 24.4675
R9339 CS_BIAS.n803 CS_BIAS.n763 24.4675
R9340 CS_BIAS.n832 CS_BIAS.n752 24.4675
R9341 CS_BIAS.n832 CS_BIAS.n831 24.4675
R9342 CS_BIAS.n831 CS_BIAS.n830 24.4675
R9343 CS_BIAS.n830 CS_BIAS.n754 24.4675
R9344 CS_BIAS.n826 CS_BIAS.n825 24.4675
R9345 CS_BIAS.n825 CS_BIAS.n824 24.4675
R9346 CS_BIAS.n824 CS_BIAS.n757 24.4675
R9347 CS_BIAS.n820 CS_BIAS.n757 24.4675
R9348 CS_BIAS.n853 CS_BIAS.n746 24.4675
R9349 CS_BIAS.n849 CS_BIAS.n746 24.4675
R9350 CS_BIAS.n849 CS_BIAS.n848 24.4675
R9351 CS_BIAS.n848 CS_BIAS.n847 24.4675
R9352 CS_BIAS.n844 CS_BIAS.n843 24.4675
R9353 CS_BIAS.n843 CS_BIAS.n842 24.4675
R9354 CS_BIAS.n842 CS_BIAS.n750 24.4675
R9355 CS_BIAS.n838 CS_BIAS.n750 24.4675
R9356 CS_BIAS.n870 CS_BIAS.n740 24.4675
R9357 CS_BIAS.n866 CS_BIAS.n740 24.4675
R9358 CS_BIAS.n866 CS_BIAS.n865 24.4675
R9359 CS_BIAS.n865 CS_BIAS.n864 24.4675
R9360 CS_BIAS.n861 CS_BIAS.n860 24.4675
R9361 CS_BIAS.n860 CS_BIAS.n859 24.4675
R9362 CS_BIAS.n859 CS_BIAS.n744 24.4675
R9363 CS_BIAS.n855 CS_BIAS.n744 24.4675
R9364 CS_BIAS.n878 CS_BIAS.n877 24.4675
R9365 CS_BIAS.n877 CS_BIAS.n876 24.4675
R9366 CS_BIAS.n876 CS_BIAS.n738 24.4675
R9367 CS_BIAS.n872 CS_BIAS.n738 24.4675
R9368 CS_BIAS.n732 CS_BIAS.n731 24.4675
R9369 CS_BIAS.n731 CS_BIAS.n730 24.4675
R9370 CS_BIAS.n730 CS_BIAS.n592 24.4675
R9371 CS_BIAS.n726 CS_BIAS.n592 24.4675
R9372 CS_BIAS.n724 CS_BIAS.n594 24.4675
R9373 CS_BIAS.n720 CS_BIAS.n594 24.4675
R9374 CS_BIAS.n720 CS_BIAS.n719 24.4675
R9375 CS_BIAS.n719 CS_BIAS.n718 24.4675
R9376 CS_BIAS.n715 CS_BIAS.n714 24.4675
R9377 CS_BIAS.n714 CS_BIAS.n713 24.4675
R9378 CS_BIAS.n713 CS_BIAS.n598 24.4675
R9379 CS_BIAS.n709 CS_BIAS.n598 24.4675
R9380 CS_BIAS.n707 CS_BIAS.n600 24.4675
R9381 CS_BIAS.n703 CS_BIAS.n600 24.4675
R9382 CS_BIAS.n703 CS_BIAS.n702 24.4675
R9383 CS_BIAS.n702 CS_BIAS.n701 24.4675
R9384 CS_BIAS.n698 CS_BIAS.n697 24.4675
R9385 CS_BIAS.n697 CS_BIAS.n696 24.4675
R9386 CS_BIAS.n696 CS_BIAS.n604 24.4675
R9387 CS_BIAS.n692 CS_BIAS.n604 24.4675
R9388 CS_BIAS.n686 CS_BIAS.n606 24.4675
R9389 CS_BIAS.n686 CS_BIAS.n685 24.4675
R9390 CS_BIAS.n685 CS_BIAS.n684 24.4675
R9391 CS_BIAS.n684 CS_BIAS.n608 24.4675
R9392 CS_BIAS.n680 CS_BIAS.n679 24.4675
R9393 CS_BIAS.n679 CS_BIAS.n678 24.4675
R9394 CS_BIAS.n678 CS_BIAS.n611 24.4675
R9395 CS_BIAS.n674 CS_BIAS.n611 24.4675
R9396 CS_BIAS.n672 CS_BIAS.n613 24.4675
R9397 CS_BIAS.n668 CS_BIAS.n613 24.4675
R9398 CS_BIAS.n668 CS_BIAS.n667 24.4675
R9399 CS_BIAS.n667 CS_BIAS.n666 24.4675
R9400 CS_BIAS.n663 CS_BIAS.n662 24.4675
R9401 CS_BIAS.n662 CS_BIAS.n661 24.4675
R9402 CS_BIAS.n661 CS_BIAS.n617 24.4675
R9403 CS_BIAS.n657 CS_BIAS.n617 24.4675
R9404 CS_BIAS.n651 CS_BIAS.n619 24.4675
R9405 CS_BIAS.n651 CS_BIAS.n650 24.4675
R9406 CS_BIAS.n650 CS_BIAS.n649 24.4675
R9407 CS_BIAS.n649 CS_BIAS.n621 24.4675
R9408 CS_BIAS.n645 CS_BIAS.n644 24.4675
R9409 CS_BIAS.n644 CS_BIAS.n643 24.4675
R9410 CS_BIAS.n643 CS_BIAS.n624 24.4675
R9411 CS_BIAS.n639 CS_BIAS.n624 24.4675
R9412 CS_BIAS.n637 CS_BIAS.n626 24.4675
R9413 CS_BIAS.n633 CS_BIAS.n626 24.4675
R9414 CS_BIAS.n633 CS_BIAS.n632 24.4675
R9415 CS_BIAS.n632 CS_BIAS.n631 24.4675
R9416 CS_BIAS.n586 CS_BIAS.n585 24.4675
R9417 CS_BIAS.n585 CS_BIAS.n584 24.4675
R9418 CS_BIAS.n584 CS_BIAS.n446 24.4675
R9419 CS_BIAS.n580 CS_BIAS.n446 24.4675
R9420 CS_BIAS.n578 CS_BIAS.n448 24.4675
R9421 CS_BIAS.n574 CS_BIAS.n448 24.4675
R9422 CS_BIAS.n574 CS_BIAS.n573 24.4675
R9423 CS_BIAS.n573 CS_BIAS.n572 24.4675
R9424 CS_BIAS.n569 CS_BIAS.n568 24.4675
R9425 CS_BIAS.n568 CS_BIAS.n567 24.4675
R9426 CS_BIAS.n567 CS_BIAS.n452 24.4675
R9427 CS_BIAS.n563 CS_BIAS.n452 24.4675
R9428 CS_BIAS.n561 CS_BIAS.n454 24.4675
R9429 CS_BIAS.n557 CS_BIAS.n454 24.4675
R9430 CS_BIAS.n557 CS_BIAS.n556 24.4675
R9431 CS_BIAS.n556 CS_BIAS.n555 24.4675
R9432 CS_BIAS.n552 CS_BIAS.n551 24.4675
R9433 CS_BIAS.n551 CS_BIAS.n550 24.4675
R9434 CS_BIAS.n550 CS_BIAS.n458 24.4675
R9435 CS_BIAS.n546 CS_BIAS.n458 24.4675
R9436 CS_BIAS.n540 CS_BIAS.n460 24.4675
R9437 CS_BIAS.n540 CS_BIAS.n539 24.4675
R9438 CS_BIAS.n539 CS_BIAS.n538 24.4675
R9439 CS_BIAS.n538 CS_BIAS.n462 24.4675
R9440 CS_BIAS.n534 CS_BIAS.n533 24.4675
R9441 CS_BIAS.n533 CS_BIAS.n532 24.4675
R9442 CS_BIAS.n532 CS_BIAS.n465 24.4675
R9443 CS_BIAS.n528 CS_BIAS.n465 24.4675
R9444 CS_BIAS.n526 CS_BIAS.n467 24.4675
R9445 CS_BIAS.n522 CS_BIAS.n467 24.4675
R9446 CS_BIAS.n522 CS_BIAS.n521 24.4675
R9447 CS_BIAS.n521 CS_BIAS.n520 24.4675
R9448 CS_BIAS.n517 CS_BIAS.n516 24.4675
R9449 CS_BIAS.n516 CS_BIAS.n515 24.4675
R9450 CS_BIAS.n515 CS_BIAS.n471 24.4675
R9451 CS_BIAS.n511 CS_BIAS.n471 24.4675
R9452 CS_BIAS.n505 CS_BIAS.n473 24.4675
R9453 CS_BIAS.n505 CS_BIAS.n504 24.4675
R9454 CS_BIAS.n504 CS_BIAS.n503 24.4675
R9455 CS_BIAS.n503 CS_BIAS.n475 24.4675
R9456 CS_BIAS.n499 CS_BIAS.n498 24.4675
R9457 CS_BIAS.n498 CS_BIAS.n497 24.4675
R9458 CS_BIAS.n497 CS_BIAS.n478 24.4675
R9459 CS_BIAS.n493 CS_BIAS.n478 24.4675
R9460 CS_BIAS.n491 CS_BIAS.n480 24.4675
R9461 CS_BIAS.n487 CS_BIAS.n480 24.4675
R9462 CS_BIAS.n487 CS_BIAS.n486 24.4675
R9463 CS_BIAS.n486 CS_BIAS.n485 24.4675
R9464 CS_BIAS.n440 CS_BIAS.n439 24.4675
R9465 CS_BIAS.n439 CS_BIAS.n438 24.4675
R9466 CS_BIAS.n438 CS_BIAS.n300 24.4675
R9467 CS_BIAS.n434 CS_BIAS.n300 24.4675
R9468 CS_BIAS.n432 CS_BIAS.n302 24.4675
R9469 CS_BIAS.n428 CS_BIAS.n302 24.4675
R9470 CS_BIAS.n428 CS_BIAS.n427 24.4675
R9471 CS_BIAS.n427 CS_BIAS.n426 24.4675
R9472 CS_BIAS.n423 CS_BIAS.n422 24.4675
R9473 CS_BIAS.n422 CS_BIAS.n421 24.4675
R9474 CS_BIAS.n421 CS_BIAS.n306 24.4675
R9475 CS_BIAS.n417 CS_BIAS.n306 24.4675
R9476 CS_BIAS.n415 CS_BIAS.n308 24.4675
R9477 CS_BIAS.n411 CS_BIAS.n308 24.4675
R9478 CS_BIAS.n411 CS_BIAS.n410 24.4675
R9479 CS_BIAS.n410 CS_BIAS.n409 24.4675
R9480 CS_BIAS.n406 CS_BIAS.n405 24.4675
R9481 CS_BIAS.n405 CS_BIAS.n404 24.4675
R9482 CS_BIAS.n404 CS_BIAS.n312 24.4675
R9483 CS_BIAS.n400 CS_BIAS.n312 24.4675
R9484 CS_BIAS.n394 CS_BIAS.n314 24.4675
R9485 CS_BIAS.n394 CS_BIAS.n393 24.4675
R9486 CS_BIAS.n393 CS_BIAS.n392 24.4675
R9487 CS_BIAS.n392 CS_BIAS.n316 24.4675
R9488 CS_BIAS.n388 CS_BIAS.n387 24.4675
R9489 CS_BIAS.n387 CS_BIAS.n386 24.4675
R9490 CS_BIAS.n386 CS_BIAS.n319 24.4675
R9491 CS_BIAS.n382 CS_BIAS.n319 24.4675
R9492 CS_BIAS.n380 CS_BIAS.n321 24.4675
R9493 CS_BIAS.n376 CS_BIAS.n321 24.4675
R9494 CS_BIAS.n376 CS_BIAS.n375 24.4675
R9495 CS_BIAS.n375 CS_BIAS.n374 24.4675
R9496 CS_BIAS.n371 CS_BIAS.n370 24.4675
R9497 CS_BIAS.n370 CS_BIAS.n369 24.4675
R9498 CS_BIAS.n369 CS_BIAS.n325 24.4675
R9499 CS_BIAS.n365 CS_BIAS.n325 24.4675
R9500 CS_BIAS.n359 CS_BIAS.n327 24.4675
R9501 CS_BIAS.n359 CS_BIAS.n358 24.4675
R9502 CS_BIAS.n358 CS_BIAS.n357 24.4675
R9503 CS_BIAS.n357 CS_BIAS.n329 24.4675
R9504 CS_BIAS.n353 CS_BIAS.n352 24.4675
R9505 CS_BIAS.n352 CS_BIAS.n351 24.4675
R9506 CS_BIAS.n351 CS_BIAS.n332 24.4675
R9507 CS_BIAS.n347 CS_BIAS.n332 24.4675
R9508 CS_BIAS.n345 CS_BIAS.n334 24.4675
R9509 CS_BIAS.n341 CS_BIAS.n334 24.4675
R9510 CS_BIAS.n341 CS_BIAS.n340 24.4675
R9511 CS_BIAS.n340 CS_BIAS.n339 24.4675
R9512 CS_BIAS.n164 CS_BIAS.n163 24.4675
R9513 CS_BIAS.n163 CS_BIAS.n162 24.4675
R9514 CS_BIAS.n162 CS_BIAS.n24 24.4675
R9515 CS_BIAS.n158 CS_BIAS.n24 24.4675
R9516 CS_BIAS.n156 CS_BIAS.n26 24.4675
R9517 CS_BIAS.n152 CS_BIAS.n26 24.4675
R9518 CS_BIAS.n152 CS_BIAS.n151 24.4675
R9519 CS_BIAS.n151 CS_BIAS.n150 24.4675
R9520 CS_BIAS.n147 CS_BIAS.n146 24.4675
R9521 CS_BIAS.n146 CS_BIAS.n145 24.4675
R9522 CS_BIAS.n145 CS_BIAS.n30 24.4675
R9523 CS_BIAS.n141 CS_BIAS.n30 24.4675
R9524 CS_BIAS.n139 CS_BIAS.n32 24.4675
R9525 CS_BIAS.n135 CS_BIAS.n32 24.4675
R9526 CS_BIAS.n135 CS_BIAS.n134 24.4675
R9527 CS_BIAS.n134 CS_BIAS.n133 24.4675
R9528 CS_BIAS.n130 CS_BIAS.n129 24.4675
R9529 CS_BIAS.n129 CS_BIAS.n128 24.4675
R9530 CS_BIAS.n128 CS_BIAS.n36 24.4675
R9531 CS_BIAS.n124 CS_BIAS.n36 24.4675
R9532 CS_BIAS.n118 CS_BIAS.n38 24.4675
R9533 CS_BIAS.n118 CS_BIAS.n117 24.4675
R9534 CS_BIAS.n117 CS_BIAS.n116 24.4675
R9535 CS_BIAS.n116 CS_BIAS.n40 24.4675
R9536 CS_BIAS.n112 CS_BIAS.n111 24.4675
R9537 CS_BIAS.n111 CS_BIAS.n110 24.4675
R9538 CS_BIAS.n110 CS_BIAS.n43 24.4675
R9539 CS_BIAS.n106 CS_BIAS.n43 24.4675
R9540 CS_BIAS.n104 CS_BIAS.n45 24.4675
R9541 CS_BIAS.n100 CS_BIAS.n45 24.4675
R9542 CS_BIAS.n100 CS_BIAS.n99 24.4675
R9543 CS_BIAS.n99 CS_BIAS.n98 24.4675
R9544 CS_BIAS.n95 CS_BIAS.n94 24.4675
R9545 CS_BIAS.n94 CS_BIAS.n93 24.4675
R9546 CS_BIAS.n93 CS_BIAS.n49 24.4675
R9547 CS_BIAS.n89 CS_BIAS.n49 24.4675
R9548 CS_BIAS.n83 CS_BIAS.n51 24.4675
R9549 CS_BIAS.n83 CS_BIAS.n82 24.4675
R9550 CS_BIAS.n82 CS_BIAS.n81 24.4675
R9551 CS_BIAS.n81 CS_BIAS.n53 24.4675
R9552 CS_BIAS.n77 CS_BIAS.n76 24.4675
R9553 CS_BIAS.n76 CS_BIAS.n75 24.4675
R9554 CS_BIAS.n75 CS_BIAS.n56 24.4675
R9555 CS_BIAS.n71 CS_BIAS.n56 24.4675
R9556 CS_BIAS.n69 CS_BIAS.n58 24.4675
R9557 CS_BIAS.n65 CS_BIAS.n58 24.4675
R9558 CS_BIAS.n65 CS_BIAS.n64 24.4675
R9559 CS_BIAS.n64 CS_BIAS.n63 24.4675
R9560 CS_BIAS.n295 CS_BIAS.n294 24.4675
R9561 CS_BIAS.n294 CS_BIAS.n293 24.4675
R9562 CS_BIAS.n293 CS_BIAS.n2 24.4675
R9563 CS_BIAS.n289 CS_BIAS.n2 24.4675
R9564 CS_BIAS.n287 CS_BIAS.n4 24.4675
R9565 CS_BIAS.n283 CS_BIAS.n4 24.4675
R9566 CS_BIAS.n283 CS_BIAS.n282 24.4675
R9567 CS_BIAS.n282 CS_BIAS.n281 24.4675
R9568 CS_BIAS.n278 CS_BIAS.n277 24.4675
R9569 CS_BIAS.n277 CS_BIAS.n276 24.4675
R9570 CS_BIAS.n276 CS_BIAS.n8 24.4675
R9571 CS_BIAS.n272 CS_BIAS.n8 24.4675
R9572 CS_BIAS.n270 CS_BIAS.n10 24.4675
R9573 CS_BIAS.n266 CS_BIAS.n10 24.4675
R9574 CS_BIAS.n266 CS_BIAS.n265 24.4675
R9575 CS_BIAS.n265 CS_BIAS.n264 24.4675
R9576 CS_BIAS.n261 CS_BIAS.n260 24.4675
R9577 CS_BIAS.n260 CS_BIAS.n259 24.4675
R9578 CS_BIAS.n259 CS_BIAS.n14 24.4675
R9579 CS_BIAS.n255 CS_BIAS.n14 24.4675
R9580 CS_BIAS.n249 CS_BIAS.n16 24.4675
R9581 CS_BIAS.n249 CS_BIAS.n248 24.4675
R9582 CS_BIAS.n248 CS_BIAS.n247 24.4675
R9583 CS_BIAS.n247 CS_BIAS.n18 24.4675
R9584 CS_BIAS.n243 CS_BIAS.n242 24.4675
R9585 CS_BIAS.n242 CS_BIAS.n241 24.4675
R9586 CS_BIAS.n241 CS_BIAS.n21 24.4675
R9587 CS_BIAS.n237 CS_BIAS.n21 24.4675
R9588 CS_BIAS.n235 CS_BIAS.n176 24.4675
R9589 CS_BIAS.n231 CS_BIAS.n176 24.4675
R9590 CS_BIAS.n231 CS_BIAS.n230 24.4675
R9591 CS_BIAS.n230 CS_BIAS.n229 24.4675
R9592 CS_BIAS.n226 CS_BIAS.n225 24.4675
R9593 CS_BIAS.n225 CS_BIAS.n224 24.4675
R9594 CS_BIAS.n224 CS_BIAS.n180 24.4675
R9595 CS_BIAS.n220 CS_BIAS.n180 24.4675
R9596 CS_BIAS.n214 CS_BIAS.n182 24.4675
R9597 CS_BIAS.n214 CS_BIAS.n213 24.4675
R9598 CS_BIAS.n213 CS_BIAS.n212 24.4675
R9599 CS_BIAS.n212 CS_BIAS.n184 24.4675
R9600 CS_BIAS.n208 CS_BIAS.n207 24.4675
R9601 CS_BIAS.n207 CS_BIAS.n206 24.4675
R9602 CS_BIAS.n206 CS_BIAS.n187 24.4675
R9603 CS_BIAS.n202 CS_BIAS.n187 24.4675
R9604 CS_BIAS.n200 CS_BIAS.n189 24.4675
R9605 CS_BIAS.n196 CS_BIAS.n189 24.4675
R9606 CS_BIAS.n196 CS_BIAS.n195 24.4675
R9607 CS_BIAS.n195 CS_BIAS.n194 24.4675
R9608 CS_BIAS.n1658 CS_BIAS.n1657 24.4675
R9609 CS_BIAS.n1659 CS_BIAS.n1658 24.4675
R9610 CS_BIAS.n1659 CS_BIAS.n1652 24.4675
R9611 CS_BIAS.n1663 CS_BIAS.n1652 24.4675
R9612 CS_BIAS.n1665 CS_BIAS.n1650 24.4675
R9613 CS_BIAS.n1669 CS_BIAS.n1650 24.4675
R9614 CS_BIAS.n1670 CS_BIAS.n1669 24.4675
R9615 CS_BIAS.n1672 CS_BIAS.n1670 24.4675
R9616 CS_BIAS.n1676 CS_BIAS.n1648 24.4675
R9617 CS_BIAS.n1677 CS_BIAS.n1676 24.4675
R9618 CS_BIAS.n1678 CS_BIAS.n1677 24.4675
R9619 CS_BIAS.n1678 CS_BIAS.n1646 24.4675
R9620 CS_BIAS.n1684 CS_BIAS.n1644 24.4675
R9621 CS_BIAS.n1688 CS_BIAS.n1644 24.4675
R9622 CS_BIAS.n1689 CS_BIAS.n1688 24.4675
R9623 CS_BIAS.n1690 CS_BIAS.n1689 24.4675
R9624 CS_BIAS.n1694 CS_BIAS.n1693 24.4675
R9625 CS_BIAS.n1695 CS_BIAS.n1694 24.4675
R9626 CS_BIAS.n1695 CS_BIAS.n1640 24.4675
R9627 CS_BIAS.n1699 CS_BIAS.n1640 24.4675
R9628 CS_BIAS.n1701 CS_BIAS.n1638 24.4675
R9629 CS_BIAS.n1705 CS_BIAS.n1638 24.4675
R9630 CS_BIAS.n1706 CS_BIAS.n1705 24.4675
R9631 CS_BIAS.n1708 CS_BIAS.n1706 24.4675
R9632 CS_BIAS.n1712 CS_BIAS.n1636 24.4675
R9633 CS_BIAS.n1713 CS_BIAS.n1712 24.4675
R9634 CS_BIAS.n1714 CS_BIAS.n1713 24.4675
R9635 CS_BIAS.n1714 CS_BIAS.n1634 24.4675
R9636 CS_BIAS.n1720 CS_BIAS.n1632 24.4675
R9637 CS_BIAS.n1724 CS_BIAS.n1632 24.4675
R9638 CS_BIAS.n1725 CS_BIAS.n1724 24.4675
R9639 CS_BIAS.n1726 CS_BIAS.n1725 24.4675
R9640 CS_BIAS.n1730 CS_BIAS.n1729 24.4675
R9641 CS_BIAS.n1731 CS_BIAS.n1730 24.4675
R9642 CS_BIAS.n1731 CS_BIAS.n1628 24.4675
R9643 CS_BIAS.n1735 CS_BIAS.n1628 24.4675
R9644 CS_BIAS.n1737 CS_BIAS.n1626 24.4675
R9645 CS_BIAS.n1741 CS_BIAS.n1626 24.4675
R9646 CS_BIAS.n1742 CS_BIAS.n1741 24.4675
R9647 CS_BIAS.n1743 CS_BIAS.n1742 24.4675
R9648 CS_BIAS.n1747 CS_BIAS.n1746 24.4675
R9649 CS_BIAS.n1748 CS_BIAS.n1747 24.4675
R9650 CS_BIAS.n1748 CS_BIAS.n1622 24.4675
R9651 CS_BIAS.n1752 CS_BIAS.n1622 24.4675
R9652 CS_BIAS.n1754 CS_BIAS.n1620 24.4675
R9653 CS_BIAS.n1758 CS_BIAS.n1620 24.4675
R9654 CS_BIAS.n1759 CS_BIAS.n1758 24.4675
R9655 CS_BIAS.n1760 CS_BIAS.n1759 24.4675
R9656 CS_BIAS.n1512 CS_BIAS.n1511 24.4675
R9657 CS_BIAS.n1513 CS_BIAS.n1512 24.4675
R9658 CS_BIAS.n1513 CS_BIAS.n1506 24.4675
R9659 CS_BIAS.n1517 CS_BIAS.n1506 24.4675
R9660 CS_BIAS.n1519 CS_BIAS.n1504 24.4675
R9661 CS_BIAS.n1523 CS_BIAS.n1504 24.4675
R9662 CS_BIAS.n1524 CS_BIAS.n1523 24.4675
R9663 CS_BIAS.n1526 CS_BIAS.n1524 24.4675
R9664 CS_BIAS.n1530 CS_BIAS.n1502 24.4675
R9665 CS_BIAS.n1531 CS_BIAS.n1530 24.4675
R9666 CS_BIAS.n1532 CS_BIAS.n1531 24.4675
R9667 CS_BIAS.n1532 CS_BIAS.n1500 24.4675
R9668 CS_BIAS.n1538 CS_BIAS.n1498 24.4675
R9669 CS_BIAS.n1542 CS_BIAS.n1498 24.4675
R9670 CS_BIAS.n1543 CS_BIAS.n1542 24.4675
R9671 CS_BIAS.n1544 CS_BIAS.n1543 24.4675
R9672 CS_BIAS.n1548 CS_BIAS.n1547 24.4675
R9673 CS_BIAS.n1549 CS_BIAS.n1548 24.4675
R9674 CS_BIAS.n1549 CS_BIAS.n1494 24.4675
R9675 CS_BIAS.n1553 CS_BIAS.n1494 24.4675
R9676 CS_BIAS.n1555 CS_BIAS.n1492 24.4675
R9677 CS_BIAS.n1559 CS_BIAS.n1492 24.4675
R9678 CS_BIAS.n1560 CS_BIAS.n1559 24.4675
R9679 CS_BIAS.n1562 CS_BIAS.n1560 24.4675
R9680 CS_BIAS.n1566 CS_BIAS.n1490 24.4675
R9681 CS_BIAS.n1567 CS_BIAS.n1566 24.4675
R9682 CS_BIAS.n1568 CS_BIAS.n1567 24.4675
R9683 CS_BIAS.n1568 CS_BIAS.n1488 24.4675
R9684 CS_BIAS.n1574 CS_BIAS.n1486 24.4675
R9685 CS_BIAS.n1578 CS_BIAS.n1486 24.4675
R9686 CS_BIAS.n1579 CS_BIAS.n1578 24.4675
R9687 CS_BIAS.n1580 CS_BIAS.n1579 24.4675
R9688 CS_BIAS.n1584 CS_BIAS.n1583 24.4675
R9689 CS_BIAS.n1585 CS_BIAS.n1584 24.4675
R9690 CS_BIAS.n1585 CS_BIAS.n1482 24.4675
R9691 CS_BIAS.n1589 CS_BIAS.n1482 24.4675
R9692 CS_BIAS.n1591 CS_BIAS.n1480 24.4675
R9693 CS_BIAS.n1595 CS_BIAS.n1480 24.4675
R9694 CS_BIAS.n1596 CS_BIAS.n1595 24.4675
R9695 CS_BIAS.n1597 CS_BIAS.n1596 24.4675
R9696 CS_BIAS.n1601 CS_BIAS.n1600 24.4675
R9697 CS_BIAS.n1602 CS_BIAS.n1601 24.4675
R9698 CS_BIAS.n1602 CS_BIAS.n1476 24.4675
R9699 CS_BIAS.n1606 CS_BIAS.n1476 24.4675
R9700 CS_BIAS.n1608 CS_BIAS.n1474 24.4675
R9701 CS_BIAS.n1612 CS_BIAS.n1474 24.4675
R9702 CS_BIAS.n1613 CS_BIAS.n1612 24.4675
R9703 CS_BIAS.n1614 CS_BIAS.n1613 24.4675
R9704 CS_BIAS.n1366 CS_BIAS.n1365 24.4675
R9705 CS_BIAS.n1367 CS_BIAS.n1366 24.4675
R9706 CS_BIAS.n1367 CS_BIAS.n1360 24.4675
R9707 CS_BIAS.n1371 CS_BIAS.n1360 24.4675
R9708 CS_BIAS.n1373 CS_BIAS.n1358 24.4675
R9709 CS_BIAS.n1377 CS_BIAS.n1358 24.4675
R9710 CS_BIAS.n1378 CS_BIAS.n1377 24.4675
R9711 CS_BIAS.n1380 CS_BIAS.n1378 24.4675
R9712 CS_BIAS.n1384 CS_BIAS.n1356 24.4675
R9713 CS_BIAS.n1385 CS_BIAS.n1384 24.4675
R9714 CS_BIAS.n1386 CS_BIAS.n1385 24.4675
R9715 CS_BIAS.n1386 CS_BIAS.n1354 24.4675
R9716 CS_BIAS.n1392 CS_BIAS.n1352 24.4675
R9717 CS_BIAS.n1396 CS_BIAS.n1352 24.4675
R9718 CS_BIAS.n1397 CS_BIAS.n1396 24.4675
R9719 CS_BIAS.n1398 CS_BIAS.n1397 24.4675
R9720 CS_BIAS.n1402 CS_BIAS.n1401 24.4675
R9721 CS_BIAS.n1403 CS_BIAS.n1402 24.4675
R9722 CS_BIAS.n1403 CS_BIAS.n1348 24.4675
R9723 CS_BIAS.n1407 CS_BIAS.n1348 24.4675
R9724 CS_BIAS.n1409 CS_BIAS.n1346 24.4675
R9725 CS_BIAS.n1413 CS_BIAS.n1346 24.4675
R9726 CS_BIAS.n1414 CS_BIAS.n1413 24.4675
R9727 CS_BIAS.n1416 CS_BIAS.n1414 24.4675
R9728 CS_BIAS.n1420 CS_BIAS.n1344 24.4675
R9729 CS_BIAS.n1421 CS_BIAS.n1420 24.4675
R9730 CS_BIAS.n1422 CS_BIAS.n1421 24.4675
R9731 CS_BIAS.n1422 CS_BIAS.n1342 24.4675
R9732 CS_BIAS.n1428 CS_BIAS.n1340 24.4675
R9733 CS_BIAS.n1432 CS_BIAS.n1340 24.4675
R9734 CS_BIAS.n1433 CS_BIAS.n1432 24.4675
R9735 CS_BIAS.n1434 CS_BIAS.n1433 24.4675
R9736 CS_BIAS.n1438 CS_BIAS.n1437 24.4675
R9737 CS_BIAS.n1439 CS_BIAS.n1438 24.4675
R9738 CS_BIAS.n1439 CS_BIAS.n1336 24.4675
R9739 CS_BIAS.n1443 CS_BIAS.n1336 24.4675
R9740 CS_BIAS.n1445 CS_BIAS.n1334 24.4675
R9741 CS_BIAS.n1449 CS_BIAS.n1334 24.4675
R9742 CS_BIAS.n1450 CS_BIAS.n1449 24.4675
R9743 CS_BIAS.n1451 CS_BIAS.n1450 24.4675
R9744 CS_BIAS.n1455 CS_BIAS.n1454 24.4675
R9745 CS_BIAS.n1456 CS_BIAS.n1455 24.4675
R9746 CS_BIAS.n1456 CS_BIAS.n1330 24.4675
R9747 CS_BIAS.n1460 CS_BIAS.n1330 24.4675
R9748 CS_BIAS.n1462 CS_BIAS.n1328 24.4675
R9749 CS_BIAS.n1466 CS_BIAS.n1328 24.4675
R9750 CS_BIAS.n1467 CS_BIAS.n1466 24.4675
R9751 CS_BIAS.n1468 CS_BIAS.n1467 24.4675
R9752 CS_BIAS.n1220 CS_BIAS.n1219 24.4675
R9753 CS_BIAS.n1221 CS_BIAS.n1220 24.4675
R9754 CS_BIAS.n1221 CS_BIAS.n1214 24.4675
R9755 CS_BIAS.n1225 CS_BIAS.n1214 24.4675
R9756 CS_BIAS.n1227 CS_BIAS.n1212 24.4675
R9757 CS_BIAS.n1231 CS_BIAS.n1212 24.4675
R9758 CS_BIAS.n1232 CS_BIAS.n1231 24.4675
R9759 CS_BIAS.n1234 CS_BIAS.n1232 24.4675
R9760 CS_BIAS.n1238 CS_BIAS.n1210 24.4675
R9761 CS_BIAS.n1239 CS_BIAS.n1238 24.4675
R9762 CS_BIAS.n1240 CS_BIAS.n1239 24.4675
R9763 CS_BIAS.n1240 CS_BIAS.n1208 24.4675
R9764 CS_BIAS.n1246 CS_BIAS.n1206 24.4675
R9765 CS_BIAS.n1250 CS_BIAS.n1206 24.4675
R9766 CS_BIAS.n1251 CS_BIAS.n1250 24.4675
R9767 CS_BIAS.n1252 CS_BIAS.n1251 24.4675
R9768 CS_BIAS.n1256 CS_BIAS.n1255 24.4675
R9769 CS_BIAS.n1257 CS_BIAS.n1256 24.4675
R9770 CS_BIAS.n1257 CS_BIAS.n1202 24.4675
R9771 CS_BIAS.n1261 CS_BIAS.n1202 24.4675
R9772 CS_BIAS.n1263 CS_BIAS.n1200 24.4675
R9773 CS_BIAS.n1267 CS_BIAS.n1200 24.4675
R9774 CS_BIAS.n1268 CS_BIAS.n1267 24.4675
R9775 CS_BIAS.n1270 CS_BIAS.n1268 24.4675
R9776 CS_BIAS.n1274 CS_BIAS.n1198 24.4675
R9777 CS_BIAS.n1275 CS_BIAS.n1274 24.4675
R9778 CS_BIAS.n1276 CS_BIAS.n1275 24.4675
R9779 CS_BIAS.n1276 CS_BIAS.n1196 24.4675
R9780 CS_BIAS.n1282 CS_BIAS.n1194 24.4675
R9781 CS_BIAS.n1286 CS_BIAS.n1194 24.4675
R9782 CS_BIAS.n1287 CS_BIAS.n1286 24.4675
R9783 CS_BIAS.n1288 CS_BIAS.n1287 24.4675
R9784 CS_BIAS.n1292 CS_BIAS.n1291 24.4675
R9785 CS_BIAS.n1293 CS_BIAS.n1292 24.4675
R9786 CS_BIAS.n1293 CS_BIAS.n1190 24.4675
R9787 CS_BIAS.n1297 CS_BIAS.n1190 24.4675
R9788 CS_BIAS.n1299 CS_BIAS.n1188 24.4675
R9789 CS_BIAS.n1303 CS_BIAS.n1188 24.4675
R9790 CS_BIAS.n1304 CS_BIAS.n1303 24.4675
R9791 CS_BIAS.n1305 CS_BIAS.n1304 24.4675
R9792 CS_BIAS.n1309 CS_BIAS.n1308 24.4675
R9793 CS_BIAS.n1310 CS_BIAS.n1309 24.4675
R9794 CS_BIAS.n1310 CS_BIAS.n1184 24.4675
R9795 CS_BIAS.n1314 CS_BIAS.n1184 24.4675
R9796 CS_BIAS.n1316 CS_BIAS.n1182 24.4675
R9797 CS_BIAS.n1320 CS_BIAS.n1182 24.4675
R9798 CS_BIAS.n1321 CS_BIAS.n1320 24.4675
R9799 CS_BIAS.n1322 CS_BIAS.n1321 24.4675
R9800 CS_BIAS.n946 CS_BIAS.n945 24.4675
R9801 CS_BIAS.n947 CS_BIAS.n946 24.4675
R9802 CS_BIAS.n947 CS_BIAS.n940 24.4675
R9803 CS_BIAS.n951 CS_BIAS.n940 24.4675
R9804 CS_BIAS.n953 CS_BIAS.n938 24.4675
R9805 CS_BIAS.n957 CS_BIAS.n938 24.4675
R9806 CS_BIAS.n958 CS_BIAS.n957 24.4675
R9807 CS_BIAS.n960 CS_BIAS.n958 24.4675
R9808 CS_BIAS.n964 CS_BIAS.n936 24.4675
R9809 CS_BIAS.n965 CS_BIAS.n964 24.4675
R9810 CS_BIAS.n966 CS_BIAS.n965 24.4675
R9811 CS_BIAS.n966 CS_BIAS.n934 24.4675
R9812 CS_BIAS.n972 CS_BIAS.n932 24.4675
R9813 CS_BIAS.n976 CS_BIAS.n932 24.4675
R9814 CS_BIAS.n977 CS_BIAS.n976 24.4675
R9815 CS_BIAS.n978 CS_BIAS.n977 24.4675
R9816 CS_BIAS.n982 CS_BIAS.n981 24.4675
R9817 CS_BIAS.n983 CS_BIAS.n982 24.4675
R9818 CS_BIAS.n983 CS_BIAS.n928 24.4675
R9819 CS_BIAS.n987 CS_BIAS.n928 24.4675
R9820 CS_BIAS.n989 CS_BIAS.n926 24.4675
R9821 CS_BIAS.n993 CS_BIAS.n926 24.4675
R9822 CS_BIAS.n994 CS_BIAS.n993 24.4675
R9823 CS_BIAS.n996 CS_BIAS.n994 24.4675
R9824 CS_BIAS.n1000 CS_BIAS.n924 24.4675
R9825 CS_BIAS.n1001 CS_BIAS.n1000 24.4675
R9826 CS_BIAS.n1002 CS_BIAS.n1001 24.4675
R9827 CS_BIAS.n1002 CS_BIAS.n922 24.4675
R9828 CS_BIAS.n1008 CS_BIAS.n920 24.4675
R9829 CS_BIAS.n1012 CS_BIAS.n920 24.4675
R9830 CS_BIAS.n1013 CS_BIAS.n1012 24.4675
R9831 CS_BIAS.n1014 CS_BIAS.n1013 24.4675
R9832 CS_BIAS.n1018 CS_BIAS.n1017 24.4675
R9833 CS_BIAS.n1019 CS_BIAS.n1018 24.4675
R9834 CS_BIAS.n1019 CS_BIAS.n916 24.4675
R9835 CS_BIAS.n1023 CS_BIAS.n916 24.4675
R9836 CS_BIAS.n1025 CS_BIAS.n914 24.4675
R9837 CS_BIAS.n1029 CS_BIAS.n914 24.4675
R9838 CS_BIAS.n1030 CS_BIAS.n1029 24.4675
R9839 CS_BIAS.n1031 CS_BIAS.n1030 24.4675
R9840 CS_BIAS.n1035 CS_BIAS.n1034 24.4675
R9841 CS_BIAS.n1036 CS_BIAS.n1035 24.4675
R9842 CS_BIAS.n1036 CS_BIAS.n910 24.4675
R9843 CS_BIAS.n1040 CS_BIAS.n910 24.4675
R9844 CS_BIAS.n1042 CS_BIAS.n908 24.4675
R9845 CS_BIAS.n1046 CS_BIAS.n908 24.4675
R9846 CS_BIAS.n1047 CS_BIAS.n1046 24.4675
R9847 CS_BIAS.n1048 CS_BIAS.n1047 24.4675
R9848 CS_BIAS.n1171 CS_BIAS.n884 24.4675
R9849 CS_BIAS.n1175 CS_BIAS.n884 24.4675
R9850 CS_BIAS.n1176 CS_BIAS.n1175 24.4675
R9851 CS_BIAS.n1177 CS_BIAS.n1176 24.4675
R9852 CS_BIAS.n1154 CS_BIAS.n890 24.4675
R9853 CS_BIAS.n1158 CS_BIAS.n890 24.4675
R9854 CS_BIAS.n1159 CS_BIAS.n1158 24.4675
R9855 CS_BIAS.n1160 CS_BIAS.n1159 24.4675
R9856 CS_BIAS.n1164 CS_BIAS.n1163 24.4675
R9857 CS_BIAS.n1165 CS_BIAS.n1164 24.4675
R9858 CS_BIAS.n1165 CS_BIAS.n886 24.4675
R9859 CS_BIAS.n1169 CS_BIAS.n886 24.4675
R9860 CS_BIAS.n1137 CS_BIAS.n896 24.4675
R9861 CS_BIAS.n1141 CS_BIAS.n896 24.4675
R9862 CS_BIAS.n1142 CS_BIAS.n1141 24.4675
R9863 CS_BIAS.n1143 CS_BIAS.n1142 24.4675
R9864 CS_BIAS.n1147 CS_BIAS.n1146 24.4675
R9865 CS_BIAS.n1148 CS_BIAS.n1147 24.4675
R9866 CS_BIAS.n1148 CS_BIAS.n892 24.4675
R9867 CS_BIAS.n1152 CS_BIAS.n892 24.4675
R9868 CS_BIAS.n1118 CS_BIAS.n902 24.4675
R9869 CS_BIAS.n1122 CS_BIAS.n902 24.4675
R9870 CS_BIAS.n1123 CS_BIAS.n1122 24.4675
R9871 CS_BIAS.n1125 CS_BIAS.n1123 24.4675
R9872 CS_BIAS.n1129 CS_BIAS.n900 24.4675
R9873 CS_BIAS.n1130 CS_BIAS.n1129 24.4675
R9874 CS_BIAS.n1131 CS_BIAS.n1130 24.4675
R9875 CS_BIAS.n1131 CS_BIAS.n898 24.4675
R9876 CS_BIAS.n1075 CS_BIAS.n1074 24.4675
R9877 CS_BIAS.n1076 CS_BIAS.n1075 24.4675
R9878 CS_BIAS.n1076 CS_BIAS.n1069 24.4675
R9879 CS_BIAS.n1080 CS_BIAS.n1069 24.4675
R9880 CS_BIAS.n1082 CS_BIAS.n1067 24.4675
R9881 CS_BIAS.n1086 CS_BIAS.n1067 24.4675
R9882 CS_BIAS.n1087 CS_BIAS.n1086 24.4675
R9883 CS_BIAS.n1089 CS_BIAS.n1087 24.4675
R9884 CS_BIAS.n1093 CS_BIAS.n1065 24.4675
R9885 CS_BIAS.n1094 CS_BIAS.n1093 24.4675
R9886 CS_BIAS.n1095 CS_BIAS.n1094 24.4675
R9887 CS_BIAS.n1095 CS_BIAS.n1063 24.4675
R9888 CS_BIAS.n1101 CS_BIAS.n1061 24.4675
R9889 CS_BIAS.n1105 CS_BIAS.n1061 24.4675
R9890 CS_BIAS.n1106 CS_BIAS.n1105 24.4675
R9891 CS_BIAS.n1107 CS_BIAS.n1106 24.4675
R9892 CS_BIAS.n1111 CS_BIAS.n1110 24.4675
R9893 CS_BIAS.n1112 CS_BIAS.n1111 24.4675
R9894 CS_BIAS.n1112 CS_BIAS.n1057 24.4675
R9895 CS_BIAS.n1116 CS_BIAS.n1057 24.4675
R9896 CS_BIAS.n791 CS_BIAS.n769 22.7548
R9897 CS_BIAS.n847 CS_BIAS.n748 22.7548
R9898 CS_BIAS.n701 CS_BIAS.n602 22.7548
R9899 CS_BIAS.n645 CS_BIAS.n623 22.7548
R9900 CS_BIAS.n555 CS_BIAS.n456 22.7548
R9901 CS_BIAS.n499 CS_BIAS.n477 22.7548
R9902 CS_BIAS.n409 CS_BIAS.n310 22.7548
R9903 CS_BIAS.n353 CS_BIAS.n331 22.7548
R9904 CS_BIAS.n133 CS_BIAS.n34 22.7548
R9905 CS_BIAS.n77 CS_BIAS.n55 22.7548
R9906 CS_BIAS.n264 CS_BIAS.n12 22.7548
R9907 CS_BIAS.n208 CS_BIAS.n186 22.7548
R9908 CS_BIAS.n1672 CS_BIAS.n1671 22.7548
R9909 CS_BIAS.n1729 CS_BIAS.n1630 22.7548
R9910 CS_BIAS.n1526 CS_BIAS.n1525 22.7548
R9911 CS_BIAS.n1583 CS_BIAS.n1484 22.7548
R9912 CS_BIAS.n1380 CS_BIAS.n1379 22.7548
R9913 CS_BIAS.n1437 CS_BIAS.n1338 22.7548
R9914 CS_BIAS.n1234 CS_BIAS.n1233 22.7548
R9915 CS_BIAS.n1291 CS_BIAS.n1192 22.7548
R9916 CS_BIAS.n960 CS_BIAS.n959 22.7548
R9917 CS_BIAS.n1017 CS_BIAS.n918 22.7548
R9918 CS_BIAS.n1146 CS_BIAS.n894 22.7548
R9919 CS_BIAS.n1089 CS_BIAS.n1088 22.7548
R9920 CS_BIAS.n878 CS_BIAS.n736 20.3081
R9921 CS_BIAS.n732 CS_BIAS.n590 20.3081
R9922 CS_BIAS.n586 CS_BIAS.n444 20.3081
R9923 CS_BIAS.n440 CS_BIAS.n298 20.3081
R9924 CS_BIAS.n164 CS_BIAS.n22 20.3081
R9925 CS_BIAS.n295 CS_BIAS.n0 20.3081
R9926 CS_BIAS.n1760 CS_BIAS.n1618 20.3081
R9927 CS_BIAS.n1614 CS_BIAS.n1472 20.3081
R9928 CS_BIAS.n1468 CS_BIAS.n1326 20.3081
R9929 CS_BIAS.n1322 CS_BIAS.n1180 20.3081
R9930 CS_BIAS.n1048 CS_BIAS.n906 20.3081
R9931 CS_BIAS.n1177 CS_BIAS.n882 20.3081
R9932 CS_BIAS.n812 CS_BIAS.n761 16.8827
R9933 CS_BIAS.n826 CS_BIAS.n756 16.8827
R9934 CS_BIAS.n680 CS_BIAS.n610 16.8827
R9935 CS_BIAS.n666 CS_BIAS.n615 16.8827
R9936 CS_BIAS.n534 CS_BIAS.n464 16.8827
R9937 CS_BIAS.n520 CS_BIAS.n469 16.8827
R9938 CS_BIAS.n388 CS_BIAS.n318 16.8827
R9939 CS_BIAS.n374 CS_BIAS.n323 16.8827
R9940 CS_BIAS.n112 CS_BIAS.n42 16.8827
R9941 CS_BIAS.n98 CS_BIAS.n47 16.8827
R9942 CS_BIAS.n243 CS_BIAS.n20 16.8827
R9943 CS_BIAS.n229 CS_BIAS.n178 16.8827
R9944 CS_BIAS.n1693 CS_BIAS.n1642 16.8827
R9945 CS_BIAS.n1708 CS_BIAS.n1707 16.8827
R9946 CS_BIAS.n1547 CS_BIAS.n1496 16.8827
R9947 CS_BIAS.n1562 CS_BIAS.n1561 16.8827
R9948 CS_BIAS.n1401 CS_BIAS.n1350 16.8827
R9949 CS_BIAS.n1416 CS_BIAS.n1415 16.8827
R9950 CS_BIAS.n1255 CS_BIAS.n1204 16.8827
R9951 CS_BIAS.n1270 CS_BIAS.n1269 16.8827
R9952 CS_BIAS.n981 CS_BIAS.n930 16.8827
R9953 CS_BIAS.n996 CS_BIAS.n995 16.8827
R9954 CS_BIAS.n1125 CS_BIAS.n1124 16.8827
R9955 CS_BIAS.n1110 CS_BIAS.n1059 16.8827
R9956 CS_BIAS.n171 CS_BIAS.t15 14.194
R9957 CS_BIAS.n171 CS_BIAS.t19 14.194
R9958 CS_BIAS.n172 CS_BIAS.t21 14.194
R9959 CS_BIAS.n172 CS_BIAS.t9 14.194
R9960 CS_BIAS.n169 CS_BIAS.t23 14.194
R9961 CS_BIAS.n169 CS_BIAS.t17 14.194
R9962 CS_BIAS.n167 CS_BIAS.t1 14.194
R9963 CS_BIAS.n167 CS_BIAS.t27 14.194
R9964 CS_BIAS.n1051 CS_BIAS.t3 14.194
R9965 CS_BIAS.n1051 CS_BIAS.t7 14.194
R9966 CS_BIAS.n1053 CS_BIAS.t13 14.194
R9967 CS_BIAS.n1053 CS_BIAS.t29 14.194
R9968 CS_BIAS.n904 CS_BIAS.t25 14.194
R9969 CS_BIAS.n904 CS_BIAS.t5 14.194
R9970 CS_BIAS.n903 CS_BIAS.t31 14.194
R9971 CS_BIAS.n903 CS_BIAS.t11 14.194
R9972 CS_BIAS.n864 CS_BIAS.n742 13.4574
R9973 CS_BIAS.n718 CS_BIAS.n596 13.4574
R9974 CS_BIAS.n572 CS_BIAS.n450 13.4574
R9975 CS_BIAS.n426 CS_BIAS.n304 13.4574
R9976 CS_BIAS.n150 CS_BIAS.n28 13.4574
R9977 CS_BIAS.n281 CS_BIAS.n6 13.4574
R9978 CS_BIAS.n1746 CS_BIAS.n1624 13.4574
R9979 CS_BIAS.n1600 CS_BIAS.n1478 13.4574
R9980 CS_BIAS.n1454 CS_BIAS.n1332 13.4574
R9981 CS_BIAS.n1308 CS_BIAS.n1186 13.4574
R9982 CS_BIAS.n1034 CS_BIAS.n912 13.4574
R9983 CS_BIAS.n1163 CS_BIAS.n888 13.4574
R9984 CS_BIAS.n774 CS_BIAS.t109 13.3681
R9985 CS_BIAS.n769 CS_BIAS.t54 13.3681
R9986 CS_BIAS.n761 CS_BIAS.t43 13.3681
R9987 CS_BIAS.n756 CS_BIAS.t46 13.3681
R9988 CS_BIAS.n748 CS_BIAS.t48 13.3681
R9989 CS_BIAS.n742 CS_BIAS.t76 13.3681
R9990 CS_BIAS.n736 CS_BIAS.t99 13.3681
R9991 CS_BIAS.n590 CS_BIAS.t56 13.3681
R9992 CS_BIAS.n596 CS_BIAS.t111 13.3681
R9993 CS_BIAS.n602 CS_BIAS.t96 13.3681
R9994 CS_BIAS.n610 CS_BIAS.t93 13.3681
R9995 CS_BIAS.n615 CS_BIAS.t89 13.3681
R9996 CS_BIAS.n623 CS_BIAS.t100 13.3681
R9997 CS_BIAS.n628 CS_BIAS.t77 13.3681
R9998 CS_BIAS.n444 CS_BIAS.t50 13.3681
R9999 CS_BIAS.n450 CS_BIAS.t59 13.3681
R10000 CS_BIAS.n456 CS_BIAS.t86 13.3681
R10001 CS_BIAS.n464 CS_BIAS.t98 13.3681
R10002 CS_BIAS.n469 CS_BIAS.t102 13.3681
R10003 CS_BIAS.n477 CS_BIAS.t104 13.3681
R10004 CS_BIAS.n482 CS_BIAS.t33 13.3681
R10005 CS_BIAS.n298 CS_BIAS.t32 13.3681
R10006 CS_BIAS.n304 CS_BIAS.t97 13.3681
R10007 CS_BIAS.n310 CS_BIAS.t74 13.3681
R10008 CS_BIAS.n318 CS_BIAS.t72 13.3681
R10009 CS_BIAS.n323 CS_BIAS.t68 13.3681
R10010 CS_BIAS.n331 CS_BIAS.t78 13.3681
R10011 CS_BIAS.n336 CS_BIAS.t51 13.3681
R10012 CS_BIAS.n22 CS_BIAS.t0 13.3681
R10013 CS_BIAS.n28 CS_BIAS.t26 13.3681
R10014 CS_BIAS.n34 CS_BIAS.t22 13.3681
R10015 CS_BIAS.n42 CS_BIAS.t16 13.3681
R10016 CS_BIAS.n47 CS_BIAS.t20 13.3681
R10017 CS_BIAS.n55 CS_BIAS.t8 13.3681
R10018 CS_BIAS.n60 CS_BIAS.t14 13.3681
R10019 CS_BIAS.n0 CS_BIAS.t55 13.3681
R10020 CS_BIAS.n6 CS_BIAS.t35 13.3681
R10021 CS_BIAS.n12 CS_BIAS.t103 13.3681
R10022 CS_BIAS.n20 CS_BIAS.t64 13.3681
R10023 CS_BIAS.n178 CS_BIAS.t105 13.3681
R10024 CS_BIAS.n186 CS_BIAS.t83 13.3681
R10025 CS_BIAS.n191 CS_BIAS.t67 13.3681
R10026 CS_BIAS.n1654 CS_BIAS.t44 13.3681
R10027 CS_BIAS.n1671 CS_BIAS.t47 13.3681
R10028 CS_BIAS.n1642 CS_BIAS.t41 13.3681
R10029 CS_BIAS.n1707 CS_BIAS.t65 13.3681
R10030 CS_BIAS.n1630 CS_BIAS.t69 13.3681
R10031 CS_BIAS.n1624 CS_BIAS.t90 13.3681
R10032 CS_BIAS.n1618 CS_BIAS.t94 13.3681
R10033 CS_BIAS.n1508 CS_BIAS.t92 13.3681
R10034 CS_BIAS.n1525 CS_BIAS.t95 13.3681
R10035 CS_BIAS.n1496 CS_BIAS.t82 13.3681
R10036 CS_BIAS.n1561 CS_BIAS.t106 13.3681
R10037 CS_BIAS.n1484 CS_BIAS.t107 13.3681
R10038 CS_BIAS.n1478 CS_BIAS.t49 13.3681
R10039 CS_BIAS.n1472 CS_BIAS.t53 13.3681
R10040 CS_BIAS.n1362 CS_BIAS.t63 13.3681
R10041 CS_BIAS.n1379 CS_BIAS.t58 13.3681
R10042 CS_BIAS.n1350 CS_BIAS.t52 13.3681
R10043 CS_BIAS.n1415 CS_BIAS.t40 13.3681
R10044 CS_BIAS.n1338 CS_BIAS.t36 13.3681
R10045 CS_BIAS.n1332 CS_BIAS.t91 13.3681
R10046 CS_BIAS.n1326 CS_BIAS.t81 13.3681
R10047 CS_BIAS.n1216 CS_BIAS.t70 13.3681
R10048 CS_BIAS.n1233 CS_BIAS.t73 13.3681
R10049 CS_BIAS.n1204 CS_BIAS.t62 13.3681
R10050 CS_BIAS.n1269 CS_BIAS.t84 13.3681
R10051 CS_BIAS.n1192 CS_BIAS.t87 13.3681
R10052 CS_BIAS.n1186 CS_BIAS.t108 13.3681
R10053 CS_BIAS.n1180 CS_BIAS.t110 13.3681
R10054 CS_BIAS.n942 CS_BIAS.t10 13.3681
R10055 CS_BIAS.n959 CS_BIAS.t24 13.3681
R10056 CS_BIAS.n930 CS_BIAS.t4 13.3681
R10057 CS_BIAS.n995 CS_BIAS.t12 13.3681
R10058 CS_BIAS.n918 CS_BIAS.t28 13.3681
R10059 CS_BIAS.n912 CS_BIAS.t2 13.3681
R10060 CS_BIAS.n906 CS_BIAS.t6 13.3681
R10061 CS_BIAS.n882 CS_BIAS.t85 13.3681
R10062 CS_BIAS.n888 CS_BIAS.t45 13.3681
R10063 CS_BIAS.n894 CS_BIAS.t34 13.3681
R10064 CS_BIAS.n1124 CS_BIAS.t79 13.3681
R10065 CS_BIAS.n1071 CS_BIAS.t80 13.3681
R10066 CS_BIAS.n1088 CS_BIAS.t37 13.3681
R10067 CS_BIAS.n1059 CS_BIAS.t57 13.3681
R10068 CS_BIAS.n168 CS_BIAS.n166 12.5334
R10069 CS_BIAS.n1052 CS_BIAS.n1050 12.5334
R10070 CS_BIAS.n777 CS_BIAS.n774 11.0107
R10071 CS_BIAS.n861 CS_BIAS.n742 11.0107
R10072 CS_BIAS.n715 CS_BIAS.n596 11.0107
R10073 CS_BIAS.n631 CS_BIAS.n628 11.0107
R10074 CS_BIAS.n569 CS_BIAS.n450 11.0107
R10075 CS_BIAS.n485 CS_BIAS.n482 11.0107
R10076 CS_BIAS.n423 CS_BIAS.n304 11.0107
R10077 CS_BIAS.n339 CS_BIAS.n336 11.0107
R10078 CS_BIAS.n147 CS_BIAS.n28 11.0107
R10079 CS_BIAS.n63 CS_BIAS.n60 11.0107
R10080 CS_BIAS.n278 CS_BIAS.n6 11.0107
R10081 CS_BIAS.n194 CS_BIAS.n191 11.0107
R10082 CS_BIAS.n1657 CS_BIAS.n1654 11.0107
R10083 CS_BIAS.n1743 CS_BIAS.n1624 11.0107
R10084 CS_BIAS.n1511 CS_BIAS.n1508 11.0107
R10085 CS_BIAS.n1597 CS_BIAS.n1478 11.0107
R10086 CS_BIAS.n1365 CS_BIAS.n1362 11.0107
R10087 CS_BIAS.n1451 CS_BIAS.n1332 11.0107
R10088 CS_BIAS.n1219 CS_BIAS.n1216 11.0107
R10089 CS_BIAS.n1305 CS_BIAS.n1186 11.0107
R10090 CS_BIAS.n945 CS_BIAS.n942 11.0107
R10091 CS_BIAS.n1031 CS_BIAS.n912 11.0107
R10092 CS_BIAS.n1160 CS_BIAS.n888 11.0107
R10093 CS_BIAS.n1074 CS_BIAS.n1071 11.0107
R10094 CS_BIAS.n1764 CS_BIAS.n881 9.99414
R10095 CS_BIAS.n175 CS_BIAS.n174 9.50363
R10096 CS_BIAS.n1056 CS_BIAS.n1055 9.50363
R10097 CS_BIAS.n443 CS_BIAS.n297 7.75501
R10098 CS_BIAS.n1325 CS_BIAS.n1179 7.75501
R10099 CS_BIAS.n809 CS_BIAS.n761 7.58527
R10100 CS_BIAS.n756 CS_BIAS.n754 7.58527
R10101 CS_BIAS.n610 CS_BIAS.n608 7.58527
R10102 CS_BIAS.n663 CS_BIAS.n615 7.58527
R10103 CS_BIAS.n464 CS_BIAS.n462 7.58527
R10104 CS_BIAS.n517 CS_BIAS.n469 7.58527
R10105 CS_BIAS.n318 CS_BIAS.n316 7.58527
R10106 CS_BIAS.n371 CS_BIAS.n323 7.58527
R10107 CS_BIAS.n42 CS_BIAS.n40 7.58527
R10108 CS_BIAS.n95 CS_BIAS.n47 7.58527
R10109 CS_BIAS.n20 CS_BIAS.n18 7.58527
R10110 CS_BIAS.n226 CS_BIAS.n178 7.58527
R10111 CS_BIAS.n1690 CS_BIAS.n1642 7.58527
R10112 CS_BIAS.n1707 CS_BIAS.n1636 7.58527
R10113 CS_BIAS.n1544 CS_BIAS.n1496 7.58527
R10114 CS_BIAS.n1561 CS_BIAS.n1490 7.58527
R10115 CS_BIAS.n1398 CS_BIAS.n1350 7.58527
R10116 CS_BIAS.n1415 CS_BIAS.n1344 7.58527
R10117 CS_BIAS.n1252 CS_BIAS.n1204 7.58527
R10118 CS_BIAS.n1269 CS_BIAS.n1198 7.58527
R10119 CS_BIAS.n978 CS_BIAS.n930 7.58527
R10120 CS_BIAS.n995 CS_BIAS.n924 7.58527
R10121 CS_BIAS.n1124 CS_BIAS.n900 7.58527
R10122 CS_BIAS.n1107 CS_BIAS.n1059 7.58527
R10123 CS_BIAS.n1764 CS_BIAS.n1763 6.45974
R10124 CS_BIAS.n881 CS_BIAS.n880 5.43683
R10125 CS_BIAS.n735 CS_BIAS.n734 5.43683
R10126 CS_BIAS.n589 CS_BIAS.n588 5.43683
R10127 CS_BIAS.n443 CS_BIAS.n442 5.43683
R10128 CS_BIAS.n1763 CS_BIAS.n1762 5.43683
R10129 CS_BIAS.n1617 CS_BIAS.n1616 5.43683
R10130 CS_BIAS.n1471 CS_BIAS.n1470 5.43683
R10131 CS_BIAS.n1325 CS_BIAS.n1324 5.43683
R10132 CS_BIAS CS_BIAS.n1764 4.90925
R10133 CS_BIAS.n589 CS_BIAS.n443 2.31868
R10134 CS_BIAS.n735 CS_BIAS.n589 2.31868
R10135 CS_BIAS.n881 CS_BIAS.n735 2.31868
R10136 CS_BIAS.n1471 CS_BIAS.n1325 2.31868
R10137 CS_BIAS.n1617 CS_BIAS.n1471 2.31868
R10138 CS_BIAS.n1763 CS_BIAS.n1617 2.31868
R10139 CS_BIAS.n769 CS_BIAS.n767 1.71319
R10140 CS_BIAS.n844 CS_BIAS.n748 1.71319
R10141 CS_BIAS.n698 CS_BIAS.n602 1.71319
R10142 CS_BIAS.n623 CS_BIAS.n621 1.71319
R10143 CS_BIAS.n552 CS_BIAS.n456 1.71319
R10144 CS_BIAS.n477 CS_BIAS.n475 1.71319
R10145 CS_BIAS.n406 CS_BIAS.n310 1.71319
R10146 CS_BIAS.n331 CS_BIAS.n329 1.71319
R10147 CS_BIAS.n130 CS_BIAS.n34 1.71319
R10148 CS_BIAS.n55 CS_BIAS.n53 1.71319
R10149 CS_BIAS.n261 CS_BIAS.n12 1.71319
R10150 CS_BIAS.n186 CS_BIAS.n184 1.71319
R10151 CS_BIAS.n1671 CS_BIAS.n1648 1.71319
R10152 CS_BIAS.n1726 CS_BIAS.n1630 1.71319
R10153 CS_BIAS.n1525 CS_BIAS.n1502 1.71319
R10154 CS_BIAS.n1580 CS_BIAS.n1484 1.71319
R10155 CS_BIAS.n1379 CS_BIAS.n1356 1.71319
R10156 CS_BIAS.n1434 CS_BIAS.n1338 1.71319
R10157 CS_BIAS.n1233 CS_BIAS.n1210 1.71319
R10158 CS_BIAS.n1288 CS_BIAS.n1192 1.71319
R10159 CS_BIAS.n959 CS_BIAS.n936 1.71319
R10160 CS_BIAS.n1014 CS_BIAS.n918 1.71319
R10161 CS_BIAS.n1143 CS_BIAS.n894 1.71319
R10162 CS_BIAS.n1088 CS_BIAS.n1065 1.71319
R10163 CS_BIAS.n170 CS_BIAS.n168 1.63556
R10164 CS_BIAS.n1054 CS_BIAS.n1052 1.63556
R10165 CS_BIAS.n776 CS_BIAS.n775 1.0776
R10166 CS_BIAS.n1656 CS_BIAS.n1655 1.0776
R10167 CS_BIAS.n1510 CS_BIAS.n1509 1.0776
R10168 CS_BIAS.n1364 CS_BIAS.n1363 1.0776
R10169 CS_BIAS.n1218 CS_BIAS.n1217 1.0776
R10170 CS_BIAS.n944 CS_BIAS.n943 1.0776
R10171 CS_BIAS.n1073 CS_BIAS.n1072 1.0776
R10172 CS_BIAS.n630 CS_BIAS.n629 1.0776
R10173 CS_BIAS.n484 CS_BIAS.n483 1.0776
R10174 CS_BIAS.n338 CS_BIAS.n337 1.0776
R10175 CS_BIAS.n62 CS_BIAS.n61 1.0776
R10176 CS_BIAS.n193 CS_BIAS.n192 1.0776
R10177 CS_BIAS.n174 CS_BIAS.n170 0.818029
R10178 CS_BIAS.n174 CS_BIAS.n173 0.818029
R10179 CS_BIAS.n1055 CS_BIAS.n905 0.818029
R10180 CS_BIAS.n1055 CS_BIAS.n1054 0.818029
R10181 CS_BIAS.n880 CS_BIAS.n879 0.466196
R10182 CS_BIAS.n734 CS_BIAS.n733 0.466196
R10183 CS_BIAS.n588 CS_BIAS.n587 0.466196
R10184 CS_BIAS.n442 CS_BIAS.n441 0.466196
R10185 CS_BIAS.n166 CS_BIAS.n165 0.466196
R10186 CS_BIAS.n297 CS_BIAS.n296 0.466196
R10187 CS_BIAS.n1762 CS_BIAS.n1761 0.466196
R10188 CS_BIAS.n1616 CS_BIAS.n1615 0.466196
R10189 CS_BIAS.n1470 CS_BIAS.n1469 0.466196
R10190 CS_BIAS.n1324 CS_BIAS.n1323 0.466196
R10191 CS_BIAS.n1050 CS_BIAS.n1049 0.466196
R10192 CS_BIAS.n1179 CS_BIAS.n1178 0.466196
R10193 CS_BIAS.n879 CS_BIAS.n737 0.189894
R10194 CS_BIAS.n875 CS_BIAS.n737 0.189894
R10195 CS_BIAS.n875 CS_BIAS.n874 0.189894
R10196 CS_BIAS.n874 CS_BIAS.n873 0.189894
R10197 CS_BIAS.n873 CS_BIAS.n739 0.189894
R10198 CS_BIAS.n869 CS_BIAS.n739 0.189894
R10199 CS_BIAS.n869 CS_BIAS.n868 0.189894
R10200 CS_BIAS.n868 CS_BIAS.n867 0.189894
R10201 CS_BIAS.n867 CS_BIAS.n741 0.189894
R10202 CS_BIAS.n863 CS_BIAS.n741 0.189894
R10203 CS_BIAS.n863 CS_BIAS.n862 0.189894
R10204 CS_BIAS.n862 CS_BIAS.n743 0.189894
R10205 CS_BIAS.n858 CS_BIAS.n743 0.189894
R10206 CS_BIAS.n858 CS_BIAS.n857 0.189894
R10207 CS_BIAS.n857 CS_BIAS.n856 0.189894
R10208 CS_BIAS.n856 CS_BIAS.n745 0.189894
R10209 CS_BIAS.n852 CS_BIAS.n745 0.189894
R10210 CS_BIAS.n852 CS_BIAS.n851 0.189894
R10211 CS_BIAS.n851 CS_BIAS.n850 0.189894
R10212 CS_BIAS.n850 CS_BIAS.n747 0.189894
R10213 CS_BIAS.n846 CS_BIAS.n747 0.189894
R10214 CS_BIAS.n846 CS_BIAS.n845 0.189894
R10215 CS_BIAS.n845 CS_BIAS.n749 0.189894
R10216 CS_BIAS.n841 CS_BIAS.n749 0.189894
R10217 CS_BIAS.n841 CS_BIAS.n840 0.189894
R10218 CS_BIAS.n840 CS_BIAS.n839 0.189894
R10219 CS_BIAS.n839 CS_BIAS.n751 0.189894
R10220 CS_BIAS.n835 CS_BIAS.n751 0.189894
R10221 CS_BIAS.n835 CS_BIAS.n834 0.189894
R10222 CS_BIAS.n834 CS_BIAS.n833 0.189894
R10223 CS_BIAS.n833 CS_BIAS.n753 0.189894
R10224 CS_BIAS.n829 CS_BIAS.n753 0.189894
R10225 CS_BIAS.n829 CS_BIAS.n828 0.189894
R10226 CS_BIAS.n828 CS_BIAS.n827 0.189894
R10227 CS_BIAS.n827 CS_BIAS.n755 0.189894
R10228 CS_BIAS.n823 CS_BIAS.n755 0.189894
R10229 CS_BIAS.n823 CS_BIAS.n822 0.189894
R10230 CS_BIAS.n822 CS_BIAS.n821 0.189894
R10231 CS_BIAS.n821 CS_BIAS.n758 0.189894
R10232 CS_BIAS.n817 CS_BIAS.n758 0.189894
R10233 CS_BIAS.n817 CS_BIAS.n816 0.189894
R10234 CS_BIAS.n816 CS_BIAS.n815 0.189894
R10235 CS_BIAS.n815 CS_BIAS.n760 0.189894
R10236 CS_BIAS.n811 CS_BIAS.n760 0.189894
R10237 CS_BIAS.n811 CS_BIAS.n810 0.189894
R10238 CS_BIAS.n810 CS_BIAS.n762 0.189894
R10239 CS_BIAS.n806 CS_BIAS.n762 0.189894
R10240 CS_BIAS.n806 CS_BIAS.n805 0.189894
R10241 CS_BIAS.n805 CS_BIAS.n804 0.189894
R10242 CS_BIAS.n804 CS_BIAS.n764 0.189894
R10243 CS_BIAS.n800 CS_BIAS.n764 0.189894
R10244 CS_BIAS.n800 CS_BIAS.n799 0.189894
R10245 CS_BIAS.n799 CS_BIAS.n798 0.189894
R10246 CS_BIAS.n798 CS_BIAS.n766 0.189894
R10247 CS_BIAS.n794 CS_BIAS.n766 0.189894
R10248 CS_BIAS.n794 CS_BIAS.n793 0.189894
R10249 CS_BIAS.n793 CS_BIAS.n792 0.189894
R10250 CS_BIAS.n792 CS_BIAS.n768 0.189894
R10251 CS_BIAS.n788 CS_BIAS.n768 0.189894
R10252 CS_BIAS.n788 CS_BIAS.n787 0.189894
R10253 CS_BIAS.n787 CS_BIAS.n786 0.189894
R10254 CS_BIAS.n786 CS_BIAS.n771 0.189894
R10255 CS_BIAS.n782 CS_BIAS.n771 0.189894
R10256 CS_BIAS.n782 CS_BIAS.n781 0.189894
R10257 CS_BIAS.n781 CS_BIAS.n780 0.189894
R10258 CS_BIAS.n780 CS_BIAS.n773 0.189894
R10259 CS_BIAS.n776 CS_BIAS.n773 0.189894
R10260 CS_BIAS.n733 CS_BIAS.n591 0.189894
R10261 CS_BIAS.n729 CS_BIAS.n591 0.189894
R10262 CS_BIAS.n729 CS_BIAS.n728 0.189894
R10263 CS_BIAS.n728 CS_BIAS.n727 0.189894
R10264 CS_BIAS.n727 CS_BIAS.n593 0.189894
R10265 CS_BIAS.n723 CS_BIAS.n593 0.189894
R10266 CS_BIAS.n723 CS_BIAS.n722 0.189894
R10267 CS_BIAS.n722 CS_BIAS.n721 0.189894
R10268 CS_BIAS.n721 CS_BIAS.n595 0.189894
R10269 CS_BIAS.n717 CS_BIAS.n595 0.189894
R10270 CS_BIAS.n717 CS_BIAS.n716 0.189894
R10271 CS_BIAS.n716 CS_BIAS.n597 0.189894
R10272 CS_BIAS.n712 CS_BIAS.n597 0.189894
R10273 CS_BIAS.n712 CS_BIAS.n711 0.189894
R10274 CS_BIAS.n711 CS_BIAS.n710 0.189894
R10275 CS_BIAS.n710 CS_BIAS.n599 0.189894
R10276 CS_BIAS.n706 CS_BIAS.n599 0.189894
R10277 CS_BIAS.n706 CS_BIAS.n705 0.189894
R10278 CS_BIAS.n705 CS_BIAS.n704 0.189894
R10279 CS_BIAS.n704 CS_BIAS.n601 0.189894
R10280 CS_BIAS.n700 CS_BIAS.n601 0.189894
R10281 CS_BIAS.n700 CS_BIAS.n699 0.189894
R10282 CS_BIAS.n699 CS_BIAS.n603 0.189894
R10283 CS_BIAS.n695 CS_BIAS.n603 0.189894
R10284 CS_BIAS.n695 CS_BIAS.n694 0.189894
R10285 CS_BIAS.n694 CS_BIAS.n693 0.189894
R10286 CS_BIAS.n693 CS_BIAS.n605 0.189894
R10287 CS_BIAS.n689 CS_BIAS.n605 0.189894
R10288 CS_BIAS.n689 CS_BIAS.n688 0.189894
R10289 CS_BIAS.n688 CS_BIAS.n687 0.189894
R10290 CS_BIAS.n687 CS_BIAS.n607 0.189894
R10291 CS_BIAS.n683 CS_BIAS.n607 0.189894
R10292 CS_BIAS.n683 CS_BIAS.n682 0.189894
R10293 CS_BIAS.n682 CS_BIAS.n681 0.189894
R10294 CS_BIAS.n681 CS_BIAS.n609 0.189894
R10295 CS_BIAS.n677 CS_BIAS.n609 0.189894
R10296 CS_BIAS.n677 CS_BIAS.n676 0.189894
R10297 CS_BIAS.n676 CS_BIAS.n675 0.189894
R10298 CS_BIAS.n675 CS_BIAS.n612 0.189894
R10299 CS_BIAS.n671 CS_BIAS.n612 0.189894
R10300 CS_BIAS.n671 CS_BIAS.n670 0.189894
R10301 CS_BIAS.n670 CS_BIAS.n669 0.189894
R10302 CS_BIAS.n669 CS_BIAS.n614 0.189894
R10303 CS_BIAS.n665 CS_BIAS.n614 0.189894
R10304 CS_BIAS.n665 CS_BIAS.n664 0.189894
R10305 CS_BIAS.n664 CS_BIAS.n616 0.189894
R10306 CS_BIAS.n660 CS_BIAS.n616 0.189894
R10307 CS_BIAS.n660 CS_BIAS.n659 0.189894
R10308 CS_BIAS.n659 CS_BIAS.n658 0.189894
R10309 CS_BIAS.n658 CS_BIAS.n618 0.189894
R10310 CS_BIAS.n654 CS_BIAS.n618 0.189894
R10311 CS_BIAS.n654 CS_BIAS.n653 0.189894
R10312 CS_BIAS.n653 CS_BIAS.n652 0.189894
R10313 CS_BIAS.n652 CS_BIAS.n620 0.189894
R10314 CS_BIAS.n648 CS_BIAS.n620 0.189894
R10315 CS_BIAS.n648 CS_BIAS.n647 0.189894
R10316 CS_BIAS.n647 CS_BIAS.n646 0.189894
R10317 CS_BIAS.n646 CS_BIAS.n622 0.189894
R10318 CS_BIAS.n642 CS_BIAS.n622 0.189894
R10319 CS_BIAS.n642 CS_BIAS.n641 0.189894
R10320 CS_BIAS.n641 CS_BIAS.n640 0.189894
R10321 CS_BIAS.n640 CS_BIAS.n625 0.189894
R10322 CS_BIAS.n636 CS_BIAS.n625 0.189894
R10323 CS_BIAS.n636 CS_BIAS.n635 0.189894
R10324 CS_BIAS.n635 CS_BIAS.n634 0.189894
R10325 CS_BIAS.n634 CS_BIAS.n627 0.189894
R10326 CS_BIAS.n630 CS_BIAS.n627 0.189894
R10327 CS_BIAS.n587 CS_BIAS.n445 0.189894
R10328 CS_BIAS.n583 CS_BIAS.n445 0.189894
R10329 CS_BIAS.n583 CS_BIAS.n582 0.189894
R10330 CS_BIAS.n582 CS_BIAS.n581 0.189894
R10331 CS_BIAS.n581 CS_BIAS.n447 0.189894
R10332 CS_BIAS.n577 CS_BIAS.n447 0.189894
R10333 CS_BIAS.n577 CS_BIAS.n576 0.189894
R10334 CS_BIAS.n576 CS_BIAS.n575 0.189894
R10335 CS_BIAS.n575 CS_BIAS.n449 0.189894
R10336 CS_BIAS.n571 CS_BIAS.n449 0.189894
R10337 CS_BIAS.n571 CS_BIAS.n570 0.189894
R10338 CS_BIAS.n570 CS_BIAS.n451 0.189894
R10339 CS_BIAS.n566 CS_BIAS.n451 0.189894
R10340 CS_BIAS.n566 CS_BIAS.n565 0.189894
R10341 CS_BIAS.n565 CS_BIAS.n564 0.189894
R10342 CS_BIAS.n564 CS_BIAS.n453 0.189894
R10343 CS_BIAS.n560 CS_BIAS.n453 0.189894
R10344 CS_BIAS.n560 CS_BIAS.n559 0.189894
R10345 CS_BIAS.n559 CS_BIAS.n558 0.189894
R10346 CS_BIAS.n558 CS_BIAS.n455 0.189894
R10347 CS_BIAS.n554 CS_BIAS.n455 0.189894
R10348 CS_BIAS.n554 CS_BIAS.n553 0.189894
R10349 CS_BIAS.n553 CS_BIAS.n457 0.189894
R10350 CS_BIAS.n549 CS_BIAS.n457 0.189894
R10351 CS_BIAS.n549 CS_BIAS.n548 0.189894
R10352 CS_BIAS.n548 CS_BIAS.n547 0.189894
R10353 CS_BIAS.n547 CS_BIAS.n459 0.189894
R10354 CS_BIAS.n543 CS_BIAS.n459 0.189894
R10355 CS_BIAS.n543 CS_BIAS.n542 0.189894
R10356 CS_BIAS.n542 CS_BIAS.n541 0.189894
R10357 CS_BIAS.n541 CS_BIAS.n461 0.189894
R10358 CS_BIAS.n537 CS_BIAS.n461 0.189894
R10359 CS_BIAS.n537 CS_BIAS.n536 0.189894
R10360 CS_BIAS.n536 CS_BIAS.n535 0.189894
R10361 CS_BIAS.n535 CS_BIAS.n463 0.189894
R10362 CS_BIAS.n531 CS_BIAS.n463 0.189894
R10363 CS_BIAS.n531 CS_BIAS.n530 0.189894
R10364 CS_BIAS.n530 CS_BIAS.n529 0.189894
R10365 CS_BIAS.n529 CS_BIAS.n466 0.189894
R10366 CS_BIAS.n525 CS_BIAS.n466 0.189894
R10367 CS_BIAS.n525 CS_BIAS.n524 0.189894
R10368 CS_BIAS.n524 CS_BIAS.n523 0.189894
R10369 CS_BIAS.n523 CS_BIAS.n468 0.189894
R10370 CS_BIAS.n519 CS_BIAS.n468 0.189894
R10371 CS_BIAS.n519 CS_BIAS.n518 0.189894
R10372 CS_BIAS.n518 CS_BIAS.n470 0.189894
R10373 CS_BIAS.n514 CS_BIAS.n470 0.189894
R10374 CS_BIAS.n514 CS_BIAS.n513 0.189894
R10375 CS_BIAS.n513 CS_BIAS.n512 0.189894
R10376 CS_BIAS.n512 CS_BIAS.n472 0.189894
R10377 CS_BIAS.n508 CS_BIAS.n472 0.189894
R10378 CS_BIAS.n508 CS_BIAS.n507 0.189894
R10379 CS_BIAS.n507 CS_BIAS.n506 0.189894
R10380 CS_BIAS.n506 CS_BIAS.n474 0.189894
R10381 CS_BIAS.n502 CS_BIAS.n474 0.189894
R10382 CS_BIAS.n502 CS_BIAS.n501 0.189894
R10383 CS_BIAS.n501 CS_BIAS.n500 0.189894
R10384 CS_BIAS.n500 CS_BIAS.n476 0.189894
R10385 CS_BIAS.n496 CS_BIAS.n476 0.189894
R10386 CS_BIAS.n496 CS_BIAS.n495 0.189894
R10387 CS_BIAS.n495 CS_BIAS.n494 0.189894
R10388 CS_BIAS.n494 CS_BIAS.n479 0.189894
R10389 CS_BIAS.n490 CS_BIAS.n479 0.189894
R10390 CS_BIAS.n490 CS_BIAS.n489 0.189894
R10391 CS_BIAS.n489 CS_BIAS.n488 0.189894
R10392 CS_BIAS.n488 CS_BIAS.n481 0.189894
R10393 CS_BIAS.n484 CS_BIAS.n481 0.189894
R10394 CS_BIAS.n441 CS_BIAS.n299 0.189894
R10395 CS_BIAS.n437 CS_BIAS.n299 0.189894
R10396 CS_BIAS.n437 CS_BIAS.n436 0.189894
R10397 CS_BIAS.n436 CS_BIAS.n435 0.189894
R10398 CS_BIAS.n435 CS_BIAS.n301 0.189894
R10399 CS_BIAS.n431 CS_BIAS.n301 0.189894
R10400 CS_BIAS.n431 CS_BIAS.n430 0.189894
R10401 CS_BIAS.n430 CS_BIAS.n429 0.189894
R10402 CS_BIAS.n429 CS_BIAS.n303 0.189894
R10403 CS_BIAS.n425 CS_BIAS.n303 0.189894
R10404 CS_BIAS.n425 CS_BIAS.n424 0.189894
R10405 CS_BIAS.n424 CS_BIAS.n305 0.189894
R10406 CS_BIAS.n420 CS_BIAS.n305 0.189894
R10407 CS_BIAS.n420 CS_BIAS.n419 0.189894
R10408 CS_BIAS.n419 CS_BIAS.n418 0.189894
R10409 CS_BIAS.n418 CS_BIAS.n307 0.189894
R10410 CS_BIAS.n414 CS_BIAS.n307 0.189894
R10411 CS_BIAS.n414 CS_BIAS.n413 0.189894
R10412 CS_BIAS.n413 CS_BIAS.n412 0.189894
R10413 CS_BIAS.n412 CS_BIAS.n309 0.189894
R10414 CS_BIAS.n408 CS_BIAS.n309 0.189894
R10415 CS_BIAS.n408 CS_BIAS.n407 0.189894
R10416 CS_BIAS.n407 CS_BIAS.n311 0.189894
R10417 CS_BIAS.n403 CS_BIAS.n311 0.189894
R10418 CS_BIAS.n403 CS_BIAS.n402 0.189894
R10419 CS_BIAS.n402 CS_BIAS.n401 0.189894
R10420 CS_BIAS.n401 CS_BIAS.n313 0.189894
R10421 CS_BIAS.n397 CS_BIAS.n313 0.189894
R10422 CS_BIAS.n397 CS_BIAS.n396 0.189894
R10423 CS_BIAS.n396 CS_BIAS.n395 0.189894
R10424 CS_BIAS.n395 CS_BIAS.n315 0.189894
R10425 CS_BIAS.n391 CS_BIAS.n315 0.189894
R10426 CS_BIAS.n391 CS_BIAS.n390 0.189894
R10427 CS_BIAS.n390 CS_BIAS.n389 0.189894
R10428 CS_BIAS.n389 CS_BIAS.n317 0.189894
R10429 CS_BIAS.n385 CS_BIAS.n317 0.189894
R10430 CS_BIAS.n385 CS_BIAS.n384 0.189894
R10431 CS_BIAS.n384 CS_BIAS.n383 0.189894
R10432 CS_BIAS.n383 CS_BIAS.n320 0.189894
R10433 CS_BIAS.n379 CS_BIAS.n320 0.189894
R10434 CS_BIAS.n379 CS_BIAS.n378 0.189894
R10435 CS_BIAS.n378 CS_BIAS.n377 0.189894
R10436 CS_BIAS.n377 CS_BIAS.n322 0.189894
R10437 CS_BIAS.n373 CS_BIAS.n322 0.189894
R10438 CS_BIAS.n373 CS_BIAS.n372 0.189894
R10439 CS_BIAS.n372 CS_BIAS.n324 0.189894
R10440 CS_BIAS.n368 CS_BIAS.n324 0.189894
R10441 CS_BIAS.n368 CS_BIAS.n367 0.189894
R10442 CS_BIAS.n367 CS_BIAS.n366 0.189894
R10443 CS_BIAS.n366 CS_BIAS.n326 0.189894
R10444 CS_BIAS.n362 CS_BIAS.n326 0.189894
R10445 CS_BIAS.n362 CS_BIAS.n361 0.189894
R10446 CS_BIAS.n361 CS_BIAS.n360 0.189894
R10447 CS_BIAS.n360 CS_BIAS.n328 0.189894
R10448 CS_BIAS.n356 CS_BIAS.n328 0.189894
R10449 CS_BIAS.n356 CS_BIAS.n355 0.189894
R10450 CS_BIAS.n355 CS_BIAS.n354 0.189894
R10451 CS_BIAS.n354 CS_BIAS.n330 0.189894
R10452 CS_BIAS.n350 CS_BIAS.n330 0.189894
R10453 CS_BIAS.n350 CS_BIAS.n349 0.189894
R10454 CS_BIAS.n349 CS_BIAS.n348 0.189894
R10455 CS_BIAS.n348 CS_BIAS.n333 0.189894
R10456 CS_BIAS.n344 CS_BIAS.n333 0.189894
R10457 CS_BIAS.n344 CS_BIAS.n343 0.189894
R10458 CS_BIAS.n343 CS_BIAS.n342 0.189894
R10459 CS_BIAS.n342 CS_BIAS.n335 0.189894
R10460 CS_BIAS.n338 CS_BIAS.n335 0.189894
R10461 CS_BIAS.n165 CS_BIAS.n23 0.189894
R10462 CS_BIAS.n161 CS_BIAS.n23 0.189894
R10463 CS_BIAS.n161 CS_BIAS.n160 0.189894
R10464 CS_BIAS.n160 CS_BIAS.n159 0.189894
R10465 CS_BIAS.n159 CS_BIAS.n25 0.189894
R10466 CS_BIAS.n155 CS_BIAS.n25 0.189894
R10467 CS_BIAS.n155 CS_BIAS.n154 0.189894
R10468 CS_BIAS.n154 CS_BIAS.n153 0.189894
R10469 CS_BIAS.n153 CS_BIAS.n27 0.189894
R10470 CS_BIAS.n149 CS_BIAS.n27 0.189894
R10471 CS_BIAS.n149 CS_BIAS.n148 0.189894
R10472 CS_BIAS.n148 CS_BIAS.n29 0.189894
R10473 CS_BIAS.n144 CS_BIAS.n29 0.189894
R10474 CS_BIAS.n144 CS_BIAS.n143 0.189894
R10475 CS_BIAS.n143 CS_BIAS.n142 0.189894
R10476 CS_BIAS.n142 CS_BIAS.n31 0.189894
R10477 CS_BIAS.n138 CS_BIAS.n31 0.189894
R10478 CS_BIAS.n138 CS_BIAS.n137 0.189894
R10479 CS_BIAS.n137 CS_BIAS.n136 0.189894
R10480 CS_BIAS.n136 CS_BIAS.n33 0.189894
R10481 CS_BIAS.n132 CS_BIAS.n33 0.189894
R10482 CS_BIAS.n132 CS_BIAS.n131 0.189894
R10483 CS_BIAS.n131 CS_BIAS.n35 0.189894
R10484 CS_BIAS.n127 CS_BIAS.n35 0.189894
R10485 CS_BIAS.n127 CS_BIAS.n126 0.189894
R10486 CS_BIAS.n126 CS_BIAS.n125 0.189894
R10487 CS_BIAS.n125 CS_BIAS.n37 0.189894
R10488 CS_BIAS.n121 CS_BIAS.n37 0.189894
R10489 CS_BIAS.n121 CS_BIAS.n120 0.189894
R10490 CS_BIAS.n120 CS_BIAS.n119 0.189894
R10491 CS_BIAS.n119 CS_BIAS.n39 0.189894
R10492 CS_BIAS.n115 CS_BIAS.n39 0.189894
R10493 CS_BIAS.n115 CS_BIAS.n114 0.189894
R10494 CS_BIAS.n114 CS_BIAS.n113 0.189894
R10495 CS_BIAS.n113 CS_BIAS.n41 0.189894
R10496 CS_BIAS.n109 CS_BIAS.n41 0.189894
R10497 CS_BIAS.n109 CS_BIAS.n108 0.189894
R10498 CS_BIAS.n108 CS_BIAS.n107 0.189894
R10499 CS_BIAS.n107 CS_BIAS.n44 0.189894
R10500 CS_BIAS.n103 CS_BIAS.n44 0.189894
R10501 CS_BIAS.n103 CS_BIAS.n102 0.189894
R10502 CS_BIAS.n102 CS_BIAS.n101 0.189894
R10503 CS_BIAS.n101 CS_BIAS.n46 0.189894
R10504 CS_BIAS.n97 CS_BIAS.n46 0.189894
R10505 CS_BIAS.n97 CS_BIAS.n96 0.189894
R10506 CS_BIAS.n96 CS_BIAS.n48 0.189894
R10507 CS_BIAS.n92 CS_BIAS.n48 0.189894
R10508 CS_BIAS.n92 CS_BIAS.n91 0.189894
R10509 CS_BIAS.n91 CS_BIAS.n90 0.189894
R10510 CS_BIAS.n90 CS_BIAS.n50 0.189894
R10511 CS_BIAS.n86 CS_BIAS.n50 0.189894
R10512 CS_BIAS.n86 CS_BIAS.n85 0.189894
R10513 CS_BIAS.n85 CS_BIAS.n84 0.189894
R10514 CS_BIAS.n84 CS_BIAS.n52 0.189894
R10515 CS_BIAS.n80 CS_BIAS.n52 0.189894
R10516 CS_BIAS.n80 CS_BIAS.n79 0.189894
R10517 CS_BIAS.n79 CS_BIAS.n78 0.189894
R10518 CS_BIAS.n78 CS_BIAS.n54 0.189894
R10519 CS_BIAS.n74 CS_BIAS.n54 0.189894
R10520 CS_BIAS.n74 CS_BIAS.n73 0.189894
R10521 CS_BIAS.n73 CS_BIAS.n72 0.189894
R10522 CS_BIAS.n72 CS_BIAS.n57 0.189894
R10523 CS_BIAS.n68 CS_BIAS.n57 0.189894
R10524 CS_BIAS.n68 CS_BIAS.n67 0.189894
R10525 CS_BIAS.n67 CS_BIAS.n66 0.189894
R10526 CS_BIAS.n66 CS_BIAS.n59 0.189894
R10527 CS_BIAS.n62 CS_BIAS.n59 0.189894
R10528 CS_BIAS.n234 CS_BIAS.n233 0.189894
R10529 CS_BIAS.n233 CS_BIAS.n232 0.189894
R10530 CS_BIAS.n232 CS_BIAS.n177 0.189894
R10531 CS_BIAS.n228 CS_BIAS.n177 0.189894
R10532 CS_BIAS.n228 CS_BIAS.n227 0.189894
R10533 CS_BIAS.n227 CS_BIAS.n179 0.189894
R10534 CS_BIAS.n223 CS_BIAS.n179 0.189894
R10535 CS_BIAS.n223 CS_BIAS.n222 0.189894
R10536 CS_BIAS.n222 CS_BIAS.n221 0.189894
R10537 CS_BIAS.n221 CS_BIAS.n181 0.189894
R10538 CS_BIAS.n217 CS_BIAS.n181 0.189894
R10539 CS_BIAS.n217 CS_BIAS.n216 0.189894
R10540 CS_BIAS.n216 CS_BIAS.n215 0.189894
R10541 CS_BIAS.n215 CS_BIAS.n183 0.189894
R10542 CS_BIAS.n211 CS_BIAS.n183 0.189894
R10543 CS_BIAS.n211 CS_BIAS.n210 0.189894
R10544 CS_BIAS.n210 CS_BIAS.n209 0.189894
R10545 CS_BIAS.n209 CS_BIAS.n185 0.189894
R10546 CS_BIAS.n205 CS_BIAS.n185 0.189894
R10547 CS_BIAS.n205 CS_BIAS.n204 0.189894
R10548 CS_BIAS.n204 CS_BIAS.n203 0.189894
R10549 CS_BIAS.n203 CS_BIAS.n188 0.189894
R10550 CS_BIAS.n199 CS_BIAS.n188 0.189894
R10551 CS_BIAS.n199 CS_BIAS.n198 0.189894
R10552 CS_BIAS.n198 CS_BIAS.n197 0.189894
R10553 CS_BIAS.n197 CS_BIAS.n190 0.189894
R10554 CS_BIAS.n193 CS_BIAS.n190 0.189894
R10555 CS_BIAS.n296 CS_BIAS.n1 0.189894
R10556 CS_BIAS.n292 CS_BIAS.n1 0.189894
R10557 CS_BIAS.n292 CS_BIAS.n291 0.189894
R10558 CS_BIAS.n291 CS_BIAS.n290 0.189894
R10559 CS_BIAS.n290 CS_BIAS.n3 0.189894
R10560 CS_BIAS.n286 CS_BIAS.n3 0.189894
R10561 CS_BIAS.n286 CS_BIAS.n285 0.189894
R10562 CS_BIAS.n285 CS_BIAS.n284 0.189894
R10563 CS_BIAS.n284 CS_BIAS.n5 0.189894
R10564 CS_BIAS.n280 CS_BIAS.n5 0.189894
R10565 CS_BIAS.n280 CS_BIAS.n279 0.189894
R10566 CS_BIAS.n279 CS_BIAS.n7 0.189894
R10567 CS_BIAS.n275 CS_BIAS.n7 0.189894
R10568 CS_BIAS.n275 CS_BIAS.n274 0.189894
R10569 CS_BIAS.n274 CS_BIAS.n273 0.189894
R10570 CS_BIAS.n273 CS_BIAS.n9 0.189894
R10571 CS_BIAS.n269 CS_BIAS.n9 0.189894
R10572 CS_BIAS.n269 CS_BIAS.n268 0.189894
R10573 CS_BIAS.n268 CS_BIAS.n267 0.189894
R10574 CS_BIAS.n267 CS_BIAS.n11 0.189894
R10575 CS_BIAS.n263 CS_BIAS.n11 0.189894
R10576 CS_BIAS.n263 CS_BIAS.n262 0.189894
R10577 CS_BIAS.n262 CS_BIAS.n13 0.189894
R10578 CS_BIAS.n258 CS_BIAS.n13 0.189894
R10579 CS_BIAS.n258 CS_BIAS.n257 0.189894
R10580 CS_BIAS.n257 CS_BIAS.n256 0.189894
R10581 CS_BIAS.n256 CS_BIAS.n15 0.189894
R10582 CS_BIAS.n252 CS_BIAS.n15 0.189894
R10583 CS_BIAS.n252 CS_BIAS.n251 0.189894
R10584 CS_BIAS.n251 CS_BIAS.n250 0.189894
R10585 CS_BIAS.n250 CS_BIAS.n17 0.189894
R10586 CS_BIAS.n246 CS_BIAS.n17 0.189894
R10587 CS_BIAS.n246 CS_BIAS.n245 0.189894
R10588 CS_BIAS.n245 CS_BIAS.n244 0.189894
R10589 CS_BIAS.n244 CS_BIAS.n19 0.189894
R10590 CS_BIAS.n240 CS_BIAS.n19 0.189894
R10591 CS_BIAS.n240 CS_BIAS.n239 0.189894
R10592 CS_BIAS.n239 CS_BIAS.n238 0.189894
R10593 CS_BIAS.n1656 CS_BIAS.n1653 0.189894
R10594 CS_BIAS.n1660 CS_BIAS.n1653 0.189894
R10595 CS_BIAS.n1661 CS_BIAS.n1660 0.189894
R10596 CS_BIAS.n1662 CS_BIAS.n1661 0.189894
R10597 CS_BIAS.n1662 CS_BIAS.n1651 0.189894
R10598 CS_BIAS.n1666 CS_BIAS.n1651 0.189894
R10599 CS_BIAS.n1667 CS_BIAS.n1666 0.189894
R10600 CS_BIAS.n1668 CS_BIAS.n1667 0.189894
R10601 CS_BIAS.n1668 CS_BIAS.n1649 0.189894
R10602 CS_BIAS.n1673 CS_BIAS.n1649 0.189894
R10603 CS_BIAS.n1674 CS_BIAS.n1673 0.189894
R10604 CS_BIAS.n1675 CS_BIAS.n1674 0.189894
R10605 CS_BIAS.n1675 CS_BIAS.n1647 0.189894
R10606 CS_BIAS.n1679 CS_BIAS.n1647 0.189894
R10607 CS_BIAS.n1680 CS_BIAS.n1679 0.189894
R10608 CS_BIAS.n1681 CS_BIAS.n1680 0.189894
R10609 CS_BIAS.n1681 CS_BIAS.n1645 0.189894
R10610 CS_BIAS.n1685 CS_BIAS.n1645 0.189894
R10611 CS_BIAS.n1686 CS_BIAS.n1685 0.189894
R10612 CS_BIAS.n1687 CS_BIAS.n1686 0.189894
R10613 CS_BIAS.n1687 CS_BIAS.n1643 0.189894
R10614 CS_BIAS.n1691 CS_BIAS.n1643 0.189894
R10615 CS_BIAS.n1692 CS_BIAS.n1691 0.189894
R10616 CS_BIAS.n1692 CS_BIAS.n1641 0.189894
R10617 CS_BIAS.n1696 CS_BIAS.n1641 0.189894
R10618 CS_BIAS.n1697 CS_BIAS.n1696 0.189894
R10619 CS_BIAS.n1698 CS_BIAS.n1697 0.189894
R10620 CS_BIAS.n1698 CS_BIAS.n1639 0.189894
R10621 CS_BIAS.n1702 CS_BIAS.n1639 0.189894
R10622 CS_BIAS.n1703 CS_BIAS.n1702 0.189894
R10623 CS_BIAS.n1704 CS_BIAS.n1703 0.189894
R10624 CS_BIAS.n1704 CS_BIAS.n1637 0.189894
R10625 CS_BIAS.n1709 CS_BIAS.n1637 0.189894
R10626 CS_BIAS.n1710 CS_BIAS.n1709 0.189894
R10627 CS_BIAS.n1711 CS_BIAS.n1710 0.189894
R10628 CS_BIAS.n1711 CS_BIAS.n1635 0.189894
R10629 CS_BIAS.n1715 CS_BIAS.n1635 0.189894
R10630 CS_BIAS.n1716 CS_BIAS.n1715 0.189894
R10631 CS_BIAS.n1717 CS_BIAS.n1716 0.189894
R10632 CS_BIAS.n1717 CS_BIAS.n1633 0.189894
R10633 CS_BIAS.n1721 CS_BIAS.n1633 0.189894
R10634 CS_BIAS.n1722 CS_BIAS.n1721 0.189894
R10635 CS_BIAS.n1723 CS_BIAS.n1722 0.189894
R10636 CS_BIAS.n1723 CS_BIAS.n1631 0.189894
R10637 CS_BIAS.n1727 CS_BIAS.n1631 0.189894
R10638 CS_BIAS.n1728 CS_BIAS.n1727 0.189894
R10639 CS_BIAS.n1728 CS_BIAS.n1629 0.189894
R10640 CS_BIAS.n1732 CS_BIAS.n1629 0.189894
R10641 CS_BIAS.n1733 CS_BIAS.n1732 0.189894
R10642 CS_BIAS.n1734 CS_BIAS.n1733 0.189894
R10643 CS_BIAS.n1734 CS_BIAS.n1627 0.189894
R10644 CS_BIAS.n1738 CS_BIAS.n1627 0.189894
R10645 CS_BIAS.n1739 CS_BIAS.n1738 0.189894
R10646 CS_BIAS.n1740 CS_BIAS.n1739 0.189894
R10647 CS_BIAS.n1740 CS_BIAS.n1625 0.189894
R10648 CS_BIAS.n1744 CS_BIAS.n1625 0.189894
R10649 CS_BIAS.n1745 CS_BIAS.n1744 0.189894
R10650 CS_BIAS.n1745 CS_BIAS.n1623 0.189894
R10651 CS_BIAS.n1749 CS_BIAS.n1623 0.189894
R10652 CS_BIAS.n1750 CS_BIAS.n1749 0.189894
R10653 CS_BIAS.n1751 CS_BIAS.n1750 0.189894
R10654 CS_BIAS.n1751 CS_BIAS.n1621 0.189894
R10655 CS_BIAS.n1755 CS_BIAS.n1621 0.189894
R10656 CS_BIAS.n1756 CS_BIAS.n1755 0.189894
R10657 CS_BIAS.n1757 CS_BIAS.n1756 0.189894
R10658 CS_BIAS.n1757 CS_BIAS.n1619 0.189894
R10659 CS_BIAS.n1761 CS_BIAS.n1619 0.189894
R10660 CS_BIAS.n1510 CS_BIAS.n1507 0.189894
R10661 CS_BIAS.n1514 CS_BIAS.n1507 0.189894
R10662 CS_BIAS.n1515 CS_BIAS.n1514 0.189894
R10663 CS_BIAS.n1516 CS_BIAS.n1515 0.189894
R10664 CS_BIAS.n1516 CS_BIAS.n1505 0.189894
R10665 CS_BIAS.n1520 CS_BIAS.n1505 0.189894
R10666 CS_BIAS.n1521 CS_BIAS.n1520 0.189894
R10667 CS_BIAS.n1522 CS_BIAS.n1521 0.189894
R10668 CS_BIAS.n1522 CS_BIAS.n1503 0.189894
R10669 CS_BIAS.n1527 CS_BIAS.n1503 0.189894
R10670 CS_BIAS.n1528 CS_BIAS.n1527 0.189894
R10671 CS_BIAS.n1529 CS_BIAS.n1528 0.189894
R10672 CS_BIAS.n1529 CS_BIAS.n1501 0.189894
R10673 CS_BIAS.n1533 CS_BIAS.n1501 0.189894
R10674 CS_BIAS.n1534 CS_BIAS.n1533 0.189894
R10675 CS_BIAS.n1535 CS_BIAS.n1534 0.189894
R10676 CS_BIAS.n1535 CS_BIAS.n1499 0.189894
R10677 CS_BIAS.n1539 CS_BIAS.n1499 0.189894
R10678 CS_BIAS.n1540 CS_BIAS.n1539 0.189894
R10679 CS_BIAS.n1541 CS_BIAS.n1540 0.189894
R10680 CS_BIAS.n1541 CS_BIAS.n1497 0.189894
R10681 CS_BIAS.n1545 CS_BIAS.n1497 0.189894
R10682 CS_BIAS.n1546 CS_BIAS.n1545 0.189894
R10683 CS_BIAS.n1546 CS_BIAS.n1495 0.189894
R10684 CS_BIAS.n1550 CS_BIAS.n1495 0.189894
R10685 CS_BIAS.n1551 CS_BIAS.n1550 0.189894
R10686 CS_BIAS.n1552 CS_BIAS.n1551 0.189894
R10687 CS_BIAS.n1552 CS_BIAS.n1493 0.189894
R10688 CS_BIAS.n1556 CS_BIAS.n1493 0.189894
R10689 CS_BIAS.n1557 CS_BIAS.n1556 0.189894
R10690 CS_BIAS.n1558 CS_BIAS.n1557 0.189894
R10691 CS_BIAS.n1558 CS_BIAS.n1491 0.189894
R10692 CS_BIAS.n1563 CS_BIAS.n1491 0.189894
R10693 CS_BIAS.n1564 CS_BIAS.n1563 0.189894
R10694 CS_BIAS.n1565 CS_BIAS.n1564 0.189894
R10695 CS_BIAS.n1565 CS_BIAS.n1489 0.189894
R10696 CS_BIAS.n1569 CS_BIAS.n1489 0.189894
R10697 CS_BIAS.n1570 CS_BIAS.n1569 0.189894
R10698 CS_BIAS.n1571 CS_BIAS.n1570 0.189894
R10699 CS_BIAS.n1571 CS_BIAS.n1487 0.189894
R10700 CS_BIAS.n1575 CS_BIAS.n1487 0.189894
R10701 CS_BIAS.n1576 CS_BIAS.n1575 0.189894
R10702 CS_BIAS.n1577 CS_BIAS.n1576 0.189894
R10703 CS_BIAS.n1577 CS_BIAS.n1485 0.189894
R10704 CS_BIAS.n1581 CS_BIAS.n1485 0.189894
R10705 CS_BIAS.n1582 CS_BIAS.n1581 0.189894
R10706 CS_BIAS.n1582 CS_BIAS.n1483 0.189894
R10707 CS_BIAS.n1586 CS_BIAS.n1483 0.189894
R10708 CS_BIAS.n1587 CS_BIAS.n1586 0.189894
R10709 CS_BIAS.n1588 CS_BIAS.n1587 0.189894
R10710 CS_BIAS.n1588 CS_BIAS.n1481 0.189894
R10711 CS_BIAS.n1592 CS_BIAS.n1481 0.189894
R10712 CS_BIAS.n1593 CS_BIAS.n1592 0.189894
R10713 CS_BIAS.n1594 CS_BIAS.n1593 0.189894
R10714 CS_BIAS.n1594 CS_BIAS.n1479 0.189894
R10715 CS_BIAS.n1598 CS_BIAS.n1479 0.189894
R10716 CS_BIAS.n1599 CS_BIAS.n1598 0.189894
R10717 CS_BIAS.n1599 CS_BIAS.n1477 0.189894
R10718 CS_BIAS.n1603 CS_BIAS.n1477 0.189894
R10719 CS_BIAS.n1604 CS_BIAS.n1603 0.189894
R10720 CS_BIAS.n1605 CS_BIAS.n1604 0.189894
R10721 CS_BIAS.n1605 CS_BIAS.n1475 0.189894
R10722 CS_BIAS.n1609 CS_BIAS.n1475 0.189894
R10723 CS_BIAS.n1610 CS_BIAS.n1609 0.189894
R10724 CS_BIAS.n1611 CS_BIAS.n1610 0.189894
R10725 CS_BIAS.n1611 CS_BIAS.n1473 0.189894
R10726 CS_BIAS.n1615 CS_BIAS.n1473 0.189894
R10727 CS_BIAS.n1364 CS_BIAS.n1361 0.189894
R10728 CS_BIAS.n1368 CS_BIAS.n1361 0.189894
R10729 CS_BIAS.n1369 CS_BIAS.n1368 0.189894
R10730 CS_BIAS.n1370 CS_BIAS.n1369 0.189894
R10731 CS_BIAS.n1370 CS_BIAS.n1359 0.189894
R10732 CS_BIAS.n1374 CS_BIAS.n1359 0.189894
R10733 CS_BIAS.n1375 CS_BIAS.n1374 0.189894
R10734 CS_BIAS.n1376 CS_BIAS.n1375 0.189894
R10735 CS_BIAS.n1376 CS_BIAS.n1357 0.189894
R10736 CS_BIAS.n1381 CS_BIAS.n1357 0.189894
R10737 CS_BIAS.n1382 CS_BIAS.n1381 0.189894
R10738 CS_BIAS.n1383 CS_BIAS.n1382 0.189894
R10739 CS_BIAS.n1383 CS_BIAS.n1355 0.189894
R10740 CS_BIAS.n1387 CS_BIAS.n1355 0.189894
R10741 CS_BIAS.n1388 CS_BIAS.n1387 0.189894
R10742 CS_BIAS.n1389 CS_BIAS.n1388 0.189894
R10743 CS_BIAS.n1389 CS_BIAS.n1353 0.189894
R10744 CS_BIAS.n1393 CS_BIAS.n1353 0.189894
R10745 CS_BIAS.n1394 CS_BIAS.n1393 0.189894
R10746 CS_BIAS.n1395 CS_BIAS.n1394 0.189894
R10747 CS_BIAS.n1395 CS_BIAS.n1351 0.189894
R10748 CS_BIAS.n1399 CS_BIAS.n1351 0.189894
R10749 CS_BIAS.n1400 CS_BIAS.n1399 0.189894
R10750 CS_BIAS.n1400 CS_BIAS.n1349 0.189894
R10751 CS_BIAS.n1404 CS_BIAS.n1349 0.189894
R10752 CS_BIAS.n1405 CS_BIAS.n1404 0.189894
R10753 CS_BIAS.n1406 CS_BIAS.n1405 0.189894
R10754 CS_BIAS.n1406 CS_BIAS.n1347 0.189894
R10755 CS_BIAS.n1410 CS_BIAS.n1347 0.189894
R10756 CS_BIAS.n1411 CS_BIAS.n1410 0.189894
R10757 CS_BIAS.n1412 CS_BIAS.n1411 0.189894
R10758 CS_BIAS.n1412 CS_BIAS.n1345 0.189894
R10759 CS_BIAS.n1417 CS_BIAS.n1345 0.189894
R10760 CS_BIAS.n1418 CS_BIAS.n1417 0.189894
R10761 CS_BIAS.n1419 CS_BIAS.n1418 0.189894
R10762 CS_BIAS.n1419 CS_BIAS.n1343 0.189894
R10763 CS_BIAS.n1423 CS_BIAS.n1343 0.189894
R10764 CS_BIAS.n1424 CS_BIAS.n1423 0.189894
R10765 CS_BIAS.n1425 CS_BIAS.n1424 0.189894
R10766 CS_BIAS.n1425 CS_BIAS.n1341 0.189894
R10767 CS_BIAS.n1429 CS_BIAS.n1341 0.189894
R10768 CS_BIAS.n1430 CS_BIAS.n1429 0.189894
R10769 CS_BIAS.n1431 CS_BIAS.n1430 0.189894
R10770 CS_BIAS.n1431 CS_BIAS.n1339 0.189894
R10771 CS_BIAS.n1435 CS_BIAS.n1339 0.189894
R10772 CS_BIAS.n1436 CS_BIAS.n1435 0.189894
R10773 CS_BIAS.n1436 CS_BIAS.n1337 0.189894
R10774 CS_BIAS.n1440 CS_BIAS.n1337 0.189894
R10775 CS_BIAS.n1441 CS_BIAS.n1440 0.189894
R10776 CS_BIAS.n1442 CS_BIAS.n1441 0.189894
R10777 CS_BIAS.n1442 CS_BIAS.n1335 0.189894
R10778 CS_BIAS.n1446 CS_BIAS.n1335 0.189894
R10779 CS_BIAS.n1447 CS_BIAS.n1446 0.189894
R10780 CS_BIAS.n1448 CS_BIAS.n1447 0.189894
R10781 CS_BIAS.n1448 CS_BIAS.n1333 0.189894
R10782 CS_BIAS.n1452 CS_BIAS.n1333 0.189894
R10783 CS_BIAS.n1453 CS_BIAS.n1452 0.189894
R10784 CS_BIAS.n1453 CS_BIAS.n1331 0.189894
R10785 CS_BIAS.n1457 CS_BIAS.n1331 0.189894
R10786 CS_BIAS.n1458 CS_BIAS.n1457 0.189894
R10787 CS_BIAS.n1459 CS_BIAS.n1458 0.189894
R10788 CS_BIAS.n1459 CS_BIAS.n1329 0.189894
R10789 CS_BIAS.n1463 CS_BIAS.n1329 0.189894
R10790 CS_BIAS.n1464 CS_BIAS.n1463 0.189894
R10791 CS_BIAS.n1465 CS_BIAS.n1464 0.189894
R10792 CS_BIAS.n1465 CS_BIAS.n1327 0.189894
R10793 CS_BIAS.n1469 CS_BIAS.n1327 0.189894
R10794 CS_BIAS.n1218 CS_BIAS.n1215 0.189894
R10795 CS_BIAS.n1222 CS_BIAS.n1215 0.189894
R10796 CS_BIAS.n1223 CS_BIAS.n1222 0.189894
R10797 CS_BIAS.n1224 CS_BIAS.n1223 0.189894
R10798 CS_BIAS.n1224 CS_BIAS.n1213 0.189894
R10799 CS_BIAS.n1228 CS_BIAS.n1213 0.189894
R10800 CS_BIAS.n1229 CS_BIAS.n1228 0.189894
R10801 CS_BIAS.n1230 CS_BIAS.n1229 0.189894
R10802 CS_BIAS.n1230 CS_BIAS.n1211 0.189894
R10803 CS_BIAS.n1235 CS_BIAS.n1211 0.189894
R10804 CS_BIAS.n1236 CS_BIAS.n1235 0.189894
R10805 CS_BIAS.n1237 CS_BIAS.n1236 0.189894
R10806 CS_BIAS.n1237 CS_BIAS.n1209 0.189894
R10807 CS_BIAS.n1241 CS_BIAS.n1209 0.189894
R10808 CS_BIAS.n1242 CS_BIAS.n1241 0.189894
R10809 CS_BIAS.n1243 CS_BIAS.n1242 0.189894
R10810 CS_BIAS.n1243 CS_BIAS.n1207 0.189894
R10811 CS_BIAS.n1247 CS_BIAS.n1207 0.189894
R10812 CS_BIAS.n1248 CS_BIAS.n1247 0.189894
R10813 CS_BIAS.n1249 CS_BIAS.n1248 0.189894
R10814 CS_BIAS.n1249 CS_BIAS.n1205 0.189894
R10815 CS_BIAS.n1253 CS_BIAS.n1205 0.189894
R10816 CS_BIAS.n1254 CS_BIAS.n1253 0.189894
R10817 CS_BIAS.n1254 CS_BIAS.n1203 0.189894
R10818 CS_BIAS.n1258 CS_BIAS.n1203 0.189894
R10819 CS_BIAS.n1259 CS_BIAS.n1258 0.189894
R10820 CS_BIAS.n1260 CS_BIAS.n1259 0.189894
R10821 CS_BIAS.n1260 CS_BIAS.n1201 0.189894
R10822 CS_BIAS.n1264 CS_BIAS.n1201 0.189894
R10823 CS_BIAS.n1265 CS_BIAS.n1264 0.189894
R10824 CS_BIAS.n1266 CS_BIAS.n1265 0.189894
R10825 CS_BIAS.n1266 CS_BIAS.n1199 0.189894
R10826 CS_BIAS.n1271 CS_BIAS.n1199 0.189894
R10827 CS_BIAS.n1272 CS_BIAS.n1271 0.189894
R10828 CS_BIAS.n1273 CS_BIAS.n1272 0.189894
R10829 CS_BIAS.n1273 CS_BIAS.n1197 0.189894
R10830 CS_BIAS.n1277 CS_BIAS.n1197 0.189894
R10831 CS_BIAS.n1278 CS_BIAS.n1277 0.189894
R10832 CS_BIAS.n1279 CS_BIAS.n1278 0.189894
R10833 CS_BIAS.n1279 CS_BIAS.n1195 0.189894
R10834 CS_BIAS.n1283 CS_BIAS.n1195 0.189894
R10835 CS_BIAS.n1284 CS_BIAS.n1283 0.189894
R10836 CS_BIAS.n1285 CS_BIAS.n1284 0.189894
R10837 CS_BIAS.n1285 CS_BIAS.n1193 0.189894
R10838 CS_BIAS.n1289 CS_BIAS.n1193 0.189894
R10839 CS_BIAS.n1290 CS_BIAS.n1289 0.189894
R10840 CS_BIAS.n1290 CS_BIAS.n1191 0.189894
R10841 CS_BIAS.n1294 CS_BIAS.n1191 0.189894
R10842 CS_BIAS.n1295 CS_BIAS.n1294 0.189894
R10843 CS_BIAS.n1296 CS_BIAS.n1295 0.189894
R10844 CS_BIAS.n1296 CS_BIAS.n1189 0.189894
R10845 CS_BIAS.n1300 CS_BIAS.n1189 0.189894
R10846 CS_BIAS.n1301 CS_BIAS.n1300 0.189894
R10847 CS_BIAS.n1302 CS_BIAS.n1301 0.189894
R10848 CS_BIAS.n1302 CS_BIAS.n1187 0.189894
R10849 CS_BIAS.n1306 CS_BIAS.n1187 0.189894
R10850 CS_BIAS.n1307 CS_BIAS.n1306 0.189894
R10851 CS_BIAS.n1307 CS_BIAS.n1185 0.189894
R10852 CS_BIAS.n1311 CS_BIAS.n1185 0.189894
R10853 CS_BIAS.n1312 CS_BIAS.n1311 0.189894
R10854 CS_BIAS.n1313 CS_BIAS.n1312 0.189894
R10855 CS_BIAS.n1313 CS_BIAS.n1183 0.189894
R10856 CS_BIAS.n1317 CS_BIAS.n1183 0.189894
R10857 CS_BIAS.n1318 CS_BIAS.n1317 0.189894
R10858 CS_BIAS.n1319 CS_BIAS.n1318 0.189894
R10859 CS_BIAS.n1319 CS_BIAS.n1181 0.189894
R10860 CS_BIAS.n1323 CS_BIAS.n1181 0.189894
R10861 CS_BIAS.n944 CS_BIAS.n941 0.189894
R10862 CS_BIAS.n948 CS_BIAS.n941 0.189894
R10863 CS_BIAS.n949 CS_BIAS.n948 0.189894
R10864 CS_BIAS.n950 CS_BIAS.n949 0.189894
R10865 CS_BIAS.n950 CS_BIAS.n939 0.189894
R10866 CS_BIAS.n954 CS_BIAS.n939 0.189894
R10867 CS_BIAS.n955 CS_BIAS.n954 0.189894
R10868 CS_BIAS.n956 CS_BIAS.n955 0.189894
R10869 CS_BIAS.n956 CS_BIAS.n937 0.189894
R10870 CS_BIAS.n961 CS_BIAS.n937 0.189894
R10871 CS_BIAS.n962 CS_BIAS.n961 0.189894
R10872 CS_BIAS.n963 CS_BIAS.n962 0.189894
R10873 CS_BIAS.n963 CS_BIAS.n935 0.189894
R10874 CS_BIAS.n967 CS_BIAS.n935 0.189894
R10875 CS_BIAS.n968 CS_BIAS.n967 0.189894
R10876 CS_BIAS.n969 CS_BIAS.n968 0.189894
R10877 CS_BIAS.n969 CS_BIAS.n933 0.189894
R10878 CS_BIAS.n973 CS_BIAS.n933 0.189894
R10879 CS_BIAS.n974 CS_BIAS.n973 0.189894
R10880 CS_BIAS.n975 CS_BIAS.n974 0.189894
R10881 CS_BIAS.n975 CS_BIAS.n931 0.189894
R10882 CS_BIAS.n979 CS_BIAS.n931 0.189894
R10883 CS_BIAS.n980 CS_BIAS.n979 0.189894
R10884 CS_BIAS.n980 CS_BIAS.n929 0.189894
R10885 CS_BIAS.n984 CS_BIAS.n929 0.189894
R10886 CS_BIAS.n985 CS_BIAS.n984 0.189894
R10887 CS_BIAS.n986 CS_BIAS.n985 0.189894
R10888 CS_BIAS.n986 CS_BIAS.n927 0.189894
R10889 CS_BIAS.n990 CS_BIAS.n927 0.189894
R10890 CS_BIAS.n991 CS_BIAS.n990 0.189894
R10891 CS_BIAS.n992 CS_BIAS.n991 0.189894
R10892 CS_BIAS.n992 CS_BIAS.n925 0.189894
R10893 CS_BIAS.n997 CS_BIAS.n925 0.189894
R10894 CS_BIAS.n998 CS_BIAS.n997 0.189894
R10895 CS_BIAS.n999 CS_BIAS.n998 0.189894
R10896 CS_BIAS.n999 CS_BIAS.n923 0.189894
R10897 CS_BIAS.n1003 CS_BIAS.n923 0.189894
R10898 CS_BIAS.n1004 CS_BIAS.n1003 0.189894
R10899 CS_BIAS.n1005 CS_BIAS.n1004 0.189894
R10900 CS_BIAS.n1005 CS_BIAS.n921 0.189894
R10901 CS_BIAS.n1009 CS_BIAS.n921 0.189894
R10902 CS_BIAS.n1010 CS_BIAS.n1009 0.189894
R10903 CS_BIAS.n1011 CS_BIAS.n1010 0.189894
R10904 CS_BIAS.n1011 CS_BIAS.n919 0.189894
R10905 CS_BIAS.n1015 CS_BIAS.n919 0.189894
R10906 CS_BIAS.n1016 CS_BIAS.n1015 0.189894
R10907 CS_BIAS.n1016 CS_BIAS.n917 0.189894
R10908 CS_BIAS.n1020 CS_BIAS.n917 0.189894
R10909 CS_BIAS.n1021 CS_BIAS.n1020 0.189894
R10910 CS_BIAS.n1022 CS_BIAS.n1021 0.189894
R10911 CS_BIAS.n1022 CS_BIAS.n915 0.189894
R10912 CS_BIAS.n1026 CS_BIAS.n915 0.189894
R10913 CS_BIAS.n1027 CS_BIAS.n1026 0.189894
R10914 CS_BIAS.n1028 CS_BIAS.n1027 0.189894
R10915 CS_BIAS.n1028 CS_BIAS.n913 0.189894
R10916 CS_BIAS.n1032 CS_BIAS.n913 0.189894
R10917 CS_BIAS.n1033 CS_BIAS.n1032 0.189894
R10918 CS_BIAS.n1033 CS_BIAS.n911 0.189894
R10919 CS_BIAS.n1037 CS_BIAS.n911 0.189894
R10920 CS_BIAS.n1038 CS_BIAS.n1037 0.189894
R10921 CS_BIAS.n1039 CS_BIAS.n1038 0.189894
R10922 CS_BIAS.n1039 CS_BIAS.n909 0.189894
R10923 CS_BIAS.n1043 CS_BIAS.n909 0.189894
R10924 CS_BIAS.n1044 CS_BIAS.n1043 0.189894
R10925 CS_BIAS.n1045 CS_BIAS.n1044 0.189894
R10926 CS_BIAS.n1045 CS_BIAS.n907 0.189894
R10927 CS_BIAS.n1049 CS_BIAS.n907 0.189894
R10928 CS_BIAS.n1073 CS_BIAS.n1070 0.189894
R10929 CS_BIAS.n1077 CS_BIAS.n1070 0.189894
R10930 CS_BIAS.n1078 CS_BIAS.n1077 0.189894
R10931 CS_BIAS.n1079 CS_BIAS.n1078 0.189894
R10932 CS_BIAS.n1079 CS_BIAS.n1068 0.189894
R10933 CS_BIAS.n1083 CS_BIAS.n1068 0.189894
R10934 CS_BIAS.n1084 CS_BIAS.n1083 0.189894
R10935 CS_BIAS.n1085 CS_BIAS.n1084 0.189894
R10936 CS_BIAS.n1085 CS_BIAS.n1066 0.189894
R10937 CS_BIAS.n1090 CS_BIAS.n1066 0.189894
R10938 CS_BIAS.n1091 CS_BIAS.n1090 0.189894
R10939 CS_BIAS.n1092 CS_BIAS.n1091 0.189894
R10940 CS_BIAS.n1092 CS_BIAS.n1064 0.189894
R10941 CS_BIAS.n1096 CS_BIAS.n1064 0.189894
R10942 CS_BIAS.n1097 CS_BIAS.n1096 0.189894
R10943 CS_BIAS.n1098 CS_BIAS.n1097 0.189894
R10944 CS_BIAS.n1098 CS_BIAS.n1062 0.189894
R10945 CS_BIAS.n1102 CS_BIAS.n1062 0.189894
R10946 CS_BIAS.n1103 CS_BIAS.n1102 0.189894
R10947 CS_BIAS.n1104 CS_BIAS.n1103 0.189894
R10948 CS_BIAS.n1104 CS_BIAS.n1060 0.189894
R10949 CS_BIAS.n1108 CS_BIAS.n1060 0.189894
R10950 CS_BIAS.n1109 CS_BIAS.n1108 0.189894
R10951 CS_BIAS.n1109 CS_BIAS.n1058 0.189894
R10952 CS_BIAS.n1113 CS_BIAS.n1058 0.189894
R10953 CS_BIAS.n1114 CS_BIAS.n1113 0.189894
R10954 CS_BIAS.n1115 CS_BIAS.n1114 0.189894
R10955 CS_BIAS.n1120 CS_BIAS.n1119 0.189894
R10956 CS_BIAS.n1121 CS_BIAS.n1120 0.189894
R10957 CS_BIAS.n1121 CS_BIAS.n901 0.189894
R10958 CS_BIAS.n1126 CS_BIAS.n901 0.189894
R10959 CS_BIAS.n1127 CS_BIAS.n1126 0.189894
R10960 CS_BIAS.n1128 CS_BIAS.n1127 0.189894
R10961 CS_BIAS.n1128 CS_BIAS.n899 0.189894
R10962 CS_BIAS.n1132 CS_BIAS.n899 0.189894
R10963 CS_BIAS.n1133 CS_BIAS.n1132 0.189894
R10964 CS_BIAS.n1134 CS_BIAS.n1133 0.189894
R10965 CS_BIAS.n1134 CS_BIAS.n897 0.189894
R10966 CS_BIAS.n1138 CS_BIAS.n897 0.189894
R10967 CS_BIAS.n1139 CS_BIAS.n1138 0.189894
R10968 CS_BIAS.n1140 CS_BIAS.n1139 0.189894
R10969 CS_BIAS.n1140 CS_BIAS.n895 0.189894
R10970 CS_BIAS.n1144 CS_BIAS.n895 0.189894
R10971 CS_BIAS.n1145 CS_BIAS.n1144 0.189894
R10972 CS_BIAS.n1145 CS_BIAS.n893 0.189894
R10973 CS_BIAS.n1149 CS_BIAS.n893 0.189894
R10974 CS_BIAS.n1150 CS_BIAS.n1149 0.189894
R10975 CS_BIAS.n1151 CS_BIAS.n1150 0.189894
R10976 CS_BIAS.n1151 CS_BIAS.n891 0.189894
R10977 CS_BIAS.n1155 CS_BIAS.n891 0.189894
R10978 CS_BIAS.n1156 CS_BIAS.n1155 0.189894
R10979 CS_BIAS.n1157 CS_BIAS.n1156 0.189894
R10980 CS_BIAS.n1157 CS_BIAS.n889 0.189894
R10981 CS_BIAS.n1161 CS_BIAS.n889 0.189894
R10982 CS_BIAS.n1162 CS_BIAS.n1161 0.189894
R10983 CS_BIAS.n1162 CS_BIAS.n887 0.189894
R10984 CS_BIAS.n1166 CS_BIAS.n887 0.189894
R10985 CS_BIAS.n1167 CS_BIAS.n1166 0.189894
R10986 CS_BIAS.n1168 CS_BIAS.n1167 0.189894
R10987 CS_BIAS.n1168 CS_BIAS.n885 0.189894
R10988 CS_BIAS.n1172 CS_BIAS.n885 0.189894
R10989 CS_BIAS.n1173 CS_BIAS.n1172 0.189894
R10990 CS_BIAS.n1174 CS_BIAS.n1173 0.189894
R10991 CS_BIAS.n1174 CS_BIAS.n883 0.189894
R10992 CS_BIAS.n1178 CS_BIAS.n883 0.189894
R10993 CS_BIAS.n234 CS_BIAS.n175 0.170955
R10994 CS_BIAS.n238 CS_BIAS.n175 0.170955
R10995 CS_BIAS.n1115 CS_BIAS.n1056 0.170955
R10996 CS_BIAS.n1119 CS_BIAS.n1056 0.170955
R10997 VOUT.n50 VOUT.n48 97.3561
R10998 VOUT.n44 VOUT.n42 97.3561
R10999 VOUT.n39 VOUT.n37 97.3561
R11000 VOUT.n13 VOUT.n11 97.3561
R11001 VOUT.n7 VOUT.n5 97.3561
R11002 VOUT.n2 VOUT.n0 97.3561
R11003 VOUT.n50 VOUT.n49 95.6607
R11004 VOUT.n46 VOUT.n45 95.6607
R11005 VOUT.n44 VOUT.n43 95.6607
R11006 VOUT.n41 VOUT.n40 95.6607
R11007 VOUT.n39 VOUT.n38 95.6607
R11008 VOUT.n13 VOUT.n12 95.6607
R11009 VOUT.n15 VOUT.n14 95.6607
R11010 VOUT.n7 VOUT.n6 95.6607
R11011 VOUT.n9 VOUT.n8 95.6607
R11012 VOUT.n2 VOUT.n1 95.6607
R11013 VOUT.n4 VOUT.n3 95.6607
R11014 VOUT.n52 VOUT.n51 95.6605
R11015 VOUT.n88 VOUT.n86 78.5929
R11016 VOUT.n80 VOUT.n78 78.5929
R11017 VOUT.n72 VOUT.n70 78.5929
R11018 VOUT.n64 VOUT.n62 78.5929
R11019 VOUT.n57 VOUT.n55 78.5929
R11020 VOUT.n128 VOUT.n126 78.5929
R11021 VOUT.n120 VOUT.n118 78.5929
R11022 VOUT.n112 VOUT.n110 78.5929
R11023 VOUT.n104 VOUT.n102 78.5929
R11024 VOUT.n97 VOUT.n95 78.5929
R11025 VOUT.n92 VOUT.n91 76.9579
R11026 VOUT.n90 VOUT.n89 76.9579
R11027 VOUT.n88 VOUT.n87 76.9579
R11028 VOUT.n84 VOUT.n83 76.9579
R11029 VOUT.n82 VOUT.n81 76.9579
R11030 VOUT.n80 VOUT.n79 76.9579
R11031 VOUT.n76 VOUT.n75 76.9579
R11032 VOUT.n74 VOUT.n73 76.9579
R11033 VOUT.n72 VOUT.n71 76.9579
R11034 VOUT.n68 VOUT.n67 76.9579
R11035 VOUT.n66 VOUT.n65 76.9579
R11036 VOUT.n64 VOUT.n63 76.9579
R11037 VOUT.n61 VOUT.n60 76.9579
R11038 VOUT.n59 VOUT.n58 76.9579
R11039 VOUT.n57 VOUT.n56 76.9579
R11040 VOUT.n128 VOUT.n127 76.9579
R11041 VOUT.n130 VOUT.n129 76.9579
R11042 VOUT.n132 VOUT.n131 76.9579
R11043 VOUT.n120 VOUT.n119 76.9579
R11044 VOUT.n122 VOUT.n121 76.9579
R11045 VOUT.n124 VOUT.n123 76.9579
R11046 VOUT.n112 VOUT.n111 76.9579
R11047 VOUT.n114 VOUT.n113 76.9579
R11048 VOUT.n116 VOUT.n115 76.9579
R11049 VOUT.n104 VOUT.n103 76.9579
R11050 VOUT.n106 VOUT.n105 76.9579
R11051 VOUT.n108 VOUT.n107 76.9579
R11052 VOUT.n97 VOUT.n96 76.9579
R11053 VOUT.n99 VOUT.n98 76.9579
R11054 VOUT.n101 VOUT.n100 76.9579
R11055 VOUT.n91 VOUT.t8 14.194
R11056 VOUT.n91 VOUT.t72 14.194
R11057 VOUT.n89 VOUT.t41 14.194
R11058 VOUT.n89 VOUT.t31 14.194
R11059 VOUT.n87 VOUT.t36 14.194
R11060 VOUT.n87 VOUT.t37 14.194
R11061 VOUT.n86 VOUT.t74 14.194
R11062 VOUT.n86 VOUT.t56 14.194
R11063 VOUT.n83 VOUT.t60 14.194
R11064 VOUT.n83 VOUT.t24 14.194
R11065 VOUT.n81 VOUT.t67 14.194
R11066 VOUT.n81 VOUT.t73 14.194
R11067 VOUT.n79 VOUT.t77 14.194
R11068 VOUT.n79 VOUT.t62 14.194
R11069 VOUT.n78 VOUT.t29 14.194
R11070 VOUT.n78 VOUT.t6 14.194
R11071 VOUT.n75 VOUT.t51 14.194
R11072 VOUT.n75 VOUT.t13 14.194
R11073 VOUT.n73 VOUT.t71 14.194
R11074 VOUT.n73 VOUT.t3 14.194
R11075 VOUT.n71 VOUT.t66 14.194
R11076 VOUT.n71 VOUT.t75 14.194
R11077 VOUT.n70 VOUT.t27 14.194
R11078 VOUT.n70 VOUT.t25 14.194
R11079 VOUT.n67 VOUT.t34 14.194
R11080 VOUT.n67 VOUT.t45 14.194
R11081 VOUT.n65 VOUT.t16 14.194
R11082 VOUT.n65 VOUT.t59 14.194
R11083 VOUT.n63 VOUT.t11 14.194
R11084 VOUT.n63 VOUT.t9 14.194
R11085 VOUT.n62 VOUT.t10 14.194
R11086 VOUT.n62 VOUT.t76 14.194
R11087 VOUT.n60 VOUT.t17 14.194
R11088 VOUT.n60 VOUT.t23 14.194
R11089 VOUT.n58 VOUT.t4 14.194
R11090 VOUT.n58 VOUT.t53 14.194
R11091 VOUT.n56 VOUT.t5 14.194
R11092 VOUT.n56 VOUT.t20 14.194
R11093 VOUT.n55 VOUT.t30 14.194
R11094 VOUT.n55 VOUT.t49 14.194
R11095 VOUT.n126 VOUT.t65 14.194
R11096 VOUT.n126 VOUT.t79 14.194
R11097 VOUT.n127 VOUT.t19 14.194
R11098 VOUT.n127 VOUT.t15 14.194
R11099 VOUT.n129 VOUT.t38 14.194
R11100 VOUT.n129 VOUT.t43 14.194
R11101 VOUT.n131 VOUT.t42 14.194
R11102 VOUT.n131 VOUT.t40 14.194
R11103 VOUT.n118 VOUT.t35 14.194
R11104 VOUT.n118 VOUT.t32 14.194
R11105 VOUT.n119 VOUT.t2 14.194
R11106 VOUT.n119 VOUT.t1 14.194
R11107 VOUT.n121 VOUT.t78 14.194
R11108 VOUT.n121 VOUT.t54 14.194
R11109 VOUT.n123 VOUT.t68 14.194
R11110 VOUT.n123 VOUT.t63 14.194
R11111 VOUT.n110 VOUT.t64 14.194
R11112 VOUT.n110 VOUT.t55 14.194
R11113 VOUT.n111 VOUT.t44 14.194
R11114 VOUT.n111 VOUT.t48 14.194
R11115 VOUT.n113 VOUT.t28 14.194
R11116 VOUT.n113 VOUT.t33 14.194
R11117 VOUT.n115 VOUT.t61 14.194
R11118 VOUT.n115 VOUT.t21 14.194
R11119 VOUT.n102 VOUT.t0 14.194
R11120 VOUT.n102 VOUT.t7 14.194
R11121 VOUT.n103 VOUT.t52 14.194
R11122 VOUT.n103 VOUT.t69 14.194
R11123 VOUT.n105 VOUT.t12 14.194
R11124 VOUT.n105 VOUT.t22 14.194
R11125 VOUT.n107 VOUT.t18 14.194
R11126 VOUT.n107 VOUT.t14 14.194
R11127 VOUT.n95 VOUT.t39 14.194
R11128 VOUT.n95 VOUT.t70 14.194
R11129 VOUT.n96 VOUT.t58 14.194
R11130 VOUT.n96 VOUT.t50 14.194
R11131 VOUT.n98 VOUT.t47 14.194
R11132 VOUT.n98 VOUT.t26 14.194
R11133 VOUT.n100 VOUT.t46 14.194
R11134 VOUT.n100 VOUT.t57 14.194
R11135 VOUT.n51 VOUT.t81 13.377
R11136 VOUT.n51 VOUT.t113 13.377
R11137 VOUT.n49 VOUT.t104 13.377
R11138 VOUT.n49 VOUT.t90 13.377
R11139 VOUT.n48 VOUT.t110 13.377
R11140 VOUT.n48 VOUT.t97 13.377
R11141 VOUT.n45 VOUT.t80 13.377
R11142 VOUT.n45 VOUT.t112 13.377
R11143 VOUT.n43 VOUT.t106 13.377
R11144 VOUT.n43 VOUT.t88 13.377
R11145 VOUT.n42 VOUT.t111 13.377
R11146 VOUT.n42 VOUT.t98 13.377
R11147 VOUT.n40 VOUT.t100 13.377
R11148 VOUT.n40 VOUT.t99 13.377
R11149 VOUT.n38 VOUT.t102 13.377
R11150 VOUT.n38 VOUT.t101 13.377
R11151 VOUT.n37 VOUT.t87 13.377
R11152 VOUT.n37 VOUT.t86 13.377
R11153 VOUT.n11 VOUT.t84 13.377
R11154 VOUT.n11 VOUT.t93 13.377
R11155 VOUT.n12 VOUT.t103 13.377
R11156 VOUT.n12 VOUT.t114 13.377
R11157 VOUT.n14 VOUT.t95 13.377
R11158 VOUT.n14 VOUT.t89 13.377
R11159 VOUT.n5 VOUT.t83 13.377
R11160 VOUT.n5 VOUT.t92 13.377
R11161 VOUT.n6 VOUT.t105 13.377
R11162 VOUT.n6 VOUT.t115 13.377
R11163 VOUT.n8 VOUT.t96 13.377
R11164 VOUT.n8 VOUT.t91 13.377
R11165 VOUT.n0 VOUT.t82 13.377
R11166 VOUT.n0 VOUT.t85 13.377
R11167 VOUT.n1 VOUT.t108 13.377
R11168 VOUT.n1 VOUT.t109 13.377
R11169 VOUT.n3 VOUT.t94 13.377
R11170 VOUT.n3 VOUT.t107 13.377
R11171 VOUT.n94 VOUT.n54 8.85259
R11172 VOUT.n47 VOUT.n41 6.84892
R11173 VOUT.n10 VOUT.n4 6.84892
R11174 VOUT.n69 VOUT.n61 6.52205
R11175 VOUT.n109 VOUT.n101 6.52205
R11176 VOUT.n134 VOUT.n94 6.49684
R11177 VOUT.n54 VOUT.n17 6.01681
R11178 VOUT.n53 VOUT.n52 5.65855
R11179 VOUT.n47 VOUT.n46 5.65855
R11180 VOUT.n16 VOUT.n15 5.65855
R11181 VOUT.n10 VOUT.n9 5.65855
R11182 VOUT.n93 VOUT.n92 5.62837
R11183 VOUT.n85 VOUT.n84 5.62837
R11184 VOUT.n77 VOUT.n76 5.62837
R11185 VOUT.n69 VOUT.n68 5.62837
R11186 VOUT.n133 VOUT.n132 5.62837
R11187 VOUT.n125 VOUT.n124 5.62837
R11188 VOUT.n117 VOUT.n116 5.62837
R11189 VOUT.n109 VOUT.n108 5.62837
R11190 VOUT.n135 VOUT.n17 5.11648
R11191 VOUT.n54 VOUT.n53 4.83004
R11192 VOUT.n17 VOUT.n16 4.83004
R11193 VOUT.n94 VOUT.n93 4.24958
R11194 VOUT.n134 VOUT.n133 4.24958
R11195 VOUT.n36 VOUT 3.9673
R11196 VOUT.n135 VOUT.n134 3.7171
R11197 VOUT.n52 VOUT.n50 1.6959
R11198 VOUT.n46 VOUT.n44 1.6959
R11199 VOUT.n41 VOUT.n39 1.6959
R11200 VOUT.n15 VOUT.n13 1.6959
R11201 VOUT.n9 VOUT.n7 1.6959
R11202 VOUT.n4 VOUT.n2 1.6959
R11203 VOUT.n90 VOUT.n88 1.63556
R11204 VOUT.n92 VOUT.n90 1.63556
R11205 VOUT.n82 VOUT.n80 1.63556
R11206 VOUT.n84 VOUT.n82 1.63556
R11207 VOUT.n74 VOUT.n72 1.63556
R11208 VOUT.n76 VOUT.n74 1.63556
R11209 VOUT.n66 VOUT.n64 1.63556
R11210 VOUT.n68 VOUT.n66 1.63556
R11211 VOUT.n59 VOUT.n57 1.63556
R11212 VOUT.n61 VOUT.n59 1.63556
R11213 VOUT.n132 VOUT.n130 1.63556
R11214 VOUT.n130 VOUT.n128 1.63556
R11215 VOUT.n124 VOUT.n122 1.63556
R11216 VOUT.n122 VOUT.n120 1.63556
R11217 VOUT.n116 VOUT.n114 1.63556
R11218 VOUT.n114 VOUT.n112 1.63556
R11219 VOUT.n108 VOUT.n106 1.63556
R11220 VOUT.n106 VOUT.n104 1.63556
R11221 VOUT.n101 VOUT.n99 1.63556
R11222 VOUT.n99 VOUT.n97 1.63556
R11223 VOUT.n53 VOUT.n47 1.19087
R11224 VOUT.n16 VOUT.n10 1.19087
R11225 VOUT.n93 VOUT.n85 0.894178
R11226 VOUT.n85 VOUT.n77 0.894178
R11227 VOUT.n77 VOUT.n69 0.894178
R11228 VOUT.n133 VOUT.n125 0.894178
R11229 VOUT.n125 VOUT.n117 0.894178
R11230 VOUT.n117 VOUT.n109 0.894178
R11231 VOUT.n36 VOUT.n35 0.389516
R11232 VOUT.n135 VOUT.n36 0.38778
R11233 VOUT.n28 VOUT.n27 0.0802186
R11234 VOUT.n30 VOUT.n29 0.0780158
R11235 VOUT.n22 VOUT.n21 0.077577
R11236 VOUT.n25 VOUT.n24 0.0732383
R11237 VOUT.n32 VOUT.n31 0.0732383
R11238 VOUT.n34 VOUT.n33 0.0732383
R11239 VOUT.n29 VOUT.n28 0.0704532
R11240 VOUT.n21 VOUT.n18 0.0460297
R11241 VOUT.n26 VOUT.n20 0.0391444
R11242 VOUT.n23 VOUT.n19 0.0391444
R11243 VOUT.n22 VOUT.t121 0.0335236
R11244 VOUT.n25 VOUT.t118 0.0335236
R11245 VOUT.n31 VOUT.t116 0.0335236
R11246 VOUT.n33 VOUT.t117 0.0335236
R11247 VOUT.n35 VOUT.t119 0.0335236
R11248 VOUT.n24 VOUT.t121 0.0293356
R11249 VOUT.n27 VOUT.t118 0.0293356
R11250 VOUT.t116 VOUT.n30 0.0293356
R11251 VOUT.t117 VOUT.n32 0.0293356
R11252 VOUT.t119 VOUT.n34 0.0293356
R11253 VOUT.n28 VOUT.t122 0.0173498
R11254 VOUT.n29 VOUT.t120 0.0172226
R11255 VOUT.n21 VOUT.t123 0.0166115
R11256 VOUT.n23 VOUT.n22 0.0164414
R11257 VOUT.n26 VOUT.n25 0.0164414
R11258 VOUT.n31 VOUT.n20 0.0164414
R11259 VOUT.n33 VOUT.n19 0.0164414
R11260 VOUT.n35 VOUT.n18 0.0164414
R11261 VOUT.n24 VOUT.n23 0.012294
R11262 VOUT.n27 VOUT.n26 0.012294
R11263 VOUT.n30 VOUT.n20 0.012294
R11264 VOUT.n32 VOUT.n19 0.012294
R11265 VOUT.n34 VOUT.n18 0.012294
R11266 VOUT VOUT.n135 0.0099
R11267 GND.n8498 GND.n8497 1357.48
R11268 GND.n8363 GND.n8362 1208.66
R11269 GND.n9528 GND.n571 1072.94
R11270 GND.n10134 GND.n418 754.366
R11271 GND.n10076 GND.n416 754.366
R11272 GND.n6417 GND.n6387 754.366
R11273 GND.n6361 GND.n4886 754.366
R11274 GND.n2926 GND.n1359 754.366
R11275 GND.n8025 GND.n8024 754.366
R11276 GND.n1454 GND.n1357 754.366
R11277 GND.n1706 GND.n1678 754.366
R11278 GND.n10136 GND.n414 742.355
R11279 GND.n10038 GND.n415 742.355
R11280 GND.n6415 GND.n4868 742.355
R11281 GND.n7181 GND.n4878 742.355
R11282 GND.n8022 GND.n1677 742.355
R11283 GND.n8027 GND.n1675 742.355
R11284 GND.n2929 GND.n1351 742.355
R11285 GND.n8360 GND.n1362 742.355
R11286 GND.n8496 GND.n1187 723.135
R11287 GND.n9527 GND.n572 723.135
R11288 GND.n9696 GND.n9695 723.135
R11289 GND.n8364 GND.n1321 723.135
R11290 GND.n6314 GND.n6313 687.098
R11291 GND.n7410 GND.n4416 687.098
R11292 GND.n7698 GND.n2340 687.098
R11293 GND.n7757 GND.n2344 687.098
R11294 GND.n6362 GND.n6361 589.749
R11295 GND.n8024 GND.n1682 589.749
R11296 GND.n3873 GND.n1706 588.312
R11297 GND.n6387 GND.n6386 588.312
R11298 GND.n8496 GND.n8495 585
R11299 GND.n8497 GND.n8496 585
R11300 GND.n8494 GND.n1189 585
R11301 GND.n1189 GND.n1188 585
R11302 GND.n8493 GND.n8492 585
R11303 GND.n8492 GND.n8491 585
R11304 GND.n1194 GND.n1193 585
R11305 GND.n8490 GND.n1194 585
R11306 GND.n8488 GND.n8487 585
R11307 GND.n8489 GND.n8488 585
R11308 GND.n8486 GND.n1196 585
R11309 GND.n1196 GND.n1195 585
R11310 GND.n8485 GND.n8484 585
R11311 GND.n8484 GND.n8483 585
R11312 GND.n1202 GND.n1201 585
R11313 GND.n8482 GND.n1202 585
R11314 GND.n8480 GND.n8479 585
R11315 GND.n8481 GND.n8480 585
R11316 GND.n8478 GND.n1204 585
R11317 GND.n1204 GND.n1203 585
R11318 GND.n8477 GND.n8476 585
R11319 GND.n8476 GND.n8475 585
R11320 GND.n1210 GND.n1209 585
R11321 GND.n8474 GND.n1210 585
R11322 GND.n8472 GND.n8471 585
R11323 GND.n8473 GND.n8472 585
R11324 GND.n8470 GND.n1212 585
R11325 GND.n1212 GND.n1211 585
R11326 GND.n8469 GND.n8468 585
R11327 GND.n8468 GND.n8467 585
R11328 GND.n1218 GND.n1217 585
R11329 GND.n8466 GND.n1218 585
R11330 GND.n8464 GND.n8463 585
R11331 GND.n8465 GND.n8464 585
R11332 GND.n8462 GND.n1220 585
R11333 GND.n1220 GND.n1219 585
R11334 GND.n8461 GND.n8460 585
R11335 GND.n8460 GND.n8459 585
R11336 GND.n1226 GND.n1225 585
R11337 GND.n8458 GND.n1226 585
R11338 GND.n8456 GND.n8455 585
R11339 GND.n8457 GND.n8456 585
R11340 GND.n8454 GND.n1228 585
R11341 GND.n1228 GND.n1227 585
R11342 GND.n8453 GND.n8452 585
R11343 GND.n8452 GND.n8451 585
R11344 GND.n1234 GND.n1233 585
R11345 GND.n8450 GND.n1234 585
R11346 GND.n8448 GND.n8447 585
R11347 GND.n8449 GND.n8448 585
R11348 GND.n8446 GND.n1236 585
R11349 GND.n1236 GND.n1235 585
R11350 GND.n8445 GND.n8444 585
R11351 GND.n8444 GND.n8443 585
R11352 GND.n1242 GND.n1241 585
R11353 GND.n8442 GND.n1242 585
R11354 GND.n8440 GND.n8439 585
R11355 GND.n8441 GND.n8440 585
R11356 GND.n8438 GND.n1244 585
R11357 GND.n1244 GND.n1243 585
R11358 GND.n8437 GND.n8436 585
R11359 GND.n8436 GND.n8435 585
R11360 GND.n1250 GND.n1249 585
R11361 GND.n8434 GND.n1250 585
R11362 GND.n8432 GND.n8431 585
R11363 GND.n8433 GND.n8432 585
R11364 GND.n8430 GND.n1252 585
R11365 GND.n1252 GND.n1251 585
R11366 GND.n8429 GND.n8428 585
R11367 GND.n8428 GND.n8427 585
R11368 GND.n1258 GND.n1257 585
R11369 GND.n8426 GND.n1258 585
R11370 GND.n8424 GND.n8423 585
R11371 GND.n8425 GND.n8424 585
R11372 GND.n8422 GND.n1260 585
R11373 GND.n1260 GND.n1259 585
R11374 GND.n8421 GND.n8420 585
R11375 GND.n8420 GND.n8419 585
R11376 GND.n1266 GND.n1265 585
R11377 GND.n8418 GND.n1266 585
R11378 GND.n8416 GND.n8415 585
R11379 GND.n8417 GND.n8416 585
R11380 GND.n8414 GND.n1268 585
R11381 GND.n1268 GND.n1267 585
R11382 GND.n8413 GND.n8412 585
R11383 GND.n8412 GND.n8411 585
R11384 GND.n1274 GND.n1273 585
R11385 GND.n8410 GND.n1274 585
R11386 GND.n8408 GND.n8407 585
R11387 GND.n8409 GND.n8408 585
R11388 GND.n8406 GND.n1276 585
R11389 GND.n1276 GND.n1275 585
R11390 GND.n8405 GND.n8404 585
R11391 GND.n8404 GND.n8403 585
R11392 GND.n1282 GND.n1281 585
R11393 GND.n8402 GND.n1282 585
R11394 GND.n8400 GND.n8399 585
R11395 GND.n8401 GND.n8400 585
R11396 GND.n8398 GND.n1284 585
R11397 GND.n1284 GND.n1283 585
R11398 GND.n8397 GND.n8396 585
R11399 GND.n8396 GND.n8395 585
R11400 GND.n1290 GND.n1289 585
R11401 GND.n8394 GND.n1290 585
R11402 GND.n8392 GND.n8391 585
R11403 GND.n8393 GND.n8392 585
R11404 GND.n8390 GND.n1292 585
R11405 GND.n1292 GND.n1291 585
R11406 GND.n8389 GND.n8388 585
R11407 GND.n8388 GND.n8387 585
R11408 GND.n1298 GND.n1297 585
R11409 GND.n8386 GND.n1298 585
R11410 GND.n8384 GND.n8383 585
R11411 GND.n8385 GND.n8384 585
R11412 GND.n8382 GND.n1300 585
R11413 GND.n1300 GND.n1299 585
R11414 GND.n8381 GND.n8380 585
R11415 GND.n8380 GND.n8379 585
R11416 GND.n1306 GND.n1305 585
R11417 GND.n8378 GND.n1306 585
R11418 GND.n8376 GND.n8375 585
R11419 GND.n8377 GND.n8376 585
R11420 GND.n8374 GND.n1308 585
R11421 GND.n1308 GND.n1307 585
R11422 GND.n8373 GND.n8372 585
R11423 GND.n8372 GND.n8371 585
R11424 GND.n1314 GND.n1313 585
R11425 GND.n8370 GND.n1314 585
R11426 GND.n8368 GND.n8367 585
R11427 GND.n8369 GND.n8368 585
R11428 GND.n8366 GND.n1316 585
R11429 GND.n1316 GND.n1315 585
R11430 GND.n8365 GND.n8364 585
R11431 GND.n8364 GND.n8363 585
R11432 GND.n1187 GND.n1186 585
R11433 GND.n8498 GND.n1187 585
R11434 GND.n8501 GND.n8500 585
R11435 GND.n8500 GND.n8499 585
R11436 GND.n1184 GND.n1183 585
R11437 GND.n1183 GND.n1182 585
R11438 GND.n8506 GND.n8505 585
R11439 GND.n8507 GND.n8506 585
R11440 GND.n1181 GND.n1180 585
R11441 GND.n8508 GND.n1181 585
R11442 GND.n8511 GND.n8510 585
R11443 GND.n8510 GND.n8509 585
R11444 GND.n1178 GND.n1177 585
R11445 GND.n1177 GND.n1176 585
R11446 GND.n8516 GND.n8515 585
R11447 GND.n8517 GND.n8516 585
R11448 GND.n1175 GND.n1174 585
R11449 GND.n8518 GND.n1175 585
R11450 GND.n8521 GND.n8520 585
R11451 GND.n8520 GND.n8519 585
R11452 GND.n1172 GND.n1171 585
R11453 GND.n1171 GND.n1170 585
R11454 GND.n8526 GND.n8525 585
R11455 GND.n8527 GND.n8526 585
R11456 GND.n1169 GND.n1168 585
R11457 GND.n8528 GND.n1169 585
R11458 GND.n8531 GND.n8530 585
R11459 GND.n8530 GND.n8529 585
R11460 GND.n1166 GND.n1165 585
R11461 GND.n1165 GND.n1164 585
R11462 GND.n8536 GND.n8535 585
R11463 GND.n8537 GND.n8536 585
R11464 GND.n1163 GND.n1162 585
R11465 GND.n8538 GND.n1163 585
R11466 GND.n8541 GND.n8540 585
R11467 GND.n8540 GND.n8539 585
R11468 GND.n1160 GND.n1159 585
R11469 GND.n1159 GND.n1158 585
R11470 GND.n8546 GND.n8545 585
R11471 GND.n8547 GND.n8546 585
R11472 GND.n1157 GND.n1156 585
R11473 GND.n8548 GND.n1157 585
R11474 GND.n8551 GND.n8550 585
R11475 GND.n8550 GND.n8549 585
R11476 GND.n1154 GND.n1153 585
R11477 GND.n1153 GND.n1152 585
R11478 GND.n8556 GND.n8555 585
R11479 GND.n8557 GND.n8556 585
R11480 GND.n1151 GND.n1150 585
R11481 GND.n8558 GND.n1151 585
R11482 GND.n8561 GND.n8560 585
R11483 GND.n8560 GND.n8559 585
R11484 GND.n1148 GND.n1147 585
R11485 GND.n1147 GND.n1146 585
R11486 GND.n8566 GND.n8565 585
R11487 GND.n8567 GND.n8566 585
R11488 GND.n1145 GND.n1144 585
R11489 GND.n8568 GND.n1145 585
R11490 GND.n8571 GND.n8570 585
R11491 GND.n8570 GND.n8569 585
R11492 GND.n1142 GND.n1141 585
R11493 GND.n1141 GND.n1140 585
R11494 GND.n8576 GND.n8575 585
R11495 GND.n8577 GND.n8576 585
R11496 GND.n1139 GND.n1138 585
R11497 GND.n8578 GND.n1139 585
R11498 GND.n8581 GND.n8580 585
R11499 GND.n8580 GND.n8579 585
R11500 GND.n1136 GND.n1135 585
R11501 GND.n1135 GND.n1134 585
R11502 GND.n8586 GND.n8585 585
R11503 GND.n8587 GND.n8586 585
R11504 GND.n1133 GND.n1132 585
R11505 GND.n8588 GND.n1133 585
R11506 GND.n8591 GND.n8590 585
R11507 GND.n8590 GND.n8589 585
R11508 GND.n1130 GND.n1129 585
R11509 GND.n1129 GND.n1128 585
R11510 GND.n8596 GND.n8595 585
R11511 GND.n8597 GND.n8596 585
R11512 GND.n1127 GND.n1126 585
R11513 GND.n8598 GND.n1127 585
R11514 GND.n8601 GND.n8600 585
R11515 GND.n8600 GND.n8599 585
R11516 GND.n1124 GND.n1123 585
R11517 GND.n1123 GND.n1122 585
R11518 GND.n8606 GND.n8605 585
R11519 GND.n8607 GND.n8606 585
R11520 GND.n1121 GND.n1120 585
R11521 GND.n8608 GND.n1121 585
R11522 GND.n8611 GND.n8610 585
R11523 GND.n8610 GND.n8609 585
R11524 GND.n1118 GND.n1117 585
R11525 GND.n1117 GND.n1116 585
R11526 GND.n8616 GND.n8615 585
R11527 GND.n8617 GND.n8616 585
R11528 GND.n1115 GND.n1114 585
R11529 GND.n8618 GND.n1115 585
R11530 GND.n8621 GND.n8620 585
R11531 GND.n8620 GND.n8619 585
R11532 GND.n1112 GND.n1111 585
R11533 GND.n1111 GND.n1110 585
R11534 GND.n8626 GND.n8625 585
R11535 GND.n8627 GND.n8626 585
R11536 GND.n1109 GND.n1108 585
R11537 GND.n8628 GND.n1109 585
R11538 GND.n8631 GND.n8630 585
R11539 GND.n8630 GND.n8629 585
R11540 GND.n1106 GND.n1105 585
R11541 GND.n1105 GND.n1104 585
R11542 GND.n8636 GND.n8635 585
R11543 GND.n8637 GND.n8636 585
R11544 GND.n1103 GND.n1102 585
R11545 GND.n8638 GND.n1103 585
R11546 GND.n8641 GND.n8640 585
R11547 GND.n8640 GND.n8639 585
R11548 GND.n1100 GND.n1099 585
R11549 GND.n1099 GND.n1098 585
R11550 GND.n8646 GND.n8645 585
R11551 GND.n8647 GND.n8646 585
R11552 GND.n1097 GND.n1096 585
R11553 GND.n8648 GND.n1097 585
R11554 GND.n8651 GND.n8650 585
R11555 GND.n8650 GND.n8649 585
R11556 GND.n1094 GND.n1093 585
R11557 GND.n1093 GND.n1092 585
R11558 GND.n8656 GND.n8655 585
R11559 GND.n8657 GND.n8656 585
R11560 GND.n1091 GND.n1090 585
R11561 GND.n8658 GND.n1091 585
R11562 GND.n8661 GND.n8660 585
R11563 GND.n8660 GND.n8659 585
R11564 GND.n1088 GND.n1087 585
R11565 GND.n1087 GND.n1086 585
R11566 GND.n8666 GND.n8665 585
R11567 GND.n8667 GND.n8666 585
R11568 GND.n1085 GND.n1084 585
R11569 GND.n8668 GND.n1085 585
R11570 GND.n8671 GND.n8670 585
R11571 GND.n8670 GND.n8669 585
R11572 GND.n1082 GND.n1081 585
R11573 GND.n1081 GND.n1080 585
R11574 GND.n8676 GND.n8675 585
R11575 GND.n8677 GND.n8676 585
R11576 GND.n1079 GND.n1078 585
R11577 GND.n8678 GND.n1079 585
R11578 GND.n8681 GND.n8680 585
R11579 GND.n8680 GND.n8679 585
R11580 GND.n1076 GND.n1075 585
R11581 GND.n1075 GND.n1074 585
R11582 GND.n8686 GND.n8685 585
R11583 GND.n8687 GND.n8686 585
R11584 GND.n1073 GND.n1072 585
R11585 GND.n8688 GND.n1073 585
R11586 GND.n8691 GND.n8690 585
R11587 GND.n8690 GND.n8689 585
R11588 GND.n1070 GND.n1069 585
R11589 GND.n1069 GND.n1068 585
R11590 GND.n8696 GND.n8695 585
R11591 GND.n8697 GND.n8696 585
R11592 GND.n1067 GND.n1066 585
R11593 GND.n8698 GND.n1067 585
R11594 GND.n8701 GND.n8700 585
R11595 GND.n8700 GND.n8699 585
R11596 GND.n1064 GND.n1063 585
R11597 GND.n1063 GND.n1062 585
R11598 GND.n8706 GND.n8705 585
R11599 GND.n8707 GND.n8706 585
R11600 GND.n1061 GND.n1060 585
R11601 GND.n8708 GND.n1061 585
R11602 GND.n8711 GND.n8710 585
R11603 GND.n8710 GND.n8709 585
R11604 GND.n1058 GND.n1057 585
R11605 GND.n1057 GND.n1056 585
R11606 GND.n8716 GND.n8715 585
R11607 GND.n8717 GND.n8716 585
R11608 GND.n1055 GND.n1054 585
R11609 GND.n8718 GND.n1055 585
R11610 GND.n8721 GND.n8720 585
R11611 GND.n8720 GND.n8719 585
R11612 GND.n1052 GND.n1051 585
R11613 GND.n1051 GND.n1050 585
R11614 GND.n8726 GND.n8725 585
R11615 GND.n8727 GND.n8726 585
R11616 GND.n1049 GND.n1048 585
R11617 GND.n8728 GND.n1049 585
R11618 GND.n8731 GND.n8730 585
R11619 GND.n8730 GND.n8729 585
R11620 GND.n1046 GND.n1045 585
R11621 GND.n1045 GND.n1044 585
R11622 GND.n8736 GND.n8735 585
R11623 GND.n8737 GND.n8736 585
R11624 GND.n1043 GND.n1042 585
R11625 GND.n8738 GND.n1043 585
R11626 GND.n8741 GND.n8740 585
R11627 GND.n8740 GND.n8739 585
R11628 GND.n1040 GND.n1039 585
R11629 GND.n1039 GND.n1038 585
R11630 GND.n8746 GND.n8745 585
R11631 GND.n8747 GND.n8746 585
R11632 GND.n1037 GND.n1036 585
R11633 GND.n8748 GND.n1037 585
R11634 GND.n8751 GND.n8750 585
R11635 GND.n8750 GND.n8749 585
R11636 GND.n1034 GND.n1033 585
R11637 GND.n1033 GND.n1032 585
R11638 GND.n8756 GND.n8755 585
R11639 GND.n8757 GND.n8756 585
R11640 GND.n1031 GND.n1030 585
R11641 GND.n8758 GND.n1031 585
R11642 GND.n8761 GND.n8760 585
R11643 GND.n8760 GND.n8759 585
R11644 GND.n1028 GND.n1027 585
R11645 GND.n1027 GND.n1026 585
R11646 GND.n8766 GND.n8765 585
R11647 GND.n8767 GND.n8766 585
R11648 GND.n1025 GND.n1024 585
R11649 GND.n8768 GND.n1025 585
R11650 GND.n8771 GND.n8770 585
R11651 GND.n8770 GND.n8769 585
R11652 GND.n1022 GND.n1021 585
R11653 GND.n1021 GND.n1020 585
R11654 GND.n8776 GND.n8775 585
R11655 GND.n8777 GND.n8776 585
R11656 GND.n1019 GND.n1018 585
R11657 GND.n8778 GND.n1019 585
R11658 GND.n8781 GND.n8780 585
R11659 GND.n8780 GND.n8779 585
R11660 GND.n1016 GND.n1015 585
R11661 GND.n1015 GND.n1014 585
R11662 GND.n8786 GND.n8785 585
R11663 GND.n8787 GND.n8786 585
R11664 GND.n1013 GND.n1012 585
R11665 GND.n8788 GND.n1013 585
R11666 GND.n8791 GND.n8790 585
R11667 GND.n8790 GND.n8789 585
R11668 GND.n1010 GND.n1009 585
R11669 GND.n1009 GND.n1008 585
R11670 GND.n8796 GND.n8795 585
R11671 GND.n8797 GND.n8796 585
R11672 GND.n1007 GND.n1006 585
R11673 GND.n8798 GND.n1007 585
R11674 GND.n8801 GND.n8800 585
R11675 GND.n8800 GND.n8799 585
R11676 GND.n1004 GND.n1003 585
R11677 GND.n1003 GND.n1002 585
R11678 GND.n8806 GND.n8805 585
R11679 GND.n8807 GND.n8806 585
R11680 GND.n1001 GND.n1000 585
R11681 GND.n8808 GND.n1001 585
R11682 GND.n8811 GND.n8810 585
R11683 GND.n8810 GND.n8809 585
R11684 GND.n998 GND.n997 585
R11685 GND.n997 GND.n996 585
R11686 GND.n8816 GND.n8815 585
R11687 GND.n8817 GND.n8816 585
R11688 GND.n995 GND.n994 585
R11689 GND.n8818 GND.n995 585
R11690 GND.n8821 GND.n8820 585
R11691 GND.n8820 GND.n8819 585
R11692 GND.n992 GND.n991 585
R11693 GND.n991 GND.n990 585
R11694 GND.n8826 GND.n8825 585
R11695 GND.n8827 GND.n8826 585
R11696 GND.n989 GND.n988 585
R11697 GND.n8828 GND.n989 585
R11698 GND.n8831 GND.n8830 585
R11699 GND.n8830 GND.n8829 585
R11700 GND.n986 GND.n985 585
R11701 GND.n985 GND.n984 585
R11702 GND.n8836 GND.n8835 585
R11703 GND.n8837 GND.n8836 585
R11704 GND.n983 GND.n982 585
R11705 GND.n8838 GND.n983 585
R11706 GND.n8841 GND.n8840 585
R11707 GND.n8840 GND.n8839 585
R11708 GND.n980 GND.n979 585
R11709 GND.n979 GND.n978 585
R11710 GND.n8846 GND.n8845 585
R11711 GND.n8847 GND.n8846 585
R11712 GND.n977 GND.n976 585
R11713 GND.n8848 GND.n977 585
R11714 GND.n8851 GND.n8850 585
R11715 GND.n8850 GND.n8849 585
R11716 GND.n974 GND.n973 585
R11717 GND.n973 GND.n972 585
R11718 GND.n8856 GND.n8855 585
R11719 GND.n8857 GND.n8856 585
R11720 GND.n971 GND.n970 585
R11721 GND.n8858 GND.n971 585
R11722 GND.n8861 GND.n8860 585
R11723 GND.n8860 GND.n8859 585
R11724 GND.n968 GND.n967 585
R11725 GND.n967 GND.n966 585
R11726 GND.n8866 GND.n8865 585
R11727 GND.n8867 GND.n8866 585
R11728 GND.n965 GND.n964 585
R11729 GND.n8868 GND.n965 585
R11730 GND.n8871 GND.n8870 585
R11731 GND.n8870 GND.n8869 585
R11732 GND.n962 GND.n961 585
R11733 GND.n961 GND.n960 585
R11734 GND.n8876 GND.n8875 585
R11735 GND.n8877 GND.n8876 585
R11736 GND.n959 GND.n958 585
R11737 GND.n8878 GND.n959 585
R11738 GND.n8881 GND.n8880 585
R11739 GND.n8880 GND.n8879 585
R11740 GND.n956 GND.n955 585
R11741 GND.n955 GND.n954 585
R11742 GND.n8886 GND.n8885 585
R11743 GND.n8887 GND.n8886 585
R11744 GND.n953 GND.n952 585
R11745 GND.n8888 GND.n953 585
R11746 GND.n8891 GND.n8890 585
R11747 GND.n8890 GND.n8889 585
R11748 GND.n950 GND.n949 585
R11749 GND.n949 GND.n948 585
R11750 GND.n8896 GND.n8895 585
R11751 GND.n8897 GND.n8896 585
R11752 GND.n947 GND.n946 585
R11753 GND.n8898 GND.n947 585
R11754 GND.n8901 GND.n8900 585
R11755 GND.n8900 GND.n8899 585
R11756 GND.n944 GND.n943 585
R11757 GND.n943 GND.n942 585
R11758 GND.n8906 GND.n8905 585
R11759 GND.n8907 GND.n8906 585
R11760 GND.n941 GND.n940 585
R11761 GND.n8908 GND.n941 585
R11762 GND.n8911 GND.n8910 585
R11763 GND.n8910 GND.n8909 585
R11764 GND.n938 GND.n937 585
R11765 GND.n937 GND.n936 585
R11766 GND.n8916 GND.n8915 585
R11767 GND.n8917 GND.n8916 585
R11768 GND.n935 GND.n934 585
R11769 GND.n8918 GND.n935 585
R11770 GND.n8921 GND.n8920 585
R11771 GND.n8920 GND.n8919 585
R11772 GND.n932 GND.n931 585
R11773 GND.n931 GND.n930 585
R11774 GND.n8926 GND.n8925 585
R11775 GND.n8927 GND.n8926 585
R11776 GND.n929 GND.n928 585
R11777 GND.n8928 GND.n929 585
R11778 GND.n8931 GND.n8930 585
R11779 GND.n8930 GND.n8929 585
R11780 GND.n926 GND.n925 585
R11781 GND.n925 GND.n924 585
R11782 GND.n8936 GND.n8935 585
R11783 GND.n8937 GND.n8936 585
R11784 GND.n923 GND.n922 585
R11785 GND.n8938 GND.n923 585
R11786 GND.n8941 GND.n8940 585
R11787 GND.n8940 GND.n8939 585
R11788 GND.n920 GND.n919 585
R11789 GND.n919 GND.n918 585
R11790 GND.n8946 GND.n8945 585
R11791 GND.n8947 GND.n8946 585
R11792 GND.n917 GND.n916 585
R11793 GND.n8948 GND.n917 585
R11794 GND.n8951 GND.n8950 585
R11795 GND.n8950 GND.n8949 585
R11796 GND.n914 GND.n913 585
R11797 GND.n913 GND.n912 585
R11798 GND.n8956 GND.n8955 585
R11799 GND.n8957 GND.n8956 585
R11800 GND.n911 GND.n910 585
R11801 GND.n8958 GND.n911 585
R11802 GND.n8961 GND.n8960 585
R11803 GND.n8960 GND.n8959 585
R11804 GND.n908 GND.n907 585
R11805 GND.n907 GND.n906 585
R11806 GND.n8966 GND.n8965 585
R11807 GND.n8967 GND.n8966 585
R11808 GND.n905 GND.n904 585
R11809 GND.n8968 GND.n905 585
R11810 GND.n8971 GND.n8970 585
R11811 GND.n8970 GND.n8969 585
R11812 GND.n902 GND.n901 585
R11813 GND.n901 GND.n900 585
R11814 GND.n8976 GND.n8975 585
R11815 GND.n8977 GND.n8976 585
R11816 GND.n899 GND.n898 585
R11817 GND.n8978 GND.n899 585
R11818 GND.n8981 GND.n8980 585
R11819 GND.n8980 GND.n8979 585
R11820 GND.n896 GND.n895 585
R11821 GND.n895 GND.n894 585
R11822 GND.n8986 GND.n8985 585
R11823 GND.n8987 GND.n8986 585
R11824 GND.n893 GND.n892 585
R11825 GND.n8988 GND.n893 585
R11826 GND.n8991 GND.n8990 585
R11827 GND.n8990 GND.n8989 585
R11828 GND.n890 GND.n889 585
R11829 GND.n889 GND.n888 585
R11830 GND.n8996 GND.n8995 585
R11831 GND.n8997 GND.n8996 585
R11832 GND.n887 GND.n886 585
R11833 GND.n8998 GND.n887 585
R11834 GND.n9001 GND.n9000 585
R11835 GND.n9000 GND.n8999 585
R11836 GND.n884 GND.n883 585
R11837 GND.n883 GND.n882 585
R11838 GND.n9006 GND.n9005 585
R11839 GND.n9007 GND.n9006 585
R11840 GND.n881 GND.n880 585
R11841 GND.n9008 GND.n881 585
R11842 GND.n9011 GND.n9010 585
R11843 GND.n9010 GND.n9009 585
R11844 GND.n878 GND.n877 585
R11845 GND.n877 GND.n876 585
R11846 GND.n9016 GND.n9015 585
R11847 GND.n9017 GND.n9016 585
R11848 GND.n875 GND.n874 585
R11849 GND.n9018 GND.n875 585
R11850 GND.n9021 GND.n9020 585
R11851 GND.n9020 GND.n9019 585
R11852 GND.n872 GND.n871 585
R11853 GND.n871 GND.n870 585
R11854 GND.n9026 GND.n9025 585
R11855 GND.n9027 GND.n9026 585
R11856 GND.n869 GND.n868 585
R11857 GND.n9028 GND.n869 585
R11858 GND.n9031 GND.n9030 585
R11859 GND.n9030 GND.n9029 585
R11860 GND.n866 GND.n865 585
R11861 GND.n865 GND.n864 585
R11862 GND.n9036 GND.n9035 585
R11863 GND.n9037 GND.n9036 585
R11864 GND.n863 GND.n862 585
R11865 GND.n9038 GND.n863 585
R11866 GND.n9041 GND.n9040 585
R11867 GND.n9040 GND.n9039 585
R11868 GND.n860 GND.n859 585
R11869 GND.n859 GND.n858 585
R11870 GND.n9046 GND.n9045 585
R11871 GND.n9047 GND.n9046 585
R11872 GND.n857 GND.n856 585
R11873 GND.n9048 GND.n857 585
R11874 GND.n9051 GND.n9050 585
R11875 GND.n9050 GND.n9049 585
R11876 GND.n854 GND.n853 585
R11877 GND.n853 GND.n852 585
R11878 GND.n9056 GND.n9055 585
R11879 GND.n9057 GND.n9056 585
R11880 GND.n851 GND.n850 585
R11881 GND.n9058 GND.n851 585
R11882 GND.n9061 GND.n9060 585
R11883 GND.n9060 GND.n9059 585
R11884 GND.n848 GND.n847 585
R11885 GND.n847 GND.n846 585
R11886 GND.n9066 GND.n9065 585
R11887 GND.n9067 GND.n9066 585
R11888 GND.n845 GND.n844 585
R11889 GND.n9068 GND.n845 585
R11890 GND.n9071 GND.n9070 585
R11891 GND.n9070 GND.n9069 585
R11892 GND.n842 GND.n841 585
R11893 GND.n841 GND.n840 585
R11894 GND.n9076 GND.n9075 585
R11895 GND.n9077 GND.n9076 585
R11896 GND.n839 GND.n838 585
R11897 GND.n9078 GND.n839 585
R11898 GND.n9081 GND.n9080 585
R11899 GND.n9080 GND.n9079 585
R11900 GND.n836 GND.n835 585
R11901 GND.n835 GND.n834 585
R11902 GND.n9086 GND.n9085 585
R11903 GND.n9087 GND.n9086 585
R11904 GND.n833 GND.n832 585
R11905 GND.n9088 GND.n833 585
R11906 GND.n9091 GND.n9090 585
R11907 GND.n9090 GND.n9089 585
R11908 GND.n830 GND.n829 585
R11909 GND.n829 GND.n828 585
R11910 GND.n9096 GND.n9095 585
R11911 GND.n9097 GND.n9096 585
R11912 GND.n827 GND.n826 585
R11913 GND.n9098 GND.n827 585
R11914 GND.n9101 GND.n9100 585
R11915 GND.n9100 GND.n9099 585
R11916 GND.n824 GND.n823 585
R11917 GND.n823 GND.n822 585
R11918 GND.n9106 GND.n9105 585
R11919 GND.n9107 GND.n9106 585
R11920 GND.n821 GND.n820 585
R11921 GND.n9108 GND.n821 585
R11922 GND.n9111 GND.n9110 585
R11923 GND.n9110 GND.n9109 585
R11924 GND.n818 GND.n817 585
R11925 GND.n817 GND.n816 585
R11926 GND.n9116 GND.n9115 585
R11927 GND.n9117 GND.n9116 585
R11928 GND.n815 GND.n814 585
R11929 GND.n9118 GND.n815 585
R11930 GND.n9121 GND.n9120 585
R11931 GND.n9120 GND.n9119 585
R11932 GND.n812 GND.n811 585
R11933 GND.n811 GND.n810 585
R11934 GND.n9126 GND.n9125 585
R11935 GND.n9127 GND.n9126 585
R11936 GND.n809 GND.n808 585
R11937 GND.n9128 GND.n809 585
R11938 GND.n9131 GND.n9130 585
R11939 GND.n9130 GND.n9129 585
R11940 GND.n806 GND.n805 585
R11941 GND.n805 GND.n804 585
R11942 GND.n9136 GND.n9135 585
R11943 GND.n9137 GND.n9136 585
R11944 GND.n803 GND.n802 585
R11945 GND.n9138 GND.n803 585
R11946 GND.n9141 GND.n9140 585
R11947 GND.n9140 GND.n9139 585
R11948 GND.n800 GND.n799 585
R11949 GND.n799 GND.n798 585
R11950 GND.n9146 GND.n9145 585
R11951 GND.n9147 GND.n9146 585
R11952 GND.n797 GND.n796 585
R11953 GND.n9148 GND.n797 585
R11954 GND.n9151 GND.n9150 585
R11955 GND.n9150 GND.n9149 585
R11956 GND.n794 GND.n793 585
R11957 GND.n793 GND.n792 585
R11958 GND.n9156 GND.n9155 585
R11959 GND.n9157 GND.n9156 585
R11960 GND.n791 GND.n790 585
R11961 GND.n9158 GND.n791 585
R11962 GND.n9161 GND.n9160 585
R11963 GND.n9160 GND.n9159 585
R11964 GND.n788 GND.n787 585
R11965 GND.n787 GND.n786 585
R11966 GND.n9166 GND.n9165 585
R11967 GND.n9167 GND.n9166 585
R11968 GND.n785 GND.n784 585
R11969 GND.n9168 GND.n785 585
R11970 GND.n9171 GND.n9170 585
R11971 GND.n9170 GND.n9169 585
R11972 GND.n782 GND.n781 585
R11973 GND.n781 GND.n780 585
R11974 GND.n9176 GND.n9175 585
R11975 GND.n9177 GND.n9176 585
R11976 GND.n779 GND.n778 585
R11977 GND.n9178 GND.n779 585
R11978 GND.n9181 GND.n9180 585
R11979 GND.n9180 GND.n9179 585
R11980 GND.n776 GND.n775 585
R11981 GND.n775 GND.n774 585
R11982 GND.n9186 GND.n9185 585
R11983 GND.n9187 GND.n9186 585
R11984 GND.n773 GND.n772 585
R11985 GND.n9188 GND.n773 585
R11986 GND.n9191 GND.n9190 585
R11987 GND.n9190 GND.n9189 585
R11988 GND.n770 GND.n769 585
R11989 GND.n769 GND.n768 585
R11990 GND.n9196 GND.n9195 585
R11991 GND.n9197 GND.n9196 585
R11992 GND.n767 GND.n766 585
R11993 GND.n9198 GND.n767 585
R11994 GND.n9201 GND.n9200 585
R11995 GND.n9200 GND.n9199 585
R11996 GND.n764 GND.n763 585
R11997 GND.n763 GND.n762 585
R11998 GND.n9206 GND.n9205 585
R11999 GND.n9207 GND.n9206 585
R12000 GND.n761 GND.n760 585
R12001 GND.n9208 GND.n761 585
R12002 GND.n9211 GND.n9210 585
R12003 GND.n9210 GND.n9209 585
R12004 GND.n758 GND.n757 585
R12005 GND.n757 GND.n756 585
R12006 GND.n9216 GND.n9215 585
R12007 GND.n9217 GND.n9216 585
R12008 GND.n755 GND.n754 585
R12009 GND.n9218 GND.n755 585
R12010 GND.n9221 GND.n9220 585
R12011 GND.n9220 GND.n9219 585
R12012 GND.n752 GND.n751 585
R12013 GND.n751 GND.n750 585
R12014 GND.n9226 GND.n9225 585
R12015 GND.n9227 GND.n9226 585
R12016 GND.n749 GND.n748 585
R12017 GND.n9228 GND.n749 585
R12018 GND.n9231 GND.n9230 585
R12019 GND.n9230 GND.n9229 585
R12020 GND.n746 GND.n745 585
R12021 GND.n745 GND.n744 585
R12022 GND.n9236 GND.n9235 585
R12023 GND.n9237 GND.n9236 585
R12024 GND.n743 GND.n742 585
R12025 GND.n9238 GND.n743 585
R12026 GND.n9241 GND.n9240 585
R12027 GND.n9240 GND.n9239 585
R12028 GND.n740 GND.n739 585
R12029 GND.n739 GND.n738 585
R12030 GND.n9246 GND.n9245 585
R12031 GND.n9247 GND.n9246 585
R12032 GND.n737 GND.n736 585
R12033 GND.n9248 GND.n737 585
R12034 GND.n9251 GND.n9250 585
R12035 GND.n9250 GND.n9249 585
R12036 GND.n734 GND.n733 585
R12037 GND.n733 GND.n732 585
R12038 GND.n9256 GND.n9255 585
R12039 GND.n9257 GND.n9256 585
R12040 GND.n731 GND.n730 585
R12041 GND.n9258 GND.n731 585
R12042 GND.n9261 GND.n9260 585
R12043 GND.n9260 GND.n9259 585
R12044 GND.n728 GND.n727 585
R12045 GND.n727 GND.n726 585
R12046 GND.n9266 GND.n9265 585
R12047 GND.n9267 GND.n9266 585
R12048 GND.n725 GND.n724 585
R12049 GND.n9268 GND.n725 585
R12050 GND.n9271 GND.n9270 585
R12051 GND.n9270 GND.n9269 585
R12052 GND.n722 GND.n721 585
R12053 GND.n721 GND.n720 585
R12054 GND.n9276 GND.n9275 585
R12055 GND.n9277 GND.n9276 585
R12056 GND.n719 GND.n718 585
R12057 GND.n9278 GND.n719 585
R12058 GND.n9281 GND.n9280 585
R12059 GND.n9280 GND.n9279 585
R12060 GND.n716 GND.n715 585
R12061 GND.n715 GND.n714 585
R12062 GND.n9286 GND.n9285 585
R12063 GND.n9287 GND.n9286 585
R12064 GND.n713 GND.n712 585
R12065 GND.n9288 GND.n713 585
R12066 GND.n9291 GND.n9290 585
R12067 GND.n9290 GND.n9289 585
R12068 GND.n710 GND.n709 585
R12069 GND.n709 GND.n708 585
R12070 GND.n9296 GND.n9295 585
R12071 GND.n9297 GND.n9296 585
R12072 GND.n707 GND.n706 585
R12073 GND.n9298 GND.n707 585
R12074 GND.n9301 GND.n9300 585
R12075 GND.n9300 GND.n9299 585
R12076 GND.n704 GND.n703 585
R12077 GND.n703 GND.n702 585
R12078 GND.n9306 GND.n9305 585
R12079 GND.n9307 GND.n9306 585
R12080 GND.n701 GND.n700 585
R12081 GND.n9308 GND.n701 585
R12082 GND.n9311 GND.n9310 585
R12083 GND.n9310 GND.n9309 585
R12084 GND.n698 GND.n697 585
R12085 GND.n697 GND.n696 585
R12086 GND.n9316 GND.n9315 585
R12087 GND.n9317 GND.n9316 585
R12088 GND.n695 GND.n694 585
R12089 GND.n9318 GND.n695 585
R12090 GND.n9321 GND.n9320 585
R12091 GND.n9320 GND.n9319 585
R12092 GND.n692 GND.n691 585
R12093 GND.n691 GND.n690 585
R12094 GND.n9326 GND.n9325 585
R12095 GND.n9327 GND.n9326 585
R12096 GND.n689 GND.n688 585
R12097 GND.n9328 GND.n689 585
R12098 GND.n9331 GND.n9330 585
R12099 GND.n9330 GND.n9329 585
R12100 GND.n686 GND.n685 585
R12101 GND.n685 GND.n684 585
R12102 GND.n9336 GND.n9335 585
R12103 GND.n9337 GND.n9336 585
R12104 GND.n683 GND.n682 585
R12105 GND.n9338 GND.n683 585
R12106 GND.n9341 GND.n9340 585
R12107 GND.n9340 GND.n9339 585
R12108 GND.n680 GND.n679 585
R12109 GND.n679 GND.n678 585
R12110 GND.n9346 GND.n9345 585
R12111 GND.n9347 GND.n9346 585
R12112 GND.n677 GND.n676 585
R12113 GND.n9348 GND.n677 585
R12114 GND.n9351 GND.n9350 585
R12115 GND.n9350 GND.n9349 585
R12116 GND.n674 GND.n673 585
R12117 GND.n673 GND.n672 585
R12118 GND.n9356 GND.n9355 585
R12119 GND.n9357 GND.n9356 585
R12120 GND.n671 GND.n670 585
R12121 GND.n9358 GND.n671 585
R12122 GND.n9361 GND.n9360 585
R12123 GND.n9360 GND.n9359 585
R12124 GND.n668 GND.n667 585
R12125 GND.n667 GND.n666 585
R12126 GND.n9366 GND.n9365 585
R12127 GND.n9367 GND.n9366 585
R12128 GND.n665 GND.n664 585
R12129 GND.n9368 GND.n665 585
R12130 GND.n9371 GND.n9370 585
R12131 GND.n9370 GND.n9369 585
R12132 GND.n662 GND.n661 585
R12133 GND.n661 GND.n660 585
R12134 GND.n9376 GND.n9375 585
R12135 GND.n9377 GND.n9376 585
R12136 GND.n659 GND.n658 585
R12137 GND.n9378 GND.n659 585
R12138 GND.n9381 GND.n9380 585
R12139 GND.n9380 GND.n9379 585
R12140 GND.n656 GND.n655 585
R12141 GND.n655 GND.n654 585
R12142 GND.n9386 GND.n9385 585
R12143 GND.n9387 GND.n9386 585
R12144 GND.n653 GND.n652 585
R12145 GND.n9388 GND.n653 585
R12146 GND.n9391 GND.n9390 585
R12147 GND.n9390 GND.n9389 585
R12148 GND.n650 GND.n649 585
R12149 GND.n649 GND.n648 585
R12150 GND.n9396 GND.n9395 585
R12151 GND.n9397 GND.n9396 585
R12152 GND.n647 GND.n646 585
R12153 GND.n9398 GND.n647 585
R12154 GND.n9401 GND.n9400 585
R12155 GND.n9400 GND.n9399 585
R12156 GND.n644 GND.n643 585
R12157 GND.n643 GND.n642 585
R12158 GND.n9406 GND.n9405 585
R12159 GND.n9407 GND.n9406 585
R12160 GND.n641 GND.n640 585
R12161 GND.n9408 GND.n641 585
R12162 GND.n9411 GND.n9410 585
R12163 GND.n9410 GND.n9409 585
R12164 GND.n638 GND.n637 585
R12165 GND.n637 GND.n636 585
R12166 GND.n9416 GND.n9415 585
R12167 GND.n9417 GND.n9416 585
R12168 GND.n635 GND.n634 585
R12169 GND.n9418 GND.n635 585
R12170 GND.n9421 GND.n9420 585
R12171 GND.n9420 GND.n9419 585
R12172 GND.n632 GND.n631 585
R12173 GND.n631 GND.n630 585
R12174 GND.n9426 GND.n9425 585
R12175 GND.n9427 GND.n9426 585
R12176 GND.n629 GND.n628 585
R12177 GND.n9428 GND.n629 585
R12178 GND.n9431 GND.n9430 585
R12179 GND.n9430 GND.n9429 585
R12180 GND.n626 GND.n625 585
R12181 GND.n625 GND.n624 585
R12182 GND.n9436 GND.n9435 585
R12183 GND.n9437 GND.n9436 585
R12184 GND.n623 GND.n622 585
R12185 GND.n9438 GND.n623 585
R12186 GND.n9441 GND.n9440 585
R12187 GND.n9440 GND.n9439 585
R12188 GND.n620 GND.n619 585
R12189 GND.n619 GND.n618 585
R12190 GND.n9446 GND.n9445 585
R12191 GND.n9447 GND.n9446 585
R12192 GND.n617 GND.n616 585
R12193 GND.n9448 GND.n617 585
R12194 GND.n9451 GND.n9450 585
R12195 GND.n9450 GND.n9449 585
R12196 GND.n614 GND.n613 585
R12197 GND.n613 GND.n612 585
R12198 GND.n9456 GND.n9455 585
R12199 GND.n9457 GND.n9456 585
R12200 GND.n611 GND.n610 585
R12201 GND.n9458 GND.n611 585
R12202 GND.n9461 GND.n9460 585
R12203 GND.n9460 GND.n9459 585
R12204 GND.n608 GND.n607 585
R12205 GND.n607 GND.n606 585
R12206 GND.n9466 GND.n9465 585
R12207 GND.n9467 GND.n9466 585
R12208 GND.n605 GND.n604 585
R12209 GND.n9468 GND.n605 585
R12210 GND.n9471 GND.n9470 585
R12211 GND.n9470 GND.n9469 585
R12212 GND.n602 GND.n601 585
R12213 GND.n601 GND.n600 585
R12214 GND.n9476 GND.n9475 585
R12215 GND.n9477 GND.n9476 585
R12216 GND.n599 GND.n598 585
R12217 GND.n9478 GND.n599 585
R12218 GND.n9481 GND.n9480 585
R12219 GND.n9480 GND.n9479 585
R12220 GND.n596 GND.n595 585
R12221 GND.n595 GND.n594 585
R12222 GND.n9486 GND.n9485 585
R12223 GND.n9487 GND.n9486 585
R12224 GND.n593 GND.n592 585
R12225 GND.n9488 GND.n593 585
R12226 GND.n9491 GND.n9490 585
R12227 GND.n9490 GND.n9489 585
R12228 GND.n590 GND.n589 585
R12229 GND.n589 GND.n588 585
R12230 GND.n9496 GND.n9495 585
R12231 GND.n9497 GND.n9496 585
R12232 GND.n587 GND.n586 585
R12233 GND.n9498 GND.n587 585
R12234 GND.n9501 GND.n9500 585
R12235 GND.n9500 GND.n9499 585
R12236 GND.n584 GND.n583 585
R12237 GND.n583 GND.n582 585
R12238 GND.n9506 GND.n9505 585
R12239 GND.n9507 GND.n9506 585
R12240 GND.n581 GND.n580 585
R12241 GND.n9508 GND.n581 585
R12242 GND.n9511 GND.n9510 585
R12243 GND.n9510 GND.n9509 585
R12244 GND.n578 GND.n577 585
R12245 GND.n577 GND.n576 585
R12246 GND.n9517 GND.n9516 585
R12247 GND.n9518 GND.n9517 585
R12248 GND.n575 GND.n574 585
R12249 GND.n9519 GND.n575 585
R12250 GND.n9522 GND.n9521 585
R12251 GND.n9521 GND.n9520 585
R12252 GND.n9523 GND.n572 585
R12253 GND.n572 GND.n571 585
R12254 GND.n9695 GND.n474 585
R12255 GND.n9695 GND.n9694 585
R12256 GND.n9689 GND.n473 585
R12257 GND.n9693 GND.n473 585
R12258 GND.n9691 GND.n9690 585
R12259 GND.n9692 GND.n9691 585
R12260 GND.n477 GND.n476 585
R12261 GND.n476 GND.n475 585
R12262 GND.n9682 GND.n9681 585
R12263 GND.n9681 GND.n9680 585
R12264 GND.n480 GND.n479 585
R12265 GND.n9679 GND.n480 585
R12266 GND.n9677 GND.n9676 585
R12267 GND.n9678 GND.n9677 585
R12268 GND.n483 GND.n482 585
R12269 GND.n482 GND.n481 585
R12270 GND.n9672 GND.n9671 585
R12271 GND.n9671 GND.n9670 585
R12272 GND.n486 GND.n485 585
R12273 GND.n9669 GND.n486 585
R12274 GND.n9667 GND.n9666 585
R12275 GND.n9668 GND.n9667 585
R12276 GND.n489 GND.n488 585
R12277 GND.n488 GND.n487 585
R12278 GND.n9662 GND.n9661 585
R12279 GND.n9661 GND.n9660 585
R12280 GND.n492 GND.n491 585
R12281 GND.n9659 GND.n492 585
R12282 GND.n9657 GND.n9656 585
R12283 GND.n9658 GND.n9657 585
R12284 GND.n495 GND.n494 585
R12285 GND.n494 GND.n493 585
R12286 GND.n9652 GND.n9651 585
R12287 GND.n9651 GND.n9650 585
R12288 GND.n498 GND.n497 585
R12289 GND.n9649 GND.n498 585
R12290 GND.n9647 GND.n9646 585
R12291 GND.n9648 GND.n9647 585
R12292 GND.n501 GND.n500 585
R12293 GND.n500 GND.n499 585
R12294 GND.n9642 GND.n9641 585
R12295 GND.n9641 GND.n9640 585
R12296 GND.n504 GND.n503 585
R12297 GND.n9639 GND.n504 585
R12298 GND.n9637 GND.n9636 585
R12299 GND.n9638 GND.n9637 585
R12300 GND.n507 GND.n506 585
R12301 GND.n506 GND.n505 585
R12302 GND.n9632 GND.n9631 585
R12303 GND.n9631 GND.n9630 585
R12304 GND.n510 GND.n509 585
R12305 GND.n9629 GND.n510 585
R12306 GND.n9627 GND.n9626 585
R12307 GND.n9628 GND.n9627 585
R12308 GND.n513 GND.n512 585
R12309 GND.n512 GND.n511 585
R12310 GND.n9622 GND.n9621 585
R12311 GND.n9621 GND.n9620 585
R12312 GND.n516 GND.n515 585
R12313 GND.n9619 GND.n516 585
R12314 GND.n9617 GND.n9616 585
R12315 GND.n9618 GND.n9617 585
R12316 GND.n519 GND.n518 585
R12317 GND.n518 GND.n517 585
R12318 GND.n9612 GND.n9611 585
R12319 GND.n9611 GND.n9610 585
R12320 GND.n522 GND.n521 585
R12321 GND.n9609 GND.n522 585
R12322 GND.n9607 GND.n9606 585
R12323 GND.n9608 GND.n9607 585
R12324 GND.n525 GND.n524 585
R12325 GND.n524 GND.n523 585
R12326 GND.n9602 GND.n9601 585
R12327 GND.n9601 GND.n9600 585
R12328 GND.n528 GND.n527 585
R12329 GND.n9599 GND.n528 585
R12330 GND.n9597 GND.n9596 585
R12331 GND.n9598 GND.n9597 585
R12332 GND.n531 GND.n530 585
R12333 GND.n530 GND.n529 585
R12334 GND.n9592 GND.n9591 585
R12335 GND.n9591 GND.n9590 585
R12336 GND.n534 GND.n533 585
R12337 GND.n9589 GND.n534 585
R12338 GND.n9587 GND.n9586 585
R12339 GND.n9588 GND.n9587 585
R12340 GND.n537 GND.n536 585
R12341 GND.n536 GND.n535 585
R12342 GND.n9582 GND.n9581 585
R12343 GND.n9581 GND.n9580 585
R12344 GND.n540 GND.n539 585
R12345 GND.n9579 GND.n540 585
R12346 GND.n9577 GND.n9576 585
R12347 GND.n9578 GND.n9577 585
R12348 GND.n543 GND.n542 585
R12349 GND.n542 GND.n541 585
R12350 GND.n9572 GND.n9571 585
R12351 GND.n9571 GND.n9570 585
R12352 GND.n546 GND.n545 585
R12353 GND.n9569 GND.n546 585
R12354 GND.n9567 GND.n9566 585
R12355 GND.n9568 GND.n9567 585
R12356 GND.n549 GND.n548 585
R12357 GND.n548 GND.n547 585
R12358 GND.n9562 GND.n9561 585
R12359 GND.n9561 GND.n9560 585
R12360 GND.n552 GND.n551 585
R12361 GND.n9559 GND.n552 585
R12362 GND.n9557 GND.n9556 585
R12363 GND.n9558 GND.n9557 585
R12364 GND.n555 GND.n554 585
R12365 GND.n554 GND.n553 585
R12366 GND.n9552 GND.n9551 585
R12367 GND.n9551 GND.n9550 585
R12368 GND.n558 GND.n557 585
R12369 GND.n9549 GND.n558 585
R12370 GND.n9547 GND.n9546 585
R12371 GND.n9548 GND.n9547 585
R12372 GND.n561 GND.n560 585
R12373 GND.n560 GND.n559 585
R12374 GND.n9542 GND.n9541 585
R12375 GND.n9541 GND.n9540 585
R12376 GND.n564 GND.n563 585
R12377 GND.n9539 GND.n564 585
R12378 GND.n9537 GND.n9536 585
R12379 GND.n9538 GND.n9537 585
R12380 GND.n567 GND.n566 585
R12381 GND.n566 GND.n565 585
R12382 GND.n9532 GND.n9531 585
R12383 GND.n9531 GND.n9530 585
R12384 GND.n570 GND.n569 585
R12385 GND.n9529 GND.n570 585
R12386 GND.n9527 GND.n9526 585
R12387 GND.n9528 GND.n9527 585
R12388 GND.n10134 GND.n10133 585
R12389 GND.n10135 GND.n10134 585
R12390 GND.n405 GND.n404 585
R12391 GND.n408 GND.n405 585
R12392 GND.n10143 GND.n10142 585
R12393 GND.n10142 GND.n10141 585
R12394 GND.n10144 GND.n400 585
R12395 GND.n400 GND.n399 585
R12396 GND.n10146 GND.n10145 585
R12397 GND.n10147 GND.n10146 585
R12398 GND.n386 GND.n385 585
R12399 GND.n389 GND.n386 585
R12400 GND.n10155 GND.n10154 585
R12401 GND.n10154 GND.n10153 585
R12402 GND.n10156 GND.n381 585
R12403 GND.n381 GND.n380 585
R12404 GND.n10158 GND.n10157 585
R12405 GND.n10159 GND.n10158 585
R12406 GND.n367 GND.n366 585
R12407 GND.n370 GND.n367 585
R12408 GND.n10167 GND.n10166 585
R12409 GND.n10166 GND.n10165 585
R12410 GND.n10168 GND.n362 585
R12411 GND.n362 GND.n361 585
R12412 GND.n10170 GND.n10169 585
R12413 GND.n10171 GND.n10170 585
R12414 GND.n346 GND.n345 585
R12415 GND.n358 GND.n346 585
R12416 GND.n10179 GND.n10178 585
R12417 GND.n10178 GND.n10177 585
R12418 GND.n10180 GND.n341 585
R12419 GND.n10104 GND.n341 585
R12420 GND.n10182 GND.n10181 585
R12421 GND.n10183 GND.n10182 585
R12422 GND.n325 GND.n324 585
R12423 GND.n9787 GND.n325 585
R12424 GND.n10191 GND.n10190 585
R12425 GND.n10190 GND.n10189 585
R12426 GND.n10192 GND.n320 585
R12427 GND.n9780 GND.n320 585
R12428 GND.n10194 GND.n10193 585
R12429 GND.n10195 GND.n10194 585
R12430 GND.n304 GND.n303 585
R12431 GND.n9772 GND.n304 585
R12432 GND.n10203 GND.n10202 585
R12433 GND.n10202 GND.n10201 585
R12434 GND.n10204 GND.n299 585
R12435 GND.n9765 GND.n299 585
R12436 GND.n10206 GND.n10205 585
R12437 GND.n10207 GND.n10206 585
R12438 GND.n283 GND.n282 585
R12439 GND.n9757 GND.n283 585
R12440 GND.n10215 GND.n10214 585
R12441 GND.n10214 GND.n10213 585
R12442 GND.n10216 GND.n278 585
R12443 GND.n9750 GND.n278 585
R12444 GND.n10218 GND.n10217 585
R12445 GND.n10219 GND.n10218 585
R12446 GND.n262 GND.n261 585
R12447 GND.n9742 GND.n262 585
R12448 GND.n10227 GND.n10226 585
R12449 GND.n10226 GND.n10225 585
R12450 GND.n10228 GND.n257 585
R12451 GND.n9735 GND.n257 585
R12452 GND.n10230 GND.n10229 585
R12453 GND.n10231 GND.n10230 585
R12454 GND.n242 GND.n241 585
R12455 GND.n9727 GND.n242 585
R12456 GND.n10239 GND.n10238 585
R12457 GND.n10238 GND.n10237 585
R12458 GND.n10240 GND.n237 585
R12459 GND.n6835 GND.n237 585
R12460 GND.n10242 GND.n10241 585
R12461 GND.n10243 GND.n10242 585
R12462 GND.n221 GND.n220 585
R12463 GND.n6841 GND.n221 585
R12464 GND.n10251 GND.n10250 585
R12465 GND.n10250 GND.n10249 585
R12466 GND.n10252 GND.n216 585
R12467 GND.n6847 GND.n216 585
R12468 GND.n10254 GND.n10253 585
R12469 GND.n10255 GND.n10254 585
R12470 GND.n200 GND.n199 585
R12471 GND.n6853 GND.n200 585
R12472 GND.n10263 GND.n10262 585
R12473 GND.n10262 GND.n10261 585
R12474 GND.n10264 GND.n195 585
R12475 GND.n6859 GND.n195 585
R12476 GND.n10266 GND.n10265 585
R12477 GND.n10267 GND.n10266 585
R12478 GND.n179 GND.n178 585
R12479 GND.n6865 GND.n179 585
R12480 GND.n10275 GND.n10274 585
R12481 GND.n10274 GND.n10273 585
R12482 GND.n10276 GND.n174 585
R12483 GND.n6871 GND.n174 585
R12484 GND.n10278 GND.n10277 585
R12485 GND.n10279 GND.n10278 585
R12486 GND.n158 GND.n157 585
R12487 GND.n6877 GND.n158 585
R12488 GND.n10287 GND.n10286 585
R12489 GND.n10286 GND.n10285 585
R12490 GND.n10288 GND.n153 585
R12491 GND.n6883 GND.n153 585
R12492 GND.n10290 GND.n10289 585
R12493 GND.n10291 GND.n10290 585
R12494 GND.n138 GND.n137 585
R12495 GND.n6889 GND.n138 585
R12496 GND.n10299 GND.n10298 585
R12497 GND.n10298 GND.n10297 585
R12498 GND.n10300 GND.n132 585
R12499 GND.n6895 GND.n132 585
R12500 GND.n10302 GND.n10301 585
R12501 GND.n10303 GND.n10302 585
R12502 GND.n133 GND.n131 585
R12503 GND.n6901 GND.n131 585
R12504 GND.n6791 GND.n6790 585
R12505 GND.n6790 GND.n5269 585
R12506 GND.n6789 GND.n5280 585
R12507 GND.n6789 GND.n6788 585
R12508 GND.n6782 GND.n111 585
R12509 GND.n10310 GND.n111 585
R12510 GND.n6781 GND.n6780 585
R12511 GND.n6780 GND.n6779 585
R12512 GND.n5285 GND.n5284 585
R12513 GND.n5285 GND.n5192 585
R12514 GND.n5183 GND.n5182 585
R12515 GND.n6916 GND.n5183 585
R12516 GND.n6922 GND.n6921 585
R12517 GND.n6921 GND.n6920 585
R12518 GND.n6923 GND.n5178 585
R12519 GND.n6769 GND.n5178 585
R12520 GND.n6925 GND.n6924 585
R12521 GND.n6926 GND.n6925 585
R12522 GND.n5164 GND.n5163 585
R12523 GND.n6754 GND.n5164 585
R12524 GND.n6934 GND.n6933 585
R12525 GND.n6933 GND.n6932 585
R12526 GND.n6935 GND.n5159 585
R12527 GND.n6579 GND.n5159 585
R12528 GND.n6937 GND.n6936 585
R12529 GND.n6938 GND.n6937 585
R12530 GND.n5143 GND.n5142 585
R12531 GND.n6585 GND.n5143 585
R12532 GND.n6946 GND.n6945 585
R12533 GND.n6945 GND.n6944 585
R12534 GND.n6947 GND.n5138 585
R12535 GND.n6591 GND.n5138 585
R12536 GND.n6949 GND.n6948 585
R12537 GND.n6950 GND.n6949 585
R12538 GND.n5122 GND.n5121 585
R12539 GND.n6597 GND.n5122 585
R12540 GND.n6958 GND.n6957 585
R12541 GND.n6957 GND.n6956 585
R12542 GND.n6959 GND.n5117 585
R12543 GND.n6603 GND.n5117 585
R12544 GND.n6961 GND.n6960 585
R12545 GND.n6962 GND.n6961 585
R12546 GND.n5101 GND.n5100 585
R12547 GND.n6609 GND.n5101 585
R12548 GND.n6970 GND.n6969 585
R12549 GND.n6969 GND.n6968 585
R12550 GND.n6971 GND.n5096 585
R12551 GND.n6615 GND.n5096 585
R12552 GND.n6973 GND.n6972 585
R12553 GND.n6974 GND.n6973 585
R12554 GND.n5080 GND.n5079 585
R12555 GND.n6621 GND.n5080 585
R12556 GND.n6982 GND.n6981 585
R12557 GND.n6981 GND.n6980 585
R12558 GND.n6983 GND.n5075 585
R12559 GND.n6627 GND.n5075 585
R12560 GND.n6985 GND.n6984 585
R12561 GND.n6986 GND.n6985 585
R12562 GND.n5059 GND.n5058 585
R12563 GND.n6633 GND.n5059 585
R12564 GND.n6994 GND.n6993 585
R12565 GND.n6993 GND.n6992 585
R12566 GND.n6995 GND.n5054 585
R12567 GND.n6639 GND.n5054 585
R12568 GND.n6997 GND.n6996 585
R12569 GND.n6998 GND.n6997 585
R12570 GND.n5038 GND.n5037 585
R12571 GND.n6645 GND.n5038 585
R12572 GND.n7006 GND.n7005 585
R12573 GND.n7005 GND.n7004 585
R12574 GND.n7007 GND.n5033 585
R12575 GND.n6651 GND.n5033 585
R12576 GND.n7009 GND.n7008 585
R12577 GND.n7010 GND.n7009 585
R12578 GND.n5017 GND.n5016 585
R12579 GND.n6657 GND.n5017 585
R12580 GND.n7018 GND.n7017 585
R12581 GND.n7017 GND.n7016 585
R12582 GND.n7019 GND.n5012 585
R12583 GND.n6663 GND.n5012 585
R12584 GND.n7021 GND.n7020 585
R12585 GND.n7022 GND.n7021 585
R12586 GND.n4997 GND.n4996 585
R12587 GND.n6669 GND.n4997 585
R12588 GND.n7030 GND.n7029 585
R12589 GND.n7029 GND.n7028 585
R12590 GND.n7031 GND.n4992 585
R12591 GND.n6675 GND.n4992 585
R12592 GND.n7033 GND.n7032 585
R12593 GND.n7034 GND.n7033 585
R12594 GND.n4976 GND.n4975 585
R12595 GND.n6516 GND.n4976 585
R12596 GND.n7042 GND.n7041 585
R12597 GND.n7041 GND.n7040 585
R12598 GND.n7043 GND.n4971 585
R12599 GND.n6507 GND.n4971 585
R12600 GND.n7045 GND.n7044 585
R12601 GND.n7046 GND.n7045 585
R12602 GND.n4955 GND.n4954 585
R12603 GND.n6501 GND.n4955 585
R12604 GND.n7054 GND.n7053 585
R12605 GND.n7053 GND.n7052 585
R12606 GND.n7055 GND.n4950 585
R12607 GND.n6493 GND.n4950 585
R12608 GND.n7057 GND.n7056 585
R12609 GND.n7058 GND.n7057 585
R12610 GND.n4934 GND.n4933 585
R12611 GND.n6487 GND.n4934 585
R12612 GND.n7066 GND.n7065 585
R12613 GND.n7065 GND.n7064 585
R12614 GND.n7067 GND.n4928 585
R12615 GND.n6479 GND.n4928 585
R12616 GND.n7069 GND.n7068 585
R12617 GND.n7070 GND.n7069 585
R12618 GND.n4929 GND.n4927 585
R12619 GND.n6473 GND.n4927 585
R12620 GND.n5360 GND.n4910 585
R12621 GND.n7076 GND.n4910 585
R12622 GND.n5359 GND.n5358 585
R12623 GND.n5358 GND.n4906 585
R12624 GND.n5357 GND.n5356 585
R12625 GND.n5357 GND.n4896 585
R12626 GND.n4889 GND.n4887 585
R12627 GND.n7084 GND.n4887 585
R12628 GND.n7090 GND.n7089 585
R12629 GND.n7091 GND.n7090 585
R12630 GND.n4888 GND.n4886 585
R12631 GND.n6416 GND.n4886 585
R12632 GND.n6364 GND.n6363 585
R12633 GND.n6366 GND.n6365 585
R12634 GND.n6369 GND.n6368 585
R12635 GND.n6371 GND.n6370 585
R12636 GND.n6374 GND.n6373 585
R12637 GND.n6376 GND.n6375 585
R12638 GND.n6379 GND.n6378 585
R12639 GND.n6381 GND.n6380 585
R12640 GND.n6384 GND.n6383 585
R12641 GND.n6385 GND.n6358 585
R12642 GND.n10077 GND.n10076 585
R12643 GND.n9811 GND.n9810 585
R12644 GND.n10072 GND.n10071 585
R12645 GND.n10045 GND.n10044 585
R12646 GND.n10067 GND.n10066 585
R12647 GND.n10065 GND.n10064 585
R12648 GND.n10063 GND.n10062 585
R12649 GND.n10056 GND.n10047 585
R12650 GND.n10058 GND.n10057 585
R12651 GND.n10055 GND.n10054 585
R12652 GND.n10053 GND.n10052 585
R12653 GND.n10049 GND.n418 585
R12654 GND.n10080 GND.n416 585
R12655 GND.n10135 GND.n416 585
R12656 GND.n10082 GND.n10081 585
R12657 GND.n10081 GND.n408 585
R12658 GND.n10083 GND.n407 585
R12659 GND.n10141 GND.n407 585
R12660 GND.n10085 GND.n10084 585
R12661 GND.n10084 GND.n399 585
R12662 GND.n10086 GND.n398 585
R12663 GND.n10147 GND.n398 585
R12664 GND.n10088 GND.n10087 585
R12665 GND.n10087 GND.n389 585
R12666 GND.n10089 GND.n388 585
R12667 GND.n10153 GND.n388 585
R12668 GND.n10091 GND.n10090 585
R12669 GND.n10090 GND.n380 585
R12670 GND.n10092 GND.n379 585
R12671 GND.n10159 GND.n379 585
R12672 GND.n10094 GND.n10093 585
R12673 GND.n10093 GND.n370 585
R12674 GND.n10095 GND.n369 585
R12675 GND.n10165 GND.n369 585
R12676 GND.n10097 GND.n10096 585
R12677 GND.n10096 GND.n361 585
R12678 GND.n10098 GND.n360 585
R12679 GND.n10171 GND.n360 585
R12680 GND.n10100 GND.n10099 585
R12681 GND.n10099 GND.n358 585
R12682 GND.n10101 GND.n349 585
R12683 GND.n10177 GND.n349 585
R12684 GND.n10103 GND.n10102 585
R12685 GND.n10104 GND.n10103 585
R12686 GND.n422 GND.n339 585
R12687 GND.n10183 GND.n339 585
R12688 GND.n9789 GND.n9788 585
R12689 GND.n9788 GND.n9787 585
R12690 GND.n424 GND.n328 585
R12691 GND.n10189 GND.n328 585
R12692 GND.n9779 GND.n9778 585
R12693 GND.n9780 GND.n9779 585
R12694 GND.n426 GND.n318 585
R12695 GND.n10195 GND.n318 585
R12696 GND.n9774 GND.n9773 585
R12697 GND.n9773 GND.n9772 585
R12698 GND.n428 GND.n307 585
R12699 GND.n10201 GND.n307 585
R12700 GND.n9764 GND.n9763 585
R12701 GND.n9765 GND.n9764 585
R12702 GND.n430 GND.n297 585
R12703 GND.n10207 GND.n297 585
R12704 GND.n9759 GND.n9758 585
R12705 GND.n9758 GND.n9757 585
R12706 GND.n432 GND.n286 585
R12707 GND.n10213 GND.n286 585
R12708 GND.n9749 GND.n9748 585
R12709 GND.n9750 GND.n9749 585
R12710 GND.n434 GND.n276 585
R12711 GND.n10219 GND.n276 585
R12712 GND.n9744 GND.n9743 585
R12713 GND.n9743 GND.n9742 585
R12714 GND.n436 GND.n265 585
R12715 GND.n10225 GND.n265 585
R12716 GND.n9734 GND.n9733 585
R12717 GND.n9735 GND.n9734 585
R12718 GND.n438 GND.n255 585
R12719 GND.n10231 GND.n255 585
R12720 GND.n9729 GND.n9728 585
R12721 GND.n9728 GND.n9727 585
R12722 GND.n440 GND.n245 585
R12723 GND.n10237 GND.n245 585
R12724 GND.n6837 GND.n6836 585
R12725 GND.n6836 GND.n6835 585
R12726 GND.n6838 GND.n235 585
R12727 GND.n10243 GND.n235 585
R12728 GND.n6840 GND.n6839 585
R12729 GND.n6841 GND.n6840 585
R12730 GND.n6823 GND.n224 585
R12731 GND.n10249 GND.n224 585
R12732 GND.n6849 GND.n6848 585
R12733 GND.n6848 GND.n6847 585
R12734 GND.n6850 GND.n214 585
R12735 GND.n10255 GND.n214 585
R12736 GND.n6852 GND.n6851 585
R12737 GND.n6853 GND.n6852 585
R12738 GND.n6816 GND.n203 585
R12739 GND.n10261 GND.n203 585
R12740 GND.n6861 GND.n6860 585
R12741 GND.n6860 GND.n6859 585
R12742 GND.n6862 GND.n193 585
R12743 GND.n10267 GND.n193 585
R12744 GND.n6864 GND.n6863 585
R12745 GND.n6865 GND.n6864 585
R12746 GND.n6809 GND.n182 585
R12747 GND.n10273 GND.n182 585
R12748 GND.n6873 GND.n6872 585
R12749 GND.n6872 GND.n6871 585
R12750 GND.n6874 GND.n172 585
R12751 GND.n10279 GND.n172 585
R12752 GND.n6876 GND.n6875 585
R12753 GND.n6877 GND.n6876 585
R12754 GND.n6802 GND.n161 585
R12755 GND.n10285 GND.n161 585
R12756 GND.n6885 GND.n6884 585
R12757 GND.n6884 GND.n6883 585
R12758 GND.n6886 GND.n151 585
R12759 GND.n10291 GND.n151 585
R12760 GND.n6888 GND.n6887 585
R12761 GND.n6889 GND.n6888 585
R12762 GND.n5277 GND.n141 585
R12763 GND.n10297 GND.n141 585
R12764 GND.n6897 GND.n6896 585
R12765 GND.n6896 GND.n6895 585
R12766 GND.n6898 GND.n129 585
R12767 GND.n10303 GND.n129 585
R12768 GND.n6900 GND.n6899 585
R12769 GND.n6901 GND.n6900 585
R12770 GND.n5272 GND.n5271 585
R12771 GND.n5271 GND.n5269 585
R12772 GND.n107 GND.n105 585
R12773 GND.n6788 GND.n107 585
R12774 GND.n10312 GND.n10311 585
R12775 GND.n10311 GND.n10310 585
R12776 GND.n106 GND.n104 585
R12777 GND.n6779 GND.n106 585
R12778 GND.n6764 GND.n6763 585
R12779 GND.n6763 GND.n5192 585
R12780 GND.n6765 GND.n5191 585
R12781 GND.n6916 GND.n5191 585
R12782 GND.n6766 GND.n5186 585
R12783 GND.n6920 GND.n5186 585
R12784 GND.n6768 GND.n6767 585
R12785 GND.n6769 GND.n6768 585
R12786 GND.n5288 GND.n5176 585
R12787 GND.n6926 GND.n5176 585
R12788 GND.n6756 GND.n6755 585
R12789 GND.n6755 GND.n6754 585
R12790 GND.n5290 GND.n5167 585
R12791 GND.n6932 GND.n5167 585
R12792 GND.n6578 GND.n6577 585
R12793 GND.n6579 GND.n6578 585
R12794 GND.n6570 GND.n5157 585
R12795 GND.n6938 GND.n5157 585
R12796 GND.n6587 GND.n6586 585
R12797 GND.n6586 GND.n6585 585
R12798 GND.n6588 GND.n5146 585
R12799 GND.n6944 GND.n5146 585
R12800 GND.n6590 GND.n6589 585
R12801 GND.n6591 GND.n6590 585
R12802 GND.n6563 GND.n5136 585
R12803 GND.n6950 GND.n5136 585
R12804 GND.n6599 GND.n6598 585
R12805 GND.n6598 GND.n6597 585
R12806 GND.n6600 GND.n5125 585
R12807 GND.n6956 GND.n5125 585
R12808 GND.n6602 GND.n6601 585
R12809 GND.n6603 GND.n6602 585
R12810 GND.n6556 GND.n5115 585
R12811 GND.n6962 GND.n5115 585
R12812 GND.n6611 GND.n6610 585
R12813 GND.n6610 GND.n6609 585
R12814 GND.n6612 GND.n5104 585
R12815 GND.n6968 GND.n5104 585
R12816 GND.n6614 GND.n6613 585
R12817 GND.n6615 GND.n6614 585
R12818 GND.n6549 GND.n5094 585
R12819 GND.n6974 GND.n5094 585
R12820 GND.n6623 GND.n6622 585
R12821 GND.n6622 GND.n6621 585
R12822 GND.n6624 GND.n5083 585
R12823 GND.n6980 GND.n5083 585
R12824 GND.n6626 GND.n6625 585
R12825 GND.n6627 GND.n6626 585
R12826 GND.n6542 GND.n5073 585
R12827 GND.n6986 GND.n5073 585
R12828 GND.n6635 GND.n6634 585
R12829 GND.n6634 GND.n6633 585
R12830 GND.n6636 GND.n5062 585
R12831 GND.n6992 GND.n5062 585
R12832 GND.n6638 GND.n6637 585
R12833 GND.n6639 GND.n6638 585
R12834 GND.n6535 GND.n5052 585
R12835 GND.n6998 GND.n5052 585
R12836 GND.n6647 GND.n6646 585
R12837 GND.n6646 GND.n6645 585
R12838 GND.n6648 GND.n5041 585
R12839 GND.n7004 GND.n5041 585
R12840 GND.n6650 GND.n6649 585
R12841 GND.n6651 GND.n6650 585
R12842 GND.n6528 GND.n5031 585
R12843 GND.n7010 GND.n5031 585
R12844 GND.n6659 GND.n6658 585
R12845 GND.n6658 GND.n6657 585
R12846 GND.n6660 GND.n5020 585
R12847 GND.n7016 GND.n5020 585
R12848 GND.n6662 GND.n6661 585
R12849 GND.n6663 GND.n6662 585
R12850 GND.n5335 GND.n5010 585
R12851 GND.n7022 GND.n5010 585
R12852 GND.n6671 GND.n6670 585
R12853 GND.n6670 GND.n6669 585
R12854 GND.n6672 GND.n4999 585
R12855 GND.n7028 GND.n4999 585
R12856 GND.n6674 GND.n6673 585
R12857 GND.n6675 GND.n6674 585
R12858 GND.n5331 GND.n4990 585
R12859 GND.n7034 GND.n4990 585
R12860 GND.n6515 GND.n6514 585
R12861 GND.n6516 GND.n6515 585
R12862 GND.n5338 GND.n4979 585
R12863 GND.n7040 GND.n4979 585
R12864 GND.n6509 GND.n6508 585
R12865 GND.n6508 GND.n6507 585
R12866 GND.n5340 GND.n4969 585
R12867 GND.n7046 GND.n4969 585
R12868 GND.n6500 GND.n6499 585
R12869 GND.n6501 GND.n6500 585
R12870 GND.n5343 GND.n4958 585
R12871 GND.n7052 GND.n4958 585
R12872 GND.n6495 GND.n6494 585
R12873 GND.n6494 GND.n6493 585
R12874 GND.n5345 GND.n4948 585
R12875 GND.n7058 GND.n4948 585
R12876 GND.n6486 GND.n6485 585
R12877 GND.n6487 GND.n6486 585
R12878 GND.n5348 GND.n4937 585
R12879 GND.n7064 GND.n4937 585
R12880 GND.n6481 GND.n6480 585
R12881 GND.n6480 GND.n6479 585
R12882 GND.n5350 GND.n4925 585
R12883 GND.n7070 GND.n4925 585
R12884 GND.n6431 GND.n6430 585
R12885 GND.n6473 GND.n6431 585
R12886 GND.n5363 GND.n4908 585
R12887 GND.n7076 GND.n4908 585
R12888 GND.n6426 GND.n6425 585
R12889 GND.n6425 GND.n4906 585
R12890 GND.n6424 GND.n6423 585
R12891 GND.n6424 GND.n4896 585
R12892 GND.n6422 GND.n4895 585
R12893 GND.n7084 GND.n4895 585
R12894 GND.n5365 GND.n4884 585
R12895 GND.n7091 GND.n4884 585
R12896 GND.n6418 GND.n6417 585
R12897 GND.n6417 GND.n6416 585
R12898 GND.n6313 GND.n5496 585
R12899 GND.n6313 GND.n6312 585
R12900 GND.n6193 GND.n4414 585
R12901 GND.n7417 GND.n4414 585
R12902 GND.n6196 GND.n6195 585
R12903 GND.n6195 GND.n6194 585
R12904 GND.n6197 GND.n4405 585
R12905 GND.n7423 GND.n4405 585
R12906 GND.n6199 GND.n6198 585
R12907 GND.n6198 GND.t152 585
R12908 GND.n6200 GND.n4382 585
R12909 GND.n7429 GND.n4382 585
R12910 GND.n6202 GND.n6201 585
R12911 GND.n6203 GND.n6202 585
R12912 GND.n5520 GND.n4368 585
R12913 GND.n7435 GND.n4368 585
R12914 GND.n6183 GND.n6182 585
R12915 GND.n6182 GND.n4360 585
R12916 GND.n6181 GND.n6180 585
R12917 GND.n6181 GND.n4359 585
R12918 GND.n6179 GND.n4351 585
R12919 GND.n7448 GND.n4351 585
R12920 GND.n5524 GND.n5523 585
R12921 GND.n5523 GND.n5522 585
R12922 GND.n6175 GND.n4340 585
R12923 GND.n7454 GND.n4340 585
R12924 GND.n6174 GND.n6173 585
R12925 GND.n6173 GND.n6172 585
R12926 GND.n5526 GND.n4330 585
R12927 GND.n7460 GND.n4330 585
R12928 GND.n6094 GND.n6093 585
R12929 GND.n6093 GND.n5532 585
R12930 GND.n6095 GND.n4320 585
R12931 GND.n7466 GND.n4320 585
R12932 GND.n6097 GND.n6096 585
R12933 GND.n6096 GND.n5537 585
R12934 GND.n6098 GND.n4310 585
R12935 GND.n7472 GND.n4310 585
R12936 GND.n6100 GND.n6099 585
R12937 GND.n6099 GND.n5542 585
R12938 GND.n6101 GND.n4300 585
R12939 GND.n7478 GND.n4300 585
R12940 GND.n6103 GND.n6102 585
R12941 GND.n6102 GND.n5547 585
R12942 GND.n6104 GND.n4278 585
R12943 GND.n7484 GND.n4278 585
R12944 GND.n6106 GND.n6105 585
R12945 GND.n6107 GND.n6106 585
R12946 GND.n5552 GND.n4264 585
R12947 GND.n7490 GND.n4264 585
R12948 GND.n6080 GND.n6079 585
R12949 GND.n6079 GND.n4256 585
R12950 GND.n6078 GND.n6077 585
R12951 GND.n6078 GND.n4255 585
R12952 GND.n6076 GND.n4247 585
R12953 GND.n7503 GND.n4247 585
R12954 GND.n5556 GND.n5555 585
R12955 GND.n5555 GND.n5554 585
R12956 GND.n6072 GND.n4236 585
R12957 GND.n7509 GND.n4236 585
R12958 GND.n6071 GND.n6070 585
R12959 GND.n6070 GND.n6069 585
R12960 GND.n5558 GND.n4227 585
R12961 GND.n7515 GND.n4227 585
R12962 GND.n5991 GND.n5990 585
R12963 GND.n5990 GND.n5565 585
R12964 GND.n5992 GND.n4217 585
R12965 GND.n7521 GND.n4217 585
R12966 GND.n5994 GND.n5993 585
R12967 GND.n5993 GND.n5570 585
R12968 GND.n5995 GND.n4207 585
R12969 GND.n7527 GND.n4207 585
R12970 GND.n5997 GND.n5996 585
R12971 GND.n5996 GND.n5575 585
R12972 GND.n5998 GND.n4198 585
R12973 GND.n7533 GND.n4198 585
R12974 GND.n6000 GND.n5999 585
R12975 GND.n5999 GND.n5581 585
R12976 GND.n6001 GND.n4175 585
R12977 GND.n7539 GND.n4175 585
R12978 GND.n6003 GND.n6002 585
R12979 GND.n6004 GND.n6003 585
R12980 GND.n5585 GND.n4161 585
R12981 GND.n7545 GND.n4161 585
R12982 GND.n5977 GND.n5976 585
R12983 GND.n5976 GND.n4153 585
R12984 GND.n5975 GND.n5974 585
R12985 GND.n5975 GND.n4152 585
R12986 GND.n5973 GND.n4144 585
R12987 GND.n7558 GND.n4144 585
R12988 GND.n5589 GND.n5588 585
R12989 GND.n5588 GND.n5587 585
R12990 GND.n5969 GND.n4133 585
R12991 GND.n7564 GND.n4133 585
R12992 GND.n5968 GND.n5967 585
R12993 GND.n5967 GND.n5966 585
R12994 GND.n5591 GND.n4123 585
R12995 GND.n7570 GND.n4123 585
R12996 GND.n5888 GND.n5887 585
R12997 GND.n5887 GND.n5597 585
R12998 GND.n5889 GND.n4113 585
R12999 GND.n7576 GND.n4113 585
R13000 GND.n5891 GND.n5890 585
R13001 GND.n5890 GND.n5602 585
R13002 GND.n5892 GND.n4103 585
R13003 GND.n7582 GND.n4103 585
R13004 GND.n5894 GND.n5893 585
R13005 GND.n5893 GND.n5607 585
R13006 GND.n5895 GND.n4093 585
R13007 GND.n7588 GND.n4093 585
R13008 GND.n5897 GND.n5896 585
R13009 GND.n5896 GND.n5612 585
R13010 GND.n5898 GND.n4070 585
R13011 GND.n7594 GND.n4070 585
R13012 GND.n5900 GND.n5899 585
R13013 GND.n5901 GND.n5900 585
R13014 GND.n5616 GND.n4056 585
R13015 GND.n7600 GND.n4056 585
R13016 GND.n5874 GND.n5873 585
R13017 GND.n5873 GND.n4048 585
R13018 GND.n5872 GND.n5871 585
R13019 GND.n5872 GND.n4047 585
R13020 GND.n5870 GND.n4039 585
R13021 GND.n7613 GND.n4039 585
R13022 GND.n5620 GND.n5619 585
R13023 GND.n5619 GND.n5618 585
R13024 GND.n5866 GND.n4028 585
R13025 GND.n7619 GND.n4028 585
R13026 GND.n5865 GND.n5864 585
R13027 GND.n5864 GND.n5863 585
R13028 GND.n5622 GND.n4018 585
R13029 GND.n7625 GND.n4018 585
R13030 GND.n5784 GND.n5783 585
R13031 GND.n5783 GND.n5628 585
R13032 GND.n5785 GND.n4008 585
R13033 GND.n7631 GND.n4008 585
R13034 GND.n5787 GND.n5786 585
R13035 GND.n5786 GND.n5633 585
R13036 GND.n5788 GND.n3998 585
R13037 GND.n7637 GND.n3998 585
R13038 GND.n5790 GND.n5789 585
R13039 GND.n5789 GND.n5638 585
R13040 GND.n5791 GND.n3988 585
R13041 GND.n7643 GND.n3988 585
R13042 GND.n5793 GND.n5792 585
R13043 GND.n5792 GND.n5643 585
R13044 GND.n5794 GND.n3965 585
R13045 GND.n7649 GND.n3965 585
R13046 GND.n5796 GND.n5795 585
R13047 GND.n5797 GND.n5796 585
R13048 GND.n5647 GND.n3952 585
R13049 GND.n7655 GND.n3952 585
R13050 GND.n5770 GND.n5769 585
R13051 GND.n5769 GND.n3944 585
R13052 GND.n5768 GND.n5767 585
R13053 GND.n5768 GND.n3943 585
R13054 GND.n5766 GND.n3935 585
R13055 GND.n7668 GND.n3935 585
R13056 GND.n5651 GND.n5650 585
R13057 GND.n5650 GND.n5649 585
R13058 GND.n5762 GND.n3924 585
R13059 GND.n7674 GND.n3924 585
R13060 GND.n5761 GND.n5760 585
R13061 GND.n5760 GND.n5759 585
R13062 GND.n5653 GND.n3914 585
R13063 GND.n7680 GND.n3914 585
R13064 GND.n5676 GND.n5675 585
R13065 GND.n5675 GND.n5659 585
R13066 GND.n5677 GND.n3904 585
R13067 GND.t41 GND.n3904 585
R13068 GND.n5679 GND.n5678 585
R13069 GND.n5678 GND.n5664 585
R13070 GND.n5670 GND.n3895 585
R13071 GND.n7691 GND.n3895 585
R13072 GND.n5684 GND.n5683 585
R13073 GND.n5685 GND.n5684 585
R13074 GND.n5669 GND.n2344 585
R13075 GND.n7697 GND.n2344 585
R13076 GND.n7757 GND.n7756 585
R13077 GND.n7755 GND.n2343 585
R13078 GND.n7754 GND.n2342 585
R13079 GND.n7759 GND.n2342 585
R13080 GND.n7753 GND.n7752 585
R13081 GND.n7751 GND.n7750 585
R13082 GND.n7749 GND.n7748 585
R13083 GND.n7747 GND.n7746 585
R13084 GND.n7745 GND.n7744 585
R13085 GND.n7743 GND.n7742 585
R13086 GND.n7741 GND.n7740 585
R13087 GND.n7739 GND.n2355 585
R13088 GND.n2357 GND.n2356 585
R13089 GND.n7736 GND.n7733 585
R13090 GND.n7735 GND.n7734 585
R13091 GND.n7731 GND.n7728 585
R13092 GND.n7730 GND.n7729 585
R13093 GND.n7726 GND.n7723 585
R13094 GND.n7725 GND.n7724 585
R13095 GND.n7721 GND.n7718 585
R13096 GND.n7720 GND.n7719 585
R13097 GND.n7716 GND.n7713 585
R13098 GND.n7715 GND.n7714 585
R13099 GND.n7711 GND.n3875 585
R13100 GND.n7710 GND.n7709 585
R13101 GND.n7707 GND.n7706 585
R13102 GND.n7705 GND.n7704 585
R13103 GND.n7703 GND.n3880 585
R13104 GND.n3881 GND.n2340 585
R13105 GND.n7759 GND.n2340 585
R13106 GND.n7411 GND.n7410 585
R13107 GND.n4421 GND.n4420 585
R13108 GND.n6348 GND.n6347 585
R13109 GND.n6350 GND.n6349 585
R13110 GND.n6352 GND.n6351 585
R13111 GND.n6355 GND.n6354 585
R13112 GND.n6353 GND.n6341 585
R13113 GND.n5468 GND.n5467 585
R13114 GND.n5470 GND.n5469 585
R13115 GND.n5473 GND.n5472 585
R13116 GND.n5475 GND.n5474 585
R13117 GND.n5478 GND.n5477 585
R13118 GND.n5480 GND.n5479 585
R13119 GND.n5483 GND.n5482 585
R13120 GND.n5485 GND.n5484 585
R13121 GND.n5488 GND.n5487 585
R13122 GND.n5490 GND.n5489 585
R13123 GND.n6339 GND.n6338 585
R13124 GND.n6337 GND.n6336 585
R13125 GND.n6335 GND.n6334 585
R13126 GND.n6333 GND.n5491 585
R13127 GND.n6329 GND.n6328 585
R13128 GND.n6327 GND.n6326 585
R13129 GND.n6325 GND.n6324 585
R13130 GND.n6323 GND.n5493 585
R13131 GND.n6319 GND.n6318 585
R13132 GND.n6317 GND.n6316 585
R13133 GND.n6315 GND.n6314 585
R13134 GND.n7414 GND.n4416 585
R13135 GND.n6312 GND.n4416 585
R13136 GND.n7416 GND.n7415 585
R13137 GND.n7417 GND.n7416 585
R13138 GND.n4403 GND.n4402 585
R13139 GND.n6194 GND.n4403 585
R13140 GND.n7425 GND.n7424 585
R13141 GND.n7424 GND.n7423 585
R13142 GND.n7426 GND.n4385 585
R13143 GND.t152 GND.n4385 585
R13144 GND.n7428 GND.n7427 585
R13145 GND.n7429 GND.n7428 585
R13146 GND.n4386 GND.n4384 585
R13147 GND.n6203 GND.n4384 585
R13148 GND.n4396 GND.n4370 585
R13149 GND.n7435 GND.n4370 585
R13150 GND.n4395 GND.n4394 585
R13151 GND.n4394 GND.n4360 585
R13152 GND.n4393 GND.n4392 585
R13153 GND.n4393 GND.n4359 585
R13154 GND.n4388 GND.n4353 585
R13155 GND.n7448 GND.n4353 585
R13156 GND.n4338 GND.n4337 585
R13157 GND.n5522 GND.n4338 585
R13158 GND.n7456 GND.n7455 585
R13159 GND.n7455 GND.n7454 585
R13160 GND.n7457 GND.n4332 585
R13161 GND.n6172 GND.n4332 585
R13162 GND.n7459 GND.n7458 585
R13163 GND.n7460 GND.n7459 585
R13164 GND.n4318 GND.n4317 585
R13165 GND.n5532 GND.n4318 585
R13166 GND.n7468 GND.n7467 585
R13167 GND.n7467 GND.n7466 585
R13168 GND.n7469 GND.n4312 585
R13169 GND.n5537 GND.n4312 585
R13170 GND.n7471 GND.n7470 585
R13171 GND.n7472 GND.n7471 585
R13172 GND.n4298 GND.n4297 585
R13173 GND.n5542 GND.n4298 585
R13174 GND.n7480 GND.n7479 585
R13175 GND.n7479 GND.n7478 585
R13176 GND.n7481 GND.n4280 585
R13177 GND.n5547 GND.n4280 585
R13178 GND.n7483 GND.n7482 585
R13179 GND.n7484 GND.n7483 585
R13180 GND.n4281 GND.n4279 585
R13181 GND.n6107 GND.n4279 585
R13182 GND.n4291 GND.n4266 585
R13183 GND.n7490 GND.n4266 585
R13184 GND.n4290 GND.n4289 585
R13185 GND.n4289 GND.n4256 585
R13186 GND.n4288 GND.n4287 585
R13187 GND.n4288 GND.n4255 585
R13188 GND.n4283 GND.n4249 585
R13189 GND.n7503 GND.n4249 585
R13190 GND.n4234 GND.n4233 585
R13191 GND.n5554 GND.n4234 585
R13192 GND.n7511 GND.n7510 585
R13193 GND.n7510 GND.n7509 585
R13194 GND.n7512 GND.n4228 585
R13195 GND.n6069 GND.n4228 585
R13196 GND.n7514 GND.n7513 585
R13197 GND.n7515 GND.n7514 585
R13198 GND.n4215 GND.n4214 585
R13199 GND.n5565 GND.n4215 585
R13200 GND.n7523 GND.n7522 585
R13201 GND.n7522 GND.n7521 585
R13202 GND.n7524 GND.n4209 585
R13203 GND.n5570 GND.n4209 585
R13204 GND.n7526 GND.n7525 585
R13205 GND.n7527 GND.n7526 585
R13206 GND.n4196 GND.n4195 585
R13207 GND.n5575 GND.n4196 585
R13208 GND.n7535 GND.n7534 585
R13209 GND.n7534 GND.n7533 585
R13210 GND.n7536 GND.n4178 585
R13211 GND.n5581 GND.n4178 585
R13212 GND.n7538 GND.n7537 585
R13213 GND.n7539 GND.n7538 585
R13214 GND.n4179 GND.n4177 585
R13215 GND.n6004 GND.n4177 585
R13216 GND.n4189 GND.n4163 585
R13217 GND.n7545 GND.n4163 585
R13218 GND.n4188 GND.n4187 585
R13219 GND.n4187 GND.n4153 585
R13220 GND.n4186 GND.n4185 585
R13221 GND.n4186 GND.n4152 585
R13222 GND.n4181 GND.n4146 585
R13223 GND.n7558 GND.n4146 585
R13224 GND.n4131 GND.n4130 585
R13225 GND.n5587 GND.n4131 585
R13226 GND.n7566 GND.n7565 585
R13227 GND.n7565 GND.n7564 585
R13228 GND.n7567 GND.n4125 585
R13229 GND.n5966 GND.n4125 585
R13230 GND.n7569 GND.n7568 585
R13231 GND.n7570 GND.n7569 585
R13232 GND.n4111 GND.n4110 585
R13233 GND.n5597 GND.n4111 585
R13234 GND.n7578 GND.n7577 585
R13235 GND.n7577 GND.n7576 585
R13236 GND.n7579 GND.n4105 585
R13237 GND.n5602 GND.n4105 585
R13238 GND.n7581 GND.n7580 585
R13239 GND.n7582 GND.n7581 585
R13240 GND.n4091 GND.n4090 585
R13241 GND.n5607 GND.n4091 585
R13242 GND.n7590 GND.n7589 585
R13243 GND.n7589 GND.n7588 585
R13244 GND.n7591 GND.n4073 585
R13245 GND.n5612 GND.n4073 585
R13246 GND.n7593 GND.n7592 585
R13247 GND.n7594 GND.n7593 585
R13248 GND.n4074 GND.n4072 585
R13249 GND.n5901 GND.n4072 585
R13250 GND.n4084 GND.n4058 585
R13251 GND.n7600 GND.n4058 585
R13252 GND.n4083 GND.n4082 585
R13253 GND.n4082 GND.n4048 585
R13254 GND.n4081 GND.n4080 585
R13255 GND.n4081 GND.n4047 585
R13256 GND.n4076 GND.n4041 585
R13257 GND.n7613 GND.n4041 585
R13258 GND.n4026 GND.n4025 585
R13259 GND.n5618 GND.n4026 585
R13260 GND.n7621 GND.n7620 585
R13261 GND.n7620 GND.n7619 585
R13262 GND.n7622 GND.n4020 585
R13263 GND.n5863 GND.n4020 585
R13264 GND.n7624 GND.n7623 585
R13265 GND.n7625 GND.n7624 585
R13266 GND.n4006 GND.n4005 585
R13267 GND.n5628 GND.n4006 585
R13268 GND.n7633 GND.n7632 585
R13269 GND.n7632 GND.n7631 585
R13270 GND.n7634 GND.n4000 585
R13271 GND.n5633 GND.n4000 585
R13272 GND.n7636 GND.n7635 585
R13273 GND.n7637 GND.n7636 585
R13274 GND.n3986 GND.n3985 585
R13275 GND.n5638 GND.n3986 585
R13276 GND.n7645 GND.n7644 585
R13277 GND.n7644 GND.n7643 585
R13278 GND.n7646 GND.n3968 585
R13279 GND.n5643 GND.n3968 585
R13280 GND.n7648 GND.n7647 585
R13281 GND.n7649 GND.n7648 585
R13282 GND.n3969 GND.n3967 585
R13283 GND.n5797 GND.n3967 585
R13284 GND.n3979 GND.n3953 585
R13285 GND.n7655 GND.n3953 585
R13286 GND.n3978 GND.n3977 585
R13287 GND.n3977 GND.n3944 585
R13288 GND.n3976 GND.n3975 585
R13289 GND.n3976 GND.n3943 585
R13290 GND.n3971 GND.n3937 585
R13291 GND.n7668 GND.n3937 585
R13292 GND.n3922 GND.n3921 585
R13293 GND.n5649 GND.n3922 585
R13294 GND.n7676 GND.n7675 585
R13295 GND.n7675 GND.n7674 585
R13296 GND.n7677 GND.n3916 585
R13297 GND.n5759 GND.n3916 585
R13298 GND.n7679 GND.n7678 585
R13299 GND.n7680 GND.n7679 585
R13300 GND.n3902 GND.n3901 585
R13301 GND.n5659 GND.n3902 585
R13302 GND.n7687 GND.n7686 585
R13303 GND.n7686 GND.t41 585
R13304 GND.n7688 GND.n3897 585
R13305 GND.n5664 GND.n3897 585
R13306 GND.n7690 GND.n7689 585
R13307 GND.n7691 GND.n7690 585
R13308 GND.n3884 GND.n3883 585
R13309 GND.n5685 GND.n3884 585
R13310 GND.n7699 GND.n7698 585
R13311 GND.n7698 GND.n7697 585
R13312 GND.n4769 GND.n4731 585
R13313 GND.n4731 GND.n4700 585
R13314 GND.n4771 GND.n4770 585
R13315 GND.n4772 GND.n4771 585
R13316 GND.n4686 GND.n4685 585
R13317 GND.n4689 GND.n4686 585
R13318 GND.n7260 GND.n7259 585
R13319 GND.n7259 GND.n7258 585
R13320 GND.n7261 GND.n4678 585
R13321 GND.n4687 GND.n4678 585
R13322 GND.n7263 GND.n7262 585
R13323 GND.n7264 GND.n7263 585
R13324 GND.n4684 GND.n4677 585
R13325 GND.n4677 GND.n4623 585
R13326 GND.n4683 GND.n4622 585
R13327 GND.n7270 GND.n4622 585
R13328 GND.n4682 GND.n4681 585
R13329 GND.n4681 GND.n4680 585
R13330 GND.n4612 GND.n4611 585
R13331 GND.n4614 GND.n4612 585
R13332 GND.n7279 GND.n7278 585
R13333 GND.n7278 GND.n7277 585
R13334 GND.n7280 GND.n4609 585
R13335 GND.n4666 GND.n4609 585
R13336 GND.n7282 GND.n7281 585
R13337 GND.n7283 GND.n7282 585
R13338 GND.n4610 GND.n4608 585
R13339 GND.n4608 GND.n4605 585
R13340 GND.n4660 GND.n4659 585
R13341 GND.n4661 GND.n4660 585
R13342 GND.n4594 GND.n4593 585
R13343 GND.n4597 GND.n4594 585
R13344 GND.n7293 GND.n7292 585
R13345 GND.n7292 GND.n7291 585
R13346 GND.n7294 GND.n4591 585
R13347 GND.n4595 GND.n4591 585
R13348 GND.n7296 GND.n7295 585
R13349 GND.n7297 GND.n7296 585
R13350 GND.n4592 GND.n4590 585
R13351 GND.n4590 GND.n4587 585
R13352 GND.n4647 GND.n4646 585
R13353 GND.n4648 GND.n4647 585
R13354 GND.n4576 GND.n4575 585
R13355 GND.n4579 GND.n4576 585
R13356 GND.n7307 GND.n7306 585
R13357 GND.n7306 GND.n7305 585
R13358 GND.n7308 GND.n4573 585
R13359 GND.n4577 GND.n4573 585
R13360 GND.n7310 GND.n7309 585
R13361 GND.n7311 GND.n7310 585
R13362 GND.n4574 GND.n4572 585
R13363 GND.n4572 GND.n4569 585
R13364 GND.n4634 GND.n4633 585
R13365 GND.n4635 GND.n4634 585
R13366 GND.n4555 GND.n4554 585
R13367 GND.n4558 GND.n4555 585
R13368 GND.n7321 GND.n7320 585
R13369 GND.n7320 GND.n7319 585
R13370 GND.n7322 GND.n4549 585
R13371 GND.n4556 GND.n4549 585
R13372 GND.n7324 GND.n7323 585
R13373 GND.n7325 GND.n7324 585
R13374 GND.n4553 GND.n4548 585
R13375 GND.n4548 GND.n4540 585
R13376 GND.n4552 GND.n4539 585
R13377 GND.n7331 GND.n4539 585
R13378 GND.n4551 GND.n4550 585
R13379 GND.n4550 GND.n4538 585
R13380 GND.n4526 GND.n4525 585
R13381 GND.n4529 GND.n4526 585
R13382 GND.n7340 GND.n7339 585
R13383 GND.n7339 GND.n7338 585
R13384 GND.n7341 GND.n4523 585
R13385 GND.n4527 GND.n4523 585
R13386 GND.n7343 GND.n7342 585
R13387 GND.n7344 GND.n7343 585
R13388 GND.n4524 GND.n4522 585
R13389 GND.n4522 GND.n4519 585
R13390 GND.n6252 GND.n6251 585
R13391 GND.n6253 GND.n6252 585
R13392 GND.n4508 GND.n4507 585
R13393 GND.n4511 GND.n4508 585
R13394 GND.n7354 GND.n7353 585
R13395 GND.n7353 GND.n7352 585
R13396 GND.n7355 GND.n4505 585
R13397 GND.n4509 GND.n4505 585
R13398 GND.n7357 GND.n7356 585
R13399 GND.n7358 GND.n7357 585
R13400 GND.n4506 GND.n4504 585
R13401 GND.n4504 GND.n4501 585
R13402 GND.n6265 GND.n6264 585
R13403 GND.n6266 GND.n6265 585
R13404 GND.n4490 GND.n4489 585
R13405 GND.n4493 GND.n4490 585
R13406 GND.n7368 GND.n7367 585
R13407 GND.n7367 GND.n7366 585
R13408 GND.n7369 GND.n4487 585
R13409 GND.n4491 GND.n4487 585
R13410 GND.n7371 GND.n7370 585
R13411 GND.n7372 GND.n7371 585
R13412 GND.n4488 GND.n4486 585
R13413 GND.n4486 GND.n4483 585
R13414 GND.n6278 GND.n6277 585
R13415 GND.n6279 GND.n6278 585
R13416 GND.n4472 GND.n4471 585
R13417 GND.n4475 GND.n4472 585
R13418 GND.n7382 GND.n7381 585
R13419 GND.n7381 GND.n7380 585
R13420 GND.n7383 GND.n4469 585
R13421 GND.n4473 GND.n4469 585
R13422 GND.n7385 GND.n7384 585
R13423 GND.n7386 GND.n7385 585
R13424 GND.n4470 GND.n4468 585
R13425 GND.n4468 GND.n4465 585
R13426 GND.n6290 GND.n6289 585
R13427 GND.n6291 GND.n6290 585
R13428 GND.n4454 GND.n4453 585
R13429 GND.n4457 GND.n4454 585
R13430 GND.n7396 GND.n7395 585
R13431 GND.n7395 GND.n7394 585
R13432 GND.n7397 GND.n4451 585
R13433 GND.n4451 GND.n4449 585
R13434 GND.n7399 GND.n7398 585
R13435 GND.n7400 GND.n7399 585
R13436 GND.n4452 GND.n4450 585
R13437 GND.n4450 GND.n4447 585
R13438 GND.n6304 GND.n5504 585
R13439 GND.n6304 GND.n6303 585
R13440 GND.n6305 GND.n5503 585
R13441 GND.n6305 GND.n4436 585
R13442 GND.n6307 GND.n6306 585
R13443 GND.n6306 GND.n4422 585
R13444 GND.n6308 GND.n5501 585
R13445 GND.n5501 GND.n5499 585
R13446 GND.n6310 GND.n6309 585
R13447 GND.n6311 GND.n6310 585
R13448 GND.n5502 GND.n5500 585
R13449 GND.n5500 GND.n4415 585
R13450 GND.n6227 GND.n6226 585
R13451 GND.n6228 GND.n6227 585
R13452 GND.n6225 GND.n5510 585
R13453 GND.n5510 GND.n5509 585
R13454 GND.n6224 GND.n6223 585
R13455 GND.n6223 GND.n4406 585
R13456 GND.n6222 GND.n5511 585
R13457 GND.n6222 GND.n4404 585
R13458 GND.n6221 GND.n5513 585
R13459 GND.n6221 GND.n6220 585
R13460 GND.n6205 GND.n5512 585
R13461 GND.n5512 GND.n4383 585
R13462 GND.n6206 GND.n6204 585
R13463 GND.n6204 GND.n4381 585
R13464 GND.n6208 GND.n6207 585
R13465 GND.n6209 GND.n6208 585
R13466 GND.n4365 GND.n4364 585
R13467 GND.n4369 GND.n4365 585
R13468 GND.n7438 GND.n7437 585
R13469 GND.n7437 GND.n7436 585
R13470 GND.n7439 GND.n4362 585
R13471 GND.n4366 GND.n4362 585
R13472 GND.n7441 GND.n7440 585
R13473 GND.n7442 GND.n7441 585
R13474 GND.n4363 GND.n4361 585
R13475 GND.n4361 GND.n4352 585
R13476 GND.n6163 GND.n4350 585
R13477 GND.n7448 GND.n4350 585
R13478 GND.n6165 GND.n6164 585
R13479 GND.n6165 GND.n4349 585
R13480 GND.n6167 GND.n6166 585
R13481 GND.n6166 GND.n4341 585
R13482 GND.n6168 GND.n5529 585
R13483 GND.n5529 GND.n4339 585
R13484 GND.n6170 GND.n6169 585
R13485 GND.n6171 GND.n6170 585
R13486 GND.n6162 GND.n5528 585
R13487 GND.n5528 GND.n4331 585
R13488 GND.n6161 GND.n6160 585
R13489 GND.n6160 GND.n4329 585
R13490 GND.n6159 GND.n5530 585
R13491 GND.n6159 GND.n6158 585
R13492 GND.n6139 GND.n5531 585
R13493 GND.n5531 GND.n4321 585
R13494 GND.n6140 GND.n5539 585
R13495 GND.n5539 GND.n4319 585
R13496 GND.n6142 GND.n6141 585
R13497 GND.n6143 GND.n6142 585
R13498 GND.n6138 GND.n5538 585
R13499 GND.n5538 GND.n4311 585
R13500 GND.n6137 GND.n6136 585
R13501 GND.n6136 GND.n4309 585
R13502 GND.n6135 GND.n5540 585
R13503 GND.n6135 GND.n6134 585
R13504 GND.n6121 GND.n5541 585
R13505 GND.n5541 GND.n4301 585
R13506 GND.n6122 GND.n5550 585
R13507 GND.n5550 GND.n4299 585
R13508 GND.n6124 GND.n6123 585
R13509 GND.n6125 GND.n6124 585
R13510 GND.n6120 GND.n5549 585
R13511 GND.n5549 GND.n5548 585
R13512 GND.n6119 GND.n6118 585
R13513 GND.n6118 GND.n4277 585
R13514 GND.n6117 GND.n5551 585
R13515 GND.n6117 GND.n6116 585
R13516 GND.n4261 GND.n4260 585
R13517 GND.n4265 GND.n4261 585
R13518 GND.n7493 GND.n7492 585
R13519 GND.n7492 GND.n7491 585
R13520 GND.n7494 GND.n4258 585
R13521 GND.n4262 GND.n4258 585
R13522 GND.n7496 GND.n7495 585
R13523 GND.n7497 GND.n7496 585
R13524 GND.n4259 GND.n4257 585
R13525 GND.n4257 GND.n4248 585
R13526 GND.n6060 GND.n4246 585
R13527 GND.n7503 GND.n4246 585
R13528 GND.n6062 GND.n6061 585
R13529 GND.n6062 GND.n4245 585
R13530 GND.n6064 GND.n6063 585
R13531 GND.n6063 GND.n4237 585
R13532 GND.n6065 GND.n5562 585
R13533 GND.n5562 GND.n4235 585
R13534 GND.n6067 GND.n6066 585
R13535 GND.n6068 GND.n6067 585
R13536 GND.n6059 GND.n5561 585
R13537 GND.n5561 GND.n5559 585
R13538 GND.n6058 GND.n6057 585
R13539 GND.n6057 GND.n4226 585
R13540 GND.n6056 GND.n5563 585
R13541 GND.n6056 GND.n6055 585
R13542 GND.n6036 GND.n5564 585
R13543 GND.n5564 GND.n4218 585
R13544 GND.n6037 GND.n5572 585
R13545 GND.n5572 GND.n4216 585
R13546 GND.n6039 GND.n6038 585
R13547 GND.n6040 GND.n6039 585
R13548 GND.n6035 GND.n5571 585
R13549 GND.n5571 GND.n4208 585
R13550 GND.n6034 GND.n6033 585
R13551 GND.n6033 GND.n4206 585
R13552 GND.n6032 GND.n5573 585
R13553 GND.n6032 GND.n6031 585
R13554 GND.n6018 GND.n5574 585
R13555 GND.n5576 GND.n5574 585
R13556 GND.n6019 GND.n5583 585
R13557 GND.n5583 GND.n4197 585
R13558 GND.n6021 GND.n6020 585
R13559 GND.n6022 GND.n6021 585
R13560 GND.n6017 GND.n5582 585
R13561 GND.n5582 GND.n4176 585
R13562 GND.n6016 GND.n6015 585
R13563 GND.n6015 GND.n4174 585
R13564 GND.n6014 GND.n5584 585
R13565 GND.n6014 GND.n6013 585
R13566 GND.n4158 GND.n4157 585
R13567 GND.n4162 GND.n4158 585
R13568 GND.n7548 GND.n7547 585
R13569 GND.n7547 GND.n7546 585
R13570 GND.n7549 GND.n4155 585
R13571 GND.n4159 GND.n4155 585
R13572 GND.n7551 GND.n7550 585
R13573 GND.n7552 GND.n7551 585
R13574 GND.n4156 GND.n4154 585
R13575 GND.n4154 GND.n4145 585
R13576 GND.n5957 GND.n4143 585
R13577 GND.n7558 GND.n4143 585
R13578 GND.n5959 GND.n5958 585
R13579 GND.n5959 GND.n4142 585
R13580 GND.n5961 GND.n5960 585
R13581 GND.n5960 GND.n4134 585
R13582 GND.n5962 GND.n5594 585
R13583 GND.n5594 GND.n4132 585
R13584 GND.n5964 GND.n5963 585
R13585 GND.n5965 GND.n5964 585
R13586 GND.n5956 GND.n5593 585
R13587 GND.n5593 GND.n4124 585
R13588 GND.n5955 GND.n5954 585
R13589 GND.n5954 GND.n4122 585
R13590 GND.n5953 GND.n5595 585
R13591 GND.n5953 GND.n5952 585
R13592 GND.n5933 GND.n5596 585
R13593 GND.n5596 GND.n4114 585
R13594 GND.n5934 GND.n5604 585
R13595 GND.n5604 GND.n4112 585
R13596 GND.n5936 GND.n5935 585
R13597 GND.n5937 GND.n5936 585
R13598 GND.n5932 GND.n5603 585
R13599 GND.n5603 GND.n4104 585
R13600 GND.n5931 GND.n5930 585
R13601 GND.n5930 GND.n4102 585
R13602 GND.n5929 GND.n5605 585
R13603 GND.n5929 GND.n5928 585
R13604 GND.n5915 GND.n5606 585
R13605 GND.n5606 GND.n4094 585
R13606 GND.n5916 GND.n5614 585
R13607 GND.n5614 GND.n4092 585
R13608 GND.n5918 GND.n5917 585
R13609 GND.n5919 GND.n5918 585
R13610 GND.n5914 GND.n5613 585
R13611 GND.n5613 GND.n4071 585
R13612 GND.n5913 GND.n5912 585
R13613 GND.n5912 GND.n4069 585
R13614 GND.n5911 GND.n5615 585
R13615 GND.n5911 GND.n5910 585
R13616 GND.n4053 GND.n4052 585
R13617 GND.n4057 GND.n4053 585
R13618 GND.n7603 GND.n7602 585
R13619 GND.n7602 GND.n7601 585
R13620 GND.n7604 GND.n4050 585
R13621 GND.n4054 GND.n4050 585
R13622 GND.n7606 GND.n7605 585
R13623 GND.n7607 GND.n7606 585
R13624 GND.n4051 GND.n4049 585
R13625 GND.n4049 GND.n4040 585
R13626 GND.n5854 GND.n4038 585
R13627 GND.n7613 GND.n4038 585
R13628 GND.n5856 GND.n5855 585
R13629 GND.n5856 GND.n4037 585
R13630 GND.n5858 GND.n5857 585
R13631 GND.n5857 GND.n4029 585
R13632 GND.n5859 GND.n5625 585
R13633 GND.n5625 GND.n4027 585
R13634 GND.n5861 GND.n5860 585
R13635 GND.n5862 GND.n5861 585
R13636 GND.n5853 GND.n5624 585
R13637 GND.n5624 GND.n4019 585
R13638 GND.n5852 GND.n5851 585
R13639 GND.n5851 GND.n4017 585
R13640 GND.n5850 GND.n5626 585
R13641 GND.n5850 GND.n5849 585
R13642 GND.n5830 GND.n5627 585
R13643 GND.n5627 GND.n4009 585
R13644 GND.n5831 GND.n5635 585
R13645 GND.n5635 GND.n4007 585
R13646 GND.n5833 GND.n5832 585
R13647 GND.n5834 GND.n5833 585
R13648 GND.n5829 GND.n5634 585
R13649 GND.n5634 GND.n3999 585
R13650 GND.n5828 GND.n5827 585
R13651 GND.n5827 GND.n3997 585
R13652 GND.n5826 GND.n5636 585
R13653 GND.n5826 GND.n5825 585
R13654 GND.n5812 GND.n5637 585
R13655 GND.n5637 GND.n3989 585
R13656 GND.n5813 GND.n5645 585
R13657 GND.n5645 GND.n3987 585
R13658 GND.n5815 GND.n5814 585
R13659 GND.n5816 GND.n5815 585
R13660 GND.n5811 GND.n5644 585
R13661 GND.n5644 GND.n3966 585
R13662 GND.n5810 GND.n5809 585
R13663 GND.n5809 GND.n3964 585
R13664 GND.n5808 GND.n5646 585
R13665 GND.n5808 GND.n5807 585
R13666 GND.n3949 GND.n3948 585
R13667 GND.n5798 GND.n3949 585
R13668 GND.n7658 GND.n7657 585
R13669 GND.n7657 GND.n7656 585
R13670 GND.n7659 GND.n3946 585
R13671 GND.n3950 GND.n3946 585
R13672 GND.n7661 GND.n7660 585
R13673 GND.n7662 GND.n7661 585
R13674 GND.n3947 GND.n3945 585
R13675 GND.n3945 GND.n3936 585
R13676 GND.n5750 GND.n3934 585
R13677 GND.n7668 GND.n3934 585
R13678 GND.n5752 GND.n5751 585
R13679 GND.n5752 GND.n3933 585
R13680 GND.n5754 GND.n5753 585
R13681 GND.n5753 GND.n3925 585
R13682 GND.n5755 GND.n5656 585
R13683 GND.n5656 GND.n3923 585
R13684 GND.n5757 GND.n5756 585
R13685 GND.n5758 GND.n5757 585
R13686 GND.n5749 GND.n5655 585
R13687 GND.n5655 GND.n3915 585
R13688 GND.n5748 GND.n5747 585
R13689 GND.n5747 GND.n3913 585
R13690 GND.n5746 GND.n5657 585
R13691 GND.n5746 GND.n5745 585
R13692 GND.n5726 GND.n5658 585
R13693 GND.n5658 GND.n3905 585
R13694 GND.n5727 GND.n5666 585
R13695 GND.n5666 GND.n3903 585
R13696 GND.n5729 GND.n5728 585
R13697 GND.n5730 GND.n5729 585
R13698 GND.n5725 GND.n5665 585
R13699 GND.n5665 GND.n3896 585
R13700 GND.n5724 GND.n5723 585
R13701 GND.n5723 GND.n3894 585
R13702 GND.n5722 GND.n5667 585
R13703 GND.n5722 GND.n5721 585
R13704 GND.n5708 GND.n5668 585
R13705 GND.n5668 GND.n3886 585
R13706 GND.n5709 GND.n5692 585
R13707 GND.n5692 GND.n3885 585
R13708 GND.n5711 GND.n5710 585
R13709 GND.n5712 GND.n5711 585
R13710 GND.n5707 GND.n5691 585
R13711 GND.n5691 GND.n2341 585
R13712 GND.n5706 GND.n5705 585
R13713 GND.n5705 GND.n2327 585
R13714 GND.n5704 GND.n5693 585
R13715 GND.n5704 GND.n5703 585
R13716 GND.n2313 GND.n2312 585
R13717 GND.n2316 GND.n2313 585
R13718 GND.n7769 GND.n7768 585
R13719 GND.n7768 GND.n7767 585
R13720 GND.n7770 GND.n2307 585
R13721 GND.n2314 GND.n2307 585
R13722 GND.n7772 GND.n7771 585
R13723 GND.n7773 GND.n7772 585
R13724 GND.n2311 GND.n2306 585
R13725 GND.n2306 GND.n2110 585
R13726 GND.n2310 GND.n2109 585
R13727 GND.n7779 GND.n2109 585
R13728 GND.n2309 GND.n2308 585
R13729 GND.n2308 GND.n2108 585
R13730 GND.n2096 GND.n2095 585
R13731 GND.n2099 GND.n2096 585
R13732 GND.n7788 GND.n7787 585
R13733 GND.n7787 GND.n7786 585
R13734 GND.n7789 GND.n2093 585
R13735 GND.n2097 GND.n2093 585
R13736 GND.n7791 GND.n7790 585
R13737 GND.n7792 GND.n7791 585
R13738 GND.n2094 GND.n2092 585
R13739 GND.n2092 GND.n2089 585
R13740 GND.n2290 GND.n2289 585
R13741 GND.n2291 GND.n2290 585
R13742 GND.n2078 GND.n2077 585
R13743 GND.n2081 GND.n2078 585
R13744 GND.n7802 GND.n7801 585
R13745 GND.n7801 GND.n7800 585
R13746 GND.n7803 GND.n2075 585
R13747 GND.n2079 GND.n2075 585
R13748 GND.n7805 GND.n7804 585
R13749 GND.n7806 GND.n7805 585
R13750 GND.n2076 GND.n2074 585
R13751 GND.n2074 GND.n2071 585
R13752 GND.n2277 GND.n2276 585
R13753 GND.n2278 GND.n2277 585
R13754 GND.n2060 GND.n2059 585
R13755 GND.n2063 GND.n2060 585
R13756 GND.n7816 GND.n7815 585
R13757 GND.n7815 GND.n7814 585
R13758 GND.n7817 GND.n2057 585
R13759 GND.n2061 GND.n2057 585
R13760 GND.n7819 GND.n7818 585
R13761 GND.n7820 GND.n7819 585
R13762 GND.n2058 GND.n2056 585
R13763 GND.n2056 GND.n2053 585
R13764 GND.n2264 GND.n2263 585
R13765 GND.n2265 GND.n2264 585
R13766 GND.n2042 GND.n2041 585
R13767 GND.n2045 GND.n2042 585
R13768 GND.n7830 GND.n7829 585
R13769 GND.n7829 GND.n7828 585
R13770 GND.n7831 GND.n2039 585
R13771 GND.n2043 GND.n2039 585
R13772 GND.n7833 GND.n7832 585
R13773 GND.n7834 GND.n7833 585
R13774 GND.n2040 GND.n2038 585
R13775 GND.n2038 GND.n2035 585
R13776 GND.n2251 GND.n2250 585
R13777 GND.n2252 GND.n2251 585
R13778 GND.n2024 GND.n2023 585
R13779 GND.n2027 GND.n2024 585
R13780 GND.n7844 GND.n7843 585
R13781 GND.n7843 GND.n7842 585
R13782 GND.n7845 GND.n2021 585
R13783 GND.n2021 GND.n2019 585
R13784 GND.n7847 GND.n7846 585
R13785 GND.n7848 GND.n7847 585
R13786 GND.n2022 GND.n2020 585
R13787 GND.n2020 GND.n2017 585
R13788 GND.n2239 GND.n2238 585
R13789 GND.n2240 GND.n2239 585
R13790 GND.n2006 GND.n2005 585
R13791 GND.n2009 GND.n2006 585
R13792 GND.n7858 GND.n7857 585
R13793 GND.n7857 GND.n7856 585
R13794 GND.n7859 GND.n2003 585
R13795 GND.n2003 GND.n2001 585
R13796 GND.n7861 GND.n7860 585
R13797 GND.n7862 GND.n7861 585
R13798 GND.n2004 GND.n2002 585
R13799 GND.n2002 GND.n1999 585
R13800 GND.n2226 GND.n2225 585
R13801 GND.n2227 GND.n2226 585
R13802 GND.n1988 GND.n1987 585
R13803 GND.n1991 GND.n1988 585
R13804 GND.n7872 GND.n7871 585
R13805 GND.n7871 GND.n7870 585
R13806 GND.n7873 GND.n1985 585
R13807 GND.n1985 GND.n1983 585
R13808 GND.n7875 GND.n7874 585
R13809 GND.n7876 GND.n7875 585
R13810 GND.n1986 GND.n1984 585
R13811 GND.n1984 GND.n1981 585
R13812 GND.n2213 GND.n2212 585
R13813 GND.n2214 GND.n2213 585
R13814 GND.n1970 GND.n1969 585
R13815 GND.n1973 GND.n1970 585
R13816 GND.n7886 GND.n7885 585
R13817 GND.n7885 GND.n7884 585
R13818 GND.n7887 GND.n1967 585
R13819 GND.n1967 GND.n1965 585
R13820 GND.n7889 GND.n7888 585
R13821 GND.n7890 GND.n7889 585
R13822 GND.n1968 GND.n1966 585
R13823 GND.n2202 GND.n1966 585
R13824 GND.n1954 GND.n1953 585
R13825 GND.n1955 GND.n1954 585
R13826 GND.n7899 GND.n7898 585
R13827 GND.n7898 GND.n7897 585
R13828 GND.n7900 GND.n1951 585
R13829 GND.n2195 GND.n1951 585
R13830 GND.n7902 GND.n7901 585
R13831 GND.n7903 GND.n7902 585
R13832 GND.n1952 GND.n1950 585
R13833 GND.n1950 GND.n1947 585
R13834 GND.n2189 GND.n2188 585
R13835 GND.n2190 GND.n2189 585
R13836 GND.n1935 GND.n1934 585
R13837 GND.n2186 GND.n1935 585
R13838 GND.n7913 GND.n7912 585
R13839 GND.n7912 GND.n7911 585
R13840 GND.n7914 GND.n1908 585
R13841 GND.n1936 GND.n1908 585
R13842 GND.n7970 GND.n7969 585
R13843 GND.n7968 GND.n1907 585
R13844 GND.n7967 GND.n1906 585
R13845 GND.n7972 GND.n1906 585
R13846 GND.n7966 GND.n7965 585
R13847 GND.n7964 GND.n7963 585
R13848 GND.n7962 GND.n7961 585
R13849 GND.n7960 GND.n7959 585
R13850 GND.n7958 GND.n7957 585
R13851 GND.n7956 GND.n7955 585
R13852 GND.n7954 GND.n7953 585
R13853 GND.n7952 GND.n7951 585
R13854 GND.n7950 GND.n7949 585
R13855 GND.n7948 GND.n7947 585
R13856 GND.n7946 GND.n7945 585
R13857 GND.n7944 GND.n7943 585
R13858 GND.n7942 GND.n7941 585
R13859 GND.n7940 GND.n7939 585
R13860 GND.n7938 GND.n7937 585
R13861 GND.n7936 GND.n7935 585
R13862 GND.n7934 GND.n7933 585
R13863 GND.n7932 GND.n7931 585
R13864 GND.n7930 GND.n7929 585
R13865 GND.n7928 GND.n7927 585
R13866 GND.n7926 GND.n7925 585
R13867 GND.n7924 GND.n7923 585
R13868 GND.n7922 GND.n7921 585
R13869 GND.n7919 GND.n7918 585
R13870 GND.n1875 GND.n1874 585
R13871 GND.n7975 GND.n7974 585
R13872 GND.n7976 GND.n1873 585
R13873 GND.n2124 GND.n1871 585
R13874 GND.n2126 GND.n2125 585
R13875 GND.n2128 GND.n2127 585
R13876 GND.n2130 GND.n2129 585
R13877 GND.n2132 GND.n2131 585
R13878 GND.n2134 GND.n2133 585
R13879 GND.n2136 GND.n2135 585
R13880 GND.n2138 GND.n2137 585
R13881 GND.n2140 GND.n2139 585
R13882 GND.n2142 GND.n2141 585
R13883 GND.n2144 GND.n2143 585
R13884 GND.n2146 GND.n2145 585
R13885 GND.n2148 GND.n2147 585
R13886 GND.n2150 GND.n2149 585
R13887 GND.n2152 GND.n2151 585
R13888 GND.n2154 GND.n2153 585
R13889 GND.n2156 GND.n2155 585
R13890 GND.n2158 GND.n2157 585
R13891 GND.n2160 GND.n2159 585
R13892 GND.n2162 GND.n2161 585
R13893 GND.n2164 GND.n2163 585
R13894 GND.n2166 GND.n2165 585
R13895 GND.n2168 GND.n2167 585
R13896 GND.n2170 GND.n2169 585
R13897 GND.n2172 GND.n2171 585
R13898 GND.n2174 GND.n2173 585
R13899 GND.n2176 GND.n2175 585
R13900 GND.n2178 GND.n2177 585
R13901 GND.n2180 GND.n2179 585
R13902 GND.n4776 GND.n4775 585
R13903 GND.n4778 GND.n4777 585
R13904 GND.n4780 GND.n4779 585
R13905 GND.n4782 GND.n4781 585
R13906 GND.n4784 GND.n4783 585
R13907 GND.n4786 GND.n4785 585
R13908 GND.n4788 GND.n4787 585
R13909 GND.n4790 GND.n4789 585
R13910 GND.n4792 GND.n4791 585
R13911 GND.n4794 GND.n4793 585
R13912 GND.n4796 GND.n4795 585
R13913 GND.n4798 GND.n4797 585
R13914 GND.n4800 GND.n4799 585
R13915 GND.n4802 GND.n4801 585
R13916 GND.n4804 GND.n4803 585
R13917 GND.n4806 GND.n4805 585
R13918 GND.n4808 GND.n4807 585
R13919 GND.n4810 GND.n4809 585
R13920 GND.n4812 GND.n4811 585
R13921 GND.n4814 GND.n4813 585
R13922 GND.n4816 GND.n4815 585
R13923 GND.n4818 GND.n4817 585
R13924 GND.n4820 GND.n4819 585
R13925 GND.n4822 GND.n4821 585
R13926 GND.n4824 GND.n4823 585
R13927 GND.n4826 GND.n4825 585
R13928 GND.n4828 GND.n4827 585
R13929 GND.n4830 GND.n4829 585
R13930 GND.n4832 GND.n4831 585
R13931 GND.n7190 GND.n7189 585
R13932 GND.n7192 GND.n7191 585
R13933 GND.n7194 GND.n7193 585
R13934 GND.n7196 GND.n7195 585
R13935 GND.n7199 GND.n7198 585
R13936 GND.n7201 GND.n7200 585
R13937 GND.n7203 GND.n7202 585
R13938 GND.n7205 GND.n7204 585
R13939 GND.n7207 GND.n7206 585
R13940 GND.n7209 GND.n7208 585
R13941 GND.n7211 GND.n7210 585
R13942 GND.n7213 GND.n7212 585
R13943 GND.n7215 GND.n7214 585
R13944 GND.n7217 GND.n7216 585
R13945 GND.n7219 GND.n7218 585
R13946 GND.n7221 GND.n7220 585
R13947 GND.n7223 GND.n7222 585
R13948 GND.n7225 GND.n7224 585
R13949 GND.n7227 GND.n7226 585
R13950 GND.n7229 GND.n7228 585
R13951 GND.n7231 GND.n7230 585
R13952 GND.n7233 GND.n7232 585
R13953 GND.n7235 GND.n7234 585
R13954 GND.n7237 GND.n7236 585
R13955 GND.n7239 GND.n7238 585
R13956 GND.n7241 GND.n7240 585
R13957 GND.n7243 GND.n7242 585
R13958 GND.n7245 GND.n7244 585
R13959 GND.n7246 GND.n4732 585
R13960 GND.n7248 GND.n7247 585
R13961 GND.n7249 GND.n7248 585
R13962 GND.n4774 GND.n4763 585
R13963 GND.n4774 GND.n4700 585
R13964 GND.n4773 GND.n4767 585
R13965 GND.n4773 GND.n4772 585
R13966 GND.n4766 GND.n4764 585
R13967 GND.n4764 GND.n4689 585
R13968 GND.n4765 GND.n4688 585
R13969 GND.n7258 GND.n4688 585
R13970 GND.n4674 GND.n4673 585
R13971 GND.n4687 GND.n4674 585
R13972 GND.n7266 GND.n7265 585
R13973 GND.n7265 GND.n7264 585
R13974 GND.n7267 GND.n4625 585
R13975 GND.n4625 GND.n4623 585
R13976 GND.n7269 GND.n7268 585
R13977 GND.n7270 GND.n7269 585
R13978 GND.n4672 GND.n4624 585
R13979 GND.n4680 GND.n4624 585
R13980 GND.n4671 GND.n4670 585
R13981 GND.n4670 GND.n4614 585
R13982 GND.n4669 GND.n4613 585
R13983 GND.n7277 GND.n4613 585
R13984 GND.n4668 GND.n4667 585
R13985 GND.n4667 GND.n4666 585
R13986 GND.n4665 GND.n4606 585
R13987 GND.n7283 GND.n4606 585
R13988 GND.n4664 GND.n4663 585
R13989 GND.n4663 GND.n4605 585
R13990 GND.n4662 GND.n4626 585
R13991 GND.n4662 GND.n4661 585
R13992 GND.n4657 GND.n4656 585
R13993 GND.n4657 GND.n4597 585
R13994 GND.n4655 GND.n4596 585
R13995 GND.n7291 GND.n4596 585
R13996 GND.n4654 GND.n4653 585
R13997 GND.n4653 GND.n4595 585
R13998 GND.n4652 GND.n4588 585
R13999 GND.n7297 GND.n4588 585
R14000 GND.n4651 GND.n4650 585
R14001 GND.n4650 GND.n4587 585
R14002 GND.n4649 GND.n4627 585
R14003 GND.n4649 GND.n4648 585
R14004 GND.n4644 GND.n4643 585
R14005 GND.n4644 GND.n4579 585
R14006 GND.n4642 GND.n4578 585
R14007 GND.n7305 GND.n4578 585
R14008 GND.n4641 GND.n4640 585
R14009 GND.n4640 GND.n4577 585
R14010 GND.n4639 GND.n4570 585
R14011 GND.n7311 GND.n4570 585
R14012 GND.n4638 GND.n4637 585
R14013 GND.n4637 GND.n4569 585
R14014 GND.n4636 GND.n4628 585
R14015 GND.n4636 GND.n4635 585
R14016 GND.n4631 GND.n4630 585
R14017 GND.n4631 GND.n4558 585
R14018 GND.n4629 GND.n4557 585
R14019 GND.n7319 GND.n4557 585
R14020 GND.n4545 GND.n4544 585
R14021 GND.n4556 GND.n4545 585
R14022 GND.n7327 GND.n7326 585
R14023 GND.n7326 GND.n7325 585
R14024 GND.n7328 GND.n4542 585
R14025 GND.n4542 GND.n4540 585
R14026 GND.n7330 GND.n7329 585
R14027 GND.n7331 GND.n7330 585
R14028 GND.n4543 GND.n4541 585
R14029 GND.n4541 GND.n4538 585
R14030 GND.n6243 GND.n6242 585
R14031 GND.n6242 GND.n4529 585
R14032 GND.n6244 GND.n4528 585
R14033 GND.n7338 GND.n4528 585
R14034 GND.n6246 GND.n6245 585
R14035 GND.n6245 GND.n4527 585
R14036 GND.n6247 GND.n4520 585
R14037 GND.n7344 GND.n4520 585
R14038 GND.n6249 GND.n6248 585
R14039 GND.n6249 GND.n4519 585
R14040 GND.n6254 GND.n6241 585
R14041 GND.n6254 GND.n6253 585
R14042 GND.n6256 GND.n6255 585
R14043 GND.n6255 GND.n4511 585
R14044 GND.n6257 GND.n4510 585
R14045 GND.n7352 GND.n4510 585
R14046 GND.n6259 GND.n6258 585
R14047 GND.n6258 GND.n4509 585
R14048 GND.n6260 GND.n4502 585
R14049 GND.n7358 GND.n4502 585
R14050 GND.n6262 GND.n6261 585
R14051 GND.n6262 GND.n4501 585
R14052 GND.n6267 GND.n6240 585
R14053 GND.n6267 GND.n6266 585
R14054 GND.n6269 GND.n6268 585
R14055 GND.n6268 GND.n4493 585
R14056 GND.n6270 GND.n4492 585
R14057 GND.n7366 GND.n4492 585
R14058 GND.n6272 GND.n6271 585
R14059 GND.n6271 GND.n4491 585
R14060 GND.n6273 GND.n4484 585
R14061 GND.n7372 GND.n4484 585
R14062 GND.n6275 GND.n6274 585
R14063 GND.n6275 GND.n4483 585
R14064 GND.n6280 GND.n6239 585
R14065 GND.n6280 GND.n6279 585
R14066 GND.n6282 GND.n6281 585
R14067 GND.n6281 GND.n4475 585
R14068 GND.n6283 GND.n4474 585
R14069 GND.n7380 GND.n4474 585
R14070 GND.n6285 GND.n6284 585
R14071 GND.n6284 GND.n4473 585
R14072 GND.n6286 GND.n4466 585
R14073 GND.n7386 GND.n4466 585
R14074 GND.n6288 GND.n6287 585
R14075 GND.n6288 GND.n4465 585
R14076 GND.n6292 GND.n6238 585
R14077 GND.n6292 GND.n6291 585
R14078 GND.n6294 GND.n6293 585
R14079 GND.n6293 GND.n4457 585
R14080 GND.n6295 GND.n4456 585
R14081 GND.n7394 GND.n4456 585
R14082 GND.n6297 GND.n6296 585
R14083 GND.n6296 GND.n4449 585
R14084 GND.n6298 GND.n4448 585
R14085 GND.n7400 GND.n4448 585
R14086 GND.n6299 GND.n5506 585
R14087 GND.n5506 GND.n4447 585
R14088 GND.n6301 GND.n6300 585
R14089 GND.n6303 GND.n6301 585
R14090 GND.n6237 GND.n5505 585
R14091 GND.n5505 GND.n4436 585
R14092 GND.n6236 GND.n6235 585
R14093 GND.n6235 GND.n4422 585
R14094 GND.n6234 GND.n6233 585
R14095 GND.n6234 GND.n5499 585
R14096 GND.n6232 GND.n5497 585
R14097 GND.n6311 GND.n5497 585
R14098 GND.n6231 GND.n6230 585
R14099 GND.n6230 GND.n4415 585
R14100 GND.n6229 GND.n5507 585
R14101 GND.n6229 GND.n6228 585
R14102 GND.n6214 GND.n5508 585
R14103 GND.n5509 GND.n5508 585
R14104 GND.n6216 GND.n6215 585
R14105 GND.n6215 GND.n4406 585
R14106 GND.n6217 GND.n5515 585
R14107 GND.n5515 GND.n4404 585
R14108 GND.n6219 GND.n6218 585
R14109 GND.n6220 GND.n6219 585
R14110 GND.n6213 GND.n5514 585
R14111 GND.n5514 GND.n4383 585
R14112 GND.n6212 GND.n6211 585
R14113 GND.n6211 GND.n4381 585
R14114 GND.n6210 GND.n5516 585
R14115 GND.n6210 GND.n6209 585
R14116 GND.n5519 GND.n5518 585
R14117 GND.n5519 GND.n4369 585
R14118 GND.n5517 GND.n4367 585
R14119 GND.n7436 GND.n4367 585
R14120 GND.n4358 GND.n4357 585
R14121 GND.n4366 GND.n4358 585
R14122 GND.n7444 GND.n7443 585
R14123 GND.n7443 GND.n7442 585
R14124 GND.n7445 GND.n4355 585
R14125 GND.n4355 GND.n4352 585
R14126 GND.n7447 GND.n7446 585
R14127 GND.n7448 GND.n7447 585
R14128 GND.n4356 GND.n4354 585
R14129 GND.n4354 GND.n4349 585
R14130 GND.n6149 GND.n6148 585
R14131 GND.n6149 GND.n4341 585
R14132 GND.n6151 GND.n6150 585
R14133 GND.n6150 GND.n4339 585
R14134 GND.n6152 GND.n5527 585
R14135 GND.n6171 GND.n5527 585
R14136 GND.n6154 GND.n6153 585
R14137 GND.n6153 GND.n4331 585
R14138 GND.n6155 GND.n5534 585
R14139 GND.n5534 GND.n4329 585
R14140 GND.n6157 GND.n6156 585
R14141 GND.n6158 GND.n6157 585
R14142 GND.n6147 GND.n5533 585
R14143 GND.n5533 GND.n4321 585
R14144 GND.n6146 GND.n6145 585
R14145 GND.n6145 GND.n4319 585
R14146 GND.n6144 GND.n5535 585
R14147 GND.n6144 GND.n6143 585
R14148 GND.n6130 GND.n5536 585
R14149 GND.n5536 GND.n4311 585
R14150 GND.n6131 GND.n5544 585
R14151 GND.n5544 GND.n4309 585
R14152 GND.n6133 GND.n6132 585
R14153 GND.n6134 GND.n6133 585
R14154 GND.n6129 GND.n5543 585
R14155 GND.n5543 GND.n4301 585
R14156 GND.n6128 GND.n6127 585
R14157 GND.n6127 GND.n4299 585
R14158 GND.n6126 GND.n5545 585
R14159 GND.n6126 GND.n6125 585
R14160 GND.n6112 GND.n5546 585
R14161 GND.n5548 GND.n5546 585
R14162 GND.n6113 GND.n6109 585
R14163 GND.n6109 GND.n4277 585
R14164 GND.n6115 GND.n6114 585
R14165 GND.n6116 GND.n6115 585
R14166 GND.n6111 GND.n6108 585
R14167 GND.n6108 GND.n4265 585
R14168 GND.n6110 GND.n4263 585
R14169 GND.n7491 GND.n4263 585
R14170 GND.n4254 GND.n4253 585
R14171 GND.n4262 GND.n4254 585
R14172 GND.n7499 GND.n7498 585
R14173 GND.n7498 GND.n7497 585
R14174 GND.n7500 GND.n4251 585
R14175 GND.n4251 GND.n4248 585
R14176 GND.n7502 GND.n7501 585
R14177 GND.n7503 GND.n7502 585
R14178 GND.n4252 GND.n4250 585
R14179 GND.n4250 GND.n4245 585
R14180 GND.n6046 GND.n6045 585
R14181 GND.n6046 GND.n4237 585
R14182 GND.n6048 GND.n6047 585
R14183 GND.n6047 GND.n4235 585
R14184 GND.n6049 GND.n5560 585
R14185 GND.n6068 GND.n5560 585
R14186 GND.n6051 GND.n6050 585
R14187 GND.n6050 GND.n5559 585
R14188 GND.n6052 GND.n5567 585
R14189 GND.n5567 GND.n4226 585
R14190 GND.n6054 GND.n6053 585
R14191 GND.n6055 GND.n6054 585
R14192 GND.n6044 GND.n5566 585
R14193 GND.n5566 GND.n4218 585
R14194 GND.n6043 GND.n6042 585
R14195 GND.n6042 GND.n4216 585
R14196 GND.n6041 GND.n5568 585
R14197 GND.n6041 GND.n6040 585
R14198 GND.n6027 GND.n5569 585
R14199 GND.n5569 GND.n4208 585
R14200 GND.n6028 GND.n5578 585
R14201 GND.n5578 GND.n4206 585
R14202 GND.n6030 GND.n6029 585
R14203 GND.n6031 GND.n6030 585
R14204 GND.n6026 GND.n5577 585
R14205 GND.n5577 GND.n5576 585
R14206 GND.n6025 GND.n6024 585
R14207 GND.n6024 GND.n4197 585
R14208 GND.n6023 GND.n5579 585
R14209 GND.n6023 GND.n6022 585
R14210 GND.n6009 GND.n5580 585
R14211 GND.n5580 GND.n4176 585
R14212 GND.n6010 GND.n6006 585
R14213 GND.n6006 GND.n4174 585
R14214 GND.n6012 GND.n6011 585
R14215 GND.n6013 GND.n6012 585
R14216 GND.n6008 GND.n6005 585
R14217 GND.n6005 GND.n4162 585
R14218 GND.n6007 GND.n4160 585
R14219 GND.n7546 GND.n4160 585
R14220 GND.n4151 GND.n4150 585
R14221 GND.n4159 GND.n4151 585
R14222 GND.n7554 GND.n7553 585
R14223 GND.n7553 GND.n7552 585
R14224 GND.n7555 GND.n4148 585
R14225 GND.n4148 GND.n4145 585
R14226 GND.n7557 GND.n7556 585
R14227 GND.n7558 GND.n7557 585
R14228 GND.n4149 GND.n4147 585
R14229 GND.n4147 GND.n4142 585
R14230 GND.n5943 GND.n5942 585
R14231 GND.n5943 GND.n4134 585
R14232 GND.n5945 GND.n5944 585
R14233 GND.n5944 GND.n4132 585
R14234 GND.n5946 GND.n5592 585
R14235 GND.n5965 GND.n5592 585
R14236 GND.n5948 GND.n5947 585
R14237 GND.n5947 GND.n4124 585
R14238 GND.n5949 GND.n5599 585
R14239 GND.n5599 GND.n4122 585
R14240 GND.n5951 GND.n5950 585
R14241 GND.n5952 GND.n5951 585
R14242 GND.n5941 GND.n5598 585
R14243 GND.n5598 GND.n4114 585
R14244 GND.n5940 GND.n5939 585
R14245 GND.n5939 GND.n4112 585
R14246 GND.n5938 GND.n5600 585
R14247 GND.n5938 GND.n5937 585
R14248 GND.n5924 GND.n5601 585
R14249 GND.n5601 GND.n4104 585
R14250 GND.n5925 GND.n5609 585
R14251 GND.n5609 GND.n4102 585
R14252 GND.n5927 GND.n5926 585
R14253 GND.n5928 GND.n5927 585
R14254 GND.n5923 GND.n5608 585
R14255 GND.n5608 GND.n4094 585
R14256 GND.n5922 GND.n5921 585
R14257 GND.n5921 GND.n4092 585
R14258 GND.n5920 GND.n5610 585
R14259 GND.n5920 GND.n5919 585
R14260 GND.n5906 GND.n5611 585
R14261 GND.n5611 GND.n4071 585
R14262 GND.n5907 GND.n5903 585
R14263 GND.n5903 GND.n4069 585
R14264 GND.n5909 GND.n5908 585
R14265 GND.n5910 GND.n5909 585
R14266 GND.n5905 GND.n5902 585
R14267 GND.n5902 GND.n4057 585
R14268 GND.n5904 GND.n4055 585
R14269 GND.n7601 GND.n4055 585
R14270 GND.n4046 GND.n4045 585
R14271 GND.n4054 GND.n4046 585
R14272 GND.n7609 GND.n7608 585
R14273 GND.n7608 GND.n7607 585
R14274 GND.n7610 GND.n4043 585
R14275 GND.n4043 GND.n4040 585
R14276 GND.n7612 GND.n7611 585
R14277 GND.n7613 GND.n7612 585
R14278 GND.n4044 GND.n4042 585
R14279 GND.n4042 GND.n4037 585
R14280 GND.n5840 GND.n5839 585
R14281 GND.n5840 GND.n4029 585
R14282 GND.n5842 GND.n5841 585
R14283 GND.n5841 GND.n4027 585
R14284 GND.n5843 GND.n5623 585
R14285 GND.n5862 GND.n5623 585
R14286 GND.n5845 GND.n5844 585
R14287 GND.n5844 GND.n4019 585
R14288 GND.n5846 GND.n5630 585
R14289 GND.n5630 GND.n4017 585
R14290 GND.n5848 GND.n5847 585
R14291 GND.n5849 GND.n5848 585
R14292 GND.n5838 GND.n5629 585
R14293 GND.n5629 GND.n4009 585
R14294 GND.n5837 GND.n5836 585
R14295 GND.n5836 GND.n4007 585
R14296 GND.n5835 GND.n5631 585
R14297 GND.n5835 GND.n5834 585
R14298 GND.n5821 GND.n5632 585
R14299 GND.n5632 GND.n3999 585
R14300 GND.n5822 GND.n5640 585
R14301 GND.n5640 GND.n3997 585
R14302 GND.n5824 GND.n5823 585
R14303 GND.n5825 GND.n5824 585
R14304 GND.n5820 GND.n5639 585
R14305 GND.n5639 GND.n3989 585
R14306 GND.n5819 GND.n5818 585
R14307 GND.n5818 GND.n3987 585
R14308 GND.n5817 GND.n5641 585
R14309 GND.n5817 GND.n5816 585
R14310 GND.n5803 GND.n5642 585
R14311 GND.n5642 GND.n3966 585
R14312 GND.n5804 GND.n5800 585
R14313 GND.n5800 GND.n3964 585
R14314 GND.n5806 GND.n5805 585
R14315 GND.n5807 GND.n5806 585
R14316 GND.n5802 GND.n5799 585
R14317 GND.n5799 GND.n5798 585
R14318 GND.n5801 GND.n3951 585
R14319 GND.n7656 GND.n3951 585
R14320 GND.n3942 GND.n3941 585
R14321 GND.n3950 GND.n3942 585
R14322 GND.n7664 GND.n7663 585
R14323 GND.n7663 GND.n7662 585
R14324 GND.n7665 GND.n3939 585
R14325 GND.n3939 GND.n3936 585
R14326 GND.n7667 GND.n7666 585
R14327 GND.n7668 GND.n7667 585
R14328 GND.n3940 GND.n3938 585
R14329 GND.n3938 GND.n3933 585
R14330 GND.n5736 GND.n5735 585
R14331 GND.n5736 GND.n3925 585
R14332 GND.n5738 GND.n5737 585
R14333 GND.n5737 GND.n3923 585
R14334 GND.n5739 GND.n5654 585
R14335 GND.n5758 GND.n5654 585
R14336 GND.n5741 GND.n5740 585
R14337 GND.n5740 GND.n3915 585
R14338 GND.n5742 GND.n5661 585
R14339 GND.n5661 GND.n3913 585
R14340 GND.n5744 GND.n5743 585
R14341 GND.n5745 GND.n5744 585
R14342 GND.n5734 GND.n5660 585
R14343 GND.n5660 GND.n3905 585
R14344 GND.n5733 GND.n5732 585
R14345 GND.n5732 GND.n3903 585
R14346 GND.n5731 GND.n5662 585
R14347 GND.n5731 GND.n5730 585
R14348 GND.n5717 GND.n5663 585
R14349 GND.n5663 GND.n3896 585
R14350 GND.n5718 GND.n5687 585
R14351 GND.n5687 GND.n3894 585
R14352 GND.n5720 GND.n5719 585
R14353 GND.n5721 GND.n5720 585
R14354 GND.n5716 GND.n5686 585
R14355 GND.n5686 GND.n3886 585
R14356 GND.n5715 GND.n5714 585
R14357 GND.n5714 GND.n3885 585
R14358 GND.n5713 GND.n5688 585
R14359 GND.n5713 GND.n5712 585
R14360 GND.n5699 GND.n5689 585
R14361 GND.n5689 GND.n2341 585
R14362 GND.n5700 GND.n5696 585
R14363 GND.n5696 GND.n2327 585
R14364 GND.n5702 GND.n5701 585
R14365 GND.n5703 GND.n5702 585
R14366 GND.n5698 GND.n5695 585
R14367 GND.n5695 GND.n2316 585
R14368 GND.n5697 GND.n2315 585
R14369 GND.n7767 GND.n2315 585
R14370 GND.n2303 GND.n2302 585
R14371 GND.n2314 GND.n2303 585
R14372 GND.n7775 GND.n7774 585
R14373 GND.n7774 GND.n7773 585
R14374 GND.n7776 GND.n2112 585
R14375 GND.n2112 GND.n2110 585
R14376 GND.n7778 GND.n7777 585
R14377 GND.n7779 GND.n7778 585
R14378 GND.n2301 GND.n2111 585
R14379 GND.n2111 GND.n2108 585
R14380 GND.n2300 GND.n2299 585
R14381 GND.n2299 GND.n2099 585
R14382 GND.n2298 GND.n2098 585
R14383 GND.n7786 GND.n2098 585
R14384 GND.n2297 GND.n2296 585
R14385 GND.n2296 GND.n2097 585
R14386 GND.n2295 GND.n2090 585
R14387 GND.n7792 GND.n2090 585
R14388 GND.n2294 GND.n2293 585
R14389 GND.n2293 GND.n2089 585
R14390 GND.n2292 GND.n2113 585
R14391 GND.n2292 GND.n2291 585
R14392 GND.n2287 GND.n2286 585
R14393 GND.n2287 GND.n2081 585
R14394 GND.n2285 GND.n2080 585
R14395 GND.n7800 GND.n2080 585
R14396 GND.n2284 GND.n2283 585
R14397 GND.n2283 GND.n2079 585
R14398 GND.n2282 GND.n2072 585
R14399 GND.n7806 GND.n2072 585
R14400 GND.n2281 GND.n2280 585
R14401 GND.n2280 GND.n2071 585
R14402 GND.n2279 GND.n2114 585
R14403 GND.n2279 GND.n2278 585
R14404 GND.n2274 GND.n2273 585
R14405 GND.n2274 GND.n2063 585
R14406 GND.n2272 GND.n2062 585
R14407 GND.n7814 GND.n2062 585
R14408 GND.n2271 GND.n2270 585
R14409 GND.n2270 GND.n2061 585
R14410 GND.n2269 GND.n2054 585
R14411 GND.n7820 GND.n2054 585
R14412 GND.n2268 GND.n2267 585
R14413 GND.n2267 GND.n2053 585
R14414 GND.n2266 GND.n2115 585
R14415 GND.n2266 GND.n2265 585
R14416 GND.n2261 GND.n2260 585
R14417 GND.n2261 GND.n2045 585
R14418 GND.n2259 GND.n2044 585
R14419 GND.n7828 GND.n2044 585
R14420 GND.n2258 GND.n2257 585
R14421 GND.n2257 GND.n2043 585
R14422 GND.n2256 GND.n2036 585
R14423 GND.n7834 GND.n2036 585
R14424 GND.n2255 GND.n2254 585
R14425 GND.n2254 GND.n2035 585
R14426 GND.n2253 GND.n2116 585
R14427 GND.n2253 GND.n2252 585
R14428 GND.n2249 GND.n2248 585
R14429 GND.n2249 GND.n2027 585
R14430 GND.n2247 GND.n2026 585
R14431 GND.n7842 GND.n2026 585
R14432 GND.n2246 GND.n2245 585
R14433 GND.n2245 GND.n2019 585
R14434 GND.n2244 GND.n2018 585
R14435 GND.n7848 GND.n2018 585
R14436 GND.n2243 GND.n2242 585
R14437 GND.n2242 GND.n2017 585
R14438 GND.n2241 GND.n2117 585
R14439 GND.n2241 GND.n2240 585
R14440 GND.n2236 GND.n2235 585
R14441 GND.n2236 GND.n2009 585
R14442 GND.n2234 GND.n2008 585
R14443 GND.n7856 GND.n2008 585
R14444 GND.n2233 GND.n2232 585
R14445 GND.n2232 GND.n2001 585
R14446 GND.n2231 GND.n2000 585
R14447 GND.n7862 GND.n2000 585
R14448 GND.n2230 GND.n2229 585
R14449 GND.n2229 GND.n1999 585
R14450 GND.n2228 GND.n2118 585
R14451 GND.n2228 GND.n2227 585
R14452 GND.n2223 GND.n2222 585
R14453 GND.n2223 GND.n1991 585
R14454 GND.n2221 GND.n1990 585
R14455 GND.n7870 GND.n1990 585
R14456 GND.n2220 GND.n2219 585
R14457 GND.n2219 GND.n1983 585
R14458 GND.n2218 GND.n1982 585
R14459 GND.n7876 GND.n1982 585
R14460 GND.n2217 GND.n2216 585
R14461 GND.n2216 GND.n1981 585
R14462 GND.n2215 GND.n2119 585
R14463 GND.n2215 GND.n2214 585
R14464 GND.n2210 GND.n2209 585
R14465 GND.n2210 GND.n1973 585
R14466 GND.n2208 GND.n1972 585
R14467 GND.n7884 GND.n1972 585
R14468 GND.n2207 GND.n2206 585
R14469 GND.n2206 GND.n1965 585
R14470 GND.n2205 GND.n1964 585
R14471 GND.n7890 GND.n1964 585
R14472 GND.n2204 GND.n2203 585
R14473 GND.n2203 GND.n2202 585
R14474 GND.n2200 GND.n2199 585
R14475 GND.n2200 GND.n1955 585
R14476 GND.n2198 GND.n1956 585
R14477 GND.n7897 GND.n1956 585
R14478 GND.n2197 GND.n2196 585
R14479 GND.n2196 GND.n2195 585
R14480 GND.n2194 GND.n1948 585
R14481 GND.n7903 GND.n1948 585
R14482 GND.n2193 GND.n2192 585
R14483 GND.n2192 GND.n1947 585
R14484 GND.n2191 GND.n2120 585
R14485 GND.n2191 GND.n2190 585
R14486 GND.n2185 GND.n2184 585
R14487 GND.n2186 GND.n2185 585
R14488 GND.n2183 GND.n1937 585
R14489 GND.n7911 GND.n1937 585
R14490 GND.n2182 GND.n2181 585
R14491 GND.n2181 GND.n1936 585
R14492 GND.n3840 GND.n1677 585
R14493 GND.n8026 GND.n1677 585
R14494 GND.n3842 GND.n3841 585
R14495 GND.n3843 GND.n3842 585
R14496 GND.n2364 GND.n2363 585
R14497 GND.n3830 GND.n2363 585
R14498 GND.n3836 GND.n3835 585
R14499 GND.n3835 GND.n3834 585
R14500 GND.n2367 GND.n2366 585
R14501 GND.n3828 GND.n2367 585
R14502 GND.n3814 GND.n2384 585
R14503 GND.n2384 GND.n2383 585
R14504 GND.n3816 GND.n3815 585
R14505 GND.n3817 GND.n3816 585
R14506 GND.n2385 GND.n2381 585
R14507 GND.n3804 GND.n2381 585
R14508 GND.n3809 GND.n3808 585
R14509 GND.n3808 GND.n3807 585
R14510 GND.n2388 GND.n2387 585
R14511 GND.n3801 GND.n2388 585
R14512 GND.n3788 GND.n2406 585
R14513 GND.n2406 GND.n2405 585
R14514 GND.n3790 GND.n3789 585
R14515 GND.n3791 GND.n3790 585
R14516 GND.n2407 GND.n2404 585
R14517 GND.n3778 GND.n2404 585
R14518 GND.n3783 GND.n3782 585
R14519 GND.n3782 GND.n3781 585
R14520 GND.n2410 GND.n2409 585
R14521 GND.n3776 GND.n2410 585
R14522 GND.n3763 GND.n2428 585
R14523 GND.n2428 GND.n2427 585
R14524 GND.n3765 GND.n3764 585
R14525 GND.n3766 GND.n3765 585
R14526 GND.n2429 GND.n2426 585
R14527 GND.n3753 GND.n2426 585
R14528 GND.n3758 GND.n3757 585
R14529 GND.n3757 GND.n3756 585
R14530 GND.n2432 GND.n2431 585
R14531 GND.n3750 GND.n2432 585
R14532 GND.n3737 GND.n2448 585
R14533 GND.n3473 GND.n2448 585
R14534 GND.n3739 GND.n3738 585
R14535 GND.n3740 GND.n3739 585
R14536 GND.n2449 GND.n2447 585
R14537 GND.n3726 GND.n2447 585
R14538 GND.n3732 GND.n3731 585
R14539 GND.n3731 GND.n3730 585
R14540 GND.n2452 GND.n2451 585
R14541 GND.n3724 GND.n2452 585
R14542 GND.n3711 GND.n2469 585
R14543 GND.n2469 GND.n2468 585
R14544 GND.n3713 GND.n3712 585
R14545 GND.n3714 GND.n3713 585
R14546 GND.n2470 GND.n2466 585
R14547 GND.n3701 GND.n2466 585
R14548 GND.n3706 GND.n3705 585
R14549 GND.n3705 GND.n3704 585
R14550 GND.n2473 GND.n2472 585
R14551 GND.n3698 GND.n2473 585
R14552 GND.n3685 GND.n2491 585
R14553 GND.n2491 GND.n2490 585
R14554 GND.n3687 GND.n3686 585
R14555 GND.n3688 GND.n3687 585
R14556 GND.n2492 GND.n2489 585
R14557 GND.n3675 GND.n2489 585
R14558 GND.n3680 GND.n3679 585
R14559 GND.n3679 GND.n3678 585
R14560 GND.n2495 GND.n2494 585
R14561 GND.n3673 GND.n2495 585
R14562 GND.n3660 GND.n2513 585
R14563 GND.n2513 GND.n2512 585
R14564 GND.n3662 GND.n3661 585
R14565 GND.n3663 GND.n3662 585
R14566 GND.n2514 GND.n2511 585
R14567 GND.n3650 GND.n2511 585
R14568 GND.n3655 GND.n3654 585
R14569 GND.n3654 GND.n3653 585
R14570 GND.n2517 GND.n2516 585
R14571 GND.n3647 GND.n2517 585
R14572 GND.n3634 GND.n2535 585
R14573 GND.n2535 GND.n2534 585
R14574 GND.n3636 GND.n3635 585
R14575 GND.n3637 GND.n3636 585
R14576 GND.n2536 GND.n2533 585
R14577 GND.n3623 GND.n2533 585
R14578 GND.n3629 GND.n3628 585
R14579 GND.n3628 GND.n3627 585
R14580 GND.n2539 GND.n2538 585
R14581 GND.n3621 GND.n2539 585
R14582 GND.n3608 GND.n2556 585
R14583 GND.n2556 GND.n2555 585
R14584 GND.n3610 GND.n3609 585
R14585 GND.n3611 GND.n3610 585
R14586 GND.n2557 GND.n2553 585
R14587 GND.n3598 GND.n2553 585
R14588 GND.n3603 GND.n3602 585
R14589 GND.n3602 GND.n3601 585
R14590 GND.n2560 GND.n2559 585
R14591 GND.n3595 GND.n2560 585
R14592 GND.n3582 GND.n2578 585
R14593 GND.n2578 GND.n2577 585
R14594 GND.n3584 GND.n3583 585
R14595 GND.n3585 GND.n3584 585
R14596 GND.n2579 GND.n2576 585
R14597 GND.n3572 GND.n2576 585
R14598 GND.n3577 GND.n3576 585
R14599 GND.n3576 GND.n3575 585
R14600 GND.n2582 GND.n2581 585
R14601 GND.n3570 GND.n2582 585
R14602 GND.n1551 GND.n1549 585
R14603 GND.n2588 GND.n1551 585
R14604 GND.n8118 GND.n8117 585
R14605 GND.n8117 GND.n8116 585
R14606 GND.n1550 GND.n1548 585
R14607 GND.n3559 GND.n1550 585
R14608 GND.n3555 GND.n3554 585
R14609 GND.n3556 GND.n3555 585
R14610 GND.n1540 GND.n1538 585
R14611 GND.n2600 GND.n1538 585
R14612 GND.n8122 GND.n8121 585
R14613 GND.n8123 GND.n8122 585
R14614 GND.n1539 GND.n1537 585
R14615 GND.n3542 GND.n1537 585
R14616 GND.n3325 GND.n3324 585
R14617 GND.n3325 GND.n2610 585
R14618 GND.n3326 GND.n1546 585
R14619 GND.n3327 GND.n3326 585
R14620 GND.n3323 GND.n3322 585
R14621 GND.n3323 GND.n2615 585
R14622 GND.n3321 GND.n2621 585
R14623 GND.n3321 GND.n3320 585
R14624 GND.n3291 GND.n2620 585
R14625 GND.n3308 GND.n2620 585
R14626 GND.n3292 GND.n2645 585
R14627 GND.n2645 GND.n2633 585
R14628 GND.n3294 GND.n3293 585
R14629 GND.n3295 GND.n3294 585
R14630 GND.n2646 GND.n2644 585
R14631 GND.n2644 GND.n2640 585
R14632 GND.n3286 GND.n3285 585
R14633 GND.n3285 GND.n3284 585
R14634 GND.n2649 GND.n2648 585
R14635 GND.n3269 GND.n2649 585
R14636 GND.n3254 GND.n2675 585
R14637 GND.n2675 GND.n2662 585
R14638 GND.n3256 GND.n3255 585
R14639 GND.n3257 GND.n3256 585
R14640 GND.n2676 GND.n2674 585
R14641 GND.n2674 GND.n2670 585
R14642 GND.n3249 GND.n3248 585
R14643 GND.n3248 GND.n3247 585
R14644 GND.n2679 GND.n2678 585
R14645 GND.n3232 GND.n2679 585
R14646 GND.n3217 GND.n2704 585
R14647 GND.n2704 GND.n2691 585
R14648 GND.n3219 GND.n3218 585
R14649 GND.n3220 GND.n3219 585
R14650 GND.n2705 GND.n2703 585
R14651 GND.n2703 GND.n2698 585
R14652 GND.n3212 GND.n3211 585
R14653 GND.n3211 GND.n3210 585
R14654 GND.n2708 GND.n2707 585
R14655 GND.n3195 GND.n2708 585
R14656 GND.n3180 GND.n2733 585
R14657 GND.n2733 GND.n2721 585
R14658 GND.n3182 GND.n3181 585
R14659 GND.n3183 GND.n3182 585
R14660 GND.n2734 GND.n2732 585
R14661 GND.n2732 GND.n2728 585
R14662 GND.n3175 GND.n3174 585
R14663 GND.n3174 GND.n3173 585
R14664 GND.n2737 GND.n2736 585
R14665 GND.n3158 GND.n2737 585
R14666 GND.n3142 GND.n2760 585
R14667 GND.n2760 GND.n2749 585
R14668 GND.n3144 GND.n3143 585
R14669 GND.n3145 GND.n3144 585
R14670 GND.n2761 GND.n2759 585
R14671 GND.n3122 GND.n2759 585
R14672 GND.n3137 GND.n3136 585
R14673 GND.n3136 GND.n3135 585
R14674 GND.n2764 GND.n2763 585
R14675 GND.n3119 GND.n2764 585
R14676 GND.n3104 GND.n2790 585
R14677 GND.n2790 GND.n2777 585
R14678 GND.n3106 GND.n3105 585
R14679 GND.n3107 GND.n3106 585
R14680 GND.n2791 GND.n2789 585
R14681 GND.n2789 GND.n2785 585
R14682 GND.n3099 GND.n3098 585
R14683 GND.n3098 GND.n3097 585
R14684 GND.n2794 GND.n2793 585
R14685 GND.n3082 GND.n2794 585
R14686 GND.n3067 GND.n2819 585
R14687 GND.n2819 GND.n2806 585
R14688 GND.n3069 GND.n3068 585
R14689 GND.n3070 GND.n3069 585
R14690 GND.n2820 GND.n2818 585
R14691 GND.n2818 GND.n2813 585
R14692 GND.n3062 GND.n3061 585
R14693 GND.n3061 GND.n3060 585
R14694 GND.n2823 GND.n2822 585
R14695 GND.n3045 GND.n2823 585
R14696 GND.n3034 GND.n3033 585
R14697 GND.n3035 GND.n3034 585
R14698 GND.n2844 GND.n2843 585
R14699 GND.n2843 GND.n2840 585
R14700 GND.n3029 GND.n3028 585
R14701 GND.n3028 GND.n3027 585
R14702 GND.n2847 GND.n2846 585
R14703 GND.n3018 GND.n2847 585
R14704 GND.n3001 GND.n2867 585
R14705 GND.n2867 GND.n2862 585
R14706 GND.n3003 GND.n3002 585
R14707 GND.n3004 GND.n3003 585
R14708 GND.n2868 GND.n2866 585
R14709 GND.n2875 GND.n2866 585
R14710 GND.n2996 GND.n2995 585
R14711 GND.n2995 GND.n2994 585
R14712 GND.n2871 GND.n2870 585
R14713 GND.n2873 GND.n2871 585
R14714 GND.n2977 GND.n2976 585
R14715 GND.n2978 GND.n2977 585
R14716 GND.n2887 GND.n2886 585
R14717 GND.n2886 GND.n2884 585
R14718 GND.n2972 GND.n2971 585
R14719 GND.n2971 GND.n2970 585
R14720 GND.n2890 GND.n2889 585
R14721 GND.n2892 GND.n2890 585
R14722 GND.n2960 GND.n2959 585
R14723 GND.n2961 GND.n2960 585
R14724 GND.n2907 GND.n2906 585
R14725 GND.n2906 GND.n2904 585
R14726 GND.n2955 GND.n2954 585
R14727 GND.n2954 GND.n2953 585
R14728 GND.n2910 GND.n2909 585
R14729 GND.n2912 GND.n2910 585
R14730 GND.n2943 GND.n2942 585
R14731 GND.n2944 GND.n2943 585
R14732 GND.n2937 GND.n2936 585
R14733 GND.n2936 GND.n2924 585
R14734 GND.n2938 GND.n1362 585
R14735 GND.n1362 GND.n1358 585
R14736 GND.n8360 GND.n8359 585
R14737 GND.n8358 GND.n1361 585
R14738 GND.n8357 GND.n1360 585
R14739 GND.n8362 GND.n1360 585
R14740 GND.n8356 GND.n8355 585
R14741 GND.n8354 GND.n8353 585
R14742 GND.n8352 GND.n8351 585
R14743 GND.n8350 GND.n8349 585
R14744 GND.n8348 GND.n8347 585
R14745 GND.n8346 GND.n8345 585
R14746 GND.n8344 GND.n8343 585
R14747 GND.n8342 GND.n1373 585
R14748 GND.n8341 GND.n8340 585
R14749 GND.n8339 GND.n8338 585
R14750 GND.n8337 GND.n8336 585
R14751 GND.n8335 GND.n8334 585
R14752 GND.n8333 GND.n8332 585
R14753 GND.n8331 GND.n8330 585
R14754 GND.n8329 GND.n8328 585
R14755 GND.n8327 GND.n8326 585
R14756 GND.n8325 GND.n8324 585
R14757 GND.n8323 GND.n8322 585
R14758 GND.n8321 GND.n8320 585
R14759 GND.n8319 GND.n8318 585
R14760 GND.n8317 GND.n8316 585
R14761 GND.n8315 GND.n8314 585
R14762 GND.n8313 GND.n8312 585
R14763 GND.n8311 GND.n8310 585
R14764 GND.n8309 GND.n8308 585
R14765 GND.n8307 GND.n8306 585
R14766 GND.n8305 GND.n8304 585
R14767 GND.n8303 GND.n8302 585
R14768 GND.n8301 GND.n8300 585
R14769 GND.n8299 GND.n8298 585
R14770 GND.n8297 GND.n8296 585
R14771 GND.n8295 GND.n8294 585
R14772 GND.n8293 GND.n8292 585
R14773 GND.n8291 GND.n8290 585
R14774 GND.n8289 GND.n8288 585
R14775 GND.n8287 GND.n8286 585
R14776 GND.n8285 GND.n8284 585
R14777 GND.n8283 GND.n8282 585
R14778 GND.n8281 GND.n8280 585
R14779 GND.n8279 GND.n8278 585
R14780 GND.n8277 GND.n8276 585
R14781 GND.n8275 GND.n8274 585
R14782 GND.n8273 GND.n8272 585
R14783 GND.n8271 GND.n8270 585
R14784 GND.n8269 GND.n8268 585
R14785 GND.n8266 GND.n8265 585
R14786 GND.n8264 GND.n8263 585
R14787 GND.n8262 GND.n8261 585
R14788 GND.n8260 GND.n8259 585
R14789 GND.n8258 GND.n8257 585
R14790 GND.n8256 GND.n8255 585
R14791 GND.n8254 GND.n8253 585
R14792 GND.n8252 GND.n8251 585
R14793 GND.n8250 GND.n8249 585
R14794 GND.n8248 GND.n8247 585
R14795 GND.n8246 GND.n8245 585
R14796 GND.n8244 GND.n8243 585
R14797 GND.n8242 GND.n1434 585
R14798 GND.n1433 GND.n1351 585
R14799 GND.n8362 GND.n1351 585
R14800 GND.n1821 GND.n1675 585
R14801 GND.n1822 GND.n1819 585
R14802 GND.n1823 GND.n1816 585
R14803 GND.n1814 GND.n1813 585
R14804 GND.n1827 GND.n1812 585
R14805 GND.n1828 GND.n1811 585
R14806 GND.n1829 GND.n1810 585
R14807 GND.n1808 GND.n1807 585
R14808 GND.n1833 GND.n1806 585
R14809 GND.n1834 GND.n1805 585
R14810 GND.n1835 GND.n1804 585
R14811 GND.n1802 GND.n1801 585
R14812 GND.n1839 GND.n1800 585
R14813 GND.n1840 GND.n1799 585
R14814 GND.n1842 GND.n1796 585
R14815 GND.n1794 GND.n1793 585
R14816 GND.n1846 GND.n1792 585
R14817 GND.n1847 GND.n1791 585
R14818 GND.n1848 GND.n1790 585
R14819 GND.n1788 GND.n1787 585
R14820 GND.n1852 GND.n1786 585
R14821 GND.n1853 GND.n1785 585
R14822 GND.n1854 GND.n1784 585
R14823 GND.n1782 GND.n1781 585
R14824 GND.n1858 GND.n1780 585
R14825 GND.n1859 GND.n1779 585
R14826 GND.n1860 GND.n1778 585
R14827 GND.n1774 GND.n1773 585
R14828 GND.n1864 GND.n1772 585
R14829 GND.n1865 GND.n1771 585
R14830 GND.n1866 GND.n1770 585
R14831 GND.n1768 GND.n1767 585
R14832 GND.n8023 GND.n1684 585
R14833 GND.n7979 GND.n7978 585
R14834 GND.n7980 GND.n1766 585
R14835 GND.n1764 GND.n1763 585
R14836 GND.n7984 GND.n1762 585
R14837 GND.n7985 GND.n1761 585
R14838 GND.n7987 GND.n1758 585
R14839 GND.n1756 GND.n1755 585
R14840 GND.n7991 GND.n1754 585
R14841 GND.n7992 GND.n1753 585
R14842 GND.n7993 GND.n1752 585
R14843 GND.n1750 GND.n1749 585
R14844 GND.n7997 GND.n1748 585
R14845 GND.n7998 GND.n1747 585
R14846 GND.n7999 GND.n1746 585
R14847 GND.n1744 GND.n1743 585
R14848 GND.n8003 GND.n1742 585
R14849 GND.n8004 GND.n1741 585
R14850 GND.n8005 GND.n1740 585
R14851 GND.n1736 GND.n1735 585
R14852 GND.n8009 GND.n1734 585
R14853 GND.n8010 GND.n1733 585
R14854 GND.n8011 GND.n1732 585
R14855 GND.n1730 GND.n1729 585
R14856 GND.n8015 GND.n1728 585
R14857 GND.n8016 GND.n1727 585
R14858 GND.n8017 GND.n1726 585
R14859 GND.n1723 GND.n1722 585
R14860 GND.n8022 GND.n8021 585
R14861 GND.n8023 GND.n8022 585
R14862 GND.n8028 GND.n8027 585
R14863 GND.n8027 GND.n8026 585
R14864 GND.n1674 GND.n1669 585
R14865 GND.n3843 GND.n1674 585
R14866 GND.n8032 GND.n1668 585
R14867 GND.n3830 GND.n1668 585
R14868 GND.n8033 GND.n1667 585
R14869 GND.n3834 GND.n1667 585
R14870 GND.n8034 GND.n1666 585
R14871 GND.n3828 GND.n1666 585
R14872 GND.n2382 GND.n1661 585
R14873 GND.n2383 GND.n2382 585
R14874 GND.n8038 GND.n1660 585
R14875 GND.n3817 GND.n1660 585
R14876 GND.n8039 GND.n1659 585
R14877 GND.n3804 GND.n1659 585
R14878 GND.n8040 GND.n1658 585
R14879 GND.n3807 GND.n1658 585
R14880 GND.n2394 GND.n1653 585
R14881 GND.n3801 GND.n2394 585
R14882 GND.n8044 GND.n1652 585
R14883 GND.n2405 GND.n1652 585
R14884 GND.n8045 GND.n1651 585
R14885 GND.n3791 GND.n1651 585
R14886 GND.n8046 GND.n1650 585
R14887 GND.n3778 GND.n1650 585
R14888 GND.n2412 GND.n1645 585
R14889 GND.n3781 GND.n2412 585
R14890 GND.n8050 GND.n1644 585
R14891 GND.n3776 GND.n1644 585
R14892 GND.n8051 GND.n1643 585
R14893 GND.n2427 GND.n1643 585
R14894 GND.n8052 GND.n1642 585
R14895 GND.n3766 GND.n1642 585
R14896 GND.n3752 GND.n1637 585
R14897 GND.n3753 GND.n3752 585
R14898 GND.n8056 GND.n1636 585
R14899 GND.n3756 GND.n1636 585
R14900 GND.n8057 GND.n1635 585
R14901 GND.n3750 GND.n1635 585
R14902 GND.n8058 GND.n1634 585
R14903 GND.n3473 GND.n1634 585
R14904 GND.n2445 GND.n1629 585
R14905 GND.n3740 GND.n2445 585
R14906 GND.n8062 GND.n1628 585
R14907 GND.n3726 GND.n1628 585
R14908 GND.n8063 GND.n1627 585
R14909 GND.n3730 GND.n1627 585
R14910 GND.n8064 GND.n1626 585
R14911 GND.n3724 GND.n1626 585
R14912 GND.n2467 GND.n1621 585
R14913 GND.n2468 GND.n2467 585
R14914 GND.n8068 GND.n1620 585
R14915 GND.n3714 GND.n1620 585
R14916 GND.n8069 GND.n1619 585
R14917 GND.n3701 GND.n1619 585
R14918 GND.n8070 GND.n1618 585
R14919 GND.n3704 GND.n1618 585
R14920 GND.n2479 GND.n1613 585
R14921 GND.n3698 GND.n2479 585
R14922 GND.n8074 GND.n1612 585
R14923 GND.n2490 GND.n1612 585
R14924 GND.n8075 GND.n1611 585
R14925 GND.n3688 GND.n1611 585
R14926 GND.n8076 GND.n1610 585
R14927 GND.n3675 GND.n1610 585
R14928 GND.n2497 GND.n1605 585
R14929 GND.n3678 GND.n2497 585
R14930 GND.n8080 GND.n1604 585
R14931 GND.n3673 GND.n1604 585
R14932 GND.n8081 GND.n1603 585
R14933 GND.n2512 GND.n1603 585
R14934 GND.n8082 GND.n1602 585
R14935 GND.n3663 GND.n1602 585
R14936 GND.n3649 GND.n1597 585
R14937 GND.n3650 GND.n3649 585
R14938 GND.n8086 GND.n1596 585
R14939 GND.n3653 GND.n1596 585
R14940 GND.n8087 GND.n1595 585
R14941 GND.n3647 GND.n1595 585
R14942 GND.n8088 GND.n1594 585
R14943 GND.n2534 GND.n1594 585
R14944 GND.n2530 GND.n1589 585
R14945 GND.n3637 GND.n2530 585
R14946 GND.n8092 GND.n1588 585
R14947 GND.n3623 GND.n1588 585
R14948 GND.n8093 GND.n1587 585
R14949 GND.n3627 GND.n1587 585
R14950 GND.n8094 GND.n1586 585
R14951 GND.n3621 GND.n1586 585
R14952 GND.n2554 GND.n1581 585
R14953 GND.n2555 GND.n2554 585
R14954 GND.n8098 GND.n1580 585
R14955 GND.n3611 GND.n1580 585
R14956 GND.n8099 GND.n1579 585
R14957 GND.n3598 GND.n1579 585
R14958 GND.n8100 GND.n1578 585
R14959 GND.n3601 GND.n1578 585
R14960 GND.n2566 GND.n1573 585
R14961 GND.n3595 GND.n2566 585
R14962 GND.n8104 GND.n1572 585
R14963 GND.n2577 GND.n1572 585
R14964 GND.n8105 GND.n1571 585
R14965 GND.n3585 GND.n1571 585
R14966 GND.n8106 GND.n1570 585
R14967 GND.n3572 GND.n1570 585
R14968 GND.n2584 GND.n1565 585
R14969 GND.n3575 GND.n2584 585
R14970 GND.n8110 GND.n1564 585
R14971 GND.n3570 GND.n1564 585
R14972 GND.n8111 GND.n1563 585
R14973 GND.n2588 GND.n1563 585
R14974 GND.n8112 GND.n1553 585
R14975 GND.n8116 GND.n1553 585
R14976 GND.n3558 GND.n1562 585
R14977 GND.n3559 GND.n3558 585
R14978 GND.n3557 GND.n2598 585
R14979 GND.n3557 GND.n3556 585
R14980 GND.n3549 GND.n2597 585
R14981 GND.n2600 GND.n2597 585
R14982 GND.n3548 GND.n1534 585
R14983 GND.n8123 GND.n1534 585
R14984 GND.n3547 GND.n2605 585
R14985 GND.n3542 GND.n2605 585
R14986 GND.n2616 GND.n2604 585
R14987 GND.n2616 GND.n2610 585
R14988 GND.n3314 GND.n2617 585
R14989 GND.n3327 GND.n2617 585
R14990 GND.n3315 GND.n3311 585
R14991 GND.n3311 GND.n2615 585
R14992 GND.n3316 GND.n2623 585
R14993 GND.n3320 GND.n2623 585
R14994 GND.n3310 GND.n3309 585
R14995 GND.n3309 GND.n3308 585
R14996 GND.n2632 GND.n2631 585
R14997 GND.n2633 GND.n2632 585
R14998 GND.n3278 GND.n2641 585
R14999 GND.n3295 GND.n2641 585
R15000 GND.n3279 GND.n3272 585
R15001 GND.n3272 GND.n2640 585
R15002 GND.n3280 GND.n2651 585
R15003 GND.n3284 GND.n2651 585
R15004 GND.n3271 GND.n3270 585
R15005 GND.n3270 GND.n3269 585
R15006 GND.n2661 GND.n2660 585
R15007 GND.n2662 GND.n2661 585
R15008 GND.n3241 GND.n2671 585
R15009 GND.n3257 GND.n2671 585
R15010 GND.n3242 GND.n3235 585
R15011 GND.n3235 GND.n2670 585
R15012 GND.n3243 GND.n2681 585
R15013 GND.n3247 GND.n2681 585
R15014 GND.n3234 GND.n3233 585
R15015 GND.n3233 GND.n3232 585
R15016 GND.n2690 GND.n2689 585
R15017 GND.n2691 GND.n2690 585
R15018 GND.n3204 GND.n2699 585
R15019 GND.n3220 GND.n2699 585
R15020 GND.n3205 GND.n3198 585
R15021 GND.n3198 GND.n2698 585
R15022 GND.n3206 GND.n2710 585
R15023 GND.n3210 GND.n2710 585
R15024 GND.n3197 GND.n3196 585
R15025 GND.n3196 GND.n3195 585
R15026 GND.n2719 GND.n2718 585
R15027 GND.n2721 GND.n2719 585
R15028 GND.n3167 GND.n2729 585
R15029 GND.n3183 GND.n2729 585
R15030 GND.n3168 GND.n3161 585
R15031 GND.n3161 GND.n2728 585
R15032 GND.n3169 GND.n2739 585
R15033 GND.n3173 GND.n2739 585
R15034 GND.n3160 GND.n3159 585
R15035 GND.n3159 GND.n3158 585
R15036 GND.n2748 GND.n2747 585
R15037 GND.n2749 GND.n2748 585
R15038 GND.n3129 GND.n2756 585
R15039 GND.n3145 GND.n2756 585
R15040 GND.n3130 GND.n3123 585
R15041 GND.n3123 GND.n3122 585
R15042 GND.n3131 GND.n2766 585
R15043 GND.n3135 GND.n2766 585
R15044 GND.n3121 GND.n3120 585
R15045 GND.n3120 GND.n3119 585
R15046 GND.n2776 GND.n2775 585
R15047 GND.n2777 GND.n2776 585
R15048 GND.n3091 GND.n2786 585
R15049 GND.n3107 GND.n2786 585
R15050 GND.n3092 GND.n3085 585
R15051 GND.n3085 GND.n2785 585
R15052 GND.n3093 GND.n2796 585
R15053 GND.n3097 GND.n2796 585
R15054 GND.n3084 GND.n3083 585
R15055 GND.n3083 GND.n3082 585
R15056 GND.n2805 GND.n2804 585
R15057 GND.n2806 GND.n2805 585
R15058 GND.n3054 GND.n2814 585
R15059 GND.n3070 GND.n2814 585
R15060 GND.n3055 GND.n3048 585
R15061 GND.n3048 GND.n2813 585
R15062 GND.n3056 GND.n2824 585
R15063 GND.n3060 GND.n2824 585
R15064 GND.n3047 GND.n3046 585
R15065 GND.n3046 GND.n3045 585
R15066 GND.n2833 GND.n2832 585
R15067 GND.n3035 GND.n2833 585
R15068 GND.n3022 GND.n3021 585
R15069 GND.n3021 GND.n2840 585
R15070 GND.n3023 GND.n2849 585
R15071 GND.n3027 GND.n2849 585
R15072 GND.n3020 GND.n3019 585
R15073 GND.n3019 GND.n3018 585
R15074 GND.n2860 GND.n2859 585
R15075 GND.n2862 GND.n2860 585
R15076 GND.n2988 GND.n2864 585
R15077 GND.n3004 GND.n2864 585
R15078 GND.n2989 GND.n2982 585
R15079 GND.n2982 GND.n2875 585
R15080 GND.n2990 GND.n2874 585
R15081 GND.n2994 GND.n2874 585
R15082 GND.n2981 GND.n2980 585
R15083 GND.n2980 GND.n2873 585
R15084 GND.n2979 GND.n2882 585
R15085 GND.n2979 GND.n2978 585
R15086 GND.n2965 GND.n2883 585
R15087 GND.n2884 GND.n2883 585
R15088 GND.n2966 GND.n2893 585
R15089 GND.n2970 GND.n2893 585
R15090 GND.n2964 GND.n2963 585
R15091 GND.n2963 GND.n2892 585
R15092 GND.n2962 GND.n2902 585
R15093 GND.n2962 GND.n2961 585
R15094 GND.n2948 GND.n2903 585
R15095 GND.n2904 GND.n2903 585
R15096 GND.n2949 GND.n2913 585
R15097 GND.n2953 GND.n2913 585
R15098 GND.n2947 GND.n2946 585
R15099 GND.n2946 GND.n2912 585
R15100 GND.n2945 GND.n2922 585
R15101 GND.n2945 GND.n2944 585
R15102 GND.n2931 GND.n2923 585
R15103 GND.n2924 GND.n2923 585
R15104 GND.n2930 GND.n2929 585
R15105 GND.n2929 GND.n1358 585
R15106 GND.n10137 GND.n10136 585
R15107 GND.n10136 GND.n10135 585
R15108 GND.n10138 GND.n409 585
R15109 GND.n409 GND.n408 585
R15110 GND.n10140 GND.n10139 585
R15111 GND.n10141 GND.n10140 585
R15112 GND.n396 GND.n395 585
R15113 GND.n399 GND.n396 585
R15114 GND.n10149 GND.n10148 585
R15115 GND.n10148 GND.n10147 585
R15116 GND.n10150 GND.n390 585
R15117 GND.n390 GND.n389 585
R15118 GND.n10152 GND.n10151 585
R15119 GND.n10153 GND.n10152 585
R15120 GND.n377 GND.n376 585
R15121 GND.n380 GND.n377 585
R15122 GND.n10161 GND.n10160 585
R15123 GND.n10160 GND.n10159 585
R15124 GND.n10162 GND.n371 585
R15125 GND.n371 GND.n370 585
R15126 GND.n10164 GND.n10163 585
R15127 GND.n10165 GND.n10164 585
R15128 GND.n357 GND.n356 585
R15129 GND.n361 GND.n357 585
R15130 GND.n10173 GND.n10172 585
R15131 GND.n10172 GND.n10171 585
R15132 GND.n10174 GND.n351 585
R15133 GND.n358 GND.n351 585
R15134 GND.n10176 GND.n10175 585
R15135 GND.n10177 GND.n10176 585
R15136 GND.n336 GND.n335 585
R15137 GND.n10104 GND.n336 585
R15138 GND.n10185 GND.n10184 585
R15139 GND.n10184 GND.n10183 585
R15140 GND.n10186 GND.n330 585
R15141 GND.n9787 GND.n330 585
R15142 GND.n10188 GND.n10187 585
R15143 GND.n10189 GND.n10188 585
R15144 GND.n315 GND.n314 585
R15145 GND.n9780 GND.n315 585
R15146 GND.n10197 GND.n10196 585
R15147 GND.n10196 GND.n10195 585
R15148 GND.n10198 GND.n309 585
R15149 GND.n9772 GND.n309 585
R15150 GND.n10200 GND.n10199 585
R15151 GND.n10201 GND.n10200 585
R15152 GND.n294 GND.n293 585
R15153 GND.n9765 GND.n294 585
R15154 GND.n10209 GND.n10208 585
R15155 GND.n10208 GND.n10207 585
R15156 GND.n10210 GND.n288 585
R15157 GND.n9757 GND.n288 585
R15158 GND.n10212 GND.n10211 585
R15159 GND.n10213 GND.n10212 585
R15160 GND.n273 GND.n272 585
R15161 GND.n9750 GND.n273 585
R15162 GND.n10221 GND.n10220 585
R15163 GND.n10220 GND.n10219 585
R15164 GND.n10222 GND.n267 585
R15165 GND.n9742 GND.n267 585
R15166 GND.n10224 GND.n10223 585
R15167 GND.n10225 GND.n10224 585
R15168 GND.n253 GND.n252 585
R15169 GND.n9735 GND.n253 585
R15170 GND.n10233 GND.n10232 585
R15171 GND.n10232 GND.n10231 585
R15172 GND.n10234 GND.n247 585
R15173 GND.n9727 GND.n247 585
R15174 GND.n10236 GND.n10235 585
R15175 GND.n10237 GND.n10236 585
R15176 GND.n232 GND.n231 585
R15177 GND.n6835 GND.n232 585
R15178 GND.n10245 GND.n10244 585
R15179 GND.n10244 GND.n10243 585
R15180 GND.n10246 GND.n226 585
R15181 GND.n6841 GND.n226 585
R15182 GND.n10248 GND.n10247 585
R15183 GND.n10249 GND.n10248 585
R15184 GND.n211 GND.n210 585
R15185 GND.n6847 GND.n211 585
R15186 GND.n10257 GND.n10256 585
R15187 GND.n10256 GND.n10255 585
R15188 GND.n10258 GND.n205 585
R15189 GND.n6853 GND.n205 585
R15190 GND.n10260 GND.n10259 585
R15191 GND.n10261 GND.n10260 585
R15192 GND.n190 GND.n189 585
R15193 GND.n6859 GND.n190 585
R15194 GND.n10269 GND.n10268 585
R15195 GND.n10268 GND.n10267 585
R15196 GND.n10270 GND.n184 585
R15197 GND.n6865 GND.n184 585
R15198 GND.n10272 GND.n10271 585
R15199 GND.n10273 GND.n10272 585
R15200 GND.n169 GND.n168 585
R15201 GND.n6871 GND.n169 585
R15202 GND.n10281 GND.n10280 585
R15203 GND.n10280 GND.n10279 585
R15204 GND.n10282 GND.n163 585
R15205 GND.n6877 GND.n163 585
R15206 GND.n10284 GND.n10283 585
R15207 GND.n10285 GND.n10284 585
R15208 GND.n148 GND.n147 585
R15209 GND.n6883 GND.n148 585
R15210 GND.n10293 GND.n10292 585
R15211 GND.n10292 GND.n10291 585
R15212 GND.n10294 GND.n143 585
R15213 GND.n6889 GND.n143 585
R15214 GND.n10296 GND.n10295 585
R15215 GND.n10297 GND.n10296 585
R15216 GND.n126 GND.n124 585
R15217 GND.n6895 GND.n126 585
R15218 GND.n10305 GND.n10304 585
R15219 GND.n10304 GND.n10303 585
R15220 GND.n125 GND.n123 585
R15221 GND.n6901 GND.n125 585
R15222 GND.n5268 GND.n5267 585
R15223 GND.n5269 GND.n5268 585
R15224 GND.n115 GND.n113 585
R15225 GND.n6788 GND.n113 585
R15226 GND.n10309 GND.n10308 585
R15227 GND.n10310 GND.n10309 585
R15228 GND.n114 GND.n112 585
R15229 GND.n6779 GND.n112 585
R15230 GND.n5189 GND.n5188 585
R15231 GND.n5192 GND.n5189 585
R15232 GND.n6917 GND.n121 585
R15233 GND.n6917 GND.n6916 585
R15234 GND.n6919 GND.n6918 585
R15235 GND.n6920 GND.n6919 585
R15236 GND.n5174 GND.n5173 585
R15237 GND.n6769 GND.n5174 585
R15238 GND.n6928 GND.n6927 585
R15239 GND.n6927 GND.n6926 585
R15240 GND.n6929 GND.n5169 585
R15241 GND.n6754 GND.n5169 585
R15242 GND.n6931 GND.n6930 585
R15243 GND.n6932 GND.n6931 585
R15244 GND.n5154 GND.n5153 585
R15245 GND.n6579 GND.n5154 585
R15246 GND.n6940 GND.n6939 585
R15247 GND.n6939 GND.n6938 585
R15248 GND.n6941 GND.n5148 585
R15249 GND.n6585 GND.n5148 585
R15250 GND.n6943 GND.n6942 585
R15251 GND.n6944 GND.n6943 585
R15252 GND.n5133 GND.n5132 585
R15253 GND.n6591 GND.n5133 585
R15254 GND.n6952 GND.n6951 585
R15255 GND.n6951 GND.n6950 585
R15256 GND.n6953 GND.n5127 585
R15257 GND.n6597 GND.n5127 585
R15258 GND.n6955 GND.n6954 585
R15259 GND.n6956 GND.n6955 585
R15260 GND.n5112 GND.n5111 585
R15261 GND.n6603 GND.n5112 585
R15262 GND.n6964 GND.n6963 585
R15263 GND.n6963 GND.n6962 585
R15264 GND.n6965 GND.n5106 585
R15265 GND.n6609 GND.n5106 585
R15266 GND.n6967 GND.n6966 585
R15267 GND.n6968 GND.n6967 585
R15268 GND.n5091 GND.n5090 585
R15269 GND.n6615 GND.n5091 585
R15270 GND.n6976 GND.n6975 585
R15271 GND.n6975 GND.n6974 585
R15272 GND.n6977 GND.n5085 585
R15273 GND.n6621 GND.n5085 585
R15274 GND.n6979 GND.n6978 585
R15275 GND.n6980 GND.n6979 585
R15276 GND.n5070 GND.n5069 585
R15277 GND.n6627 GND.n5070 585
R15278 GND.n6988 GND.n6987 585
R15279 GND.n6987 GND.n6986 585
R15280 GND.n6989 GND.n5064 585
R15281 GND.n6633 GND.n5064 585
R15282 GND.n6991 GND.n6990 585
R15283 GND.n6992 GND.n6991 585
R15284 GND.n5049 GND.n5048 585
R15285 GND.n6639 GND.n5049 585
R15286 GND.n7000 GND.n6999 585
R15287 GND.n6999 GND.n6998 585
R15288 GND.n7001 GND.n5043 585
R15289 GND.n6645 GND.n5043 585
R15290 GND.n7003 GND.n7002 585
R15291 GND.n7004 GND.n7003 585
R15292 GND.n5028 GND.n5027 585
R15293 GND.n6651 GND.n5028 585
R15294 GND.n7012 GND.n7011 585
R15295 GND.n7011 GND.n7010 585
R15296 GND.n7013 GND.n5022 585
R15297 GND.n6657 GND.n5022 585
R15298 GND.n7015 GND.n7014 585
R15299 GND.n7016 GND.n7015 585
R15300 GND.n5007 GND.n5006 585
R15301 GND.n6663 GND.n5007 585
R15302 GND.n7024 GND.n7023 585
R15303 GND.n7023 GND.n7022 585
R15304 GND.n7025 GND.n5001 585
R15305 GND.n6669 GND.n5001 585
R15306 GND.n7027 GND.n7026 585
R15307 GND.n7028 GND.n7027 585
R15308 GND.n4987 GND.n4986 585
R15309 GND.n6675 GND.n4987 585
R15310 GND.n7036 GND.n7035 585
R15311 GND.n7035 GND.n7034 585
R15312 GND.n7037 GND.n4981 585
R15313 GND.n6516 GND.n4981 585
R15314 GND.n7039 GND.n7038 585
R15315 GND.n7040 GND.n7039 585
R15316 GND.n4966 GND.n4965 585
R15317 GND.n6507 GND.n4966 585
R15318 GND.n7048 GND.n7047 585
R15319 GND.n7047 GND.n7046 585
R15320 GND.n7049 GND.n4960 585
R15321 GND.n6501 GND.n4960 585
R15322 GND.n7051 GND.n7050 585
R15323 GND.n7052 GND.n7051 585
R15324 GND.n4945 GND.n4944 585
R15325 GND.n6493 GND.n4945 585
R15326 GND.n7060 GND.n7059 585
R15327 GND.n7059 GND.n7058 585
R15328 GND.n7061 GND.n4939 585
R15329 GND.n6487 GND.n4939 585
R15330 GND.n7063 GND.n7062 585
R15331 GND.n7064 GND.n7063 585
R15332 GND.n4923 GND.n4922 585
R15333 GND.n6479 GND.n4923 585
R15334 GND.n7072 GND.n7071 585
R15335 GND.n7071 GND.n7070 585
R15336 GND.n7073 GND.n4912 585
R15337 GND.n6473 GND.n4912 585
R15338 GND.n7075 GND.n7074 585
R15339 GND.n7076 GND.n7075 585
R15340 GND.n4913 GND.n4911 585
R15341 GND.n4911 GND.n4906 585
R15342 GND.n4916 GND.n4915 585
R15343 GND.n4915 GND.n4896 585
R15344 GND.n4881 GND.n4880 585
R15345 GND.n7084 GND.n4881 585
R15346 GND.n7093 GND.n7092 585
R15347 GND.n7092 GND.n7091 585
R15348 GND.n7094 GND.n4878 585
R15349 GND.n6416 GND.n4878 585
R15350 GND.n7181 GND.n7180 585
R15351 GND.n7179 GND.n4877 585
R15352 GND.n7178 GND.n4876 585
R15353 GND.n7183 GND.n4876 585
R15354 GND.n7177 GND.n7176 585
R15355 GND.n7175 GND.n7174 585
R15356 GND.n7173 GND.n7172 585
R15357 GND.n7171 GND.n7170 585
R15358 GND.n7169 GND.n7168 585
R15359 GND.n7167 GND.n7166 585
R15360 GND.n7165 GND.n7164 585
R15361 GND.n7163 GND.n7106 585
R15362 GND.n7162 GND.n7161 585
R15363 GND.n7160 GND.n7159 585
R15364 GND.n7158 GND.n7157 585
R15365 GND.n7156 GND.n7155 585
R15366 GND.n7154 GND.n7153 585
R15367 GND.n7152 GND.n7151 585
R15368 GND.n7150 GND.n7149 585
R15369 GND.n7148 GND.n7147 585
R15370 GND.n7146 GND.n7145 585
R15371 GND.n7144 GND.n7143 585
R15372 GND.n7142 GND.n7141 585
R15373 GND.n7140 GND.n7139 585
R15374 GND.n7138 GND.n7137 585
R15375 GND.n7136 GND.n7135 585
R15376 GND.n7134 GND.n7133 585
R15377 GND.n7132 GND.n7131 585
R15378 GND.n7130 GND.n4833 585
R15379 GND.n7186 GND.n7185 585
R15380 GND.n4838 GND.n4837 585
R15381 GND.n5385 GND.n5384 585
R15382 GND.n5387 GND.n5386 585
R15383 GND.n5380 GND.n5379 585
R15384 GND.n5393 GND.n5381 585
R15385 GND.n5395 GND.n5394 585
R15386 GND.n5397 GND.n5396 585
R15387 GND.n5401 GND.n5377 585
R15388 GND.n5403 GND.n5402 585
R15389 GND.n5405 GND.n5404 585
R15390 GND.n5407 GND.n5406 585
R15391 GND.n5411 GND.n5375 585
R15392 GND.n5413 GND.n5412 585
R15393 GND.n5415 GND.n5414 585
R15394 GND.n5417 GND.n5416 585
R15395 GND.n5421 GND.n5373 585
R15396 GND.n5423 GND.n5422 585
R15397 GND.n5428 GND.n5427 585
R15398 GND.n5430 GND.n5429 585
R15399 GND.n5434 GND.n5371 585
R15400 GND.n5436 GND.n5435 585
R15401 GND.n5438 GND.n5437 585
R15402 GND.n5440 GND.n5439 585
R15403 GND.n5444 GND.n5369 585
R15404 GND.n5446 GND.n5445 585
R15405 GND.n5448 GND.n5447 585
R15406 GND.n5450 GND.n5449 585
R15407 GND.n5454 GND.n5367 585
R15408 GND.n5456 GND.n5455 585
R15409 GND.n5460 GND.n5457 585
R15410 GND.n5461 GND.n4868 585
R15411 GND.n7183 GND.n4868 585
R15412 GND.n10038 GND.n10037 585
R15413 GND.n9845 GND.n9842 585
R15414 GND.n10033 GND.n10032 585
R15415 GND.n10031 GND.n10030 585
R15416 GND.n10029 GND.n10028 585
R15417 GND.n10022 GND.n9847 585
R15418 GND.n10024 GND.n10023 585
R15419 GND.n10021 GND.n10020 585
R15420 GND.n10019 GND.n10018 585
R15421 GND.n10012 GND.n9849 585
R15422 GND.n10014 GND.n10013 585
R15423 GND.n10011 GND.n10010 585
R15424 GND.n10009 GND.n10008 585
R15425 GND.n10002 GND.n9851 585
R15426 GND.n10004 GND.n10003 585
R15427 GND.n9998 GND.n9997 585
R15428 GND.n9996 GND.n9995 585
R15429 GND.n9989 GND.n9853 585
R15430 GND.n9991 GND.n9990 585
R15431 GND.n9988 GND.n9987 585
R15432 GND.n9986 GND.n9985 585
R15433 GND.n9979 GND.n9855 585
R15434 GND.n9981 GND.n9980 585
R15435 GND.n9978 GND.n9977 585
R15436 GND.n9976 GND.n9975 585
R15437 GND.n9861 GND.n9857 585
R15438 GND.n9971 GND.n9862 585
R15439 GND.n9970 GND.n9969 585
R15440 GND.n9968 GND.n9967 585
R15441 GND.n9961 GND.n9863 585
R15442 GND.n9963 GND.n9962 585
R15443 GND.n9960 GND.n9959 585
R15444 GND.n9958 GND.n9957 585
R15445 GND.n9951 GND.n9865 585
R15446 GND.n9953 GND.n9952 585
R15447 GND.n9950 GND.n9949 585
R15448 GND.n9948 GND.n9947 585
R15449 GND.n9941 GND.n9867 585
R15450 GND.n9943 GND.n9942 585
R15451 GND.n9939 GND.n9938 585
R15452 GND.n9937 GND.n9936 585
R15453 GND.n9930 GND.n9871 585
R15454 GND.n9932 GND.n9931 585
R15455 GND.n9929 GND.n9928 585
R15456 GND.n9927 GND.n9926 585
R15457 GND.n9920 GND.n9873 585
R15458 GND.n9922 GND.n9921 585
R15459 GND.n9919 GND.n9918 585
R15460 GND.n9917 GND.n9916 585
R15461 GND.n9910 GND.n9875 585
R15462 GND.n9912 GND.n9911 585
R15463 GND.n9909 GND.n9879 585
R15464 GND.n9908 GND.n9907 585
R15465 GND.n9901 GND.n9880 585
R15466 GND.n9903 GND.n9902 585
R15467 GND.n9900 GND.n9899 585
R15468 GND.n9898 GND.n9897 585
R15469 GND.n9891 GND.n9882 585
R15470 GND.n9893 GND.n9892 585
R15471 GND.n9890 GND.n9889 585
R15472 GND.n9888 GND.n9887 585
R15473 GND.n9884 GND.n414 585
R15474 GND.n10131 GND.n415 585
R15475 GND.n10135 GND.n415 585
R15476 GND.n10130 GND.n10129 585
R15477 GND.n10129 GND.n408 585
R15478 GND.n10128 GND.n406 585
R15479 GND.n10141 GND.n406 585
R15480 GND.n10127 GND.n10126 585
R15481 GND.n10126 GND.n399 585
R15482 GND.n10125 GND.n397 585
R15483 GND.n10147 GND.n397 585
R15484 GND.n10124 GND.n10123 585
R15485 GND.n10123 GND.n389 585
R15486 GND.n10121 GND.n387 585
R15487 GND.n10153 GND.n387 585
R15488 GND.n10120 GND.n10119 585
R15489 GND.n10119 GND.n380 585
R15490 GND.n10118 GND.n378 585
R15491 GND.n10159 GND.n378 585
R15492 GND.n10117 GND.n10116 585
R15493 GND.n10116 GND.n370 585
R15494 GND.n10114 GND.n368 585
R15495 GND.n10165 GND.n368 585
R15496 GND.n10113 GND.n10112 585
R15497 GND.n10112 GND.n361 585
R15498 GND.n10111 GND.n359 585
R15499 GND.n10171 GND.n359 585
R15500 GND.n10110 GND.n10109 585
R15501 GND.n10109 GND.n358 585
R15502 GND.n10107 GND.n348 585
R15503 GND.n10177 GND.n348 585
R15504 GND.n10106 GND.n10105 585
R15505 GND.n10105 GND.n10104 585
R15506 GND.n421 GND.n338 585
R15507 GND.n10183 GND.n338 585
R15508 GND.n9786 GND.n9785 585
R15509 GND.n9787 GND.n9786 585
R15510 GND.n9783 GND.n327 585
R15511 GND.n10189 GND.n327 585
R15512 GND.n9782 GND.n9781 585
R15513 GND.n9781 GND.n9780 585
R15514 GND.n425 GND.n317 585
R15515 GND.n10195 GND.n317 585
R15516 GND.n9771 GND.n9770 585
R15517 GND.n9772 GND.n9771 585
R15518 GND.n9768 GND.n306 585
R15519 GND.n10201 GND.n306 585
R15520 GND.n9767 GND.n9766 585
R15521 GND.n9766 GND.n9765 585
R15522 GND.n429 GND.n296 585
R15523 GND.n10207 GND.n296 585
R15524 GND.n9756 GND.n9755 585
R15525 GND.n9757 GND.n9756 585
R15526 GND.n9753 GND.n285 585
R15527 GND.n10213 GND.n285 585
R15528 GND.n9752 GND.n9751 585
R15529 GND.n9751 GND.n9750 585
R15530 GND.n433 GND.n275 585
R15531 GND.n10219 GND.n275 585
R15532 GND.n9741 GND.n9740 585
R15533 GND.n9742 GND.n9741 585
R15534 GND.n9738 GND.n264 585
R15535 GND.n10225 GND.n264 585
R15536 GND.n9737 GND.n9736 585
R15537 GND.n9736 GND.n9735 585
R15538 GND.n437 GND.n254 585
R15539 GND.n10231 GND.n254 585
R15540 GND.n6831 GND.n441 585
R15541 GND.n9727 GND.n441 585
R15542 GND.n6832 GND.n244 585
R15543 GND.n10237 GND.n244 585
R15544 GND.n6834 GND.n6833 585
R15545 GND.n6835 GND.n6834 585
R15546 GND.n6825 GND.n234 585
R15547 GND.n10243 GND.n234 585
R15548 GND.n6843 GND.n6842 585
R15549 GND.n6842 GND.n6841 585
R15550 GND.n6844 GND.n223 585
R15551 GND.n10249 GND.n223 585
R15552 GND.n6846 GND.n6845 585
R15553 GND.n6847 GND.n6846 585
R15554 GND.n6818 GND.n213 585
R15555 GND.n10255 GND.n213 585
R15556 GND.n6855 GND.n6854 585
R15557 GND.n6854 GND.n6853 585
R15558 GND.n6856 GND.n202 585
R15559 GND.n10261 GND.n202 585
R15560 GND.n6858 GND.n6857 585
R15561 GND.n6859 GND.n6858 585
R15562 GND.n6811 GND.n192 585
R15563 GND.n10267 GND.n192 585
R15564 GND.n6867 GND.n6866 585
R15565 GND.n6866 GND.n6865 585
R15566 GND.n6868 GND.n181 585
R15567 GND.n10273 GND.n181 585
R15568 GND.n6870 GND.n6869 585
R15569 GND.n6871 GND.n6870 585
R15570 GND.n6804 GND.n171 585
R15571 GND.n10279 GND.n171 585
R15572 GND.n6879 GND.n6878 585
R15573 GND.n6878 GND.n6877 585
R15574 GND.n6880 GND.n160 585
R15575 GND.n10285 GND.n160 585
R15576 GND.n6882 GND.n6881 585
R15577 GND.n6883 GND.n6882 585
R15578 GND.n6797 GND.n150 585
R15579 GND.n10291 GND.n150 585
R15580 GND.n6891 GND.n6890 585
R15581 GND.n6890 GND.n6889 585
R15582 GND.n6892 GND.n140 585
R15583 GND.n10297 GND.n140 585
R15584 GND.n6894 GND.n6893 585
R15585 GND.n6895 GND.n6894 585
R15586 GND.n6795 GND.n128 585
R15587 GND.n10303 GND.n128 585
R15588 GND.n6794 GND.n5270 585
R15589 GND.n6901 GND.n5270 585
R15590 GND.n5281 GND.n5278 585
R15591 GND.n5281 GND.n5269 585
R15592 GND.n6786 GND.n6785 585
R15593 GND.n6788 GND.n6786 585
R15594 GND.n6784 GND.n109 585
R15595 GND.n10310 GND.n109 585
R15596 GND.n6778 GND.n5282 585
R15597 GND.n6779 GND.n6778 585
R15598 GND.n6777 GND.n6776 585
R15599 GND.n6777 GND.n5192 585
R15600 GND.n6773 GND.n5190 585
R15601 GND.n6916 GND.n5190 585
R15602 GND.n6772 GND.n5185 585
R15603 GND.n6920 GND.n5185 585
R15604 GND.n6771 GND.n6770 585
R15605 GND.n6770 GND.n6769 585
R15606 GND.n5287 GND.n5175 585
R15607 GND.n6926 GND.n5175 585
R15608 GND.n6573 GND.n5291 585
R15609 GND.n6754 GND.n5291 585
R15610 GND.n6574 GND.n5166 585
R15611 GND.n6932 GND.n5166 585
R15612 GND.n6581 GND.n6580 585
R15613 GND.n6580 GND.n6579 585
R15614 GND.n6582 GND.n5156 585
R15615 GND.n6938 GND.n5156 585
R15616 GND.n6584 GND.n6583 585
R15617 GND.n6585 GND.n6584 585
R15618 GND.n6565 GND.n5145 585
R15619 GND.n6944 GND.n5145 585
R15620 GND.n6593 GND.n6592 585
R15621 GND.n6592 GND.n6591 585
R15622 GND.n6594 GND.n5135 585
R15623 GND.n6950 GND.n5135 585
R15624 GND.n6596 GND.n6595 585
R15625 GND.n6597 GND.n6596 585
R15626 GND.n6558 GND.n5124 585
R15627 GND.n6956 GND.n5124 585
R15628 GND.n6605 GND.n6604 585
R15629 GND.n6604 GND.n6603 585
R15630 GND.n6606 GND.n5114 585
R15631 GND.n6962 GND.n5114 585
R15632 GND.n6608 GND.n6607 585
R15633 GND.n6609 GND.n6608 585
R15634 GND.n6551 GND.n5103 585
R15635 GND.n6968 GND.n5103 585
R15636 GND.n6617 GND.n6616 585
R15637 GND.n6616 GND.n6615 585
R15638 GND.n6618 GND.n5093 585
R15639 GND.n6974 GND.n5093 585
R15640 GND.n6620 GND.n6619 585
R15641 GND.n6621 GND.n6620 585
R15642 GND.n6544 GND.n5082 585
R15643 GND.n6980 GND.n5082 585
R15644 GND.n6629 GND.n6628 585
R15645 GND.n6628 GND.n6627 585
R15646 GND.n6630 GND.n5072 585
R15647 GND.n6986 GND.n5072 585
R15648 GND.n6632 GND.n6631 585
R15649 GND.n6633 GND.n6632 585
R15650 GND.n6537 GND.n5061 585
R15651 GND.n6992 GND.n5061 585
R15652 GND.n6641 GND.n6640 585
R15653 GND.n6640 GND.n6639 585
R15654 GND.n6642 GND.n5051 585
R15655 GND.n6998 GND.n5051 585
R15656 GND.n6644 GND.n6643 585
R15657 GND.n6645 GND.n6644 585
R15658 GND.n6530 GND.n5040 585
R15659 GND.n7004 GND.n5040 585
R15660 GND.n6653 GND.n6652 585
R15661 GND.n6652 GND.n6651 585
R15662 GND.n6654 GND.n5030 585
R15663 GND.n7010 GND.n5030 585
R15664 GND.n6656 GND.n6655 585
R15665 GND.n6657 GND.n6656 585
R15666 GND.n6523 GND.n5019 585
R15667 GND.n7016 GND.n5019 585
R15668 GND.n6665 GND.n6664 585
R15669 GND.n6664 GND.n6663 585
R15670 GND.n6666 GND.n5009 585
R15671 GND.n7022 GND.n5009 585
R15672 GND.n6668 GND.n6667 585
R15673 GND.n6669 GND.n6668 585
R15674 GND.n6521 GND.n4998 585
R15675 GND.n7028 GND.n4998 585
R15676 GND.n6520 GND.n5330 585
R15677 GND.n6675 GND.n5330 585
R15678 GND.n6519 GND.n4989 585
R15679 GND.n7034 GND.n4989 585
R15680 GND.n6518 GND.n6517 585
R15681 GND.n6517 GND.n6516 585
R15682 GND.n5336 GND.n4978 585
R15683 GND.n7040 GND.n4978 585
R15684 GND.n6506 GND.n6505 585
R15685 GND.n6507 GND.n6506 585
R15686 GND.n6504 GND.n4968 585
R15687 GND.n7046 GND.n4968 585
R15688 GND.n6503 GND.n6502 585
R15689 GND.n6502 GND.n6501 585
R15690 GND.n5341 GND.n4957 585
R15691 GND.n7052 GND.n4957 585
R15692 GND.n6492 GND.n6491 585
R15693 GND.n6493 GND.n6492 585
R15694 GND.n6490 GND.n4947 585
R15695 GND.n7058 GND.n4947 585
R15696 GND.n6489 GND.n6488 585
R15697 GND.n6488 GND.n6487 585
R15698 GND.n5346 GND.n4936 585
R15699 GND.n7064 GND.n4936 585
R15700 GND.n6478 GND.n6477 585
R15701 GND.n6479 GND.n6478 585
R15702 GND.n6476 GND.n4924 585
R15703 GND.n7070 GND.n4924 585
R15704 GND.n6475 GND.n6474 585
R15705 GND.n6474 GND.n6473 585
R15706 GND.n5351 GND.n4907 585
R15707 GND.n7076 GND.n4907 585
R15708 GND.n5353 GND.n5352 585
R15709 GND.n5352 GND.n4906 585
R15710 GND.n4894 GND.n4893 585
R15711 GND.n4896 GND.n4894 585
R15712 GND.n7086 GND.n7085 585
R15713 GND.n7085 GND.n7084 585
R15714 GND.n7087 GND.n4883 585
R15715 GND.n7091 GND.n4883 585
R15716 GND.n6415 GND.n4892 585
R15717 GND.n6416 GND.n6415 585
R15718 GND.n9696 GND.n472 585
R15719 GND.n9696 GND.n350 585
R15720 GND.n9698 GND.n9697 585
R15721 GND.n9697 GND.n347 585
R15722 GND.n9699 GND.n467 585
R15723 GND.n467 GND.n340 585
R15724 GND.n9701 GND.n9700 585
R15725 GND.n9701 GND.n337 585
R15726 GND.n9702 GND.n466 585
R15727 GND.n9702 GND.n329 585
R15728 GND.n9704 GND.n9703 585
R15729 GND.n9703 GND.n326 585
R15730 GND.n9705 GND.n461 585
R15731 GND.n461 GND.n319 585
R15732 GND.n9707 GND.n9706 585
R15733 GND.n9707 GND.n316 585
R15734 GND.n9708 GND.n460 585
R15735 GND.n9708 GND.n308 585
R15736 GND.n9710 GND.n9709 585
R15737 GND.n9709 GND.n305 585
R15738 GND.n9711 GND.n455 585
R15739 GND.n455 GND.n298 585
R15740 GND.n9713 GND.n9712 585
R15741 GND.n9713 GND.n295 585
R15742 GND.n9714 GND.n454 585
R15743 GND.n9714 GND.n287 585
R15744 GND.n9716 GND.n9715 585
R15745 GND.n9715 GND.n284 585
R15746 GND.n9717 GND.n449 585
R15747 GND.n449 GND.n277 585
R15748 GND.n9719 GND.n9718 585
R15749 GND.n9719 GND.n274 585
R15750 GND.n9720 GND.n448 585
R15751 GND.n9720 GND.n266 585
R15752 GND.n9722 GND.n9721 585
R15753 GND.n9721 GND.n263 585
R15754 GND.n9723 GND.n443 585
R15755 GND.n443 GND.n256 585
R15756 GND.n9725 GND.n9724 585
R15757 GND.n9726 GND.n9725 585
R15758 GND.n444 GND.n442 585
R15759 GND.n442 GND.n246 585
R15760 GND.n5233 GND.n5228 585
R15761 GND.n5228 GND.n243 585
R15762 GND.n5235 GND.n5234 585
R15763 GND.n5235 GND.n236 585
R15764 GND.n5236 GND.n5227 585
R15765 GND.n5236 GND.n233 585
R15766 GND.n5238 GND.n5237 585
R15767 GND.n5237 GND.n225 585
R15768 GND.n5239 GND.n5222 585
R15769 GND.n5222 GND.n222 585
R15770 GND.n5241 GND.n5240 585
R15771 GND.n5241 GND.n215 585
R15772 GND.n5242 GND.n5221 585
R15773 GND.n5242 GND.n212 585
R15774 GND.n5244 GND.n5243 585
R15775 GND.n5243 GND.n204 585
R15776 GND.n5245 GND.n5216 585
R15777 GND.n5216 GND.n201 585
R15778 GND.n5247 GND.n5246 585
R15779 GND.n5247 GND.n194 585
R15780 GND.n5248 GND.n5215 585
R15781 GND.n5248 GND.n191 585
R15782 GND.n5250 GND.n5249 585
R15783 GND.n5249 GND.n183 585
R15784 GND.n5251 GND.n5210 585
R15785 GND.n5210 GND.n180 585
R15786 GND.n5253 GND.n5252 585
R15787 GND.n5253 GND.n173 585
R15788 GND.n5254 GND.n5209 585
R15789 GND.n5254 GND.n170 585
R15790 GND.n5256 GND.n5255 585
R15791 GND.n5255 GND.n162 585
R15792 GND.n5257 GND.n5204 585
R15793 GND.n5204 GND.n159 585
R15794 GND.n5259 GND.n5258 585
R15795 GND.n5259 GND.n152 585
R15796 GND.n5260 GND.n5203 585
R15797 GND.n5260 GND.n149 585
R15798 GND.n5262 GND.n5261 585
R15799 GND.n5261 GND.n142 585
R15800 GND.n5263 GND.n5199 585
R15801 GND.n5199 GND.n139 585
R15802 GND.n5265 GND.n5264 585
R15803 GND.n5265 GND.n130 585
R15804 GND.n5266 GND.n5198 585
R15805 GND.n5266 GND.n127 585
R15806 GND.n6904 GND.n6903 585
R15807 GND.n6903 GND.n6902 585
R15808 GND.n6906 GND.n5197 585
R15809 GND.n6787 GND.n5197 585
R15810 GND.n6908 GND.n6907 585
R15811 GND.n6908 GND.n110 585
R15812 GND.n6910 GND.n6909 585
R15813 GND.n6909 GND.n108 585
R15814 GND.n6911 GND.n5194 585
R15815 GND.n5286 GND.n5194 585
R15816 GND.n6914 GND.n6913 585
R15817 GND.n6915 GND.n6914 585
R15818 GND.n5195 GND.n5193 585
R15819 GND.n5193 GND.n5187 585
R15820 GND.n6749 GND.n6748 585
R15821 GND.n6748 GND.n5184 585
R15822 GND.n6750 GND.n5293 585
R15823 GND.n5293 GND.n5177 585
R15824 GND.n6752 GND.n6751 585
R15825 GND.n6753 GND.n6752 585
R15826 GND.n5294 GND.n5292 585
R15827 GND.n5292 GND.n5168 585
R15828 GND.n6742 GND.n6741 585
R15829 GND.n6741 GND.n5165 585
R15830 GND.n6740 GND.n5296 585
R15831 GND.n6740 GND.n5158 585
R15832 GND.n6739 GND.n6738 585
R15833 GND.n6739 GND.n5155 585
R15834 GND.n5298 GND.n5297 585
R15835 GND.n5297 GND.n5147 585
R15836 GND.n6734 GND.n6733 585
R15837 GND.n6733 GND.n5144 585
R15838 GND.n6732 GND.n5300 585
R15839 GND.n6732 GND.n5137 585
R15840 GND.n6731 GND.n6730 585
R15841 GND.n6731 GND.n5134 585
R15842 GND.n5302 GND.n5301 585
R15843 GND.n5301 GND.n5126 585
R15844 GND.n6726 GND.n6725 585
R15845 GND.n6725 GND.n5123 585
R15846 GND.n6724 GND.n5304 585
R15847 GND.n6724 GND.n5116 585
R15848 GND.n6723 GND.n6722 585
R15849 GND.n6723 GND.n5113 585
R15850 GND.n5306 GND.n5305 585
R15851 GND.n5305 GND.n5105 585
R15852 GND.n6718 GND.n6717 585
R15853 GND.n6717 GND.n5102 585
R15854 GND.n6716 GND.n5308 585
R15855 GND.n6716 GND.n5095 585
R15856 GND.n6715 GND.n6714 585
R15857 GND.n6715 GND.n5092 585
R15858 GND.n5310 GND.n5309 585
R15859 GND.n5309 GND.n5084 585
R15860 GND.n6710 GND.n6709 585
R15861 GND.n6709 GND.n5081 585
R15862 GND.n6708 GND.n5312 585
R15863 GND.n6708 GND.n5074 585
R15864 GND.n6707 GND.n6706 585
R15865 GND.n6707 GND.n5071 585
R15866 GND.n5314 GND.n5313 585
R15867 GND.n5313 GND.n5063 585
R15868 GND.n6702 GND.n6701 585
R15869 GND.n6701 GND.n5060 585
R15870 GND.n6700 GND.n5316 585
R15871 GND.n6700 GND.n5053 585
R15872 GND.n6699 GND.n6698 585
R15873 GND.n6699 GND.n5050 585
R15874 GND.n5318 GND.n5317 585
R15875 GND.n5317 GND.n5042 585
R15876 GND.n6694 GND.n6693 585
R15877 GND.n6693 GND.n5039 585
R15878 GND.n6692 GND.n5320 585
R15879 GND.n6692 GND.n5032 585
R15880 GND.n6691 GND.n6690 585
R15881 GND.n6691 GND.n5029 585
R15882 GND.n5322 GND.n5321 585
R15883 GND.n5321 GND.n5021 585
R15884 GND.n6686 GND.n6685 585
R15885 GND.n6685 GND.n5018 585
R15886 GND.n6684 GND.n5324 585
R15887 GND.n6684 GND.n5011 585
R15888 GND.n6683 GND.n6682 585
R15889 GND.n6683 GND.n5008 585
R15890 GND.n5326 GND.n5325 585
R15891 GND.n5325 GND.n5000 585
R15892 GND.n6678 GND.n6677 585
R15893 GND.n6677 GND.n6676 585
R15894 GND.n5329 GND.n5328 585
R15895 GND.n5329 GND.n4991 585
R15896 GND.n6453 GND.n6452 585
R15897 GND.n6453 GND.n4988 585
R15898 GND.n6454 GND.n6449 585
R15899 GND.n6454 GND.n4980 585
R15900 GND.n6456 GND.n6455 585
R15901 GND.n6455 GND.n4977 585
R15902 GND.n6457 GND.n6444 585
R15903 GND.n6444 GND.n4970 585
R15904 GND.n6459 GND.n6458 585
R15905 GND.n6459 GND.n4967 585
R15906 GND.n6460 GND.n6443 585
R15907 GND.n6460 GND.n4959 585
R15908 GND.n6462 GND.n6461 585
R15909 GND.n6461 GND.n4956 585
R15910 GND.n6463 GND.n6438 585
R15911 GND.n6438 GND.n4949 585
R15912 GND.n6465 GND.n6464 585
R15913 GND.n6465 GND.n4946 585
R15914 GND.n6466 GND.n6437 585
R15915 GND.n6466 GND.n4938 585
R15916 GND.n6468 GND.n6467 585
R15917 GND.n6467 GND.n4935 585
R15918 GND.n6469 GND.n6432 585
R15919 GND.n6432 GND.n4926 585
R15920 GND.n6471 GND.n6470 585
R15921 GND.n6472 GND.n6471 585
R15922 GND.n4904 GND.n4903 585
R15923 GND.n4909 GND.n4904 585
R15924 GND.n7079 GND.n7078 585
R15925 GND.n7078 GND.n7077 585
R15926 GND.n7080 GND.n4898 585
R15927 GND.n4905 GND.n4898 585
R15928 GND.n7082 GND.n7081 585
R15929 GND.n7083 GND.n7082 585
R15930 GND.n4899 GND.n4897 585
R15931 GND.n4897 GND.n4885 585
R15932 GND.n6411 GND.n6389 585
R15933 GND.n6389 GND.n4882 585
R15934 GND.n6413 GND.n6412 585
R15935 GND.n6414 GND.n6413 585
R15936 GND.n6390 GND.n6388 585
R15937 GND.n6388 GND.n4869 585
R15938 GND.n6405 GND.n6404 585
R15939 GND.n6404 GND.n4839 585
R15940 GND.n6403 GND.n6392 585
R15941 GND.n6403 GND.n6402 585
R15942 GND.n6397 GND.n6393 585
R15943 GND.n6401 GND.n6393 585
R15944 GND.n6399 GND.n6398 585
R15945 GND.n6400 GND.n6399 585
R15946 GND.n4699 GND.n4698 585
R15947 GND.n7250 GND.n4699 585
R15948 GND.n7253 GND.n7252 585
R15949 GND.n7252 GND.n7251 585
R15950 GND.n7254 GND.n4691 585
R15951 GND.n4768 GND.n4691 585
R15952 GND.n7256 GND.n7255 585
R15953 GND.n7257 GND.n7256 585
R15954 GND.n4692 GND.n4690 585
R15955 GND.n4690 GND.n4676 585
R15956 GND.n4621 GND.n4620 585
R15957 GND.n4675 GND.n4621 585
R15958 GND.n7272 GND.n7271 585
R15959 GND.n7271 GND.n7270 585
R15960 GND.n7273 GND.n4615 585
R15961 GND.n4679 GND.n4615 585
R15962 GND.n7275 GND.n7274 585
R15963 GND.n7276 GND.n7275 585
R15964 GND.n4604 GND.n4603 585
R15965 GND.n4607 GND.n4604 585
R15966 GND.n7286 GND.n7285 585
R15967 GND.n7285 GND.n7284 585
R15968 GND.n7287 GND.n4598 585
R15969 GND.n4658 GND.n4598 585
R15970 GND.n7289 GND.n7288 585
R15971 GND.n7290 GND.n7289 585
R15972 GND.n4586 GND.n4585 585
R15973 GND.n4589 GND.n4586 585
R15974 GND.n7300 GND.n7299 585
R15975 GND.n7299 GND.n7298 585
R15976 GND.n7301 GND.n4580 585
R15977 GND.n4645 GND.n4580 585
R15978 GND.n7303 GND.n7302 585
R15979 GND.n7304 GND.n7303 585
R15980 GND.n4568 GND.n4567 585
R15981 GND.n4571 GND.n4568 585
R15982 GND.n7314 GND.n7313 585
R15983 GND.n7313 GND.n7312 585
R15984 GND.n7315 GND.n4560 585
R15985 GND.n4632 GND.n4560 585
R15986 GND.n7317 GND.n7316 585
R15987 GND.n7318 GND.n7317 585
R15988 GND.n4561 GND.n4559 585
R15989 GND.n4559 GND.n4547 585
R15990 GND.n4536 GND.n4535 585
R15991 GND.n4546 GND.n4536 585
R15992 GND.n7333 GND.n7332 585
R15993 GND.n7332 GND.n7331 585
R15994 GND.n7334 GND.n4530 585
R15995 GND.n4537 GND.n4530 585
R15996 GND.n7336 GND.n7335 585
R15997 GND.n7337 GND.n7336 585
R15998 GND.n4518 GND.n4517 585
R15999 GND.n4521 GND.n4518 585
R16000 GND.n7347 GND.n7346 585
R16001 GND.n7346 GND.n7345 585
R16002 GND.n7348 GND.n4512 585
R16003 GND.n6250 GND.n4512 585
R16004 GND.n7350 GND.n7349 585
R16005 GND.n7351 GND.n7350 585
R16006 GND.n4500 GND.n4499 585
R16007 GND.n4503 GND.n4500 585
R16008 GND.n7361 GND.n7360 585
R16009 GND.n7360 GND.n7359 585
R16010 GND.n7362 GND.n4494 585
R16011 GND.n6263 GND.n4494 585
R16012 GND.n7364 GND.n7363 585
R16013 GND.n7365 GND.n7364 585
R16014 GND.n4482 GND.n4481 585
R16015 GND.n4485 GND.n4482 585
R16016 GND.n7375 GND.n7374 585
R16017 GND.n7374 GND.n7373 585
R16018 GND.n7376 GND.n4476 585
R16019 GND.n6276 GND.n4476 585
R16020 GND.n7378 GND.n7377 585
R16021 GND.n7379 GND.n7378 585
R16022 GND.n4464 GND.n4463 585
R16023 GND.n4467 GND.n4464 585
R16024 GND.n7389 GND.n7388 585
R16025 GND.n7388 GND.n7387 585
R16026 GND.n7390 GND.n4458 585
R16027 GND.n6291 GND.n4458 585
R16028 GND.n7392 GND.n7391 585
R16029 GND.n7393 GND.n7392 585
R16030 GND.n4446 GND.n4445 585
R16031 GND.n4455 GND.n4446 585
R16032 GND.n7403 GND.n7402 585
R16033 GND.n7402 GND.n7401 585
R16034 GND.n7404 GND.n4438 585
R16035 GND.n6302 GND.n4438 585
R16036 GND.n7406 GND.n7405 585
R16037 GND.n7407 GND.n7406 585
R16038 GND.n4439 GND.n4437 585
R16039 GND.n5498 GND.n4437 585
R16040 GND.n4413 GND.n4412 585
R16041 GND.n6312 GND.n4413 585
R16042 GND.n7419 GND.n7418 585
R16043 GND.n7418 GND.n7417 585
R16044 GND.n7420 GND.n4407 585
R16045 GND.n6194 GND.n4407 585
R16046 GND.n7422 GND.n7421 585
R16047 GND.n7423 GND.n7422 585
R16048 GND.n4380 GND.n4379 585
R16049 GND.t152 GND.n4380 585
R16050 GND.n7431 GND.n7430 585
R16051 GND.n7430 GND.n7429 585
R16052 GND.n7432 GND.n4372 585
R16053 GND.n6203 GND.n4372 585
R16054 GND.n7434 GND.n7433 585
R16055 GND.n7435 GND.n7434 585
R16056 GND.n4373 GND.n4371 585
R16057 GND.n4371 GND.n4360 585
R16058 GND.n4348 GND.n4347 585
R16059 GND.n4359 GND.n4348 585
R16060 GND.n7450 GND.n7449 585
R16061 GND.n7449 GND.n7448 585
R16062 GND.n7451 GND.n4342 585
R16063 GND.n5522 GND.n4342 585
R16064 GND.n7453 GND.n7452 585
R16065 GND.n7454 GND.n7453 585
R16066 GND.n4328 GND.n4327 585
R16067 GND.n6172 GND.n4328 585
R16068 GND.n7462 GND.n7461 585
R16069 GND.n7461 GND.n7460 585
R16070 GND.n7463 GND.n4322 585
R16071 GND.n5532 GND.n4322 585
R16072 GND.n7465 GND.n7464 585
R16073 GND.n7466 GND.n7465 585
R16074 GND.n4308 GND.n4307 585
R16075 GND.n5537 GND.n4308 585
R16076 GND.n7474 GND.n7473 585
R16077 GND.n7473 GND.n7472 585
R16078 GND.n7475 GND.n4302 585
R16079 GND.n5542 GND.n4302 585
R16080 GND.n7477 GND.n7476 585
R16081 GND.n7478 GND.n7477 585
R16082 GND.n4276 GND.n4275 585
R16083 GND.n5547 GND.n4276 585
R16084 GND.n7486 GND.n7485 585
R16085 GND.n7485 GND.n7484 585
R16086 GND.n7487 GND.n4268 585
R16087 GND.n6107 GND.n4268 585
R16088 GND.n7489 GND.n7488 585
R16089 GND.n7490 GND.n7489 585
R16090 GND.n4269 GND.n4267 585
R16091 GND.n4267 GND.n4256 585
R16092 GND.n4244 GND.n4243 585
R16093 GND.n4255 GND.n4244 585
R16094 GND.n7505 GND.n7504 585
R16095 GND.n7504 GND.n7503 585
R16096 GND.n7506 GND.n4238 585
R16097 GND.n5554 GND.n4238 585
R16098 GND.n7508 GND.n7507 585
R16099 GND.n7509 GND.n7508 585
R16100 GND.n4225 GND.n4224 585
R16101 GND.n6069 GND.n4225 585
R16102 GND.n7517 GND.n7516 585
R16103 GND.n7516 GND.n7515 585
R16104 GND.n7518 GND.n4219 585
R16105 GND.n5565 GND.n4219 585
R16106 GND.n7520 GND.n7519 585
R16107 GND.n7521 GND.n7520 585
R16108 GND.n4205 GND.n4204 585
R16109 GND.n5570 GND.n4205 585
R16110 GND.n7529 GND.n7528 585
R16111 GND.n7528 GND.n7527 585
R16112 GND.n7530 GND.n4199 585
R16113 GND.n5575 GND.n4199 585
R16114 GND.n7532 GND.n7531 585
R16115 GND.n7533 GND.n7532 585
R16116 GND.n4173 GND.n4172 585
R16117 GND.n5581 GND.n4173 585
R16118 GND.n7541 GND.n7540 585
R16119 GND.n7540 GND.n7539 585
R16120 GND.n7542 GND.n4165 585
R16121 GND.n6004 GND.n4165 585
R16122 GND.n7544 GND.n7543 585
R16123 GND.n7545 GND.n7544 585
R16124 GND.n4166 GND.n4164 585
R16125 GND.n4164 GND.n4153 585
R16126 GND.n4141 GND.n4140 585
R16127 GND.n4152 GND.n4141 585
R16128 GND.n7560 GND.n7559 585
R16129 GND.n7559 GND.n7558 585
R16130 GND.n7561 GND.n4135 585
R16131 GND.n5587 GND.n4135 585
R16132 GND.n7563 GND.n7562 585
R16133 GND.n7564 GND.n7563 585
R16134 GND.n4121 GND.n4120 585
R16135 GND.n5966 GND.n4121 585
R16136 GND.n7572 GND.n7571 585
R16137 GND.n7571 GND.n7570 585
R16138 GND.n7573 GND.n4115 585
R16139 GND.n5597 GND.n4115 585
R16140 GND.n7575 GND.n7574 585
R16141 GND.n7576 GND.n7575 585
R16142 GND.n4101 GND.n4100 585
R16143 GND.n5602 GND.n4101 585
R16144 GND.n7584 GND.n7583 585
R16145 GND.n7583 GND.n7582 585
R16146 GND.n7585 GND.n4095 585
R16147 GND.n5607 GND.n4095 585
R16148 GND.n7587 GND.n7586 585
R16149 GND.n7588 GND.n7587 585
R16150 GND.n4068 GND.n4067 585
R16151 GND.n5612 GND.n4068 585
R16152 GND.n7596 GND.n7595 585
R16153 GND.n7595 GND.n7594 585
R16154 GND.n7597 GND.n4060 585
R16155 GND.n5901 GND.n4060 585
R16156 GND.n7599 GND.n7598 585
R16157 GND.n7600 GND.n7599 585
R16158 GND.n4061 GND.n4059 585
R16159 GND.n4059 GND.n4048 585
R16160 GND.n4036 GND.n4035 585
R16161 GND.n4047 GND.n4036 585
R16162 GND.n7615 GND.n7614 585
R16163 GND.n7614 GND.n7613 585
R16164 GND.n7616 GND.n4030 585
R16165 GND.n5618 GND.n4030 585
R16166 GND.n7618 GND.n7617 585
R16167 GND.n7619 GND.n7618 585
R16168 GND.n4016 GND.n4015 585
R16169 GND.n5863 GND.n4016 585
R16170 GND.n7627 GND.n7626 585
R16171 GND.n7626 GND.n7625 585
R16172 GND.n7628 GND.n4010 585
R16173 GND.n5628 GND.n4010 585
R16174 GND.n7630 GND.n7629 585
R16175 GND.n7631 GND.n7630 585
R16176 GND.n3996 GND.n3995 585
R16177 GND.n5633 GND.n3996 585
R16178 GND.n7639 GND.n7638 585
R16179 GND.n7638 GND.n7637 585
R16180 GND.n7640 GND.n3990 585
R16181 GND.n5638 GND.n3990 585
R16182 GND.n7642 GND.n7641 585
R16183 GND.n7643 GND.n7642 585
R16184 GND.n3963 GND.n3962 585
R16185 GND.n5643 GND.n3963 585
R16186 GND.n7651 GND.n7650 585
R16187 GND.n7650 GND.n7649 585
R16188 GND.n7652 GND.n3955 585
R16189 GND.n5797 GND.n3955 585
R16190 GND.n7654 GND.n7653 585
R16191 GND.n7655 GND.n7654 585
R16192 GND.n3956 GND.n3954 585
R16193 GND.n3954 GND.n3944 585
R16194 GND.n3932 GND.n3931 585
R16195 GND.n3943 GND.n3932 585
R16196 GND.n7670 GND.n7669 585
R16197 GND.n7669 GND.n7668 585
R16198 GND.n7671 GND.n3926 585
R16199 GND.n5649 GND.n3926 585
R16200 GND.n7673 GND.n7672 585
R16201 GND.n7674 GND.n7673 585
R16202 GND.n3912 GND.n3911 585
R16203 GND.n5759 GND.n3912 585
R16204 GND.n7682 GND.n7681 585
R16205 GND.n7681 GND.n7680 585
R16206 GND.n7683 GND.n3906 585
R16207 GND.n5659 GND.n3906 585
R16208 GND.n7685 GND.n7684 585
R16209 GND.t41 GND.n7685 585
R16210 GND.n3893 GND.n3892 585
R16211 GND.n5664 GND.n3893 585
R16212 GND.n7693 GND.n7692 585
R16213 GND.n7692 GND.n7691 585
R16214 GND.n7694 GND.n3887 585
R16215 GND.n5685 GND.n3887 585
R16216 GND.n7696 GND.n7695 585
R16217 GND.n7697 GND.n7696 585
R16218 GND.n2326 GND.n2325 585
R16219 GND.n5690 GND.n2326 585
R16220 GND.n7762 GND.n7761 585
R16221 GND.n7761 GND.n7760 585
R16222 GND.n7763 GND.n2318 585
R16223 GND.n5694 GND.n2318 585
R16224 GND.n7765 GND.n7764 585
R16225 GND.n7766 GND.n7765 585
R16226 GND.n2319 GND.n2317 585
R16227 GND.n2317 GND.n2305 585
R16228 GND.n2106 GND.n2105 585
R16229 GND.n2304 GND.n2106 585
R16230 GND.n7781 GND.n7780 585
R16231 GND.n7780 GND.n7779 585
R16232 GND.n7782 GND.n2100 585
R16233 GND.n2107 GND.n2100 585
R16234 GND.n7784 GND.n7783 585
R16235 GND.n7785 GND.n7784 585
R16236 GND.n2088 GND.n2087 585
R16237 GND.n2091 GND.n2088 585
R16238 GND.n7795 GND.n7794 585
R16239 GND.n7794 GND.n7793 585
R16240 GND.n7796 GND.n2082 585
R16241 GND.n2288 GND.n2082 585
R16242 GND.n7798 GND.n7797 585
R16243 GND.n7799 GND.n7798 585
R16244 GND.n2070 GND.n2069 585
R16245 GND.n2073 GND.n2070 585
R16246 GND.n7809 GND.n7808 585
R16247 GND.n7808 GND.n7807 585
R16248 GND.n7810 GND.n2064 585
R16249 GND.n2275 GND.n2064 585
R16250 GND.n7812 GND.n7811 585
R16251 GND.n7813 GND.n7812 585
R16252 GND.n2052 GND.n2051 585
R16253 GND.n2055 GND.n2052 585
R16254 GND.n7823 GND.n7822 585
R16255 GND.n7822 GND.n7821 585
R16256 GND.n7824 GND.n2046 585
R16257 GND.n2262 GND.n2046 585
R16258 GND.n7826 GND.n7825 585
R16259 GND.n7827 GND.n7826 585
R16260 GND.n2034 GND.n2033 585
R16261 GND.n2037 GND.n2034 585
R16262 GND.n7837 GND.n7836 585
R16263 GND.n7836 GND.n7835 585
R16264 GND.n7838 GND.n2028 585
R16265 GND.n2252 GND.n2028 585
R16266 GND.n7840 GND.n7839 585
R16267 GND.n7841 GND.n7840 585
R16268 GND.n2016 GND.n2015 585
R16269 GND.n2025 GND.n2016 585
R16270 GND.n7851 GND.n7850 585
R16271 GND.n7850 GND.n7849 585
R16272 GND.n7852 GND.n2010 585
R16273 GND.n2237 GND.n2010 585
R16274 GND.n7854 GND.n7853 585
R16275 GND.n7855 GND.n7854 585
R16276 GND.n1998 GND.n1997 585
R16277 GND.n2007 GND.n1998 585
R16278 GND.n7865 GND.n7864 585
R16279 GND.n7864 GND.n7863 585
R16280 GND.n7866 GND.n1992 585
R16281 GND.n2224 GND.n1992 585
R16282 GND.n7868 GND.n7867 585
R16283 GND.n7869 GND.n7868 585
R16284 GND.n1980 GND.n1979 585
R16285 GND.n1989 GND.n1980 585
R16286 GND.n7879 GND.n7878 585
R16287 GND.n7878 GND.n7877 585
R16288 GND.n7880 GND.n1974 585
R16289 GND.n2211 GND.n1974 585
R16290 GND.n7882 GND.n7881 585
R16291 GND.n7883 GND.n7882 585
R16292 GND.n1963 GND.n1962 585
R16293 GND.n1971 GND.n1963 585
R16294 GND.n7893 GND.n7892 585
R16295 GND.n7892 GND.n7891 585
R16296 GND.n7894 GND.n1957 585
R16297 GND.n2201 GND.n1957 585
R16298 GND.n7896 GND.n7895 585
R16299 GND.n7897 GND.n7896 585
R16300 GND.n1946 GND.n1945 585
R16301 GND.n1949 GND.n1946 585
R16302 GND.n7906 GND.n7905 585
R16303 GND.n7905 GND.n7904 585
R16304 GND.n7907 GND.n1940 585
R16305 GND.n2187 GND.n1940 585
R16306 GND.n7909 GND.n7908 585
R16307 GND.n7910 GND.n7909 585
R16308 GND.n1941 GND.n1939 585
R16309 GND.n1939 GND.n1938 585
R16310 GND.n3431 GND.n3426 585
R16311 GND.n3426 GND.n1905 585
R16312 GND.n3433 GND.n3432 585
R16313 GND.n3433 GND.n1876 585
R16314 GND.n3434 GND.n3425 585
R16315 GND.n3435 GND.n3434 585
R16316 GND.n3438 GND.n3437 585
R16317 GND.n3437 GND.n3436 585
R16318 GND.n3439 GND.n3420 585
R16319 GND.n3420 GND.n1707 585
R16320 GND.n3441 GND.n3440 585
R16321 GND.n3441 GND.n1683 585
R16322 GND.n3442 GND.n3419 585
R16323 GND.n3442 GND.n1679 585
R16324 GND.n3444 GND.n3443 585
R16325 GND.n3443 GND.n1676 585
R16326 GND.n3445 GND.n3414 585
R16327 GND.n3414 GND.n2362 585
R16328 GND.n3447 GND.n3446 585
R16329 GND.n3447 GND.n2370 585
R16330 GND.n3448 GND.n3413 585
R16331 GND.n3448 GND.n2368 585
R16332 GND.n3450 GND.n3449 585
R16333 GND.n3449 GND.n2372 585
R16334 GND.n3451 GND.n3408 585
R16335 GND.n3408 GND.n2379 585
R16336 GND.n3453 GND.n3452 585
R16337 GND.n3453 GND.n2378 585
R16338 GND.n3454 GND.n3407 585
R16339 GND.n3454 GND.n2391 585
R16340 GND.n3456 GND.n3455 585
R16341 GND.n3455 GND.n2389 585
R16342 GND.n3457 GND.n3402 585
R16343 GND.n3402 GND.n2393 585
R16344 GND.n3459 GND.n3458 585
R16345 GND.n3459 GND.n2401 585
R16346 GND.n3460 GND.n3401 585
R16347 GND.n3460 GND.n2400 585
R16348 GND.n3462 GND.n3461 585
R16349 GND.n3461 GND.n2414 585
R16350 GND.n3463 GND.n3396 585
R16351 GND.n3396 GND.n2411 585
R16352 GND.n3465 GND.n3464 585
R16353 GND.n3465 GND.n2417 585
R16354 GND.n3466 GND.n3395 585
R16355 GND.n3466 GND.n2424 585
R16356 GND.n3468 GND.n3467 585
R16357 GND.n3467 GND.n2423 585
R16358 GND.n3469 GND.n3390 585
R16359 GND.n3390 GND.n2435 585
R16360 GND.n3471 GND.n3470 585
R16361 GND.n3471 GND.n2433 585
R16362 GND.n3472 GND.n3389 585
R16363 GND.n3472 GND.n2438 585
R16364 GND.n3476 GND.n3475 585
R16365 GND.n3475 GND.n3474 585
R16366 GND.n3477 GND.n3384 585
R16367 GND.n3384 GND.n2444 585
R16368 GND.n3479 GND.n3478 585
R16369 GND.n3479 GND.n2455 585
R16370 GND.n3480 GND.n3383 585
R16371 GND.n3480 GND.n2453 585
R16372 GND.n3482 GND.n3481 585
R16373 GND.n3481 GND.n2457 585
R16374 GND.n3483 GND.n3378 585
R16375 GND.n3378 GND.n2464 585
R16376 GND.n3485 GND.n3484 585
R16377 GND.n3485 GND.n2463 585
R16378 GND.n3486 GND.n3377 585
R16379 GND.n3486 GND.n2476 585
R16380 GND.n3488 GND.n3487 585
R16381 GND.n3487 GND.n2474 585
R16382 GND.n3489 GND.n3372 585
R16383 GND.n3372 GND.n2478 585
R16384 GND.n3491 GND.n3490 585
R16385 GND.n3491 GND.n2486 585
R16386 GND.n3492 GND.n3371 585
R16387 GND.n3492 GND.n2485 585
R16388 GND.n3494 GND.n3493 585
R16389 GND.n3493 GND.n2499 585
R16390 GND.n3495 GND.n3366 585
R16391 GND.n3366 GND.n2496 585
R16392 GND.n3497 GND.n3496 585
R16393 GND.n3497 GND.n2502 585
R16394 GND.n3498 GND.n3365 585
R16395 GND.n3498 GND.n2509 585
R16396 GND.n3500 GND.n3499 585
R16397 GND.n3499 GND.n2508 585
R16398 GND.n3501 GND.n3360 585
R16399 GND.n3360 GND.n2520 585
R16400 GND.n3503 GND.n3502 585
R16401 GND.n3503 GND.n2518 585
R16402 GND.n3504 GND.n3359 585
R16403 GND.n3504 GND.n2523 585
R16404 GND.n3506 GND.n3505 585
R16405 GND.n3505 GND.n2531 585
R16406 GND.n3507 GND.n3354 585
R16407 GND.n3354 GND.n2529 585
R16408 GND.n3509 GND.n3508 585
R16409 GND.n3509 GND.n2542 585
R16410 GND.n3510 GND.n3353 585
R16411 GND.n3510 GND.n2540 585
R16412 GND.n3512 GND.n3511 585
R16413 GND.n3511 GND.n2544 585
R16414 GND.n3513 GND.n3348 585
R16415 GND.n3348 GND.n2551 585
R16416 GND.n3515 GND.n3514 585
R16417 GND.n3515 GND.n2550 585
R16418 GND.n3516 GND.n3347 585
R16419 GND.n3516 GND.n2563 585
R16420 GND.n3518 GND.n3517 585
R16421 GND.n3517 GND.n2561 585
R16422 GND.n3519 GND.n3342 585
R16423 GND.n3342 GND.n2565 585
R16424 GND.n3521 GND.n3520 585
R16425 GND.n3521 GND.n2573 585
R16426 GND.n3522 GND.n3341 585
R16427 GND.n3522 GND.n2572 585
R16428 GND.n3524 GND.n3523 585
R16429 GND.n3523 GND.n2586 585
R16430 GND.n3525 GND.n3336 585
R16431 GND.n3336 GND.n2583 585
R16432 GND.n3527 GND.n3526 585
R16433 GND.n3527 GND.n2587 585
R16434 GND.n3528 GND.n3335 585
R16435 GND.n3528 GND.n1555 585
R16436 GND.n3530 GND.n3529 585
R16437 GND.n3529 GND.n1552 585
R16438 GND.n3532 GND.n3334 585
R16439 GND.n3334 GND.n2596 585
R16440 GND.n3534 GND.n3533 585
R16441 GND.n3534 GND.n2599 585
R16442 GND.n3536 GND.n3535 585
R16443 GND.n3535 GND.n1535 585
R16444 GND.n3537 GND.n2612 585
R16445 GND.n2612 GND.n1533 585
R16446 GND.n3540 GND.n3539 585
R16447 GND.n3541 GND.n3540 585
R16448 GND.n3332 GND.n2611 585
R16449 GND.n2618 GND.n2611 585
R16450 GND.n3330 GND.n3329 585
R16451 GND.n3329 GND.n3328 585
R16452 GND.n2614 GND.n2613 585
R16453 GND.n2624 GND.n2614 585
R16454 GND.n3303 GND.n2635 585
R16455 GND.n2635 GND.n2622 585
R16456 GND.n3305 GND.n3304 585
R16457 GND.n3306 GND.n3305 585
R16458 GND.n2636 GND.n2634 585
R16459 GND.n2642 GND.n2634 585
R16460 GND.n3298 GND.n3297 585
R16461 GND.n3297 GND.n3296 585
R16462 GND.n2639 GND.n2638 585
R16463 GND.n2653 GND.n2639 585
R16464 GND.n3265 GND.n2664 585
R16465 GND.n2664 GND.n2650 585
R16466 GND.n3267 GND.n3266 585
R16467 GND.n3268 GND.n3267 585
R16468 GND.n2665 GND.n2663 585
R16469 GND.n2672 GND.n2663 585
R16470 GND.n3260 GND.n3259 585
R16471 GND.n3259 GND.n3258 585
R16472 GND.n2668 GND.n2667 585
R16473 GND.n2682 GND.n2668 585
R16474 GND.n3228 GND.n2693 585
R16475 GND.n2693 GND.n2680 585
R16476 GND.n3230 GND.n3229 585
R16477 GND.n3231 GND.n3230 585
R16478 GND.n2694 GND.n2692 585
R16479 GND.n2701 GND.n2692 585
R16480 GND.n3223 GND.n3222 585
R16481 GND.n3222 GND.n3221 585
R16482 GND.n2697 GND.n2696 585
R16483 GND.n2711 GND.n2697 585
R16484 GND.n3191 GND.n2723 585
R16485 GND.n2723 GND.n2709 585
R16486 GND.n3193 GND.n3192 585
R16487 GND.n3194 GND.n3193 585
R16488 GND.n2724 GND.n2722 585
R16489 GND.n2730 GND.n2722 585
R16490 GND.n3186 GND.n3185 585
R16491 GND.n3185 GND.n3184 585
R16492 GND.n2727 GND.n2726 585
R16493 GND.n2740 GND.n2727 585
R16494 GND.n3153 GND.n2751 585
R16495 GND.n2751 GND.n2738 585
R16496 GND.n3155 GND.n3154 585
R16497 GND.n3156 GND.n3155 585
R16498 GND.n2752 GND.n2750 585
R16499 GND.n2757 GND.n2750 585
R16500 GND.n3148 GND.n3147 585
R16501 GND.n3147 GND.n3146 585
R16502 GND.n2755 GND.n2754 585
R16503 GND.n2768 GND.n2755 585
R16504 GND.n3115 GND.n2779 585
R16505 GND.n2779 GND.n2765 585
R16506 GND.n3117 GND.n3116 585
R16507 GND.n3118 GND.n3117 585
R16508 GND.n2780 GND.n2778 585
R16509 GND.n2787 GND.n2778 585
R16510 GND.n3110 GND.n3109 585
R16511 GND.n3109 GND.n3108 585
R16512 GND.n2783 GND.n2782 585
R16513 GND.n2797 GND.n2783 585
R16514 GND.n3078 GND.n2808 585
R16515 GND.n2808 GND.n2795 585
R16516 GND.n3080 GND.n3079 585
R16517 GND.n3081 GND.n3080 585
R16518 GND.n2809 GND.n2807 585
R16519 GND.n2816 GND.n2807 585
R16520 GND.n3073 GND.n3072 585
R16521 GND.n3072 GND.n3071 585
R16522 GND.n2812 GND.n2811 585
R16523 GND.n2825 GND.n2812 585
R16524 GND.n3043 GND.n3042 585
R16525 GND.n3044 GND.n3043 585
R16526 GND.n2836 GND.n2835 585
R16527 GND.n2835 GND.n2834 585
R16528 GND.n3038 GND.n3037 585
R16529 GND.n3037 GND.n3036 585
R16530 GND.n2839 GND.n2838 585
R16531 GND.n2850 GND.n2839 585
R16532 GND.n3014 GND.n3007 585
R16533 GND.n3007 GND.n2848 585
R16534 GND.n3016 GND.n3015 585
R16535 GND.n3017 GND.n3016 585
R16536 GND.n3008 GND.n3006 585
R16537 GND.n3006 GND.n3005 585
R16538 GND.n3009 GND.n1321 585
R16539 GND.n2863 GND.n1321 585
R16540 GND.n8025 GND.n1672 585
R16541 GND.n8026 GND.n8025 585
R16542 GND.n1680 GND.n1671 585
R16543 GND.n3843 GND.n1680 585
R16544 GND.n3831 GND.n1670 585
R16545 GND.n3831 GND.n3830 585
R16546 GND.n3833 GND.n3832 585
R16547 GND.n3834 GND.n3833 585
R16548 GND.n3829 GND.n1664 585
R16549 GND.n3829 GND.n3828 585
R16550 GND.n2371 GND.n1663 585
R16551 GND.n2383 GND.n2371 585
R16552 GND.n2380 GND.n1662 585
R16553 GND.n3817 GND.n2380 585
R16554 GND.n3805 GND.n3803 585
R16555 GND.n3805 GND.n3804 585
R16556 GND.n3806 GND.n1656 585
R16557 GND.n3807 GND.n3806 585
R16558 GND.n3802 GND.n1655 585
R16559 GND.n3802 GND.n3801 585
R16560 GND.n2392 GND.n1654 585
R16561 GND.n2405 GND.n2392 585
R16562 GND.n2403 GND.n2402 585
R16563 GND.n3791 GND.n2403 585
R16564 GND.n3779 GND.n1648 585
R16565 GND.n3779 GND.n3778 585
R16566 GND.n3780 GND.n1647 585
R16567 GND.n3781 GND.n3780 585
R16568 GND.n3777 GND.n1646 585
R16569 GND.n3777 GND.n3776 585
R16570 GND.n2416 GND.n2415 585
R16571 GND.n2427 GND.n2416 585
R16572 GND.n2425 GND.n1640 585
R16573 GND.n3766 GND.n2425 585
R16574 GND.n3754 GND.n1639 585
R16575 GND.n3754 GND.n3753 585
R16576 GND.n3755 GND.n1638 585
R16577 GND.n3756 GND.n3755 585
R16578 GND.n3751 GND.n2437 585
R16579 GND.n3751 GND.n3750 585
R16580 GND.n2436 GND.n1632 585
R16581 GND.n3473 GND.n2436 585
R16582 GND.n2446 GND.n1631 585
R16583 GND.n3740 GND.n2446 585
R16584 GND.n3727 GND.n1630 585
R16585 GND.n3727 GND.n3726 585
R16586 GND.n3729 GND.n3728 585
R16587 GND.n3730 GND.n3729 585
R16588 GND.n3725 GND.n1624 585
R16589 GND.n3725 GND.n3724 585
R16590 GND.n2456 GND.n1623 585
R16591 GND.n2468 GND.n2456 585
R16592 GND.n2465 GND.n1622 585
R16593 GND.n3714 GND.n2465 585
R16594 GND.n3702 GND.n3700 585
R16595 GND.n3702 GND.n3701 585
R16596 GND.n3703 GND.n1616 585
R16597 GND.n3704 GND.n3703 585
R16598 GND.n3699 GND.n1615 585
R16599 GND.n3699 GND.n3698 585
R16600 GND.n2477 GND.n1614 585
R16601 GND.n2490 GND.n2477 585
R16602 GND.n2488 GND.n2487 585
R16603 GND.n3688 GND.n2488 585
R16604 GND.n3676 GND.n1608 585
R16605 GND.n3676 GND.n3675 585
R16606 GND.n3677 GND.n1607 585
R16607 GND.n3678 GND.n3677 585
R16608 GND.n3674 GND.n1606 585
R16609 GND.n3674 GND.n3673 585
R16610 GND.n2501 GND.n2500 585
R16611 GND.n2512 GND.n2501 585
R16612 GND.n2510 GND.n1600 585
R16613 GND.n3663 GND.n2510 585
R16614 GND.n3651 GND.n1599 585
R16615 GND.n3651 GND.n3650 585
R16616 GND.n3652 GND.n1598 585
R16617 GND.n3653 GND.n3652 585
R16618 GND.n3648 GND.n2522 585
R16619 GND.n3648 GND.n3647 585
R16620 GND.n2521 GND.n1592 585
R16621 GND.n2534 GND.n2521 585
R16622 GND.n2532 GND.n1591 585
R16623 GND.n3637 GND.n2532 585
R16624 GND.n3624 GND.n1590 585
R16625 GND.n3624 GND.n3623 585
R16626 GND.n3626 GND.n3625 585
R16627 GND.n3627 GND.n3626 585
R16628 GND.n3622 GND.n1584 585
R16629 GND.n3622 GND.n3621 585
R16630 GND.n2543 GND.n1583 585
R16631 GND.n2555 GND.n2543 585
R16632 GND.n2552 GND.n1582 585
R16633 GND.n3611 GND.n2552 585
R16634 GND.n3599 GND.n3597 585
R16635 GND.n3599 GND.n3598 585
R16636 GND.n3600 GND.n1576 585
R16637 GND.n3601 GND.n3600 585
R16638 GND.n3596 GND.n1575 585
R16639 GND.n3596 GND.n3595 585
R16640 GND.n2564 GND.n1574 585
R16641 GND.n2577 GND.n2564 585
R16642 GND.n2575 GND.n2574 585
R16643 GND.n3585 GND.n2575 585
R16644 GND.n3573 GND.n1568 585
R16645 GND.n3573 GND.n3572 585
R16646 GND.n3574 GND.n1567 585
R16647 GND.n3575 GND.n3574 585
R16648 GND.n3571 GND.n1566 585
R16649 GND.n3571 GND.n3570 585
R16650 GND.n1559 GND.n1557 585
R16651 GND.n2588 GND.n1557 585
R16652 GND.n8115 GND.n8114 585
R16653 GND.n8116 GND.n8115 585
R16654 GND.n1558 GND.n1556 585
R16655 GND.n3559 GND.n1556 585
R16656 GND.n3553 GND.n3552 585
R16657 GND.n3556 GND.n3553 585
R16658 GND.n2602 GND.n2601 585
R16659 GND.n2601 GND.n2600 585
R16660 GND.n3544 GND.n1536 585
R16661 GND.n8123 GND.n1536 585
R16662 GND.n3545 GND.n3543 585
R16663 GND.n3543 GND.n3542 585
R16664 GND.n2608 GND.n2607 585
R16665 GND.n2610 GND.n2608 585
R16666 GND.n3312 GND.n2619 585
R16667 GND.n3327 GND.n2619 585
R16668 GND.n2628 GND.n2626 585
R16669 GND.n2626 GND.n2615 585
R16670 GND.n3319 GND.n3318 585
R16671 GND.n3320 GND.n3319 585
R16672 GND.n2627 GND.n2625 585
R16673 GND.n3308 GND.n2625 585
R16674 GND.n3275 GND.n3274 585
R16675 GND.n3274 GND.n2633 585
R16676 GND.n3273 GND.n2643 585
R16677 GND.n3295 GND.n2643 585
R16678 GND.n2657 GND.n2655 585
R16679 GND.n2655 GND.n2640 585
R16680 GND.n3283 GND.n3282 585
R16681 GND.n3284 GND.n3283 585
R16682 GND.n2656 GND.n2654 585
R16683 GND.n3269 GND.n2654 585
R16684 GND.n3238 GND.n3237 585
R16685 GND.n3237 GND.n2662 585
R16686 GND.n3236 GND.n2673 585
R16687 GND.n3257 GND.n2673 585
R16688 GND.n2686 GND.n2684 585
R16689 GND.n2684 GND.n2670 585
R16690 GND.n3246 GND.n3245 585
R16691 GND.n3247 GND.n3246 585
R16692 GND.n2685 GND.n2683 585
R16693 GND.n3232 GND.n2683 585
R16694 GND.n3201 GND.n3200 585
R16695 GND.n3200 GND.n2691 585
R16696 GND.n3199 GND.n2702 585
R16697 GND.n3220 GND.n2702 585
R16698 GND.n2715 GND.n2713 585
R16699 GND.n2713 GND.n2698 585
R16700 GND.n3209 GND.n3208 585
R16701 GND.n3210 GND.n3209 585
R16702 GND.n2714 GND.n2712 585
R16703 GND.n3195 GND.n2712 585
R16704 GND.n3164 GND.n3163 585
R16705 GND.n3163 GND.n2721 585
R16706 GND.n3162 GND.n2731 585
R16707 GND.n3183 GND.n2731 585
R16708 GND.n2744 GND.n2742 585
R16709 GND.n2742 GND.n2728 585
R16710 GND.n3172 GND.n3171 585
R16711 GND.n3173 GND.n3172 585
R16712 GND.n2743 GND.n2741 585
R16713 GND.n3158 GND.n2741 585
R16714 GND.n3126 GND.n3125 585
R16715 GND.n3125 GND.n2749 585
R16716 GND.n3124 GND.n2758 585
R16717 GND.n3145 GND.n2758 585
R16718 GND.n2772 GND.n2770 585
R16719 GND.n3122 GND.n2770 585
R16720 GND.n3134 GND.n3133 585
R16721 GND.n3135 GND.n3134 585
R16722 GND.n2771 GND.n2769 585
R16723 GND.n3119 GND.n2769 585
R16724 GND.n3088 GND.n3087 585
R16725 GND.n3087 GND.n2777 585
R16726 GND.n3086 GND.n2788 585
R16727 GND.n3107 GND.n2788 585
R16728 GND.n2801 GND.n2799 585
R16729 GND.n2799 GND.n2785 585
R16730 GND.n3096 GND.n3095 585
R16731 GND.n3097 GND.n3096 585
R16732 GND.n2800 GND.n2798 585
R16733 GND.n3082 GND.n2798 585
R16734 GND.n3051 GND.n3050 585
R16735 GND.n3050 GND.n2806 585
R16736 GND.n3049 GND.n2817 585
R16737 GND.n3070 GND.n2817 585
R16738 GND.n2829 GND.n2827 585
R16739 GND.n2827 GND.n2813 585
R16740 GND.n3059 GND.n3058 585
R16741 GND.n3060 GND.n3059 585
R16742 GND.n2828 GND.n2826 585
R16743 GND.n3045 GND.n2826 585
R16744 GND.n2856 GND.n2842 585
R16745 GND.n3035 GND.n2842 585
R16746 GND.n2854 GND.n2852 585
R16747 GND.n2852 GND.n2840 585
R16748 GND.n3026 GND.n3025 585
R16749 GND.n3027 GND.n3026 585
R16750 GND.n2853 GND.n2851 585
R16751 GND.n3018 GND.n2851 585
R16752 GND.n2985 GND.n2984 585
R16753 GND.n2984 GND.n2862 585
R16754 GND.n2983 GND.n2865 585
R16755 GND.n3004 GND.n2865 585
R16756 GND.n2879 GND.n2877 585
R16757 GND.n2877 GND.n2875 585
R16758 GND.n2993 GND.n2992 585
R16759 GND.n2994 GND.n2993 585
R16760 GND.n2878 GND.n2876 585
R16761 GND.n2876 GND.n2873 585
R16762 GND.n2899 GND.n2885 585
R16763 GND.n2978 GND.n2885 585
R16764 GND.n2897 GND.n2895 585
R16765 GND.n2895 GND.n2884 585
R16766 GND.n2969 GND.n2968 585
R16767 GND.n2970 GND.n2969 585
R16768 GND.n2896 GND.n2894 585
R16769 GND.n2894 GND.n2892 585
R16770 GND.n2919 GND.n2905 585
R16771 GND.n2961 GND.n2905 585
R16772 GND.n2917 GND.n2915 585
R16773 GND.n2915 GND.n2904 585
R16774 GND.n2952 GND.n2951 585
R16775 GND.n2953 GND.n2952 585
R16776 GND.n2916 GND.n2914 585
R16777 GND.n2914 GND.n2912 585
R16778 GND.n2935 GND.n2934 585
R16779 GND.n2944 GND.n2935 585
R16780 GND.n2928 GND.n2925 585
R16781 GND.n2925 GND.n2924 585
R16782 GND.n2927 GND.n2926 585
R16783 GND.n2926 GND.n1358 585
R16784 GND.n8237 GND.n1359 585
R16785 GND.n8362 GND.n1359 585
R16786 GND.n8236 GND.n1439 585
R16787 GND.n8235 GND.n1440 585
R16788 GND.n1442 GND.n1441 585
R16789 GND.n8231 GND.n1444 585
R16790 GND.n8230 GND.n1445 585
R16791 GND.n8229 GND.n1446 585
R16792 GND.n1448 GND.n1447 585
R16793 GND.n8225 GND.n1450 585
R16794 GND.n8224 GND.n1451 585
R16795 GND.n8223 GND.n8220 585
R16796 GND.n1452 GND.n1357 585
R16797 GND.n8362 GND.n1357 585
R16798 GND.n3846 GND.n1678 585
R16799 GND.n8026 GND.n1678 585
R16800 GND.n3845 GND.n3844 585
R16801 GND.n3844 GND.n3843 585
R16802 GND.n2361 GND.n2360 585
R16803 GND.n3830 GND.n2361 585
R16804 GND.n3825 GND.n2369 585
R16805 GND.n3834 GND.n2369 585
R16806 GND.n3827 GND.n3826 585
R16807 GND.n3828 GND.n3827 585
R16808 GND.n2374 GND.n2373 585
R16809 GND.n2383 GND.n2373 585
R16810 GND.n3819 GND.n3818 585
R16811 GND.n3818 GND.n3817 585
R16812 GND.n2377 GND.n2376 585
R16813 GND.n3804 GND.n2377 585
R16814 GND.n3798 GND.n2390 585
R16815 GND.n3807 GND.n2390 585
R16816 GND.n3800 GND.n3799 585
R16817 GND.n3801 GND.n3800 585
R16818 GND.n2396 GND.n2395 585
R16819 GND.n2405 GND.n2395 585
R16820 GND.n3793 GND.n3792 585
R16821 GND.n3792 GND.n3791 585
R16822 GND.n2399 GND.n2398 585
R16823 GND.n3778 GND.n2399 585
R16824 GND.n3773 GND.n2413 585
R16825 GND.n3781 GND.n2413 585
R16826 GND.n3775 GND.n3774 585
R16827 GND.n3776 GND.n3775 585
R16828 GND.n2419 GND.n2418 585
R16829 GND.n2427 GND.n2418 585
R16830 GND.n3768 GND.n3767 585
R16831 GND.n3767 GND.n3766 585
R16832 GND.n2422 GND.n2421 585
R16833 GND.n3753 GND.n2422 585
R16834 GND.n3747 GND.n2434 585
R16835 GND.n3756 GND.n2434 585
R16836 GND.n3749 GND.n3748 585
R16837 GND.n3750 GND.n3749 585
R16838 GND.n2440 GND.n2439 585
R16839 GND.n3473 GND.n2439 585
R16840 GND.n3742 GND.n3741 585
R16841 GND.n3741 GND.n3740 585
R16842 GND.n2443 GND.n2442 585
R16843 GND.n3726 GND.n2443 585
R16844 GND.n3721 GND.n2454 585
R16845 GND.n3730 GND.n2454 585
R16846 GND.n3723 GND.n3722 585
R16847 GND.n3724 GND.n3723 585
R16848 GND.n2459 GND.n2458 585
R16849 GND.n2468 GND.n2458 585
R16850 GND.n3716 GND.n3715 585
R16851 GND.n3715 GND.n3714 585
R16852 GND.n2462 GND.n2461 585
R16853 GND.n3701 GND.n2462 585
R16854 GND.n3695 GND.n2475 585
R16855 GND.n3704 GND.n2475 585
R16856 GND.n3697 GND.n3696 585
R16857 GND.n3698 GND.n3697 585
R16858 GND.n2481 GND.n2480 585
R16859 GND.n2490 GND.n2480 585
R16860 GND.n3690 GND.n3689 585
R16861 GND.n3689 GND.n3688 585
R16862 GND.n2484 GND.n2483 585
R16863 GND.n3675 GND.n2484 585
R16864 GND.n3670 GND.n2498 585
R16865 GND.n3678 GND.n2498 585
R16866 GND.n3672 GND.n3671 585
R16867 GND.n3673 GND.n3672 585
R16868 GND.n2504 GND.n2503 585
R16869 GND.n2512 GND.n2503 585
R16870 GND.n3665 GND.n3664 585
R16871 GND.n3664 GND.n3663 585
R16872 GND.n2507 GND.n2506 585
R16873 GND.n3650 GND.n2507 585
R16874 GND.n3644 GND.n2519 585
R16875 GND.n3653 GND.n2519 585
R16876 GND.n3646 GND.n3645 585
R16877 GND.n3647 GND.n3646 585
R16878 GND.n2525 GND.n2524 585
R16879 GND.n2534 GND.n2524 585
R16880 GND.n3639 GND.n3638 585
R16881 GND.n3638 GND.n3637 585
R16882 GND.n2528 GND.n2527 585
R16883 GND.n3623 GND.n2528 585
R16884 GND.n3618 GND.n2541 585
R16885 GND.n3627 GND.n2541 585
R16886 GND.n3620 GND.n3619 585
R16887 GND.n3621 GND.n3620 585
R16888 GND.n2546 GND.n2545 585
R16889 GND.n2555 GND.n2545 585
R16890 GND.n3613 GND.n3612 585
R16891 GND.n3612 GND.n3611 585
R16892 GND.n2549 GND.n2548 585
R16893 GND.n3598 GND.n2549 585
R16894 GND.n3592 GND.n2562 585
R16895 GND.n3601 GND.n2562 585
R16896 GND.n3594 GND.n3593 585
R16897 GND.n3595 GND.n3594 585
R16898 GND.n2568 GND.n2567 585
R16899 GND.n2577 GND.n2567 585
R16900 GND.n3587 GND.n3586 585
R16901 GND.n3586 GND.n3585 585
R16902 GND.n2571 GND.n2570 585
R16903 GND.n3572 GND.n2571 585
R16904 GND.n3567 GND.n2585 585
R16905 GND.n3575 GND.n2585 585
R16906 GND.n3569 GND.n3568 585
R16907 GND.n3570 GND.n3569 585
R16908 GND.n2590 GND.n2589 585
R16909 GND.n2589 GND.n2588 585
R16910 GND.n3562 GND.n1554 585
R16911 GND.n8116 GND.n1554 585
R16912 GND.n3561 GND.n3560 585
R16913 GND.n3560 GND.n3559 585
R16914 GND.n2595 GND.n2594 585
R16915 GND.n3556 GND.n2595 585
R16916 GND.n1532 GND.n1531 585
R16917 GND.n2600 GND.n1532 585
R16918 GND.n8125 GND.n8124 585
R16919 GND.n8124 GND.n8123 585
R16920 GND.n8126 GND.n1529 585
R16921 GND.n3542 GND.n1529 585
R16922 GND.n2609 GND.n1527 585
R16923 GND.n2610 GND.n2609 585
R16924 GND.n8130 GND.n1526 585
R16925 GND.n3327 GND.n1526 585
R16926 GND.n8131 GND.n1525 585
R16927 GND.n2615 GND.n1525 585
R16928 GND.n8132 GND.n1524 585
R16929 GND.n3320 GND.n1524 585
R16930 GND.n3307 GND.n1522 585
R16931 GND.n3308 GND.n3307 585
R16932 GND.n8136 GND.n1521 585
R16933 GND.n2633 GND.n1521 585
R16934 GND.n8137 GND.n1520 585
R16935 GND.n3295 GND.n1520 585
R16936 GND.n8138 GND.n1519 585
R16937 GND.n2640 GND.n1519 585
R16938 GND.n2652 GND.n1517 585
R16939 GND.n3284 GND.n2652 585
R16940 GND.n8142 GND.n1516 585
R16941 GND.n3269 GND.n1516 585
R16942 GND.n8143 GND.n1515 585
R16943 GND.n2662 GND.n1515 585
R16944 GND.n8144 GND.n1514 585
R16945 GND.n3257 GND.n1514 585
R16946 GND.n2669 GND.n1512 585
R16947 GND.n2670 GND.n2669 585
R16948 GND.n8148 GND.n1511 585
R16949 GND.n3247 GND.n1511 585
R16950 GND.n8149 GND.n1510 585
R16951 GND.n3232 GND.n1510 585
R16952 GND.n8150 GND.n1509 585
R16953 GND.n2691 GND.n1509 585
R16954 GND.n2700 GND.n1507 585
R16955 GND.n3220 GND.n2700 585
R16956 GND.n8154 GND.n1506 585
R16957 GND.n2698 GND.n1506 585
R16958 GND.n8155 GND.n1505 585
R16959 GND.n3210 GND.n1505 585
R16960 GND.n8156 GND.n1504 585
R16961 GND.n3195 GND.n1504 585
R16962 GND.n2720 GND.n1502 585
R16963 GND.n2721 GND.n2720 585
R16964 GND.n8160 GND.n1501 585
R16965 GND.n3183 GND.n1501 585
R16966 GND.n8161 GND.n1500 585
R16967 GND.n2728 GND.n1500 585
R16968 GND.n8162 GND.n1499 585
R16969 GND.n3173 GND.n1499 585
R16970 GND.n3157 GND.n1497 585
R16971 GND.n3158 GND.n3157 585
R16972 GND.n8166 GND.n1496 585
R16973 GND.n2749 GND.n1496 585
R16974 GND.n8167 GND.n1495 585
R16975 GND.n3145 GND.n1495 585
R16976 GND.n8168 GND.n1494 585
R16977 GND.n3122 GND.n1494 585
R16978 GND.n2767 GND.n1492 585
R16979 GND.n3135 GND.n2767 585
R16980 GND.n8172 GND.n1491 585
R16981 GND.n3119 GND.n1491 585
R16982 GND.n8173 GND.n1490 585
R16983 GND.n2777 GND.n1490 585
R16984 GND.n8174 GND.n1489 585
R16985 GND.n3107 GND.n1489 585
R16986 GND.n2784 GND.n1487 585
R16987 GND.n2785 GND.n2784 585
R16988 GND.n8178 GND.n1486 585
R16989 GND.n3097 GND.n1486 585
R16990 GND.n8179 GND.n1485 585
R16991 GND.n3082 GND.n1485 585
R16992 GND.n8180 GND.n1484 585
R16993 GND.n2806 GND.n1484 585
R16994 GND.n2815 GND.n1482 585
R16995 GND.n3070 GND.n2815 585
R16996 GND.n8184 GND.n1481 585
R16997 GND.n2813 GND.n1481 585
R16998 GND.n8185 GND.n1480 585
R16999 GND.n3060 GND.n1480 585
R17000 GND.n8186 GND.n1479 585
R17001 GND.n3045 GND.n1479 585
R17002 GND.n2841 GND.n1477 585
R17003 GND.n3035 GND.n2841 585
R17004 GND.n8190 GND.n1476 585
R17005 GND.n2840 GND.n1476 585
R17006 GND.n8191 GND.n1475 585
R17007 GND.n3027 GND.n1475 585
R17008 GND.n8192 GND.n1474 585
R17009 GND.n3018 GND.n1474 585
R17010 GND.n2861 GND.n1472 585
R17011 GND.n2862 GND.n2861 585
R17012 GND.n8196 GND.n1471 585
R17013 GND.n3004 GND.n1471 585
R17014 GND.n8197 GND.n1470 585
R17015 GND.n2875 GND.n1470 585
R17016 GND.n8198 GND.n1469 585
R17017 GND.n2994 GND.n1469 585
R17018 GND.n2872 GND.n1467 585
R17019 GND.n2873 GND.n2872 585
R17020 GND.n8202 GND.n1466 585
R17021 GND.n2978 GND.n1466 585
R17022 GND.n8203 GND.n1465 585
R17023 GND.n2884 GND.n1465 585
R17024 GND.n8204 GND.n1464 585
R17025 GND.n2970 GND.n1464 585
R17026 GND.n2891 GND.n1462 585
R17027 GND.n2892 GND.n2891 585
R17028 GND.n8208 GND.n1461 585
R17029 GND.n2961 GND.n1461 585
R17030 GND.n8209 GND.n1460 585
R17031 GND.n2904 GND.n1460 585
R17032 GND.n8210 GND.n1459 585
R17033 GND.n2953 GND.n1459 585
R17034 GND.n2911 GND.n1457 585
R17035 GND.n2912 GND.n2911 585
R17036 GND.n8214 GND.n1456 585
R17037 GND.n2944 GND.n1456 585
R17038 GND.n8215 GND.n1455 585
R17039 GND.n2924 GND.n1455 585
R17040 GND.n8216 GND.n1454 585
R17041 GND.n1454 GND.n1358 585
R17042 GND.n8023 GND.n1706 585
R17043 GND.n3872 GND.n3854 585
R17044 GND.n3871 GND.n3870 585
R17045 GND.n3869 GND.n3868 585
R17046 GND.n3867 GND.n3866 585
R17047 GND.n3865 GND.n3864 585
R17048 GND.n3863 GND.n3862 585
R17049 GND.n3861 GND.n3860 585
R17050 GND.n3859 GND.n3858 585
R17051 GND.n3857 GND.n3856 585
R17052 GND.n3855 GND.n1681 585
R17053 GND.n8024 GND.n8023 585
R17054 GND.n7248 GND.n4731 526.135
R17055 GND.n4775 GND.n4774 526.135
R17056 GND.n2181 GND.n2180 526.135
R17057 GND.n7970 GND.n1908 526.135
R17058 GND.n7972 GND.n7971 256.663
R17059 GND.n7972 GND.n1877 256.663
R17060 GND.n7972 GND.n1878 256.663
R17061 GND.n7972 GND.n1879 256.663
R17062 GND.n7972 GND.n1880 256.663
R17063 GND.n7972 GND.n1881 256.663
R17064 GND.n7972 GND.n1882 256.663
R17065 GND.n7972 GND.n1883 256.663
R17066 GND.n7972 GND.n1884 256.663
R17067 GND.n7972 GND.n1885 256.663
R17068 GND.n7972 GND.n1886 256.663
R17069 GND.n7972 GND.n1887 256.663
R17070 GND.n7972 GND.n1888 256.663
R17071 GND.n7973 GND.n7972 256.663
R17072 GND.n7972 GND.n1889 256.663
R17073 GND.n7976 GND.n1872 256.663
R17074 GND.n7972 GND.n1890 256.663
R17075 GND.n7972 GND.n1891 256.663
R17076 GND.n7972 GND.n1892 256.663
R17077 GND.n7972 GND.n1893 256.663
R17078 GND.n7972 GND.n1894 256.663
R17079 GND.n7972 GND.n1895 256.663
R17080 GND.n7972 GND.n1896 256.663
R17081 GND.n7972 GND.n1897 256.663
R17082 GND.n7972 GND.n1898 256.663
R17083 GND.n7972 GND.n1899 256.663
R17084 GND.n7972 GND.n1900 256.663
R17085 GND.n7972 GND.n1901 256.663
R17086 GND.n7972 GND.n1902 256.663
R17087 GND.n7972 GND.n1903 256.663
R17088 GND.n7972 GND.n1904 256.663
R17089 GND.n7249 GND.n4701 256.663
R17090 GND.n7249 GND.n4702 256.663
R17091 GND.n7249 GND.n4703 256.663
R17092 GND.n7249 GND.n4704 256.663
R17093 GND.n7249 GND.n4705 256.663
R17094 GND.n7249 GND.n4706 256.663
R17095 GND.n7249 GND.n4707 256.663
R17096 GND.n7249 GND.n4708 256.663
R17097 GND.n7249 GND.n4709 256.663
R17098 GND.n7249 GND.n4710 256.663
R17099 GND.n7249 GND.n4711 256.663
R17100 GND.n7249 GND.n4712 256.663
R17101 GND.n7249 GND.n4713 256.663
R17102 GND.n7249 GND.n4714 256.663
R17103 GND.n7249 GND.n4715 256.663
R17104 GND.n7189 GND.n7188 256.663
R17105 GND.n7249 GND.n4716 256.663
R17106 GND.n7249 GND.n4717 256.663
R17107 GND.n7249 GND.n4718 256.663
R17108 GND.n7249 GND.n4719 256.663
R17109 GND.n7249 GND.n4720 256.663
R17110 GND.n7249 GND.n4721 256.663
R17111 GND.n7249 GND.n4722 256.663
R17112 GND.n7249 GND.n4723 256.663
R17113 GND.n7249 GND.n4724 256.663
R17114 GND.n7249 GND.n4725 256.663
R17115 GND.n7249 GND.n4726 256.663
R17116 GND.n7249 GND.n4727 256.663
R17117 GND.n7249 GND.n4728 256.663
R17118 GND.n7249 GND.n4729 256.663
R17119 GND.n7249 GND.n4730 256.663
R17120 GND.n3876 GND.t40 255.518
R17121 GND.n6342 GND.t151 255.518
R17122 GND.n7183 GND.n4875 242.672
R17123 GND.n7183 GND.n4874 242.672
R17124 GND.n7183 GND.n4873 242.672
R17125 GND.n7183 GND.n4872 242.672
R17126 GND.n7183 GND.n4871 242.672
R17127 GND.n7183 GND.n4870 242.672
R17128 GND.n10075 GND.n10074 242.672
R17129 GND.n10074 GND.n10073 242.672
R17130 GND.n10074 GND.n10043 242.672
R17131 GND.n10074 GND.n10042 242.672
R17132 GND.n10074 GND.n10041 242.672
R17133 GND.n10074 GND.n10040 242.672
R17134 GND.n7759 GND.n7758 242.672
R17135 GND.n7759 GND.n2328 242.672
R17136 GND.n7759 GND.n2329 242.672
R17137 GND.n7759 GND.n2330 242.672
R17138 GND.n7759 GND.n2331 242.672
R17139 GND.n7759 GND.n2332 242.672
R17140 GND.n7759 GND.n2333 242.672
R17141 GND.n7759 GND.n2334 242.672
R17142 GND.n7759 GND.n2335 242.672
R17143 GND.n7759 GND.n2336 242.672
R17144 GND.n7759 GND.n2337 242.672
R17145 GND.n7759 GND.n2338 242.672
R17146 GND.n7759 GND.n2339 242.672
R17147 GND.n7409 GND.n7408 242.672
R17148 GND.n7408 GND.n4435 242.672
R17149 GND.n7408 GND.n4434 242.672
R17150 GND.n7408 GND.n4433 242.672
R17151 GND.n7408 GND.n4432 242.672
R17152 GND.n7408 GND.n4431 242.672
R17153 GND.n7408 GND.n4430 242.672
R17154 GND.n7408 GND.n4429 242.672
R17155 GND.n7408 GND.n4428 242.672
R17156 GND.n7408 GND.n4427 242.672
R17157 GND.n7408 GND.n4426 242.672
R17158 GND.n7408 GND.n4425 242.672
R17159 GND.n7408 GND.n4424 242.672
R17160 GND.n7408 GND.n4423 242.672
R17161 GND.n8362 GND.n8361 242.672
R17162 GND.n8362 GND.n1322 242.672
R17163 GND.n8362 GND.n1323 242.672
R17164 GND.n8362 GND.n1324 242.672
R17165 GND.n8362 GND.n1325 242.672
R17166 GND.n8362 GND.n1326 242.672
R17167 GND.n8362 GND.n1327 242.672
R17168 GND.n8362 GND.n1328 242.672
R17169 GND.n8362 GND.n1329 242.672
R17170 GND.n8362 GND.n1330 242.672
R17171 GND.n8362 GND.n1331 242.672
R17172 GND.n8362 GND.n1332 242.672
R17173 GND.n8362 GND.n1333 242.672
R17174 GND.n8362 GND.n1334 242.672
R17175 GND.n8362 GND.n1335 242.672
R17176 GND.n8362 GND.n1336 242.672
R17177 GND.n8362 GND.n1337 242.672
R17178 GND.n8362 GND.n1338 242.672
R17179 GND.n8362 GND.n1339 242.672
R17180 GND.n8362 GND.n1340 242.672
R17181 GND.n8362 GND.n1341 242.672
R17182 GND.n8362 GND.n1342 242.672
R17183 GND.n8362 GND.n1343 242.672
R17184 GND.n8362 GND.n1344 242.672
R17185 GND.n8362 GND.n1345 242.672
R17186 GND.n8362 GND.n1346 242.672
R17187 GND.n8362 GND.n1347 242.672
R17188 GND.n8362 GND.n1348 242.672
R17189 GND.n8362 GND.n1349 242.672
R17190 GND.n8362 GND.n1350 242.672
R17191 GND.n8023 GND.n1700 242.672
R17192 GND.n8023 GND.n1699 242.672
R17193 GND.n8023 GND.n1698 242.672
R17194 GND.n8023 GND.n1697 242.672
R17195 GND.n8023 GND.n1696 242.672
R17196 GND.n8023 GND.n1695 242.672
R17197 GND.n8023 GND.n1694 242.672
R17198 GND.n8023 GND.n1693 242.672
R17199 GND.n8023 GND.n1692 242.672
R17200 GND.n8023 GND.n1691 242.672
R17201 GND.n8023 GND.n1690 242.672
R17202 GND.n8023 GND.n1689 242.672
R17203 GND.n8023 GND.n1688 242.672
R17204 GND.n8023 GND.n1687 242.672
R17205 GND.n8023 GND.n1686 242.672
R17206 GND.n8023 GND.n1685 242.672
R17207 GND.n7977 GND.n1870 242.672
R17208 GND.n8023 GND.n1708 242.672
R17209 GND.n8023 GND.n1709 242.672
R17210 GND.n8023 GND.n1710 242.672
R17211 GND.n8023 GND.n1711 242.672
R17212 GND.n8023 GND.n1712 242.672
R17213 GND.n8023 GND.n1713 242.672
R17214 GND.n8023 GND.n1714 242.672
R17215 GND.n8023 GND.n1715 242.672
R17216 GND.n8023 GND.n1716 242.672
R17217 GND.n8023 GND.n1717 242.672
R17218 GND.n8023 GND.n1718 242.672
R17219 GND.n8023 GND.n1719 242.672
R17220 GND.n8023 GND.n1720 242.672
R17221 GND.n8023 GND.n1721 242.672
R17222 GND.n7183 GND.n7182 242.672
R17223 GND.n7183 GND.n4840 242.672
R17224 GND.n7183 GND.n4841 242.672
R17225 GND.n7183 GND.n4842 242.672
R17226 GND.n7183 GND.n4843 242.672
R17227 GND.n7183 GND.n4844 242.672
R17228 GND.n7183 GND.n4845 242.672
R17229 GND.n7183 GND.n4846 242.672
R17230 GND.n7183 GND.n4847 242.672
R17231 GND.n7183 GND.n4848 242.672
R17232 GND.n7183 GND.n4849 242.672
R17233 GND.n7183 GND.n4850 242.672
R17234 GND.n7183 GND.n4851 242.672
R17235 GND.n7183 GND.n4852 242.672
R17236 GND.n7187 GND.n4834 242.672
R17237 GND.n7184 GND.n7183 242.672
R17238 GND.n7183 GND.n4853 242.672
R17239 GND.n7183 GND.n4854 242.672
R17240 GND.n7183 GND.n4855 242.672
R17241 GND.n7183 GND.n4856 242.672
R17242 GND.n7183 GND.n4857 242.672
R17243 GND.n7183 GND.n4858 242.672
R17244 GND.n7183 GND.n4859 242.672
R17245 GND.n7183 GND.n4860 242.672
R17246 GND.n7183 GND.n4861 242.672
R17247 GND.n7183 GND.n4862 242.672
R17248 GND.n7183 GND.n4863 242.672
R17249 GND.n7183 GND.n4864 242.672
R17250 GND.n7183 GND.n4865 242.672
R17251 GND.n7183 GND.n4866 242.672
R17252 GND.n7183 GND.n4867 242.672
R17253 GND.n10074 GND.n10039 242.672
R17254 GND.n10074 GND.n9841 242.672
R17255 GND.n10074 GND.n9840 242.672
R17256 GND.n10074 GND.n9839 242.672
R17257 GND.n10074 GND.n9838 242.672
R17258 GND.n10074 GND.n9837 242.672
R17259 GND.n10074 GND.n9836 242.672
R17260 GND.n10074 GND.n9835 242.672
R17261 GND.n10074 GND.n9834 242.672
R17262 GND.n10074 GND.n9833 242.672
R17263 GND.n10074 GND.n9832 242.672
R17264 GND.n10074 GND.n9831 242.672
R17265 GND.n10074 GND.n9830 242.672
R17266 GND.n10074 GND.n9829 242.672
R17267 GND.n10074 GND.n9828 242.672
R17268 GND.n10074 GND.n9827 242.672
R17269 GND.n10074 GND.n9826 242.672
R17270 GND.n10074 GND.n9825 242.672
R17271 GND.n10074 GND.n9824 242.672
R17272 GND.n10074 GND.n9823 242.672
R17273 GND.n10074 GND.n9822 242.672
R17274 GND.n10074 GND.n9821 242.672
R17275 GND.n10074 GND.n9820 242.672
R17276 GND.n10074 GND.n9819 242.672
R17277 GND.n10074 GND.n9818 242.672
R17278 GND.n10074 GND.n9817 242.672
R17279 GND.n10074 GND.n9816 242.672
R17280 GND.n10074 GND.n9815 242.672
R17281 GND.n10074 GND.n9814 242.672
R17282 GND.n10074 GND.n9813 242.672
R17283 GND.n10074 GND.n9812 242.672
R17284 GND.n8362 GND.n1352 242.672
R17285 GND.n8362 GND.n1353 242.672
R17286 GND.n8362 GND.n1354 242.672
R17287 GND.n8362 GND.n1355 242.672
R17288 GND.n8362 GND.n1356 242.672
R17289 GND.n8023 GND.n1705 242.672
R17290 GND.n8023 GND.n1704 242.672
R17291 GND.n8023 GND.n1703 242.672
R17292 GND.n8023 GND.n1702 242.672
R17293 GND.n8023 GND.n1701 242.672
R17294 GND.n1917 GND.n1915 240.849
R17295 GND.n4749 GND.n4747 240.849
R17296 GND.n9889 GND.n9888 240.244
R17297 GND.n9892 GND.n9891 240.244
R17298 GND.n9899 GND.n9898 240.244
R17299 GND.n9902 GND.n9901 240.244
R17300 GND.n9907 GND.n9879 240.244
R17301 GND.n9911 GND.n9910 240.244
R17302 GND.n9918 GND.n9917 240.244
R17303 GND.n9921 GND.n9920 240.244
R17304 GND.n9928 GND.n9927 240.244
R17305 GND.n9931 GND.n9930 240.244
R17306 GND.n9938 GND.n9937 240.244
R17307 GND.n9942 GND.n9941 240.244
R17308 GND.n9949 GND.n9948 240.244
R17309 GND.n9952 GND.n9951 240.244
R17310 GND.n9959 GND.n9958 240.244
R17311 GND.n9962 GND.n9961 240.244
R17312 GND.n9969 GND.n9968 240.244
R17313 GND.n9862 GND.n9861 240.244
R17314 GND.n9977 GND.n9976 240.244
R17315 GND.n9980 GND.n9979 240.244
R17316 GND.n9987 GND.n9986 240.244
R17317 GND.n9990 GND.n9989 240.244
R17318 GND.n9997 GND.n9996 240.244
R17319 GND.n10003 GND.n10002 240.244
R17320 GND.n10010 GND.n10009 240.244
R17321 GND.n10013 GND.n10012 240.244
R17322 GND.n10020 GND.n10019 240.244
R17323 GND.n10023 GND.n10022 240.244
R17324 GND.n10030 GND.n10029 240.244
R17325 GND.n10032 GND.n9842 240.244
R17326 GND.n6415 GND.n4883 240.244
R17327 GND.n7085 GND.n4883 240.244
R17328 GND.n7085 GND.n4894 240.244
R17329 GND.n5352 GND.n4894 240.244
R17330 GND.n5352 GND.n4907 240.244
R17331 GND.n6474 GND.n4907 240.244
R17332 GND.n6474 GND.n4924 240.244
R17333 GND.n6478 GND.n4924 240.244
R17334 GND.n6478 GND.n4936 240.244
R17335 GND.n6488 GND.n4936 240.244
R17336 GND.n6488 GND.n4947 240.244
R17337 GND.n6492 GND.n4947 240.244
R17338 GND.n6492 GND.n4957 240.244
R17339 GND.n6502 GND.n4957 240.244
R17340 GND.n6502 GND.n4968 240.244
R17341 GND.n6506 GND.n4968 240.244
R17342 GND.n6506 GND.n4978 240.244
R17343 GND.n6517 GND.n4978 240.244
R17344 GND.n6517 GND.n4989 240.244
R17345 GND.n5330 GND.n4989 240.244
R17346 GND.n5330 GND.n4998 240.244
R17347 GND.n6668 GND.n4998 240.244
R17348 GND.n6668 GND.n5009 240.244
R17349 GND.n6664 GND.n5009 240.244
R17350 GND.n6664 GND.n5019 240.244
R17351 GND.n6656 GND.n5019 240.244
R17352 GND.n6656 GND.n5030 240.244
R17353 GND.n6652 GND.n5030 240.244
R17354 GND.n6652 GND.n5040 240.244
R17355 GND.n6644 GND.n5040 240.244
R17356 GND.n6644 GND.n5051 240.244
R17357 GND.n6640 GND.n5051 240.244
R17358 GND.n6640 GND.n5061 240.244
R17359 GND.n6632 GND.n5061 240.244
R17360 GND.n6632 GND.n5072 240.244
R17361 GND.n6628 GND.n5072 240.244
R17362 GND.n6628 GND.n5082 240.244
R17363 GND.n6620 GND.n5082 240.244
R17364 GND.n6620 GND.n5093 240.244
R17365 GND.n6616 GND.n5093 240.244
R17366 GND.n6616 GND.n5103 240.244
R17367 GND.n6608 GND.n5103 240.244
R17368 GND.n6608 GND.n5114 240.244
R17369 GND.n6604 GND.n5114 240.244
R17370 GND.n6604 GND.n5124 240.244
R17371 GND.n6596 GND.n5124 240.244
R17372 GND.n6596 GND.n5135 240.244
R17373 GND.n6592 GND.n5135 240.244
R17374 GND.n6592 GND.n5145 240.244
R17375 GND.n6584 GND.n5145 240.244
R17376 GND.n6584 GND.n5156 240.244
R17377 GND.n6580 GND.n5156 240.244
R17378 GND.n6580 GND.n5166 240.244
R17379 GND.n5291 GND.n5166 240.244
R17380 GND.n5291 GND.n5175 240.244
R17381 GND.n6770 GND.n5175 240.244
R17382 GND.n6770 GND.n5185 240.244
R17383 GND.n5190 GND.n5185 240.244
R17384 GND.n6777 GND.n5190 240.244
R17385 GND.n6778 GND.n6777 240.244
R17386 GND.n6778 GND.n109 240.244
R17387 GND.n6786 GND.n109 240.244
R17388 GND.n6786 GND.n5281 240.244
R17389 GND.n5281 GND.n5270 240.244
R17390 GND.n5270 GND.n128 240.244
R17391 GND.n6894 GND.n128 240.244
R17392 GND.n6894 GND.n140 240.244
R17393 GND.n6890 GND.n140 240.244
R17394 GND.n6890 GND.n150 240.244
R17395 GND.n6882 GND.n150 240.244
R17396 GND.n6882 GND.n160 240.244
R17397 GND.n6878 GND.n160 240.244
R17398 GND.n6878 GND.n171 240.244
R17399 GND.n6870 GND.n171 240.244
R17400 GND.n6870 GND.n181 240.244
R17401 GND.n6866 GND.n181 240.244
R17402 GND.n6866 GND.n192 240.244
R17403 GND.n6858 GND.n192 240.244
R17404 GND.n6858 GND.n202 240.244
R17405 GND.n6854 GND.n202 240.244
R17406 GND.n6854 GND.n213 240.244
R17407 GND.n6846 GND.n213 240.244
R17408 GND.n6846 GND.n223 240.244
R17409 GND.n6842 GND.n223 240.244
R17410 GND.n6842 GND.n234 240.244
R17411 GND.n6834 GND.n234 240.244
R17412 GND.n6834 GND.n244 240.244
R17413 GND.n441 GND.n244 240.244
R17414 GND.n441 GND.n254 240.244
R17415 GND.n9736 GND.n254 240.244
R17416 GND.n9736 GND.n264 240.244
R17417 GND.n9741 GND.n264 240.244
R17418 GND.n9741 GND.n275 240.244
R17419 GND.n9751 GND.n275 240.244
R17420 GND.n9751 GND.n285 240.244
R17421 GND.n9756 GND.n285 240.244
R17422 GND.n9756 GND.n296 240.244
R17423 GND.n9766 GND.n296 240.244
R17424 GND.n9766 GND.n306 240.244
R17425 GND.n9771 GND.n306 240.244
R17426 GND.n9771 GND.n317 240.244
R17427 GND.n9781 GND.n317 240.244
R17428 GND.n9781 GND.n327 240.244
R17429 GND.n9786 GND.n327 240.244
R17430 GND.n9786 GND.n338 240.244
R17431 GND.n10105 GND.n338 240.244
R17432 GND.n10105 GND.n348 240.244
R17433 GND.n10109 GND.n348 240.244
R17434 GND.n10109 GND.n359 240.244
R17435 GND.n10112 GND.n359 240.244
R17436 GND.n10112 GND.n368 240.244
R17437 GND.n10116 GND.n368 240.244
R17438 GND.n10116 GND.n378 240.244
R17439 GND.n10119 GND.n378 240.244
R17440 GND.n10119 GND.n387 240.244
R17441 GND.n10123 GND.n387 240.244
R17442 GND.n10123 GND.n397 240.244
R17443 GND.n10126 GND.n397 240.244
R17444 GND.n10126 GND.n406 240.244
R17445 GND.n10129 GND.n406 240.244
R17446 GND.n10129 GND.n415 240.244
R17447 GND.n4877 GND.n4876 240.244
R17448 GND.n7176 GND.n4876 240.244
R17449 GND.n7174 GND.n7173 240.244
R17450 GND.n7170 GND.n7169 240.244
R17451 GND.n7166 GND.n7165 240.244
R17452 GND.n7161 GND.n7106 240.244
R17453 GND.n7159 GND.n7158 240.244
R17454 GND.n7155 GND.n7154 240.244
R17455 GND.n7151 GND.n7150 240.244
R17456 GND.n7147 GND.n7146 240.244
R17457 GND.n7143 GND.n7142 240.244
R17458 GND.n7139 GND.n7138 240.244
R17459 GND.n7135 GND.n7134 240.244
R17460 GND.n7131 GND.n7130 240.244
R17461 GND.n7185 GND.n4838 240.244
R17462 GND.n5386 GND.n5385 240.244
R17463 GND.n5381 GND.n5380 240.244
R17464 GND.n5396 GND.n5395 240.244
R17465 GND.n5402 GND.n5401 240.244
R17466 GND.n5406 GND.n5405 240.244
R17467 GND.n5412 GND.n5411 240.244
R17468 GND.n5416 GND.n5415 240.244
R17469 GND.n5422 GND.n5421 240.244
R17470 GND.n5429 GND.n5428 240.244
R17471 GND.n5435 GND.n5434 240.244
R17472 GND.n5439 GND.n5438 240.244
R17473 GND.n5445 GND.n5444 240.244
R17474 GND.n5449 GND.n5448 240.244
R17475 GND.n5455 GND.n5454 240.244
R17476 GND.n5457 GND.n4868 240.244
R17477 GND.n7092 GND.n4878 240.244
R17478 GND.n7092 GND.n4881 240.244
R17479 GND.n4915 GND.n4881 240.244
R17480 GND.n4915 GND.n4911 240.244
R17481 GND.n7075 GND.n4911 240.244
R17482 GND.n7075 GND.n4912 240.244
R17483 GND.n7071 GND.n4912 240.244
R17484 GND.n7071 GND.n4923 240.244
R17485 GND.n7063 GND.n4923 240.244
R17486 GND.n7063 GND.n4939 240.244
R17487 GND.n7059 GND.n4939 240.244
R17488 GND.n7059 GND.n4945 240.244
R17489 GND.n7051 GND.n4945 240.244
R17490 GND.n7051 GND.n4960 240.244
R17491 GND.n7047 GND.n4960 240.244
R17492 GND.n7047 GND.n4966 240.244
R17493 GND.n7039 GND.n4966 240.244
R17494 GND.n7039 GND.n4981 240.244
R17495 GND.n7035 GND.n4981 240.244
R17496 GND.n7035 GND.n4987 240.244
R17497 GND.n7027 GND.n4987 240.244
R17498 GND.n7027 GND.n5001 240.244
R17499 GND.n7023 GND.n5001 240.244
R17500 GND.n7023 GND.n5007 240.244
R17501 GND.n7015 GND.n5007 240.244
R17502 GND.n7015 GND.n5022 240.244
R17503 GND.n7011 GND.n5022 240.244
R17504 GND.n7011 GND.n5028 240.244
R17505 GND.n7003 GND.n5028 240.244
R17506 GND.n7003 GND.n5043 240.244
R17507 GND.n6999 GND.n5043 240.244
R17508 GND.n6999 GND.n5049 240.244
R17509 GND.n6991 GND.n5049 240.244
R17510 GND.n6991 GND.n5064 240.244
R17511 GND.n6987 GND.n5064 240.244
R17512 GND.n6987 GND.n5070 240.244
R17513 GND.n6979 GND.n5070 240.244
R17514 GND.n6979 GND.n5085 240.244
R17515 GND.n6975 GND.n5085 240.244
R17516 GND.n6975 GND.n5091 240.244
R17517 GND.n6967 GND.n5091 240.244
R17518 GND.n6967 GND.n5106 240.244
R17519 GND.n6963 GND.n5106 240.244
R17520 GND.n6963 GND.n5112 240.244
R17521 GND.n6955 GND.n5112 240.244
R17522 GND.n6955 GND.n5127 240.244
R17523 GND.n6951 GND.n5127 240.244
R17524 GND.n6951 GND.n5133 240.244
R17525 GND.n6943 GND.n5133 240.244
R17526 GND.n6943 GND.n5148 240.244
R17527 GND.n6939 GND.n5148 240.244
R17528 GND.n6939 GND.n5154 240.244
R17529 GND.n6931 GND.n5154 240.244
R17530 GND.n6931 GND.n5169 240.244
R17531 GND.n6927 GND.n5169 240.244
R17532 GND.n6927 GND.n5174 240.244
R17533 GND.n6919 GND.n5174 240.244
R17534 GND.n6919 GND.n6917 240.244
R17535 GND.n6917 GND.n5189 240.244
R17536 GND.n5189 GND.n112 240.244
R17537 GND.n10309 GND.n112 240.244
R17538 GND.n10309 GND.n113 240.244
R17539 GND.n5268 GND.n113 240.244
R17540 GND.n5268 GND.n125 240.244
R17541 GND.n10304 GND.n125 240.244
R17542 GND.n10304 GND.n126 240.244
R17543 GND.n10296 GND.n126 240.244
R17544 GND.n10296 GND.n143 240.244
R17545 GND.n10292 GND.n143 240.244
R17546 GND.n10292 GND.n148 240.244
R17547 GND.n10284 GND.n148 240.244
R17548 GND.n10284 GND.n163 240.244
R17549 GND.n10280 GND.n163 240.244
R17550 GND.n10280 GND.n169 240.244
R17551 GND.n10272 GND.n169 240.244
R17552 GND.n10272 GND.n184 240.244
R17553 GND.n10268 GND.n184 240.244
R17554 GND.n10268 GND.n190 240.244
R17555 GND.n10260 GND.n190 240.244
R17556 GND.n10260 GND.n205 240.244
R17557 GND.n10256 GND.n205 240.244
R17558 GND.n10256 GND.n211 240.244
R17559 GND.n10248 GND.n211 240.244
R17560 GND.n10248 GND.n226 240.244
R17561 GND.n10244 GND.n226 240.244
R17562 GND.n10244 GND.n232 240.244
R17563 GND.n10236 GND.n232 240.244
R17564 GND.n10236 GND.n247 240.244
R17565 GND.n10232 GND.n247 240.244
R17566 GND.n10232 GND.n253 240.244
R17567 GND.n10224 GND.n253 240.244
R17568 GND.n10224 GND.n267 240.244
R17569 GND.n10220 GND.n267 240.244
R17570 GND.n10220 GND.n273 240.244
R17571 GND.n10212 GND.n273 240.244
R17572 GND.n10212 GND.n288 240.244
R17573 GND.n10208 GND.n288 240.244
R17574 GND.n10208 GND.n294 240.244
R17575 GND.n10200 GND.n294 240.244
R17576 GND.n10200 GND.n309 240.244
R17577 GND.n10196 GND.n309 240.244
R17578 GND.n10196 GND.n315 240.244
R17579 GND.n10188 GND.n315 240.244
R17580 GND.n10188 GND.n330 240.244
R17581 GND.n10184 GND.n330 240.244
R17582 GND.n10184 GND.n336 240.244
R17583 GND.n10176 GND.n336 240.244
R17584 GND.n10176 GND.n351 240.244
R17585 GND.n10172 GND.n351 240.244
R17586 GND.n10172 GND.n357 240.244
R17587 GND.n10164 GND.n357 240.244
R17588 GND.n10164 GND.n371 240.244
R17589 GND.n10160 GND.n371 240.244
R17590 GND.n10160 GND.n377 240.244
R17591 GND.n10152 GND.n377 240.244
R17592 GND.n10152 GND.n390 240.244
R17593 GND.n10148 GND.n390 240.244
R17594 GND.n10148 GND.n396 240.244
R17595 GND.n10140 GND.n396 240.244
R17596 GND.n10140 GND.n409 240.244
R17597 GND.n10136 GND.n409 240.244
R17598 GND.n8022 GND.n1722 240.244
R17599 GND.n1727 GND.n1726 240.244
R17600 GND.n1729 GND.n1728 240.244
R17601 GND.n1733 GND.n1732 240.244
R17602 GND.n1735 GND.n1734 240.244
R17603 GND.n1741 GND.n1740 240.244
R17604 GND.n1743 GND.n1742 240.244
R17605 GND.n1747 GND.n1746 240.244
R17606 GND.n1749 GND.n1748 240.244
R17607 GND.n1753 GND.n1752 240.244
R17608 GND.n1755 GND.n1754 240.244
R17609 GND.n1761 GND.n1758 240.244
R17610 GND.n1763 GND.n1762 240.244
R17611 GND.n7978 GND.n1766 240.244
R17612 GND.n1767 GND.n1684 240.244
R17613 GND.n1771 GND.n1770 240.244
R17614 GND.n1773 GND.n1772 240.244
R17615 GND.n1779 GND.n1778 240.244
R17616 GND.n1781 GND.n1780 240.244
R17617 GND.n1785 GND.n1784 240.244
R17618 GND.n1787 GND.n1786 240.244
R17619 GND.n1791 GND.n1790 240.244
R17620 GND.n1793 GND.n1792 240.244
R17621 GND.n1799 GND.n1796 240.244
R17622 GND.n1801 GND.n1800 240.244
R17623 GND.n1805 GND.n1804 240.244
R17624 GND.n1807 GND.n1806 240.244
R17625 GND.n1811 GND.n1810 240.244
R17626 GND.n1813 GND.n1812 240.244
R17627 GND.n1819 GND.n1816 240.244
R17628 GND.n2929 GND.n2923 240.244
R17629 GND.n2945 GND.n2923 240.244
R17630 GND.n2946 GND.n2945 240.244
R17631 GND.n2946 GND.n2913 240.244
R17632 GND.n2913 GND.n2903 240.244
R17633 GND.n2962 GND.n2903 240.244
R17634 GND.n2963 GND.n2962 240.244
R17635 GND.n2963 GND.n2893 240.244
R17636 GND.n2893 GND.n2883 240.244
R17637 GND.n2979 GND.n2883 240.244
R17638 GND.n2980 GND.n2979 240.244
R17639 GND.n2980 GND.n2874 240.244
R17640 GND.n2982 GND.n2874 240.244
R17641 GND.n2982 GND.n2864 240.244
R17642 GND.n2864 GND.n2860 240.244
R17643 GND.n3019 GND.n2860 240.244
R17644 GND.n3019 GND.n2849 240.244
R17645 GND.n3021 GND.n2849 240.244
R17646 GND.n3021 GND.n2833 240.244
R17647 GND.n3046 GND.n2833 240.244
R17648 GND.n3046 GND.n2824 240.244
R17649 GND.n3048 GND.n2824 240.244
R17650 GND.n3048 GND.n2814 240.244
R17651 GND.n2814 GND.n2805 240.244
R17652 GND.n3083 GND.n2805 240.244
R17653 GND.n3083 GND.n2796 240.244
R17654 GND.n3085 GND.n2796 240.244
R17655 GND.n3085 GND.n2786 240.244
R17656 GND.n2786 GND.n2776 240.244
R17657 GND.n3120 GND.n2776 240.244
R17658 GND.n3120 GND.n2766 240.244
R17659 GND.n3123 GND.n2766 240.244
R17660 GND.n3123 GND.n2756 240.244
R17661 GND.n2756 GND.n2748 240.244
R17662 GND.n3159 GND.n2748 240.244
R17663 GND.n3159 GND.n2739 240.244
R17664 GND.n3161 GND.n2739 240.244
R17665 GND.n3161 GND.n2729 240.244
R17666 GND.n2729 GND.n2719 240.244
R17667 GND.n3196 GND.n2719 240.244
R17668 GND.n3196 GND.n2710 240.244
R17669 GND.n3198 GND.n2710 240.244
R17670 GND.n3198 GND.n2699 240.244
R17671 GND.n2699 GND.n2690 240.244
R17672 GND.n3233 GND.n2690 240.244
R17673 GND.n3233 GND.n2681 240.244
R17674 GND.n3235 GND.n2681 240.244
R17675 GND.n3235 GND.n2671 240.244
R17676 GND.n2671 GND.n2661 240.244
R17677 GND.n3270 GND.n2661 240.244
R17678 GND.n3270 GND.n2651 240.244
R17679 GND.n3272 GND.n2651 240.244
R17680 GND.n3272 GND.n2641 240.244
R17681 GND.n2641 GND.n2632 240.244
R17682 GND.n3309 GND.n2632 240.244
R17683 GND.n3309 GND.n2623 240.244
R17684 GND.n3311 GND.n2623 240.244
R17685 GND.n3311 GND.n2617 240.244
R17686 GND.n2617 GND.n2616 240.244
R17687 GND.n2616 GND.n2605 240.244
R17688 GND.n2605 GND.n1534 240.244
R17689 GND.n2597 GND.n1534 240.244
R17690 GND.n3557 GND.n2597 240.244
R17691 GND.n3558 GND.n3557 240.244
R17692 GND.n3558 GND.n1553 240.244
R17693 GND.n1563 GND.n1553 240.244
R17694 GND.n1564 GND.n1563 240.244
R17695 GND.n2584 GND.n1564 240.244
R17696 GND.n2584 GND.n1570 240.244
R17697 GND.n1571 GND.n1570 240.244
R17698 GND.n1572 GND.n1571 240.244
R17699 GND.n2566 GND.n1572 240.244
R17700 GND.n2566 GND.n1578 240.244
R17701 GND.n1579 GND.n1578 240.244
R17702 GND.n1580 GND.n1579 240.244
R17703 GND.n2554 GND.n1580 240.244
R17704 GND.n2554 GND.n1586 240.244
R17705 GND.n1587 GND.n1586 240.244
R17706 GND.n1588 GND.n1587 240.244
R17707 GND.n2530 GND.n1588 240.244
R17708 GND.n2530 GND.n1594 240.244
R17709 GND.n1595 GND.n1594 240.244
R17710 GND.n1596 GND.n1595 240.244
R17711 GND.n3649 GND.n1596 240.244
R17712 GND.n3649 GND.n1602 240.244
R17713 GND.n1603 GND.n1602 240.244
R17714 GND.n1604 GND.n1603 240.244
R17715 GND.n2497 GND.n1604 240.244
R17716 GND.n2497 GND.n1610 240.244
R17717 GND.n1611 GND.n1610 240.244
R17718 GND.n1612 GND.n1611 240.244
R17719 GND.n2479 GND.n1612 240.244
R17720 GND.n2479 GND.n1618 240.244
R17721 GND.n1619 GND.n1618 240.244
R17722 GND.n1620 GND.n1619 240.244
R17723 GND.n2467 GND.n1620 240.244
R17724 GND.n2467 GND.n1626 240.244
R17725 GND.n1627 GND.n1626 240.244
R17726 GND.n1628 GND.n1627 240.244
R17727 GND.n2445 GND.n1628 240.244
R17728 GND.n2445 GND.n1634 240.244
R17729 GND.n1635 GND.n1634 240.244
R17730 GND.n1636 GND.n1635 240.244
R17731 GND.n3752 GND.n1636 240.244
R17732 GND.n3752 GND.n1642 240.244
R17733 GND.n1643 GND.n1642 240.244
R17734 GND.n1644 GND.n1643 240.244
R17735 GND.n2412 GND.n1644 240.244
R17736 GND.n2412 GND.n1650 240.244
R17737 GND.n1651 GND.n1650 240.244
R17738 GND.n1652 GND.n1651 240.244
R17739 GND.n2394 GND.n1652 240.244
R17740 GND.n2394 GND.n1658 240.244
R17741 GND.n1659 GND.n1658 240.244
R17742 GND.n1660 GND.n1659 240.244
R17743 GND.n2382 GND.n1660 240.244
R17744 GND.n2382 GND.n1666 240.244
R17745 GND.n1667 GND.n1666 240.244
R17746 GND.n1668 GND.n1667 240.244
R17747 GND.n1674 GND.n1668 240.244
R17748 GND.n8027 GND.n1674 240.244
R17749 GND.n1361 GND.n1360 240.244
R17750 GND.n8355 GND.n1360 240.244
R17751 GND.n8353 GND.n8352 240.244
R17752 GND.n8349 GND.n8348 240.244
R17753 GND.n8345 GND.n8344 240.244
R17754 GND.n8340 GND.n1373 240.244
R17755 GND.n8338 GND.n8337 240.244
R17756 GND.n8334 GND.n8333 240.244
R17757 GND.n8330 GND.n8329 240.244
R17758 GND.n8326 GND.n8325 240.244
R17759 GND.n8322 GND.n8321 240.244
R17760 GND.n8318 GND.n8317 240.244
R17761 GND.n8314 GND.n8313 240.244
R17762 GND.n8310 GND.n8309 240.244
R17763 GND.n8306 GND.n8305 240.244
R17764 GND.n8302 GND.n8301 240.244
R17765 GND.n8298 GND.n8297 240.244
R17766 GND.n8294 GND.n8293 240.244
R17767 GND.n8290 GND.n8289 240.244
R17768 GND.n8286 GND.n8285 240.244
R17769 GND.n8282 GND.n8281 240.244
R17770 GND.n8278 GND.n8277 240.244
R17771 GND.n8274 GND.n8273 240.244
R17772 GND.n8270 GND.n8269 240.244
R17773 GND.n8265 GND.n8264 240.244
R17774 GND.n8261 GND.n8260 240.244
R17775 GND.n8257 GND.n8256 240.244
R17776 GND.n8253 GND.n8252 240.244
R17777 GND.n8249 GND.n8248 240.244
R17778 GND.n8245 GND.n8244 240.244
R17779 GND.n1434 GND.n1351 240.244
R17780 GND.n2936 GND.n1362 240.244
R17781 GND.n2943 GND.n2936 240.244
R17782 GND.n2943 GND.n2910 240.244
R17783 GND.n2954 GND.n2910 240.244
R17784 GND.n2954 GND.n2906 240.244
R17785 GND.n2960 GND.n2906 240.244
R17786 GND.n2960 GND.n2890 240.244
R17787 GND.n2971 GND.n2890 240.244
R17788 GND.n2971 GND.n2886 240.244
R17789 GND.n2977 GND.n2886 240.244
R17790 GND.n2977 GND.n2871 240.244
R17791 GND.n2995 GND.n2871 240.244
R17792 GND.n2995 GND.n2866 240.244
R17793 GND.n3003 GND.n2866 240.244
R17794 GND.n3003 GND.n2867 240.244
R17795 GND.n2867 GND.n2847 240.244
R17796 GND.n3028 GND.n2847 240.244
R17797 GND.n3028 GND.n2843 240.244
R17798 GND.n3034 GND.n2843 240.244
R17799 GND.n3034 GND.n2823 240.244
R17800 GND.n3061 GND.n2823 240.244
R17801 GND.n3061 GND.n2818 240.244
R17802 GND.n3069 GND.n2818 240.244
R17803 GND.n3069 GND.n2819 240.244
R17804 GND.n2819 GND.n2794 240.244
R17805 GND.n3098 GND.n2794 240.244
R17806 GND.n3098 GND.n2789 240.244
R17807 GND.n3106 GND.n2789 240.244
R17808 GND.n3106 GND.n2790 240.244
R17809 GND.n2790 GND.n2764 240.244
R17810 GND.n3136 GND.n2764 240.244
R17811 GND.n3136 GND.n2759 240.244
R17812 GND.n3144 GND.n2759 240.244
R17813 GND.n3144 GND.n2760 240.244
R17814 GND.n2760 GND.n2737 240.244
R17815 GND.n3174 GND.n2737 240.244
R17816 GND.n3174 GND.n2732 240.244
R17817 GND.n3182 GND.n2732 240.244
R17818 GND.n3182 GND.n2733 240.244
R17819 GND.n2733 GND.n2708 240.244
R17820 GND.n3211 GND.n2708 240.244
R17821 GND.n3211 GND.n2703 240.244
R17822 GND.n3219 GND.n2703 240.244
R17823 GND.n3219 GND.n2704 240.244
R17824 GND.n2704 GND.n2679 240.244
R17825 GND.n3248 GND.n2679 240.244
R17826 GND.n3248 GND.n2674 240.244
R17827 GND.n3256 GND.n2674 240.244
R17828 GND.n3256 GND.n2675 240.244
R17829 GND.n2675 GND.n2649 240.244
R17830 GND.n3285 GND.n2649 240.244
R17831 GND.n3285 GND.n2644 240.244
R17832 GND.n3294 GND.n2644 240.244
R17833 GND.n3294 GND.n2645 240.244
R17834 GND.n2645 GND.n2620 240.244
R17835 GND.n3321 GND.n2620 240.244
R17836 GND.n3323 GND.n3321 240.244
R17837 GND.n3326 GND.n3323 240.244
R17838 GND.n3326 GND.n3325 240.244
R17839 GND.n3325 GND.n1537 240.244
R17840 GND.n8122 GND.n1537 240.244
R17841 GND.n8122 GND.n1538 240.244
R17842 GND.n3555 GND.n1538 240.244
R17843 GND.n3555 GND.n1550 240.244
R17844 GND.n8117 GND.n1550 240.244
R17845 GND.n8117 GND.n1551 240.244
R17846 GND.n2582 GND.n1551 240.244
R17847 GND.n3576 GND.n2582 240.244
R17848 GND.n3576 GND.n2576 240.244
R17849 GND.n3584 GND.n2576 240.244
R17850 GND.n3584 GND.n2578 240.244
R17851 GND.n2578 GND.n2560 240.244
R17852 GND.n3602 GND.n2560 240.244
R17853 GND.n3602 GND.n2553 240.244
R17854 GND.n3610 GND.n2553 240.244
R17855 GND.n3610 GND.n2556 240.244
R17856 GND.n2556 GND.n2539 240.244
R17857 GND.n3628 GND.n2539 240.244
R17858 GND.n3628 GND.n2533 240.244
R17859 GND.n3636 GND.n2533 240.244
R17860 GND.n3636 GND.n2535 240.244
R17861 GND.n2535 GND.n2517 240.244
R17862 GND.n3654 GND.n2517 240.244
R17863 GND.n3654 GND.n2511 240.244
R17864 GND.n3662 GND.n2511 240.244
R17865 GND.n3662 GND.n2513 240.244
R17866 GND.n2513 GND.n2495 240.244
R17867 GND.n3679 GND.n2495 240.244
R17868 GND.n3679 GND.n2489 240.244
R17869 GND.n3687 GND.n2489 240.244
R17870 GND.n3687 GND.n2491 240.244
R17871 GND.n2491 GND.n2473 240.244
R17872 GND.n3705 GND.n2473 240.244
R17873 GND.n3705 GND.n2466 240.244
R17874 GND.n3713 GND.n2466 240.244
R17875 GND.n3713 GND.n2469 240.244
R17876 GND.n2469 GND.n2452 240.244
R17877 GND.n3731 GND.n2452 240.244
R17878 GND.n3731 GND.n2447 240.244
R17879 GND.n3739 GND.n2447 240.244
R17880 GND.n3739 GND.n2448 240.244
R17881 GND.n2448 GND.n2432 240.244
R17882 GND.n3757 GND.n2432 240.244
R17883 GND.n3757 GND.n2426 240.244
R17884 GND.n3765 GND.n2426 240.244
R17885 GND.n3765 GND.n2428 240.244
R17886 GND.n2428 GND.n2410 240.244
R17887 GND.n3782 GND.n2410 240.244
R17888 GND.n3782 GND.n2404 240.244
R17889 GND.n3790 GND.n2404 240.244
R17890 GND.n3790 GND.n2406 240.244
R17891 GND.n2406 GND.n2388 240.244
R17892 GND.n3808 GND.n2388 240.244
R17893 GND.n3808 GND.n2381 240.244
R17894 GND.n3816 GND.n2381 240.244
R17895 GND.n3816 GND.n2384 240.244
R17896 GND.n2384 GND.n2367 240.244
R17897 GND.n3835 GND.n2367 240.244
R17898 GND.n3835 GND.n2363 240.244
R17899 GND.n3842 GND.n2363 240.244
R17900 GND.n3842 GND.n1677 240.244
R17901 GND.n6318 GND.n6317 240.244
R17902 GND.n6324 GND.n6323 240.244
R17903 GND.n6328 GND.n6327 240.244
R17904 GND.n6334 GND.n6333 240.244
R17905 GND.n6338 GND.n6337 240.244
R17906 GND.n5489 GND.n5488 240.244
R17907 GND.n5484 GND.n5483 240.244
R17908 GND.n5479 GND.n5478 240.244
R17909 GND.n5474 GND.n5473 240.244
R17910 GND.n5469 GND.n5468 240.244
R17911 GND.n6354 GND.n6353 240.244
R17912 GND.n6351 GND.n6350 240.244
R17913 GND.n6347 GND.n4421 240.244
R17914 GND.n7698 GND.n3884 240.244
R17915 GND.n7690 GND.n3884 240.244
R17916 GND.n7690 GND.n3897 240.244
R17917 GND.n7686 GND.n3897 240.244
R17918 GND.n7686 GND.n3902 240.244
R17919 GND.n7679 GND.n3902 240.244
R17920 GND.n7679 GND.n3916 240.244
R17921 GND.n7675 GND.n3916 240.244
R17922 GND.n7675 GND.n3922 240.244
R17923 GND.n3937 GND.n3922 240.244
R17924 GND.n3976 GND.n3937 240.244
R17925 GND.n3977 GND.n3976 240.244
R17926 GND.n3977 GND.n3953 240.244
R17927 GND.n3967 GND.n3953 240.244
R17928 GND.n7648 GND.n3967 240.244
R17929 GND.n7648 GND.n3968 240.244
R17930 GND.n7644 GND.n3968 240.244
R17931 GND.n7644 GND.n3986 240.244
R17932 GND.n7636 GND.n3986 240.244
R17933 GND.n7636 GND.n4000 240.244
R17934 GND.n7632 GND.n4000 240.244
R17935 GND.n7632 GND.n4006 240.244
R17936 GND.n7624 GND.n4006 240.244
R17937 GND.n7624 GND.n4020 240.244
R17938 GND.n7620 GND.n4020 240.244
R17939 GND.n7620 GND.n4026 240.244
R17940 GND.n4041 GND.n4026 240.244
R17941 GND.n4081 GND.n4041 240.244
R17942 GND.n4082 GND.n4081 240.244
R17943 GND.n4082 GND.n4058 240.244
R17944 GND.n4072 GND.n4058 240.244
R17945 GND.n7593 GND.n4072 240.244
R17946 GND.n7593 GND.n4073 240.244
R17947 GND.n7589 GND.n4073 240.244
R17948 GND.n7589 GND.n4091 240.244
R17949 GND.n7581 GND.n4091 240.244
R17950 GND.n7581 GND.n4105 240.244
R17951 GND.n7577 GND.n4105 240.244
R17952 GND.n7577 GND.n4111 240.244
R17953 GND.n7569 GND.n4111 240.244
R17954 GND.n7569 GND.n4125 240.244
R17955 GND.n7565 GND.n4125 240.244
R17956 GND.n7565 GND.n4131 240.244
R17957 GND.n4146 GND.n4131 240.244
R17958 GND.n4186 GND.n4146 240.244
R17959 GND.n4187 GND.n4186 240.244
R17960 GND.n4187 GND.n4163 240.244
R17961 GND.n4177 GND.n4163 240.244
R17962 GND.n7538 GND.n4177 240.244
R17963 GND.n7538 GND.n4178 240.244
R17964 GND.n7534 GND.n4178 240.244
R17965 GND.n7534 GND.n4196 240.244
R17966 GND.n7526 GND.n4196 240.244
R17967 GND.n7526 GND.n4209 240.244
R17968 GND.n7522 GND.n4209 240.244
R17969 GND.n7522 GND.n4215 240.244
R17970 GND.n7514 GND.n4215 240.244
R17971 GND.n7514 GND.n4228 240.244
R17972 GND.n7510 GND.n4228 240.244
R17973 GND.n7510 GND.n4234 240.244
R17974 GND.n4249 GND.n4234 240.244
R17975 GND.n4288 GND.n4249 240.244
R17976 GND.n4289 GND.n4288 240.244
R17977 GND.n4289 GND.n4266 240.244
R17978 GND.n4279 GND.n4266 240.244
R17979 GND.n7483 GND.n4279 240.244
R17980 GND.n7483 GND.n4280 240.244
R17981 GND.n7479 GND.n4280 240.244
R17982 GND.n7479 GND.n4298 240.244
R17983 GND.n7471 GND.n4298 240.244
R17984 GND.n7471 GND.n4312 240.244
R17985 GND.n7467 GND.n4312 240.244
R17986 GND.n7467 GND.n4318 240.244
R17987 GND.n7459 GND.n4318 240.244
R17988 GND.n7459 GND.n4332 240.244
R17989 GND.n7455 GND.n4332 240.244
R17990 GND.n7455 GND.n4338 240.244
R17991 GND.n4353 GND.n4338 240.244
R17992 GND.n4393 GND.n4353 240.244
R17993 GND.n4394 GND.n4393 240.244
R17994 GND.n4394 GND.n4370 240.244
R17995 GND.n4384 GND.n4370 240.244
R17996 GND.n7428 GND.n4384 240.244
R17997 GND.n7428 GND.n4385 240.244
R17998 GND.n7424 GND.n4385 240.244
R17999 GND.n7424 GND.n4403 240.244
R18000 GND.n7416 GND.n4403 240.244
R18001 GND.n7416 GND.n4416 240.244
R18002 GND.n2343 GND.n2342 240.244
R18003 GND.n7752 GND.n2342 240.244
R18004 GND.n7750 GND.n7749 240.244
R18005 GND.n7746 GND.n7745 240.244
R18006 GND.n7742 GND.n7741 240.244
R18007 GND.n2356 GND.n2355 240.244
R18008 GND.n7734 GND.n7733 240.244
R18009 GND.n7729 GND.n7728 240.244
R18010 GND.n7724 GND.n7723 240.244
R18011 GND.n7719 GND.n7718 240.244
R18012 GND.n7714 GND.n7713 240.244
R18013 GND.n7709 GND.n3875 240.244
R18014 GND.n7706 GND.n7705 240.244
R18015 GND.n3880 GND.n2340 240.244
R18016 GND.n5684 GND.n2344 240.244
R18017 GND.n5684 GND.n3895 240.244
R18018 GND.n5678 GND.n3895 240.244
R18019 GND.n5678 GND.n3904 240.244
R18020 GND.n5675 GND.n3904 240.244
R18021 GND.n5675 GND.n3914 240.244
R18022 GND.n5760 GND.n3914 240.244
R18023 GND.n5760 GND.n3924 240.244
R18024 GND.n5650 GND.n3924 240.244
R18025 GND.n5650 GND.n3935 240.244
R18026 GND.n5768 GND.n3935 240.244
R18027 GND.n5769 GND.n5768 240.244
R18028 GND.n5769 GND.n3952 240.244
R18029 GND.n5796 GND.n3952 240.244
R18030 GND.n5796 GND.n3965 240.244
R18031 GND.n5792 GND.n3965 240.244
R18032 GND.n5792 GND.n3988 240.244
R18033 GND.n5789 GND.n3988 240.244
R18034 GND.n5789 GND.n3998 240.244
R18035 GND.n5786 GND.n3998 240.244
R18036 GND.n5786 GND.n4008 240.244
R18037 GND.n5783 GND.n4008 240.244
R18038 GND.n5783 GND.n4018 240.244
R18039 GND.n5864 GND.n4018 240.244
R18040 GND.n5864 GND.n4028 240.244
R18041 GND.n5619 GND.n4028 240.244
R18042 GND.n5619 GND.n4039 240.244
R18043 GND.n5872 GND.n4039 240.244
R18044 GND.n5873 GND.n5872 240.244
R18045 GND.n5873 GND.n4056 240.244
R18046 GND.n5900 GND.n4056 240.244
R18047 GND.n5900 GND.n4070 240.244
R18048 GND.n5896 GND.n4070 240.244
R18049 GND.n5896 GND.n4093 240.244
R18050 GND.n5893 GND.n4093 240.244
R18051 GND.n5893 GND.n4103 240.244
R18052 GND.n5890 GND.n4103 240.244
R18053 GND.n5890 GND.n4113 240.244
R18054 GND.n5887 GND.n4113 240.244
R18055 GND.n5887 GND.n4123 240.244
R18056 GND.n5967 GND.n4123 240.244
R18057 GND.n5967 GND.n4133 240.244
R18058 GND.n5588 GND.n4133 240.244
R18059 GND.n5588 GND.n4144 240.244
R18060 GND.n5975 GND.n4144 240.244
R18061 GND.n5976 GND.n5975 240.244
R18062 GND.n5976 GND.n4161 240.244
R18063 GND.n6003 GND.n4161 240.244
R18064 GND.n6003 GND.n4175 240.244
R18065 GND.n5999 GND.n4175 240.244
R18066 GND.n5999 GND.n4198 240.244
R18067 GND.n5996 GND.n4198 240.244
R18068 GND.n5996 GND.n4207 240.244
R18069 GND.n5993 GND.n4207 240.244
R18070 GND.n5993 GND.n4217 240.244
R18071 GND.n5990 GND.n4217 240.244
R18072 GND.n5990 GND.n4227 240.244
R18073 GND.n6070 GND.n4227 240.244
R18074 GND.n6070 GND.n4236 240.244
R18075 GND.n5555 GND.n4236 240.244
R18076 GND.n5555 GND.n4247 240.244
R18077 GND.n6078 GND.n4247 240.244
R18078 GND.n6079 GND.n6078 240.244
R18079 GND.n6079 GND.n4264 240.244
R18080 GND.n6106 GND.n4264 240.244
R18081 GND.n6106 GND.n4278 240.244
R18082 GND.n6102 GND.n4278 240.244
R18083 GND.n6102 GND.n4300 240.244
R18084 GND.n6099 GND.n4300 240.244
R18085 GND.n6099 GND.n4310 240.244
R18086 GND.n6096 GND.n4310 240.244
R18087 GND.n6096 GND.n4320 240.244
R18088 GND.n6093 GND.n4320 240.244
R18089 GND.n6093 GND.n4330 240.244
R18090 GND.n6173 GND.n4330 240.244
R18091 GND.n6173 GND.n4340 240.244
R18092 GND.n5523 GND.n4340 240.244
R18093 GND.n5523 GND.n4351 240.244
R18094 GND.n6181 GND.n4351 240.244
R18095 GND.n6182 GND.n6181 240.244
R18096 GND.n6182 GND.n4368 240.244
R18097 GND.n6202 GND.n4368 240.244
R18098 GND.n6202 GND.n4382 240.244
R18099 GND.n6198 GND.n4382 240.244
R18100 GND.n6198 GND.n4405 240.244
R18101 GND.n6195 GND.n4405 240.244
R18102 GND.n6195 GND.n4414 240.244
R18103 GND.n6313 GND.n4414 240.244
R18104 GND.n10054 GND.n10053 240.244
R18105 GND.n10057 GND.n10056 240.244
R18106 GND.n10064 GND.n10063 240.244
R18107 GND.n10066 GND.n10044 240.244
R18108 GND.n10072 GND.n9811 240.244
R18109 GND.n6417 GND.n4884 240.244
R18110 GND.n4895 GND.n4884 240.244
R18111 GND.n6424 GND.n4895 240.244
R18112 GND.n6425 GND.n6424 240.244
R18113 GND.n6425 GND.n4908 240.244
R18114 GND.n6431 GND.n4908 240.244
R18115 GND.n6431 GND.n4925 240.244
R18116 GND.n6480 GND.n4925 240.244
R18117 GND.n6480 GND.n4937 240.244
R18118 GND.n6486 GND.n4937 240.244
R18119 GND.n6486 GND.n4948 240.244
R18120 GND.n6494 GND.n4948 240.244
R18121 GND.n6494 GND.n4958 240.244
R18122 GND.n6500 GND.n4958 240.244
R18123 GND.n6500 GND.n4969 240.244
R18124 GND.n6508 GND.n4969 240.244
R18125 GND.n6508 GND.n4979 240.244
R18126 GND.n6515 GND.n4979 240.244
R18127 GND.n6515 GND.n4990 240.244
R18128 GND.n6674 GND.n4990 240.244
R18129 GND.n6674 GND.n4999 240.244
R18130 GND.n6670 GND.n4999 240.244
R18131 GND.n6670 GND.n5010 240.244
R18132 GND.n6662 GND.n5010 240.244
R18133 GND.n6662 GND.n5020 240.244
R18134 GND.n6658 GND.n5020 240.244
R18135 GND.n6658 GND.n5031 240.244
R18136 GND.n6650 GND.n5031 240.244
R18137 GND.n6650 GND.n5041 240.244
R18138 GND.n6646 GND.n5041 240.244
R18139 GND.n6646 GND.n5052 240.244
R18140 GND.n6638 GND.n5052 240.244
R18141 GND.n6638 GND.n5062 240.244
R18142 GND.n6634 GND.n5062 240.244
R18143 GND.n6634 GND.n5073 240.244
R18144 GND.n6626 GND.n5073 240.244
R18145 GND.n6626 GND.n5083 240.244
R18146 GND.n6622 GND.n5083 240.244
R18147 GND.n6622 GND.n5094 240.244
R18148 GND.n6614 GND.n5094 240.244
R18149 GND.n6614 GND.n5104 240.244
R18150 GND.n6610 GND.n5104 240.244
R18151 GND.n6610 GND.n5115 240.244
R18152 GND.n6602 GND.n5115 240.244
R18153 GND.n6602 GND.n5125 240.244
R18154 GND.n6598 GND.n5125 240.244
R18155 GND.n6598 GND.n5136 240.244
R18156 GND.n6590 GND.n5136 240.244
R18157 GND.n6590 GND.n5146 240.244
R18158 GND.n6586 GND.n5146 240.244
R18159 GND.n6586 GND.n5157 240.244
R18160 GND.n6578 GND.n5157 240.244
R18161 GND.n6578 GND.n5167 240.244
R18162 GND.n6755 GND.n5167 240.244
R18163 GND.n6755 GND.n5176 240.244
R18164 GND.n6768 GND.n5176 240.244
R18165 GND.n6768 GND.n5186 240.244
R18166 GND.n5191 GND.n5186 240.244
R18167 GND.n6763 GND.n5191 240.244
R18168 GND.n6763 GND.n106 240.244
R18169 GND.n10311 GND.n106 240.244
R18170 GND.n10311 GND.n107 240.244
R18171 GND.n5271 GND.n107 240.244
R18172 GND.n6900 GND.n5271 240.244
R18173 GND.n6900 GND.n129 240.244
R18174 GND.n6896 GND.n129 240.244
R18175 GND.n6896 GND.n141 240.244
R18176 GND.n6888 GND.n141 240.244
R18177 GND.n6888 GND.n151 240.244
R18178 GND.n6884 GND.n151 240.244
R18179 GND.n6884 GND.n161 240.244
R18180 GND.n6876 GND.n161 240.244
R18181 GND.n6876 GND.n172 240.244
R18182 GND.n6872 GND.n172 240.244
R18183 GND.n6872 GND.n182 240.244
R18184 GND.n6864 GND.n182 240.244
R18185 GND.n6864 GND.n193 240.244
R18186 GND.n6860 GND.n193 240.244
R18187 GND.n6860 GND.n203 240.244
R18188 GND.n6852 GND.n203 240.244
R18189 GND.n6852 GND.n214 240.244
R18190 GND.n6848 GND.n214 240.244
R18191 GND.n6848 GND.n224 240.244
R18192 GND.n6840 GND.n224 240.244
R18193 GND.n6840 GND.n235 240.244
R18194 GND.n6836 GND.n235 240.244
R18195 GND.n6836 GND.n245 240.244
R18196 GND.n9728 GND.n245 240.244
R18197 GND.n9728 GND.n255 240.244
R18198 GND.n9734 GND.n255 240.244
R18199 GND.n9734 GND.n265 240.244
R18200 GND.n9743 GND.n265 240.244
R18201 GND.n9743 GND.n276 240.244
R18202 GND.n9749 GND.n276 240.244
R18203 GND.n9749 GND.n286 240.244
R18204 GND.n9758 GND.n286 240.244
R18205 GND.n9758 GND.n297 240.244
R18206 GND.n9764 GND.n297 240.244
R18207 GND.n9764 GND.n307 240.244
R18208 GND.n9773 GND.n307 240.244
R18209 GND.n9773 GND.n318 240.244
R18210 GND.n9779 GND.n318 240.244
R18211 GND.n9779 GND.n328 240.244
R18212 GND.n9788 GND.n328 240.244
R18213 GND.n9788 GND.n339 240.244
R18214 GND.n10103 GND.n339 240.244
R18215 GND.n10103 GND.n349 240.244
R18216 GND.n10099 GND.n349 240.244
R18217 GND.n10099 GND.n360 240.244
R18218 GND.n10096 GND.n360 240.244
R18219 GND.n10096 GND.n369 240.244
R18220 GND.n10093 GND.n369 240.244
R18221 GND.n10093 GND.n379 240.244
R18222 GND.n10090 GND.n379 240.244
R18223 GND.n10090 GND.n388 240.244
R18224 GND.n10087 GND.n388 240.244
R18225 GND.n10087 GND.n398 240.244
R18226 GND.n10084 GND.n398 240.244
R18227 GND.n10084 GND.n407 240.244
R18228 GND.n10081 GND.n407 240.244
R18229 GND.n10081 GND.n416 240.244
R18230 GND.n6365 GND.n6364 240.244
R18231 GND.n6370 GND.n6369 240.244
R18232 GND.n6375 GND.n6374 240.244
R18233 GND.n6380 GND.n6379 240.244
R18234 GND.n6383 GND.n6358 240.244
R18235 GND.n7090 GND.n4886 240.244
R18236 GND.n7090 GND.n4887 240.244
R18237 GND.n5357 GND.n4887 240.244
R18238 GND.n5358 GND.n5357 240.244
R18239 GND.n5358 GND.n4910 240.244
R18240 GND.n4927 GND.n4910 240.244
R18241 GND.n7069 GND.n4927 240.244
R18242 GND.n7069 GND.n4928 240.244
R18243 GND.n7065 GND.n4928 240.244
R18244 GND.n7065 GND.n4934 240.244
R18245 GND.n7057 GND.n4934 240.244
R18246 GND.n7057 GND.n4950 240.244
R18247 GND.n7053 GND.n4950 240.244
R18248 GND.n7053 GND.n4955 240.244
R18249 GND.n7045 GND.n4955 240.244
R18250 GND.n7045 GND.n4971 240.244
R18251 GND.n7041 GND.n4971 240.244
R18252 GND.n7041 GND.n4976 240.244
R18253 GND.n7033 GND.n4976 240.244
R18254 GND.n7033 GND.n4992 240.244
R18255 GND.n7029 GND.n4992 240.244
R18256 GND.n7029 GND.n4997 240.244
R18257 GND.n7021 GND.n4997 240.244
R18258 GND.n7021 GND.n5012 240.244
R18259 GND.n7017 GND.n5012 240.244
R18260 GND.n7017 GND.n5017 240.244
R18261 GND.n7009 GND.n5017 240.244
R18262 GND.n7009 GND.n5033 240.244
R18263 GND.n7005 GND.n5033 240.244
R18264 GND.n7005 GND.n5038 240.244
R18265 GND.n6997 GND.n5038 240.244
R18266 GND.n6997 GND.n5054 240.244
R18267 GND.n6993 GND.n5054 240.244
R18268 GND.n6993 GND.n5059 240.244
R18269 GND.n6985 GND.n5059 240.244
R18270 GND.n6985 GND.n5075 240.244
R18271 GND.n6981 GND.n5075 240.244
R18272 GND.n6981 GND.n5080 240.244
R18273 GND.n6973 GND.n5080 240.244
R18274 GND.n6973 GND.n5096 240.244
R18275 GND.n6969 GND.n5096 240.244
R18276 GND.n6969 GND.n5101 240.244
R18277 GND.n6961 GND.n5101 240.244
R18278 GND.n6961 GND.n5117 240.244
R18279 GND.n6957 GND.n5117 240.244
R18280 GND.n6957 GND.n5122 240.244
R18281 GND.n6949 GND.n5122 240.244
R18282 GND.n6949 GND.n5138 240.244
R18283 GND.n6945 GND.n5138 240.244
R18284 GND.n6945 GND.n5143 240.244
R18285 GND.n6937 GND.n5143 240.244
R18286 GND.n6937 GND.n5159 240.244
R18287 GND.n6933 GND.n5159 240.244
R18288 GND.n6933 GND.n5164 240.244
R18289 GND.n6925 GND.n5164 240.244
R18290 GND.n6925 GND.n5178 240.244
R18291 GND.n6921 GND.n5178 240.244
R18292 GND.n6921 GND.n5183 240.244
R18293 GND.n5285 GND.n5183 240.244
R18294 GND.n6780 GND.n5285 240.244
R18295 GND.n6780 GND.n111 240.244
R18296 GND.n6789 GND.n111 240.244
R18297 GND.n6790 GND.n6789 240.244
R18298 GND.n6790 GND.n131 240.244
R18299 GND.n10302 GND.n131 240.244
R18300 GND.n10302 GND.n132 240.244
R18301 GND.n10298 GND.n132 240.244
R18302 GND.n10298 GND.n138 240.244
R18303 GND.n10290 GND.n138 240.244
R18304 GND.n10290 GND.n153 240.244
R18305 GND.n10286 GND.n153 240.244
R18306 GND.n10286 GND.n158 240.244
R18307 GND.n10278 GND.n158 240.244
R18308 GND.n10278 GND.n174 240.244
R18309 GND.n10274 GND.n174 240.244
R18310 GND.n10274 GND.n179 240.244
R18311 GND.n10266 GND.n179 240.244
R18312 GND.n10266 GND.n195 240.244
R18313 GND.n10262 GND.n195 240.244
R18314 GND.n10262 GND.n200 240.244
R18315 GND.n10254 GND.n200 240.244
R18316 GND.n10254 GND.n216 240.244
R18317 GND.n10250 GND.n216 240.244
R18318 GND.n10250 GND.n221 240.244
R18319 GND.n10242 GND.n221 240.244
R18320 GND.n10242 GND.n237 240.244
R18321 GND.n10238 GND.n237 240.244
R18322 GND.n10238 GND.n242 240.244
R18323 GND.n10230 GND.n242 240.244
R18324 GND.n10230 GND.n257 240.244
R18325 GND.n10226 GND.n257 240.244
R18326 GND.n10226 GND.n262 240.244
R18327 GND.n10218 GND.n262 240.244
R18328 GND.n10218 GND.n278 240.244
R18329 GND.n10214 GND.n278 240.244
R18330 GND.n10214 GND.n283 240.244
R18331 GND.n10206 GND.n283 240.244
R18332 GND.n10206 GND.n299 240.244
R18333 GND.n10202 GND.n299 240.244
R18334 GND.n10202 GND.n304 240.244
R18335 GND.n10194 GND.n304 240.244
R18336 GND.n10194 GND.n320 240.244
R18337 GND.n10190 GND.n320 240.244
R18338 GND.n10190 GND.n325 240.244
R18339 GND.n10182 GND.n325 240.244
R18340 GND.n10182 GND.n341 240.244
R18341 GND.n10178 GND.n341 240.244
R18342 GND.n10178 GND.n346 240.244
R18343 GND.n10170 GND.n346 240.244
R18344 GND.n10170 GND.n362 240.244
R18345 GND.n10166 GND.n362 240.244
R18346 GND.n10166 GND.n367 240.244
R18347 GND.n10158 GND.n367 240.244
R18348 GND.n10158 GND.n381 240.244
R18349 GND.n10154 GND.n381 240.244
R18350 GND.n10154 GND.n386 240.244
R18351 GND.n10146 GND.n386 240.244
R18352 GND.n10146 GND.n400 240.244
R18353 GND.n10142 GND.n400 240.244
R18354 GND.n10142 GND.n405 240.244
R18355 GND.n10134 GND.n405 240.244
R18356 GND.n8500 GND.n1187 240.244
R18357 GND.n8500 GND.n1183 240.244
R18358 GND.n8506 GND.n1183 240.244
R18359 GND.n8506 GND.n1181 240.244
R18360 GND.n8510 GND.n1181 240.244
R18361 GND.n8510 GND.n1177 240.244
R18362 GND.n8516 GND.n1177 240.244
R18363 GND.n8516 GND.n1175 240.244
R18364 GND.n8520 GND.n1175 240.244
R18365 GND.n8520 GND.n1171 240.244
R18366 GND.n8526 GND.n1171 240.244
R18367 GND.n8526 GND.n1169 240.244
R18368 GND.n8530 GND.n1169 240.244
R18369 GND.n8530 GND.n1165 240.244
R18370 GND.n8536 GND.n1165 240.244
R18371 GND.n8536 GND.n1163 240.244
R18372 GND.n8540 GND.n1163 240.244
R18373 GND.n8540 GND.n1159 240.244
R18374 GND.n8546 GND.n1159 240.244
R18375 GND.n8546 GND.n1157 240.244
R18376 GND.n8550 GND.n1157 240.244
R18377 GND.n8550 GND.n1153 240.244
R18378 GND.n8556 GND.n1153 240.244
R18379 GND.n8556 GND.n1151 240.244
R18380 GND.n8560 GND.n1151 240.244
R18381 GND.n8560 GND.n1147 240.244
R18382 GND.n8566 GND.n1147 240.244
R18383 GND.n8566 GND.n1145 240.244
R18384 GND.n8570 GND.n1145 240.244
R18385 GND.n8570 GND.n1141 240.244
R18386 GND.n8576 GND.n1141 240.244
R18387 GND.n8576 GND.n1139 240.244
R18388 GND.n8580 GND.n1139 240.244
R18389 GND.n8580 GND.n1135 240.244
R18390 GND.n8586 GND.n1135 240.244
R18391 GND.n8586 GND.n1133 240.244
R18392 GND.n8590 GND.n1133 240.244
R18393 GND.n8590 GND.n1129 240.244
R18394 GND.n8596 GND.n1129 240.244
R18395 GND.n8596 GND.n1127 240.244
R18396 GND.n8600 GND.n1127 240.244
R18397 GND.n8600 GND.n1123 240.244
R18398 GND.n8606 GND.n1123 240.244
R18399 GND.n8606 GND.n1121 240.244
R18400 GND.n8610 GND.n1121 240.244
R18401 GND.n8610 GND.n1117 240.244
R18402 GND.n8616 GND.n1117 240.244
R18403 GND.n8616 GND.n1115 240.244
R18404 GND.n8620 GND.n1115 240.244
R18405 GND.n8620 GND.n1111 240.244
R18406 GND.n8626 GND.n1111 240.244
R18407 GND.n8626 GND.n1109 240.244
R18408 GND.n8630 GND.n1109 240.244
R18409 GND.n8630 GND.n1105 240.244
R18410 GND.n8636 GND.n1105 240.244
R18411 GND.n8636 GND.n1103 240.244
R18412 GND.n8640 GND.n1103 240.244
R18413 GND.n8640 GND.n1099 240.244
R18414 GND.n8646 GND.n1099 240.244
R18415 GND.n8646 GND.n1097 240.244
R18416 GND.n8650 GND.n1097 240.244
R18417 GND.n8650 GND.n1093 240.244
R18418 GND.n8656 GND.n1093 240.244
R18419 GND.n8656 GND.n1091 240.244
R18420 GND.n8660 GND.n1091 240.244
R18421 GND.n8660 GND.n1087 240.244
R18422 GND.n8666 GND.n1087 240.244
R18423 GND.n8666 GND.n1085 240.244
R18424 GND.n8670 GND.n1085 240.244
R18425 GND.n8670 GND.n1081 240.244
R18426 GND.n8676 GND.n1081 240.244
R18427 GND.n8676 GND.n1079 240.244
R18428 GND.n8680 GND.n1079 240.244
R18429 GND.n8680 GND.n1075 240.244
R18430 GND.n8686 GND.n1075 240.244
R18431 GND.n8686 GND.n1073 240.244
R18432 GND.n8690 GND.n1073 240.244
R18433 GND.n8690 GND.n1069 240.244
R18434 GND.n8696 GND.n1069 240.244
R18435 GND.n8696 GND.n1067 240.244
R18436 GND.n8700 GND.n1067 240.244
R18437 GND.n8700 GND.n1063 240.244
R18438 GND.n8706 GND.n1063 240.244
R18439 GND.n8706 GND.n1061 240.244
R18440 GND.n8710 GND.n1061 240.244
R18441 GND.n8710 GND.n1057 240.244
R18442 GND.n8716 GND.n1057 240.244
R18443 GND.n8716 GND.n1055 240.244
R18444 GND.n8720 GND.n1055 240.244
R18445 GND.n8720 GND.n1051 240.244
R18446 GND.n8726 GND.n1051 240.244
R18447 GND.n8726 GND.n1049 240.244
R18448 GND.n8730 GND.n1049 240.244
R18449 GND.n8730 GND.n1045 240.244
R18450 GND.n8736 GND.n1045 240.244
R18451 GND.n8736 GND.n1043 240.244
R18452 GND.n8740 GND.n1043 240.244
R18453 GND.n8740 GND.n1039 240.244
R18454 GND.n8746 GND.n1039 240.244
R18455 GND.n8746 GND.n1037 240.244
R18456 GND.n8750 GND.n1037 240.244
R18457 GND.n8750 GND.n1033 240.244
R18458 GND.n8756 GND.n1033 240.244
R18459 GND.n8756 GND.n1031 240.244
R18460 GND.n8760 GND.n1031 240.244
R18461 GND.n8760 GND.n1027 240.244
R18462 GND.n8766 GND.n1027 240.244
R18463 GND.n8766 GND.n1025 240.244
R18464 GND.n8770 GND.n1025 240.244
R18465 GND.n8770 GND.n1021 240.244
R18466 GND.n8776 GND.n1021 240.244
R18467 GND.n8776 GND.n1019 240.244
R18468 GND.n8780 GND.n1019 240.244
R18469 GND.n8780 GND.n1015 240.244
R18470 GND.n8786 GND.n1015 240.244
R18471 GND.n8786 GND.n1013 240.244
R18472 GND.n8790 GND.n1013 240.244
R18473 GND.n8790 GND.n1009 240.244
R18474 GND.n8796 GND.n1009 240.244
R18475 GND.n8796 GND.n1007 240.244
R18476 GND.n8800 GND.n1007 240.244
R18477 GND.n8800 GND.n1003 240.244
R18478 GND.n8806 GND.n1003 240.244
R18479 GND.n8806 GND.n1001 240.244
R18480 GND.n8810 GND.n1001 240.244
R18481 GND.n8810 GND.n997 240.244
R18482 GND.n8816 GND.n997 240.244
R18483 GND.n8816 GND.n995 240.244
R18484 GND.n8820 GND.n995 240.244
R18485 GND.n8820 GND.n991 240.244
R18486 GND.n8826 GND.n991 240.244
R18487 GND.n8826 GND.n989 240.244
R18488 GND.n8830 GND.n989 240.244
R18489 GND.n8830 GND.n985 240.244
R18490 GND.n8836 GND.n985 240.244
R18491 GND.n8836 GND.n983 240.244
R18492 GND.n8840 GND.n983 240.244
R18493 GND.n8840 GND.n979 240.244
R18494 GND.n8846 GND.n979 240.244
R18495 GND.n8846 GND.n977 240.244
R18496 GND.n8850 GND.n977 240.244
R18497 GND.n8850 GND.n973 240.244
R18498 GND.n8856 GND.n973 240.244
R18499 GND.n8856 GND.n971 240.244
R18500 GND.n8860 GND.n971 240.244
R18501 GND.n8860 GND.n967 240.244
R18502 GND.n8866 GND.n967 240.244
R18503 GND.n8866 GND.n965 240.244
R18504 GND.n8870 GND.n965 240.244
R18505 GND.n8870 GND.n961 240.244
R18506 GND.n8876 GND.n961 240.244
R18507 GND.n8876 GND.n959 240.244
R18508 GND.n8880 GND.n959 240.244
R18509 GND.n8880 GND.n955 240.244
R18510 GND.n8886 GND.n955 240.244
R18511 GND.n8886 GND.n953 240.244
R18512 GND.n8890 GND.n953 240.244
R18513 GND.n8890 GND.n949 240.244
R18514 GND.n8896 GND.n949 240.244
R18515 GND.n8896 GND.n947 240.244
R18516 GND.n8900 GND.n947 240.244
R18517 GND.n8900 GND.n943 240.244
R18518 GND.n8906 GND.n943 240.244
R18519 GND.n8906 GND.n941 240.244
R18520 GND.n8910 GND.n941 240.244
R18521 GND.n8910 GND.n937 240.244
R18522 GND.n8916 GND.n937 240.244
R18523 GND.n8916 GND.n935 240.244
R18524 GND.n8920 GND.n935 240.244
R18525 GND.n8920 GND.n931 240.244
R18526 GND.n8926 GND.n931 240.244
R18527 GND.n8926 GND.n929 240.244
R18528 GND.n8930 GND.n929 240.244
R18529 GND.n8930 GND.n925 240.244
R18530 GND.n8936 GND.n925 240.244
R18531 GND.n8936 GND.n923 240.244
R18532 GND.n8940 GND.n923 240.244
R18533 GND.n8940 GND.n919 240.244
R18534 GND.n8946 GND.n919 240.244
R18535 GND.n8946 GND.n917 240.244
R18536 GND.n8950 GND.n917 240.244
R18537 GND.n8950 GND.n913 240.244
R18538 GND.n8956 GND.n913 240.244
R18539 GND.n8956 GND.n911 240.244
R18540 GND.n8960 GND.n911 240.244
R18541 GND.n8960 GND.n907 240.244
R18542 GND.n8966 GND.n907 240.244
R18543 GND.n8966 GND.n905 240.244
R18544 GND.n8970 GND.n905 240.244
R18545 GND.n8970 GND.n901 240.244
R18546 GND.n8976 GND.n901 240.244
R18547 GND.n8976 GND.n899 240.244
R18548 GND.n8980 GND.n899 240.244
R18549 GND.n8980 GND.n895 240.244
R18550 GND.n8986 GND.n895 240.244
R18551 GND.n8986 GND.n893 240.244
R18552 GND.n8990 GND.n893 240.244
R18553 GND.n8990 GND.n889 240.244
R18554 GND.n8996 GND.n889 240.244
R18555 GND.n8996 GND.n887 240.244
R18556 GND.n9000 GND.n887 240.244
R18557 GND.n9000 GND.n883 240.244
R18558 GND.n9006 GND.n883 240.244
R18559 GND.n9006 GND.n881 240.244
R18560 GND.n9010 GND.n881 240.244
R18561 GND.n9010 GND.n877 240.244
R18562 GND.n9016 GND.n877 240.244
R18563 GND.n9016 GND.n875 240.244
R18564 GND.n9020 GND.n875 240.244
R18565 GND.n9020 GND.n871 240.244
R18566 GND.n9026 GND.n871 240.244
R18567 GND.n9026 GND.n869 240.244
R18568 GND.n9030 GND.n869 240.244
R18569 GND.n9030 GND.n865 240.244
R18570 GND.n9036 GND.n865 240.244
R18571 GND.n9036 GND.n863 240.244
R18572 GND.n9040 GND.n863 240.244
R18573 GND.n9040 GND.n859 240.244
R18574 GND.n9046 GND.n859 240.244
R18575 GND.n9046 GND.n857 240.244
R18576 GND.n9050 GND.n857 240.244
R18577 GND.n9050 GND.n853 240.244
R18578 GND.n9056 GND.n853 240.244
R18579 GND.n9056 GND.n851 240.244
R18580 GND.n9060 GND.n851 240.244
R18581 GND.n9060 GND.n847 240.244
R18582 GND.n9066 GND.n847 240.244
R18583 GND.n9066 GND.n845 240.244
R18584 GND.n9070 GND.n845 240.244
R18585 GND.n9070 GND.n841 240.244
R18586 GND.n9076 GND.n841 240.244
R18587 GND.n9076 GND.n839 240.244
R18588 GND.n9080 GND.n839 240.244
R18589 GND.n9080 GND.n835 240.244
R18590 GND.n9086 GND.n835 240.244
R18591 GND.n9086 GND.n833 240.244
R18592 GND.n9090 GND.n833 240.244
R18593 GND.n9090 GND.n829 240.244
R18594 GND.n9096 GND.n829 240.244
R18595 GND.n9096 GND.n827 240.244
R18596 GND.n9100 GND.n827 240.244
R18597 GND.n9100 GND.n823 240.244
R18598 GND.n9106 GND.n823 240.244
R18599 GND.n9106 GND.n821 240.244
R18600 GND.n9110 GND.n821 240.244
R18601 GND.n9110 GND.n817 240.244
R18602 GND.n9116 GND.n817 240.244
R18603 GND.n9116 GND.n815 240.244
R18604 GND.n9120 GND.n815 240.244
R18605 GND.n9120 GND.n811 240.244
R18606 GND.n9126 GND.n811 240.244
R18607 GND.n9126 GND.n809 240.244
R18608 GND.n9130 GND.n809 240.244
R18609 GND.n9130 GND.n805 240.244
R18610 GND.n9136 GND.n805 240.244
R18611 GND.n9136 GND.n803 240.244
R18612 GND.n9140 GND.n803 240.244
R18613 GND.n9140 GND.n799 240.244
R18614 GND.n9146 GND.n799 240.244
R18615 GND.n9146 GND.n797 240.244
R18616 GND.n9150 GND.n797 240.244
R18617 GND.n9150 GND.n793 240.244
R18618 GND.n9156 GND.n793 240.244
R18619 GND.n9156 GND.n791 240.244
R18620 GND.n9160 GND.n791 240.244
R18621 GND.n9160 GND.n787 240.244
R18622 GND.n9166 GND.n787 240.244
R18623 GND.n9166 GND.n785 240.244
R18624 GND.n9170 GND.n785 240.244
R18625 GND.n9170 GND.n781 240.244
R18626 GND.n9176 GND.n781 240.244
R18627 GND.n9176 GND.n779 240.244
R18628 GND.n9180 GND.n779 240.244
R18629 GND.n9180 GND.n775 240.244
R18630 GND.n9186 GND.n775 240.244
R18631 GND.n9186 GND.n773 240.244
R18632 GND.n9190 GND.n773 240.244
R18633 GND.n9190 GND.n769 240.244
R18634 GND.n9196 GND.n769 240.244
R18635 GND.n9196 GND.n767 240.244
R18636 GND.n9200 GND.n767 240.244
R18637 GND.n9200 GND.n763 240.244
R18638 GND.n9206 GND.n763 240.244
R18639 GND.n9206 GND.n761 240.244
R18640 GND.n9210 GND.n761 240.244
R18641 GND.n9210 GND.n757 240.244
R18642 GND.n9216 GND.n757 240.244
R18643 GND.n9216 GND.n755 240.244
R18644 GND.n9220 GND.n755 240.244
R18645 GND.n9220 GND.n751 240.244
R18646 GND.n9226 GND.n751 240.244
R18647 GND.n9226 GND.n749 240.244
R18648 GND.n9230 GND.n749 240.244
R18649 GND.n9230 GND.n745 240.244
R18650 GND.n9236 GND.n745 240.244
R18651 GND.n9236 GND.n743 240.244
R18652 GND.n9240 GND.n743 240.244
R18653 GND.n9240 GND.n739 240.244
R18654 GND.n9246 GND.n739 240.244
R18655 GND.n9246 GND.n737 240.244
R18656 GND.n9250 GND.n737 240.244
R18657 GND.n9250 GND.n733 240.244
R18658 GND.n9256 GND.n733 240.244
R18659 GND.n9256 GND.n731 240.244
R18660 GND.n9260 GND.n731 240.244
R18661 GND.n9260 GND.n727 240.244
R18662 GND.n9266 GND.n727 240.244
R18663 GND.n9266 GND.n725 240.244
R18664 GND.n9270 GND.n725 240.244
R18665 GND.n9270 GND.n721 240.244
R18666 GND.n9276 GND.n721 240.244
R18667 GND.n9276 GND.n719 240.244
R18668 GND.n9280 GND.n719 240.244
R18669 GND.n9280 GND.n715 240.244
R18670 GND.n9286 GND.n715 240.244
R18671 GND.n9286 GND.n713 240.244
R18672 GND.n9290 GND.n713 240.244
R18673 GND.n9290 GND.n709 240.244
R18674 GND.n9296 GND.n709 240.244
R18675 GND.n9296 GND.n707 240.244
R18676 GND.n9300 GND.n707 240.244
R18677 GND.n9300 GND.n703 240.244
R18678 GND.n9306 GND.n703 240.244
R18679 GND.n9306 GND.n701 240.244
R18680 GND.n9310 GND.n701 240.244
R18681 GND.n9310 GND.n697 240.244
R18682 GND.n9316 GND.n697 240.244
R18683 GND.n9316 GND.n695 240.244
R18684 GND.n9320 GND.n695 240.244
R18685 GND.n9320 GND.n691 240.244
R18686 GND.n9326 GND.n691 240.244
R18687 GND.n9326 GND.n689 240.244
R18688 GND.n9330 GND.n689 240.244
R18689 GND.n9330 GND.n685 240.244
R18690 GND.n9336 GND.n685 240.244
R18691 GND.n9336 GND.n683 240.244
R18692 GND.n9340 GND.n683 240.244
R18693 GND.n9340 GND.n679 240.244
R18694 GND.n9346 GND.n679 240.244
R18695 GND.n9346 GND.n677 240.244
R18696 GND.n9350 GND.n677 240.244
R18697 GND.n9350 GND.n673 240.244
R18698 GND.n9356 GND.n673 240.244
R18699 GND.n9356 GND.n671 240.244
R18700 GND.n9360 GND.n671 240.244
R18701 GND.n9360 GND.n667 240.244
R18702 GND.n9366 GND.n667 240.244
R18703 GND.n9366 GND.n665 240.244
R18704 GND.n9370 GND.n665 240.244
R18705 GND.n9370 GND.n661 240.244
R18706 GND.n9376 GND.n661 240.244
R18707 GND.n9376 GND.n659 240.244
R18708 GND.n9380 GND.n659 240.244
R18709 GND.n9380 GND.n655 240.244
R18710 GND.n9386 GND.n655 240.244
R18711 GND.n9386 GND.n653 240.244
R18712 GND.n9390 GND.n653 240.244
R18713 GND.n9390 GND.n649 240.244
R18714 GND.n9396 GND.n649 240.244
R18715 GND.n9396 GND.n647 240.244
R18716 GND.n9400 GND.n647 240.244
R18717 GND.n9400 GND.n643 240.244
R18718 GND.n9406 GND.n643 240.244
R18719 GND.n9406 GND.n641 240.244
R18720 GND.n9410 GND.n641 240.244
R18721 GND.n9410 GND.n637 240.244
R18722 GND.n9416 GND.n637 240.244
R18723 GND.n9416 GND.n635 240.244
R18724 GND.n9420 GND.n635 240.244
R18725 GND.n9420 GND.n631 240.244
R18726 GND.n9426 GND.n631 240.244
R18727 GND.n9426 GND.n629 240.244
R18728 GND.n9430 GND.n629 240.244
R18729 GND.n9430 GND.n625 240.244
R18730 GND.n9436 GND.n625 240.244
R18731 GND.n9436 GND.n623 240.244
R18732 GND.n9440 GND.n623 240.244
R18733 GND.n9440 GND.n619 240.244
R18734 GND.n9446 GND.n619 240.244
R18735 GND.n9446 GND.n617 240.244
R18736 GND.n9450 GND.n617 240.244
R18737 GND.n9450 GND.n613 240.244
R18738 GND.n9456 GND.n613 240.244
R18739 GND.n9456 GND.n611 240.244
R18740 GND.n9460 GND.n611 240.244
R18741 GND.n9460 GND.n607 240.244
R18742 GND.n9466 GND.n607 240.244
R18743 GND.n9466 GND.n605 240.244
R18744 GND.n9470 GND.n605 240.244
R18745 GND.n9470 GND.n601 240.244
R18746 GND.n9476 GND.n601 240.244
R18747 GND.n9476 GND.n599 240.244
R18748 GND.n9480 GND.n599 240.244
R18749 GND.n9480 GND.n595 240.244
R18750 GND.n9486 GND.n595 240.244
R18751 GND.n9486 GND.n593 240.244
R18752 GND.n9490 GND.n593 240.244
R18753 GND.n9490 GND.n589 240.244
R18754 GND.n9496 GND.n589 240.244
R18755 GND.n9496 GND.n587 240.244
R18756 GND.n9500 GND.n587 240.244
R18757 GND.n9500 GND.n583 240.244
R18758 GND.n9506 GND.n583 240.244
R18759 GND.n9506 GND.n581 240.244
R18760 GND.n9510 GND.n581 240.244
R18761 GND.n9510 GND.n577 240.244
R18762 GND.n9517 GND.n577 240.244
R18763 GND.n9517 GND.n575 240.244
R18764 GND.n9521 GND.n575 240.244
R18765 GND.n9521 GND.n572 240.244
R18766 GND.n9527 GND.n570 240.244
R18767 GND.n9531 GND.n570 240.244
R18768 GND.n9531 GND.n566 240.244
R18769 GND.n9537 GND.n566 240.244
R18770 GND.n9537 GND.n564 240.244
R18771 GND.n9541 GND.n564 240.244
R18772 GND.n9541 GND.n560 240.244
R18773 GND.n9547 GND.n560 240.244
R18774 GND.n9547 GND.n558 240.244
R18775 GND.n9551 GND.n558 240.244
R18776 GND.n9551 GND.n554 240.244
R18777 GND.n9557 GND.n554 240.244
R18778 GND.n9557 GND.n552 240.244
R18779 GND.n9561 GND.n552 240.244
R18780 GND.n9561 GND.n548 240.244
R18781 GND.n9567 GND.n548 240.244
R18782 GND.n9567 GND.n546 240.244
R18783 GND.n9571 GND.n546 240.244
R18784 GND.n9571 GND.n542 240.244
R18785 GND.n9577 GND.n542 240.244
R18786 GND.n9577 GND.n540 240.244
R18787 GND.n9581 GND.n540 240.244
R18788 GND.n9581 GND.n536 240.244
R18789 GND.n9587 GND.n536 240.244
R18790 GND.n9587 GND.n534 240.244
R18791 GND.n9591 GND.n534 240.244
R18792 GND.n9591 GND.n530 240.244
R18793 GND.n9597 GND.n530 240.244
R18794 GND.n9597 GND.n528 240.244
R18795 GND.n9601 GND.n528 240.244
R18796 GND.n9601 GND.n524 240.244
R18797 GND.n9607 GND.n524 240.244
R18798 GND.n9607 GND.n522 240.244
R18799 GND.n9611 GND.n522 240.244
R18800 GND.n9611 GND.n518 240.244
R18801 GND.n9617 GND.n518 240.244
R18802 GND.n9617 GND.n516 240.244
R18803 GND.n9621 GND.n516 240.244
R18804 GND.n9621 GND.n512 240.244
R18805 GND.n9627 GND.n512 240.244
R18806 GND.n9627 GND.n510 240.244
R18807 GND.n9631 GND.n510 240.244
R18808 GND.n9631 GND.n506 240.244
R18809 GND.n9637 GND.n506 240.244
R18810 GND.n9637 GND.n504 240.244
R18811 GND.n9641 GND.n504 240.244
R18812 GND.n9641 GND.n500 240.244
R18813 GND.n9647 GND.n500 240.244
R18814 GND.n9647 GND.n498 240.244
R18815 GND.n9651 GND.n498 240.244
R18816 GND.n9651 GND.n494 240.244
R18817 GND.n9657 GND.n494 240.244
R18818 GND.n9657 GND.n492 240.244
R18819 GND.n9661 GND.n492 240.244
R18820 GND.n9661 GND.n488 240.244
R18821 GND.n9667 GND.n488 240.244
R18822 GND.n9667 GND.n486 240.244
R18823 GND.n9671 GND.n486 240.244
R18824 GND.n9671 GND.n482 240.244
R18825 GND.n9677 GND.n482 240.244
R18826 GND.n9677 GND.n480 240.244
R18827 GND.n9681 GND.n480 240.244
R18828 GND.n9681 GND.n476 240.244
R18829 GND.n9691 GND.n476 240.244
R18830 GND.n9691 GND.n473 240.244
R18831 GND.n9695 GND.n473 240.244
R18832 GND.n3006 GND.n1321 240.244
R18833 GND.n3016 GND.n3006 240.244
R18834 GND.n3016 GND.n3007 240.244
R18835 GND.n3007 GND.n2839 240.244
R18836 GND.n3037 GND.n2839 240.244
R18837 GND.n3037 GND.n2835 240.244
R18838 GND.n3043 GND.n2835 240.244
R18839 GND.n3043 GND.n2812 240.244
R18840 GND.n3072 GND.n2812 240.244
R18841 GND.n3072 GND.n2807 240.244
R18842 GND.n3080 GND.n2807 240.244
R18843 GND.n3080 GND.n2808 240.244
R18844 GND.n2808 GND.n2783 240.244
R18845 GND.n3109 GND.n2783 240.244
R18846 GND.n3109 GND.n2778 240.244
R18847 GND.n3117 GND.n2778 240.244
R18848 GND.n3117 GND.n2779 240.244
R18849 GND.n2779 GND.n2755 240.244
R18850 GND.n3147 GND.n2755 240.244
R18851 GND.n3147 GND.n2750 240.244
R18852 GND.n3155 GND.n2750 240.244
R18853 GND.n3155 GND.n2751 240.244
R18854 GND.n2751 GND.n2727 240.244
R18855 GND.n3185 GND.n2727 240.244
R18856 GND.n3185 GND.n2722 240.244
R18857 GND.n3193 GND.n2722 240.244
R18858 GND.n3193 GND.n2723 240.244
R18859 GND.n2723 GND.n2697 240.244
R18860 GND.n3222 GND.n2697 240.244
R18861 GND.n3222 GND.n2692 240.244
R18862 GND.n3230 GND.n2692 240.244
R18863 GND.n3230 GND.n2693 240.244
R18864 GND.n2693 GND.n2668 240.244
R18865 GND.n3259 GND.n2668 240.244
R18866 GND.n3259 GND.n2663 240.244
R18867 GND.n3267 GND.n2663 240.244
R18868 GND.n3267 GND.n2664 240.244
R18869 GND.n2664 GND.n2639 240.244
R18870 GND.n3297 GND.n2639 240.244
R18871 GND.n3297 GND.n2634 240.244
R18872 GND.n3305 GND.n2634 240.244
R18873 GND.n3305 GND.n2635 240.244
R18874 GND.n2635 GND.n2614 240.244
R18875 GND.n3329 GND.n2614 240.244
R18876 GND.n3329 GND.n2611 240.244
R18877 GND.n3540 GND.n2611 240.244
R18878 GND.n3540 GND.n2612 240.244
R18879 GND.n3535 GND.n2612 240.244
R18880 GND.n3535 GND.n3534 240.244
R18881 GND.n3534 GND.n3334 240.244
R18882 GND.n3529 GND.n3334 240.244
R18883 GND.n3529 GND.n3528 240.244
R18884 GND.n3528 GND.n3527 240.244
R18885 GND.n3527 GND.n3336 240.244
R18886 GND.n3523 GND.n3336 240.244
R18887 GND.n3523 GND.n3522 240.244
R18888 GND.n3522 GND.n3521 240.244
R18889 GND.n3521 GND.n3342 240.244
R18890 GND.n3517 GND.n3342 240.244
R18891 GND.n3517 GND.n3516 240.244
R18892 GND.n3516 GND.n3515 240.244
R18893 GND.n3515 GND.n3348 240.244
R18894 GND.n3511 GND.n3348 240.244
R18895 GND.n3511 GND.n3510 240.244
R18896 GND.n3510 GND.n3509 240.244
R18897 GND.n3509 GND.n3354 240.244
R18898 GND.n3505 GND.n3354 240.244
R18899 GND.n3505 GND.n3504 240.244
R18900 GND.n3504 GND.n3503 240.244
R18901 GND.n3503 GND.n3360 240.244
R18902 GND.n3499 GND.n3360 240.244
R18903 GND.n3499 GND.n3498 240.244
R18904 GND.n3498 GND.n3497 240.244
R18905 GND.n3497 GND.n3366 240.244
R18906 GND.n3493 GND.n3366 240.244
R18907 GND.n3493 GND.n3492 240.244
R18908 GND.n3492 GND.n3491 240.244
R18909 GND.n3491 GND.n3372 240.244
R18910 GND.n3487 GND.n3372 240.244
R18911 GND.n3487 GND.n3486 240.244
R18912 GND.n3486 GND.n3485 240.244
R18913 GND.n3485 GND.n3378 240.244
R18914 GND.n3481 GND.n3378 240.244
R18915 GND.n3481 GND.n3480 240.244
R18916 GND.n3480 GND.n3479 240.244
R18917 GND.n3479 GND.n3384 240.244
R18918 GND.n3475 GND.n3384 240.244
R18919 GND.n3475 GND.n3472 240.244
R18920 GND.n3472 GND.n3471 240.244
R18921 GND.n3471 GND.n3390 240.244
R18922 GND.n3467 GND.n3390 240.244
R18923 GND.n3467 GND.n3466 240.244
R18924 GND.n3466 GND.n3465 240.244
R18925 GND.n3465 GND.n3396 240.244
R18926 GND.n3461 GND.n3396 240.244
R18927 GND.n3461 GND.n3460 240.244
R18928 GND.n3460 GND.n3459 240.244
R18929 GND.n3459 GND.n3402 240.244
R18930 GND.n3455 GND.n3402 240.244
R18931 GND.n3455 GND.n3454 240.244
R18932 GND.n3454 GND.n3453 240.244
R18933 GND.n3453 GND.n3408 240.244
R18934 GND.n3449 GND.n3408 240.244
R18935 GND.n3449 GND.n3448 240.244
R18936 GND.n3448 GND.n3447 240.244
R18937 GND.n3447 GND.n3414 240.244
R18938 GND.n3443 GND.n3414 240.244
R18939 GND.n3443 GND.n3442 240.244
R18940 GND.n3442 GND.n3441 240.244
R18941 GND.n3441 GND.n3420 240.244
R18942 GND.n3437 GND.n3420 240.244
R18943 GND.n3437 GND.n3434 240.244
R18944 GND.n3434 GND.n3433 240.244
R18945 GND.n3433 GND.n3426 240.244
R18946 GND.n3426 GND.n1939 240.244
R18947 GND.n7909 GND.n1939 240.244
R18948 GND.n7909 GND.n1940 240.244
R18949 GND.n7905 GND.n1940 240.244
R18950 GND.n7905 GND.n1946 240.244
R18951 GND.n7896 GND.n1946 240.244
R18952 GND.n7896 GND.n1957 240.244
R18953 GND.n7892 GND.n1957 240.244
R18954 GND.n7892 GND.n1963 240.244
R18955 GND.n7882 GND.n1963 240.244
R18956 GND.n7882 GND.n1974 240.244
R18957 GND.n7878 GND.n1974 240.244
R18958 GND.n7878 GND.n1980 240.244
R18959 GND.n7868 GND.n1980 240.244
R18960 GND.n7868 GND.n1992 240.244
R18961 GND.n7864 GND.n1992 240.244
R18962 GND.n7864 GND.n1998 240.244
R18963 GND.n7854 GND.n1998 240.244
R18964 GND.n7854 GND.n2010 240.244
R18965 GND.n7850 GND.n2010 240.244
R18966 GND.n7850 GND.n2016 240.244
R18967 GND.n7840 GND.n2016 240.244
R18968 GND.n7840 GND.n2028 240.244
R18969 GND.n7836 GND.n2028 240.244
R18970 GND.n7836 GND.n2034 240.244
R18971 GND.n7826 GND.n2034 240.244
R18972 GND.n7826 GND.n2046 240.244
R18973 GND.n7822 GND.n2046 240.244
R18974 GND.n7822 GND.n2052 240.244
R18975 GND.n7812 GND.n2052 240.244
R18976 GND.n7812 GND.n2064 240.244
R18977 GND.n7808 GND.n2064 240.244
R18978 GND.n7808 GND.n2070 240.244
R18979 GND.n7798 GND.n2070 240.244
R18980 GND.n7798 GND.n2082 240.244
R18981 GND.n7794 GND.n2082 240.244
R18982 GND.n7794 GND.n2088 240.244
R18983 GND.n7784 GND.n2088 240.244
R18984 GND.n7784 GND.n2100 240.244
R18985 GND.n7780 GND.n2100 240.244
R18986 GND.n7780 GND.n2106 240.244
R18987 GND.n2317 GND.n2106 240.244
R18988 GND.n7765 GND.n2317 240.244
R18989 GND.n7765 GND.n2318 240.244
R18990 GND.n7761 GND.n2318 240.244
R18991 GND.n7761 GND.n2326 240.244
R18992 GND.n7696 GND.n2326 240.244
R18993 GND.n7696 GND.n3887 240.244
R18994 GND.n7692 GND.n3887 240.244
R18995 GND.n7692 GND.n3893 240.244
R18996 GND.n7685 GND.n3893 240.244
R18997 GND.n7685 GND.n3906 240.244
R18998 GND.n7681 GND.n3906 240.244
R18999 GND.n7681 GND.n3912 240.244
R19000 GND.n7673 GND.n3912 240.244
R19001 GND.n7673 GND.n3926 240.244
R19002 GND.n7669 GND.n3926 240.244
R19003 GND.n7669 GND.n3932 240.244
R19004 GND.n3954 GND.n3932 240.244
R19005 GND.n7654 GND.n3954 240.244
R19006 GND.n7654 GND.n3955 240.244
R19007 GND.n7650 GND.n3955 240.244
R19008 GND.n7650 GND.n3963 240.244
R19009 GND.n7642 GND.n3963 240.244
R19010 GND.n7642 GND.n3990 240.244
R19011 GND.n7638 GND.n3990 240.244
R19012 GND.n7638 GND.n3996 240.244
R19013 GND.n7630 GND.n3996 240.244
R19014 GND.n7630 GND.n4010 240.244
R19015 GND.n7626 GND.n4010 240.244
R19016 GND.n7626 GND.n4016 240.244
R19017 GND.n7618 GND.n4016 240.244
R19018 GND.n7618 GND.n4030 240.244
R19019 GND.n7614 GND.n4030 240.244
R19020 GND.n7614 GND.n4036 240.244
R19021 GND.n4059 GND.n4036 240.244
R19022 GND.n7599 GND.n4059 240.244
R19023 GND.n7599 GND.n4060 240.244
R19024 GND.n7595 GND.n4060 240.244
R19025 GND.n7595 GND.n4068 240.244
R19026 GND.n7587 GND.n4068 240.244
R19027 GND.n7587 GND.n4095 240.244
R19028 GND.n7583 GND.n4095 240.244
R19029 GND.n7583 GND.n4101 240.244
R19030 GND.n7575 GND.n4101 240.244
R19031 GND.n7575 GND.n4115 240.244
R19032 GND.n7571 GND.n4115 240.244
R19033 GND.n7571 GND.n4121 240.244
R19034 GND.n7563 GND.n4121 240.244
R19035 GND.n7563 GND.n4135 240.244
R19036 GND.n7559 GND.n4135 240.244
R19037 GND.n7559 GND.n4141 240.244
R19038 GND.n4164 GND.n4141 240.244
R19039 GND.n7544 GND.n4164 240.244
R19040 GND.n7544 GND.n4165 240.244
R19041 GND.n7540 GND.n4165 240.244
R19042 GND.n7540 GND.n4173 240.244
R19043 GND.n7532 GND.n4173 240.244
R19044 GND.n7532 GND.n4199 240.244
R19045 GND.n7528 GND.n4199 240.244
R19046 GND.n7528 GND.n4205 240.244
R19047 GND.n7520 GND.n4205 240.244
R19048 GND.n7520 GND.n4219 240.244
R19049 GND.n7516 GND.n4219 240.244
R19050 GND.n7516 GND.n4225 240.244
R19051 GND.n7508 GND.n4225 240.244
R19052 GND.n7508 GND.n4238 240.244
R19053 GND.n7504 GND.n4238 240.244
R19054 GND.n7504 GND.n4244 240.244
R19055 GND.n4267 GND.n4244 240.244
R19056 GND.n7489 GND.n4267 240.244
R19057 GND.n7489 GND.n4268 240.244
R19058 GND.n7485 GND.n4268 240.244
R19059 GND.n7485 GND.n4276 240.244
R19060 GND.n7477 GND.n4276 240.244
R19061 GND.n7477 GND.n4302 240.244
R19062 GND.n7473 GND.n4302 240.244
R19063 GND.n7473 GND.n4308 240.244
R19064 GND.n7465 GND.n4308 240.244
R19065 GND.n7465 GND.n4322 240.244
R19066 GND.n7461 GND.n4322 240.244
R19067 GND.n7461 GND.n4328 240.244
R19068 GND.n7453 GND.n4328 240.244
R19069 GND.n7453 GND.n4342 240.244
R19070 GND.n7449 GND.n4342 240.244
R19071 GND.n7449 GND.n4348 240.244
R19072 GND.n4371 GND.n4348 240.244
R19073 GND.n7434 GND.n4371 240.244
R19074 GND.n7434 GND.n4372 240.244
R19075 GND.n7430 GND.n4372 240.244
R19076 GND.n7430 GND.n4380 240.244
R19077 GND.n7422 GND.n4380 240.244
R19078 GND.n7422 GND.n4407 240.244
R19079 GND.n7418 GND.n4407 240.244
R19080 GND.n7418 GND.n4413 240.244
R19081 GND.n4437 GND.n4413 240.244
R19082 GND.n7406 GND.n4437 240.244
R19083 GND.n7406 GND.n4438 240.244
R19084 GND.n7402 GND.n4438 240.244
R19085 GND.n7402 GND.n4446 240.244
R19086 GND.n7392 GND.n4446 240.244
R19087 GND.n7392 GND.n4458 240.244
R19088 GND.n7388 GND.n4458 240.244
R19089 GND.n7388 GND.n4464 240.244
R19090 GND.n7378 GND.n4464 240.244
R19091 GND.n7378 GND.n4476 240.244
R19092 GND.n7374 GND.n4476 240.244
R19093 GND.n7374 GND.n4482 240.244
R19094 GND.n7364 GND.n4482 240.244
R19095 GND.n7364 GND.n4494 240.244
R19096 GND.n7360 GND.n4494 240.244
R19097 GND.n7360 GND.n4500 240.244
R19098 GND.n7350 GND.n4500 240.244
R19099 GND.n7350 GND.n4512 240.244
R19100 GND.n7346 GND.n4512 240.244
R19101 GND.n7346 GND.n4518 240.244
R19102 GND.n7336 GND.n4518 240.244
R19103 GND.n7336 GND.n4530 240.244
R19104 GND.n7332 GND.n4530 240.244
R19105 GND.n7332 GND.n4536 240.244
R19106 GND.n4559 GND.n4536 240.244
R19107 GND.n7317 GND.n4559 240.244
R19108 GND.n7317 GND.n4560 240.244
R19109 GND.n7313 GND.n4560 240.244
R19110 GND.n7313 GND.n4568 240.244
R19111 GND.n7303 GND.n4568 240.244
R19112 GND.n7303 GND.n4580 240.244
R19113 GND.n7299 GND.n4580 240.244
R19114 GND.n7299 GND.n4586 240.244
R19115 GND.n7289 GND.n4586 240.244
R19116 GND.n7289 GND.n4598 240.244
R19117 GND.n7285 GND.n4598 240.244
R19118 GND.n7285 GND.n4604 240.244
R19119 GND.n7275 GND.n4604 240.244
R19120 GND.n7275 GND.n4615 240.244
R19121 GND.n7271 GND.n4615 240.244
R19122 GND.n7271 GND.n4621 240.244
R19123 GND.n4690 GND.n4621 240.244
R19124 GND.n7256 GND.n4690 240.244
R19125 GND.n7256 GND.n4691 240.244
R19126 GND.n7252 GND.n4691 240.244
R19127 GND.n7252 GND.n4699 240.244
R19128 GND.n6399 GND.n4699 240.244
R19129 GND.n6399 GND.n6393 240.244
R19130 GND.n6403 GND.n6393 240.244
R19131 GND.n6404 GND.n6403 240.244
R19132 GND.n6404 GND.n6388 240.244
R19133 GND.n6413 GND.n6388 240.244
R19134 GND.n6413 GND.n6389 240.244
R19135 GND.n6389 GND.n4897 240.244
R19136 GND.n7082 GND.n4897 240.244
R19137 GND.n7082 GND.n4898 240.244
R19138 GND.n7078 GND.n4898 240.244
R19139 GND.n7078 GND.n4904 240.244
R19140 GND.n6471 GND.n4904 240.244
R19141 GND.n6471 GND.n6432 240.244
R19142 GND.n6467 GND.n6432 240.244
R19143 GND.n6467 GND.n6466 240.244
R19144 GND.n6466 GND.n6465 240.244
R19145 GND.n6465 GND.n6438 240.244
R19146 GND.n6461 GND.n6438 240.244
R19147 GND.n6461 GND.n6460 240.244
R19148 GND.n6460 GND.n6459 240.244
R19149 GND.n6459 GND.n6444 240.244
R19150 GND.n6455 GND.n6444 240.244
R19151 GND.n6455 GND.n6454 240.244
R19152 GND.n6454 GND.n6453 240.244
R19153 GND.n6453 GND.n5329 240.244
R19154 GND.n6677 GND.n5329 240.244
R19155 GND.n6677 GND.n5325 240.244
R19156 GND.n6683 GND.n5325 240.244
R19157 GND.n6684 GND.n6683 240.244
R19158 GND.n6685 GND.n6684 240.244
R19159 GND.n6685 GND.n5321 240.244
R19160 GND.n6691 GND.n5321 240.244
R19161 GND.n6692 GND.n6691 240.244
R19162 GND.n6693 GND.n6692 240.244
R19163 GND.n6693 GND.n5317 240.244
R19164 GND.n6699 GND.n5317 240.244
R19165 GND.n6700 GND.n6699 240.244
R19166 GND.n6701 GND.n6700 240.244
R19167 GND.n6701 GND.n5313 240.244
R19168 GND.n6707 GND.n5313 240.244
R19169 GND.n6708 GND.n6707 240.244
R19170 GND.n6709 GND.n6708 240.244
R19171 GND.n6709 GND.n5309 240.244
R19172 GND.n6715 GND.n5309 240.244
R19173 GND.n6716 GND.n6715 240.244
R19174 GND.n6717 GND.n6716 240.244
R19175 GND.n6717 GND.n5305 240.244
R19176 GND.n6723 GND.n5305 240.244
R19177 GND.n6724 GND.n6723 240.244
R19178 GND.n6725 GND.n6724 240.244
R19179 GND.n6725 GND.n5301 240.244
R19180 GND.n6731 GND.n5301 240.244
R19181 GND.n6732 GND.n6731 240.244
R19182 GND.n6733 GND.n6732 240.244
R19183 GND.n6733 GND.n5297 240.244
R19184 GND.n6739 GND.n5297 240.244
R19185 GND.n6740 GND.n6739 240.244
R19186 GND.n6741 GND.n6740 240.244
R19187 GND.n6741 GND.n5292 240.244
R19188 GND.n6752 GND.n5292 240.244
R19189 GND.n6752 GND.n5293 240.244
R19190 GND.n6748 GND.n5293 240.244
R19191 GND.n6748 GND.n5193 240.244
R19192 GND.n6914 GND.n5193 240.244
R19193 GND.n6914 GND.n5194 240.244
R19194 GND.n6909 GND.n5194 240.244
R19195 GND.n6909 GND.n6908 240.244
R19196 GND.n6908 GND.n5197 240.244
R19197 GND.n6903 GND.n5197 240.244
R19198 GND.n6903 GND.n5266 240.244
R19199 GND.n5266 GND.n5265 240.244
R19200 GND.n5265 GND.n5199 240.244
R19201 GND.n5261 GND.n5199 240.244
R19202 GND.n5261 GND.n5260 240.244
R19203 GND.n5260 GND.n5259 240.244
R19204 GND.n5259 GND.n5204 240.244
R19205 GND.n5255 GND.n5204 240.244
R19206 GND.n5255 GND.n5254 240.244
R19207 GND.n5254 GND.n5253 240.244
R19208 GND.n5253 GND.n5210 240.244
R19209 GND.n5249 GND.n5210 240.244
R19210 GND.n5249 GND.n5248 240.244
R19211 GND.n5248 GND.n5247 240.244
R19212 GND.n5247 GND.n5216 240.244
R19213 GND.n5243 GND.n5216 240.244
R19214 GND.n5243 GND.n5242 240.244
R19215 GND.n5242 GND.n5241 240.244
R19216 GND.n5241 GND.n5222 240.244
R19217 GND.n5237 GND.n5222 240.244
R19218 GND.n5237 GND.n5236 240.244
R19219 GND.n5236 GND.n5235 240.244
R19220 GND.n5235 GND.n5228 240.244
R19221 GND.n5228 GND.n442 240.244
R19222 GND.n9725 GND.n442 240.244
R19223 GND.n9725 GND.n443 240.244
R19224 GND.n9721 GND.n443 240.244
R19225 GND.n9721 GND.n9720 240.244
R19226 GND.n9720 GND.n9719 240.244
R19227 GND.n9719 GND.n449 240.244
R19228 GND.n9715 GND.n449 240.244
R19229 GND.n9715 GND.n9714 240.244
R19230 GND.n9714 GND.n9713 240.244
R19231 GND.n9713 GND.n455 240.244
R19232 GND.n9709 GND.n455 240.244
R19233 GND.n9709 GND.n9708 240.244
R19234 GND.n9708 GND.n9707 240.244
R19235 GND.n9707 GND.n461 240.244
R19236 GND.n9703 GND.n461 240.244
R19237 GND.n9703 GND.n9702 240.244
R19238 GND.n9702 GND.n9701 240.244
R19239 GND.n9701 GND.n467 240.244
R19240 GND.n9697 GND.n467 240.244
R19241 GND.n9697 GND.n9696 240.244
R19242 GND.n8496 GND.n1189 240.244
R19243 GND.n8492 GND.n1189 240.244
R19244 GND.n8492 GND.n1194 240.244
R19245 GND.n8488 GND.n1194 240.244
R19246 GND.n8488 GND.n1196 240.244
R19247 GND.n8484 GND.n1196 240.244
R19248 GND.n8484 GND.n1202 240.244
R19249 GND.n8480 GND.n1202 240.244
R19250 GND.n8480 GND.n1204 240.244
R19251 GND.n8476 GND.n1204 240.244
R19252 GND.n8476 GND.n1210 240.244
R19253 GND.n8472 GND.n1210 240.244
R19254 GND.n8472 GND.n1212 240.244
R19255 GND.n8468 GND.n1212 240.244
R19256 GND.n8468 GND.n1218 240.244
R19257 GND.n8464 GND.n1218 240.244
R19258 GND.n8464 GND.n1220 240.244
R19259 GND.n8460 GND.n1220 240.244
R19260 GND.n8460 GND.n1226 240.244
R19261 GND.n8456 GND.n1226 240.244
R19262 GND.n8456 GND.n1228 240.244
R19263 GND.n8452 GND.n1228 240.244
R19264 GND.n8452 GND.n1234 240.244
R19265 GND.n8448 GND.n1234 240.244
R19266 GND.n8448 GND.n1236 240.244
R19267 GND.n8444 GND.n1236 240.244
R19268 GND.n8444 GND.n1242 240.244
R19269 GND.n8440 GND.n1242 240.244
R19270 GND.n8440 GND.n1244 240.244
R19271 GND.n8436 GND.n1244 240.244
R19272 GND.n8436 GND.n1250 240.244
R19273 GND.n8432 GND.n1250 240.244
R19274 GND.n8432 GND.n1252 240.244
R19275 GND.n8428 GND.n1252 240.244
R19276 GND.n8428 GND.n1258 240.244
R19277 GND.n8424 GND.n1258 240.244
R19278 GND.n8424 GND.n1260 240.244
R19279 GND.n8420 GND.n1260 240.244
R19280 GND.n8420 GND.n1266 240.244
R19281 GND.n8416 GND.n1266 240.244
R19282 GND.n8416 GND.n1268 240.244
R19283 GND.n8412 GND.n1268 240.244
R19284 GND.n8412 GND.n1274 240.244
R19285 GND.n8408 GND.n1274 240.244
R19286 GND.n8408 GND.n1276 240.244
R19287 GND.n8404 GND.n1276 240.244
R19288 GND.n8404 GND.n1282 240.244
R19289 GND.n8400 GND.n1282 240.244
R19290 GND.n8400 GND.n1284 240.244
R19291 GND.n8396 GND.n1284 240.244
R19292 GND.n8396 GND.n1290 240.244
R19293 GND.n8392 GND.n1290 240.244
R19294 GND.n8392 GND.n1292 240.244
R19295 GND.n8388 GND.n1292 240.244
R19296 GND.n8388 GND.n1298 240.244
R19297 GND.n8384 GND.n1298 240.244
R19298 GND.n8384 GND.n1300 240.244
R19299 GND.n8380 GND.n1300 240.244
R19300 GND.n8380 GND.n1306 240.244
R19301 GND.n8376 GND.n1306 240.244
R19302 GND.n8376 GND.n1308 240.244
R19303 GND.n8372 GND.n1308 240.244
R19304 GND.n8372 GND.n1314 240.244
R19305 GND.n8368 GND.n1314 240.244
R19306 GND.n8368 GND.n1316 240.244
R19307 GND.n8364 GND.n1316 240.244
R19308 GND.n2926 GND.n2925 240.244
R19309 GND.n2935 GND.n2925 240.244
R19310 GND.n2935 GND.n2914 240.244
R19311 GND.n2952 GND.n2914 240.244
R19312 GND.n2952 GND.n2915 240.244
R19313 GND.n2915 GND.n2905 240.244
R19314 GND.n2905 GND.n2894 240.244
R19315 GND.n2969 GND.n2894 240.244
R19316 GND.n2969 GND.n2895 240.244
R19317 GND.n2895 GND.n2885 240.244
R19318 GND.n2885 GND.n2876 240.244
R19319 GND.n2993 GND.n2876 240.244
R19320 GND.n2993 GND.n2877 240.244
R19321 GND.n2877 GND.n2865 240.244
R19322 GND.n2984 GND.n2865 240.244
R19323 GND.n2984 GND.n2851 240.244
R19324 GND.n3026 GND.n2851 240.244
R19325 GND.n3026 GND.n2852 240.244
R19326 GND.n2852 GND.n2842 240.244
R19327 GND.n2842 GND.n2826 240.244
R19328 GND.n3059 GND.n2826 240.244
R19329 GND.n3059 GND.n2827 240.244
R19330 GND.n2827 GND.n2817 240.244
R19331 GND.n3050 GND.n2817 240.244
R19332 GND.n3050 GND.n2798 240.244
R19333 GND.n3096 GND.n2798 240.244
R19334 GND.n3096 GND.n2799 240.244
R19335 GND.n2799 GND.n2788 240.244
R19336 GND.n3087 GND.n2788 240.244
R19337 GND.n3087 GND.n2769 240.244
R19338 GND.n3134 GND.n2769 240.244
R19339 GND.n3134 GND.n2770 240.244
R19340 GND.n2770 GND.n2758 240.244
R19341 GND.n3125 GND.n2758 240.244
R19342 GND.n3125 GND.n2741 240.244
R19343 GND.n3172 GND.n2741 240.244
R19344 GND.n3172 GND.n2742 240.244
R19345 GND.n2742 GND.n2731 240.244
R19346 GND.n3163 GND.n2731 240.244
R19347 GND.n3163 GND.n2712 240.244
R19348 GND.n3209 GND.n2712 240.244
R19349 GND.n3209 GND.n2713 240.244
R19350 GND.n2713 GND.n2702 240.244
R19351 GND.n3200 GND.n2702 240.244
R19352 GND.n3200 GND.n2683 240.244
R19353 GND.n3246 GND.n2683 240.244
R19354 GND.n3246 GND.n2684 240.244
R19355 GND.n2684 GND.n2673 240.244
R19356 GND.n3237 GND.n2673 240.244
R19357 GND.n3237 GND.n2654 240.244
R19358 GND.n3283 GND.n2654 240.244
R19359 GND.n3283 GND.n2655 240.244
R19360 GND.n2655 GND.n2643 240.244
R19361 GND.n3274 GND.n2643 240.244
R19362 GND.n3274 GND.n2625 240.244
R19363 GND.n3319 GND.n2625 240.244
R19364 GND.n3319 GND.n2626 240.244
R19365 GND.n2626 GND.n2619 240.244
R19366 GND.n2619 GND.n2608 240.244
R19367 GND.n3543 GND.n2608 240.244
R19368 GND.n3543 GND.n1536 240.244
R19369 GND.n2601 GND.n1536 240.244
R19370 GND.n3553 GND.n2601 240.244
R19371 GND.n3553 GND.n1556 240.244
R19372 GND.n8115 GND.n1556 240.244
R19373 GND.n8115 GND.n1557 240.244
R19374 GND.n3571 GND.n1557 240.244
R19375 GND.n3574 GND.n3571 240.244
R19376 GND.n3574 GND.n3573 240.244
R19377 GND.n3573 GND.n2575 240.244
R19378 GND.n2575 GND.n2564 240.244
R19379 GND.n3596 GND.n2564 240.244
R19380 GND.n3600 GND.n3596 240.244
R19381 GND.n3600 GND.n3599 240.244
R19382 GND.n3599 GND.n2552 240.244
R19383 GND.n2552 GND.n2543 240.244
R19384 GND.n3622 GND.n2543 240.244
R19385 GND.n3626 GND.n3622 240.244
R19386 GND.n3626 GND.n3624 240.244
R19387 GND.n3624 GND.n2532 240.244
R19388 GND.n2532 GND.n2521 240.244
R19389 GND.n3648 GND.n2521 240.244
R19390 GND.n3652 GND.n3648 240.244
R19391 GND.n3652 GND.n3651 240.244
R19392 GND.n3651 GND.n2510 240.244
R19393 GND.n2510 GND.n2501 240.244
R19394 GND.n3674 GND.n2501 240.244
R19395 GND.n3677 GND.n3674 240.244
R19396 GND.n3677 GND.n3676 240.244
R19397 GND.n3676 GND.n2488 240.244
R19398 GND.n2488 GND.n2477 240.244
R19399 GND.n3699 GND.n2477 240.244
R19400 GND.n3703 GND.n3699 240.244
R19401 GND.n3703 GND.n3702 240.244
R19402 GND.n3702 GND.n2465 240.244
R19403 GND.n2465 GND.n2456 240.244
R19404 GND.n3725 GND.n2456 240.244
R19405 GND.n3729 GND.n3725 240.244
R19406 GND.n3729 GND.n3727 240.244
R19407 GND.n3727 GND.n2446 240.244
R19408 GND.n2446 GND.n2436 240.244
R19409 GND.n3751 GND.n2436 240.244
R19410 GND.n3755 GND.n3751 240.244
R19411 GND.n3755 GND.n3754 240.244
R19412 GND.n3754 GND.n2425 240.244
R19413 GND.n2425 GND.n2416 240.244
R19414 GND.n3777 GND.n2416 240.244
R19415 GND.n3780 GND.n3777 240.244
R19416 GND.n3780 GND.n3779 240.244
R19417 GND.n3779 GND.n2403 240.244
R19418 GND.n2403 GND.n2392 240.244
R19419 GND.n3802 GND.n2392 240.244
R19420 GND.n3806 GND.n3802 240.244
R19421 GND.n3806 GND.n3805 240.244
R19422 GND.n3805 GND.n2380 240.244
R19423 GND.n2380 GND.n2371 240.244
R19424 GND.n3829 GND.n2371 240.244
R19425 GND.n3833 GND.n3829 240.244
R19426 GND.n3833 GND.n3831 240.244
R19427 GND.n3831 GND.n1680 240.244
R19428 GND.n8025 GND.n1680 240.244
R19429 GND.n1439 GND.n1359 240.244
R19430 GND.n1441 GND.n1440 240.244
R19431 GND.n1445 GND.n1444 240.244
R19432 GND.n1447 GND.n1446 240.244
R19433 GND.n1451 GND.n1450 240.244
R19434 GND.n8220 GND.n1357 240.244
R19435 GND.n1455 GND.n1454 240.244
R19436 GND.n1456 GND.n1455 240.244
R19437 GND.n2911 GND.n1456 240.244
R19438 GND.n2911 GND.n1459 240.244
R19439 GND.n1460 GND.n1459 240.244
R19440 GND.n1461 GND.n1460 240.244
R19441 GND.n2891 GND.n1461 240.244
R19442 GND.n2891 GND.n1464 240.244
R19443 GND.n1465 GND.n1464 240.244
R19444 GND.n1466 GND.n1465 240.244
R19445 GND.n2872 GND.n1466 240.244
R19446 GND.n2872 GND.n1469 240.244
R19447 GND.n1470 GND.n1469 240.244
R19448 GND.n1471 GND.n1470 240.244
R19449 GND.n2861 GND.n1471 240.244
R19450 GND.n2861 GND.n1474 240.244
R19451 GND.n1475 GND.n1474 240.244
R19452 GND.n1476 GND.n1475 240.244
R19453 GND.n2841 GND.n1476 240.244
R19454 GND.n2841 GND.n1479 240.244
R19455 GND.n1480 GND.n1479 240.244
R19456 GND.n1481 GND.n1480 240.244
R19457 GND.n2815 GND.n1481 240.244
R19458 GND.n2815 GND.n1484 240.244
R19459 GND.n1485 GND.n1484 240.244
R19460 GND.n1486 GND.n1485 240.244
R19461 GND.n2784 GND.n1486 240.244
R19462 GND.n2784 GND.n1489 240.244
R19463 GND.n1490 GND.n1489 240.244
R19464 GND.n1491 GND.n1490 240.244
R19465 GND.n2767 GND.n1491 240.244
R19466 GND.n2767 GND.n1494 240.244
R19467 GND.n1495 GND.n1494 240.244
R19468 GND.n1496 GND.n1495 240.244
R19469 GND.n3157 GND.n1496 240.244
R19470 GND.n3157 GND.n1499 240.244
R19471 GND.n1500 GND.n1499 240.244
R19472 GND.n1501 GND.n1500 240.244
R19473 GND.n2720 GND.n1501 240.244
R19474 GND.n2720 GND.n1504 240.244
R19475 GND.n1505 GND.n1504 240.244
R19476 GND.n1506 GND.n1505 240.244
R19477 GND.n2700 GND.n1506 240.244
R19478 GND.n2700 GND.n1509 240.244
R19479 GND.n1510 GND.n1509 240.244
R19480 GND.n1511 GND.n1510 240.244
R19481 GND.n2669 GND.n1511 240.244
R19482 GND.n2669 GND.n1514 240.244
R19483 GND.n1515 GND.n1514 240.244
R19484 GND.n1516 GND.n1515 240.244
R19485 GND.n2652 GND.n1516 240.244
R19486 GND.n2652 GND.n1519 240.244
R19487 GND.n1520 GND.n1519 240.244
R19488 GND.n1521 GND.n1520 240.244
R19489 GND.n3307 GND.n1521 240.244
R19490 GND.n3307 GND.n1524 240.244
R19491 GND.n1525 GND.n1524 240.244
R19492 GND.n1526 GND.n1525 240.244
R19493 GND.n2609 GND.n1526 240.244
R19494 GND.n2609 GND.n1529 240.244
R19495 GND.n8124 GND.n1529 240.244
R19496 GND.n8124 GND.n1532 240.244
R19497 GND.n2595 GND.n1532 240.244
R19498 GND.n3560 GND.n2595 240.244
R19499 GND.n3560 GND.n1554 240.244
R19500 GND.n2589 GND.n1554 240.244
R19501 GND.n3569 GND.n2589 240.244
R19502 GND.n3569 GND.n2585 240.244
R19503 GND.n2585 GND.n2571 240.244
R19504 GND.n3586 GND.n2571 240.244
R19505 GND.n3586 GND.n2567 240.244
R19506 GND.n3594 GND.n2567 240.244
R19507 GND.n3594 GND.n2562 240.244
R19508 GND.n2562 GND.n2549 240.244
R19509 GND.n3612 GND.n2549 240.244
R19510 GND.n3612 GND.n2545 240.244
R19511 GND.n3620 GND.n2545 240.244
R19512 GND.n3620 GND.n2541 240.244
R19513 GND.n2541 GND.n2528 240.244
R19514 GND.n3638 GND.n2528 240.244
R19515 GND.n3638 GND.n2524 240.244
R19516 GND.n3646 GND.n2524 240.244
R19517 GND.n3646 GND.n2519 240.244
R19518 GND.n2519 GND.n2507 240.244
R19519 GND.n3664 GND.n2507 240.244
R19520 GND.n3664 GND.n2503 240.244
R19521 GND.n3672 GND.n2503 240.244
R19522 GND.n3672 GND.n2498 240.244
R19523 GND.n2498 GND.n2484 240.244
R19524 GND.n3689 GND.n2484 240.244
R19525 GND.n3689 GND.n2480 240.244
R19526 GND.n3697 GND.n2480 240.244
R19527 GND.n3697 GND.n2475 240.244
R19528 GND.n2475 GND.n2462 240.244
R19529 GND.n3715 GND.n2462 240.244
R19530 GND.n3715 GND.n2458 240.244
R19531 GND.n3723 GND.n2458 240.244
R19532 GND.n3723 GND.n2454 240.244
R19533 GND.n2454 GND.n2443 240.244
R19534 GND.n3741 GND.n2443 240.244
R19535 GND.n3741 GND.n2439 240.244
R19536 GND.n3749 GND.n2439 240.244
R19537 GND.n3749 GND.n2434 240.244
R19538 GND.n2434 GND.n2422 240.244
R19539 GND.n3767 GND.n2422 240.244
R19540 GND.n3767 GND.n2418 240.244
R19541 GND.n3775 GND.n2418 240.244
R19542 GND.n3775 GND.n2413 240.244
R19543 GND.n2413 GND.n2399 240.244
R19544 GND.n3792 GND.n2399 240.244
R19545 GND.n3792 GND.n2395 240.244
R19546 GND.n3800 GND.n2395 240.244
R19547 GND.n3800 GND.n2390 240.244
R19548 GND.n2390 GND.n2377 240.244
R19549 GND.n3818 GND.n2377 240.244
R19550 GND.n3818 GND.n2373 240.244
R19551 GND.n3827 GND.n2373 240.244
R19552 GND.n3827 GND.n2369 240.244
R19553 GND.n2369 GND.n2361 240.244
R19554 GND.n3844 GND.n2361 240.244
R19555 GND.n3844 GND.n1678 240.244
R19556 GND.n8024 GND.n1681 240.244
R19557 GND.n3858 GND.n3857 240.244
R19558 GND.n3862 GND.n3861 240.244
R19559 GND.n3866 GND.n3865 240.244
R19560 GND.n3870 GND.n3869 240.244
R19561 GND.n3854 GND.n1706 240.244
R19562 GND.n1917 GND.n1916 240.132
R19563 GND.n4749 GND.n4748 240.132
R19564 GND.n7916 GND.t96 235.065
R19565 GND.n2121 GND.t142 235.065
R19566 GND.n4760 GND.t25 235.065
R19567 GND.n4758 GND.t106 235.065
R19568 GND.n8221 GND.t145 223.448
R19569 GND.n1738 GND.t57 223.448
R19570 GND.n1759 GND.t115 223.448
R19571 GND.n1776 GND.t81 223.448
R19572 GND.n1797 GND.t21 223.448
R19573 GND.n1817 GND.t139 223.448
R19574 GND.n7108 GND.t109 223.448
R19575 GND.n7122 GND.t44 223.448
R19576 GND.n5391 GND.t136 223.448
R19577 GND.n5424 GND.t75 223.448
R19578 GND.n5458 GND.t133 223.448
R19579 GND.n9843 GND.t118 223.448
R19580 GND.n9999 GND.t66 223.448
R19581 GND.n9859 GND.t130 223.448
R19582 GND.n9869 GND.t29 223.448
R19583 GND.n9877 GND.t93 223.448
R19584 GND.n9808 GND.t37 223.448
R19585 GND.n6359 GND.t54 223.448
R19586 GND.n1375 GND.t72 223.448
R19587 GND.n1389 GND.t121 223.448
R19588 GND.n1405 GND.t84 223.448
R19589 GND.n1419 GND.t33 223.448
R19590 GND.n1435 GND.t100 223.448
R19591 GND.n3852 GND.t63 223.448
R19592 GND.n4852 GND.n4834 199.319
R19593 GND.n7184 GND.n4834 199.319
R19594 GND.n1870 GND.n1708 199.319
R19595 GND.n1918 GND.n1914 186.49
R19596 GND.n4750 GND.n4746 186.49
R19597 GND.n5391 GND.t138 173.85
R19598 GND.n5424 GND.t77 173.85
R19599 GND.n9843 GND.t119 173.85
R19600 GND.n9999 GND.t67 173.85
R19601 GND.n8221 GND.t147 164.25
R19602 GND.n1738 GND.t58 164.25
R19603 GND.n1759 GND.t116 164.25
R19604 GND.n1776 GND.t82 164.25
R19605 GND.n1797 GND.t23 164.25
R19606 GND.n1817 GND.t140 164.25
R19607 GND.n7108 GND.t111 164.25
R19608 GND.n7122 GND.t47 164.25
R19609 GND.n5458 GND.t135 164.25
R19610 GND.n9859 GND.t131 164.25
R19611 GND.n9869 GND.t31 164.25
R19612 GND.n9877 GND.t94 164.25
R19613 GND.n9808 GND.t38 164.25
R19614 GND.n6359 GND.t56 164.25
R19615 GND.n1375 GND.t74 164.25
R19616 GND.n1389 GND.t123 164.25
R19617 GND.n1405 GND.t86 164.25
R19618 GND.n1419 GND.t36 164.25
R19619 GND.n1435 GND.t102 164.25
R19620 GND.n3852 GND.t64 164.25
R19621 GND.n7248 GND.n4732 163.367
R19622 GND.n7244 GND.n7243 163.367
R19623 GND.n7240 GND.n7239 163.367
R19624 GND.n7236 GND.n7235 163.367
R19625 GND.n7232 GND.n7231 163.367
R19626 GND.n7228 GND.n7227 163.367
R19627 GND.n7224 GND.n7223 163.367
R19628 GND.n7220 GND.n7219 163.367
R19629 GND.n7216 GND.n7215 163.367
R19630 GND.n7212 GND.n7211 163.367
R19631 GND.n7208 GND.n7207 163.367
R19632 GND.n7204 GND.n7203 163.367
R19633 GND.n7200 GND.n7199 163.367
R19634 GND.n7195 GND.n7194 163.367
R19635 GND.n7191 GND.n7190 163.367
R19636 GND.n4831 GND.n4830 163.367
R19637 GND.n4827 GND.n4826 163.367
R19638 GND.n4823 GND.n4822 163.367
R19639 GND.n4819 GND.n4818 163.367
R19640 GND.n4815 GND.n4814 163.367
R19641 GND.n4811 GND.n4810 163.367
R19642 GND.n4807 GND.n4806 163.367
R19643 GND.n4803 GND.n4802 163.367
R19644 GND.n4799 GND.n4798 163.367
R19645 GND.n4795 GND.n4794 163.367
R19646 GND.n4791 GND.n4790 163.367
R19647 GND.n4787 GND.n4786 163.367
R19648 GND.n4783 GND.n4782 163.367
R19649 GND.n4779 GND.n4778 163.367
R19650 GND.n2181 GND.n1937 163.367
R19651 GND.n2185 GND.n1937 163.367
R19652 GND.n2191 GND.n2185 163.367
R19653 GND.n2192 GND.n2191 163.367
R19654 GND.n2192 GND.n1948 163.367
R19655 GND.n2196 GND.n1948 163.367
R19656 GND.n2196 GND.n1956 163.367
R19657 GND.n2200 GND.n1956 163.367
R19658 GND.n2203 GND.n2200 163.367
R19659 GND.n2203 GND.n1964 163.367
R19660 GND.n2206 GND.n1964 163.367
R19661 GND.n2206 GND.n1972 163.367
R19662 GND.n2210 GND.n1972 163.367
R19663 GND.n2215 GND.n2210 163.367
R19664 GND.n2216 GND.n2215 163.367
R19665 GND.n2216 GND.n1982 163.367
R19666 GND.n2219 GND.n1982 163.367
R19667 GND.n2219 GND.n1990 163.367
R19668 GND.n2223 GND.n1990 163.367
R19669 GND.n2228 GND.n2223 163.367
R19670 GND.n2229 GND.n2228 163.367
R19671 GND.n2229 GND.n2000 163.367
R19672 GND.n2232 GND.n2000 163.367
R19673 GND.n2232 GND.n2008 163.367
R19674 GND.n2236 GND.n2008 163.367
R19675 GND.n2241 GND.n2236 163.367
R19676 GND.n2242 GND.n2241 163.367
R19677 GND.n2242 GND.n2018 163.367
R19678 GND.n2245 GND.n2018 163.367
R19679 GND.n2245 GND.n2026 163.367
R19680 GND.n2249 GND.n2026 163.367
R19681 GND.n2253 GND.n2249 163.367
R19682 GND.n2254 GND.n2253 163.367
R19683 GND.n2254 GND.n2036 163.367
R19684 GND.n2257 GND.n2036 163.367
R19685 GND.n2257 GND.n2044 163.367
R19686 GND.n2261 GND.n2044 163.367
R19687 GND.n2266 GND.n2261 163.367
R19688 GND.n2267 GND.n2266 163.367
R19689 GND.n2267 GND.n2054 163.367
R19690 GND.n2270 GND.n2054 163.367
R19691 GND.n2270 GND.n2062 163.367
R19692 GND.n2274 GND.n2062 163.367
R19693 GND.n2279 GND.n2274 163.367
R19694 GND.n2280 GND.n2279 163.367
R19695 GND.n2280 GND.n2072 163.367
R19696 GND.n2283 GND.n2072 163.367
R19697 GND.n2283 GND.n2080 163.367
R19698 GND.n2287 GND.n2080 163.367
R19699 GND.n2292 GND.n2287 163.367
R19700 GND.n2293 GND.n2292 163.367
R19701 GND.n2293 GND.n2090 163.367
R19702 GND.n2296 GND.n2090 163.367
R19703 GND.n2296 GND.n2098 163.367
R19704 GND.n2299 GND.n2098 163.367
R19705 GND.n2299 GND.n2111 163.367
R19706 GND.n7778 GND.n2111 163.367
R19707 GND.n7778 GND.n2112 163.367
R19708 GND.n7774 GND.n2112 163.367
R19709 GND.n7774 GND.n2303 163.367
R19710 GND.n2315 GND.n2303 163.367
R19711 GND.n5695 GND.n2315 163.367
R19712 GND.n5702 GND.n5695 163.367
R19713 GND.n5702 GND.n5696 163.367
R19714 GND.n5696 GND.n5689 163.367
R19715 GND.n5713 GND.n5689 163.367
R19716 GND.n5714 GND.n5713 163.367
R19717 GND.n5714 GND.n5686 163.367
R19718 GND.n5720 GND.n5686 163.367
R19719 GND.n5720 GND.n5687 163.367
R19720 GND.n5687 GND.n5663 163.367
R19721 GND.n5731 GND.n5663 163.367
R19722 GND.n5732 GND.n5731 163.367
R19723 GND.n5732 GND.n5660 163.367
R19724 GND.n5744 GND.n5660 163.367
R19725 GND.n5744 GND.n5661 163.367
R19726 GND.n5740 GND.n5661 163.367
R19727 GND.n5740 GND.n5654 163.367
R19728 GND.n5737 GND.n5654 163.367
R19729 GND.n5737 GND.n5736 163.367
R19730 GND.n5736 GND.n3938 163.367
R19731 GND.n7667 GND.n3938 163.367
R19732 GND.n7667 GND.n3939 163.367
R19733 GND.n7663 GND.n3939 163.367
R19734 GND.n7663 GND.n3942 163.367
R19735 GND.n3951 GND.n3942 163.367
R19736 GND.n5799 GND.n3951 163.367
R19737 GND.n5806 GND.n5799 163.367
R19738 GND.n5806 GND.n5800 163.367
R19739 GND.n5800 GND.n5642 163.367
R19740 GND.n5817 GND.n5642 163.367
R19741 GND.n5818 GND.n5817 163.367
R19742 GND.n5818 GND.n5639 163.367
R19743 GND.n5824 GND.n5639 163.367
R19744 GND.n5824 GND.n5640 163.367
R19745 GND.n5640 GND.n5632 163.367
R19746 GND.n5835 GND.n5632 163.367
R19747 GND.n5836 GND.n5835 163.367
R19748 GND.n5836 GND.n5629 163.367
R19749 GND.n5848 GND.n5629 163.367
R19750 GND.n5848 GND.n5630 163.367
R19751 GND.n5844 GND.n5630 163.367
R19752 GND.n5844 GND.n5623 163.367
R19753 GND.n5841 GND.n5623 163.367
R19754 GND.n5841 GND.n5840 163.367
R19755 GND.n5840 GND.n4042 163.367
R19756 GND.n7612 GND.n4042 163.367
R19757 GND.n7612 GND.n4043 163.367
R19758 GND.n7608 GND.n4043 163.367
R19759 GND.n7608 GND.n4046 163.367
R19760 GND.n4055 GND.n4046 163.367
R19761 GND.n5902 GND.n4055 163.367
R19762 GND.n5909 GND.n5902 163.367
R19763 GND.n5909 GND.n5903 163.367
R19764 GND.n5903 GND.n5611 163.367
R19765 GND.n5920 GND.n5611 163.367
R19766 GND.n5921 GND.n5920 163.367
R19767 GND.n5921 GND.n5608 163.367
R19768 GND.n5927 GND.n5608 163.367
R19769 GND.n5927 GND.n5609 163.367
R19770 GND.n5609 GND.n5601 163.367
R19771 GND.n5938 GND.n5601 163.367
R19772 GND.n5939 GND.n5938 163.367
R19773 GND.n5939 GND.n5598 163.367
R19774 GND.n5951 GND.n5598 163.367
R19775 GND.n5951 GND.n5599 163.367
R19776 GND.n5947 GND.n5599 163.367
R19777 GND.n5947 GND.n5592 163.367
R19778 GND.n5944 GND.n5592 163.367
R19779 GND.n5944 GND.n5943 163.367
R19780 GND.n5943 GND.n4147 163.367
R19781 GND.n7557 GND.n4147 163.367
R19782 GND.n7557 GND.n4148 163.367
R19783 GND.n7553 GND.n4148 163.367
R19784 GND.n7553 GND.n4151 163.367
R19785 GND.n4160 GND.n4151 163.367
R19786 GND.n6005 GND.n4160 163.367
R19787 GND.n6012 GND.n6005 163.367
R19788 GND.n6012 GND.n6006 163.367
R19789 GND.n6006 GND.n5580 163.367
R19790 GND.n6023 GND.n5580 163.367
R19791 GND.n6024 GND.n6023 163.367
R19792 GND.n6024 GND.n5577 163.367
R19793 GND.n6030 GND.n5577 163.367
R19794 GND.n6030 GND.n5578 163.367
R19795 GND.n5578 GND.n5569 163.367
R19796 GND.n6041 GND.n5569 163.367
R19797 GND.n6042 GND.n6041 163.367
R19798 GND.n6042 GND.n5566 163.367
R19799 GND.n6054 GND.n5566 163.367
R19800 GND.n6054 GND.n5567 163.367
R19801 GND.n6050 GND.n5567 163.367
R19802 GND.n6050 GND.n5560 163.367
R19803 GND.n6047 GND.n5560 163.367
R19804 GND.n6047 GND.n6046 163.367
R19805 GND.n6046 GND.n4250 163.367
R19806 GND.n7502 GND.n4250 163.367
R19807 GND.n7502 GND.n4251 163.367
R19808 GND.n7498 GND.n4251 163.367
R19809 GND.n7498 GND.n4254 163.367
R19810 GND.n4263 GND.n4254 163.367
R19811 GND.n6108 GND.n4263 163.367
R19812 GND.n6115 GND.n6108 163.367
R19813 GND.n6115 GND.n6109 163.367
R19814 GND.n6109 GND.n5546 163.367
R19815 GND.n6126 GND.n5546 163.367
R19816 GND.n6127 GND.n6126 163.367
R19817 GND.n6127 GND.n5543 163.367
R19818 GND.n6133 GND.n5543 163.367
R19819 GND.n6133 GND.n5544 163.367
R19820 GND.n5544 GND.n5536 163.367
R19821 GND.n6144 GND.n5536 163.367
R19822 GND.n6145 GND.n6144 163.367
R19823 GND.n6145 GND.n5533 163.367
R19824 GND.n6157 GND.n5533 163.367
R19825 GND.n6157 GND.n5534 163.367
R19826 GND.n6153 GND.n5534 163.367
R19827 GND.n6153 GND.n5527 163.367
R19828 GND.n6150 GND.n5527 163.367
R19829 GND.n6150 GND.n6149 163.367
R19830 GND.n6149 GND.n4354 163.367
R19831 GND.n7447 GND.n4354 163.367
R19832 GND.n7447 GND.n4355 163.367
R19833 GND.n7443 GND.n4355 163.367
R19834 GND.n7443 GND.n4358 163.367
R19835 GND.n4367 GND.n4358 163.367
R19836 GND.n5519 GND.n4367 163.367
R19837 GND.n6210 GND.n5519 163.367
R19838 GND.n6211 GND.n6210 163.367
R19839 GND.n6211 GND.n5514 163.367
R19840 GND.n6219 GND.n5514 163.367
R19841 GND.n6219 GND.n5515 163.367
R19842 GND.n6215 GND.n5515 163.367
R19843 GND.n6215 GND.n5508 163.367
R19844 GND.n6229 GND.n5508 163.367
R19845 GND.n6230 GND.n6229 163.367
R19846 GND.n6230 GND.n5497 163.367
R19847 GND.n6234 GND.n5497 163.367
R19848 GND.n6235 GND.n6234 163.367
R19849 GND.n6235 GND.n5505 163.367
R19850 GND.n6301 GND.n5505 163.367
R19851 GND.n6301 GND.n5506 163.367
R19852 GND.n5506 GND.n4448 163.367
R19853 GND.n6296 GND.n4448 163.367
R19854 GND.n6296 GND.n4456 163.367
R19855 GND.n6293 GND.n4456 163.367
R19856 GND.n6293 GND.n6292 163.367
R19857 GND.n6292 GND.n6288 163.367
R19858 GND.n6288 GND.n4466 163.367
R19859 GND.n6284 GND.n4466 163.367
R19860 GND.n6284 GND.n4474 163.367
R19861 GND.n6281 GND.n4474 163.367
R19862 GND.n6281 GND.n6280 163.367
R19863 GND.n6280 GND.n6275 163.367
R19864 GND.n6275 GND.n4484 163.367
R19865 GND.n6271 GND.n4484 163.367
R19866 GND.n6271 GND.n4492 163.367
R19867 GND.n6268 GND.n4492 163.367
R19868 GND.n6268 GND.n6267 163.367
R19869 GND.n6267 GND.n6262 163.367
R19870 GND.n6262 GND.n4502 163.367
R19871 GND.n6258 GND.n4502 163.367
R19872 GND.n6258 GND.n4510 163.367
R19873 GND.n6255 GND.n4510 163.367
R19874 GND.n6255 GND.n6254 163.367
R19875 GND.n6254 GND.n6249 163.367
R19876 GND.n6249 GND.n4520 163.367
R19877 GND.n6245 GND.n4520 163.367
R19878 GND.n6245 GND.n4528 163.367
R19879 GND.n6242 GND.n4528 163.367
R19880 GND.n6242 GND.n4541 163.367
R19881 GND.n7330 GND.n4541 163.367
R19882 GND.n7330 GND.n4542 163.367
R19883 GND.n7326 GND.n4542 163.367
R19884 GND.n7326 GND.n4545 163.367
R19885 GND.n4557 GND.n4545 163.367
R19886 GND.n4631 GND.n4557 163.367
R19887 GND.n4636 GND.n4631 163.367
R19888 GND.n4637 GND.n4636 163.367
R19889 GND.n4637 GND.n4570 163.367
R19890 GND.n4640 GND.n4570 163.367
R19891 GND.n4640 GND.n4578 163.367
R19892 GND.n4644 GND.n4578 163.367
R19893 GND.n4649 GND.n4644 163.367
R19894 GND.n4650 GND.n4649 163.367
R19895 GND.n4650 GND.n4588 163.367
R19896 GND.n4653 GND.n4588 163.367
R19897 GND.n4653 GND.n4596 163.367
R19898 GND.n4657 GND.n4596 163.367
R19899 GND.n4662 GND.n4657 163.367
R19900 GND.n4663 GND.n4662 163.367
R19901 GND.n4663 GND.n4606 163.367
R19902 GND.n4667 GND.n4606 163.367
R19903 GND.n4667 GND.n4613 163.367
R19904 GND.n4670 GND.n4613 163.367
R19905 GND.n4670 GND.n4624 163.367
R19906 GND.n7269 GND.n4624 163.367
R19907 GND.n7269 GND.n4625 163.367
R19908 GND.n7265 GND.n4625 163.367
R19909 GND.n7265 GND.n4674 163.367
R19910 GND.n4688 GND.n4674 163.367
R19911 GND.n4764 GND.n4688 163.367
R19912 GND.n4773 GND.n4764 163.367
R19913 GND.n4774 GND.n4773 163.367
R19914 GND.n1907 GND.n1906 163.367
R19915 GND.n7965 GND.n1906 163.367
R19916 GND.n7963 GND.n7962 163.367
R19917 GND.n7959 GND.n7958 163.367
R19918 GND.n7955 GND.n7954 163.367
R19919 GND.n7951 GND.n7950 163.367
R19920 GND.n7947 GND.n7946 163.367
R19921 GND.n7943 GND.n7942 163.367
R19922 GND.n7939 GND.n7938 163.367
R19923 GND.n7935 GND.n7934 163.367
R19924 GND.n7931 GND.n7930 163.367
R19925 GND.n7927 GND.n7926 163.367
R19926 GND.n7923 GND.n7922 163.367
R19927 GND.n7918 GND.n1875 163.367
R19928 GND.n7974 GND.n1873 163.367
R19929 GND.n2125 GND.n2124 163.367
R19930 GND.n2129 GND.n2128 163.367
R19931 GND.n2133 GND.n2132 163.367
R19932 GND.n2137 GND.n2136 163.367
R19933 GND.n2141 GND.n2140 163.367
R19934 GND.n2145 GND.n2144 163.367
R19935 GND.n2149 GND.n2148 163.367
R19936 GND.n2153 GND.n2152 163.367
R19937 GND.n2157 GND.n2156 163.367
R19938 GND.n2161 GND.n2160 163.367
R19939 GND.n2165 GND.n2164 163.367
R19940 GND.n2169 GND.n2168 163.367
R19941 GND.n2173 GND.n2172 163.367
R19942 GND.n2177 GND.n2176 163.367
R19943 GND.n7912 GND.n1908 163.367
R19944 GND.n7912 GND.n1935 163.367
R19945 GND.n2189 GND.n1935 163.367
R19946 GND.n2189 GND.n1950 163.367
R19947 GND.n7902 GND.n1950 163.367
R19948 GND.n7902 GND.n1951 163.367
R19949 GND.n7898 GND.n1951 163.367
R19950 GND.n7898 GND.n1954 163.367
R19951 GND.n1966 GND.n1954 163.367
R19952 GND.n7889 GND.n1966 163.367
R19953 GND.n7889 GND.n1967 163.367
R19954 GND.n7885 GND.n1967 163.367
R19955 GND.n7885 GND.n1970 163.367
R19956 GND.n2213 GND.n1970 163.367
R19957 GND.n2213 GND.n1984 163.367
R19958 GND.n7875 GND.n1984 163.367
R19959 GND.n7875 GND.n1985 163.367
R19960 GND.n7871 GND.n1985 163.367
R19961 GND.n7871 GND.n1988 163.367
R19962 GND.n2226 GND.n1988 163.367
R19963 GND.n2226 GND.n2002 163.367
R19964 GND.n7861 GND.n2002 163.367
R19965 GND.n7861 GND.n2003 163.367
R19966 GND.n7857 GND.n2003 163.367
R19967 GND.n7857 GND.n2006 163.367
R19968 GND.n2239 GND.n2006 163.367
R19969 GND.n2239 GND.n2020 163.367
R19970 GND.n7847 GND.n2020 163.367
R19971 GND.n7847 GND.n2021 163.367
R19972 GND.n7843 GND.n2021 163.367
R19973 GND.n7843 GND.n2024 163.367
R19974 GND.n2251 GND.n2024 163.367
R19975 GND.n2251 GND.n2038 163.367
R19976 GND.n7833 GND.n2038 163.367
R19977 GND.n7833 GND.n2039 163.367
R19978 GND.n7829 GND.n2039 163.367
R19979 GND.n7829 GND.n2042 163.367
R19980 GND.n2264 GND.n2042 163.367
R19981 GND.n2264 GND.n2056 163.367
R19982 GND.n7819 GND.n2056 163.367
R19983 GND.n7819 GND.n2057 163.367
R19984 GND.n7815 GND.n2057 163.367
R19985 GND.n7815 GND.n2060 163.367
R19986 GND.n2277 GND.n2060 163.367
R19987 GND.n2277 GND.n2074 163.367
R19988 GND.n7805 GND.n2074 163.367
R19989 GND.n7805 GND.n2075 163.367
R19990 GND.n7801 GND.n2075 163.367
R19991 GND.n7801 GND.n2078 163.367
R19992 GND.n2290 GND.n2078 163.367
R19993 GND.n2290 GND.n2092 163.367
R19994 GND.n7791 GND.n2092 163.367
R19995 GND.n7791 GND.n2093 163.367
R19996 GND.n7787 GND.n2093 163.367
R19997 GND.n7787 GND.n2096 163.367
R19998 GND.n2308 GND.n2096 163.367
R19999 GND.n2308 GND.n2109 163.367
R20000 GND.n2306 GND.n2109 163.367
R20001 GND.n7772 GND.n2306 163.367
R20002 GND.n7772 GND.n2307 163.367
R20003 GND.n7768 GND.n2307 163.367
R20004 GND.n7768 GND.n2313 163.367
R20005 GND.n5704 GND.n2313 163.367
R20006 GND.n5705 GND.n5704 163.367
R20007 GND.n5705 GND.n5691 163.367
R20008 GND.n5711 GND.n5691 163.367
R20009 GND.n5711 GND.n5692 163.367
R20010 GND.n5692 GND.n5668 163.367
R20011 GND.n5722 GND.n5668 163.367
R20012 GND.n5723 GND.n5722 163.367
R20013 GND.n5723 GND.n5665 163.367
R20014 GND.n5729 GND.n5665 163.367
R20015 GND.n5729 GND.n5666 163.367
R20016 GND.n5666 GND.n5658 163.367
R20017 GND.n5746 GND.n5658 163.367
R20018 GND.n5747 GND.n5746 163.367
R20019 GND.n5747 GND.n5655 163.367
R20020 GND.n5757 GND.n5655 163.367
R20021 GND.n5757 GND.n5656 163.367
R20022 GND.n5753 GND.n5656 163.367
R20023 GND.n5753 GND.n5752 163.367
R20024 GND.n5752 GND.n3934 163.367
R20025 GND.n3945 GND.n3934 163.367
R20026 GND.n7661 GND.n3945 163.367
R20027 GND.n7661 GND.n3946 163.367
R20028 GND.n7657 GND.n3946 163.367
R20029 GND.n7657 GND.n3949 163.367
R20030 GND.n5808 GND.n3949 163.367
R20031 GND.n5809 GND.n5808 163.367
R20032 GND.n5809 GND.n5644 163.367
R20033 GND.n5815 GND.n5644 163.367
R20034 GND.n5815 GND.n5645 163.367
R20035 GND.n5645 GND.n5637 163.367
R20036 GND.n5826 GND.n5637 163.367
R20037 GND.n5827 GND.n5826 163.367
R20038 GND.n5827 GND.n5634 163.367
R20039 GND.n5833 GND.n5634 163.367
R20040 GND.n5833 GND.n5635 163.367
R20041 GND.n5635 GND.n5627 163.367
R20042 GND.n5850 GND.n5627 163.367
R20043 GND.n5851 GND.n5850 163.367
R20044 GND.n5851 GND.n5624 163.367
R20045 GND.n5861 GND.n5624 163.367
R20046 GND.n5861 GND.n5625 163.367
R20047 GND.n5857 GND.n5625 163.367
R20048 GND.n5857 GND.n5856 163.367
R20049 GND.n5856 GND.n4038 163.367
R20050 GND.n4049 GND.n4038 163.367
R20051 GND.n7606 GND.n4049 163.367
R20052 GND.n7606 GND.n4050 163.367
R20053 GND.n7602 GND.n4050 163.367
R20054 GND.n7602 GND.n4053 163.367
R20055 GND.n5911 GND.n4053 163.367
R20056 GND.n5912 GND.n5911 163.367
R20057 GND.n5912 GND.n5613 163.367
R20058 GND.n5918 GND.n5613 163.367
R20059 GND.n5918 GND.n5614 163.367
R20060 GND.n5614 GND.n5606 163.367
R20061 GND.n5929 GND.n5606 163.367
R20062 GND.n5930 GND.n5929 163.367
R20063 GND.n5930 GND.n5603 163.367
R20064 GND.n5936 GND.n5603 163.367
R20065 GND.n5936 GND.n5604 163.367
R20066 GND.n5604 GND.n5596 163.367
R20067 GND.n5953 GND.n5596 163.367
R20068 GND.n5954 GND.n5953 163.367
R20069 GND.n5954 GND.n5593 163.367
R20070 GND.n5964 GND.n5593 163.367
R20071 GND.n5964 GND.n5594 163.367
R20072 GND.n5960 GND.n5594 163.367
R20073 GND.n5960 GND.n5959 163.367
R20074 GND.n5959 GND.n4143 163.367
R20075 GND.n4154 GND.n4143 163.367
R20076 GND.n7551 GND.n4154 163.367
R20077 GND.n7551 GND.n4155 163.367
R20078 GND.n7547 GND.n4155 163.367
R20079 GND.n7547 GND.n4158 163.367
R20080 GND.n6014 GND.n4158 163.367
R20081 GND.n6015 GND.n6014 163.367
R20082 GND.n6015 GND.n5582 163.367
R20083 GND.n6021 GND.n5582 163.367
R20084 GND.n6021 GND.n5583 163.367
R20085 GND.n5583 GND.n5574 163.367
R20086 GND.n6032 GND.n5574 163.367
R20087 GND.n6033 GND.n6032 163.367
R20088 GND.n6033 GND.n5571 163.367
R20089 GND.n6039 GND.n5571 163.367
R20090 GND.n6039 GND.n5572 163.367
R20091 GND.n5572 GND.n5564 163.367
R20092 GND.n6056 GND.n5564 163.367
R20093 GND.n6057 GND.n6056 163.367
R20094 GND.n6057 GND.n5561 163.367
R20095 GND.n6067 GND.n5561 163.367
R20096 GND.n6067 GND.n5562 163.367
R20097 GND.n6063 GND.n5562 163.367
R20098 GND.n6063 GND.n6062 163.367
R20099 GND.n6062 GND.n4246 163.367
R20100 GND.n4257 GND.n4246 163.367
R20101 GND.n7496 GND.n4257 163.367
R20102 GND.n7496 GND.n4258 163.367
R20103 GND.n7492 GND.n4258 163.367
R20104 GND.n7492 GND.n4261 163.367
R20105 GND.n6117 GND.n4261 163.367
R20106 GND.n6118 GND.n6117 163.367
R20107 GND.n6118 GND.n5549 163.367
R20108 GND.n6124 GND.n5549 163.367
R20109 GND.n6124 GND.n5550 163.367
R20110 GND.n5550 GND.n5541 163.367
R20111 GND.n6135 GND.n5541 163.367
R20112 GND.n6136 GND.n6135 163.367
R20113 GND.n6136 GND.n5538 163.367
R20114 GND.n6142 GND.n5538 163.367
R20115 GND.n6142 GND.n5539 163.367
R20116 GND.n5539 GND.n5531 163.367
R20117 GND.n6159 GND.n5531 163.367
R20118 GND.n6160 GND.n6159 163.367
R20119 GND.n6160 GND.n5528 163.367
R20120 GND.n6170 GND.n5528 163.367
R20121 GND.n6170 GND.n5529 163.367
R20122 GND.n6166 GND.n5529 163.367
R20123 GND.n6166 GND.n6165 163.367
R20124 GND.n6165 GND.n4350 163.367
R20125 GND.n4361 GND.n4350 163.367
R20126 GND.n7441 GND.n4361 163.367
R20127 GND.n7441 GND.n4362 163.367
R20128 GND.n7437 GND.n4362 163.367
R20129 GND.n7437 GND.n4365 163.367
R20130 GND.n6208 GND.n4365 163.367
R20131 GND.n6208 GND.n6204 163.367
R20132 GND.n6204 GND.n5512 163.367
R20133 GND.n6221 GND.n5512 163.367
R20134 GND.n6222 GND.n6221 163.367
R20135 GND.n6223 GND.n6222 163.367
R20136 GND.n6223 GND.n5510 163.367
R20137 GND.n6227 GND.n5510 163.367
R20138 GND.n6227 GND.n5500 163.367
R20139 GND.n6310 GND.n5500 163.367
R20140 GND.n6310 GND.n5501 163.367
R20141 GND.n6306 GND.n5501 163.367
R20142 GND.n6306 GND.n6305 163.367
R20143 GND.n6305 GND.n6304 163.367
R20144 GND.n6304 GND.n4450 163.367
R20145 GND.n7399 GND.n4450 163.367
R20146 GND.n7399 GND.n4451 163.367
R20147 GND.n7395 GND.n4451 163.367
R20148 GND.n7395 GND.n4454 163.367
R20149 GND.n6290 GND.n4454 163.367
R20150 GND.n6290 GND.n4468 163.367
R20151 GND.n7385 GND.n4468 163.367
R20152 GND.n7385 GND.n4469 163.367
R20153 GND.n7381 GND.n4469 163.367
R20154 GND.n7381 GND.n4472 163.367
R20155 GND.n6278 GND.n4472 163.367
R20156 GND.n6278 GND.n4486 163.367
R20157 GND.n7371 GND.n4486 163.367
R20158 GND.n7371 GND.n4487 163.367
R20159 GND.n7367 GND.n4487 163.367
R20160 GND.n7367 GND.n4490 163.367
R20161 GND.n6265 GND.n4490 163.367
R20162 GND.n6265 GND.n4504 163.367
R20163 GND.n7357 GND.n4504 163.367
R20164 GND.n7357 GND.n4505 163.367
R20165 GND.n7353 GND.n4505 163.367
R20166 GND.n7353 GND.n4508 163.367
R20167 GND.n6252 GND.n4508 163.367
R20168 GND.n6252 GND.n4522 163.367
R20169 GND.n7343 GND.n4522 163.367
R20170 GND.n7343 GND.n4523 163.367
R20171 GND.n7339 GND.n4523 163.367
R20172 GND.n7339 GND.n4526 163.367
R20173 GND.n4550 GND.n4526 163.367
R20174 GND.n4550 GND.n4539 163.367
R20175 GND.n4548 GND.n4539 163.367
R20176 GND.n7324 GND.n4548 163.367
R20177 GND.n7324 GND.n4549 163.367
R20178 GND.n7320 GND.n4549 163.367
R20179 GND.n7320 GND.n4555 163.367
R20180 GND.n4634 GND.n4555 163.367
R20181 GND.n4634 GND.n4572 163.367
R20182 GND.n7310 GND.n4572 163.367
R20183 GND.n7310 GND.n4573 163.367
R20184 GND.n7306 GND.n4573 163.367
R20185 GND.n7306 GND.n4576 163.367
R20186 GND.n4647 GND.n4576 163.367
R20187 GND.n4647 GND.n4590 163.367
R20188 GND.n7296 GND.n4590 163.367
R20189 GND.n7296 GND.n4591 163.367
R20190 GND.n7292 GND.n4591 163.367
R20191 GND.n7292 GND.n4594 163.367
R20192 GND.n4660 GND.n4594 163.367
R20193 GND.n4660 GND.n4608 163.367
R20194 GND.n7282 GND.n4608 163.367
R20195 GND.n7282 GND.n4609 163.367
R20196 GND.n7278 GND.n4609 163.367
R20197 GND.n7278 GND.n4612 163.367
R20198 GND.n4681 GND.n4612 163.367
R20199 GND.n4681 GND.n4622 163.367
R20200 GND.n4677 GND.n4622 163.367
R20201 GND.n7263 GND.n4677 163.367
R20202 GND.n7263 GND.n4678 163.367
R20203 GND.n7259 GND.n4678 163.367
R20204 GND.n7259 GND.n4686 163.367
R20205 GND.n4771 GND.n4686 163.367
R20206 GND.n4771 GND.n4731 163.367
R20207 GND.n2121 GND.t144 156.167
R20208 GND.n4760 GND.t27 156.167
R20209 GND.n7916 GND.t99 156.161
R20210 GND.n4758 GND.t107 156.161
R20211 GND.n9529 GND.n9528 154.062
R20212 GND.n9530 GND.n9529 154.062
R20213 GND.n9530 GND.n565 154.062
R20214 GND.n9538 GND.n565 154.062
R20215 GND.n9539 GND.n9538 154.062
R20216 GND.n9540 GND.n9539 154.062
R20217 GND.n9540 GND.n559 154.062
R20218 GND.n9548 GND.n559 154.062
R20219 GND.n9549 GND.n9548 154.062
R20220 GND.n9550 GND.n9549 154.062
R20221 GND.n9550 GND.n553 154.062
R20222 GND.n9558 GND.n553 154.062
R20223 GND.n9559 GND.n9558 154.062
R20224 GND.n9560 GND.n9559 154.062
R20225 GND.n9560 GND.n547 154.062
R20226 GND.n9568 GND.n547 154.062
R20227 GND.n9569 GND.n9568 154.062
R20228 GND.n9570 GND.n9569 154.062
R20229 GND.n9570 GND.n541 154.062
R20230 GND.n9578 GND.n541 154.062
R20231 GND.n9579 GND.n9578 154.062
R20232 GND.n9580 GND.n9579 154.062
R20233 GND.n9580 GND.n535 154.062
R20234 GND.n9588 GND.n535 154.062
R20235 GND.n9589 GND.n9588 154.062
R20236 GND.n9590 GND.n9589 154.062
R20237 GND.n9590 GND.n529 154.062
R20238 GND.n9598 GND.n529 154.062
R20239 GND.n9599 GND.n9598 154.062
R20240 GND.n9600 GND.n9599 154.062
R20241 GND.n9600 GND.n523 154.062
R20242 GND.n9608 GND.n523 154.062
R20243 GND.n9609 GND.n9608 154.062
R20244 GND.n9610 GND.n9609 154.062
R20245 GND.n9610 GND.n517 154.062
R20246 GND.n9618 GND.n517 154.062
R20247 GND.n9619 GND.n9618 154.062
R20248 GND.n9620 GND.n9619 154.062
R20249 GND.n9620 GND.n511 154.062
R20250 GND.n9628 GND.n511 154.062
R20251 GND.n9629 GND.n9628 154.062
R20252 GND.n9630 GND.n9629 154.062
R20253 GND.n9630 GND.n505 154.062
R20254 GND.n9638 GND.n505 154.062
R20255 GND.n9639 GND.n9638 154.062
R20256 GND.n9640 GND.n9639 154.062
R20257 GND.n9640 GND.n499 154.062
R20258 GND.n9648 GND.n499 154.062
R20259 GND.n9649 GND.n9648 154.062
R20260 GND.n9650 GND.n9649 154.062
R20261 GND.n9650 GND.n493 154.062
R20262 GND.n9658 GND.n493 154.062
R20263 GND.n9659 GND.n9658 154.062
R20264 GND.n9660 GND.n9659 154.062
R20265 GND.n9660 GND.n487 154.062
R20266 GND.n9668 GND.n487 154.062
R20267 GND.n9669 GND.n9668 154.062
R20268 GND.n9670 GND.n9669 154.062
R20269 GND.n9670 GND.n481 154.062
R20270 GND.n9678 GND.n481 154.062
R20271 GND.n9679 GND.n9678 154.062
R20272 GND.n9680 GND.n9679 154.062
R20273 GND.n9680 GND.n475 154.062
R20274 GND.n9692 GND.n475 154.062
R20275 GND.n9693 GND.n9692 154.062
R20276 GND.n9694 GND.n9693 154.062
R20277 GND.n4756 GND.n4755 153.553
R20278 GND.n4738 GND.t48 153.314
R20279 GND.n1923 GND.n1922 152
R20280 GND.n1924 GND.n1912 152
R20281 GND.n1926 GND.n1925 152
R20282 GND.n1927 GND.n1911 152
R20283 GND.n1929 GND.n1928 152
R20284 GND.n1931 GND.n1909 152
R20285 GND.n1933 GND.n1932 152
R20286 GND.n4754 GND.n4733 152
R20287 GND.n4745 GND.n4734 152
R20288 GND.n4744 GND.n4743 152
R20289 GND.n4742 GND.n4735 152
R20290 GND.n4741 GND.n4740 152
R20291 GND.n4739 GND.n4736 152
R20292 GND.n7188 GND.n4716 143.351
R20293 GND.n7188 GND.n4715 143.351
R20294 GND.n1889 GND.n1872 143.351
R20295 GND.n1890 GND.n1872 143.351
R20296 GND.n1919 GND.t90 135.757
R20297 GND.n48 GND.t271 131.562
R20298 GND.n50 GND.t273 130.706
R20299 GND.n49 GND.t12 130.706
R20300 GND.n48 GND.t14 130.706
R20301 GND.n1932 GND.t78 126.766
R20302 GND.n1930 GND.t127 126.766
R20303 GND.n1911 GND.t87 126.766
R20304 GND.n1924 GND.t112 126.766
R20305 GND.n1913 GND.t51 126.766
R20306 GND.n4737 GND.t148 126.766
R20307 GND.n4741 GND.t60 126.766
R20308 GND.n4743 GND.t124 126.766
R20309 GND.n4753 GND.t69 126.766
R20310 GND.n4755 GND.t103 126.766
R20311 GND.n5392 GND.n5391 110.353
R20312 GND.n5425 GND.n5424 110.353
R20313 GND.n9844 GND.n9843 110.353
R20314 GND.n10000 GND.n9999 110.353
R20315 GND.n3876 GND.t43 103.507
R20316 GND.n6342 GND.t153 103.507
R20317 GND.n7917 GND.n7916 102.207
R20318 GND.n2122 GND.n2121 102.207
R20319 GND.n4761 GND.n4760 102.207
R20320 GND.n4759 GND.n4758 102.207
R20321 GND.n9888 GND.n9812 99.6594
R20322 GND.n9892 GND.n9813 99.6594
R20323 GND.n9898 GND.n9814 99.6594
R20324 GND.n9902 GND.n9815 99.6594
R20325 GND.n9907 GND.n9816 99.6594
R20326 GND.n9911 GND.n9817 99.6594
R20327 GND.n9917 GND.n9818 99.6594
R20328 GND.n9921 GND.n9819 99.6594
R20329 GND.n9927 GND.n9820 99.6594
R20330 GND.n9931 GND.n9821 99.6594
R20331 GND.n9937 GND.n9822 99.6594
R20332 GND.n9942 GND.n9823 99.6594
R20333 GND.n9948 GND.n9824 99.6594
R20334 GND.n9952 GND.n9825 99.6594
R20335 GND.n9958 GND.n9826 99.6594
R20336 GND.n9962 GND.n9827 99.6594
R20337 GND.n9968 GND.n9828 99.6594
R20338 GND.n9862 GND.n9829 99.6594
R20339 GND.n9976 GND.n9830 99.6594
R20340 GND.n9980 GND.n9831 99.6594
R20341 GND.n9986 GND.n9832 99.6594
R20342 GND.n9990 GND.n9833 99.6594
R20343 GND.n9996 GND.n9834 99.6594
R20344 GND.n10003 GND.n9835 99.6594
R20345 GND.n10009 GND.n9836 99.6594
R20346 GND.n10013 GND.n9837 99.6594
R20347 GND.n10019 GND.n9838 99.6594
R20348 GND.n10023 GND.n9839 99.6594
R20349 GND.n10029 GND.n9840 99.6594
R20350 GND.n10032 GND.n9841 99.6594
R20351 GND.n10039 GND.n10038 99.6594
R20352 GND.n7182 GND.n7181 99.6594
R20353 GND.n7176 GND.n4840 99.6594
R20354 GND.n7173 GND.n4841 99.6594
R20355 GND.n7169 GND.n4842 99.6594
R20356 GND.n7165 GND.n4843 99.6594
R20357 GND.n7161 GND.n4844 99.6594
R20358 GND.n7158 GND.n4845 99.6594
R20359 GND.n7154 GND.n4846 99.6594
R20360 GND.n7150 GND.n4847 99.6594
R20361 GND.n7146 GND.n4848 99.6594
R20362 GND.n7142 GND.n4849 99.6594
R20363 GND.n7138 GND.n4850 99.6594
R20364 GND.n7134 GND.n4851 99.6594
R20365 GND.n7130 GND.n4852 99.6594
R20366 GND.n4853 GND.n4838 99.6594
R20367 GND.n5386 GND.n4854 99.6594
R20368 GND.n5381 GND.n4855 99.6594
R20369 GND.n5396 GND.n4856 99.6594
R20370 GND.n5402 GND.n4857 99.6594
R20371 GND.n5406 GND.n4858 99.6594
R20372 GND.n5412 GND.n4859 99.6594
R20373 GND.n5416 GND.n4860 99.6594
R20374 GND.n5422 GND.n4861 99.6594
R20375 GND.n5429 GND.n4862 99.6594
R20376 GND.n5435 GND.n4863 99.6594
R20377 GND.n5439 GND.n4864 99.6594
R20378 GND.n5445 GND.n4865 99.6594
R20379 GND.n5449 GND.n4866 99.6594
R20380 GND.n5455 GND.n4867 99.6594
R20381 GND.n1726 GND.n1721 99.6594
R20382 GND.n1728 GND.n1720 99.6594
R20383 GND.n1732 GND.n1719 99.6594
R20384 GND.n1734 GND.n1718 99.6594
R20385 GND.n1740 GND.n1717 99.6594
R20386 GND.n1742 GND.n1716 99.6594
R20387 GND.n1746 GND.n1715 99.6594
R20388 GND.n1748 GND.n1714 99.6594
R20389 GND.n1752 GND.n1713 99.6594
R20390 GND.n1754 GND.n1712 99.6594
R20391 GND.n1758 GND.n1711 99.6594
R20392 GND.n1762 GND.n1710 99.6594
R20393 GND.n1766 GND.n1709 99.6594
R20394 GND.n1870 GND.n1684 99.6594
R20395 GND.n1770 GND.n1685 99.6594
R20396 GND.n1772 GND.n1686 99.6594
R20397 GND.n1778 GND.n1687 99.6594
R20398 GND.n1780 GND.n1688 99.6594
R20399 GND.n1784 GND.n1689 99.6594
R20400 GND.n1786 GND.n1690 99.6594
R20401 GND.n1790 GND.n1691 99.6594
R20402 GND.n1792 GND.n1692 99.6594
R20403 GND.n1796 GND.n1693 99.6594
R20404 GND.n1800 GND.n1694 99.6594
R20405 GND.n1804 GND.n1695 99.6594
R20406 GND.n1806 GND.n1696 99.6594
R20407 GND.n1810 GND.n1697 99.6594
R20408 GND.n1812 GND.n1698 99.6594
R20409 GND.n1816 GND.n1699 99.6594
R20410 GND.n1700 GND.n1675 99.6594
R20411 GND.n8361 GND.n8360 99.6594
R20412 GND.n8355 GND.n1322 99.6594
R20413 GND.n8352 GND.n1323 99.6594
R20414 GND.n8348 GND.n1324 99.6594
R20415 GND.n8344 GND.n1325 99.6594
R20416 GND.n8340 GND.n1326 99.6594
R20417 GND.n8337 GND.n1327 99.6594
R20418 GND.n8333 GND.n1328 99.6594
R20419 GND.n8329 GND.n1329 99.6594
R20420 GND.n8325 GND.n1330 99.6594
R20421 GND.n8321 GND.n1331 99.6594
R20422 GND.n8317 GND.n1332 99.6594
R20423 GND.n8313 GND.n1333 99.6594
R20424 GND.n8309 GND.n1334 99.6594
R20425 GND.n8305 GND.n1335 99.6594
R20426 GND.n8301 GND.n1336 99.6594
R20427 GND.n8297 GND.n1337 99.6594
R20428 GND.n8293 GND.n1338 99.6594
R20429 GND.n8289 GND.n1339 99.6594
R20430 GND.n8285 GND.n1340 99.6594
R20431 GND.n8281 GND.n1341 99.6594
R20432 GND.n8277 GND.n1342 99.6594
R20433 GND.n8273 GND.n1343 99.6594
R20434 GND.n8269 GND.n1344 99.6594
R20435 GND.n8264 GND.n1345 99.6594
R20436 GND.n8260 GND.n1346 99.6594
R20437 GND.n8256 GND.n1347 99.6594
R20438 GND.n8252 GND.n1348 99.6594
R20439 GND.n8248 GND.n1349 99.6594
R20440 GND.n8244 GND.n1350 99.6594
R20441 GND.n6317 GND.n4423 99.6594
R20442 GND.n6323 GND.n4424 99.6594
R20443 GND.n6327 GND.n4425 99.6594
R20444 GND.n6333 GND.n4426 99.6594
R20445 GND.n6337 GND.n4427 99.6594
R20446 GND.n5489 GND.n4428 99.6594
R20447 GND.n5484 GND.n4429 99.6594
R20448 GND.n5479 GND.n4430 99.6594
R20449 GND.n5474 GND.n4431 99.6594
R20450 GND.n5469 GND.n4432 99.6594
R20451 GND.n6353 GND.n4433 99.6594
R20452 GND.n6351 GND.n4434 99.6594
R20453 GND.n6347 GND.n4435 99.6594
R20454 GND.n7410 GND.n7409 99.6594
R20455 GND.n7758 GND.n7757 99.6594
R20456 GND.n7752 GND.n2328 99.6594
R20457 GND.n7749 GND.n2329 99.6594
R20458 GND.n7745 GND.n2330 99.6594
R20459 GND.n7741 GND.n2331 99.6594
R20460 GND.n2356 GND.n2332 99.6594
R20461 GND.n7734 GND.n2333 99.6594
R20462 GND.n7729 GND.n2334 99.6594
R20463 GND.n7724 GND.n2335 99.6594
R20464 GND.n7719 GND.n2336 99.6594
R20465 GND.n7714 GND.n2337 99.6594
R20466 GND.n7709 GND.n2338 99.6594
R20467 GND.n7705 GND.n2339 99.6594
R20468 GND.n10053 GND.n10040 99.6594
R20469 GND.n10057 GND.n10041 99.6594
R20470 GND.n10063 GND.n10042 99.6594
R20471 GND.n10066 GND.n10043 99.6594
R20472 GND.n10073 GND.n10072 99.6594
R20473 GND.n10076 GND.n10075 99.6594
R20474 GND.n6361 GND.n4875 99.6594
R20475 GND.n6365 GND.n4874 99.6594
R20476 GND.n6370 GND.n4873 99.6594
R20477 GND.n6375 GND.n4872 99.6594
R20478 GND.n6380 GND.n4871 99.6594
R20479 GND.n6358 GND.n4870 99.6594
R20480 GND.n6364 GND.n4875 99.6594
R20481 GND.n6369 GND.n4874 99.6594
R20482 GND.n6374 GND.n4873 99.6594
R20483 GND.n6379 GND.n4872 99.6594
R20484 GND.n6383 GND.n4871 99.6594
R20485 GND.n6387 GND.n4870 99.6594
R20486 GND.n10075 GND.n9811 99.6594
R20487 GND.n10073 GND.n10044 99.6594
R20488 GND.n10064 GND.n10043 99.6594
R20489 GND.n10056 GND.n10042 99.6594
R20490 GND.n10054 GND.n10041 99.6594
R20491 GND.n10040 GND.n418 99.6594
R20492 GND.n7758 GND.n2343 99.6594
R20493 GND.n7750 GND.n2328 99.6594
R20494 GND.n7746 GND.n2329 99.6594
R20495 GND.n7742 GND.n2330 99.6594
R20496 GND.n2355 GND.n2331 99.6594
R20497 GND.n7733 GND.n2332 99.6594
R20498 GND.n7728 GND.n2333 99.6594
R20499 GND.n7723 GND.n2334 99.6594
R20500 GND.n7718 GND.n2335 99.6594
R20501 GND.n7713 GND.n2336 99.6594
R20502 GND.n3875 GND.n2337 99.6594
R20503 GND.n7706 GND.n2338 99.6594
R20504 GND.n3880 GND.n2339 99.6594
R20505 GND.n7409 GND.n4421 99.6594
R20506 GND.n6350 GND.n4435 99.6594
R20507 GND.n6354 GND.n4434 99.6594
R20508 GND.n5468 GND.n4433 99.6594
R20509 GND.n5473 GND.n4432 99.6594
R20510 GND.n5478 GND.n4431 99.6594
R20511 GND.n5483 GND.n4430 99.6594
R20512 GND.n5488 GND.n4429 99.6594
R20513 GND.n6338 GND.n4428 99.6594
R20514 GND.n6334 GND.n4427 99.6594
R20515 GND.n6328 GND.n4426 99.6594
R20516 GND.n6324 GND.n4425 99.6594
R20517 GND.n6318 GND.n4424 99.6594
R20518 GND.n6314 GND.n4423 99.6594
R20519 GND.n8361 GND.n1361 99.6594
R20520 GND.n8353 GND.n1322 99.6594
R20521 GND.n8349 GND.n1323 99.6594
R20522 GND.n8345 GND.n1324 99.6594
R20523 GND.n1373 GND.n1325 99.6594
R20524 GND.n8338 GND.n1326 99.6594
R20525 GND.n8334 GND.n1327 99.6594
R20526 GND.n8330 GND.n1328 99.6594
R20527 GND.n8326 GND.n1329 99.6594
R20528 GND.n8322 GND.n1330 99.6594
R20529 GND.n8318 GND.n1331 99.6594
R20530 GND.n8314 GND.n1332 99.6594
R20531 GND.n8310 GND.n1333 99.6594
R20532 GND.n8306 GND.n1334 99.6594
R20533 GND.n8302 GND.n1335 99.6594
R20534 GND.n8298 GND.n1336 99.6594
R20535 GND.n8294 GND.n1337 99.6594
R20536 GND.n8290 GND.n1338 99.6594
R20537 GND.n8286 GND.n1339 99.6594
R20538 GND.n8282 GND.n1340 99.6594
R20539 GND.n8278 GND.n1341 99.6594
R20540 GND.n8274 GND.n1342 99.6594
R20541 GND.n8270 GND.n1343 99.6594
R20542 GND.n8265 GND.n1344 99.6594
R20543 GND.n8261 GND.n1345 99.6594
R20544 GND.n8257 GND.n1346 99.6594
R20545 GND.n8253 GND.n1347 99.6594
R20546 GND.n8249 GND.n1348 99.6594
R20547 GND.n8245 GND.n1349 99.6594
R20548 GND.n1434 GND.n1350 99.6594
R20549 GND.n1819 GND.n1700 99.6594
R20550 GND.n1813 GND.n1699 99.6594
R20551 GND.n1811 GND.n1698 99.6594
R20552 GND.n1807 GND.n1697 99.6594
R20553 GND.n1805 GND.n1696 99.6594
R20554 GND.n1801 GND.n1695 99.6594
R20555 GND.n1799 GND.n1694 99.6594
R20556 GND.n1793 GND.n1693 99.6594
R20557 GND.n1791 GND.n1692 99.6594
R20558 GND.n1787 GND.n1691 99.6594
R20559 GND.n1785 GND.n1690 99.6594
R20560 GND.n1781 GND.n1689 99.6594
R20561 GND.n1779 GND.n1688 99.6594
R20562 GND.n1773 GND.n1687 99.6594
R20563 GND.n1771 GND.n1686 99.6594
R20564 GND.n1767 GND.n1685 99.6594
R20565 GND.n7978 GND.n1708 99.6594
R20566 GND.n1763 GND.n1709 99.6594
R20567 GND.n1761 GND.n1710 99.6594
R20568 GND.n1755 GND.n1711 99.6594
R20569 GND.n1753 GND.n1712 99.6594
R20570 GND.n1749 GND.n1713 99.6594
R20571 GND.n1747 GND.n1714 99.6594
R20572 GND.n1743 GND.n1715 99.6594
R20573 GND.n1741 GND.n1716 99.6594
R20574 GND.n1735 GND.n1717 99.6594
R20575 GND.n1733 GND.n1718 99.6594
R20576 GND.n1729 GND.n1719 99.6594
R20577 GND.n1727 GND.n1720 99.6594
R20578 GND.n1722 GND.n1721 99.6594
R20579 GND.n7182 GND.n4877 99.6594
R20580 GND.n7174 GND.n4840 99.6594
R20581 GND.n7170 GND.n4841 99.6594
R20582 GND.n7166 GND.n4842 99.6594
R20583 GND.n7106 GND.n4843 99.6594
R20584 GND.n7159 GND.n4844 99.6594
R20585 GND.n7155 GND.n4845 99.6594
R20586 GND.n7151 GND.n4846 99.6594
R20587 GND.n7147 GND.n4847 99.6594
R20588 GND.n7143 GND.n4848 99.6594
R20589 GND.n7139 GND.n4849 99.6594
R20590 GND.n7135 GND.n4850 99.6594
R20591 GND.n7131 GND.n4851 99.6594
R20592 GND.n7185 GND.n7184 99.6594
R20593 GND.n5385 GND.n4853 99.6594
R20594 GND.n5380 GND.n4854 99.6594
R20595 GND.n5395 GND.n4855 99.6594
R20596 GND.n5401 GND.n4856 99.6594
R20597 GND.n5405 GND.n4857 99.6594
R20598 GND.n5411 GND.n4858 99.6594
R20599 GND.n5415 GND.n4859 99.6594
R20600 GND.n5421 GND.n4860 99.6594
R20601 GND.n5428 GND.n4861 99.6594
R20602 GND.n5434 GND.n4862 99.6594
R20603 GND.n5438 GND.n4863 99.6594
R20604 GND.n5444 GND.n4864 99.6594
R20605 GND.n5448 GND.n4865 99.6594
R20606 GND.n5454 GND.n4866 99.6594
R20607 GND.n5457 GND.n4867 99.6594
R20608 GND.n10039 GND.n9842 99.6594
R20609 GND.n10030 GND.n9841 99.6594
R20610 GND.n10022 GND.n9840 99.6594
R20611 GND.n10020 GND.n9839 99.6594
R20612 GND.n10012 GND.n9838 99.6594
R20613 GND.n10010 GND.n9837 99.6594
R20614 GND.n10002 GND.n9836 99.6594
R20615 GND.n9997 GND.n9835 99.6594
R20616 GND.n9989 GND.n9834 99.6594
R20617 GND.n9987 GND.n9833 99.6594
R20618 GND.n9979 GND.n9832 99.6594
R20619 GND.n9977 GND.n9831 99.6594
R20620 GND.n9861 GND.n9830 99.6594
R20621 GND.n9969 GND.n9829 99.6594
R20622 GND.n9961 GND.n9828 99.6594
R20623 GND.n9959 GND.n9827 99.6594
R20624 GND.n9951 GND.n9826 99.6594
R20625 GND.n9949 GND.n9825 99.6594
R20626 GND.n9941 GND.n9824 99.6594
R20627 GND.n9938 GND.n9823 99.6594
R20628 GND.n9930 GND.n9822 99.6594
R20629 GND.n9928 GND.n9821 99.6594
R20630 GND.n9920 GND.n9820 99.6594
R20631 GND.n9918 GND.n9819 99.6594
R20632 GND.n9910 GND.n9818 99.6594
R20633 GND.n9879 GND.n9817 99.6594
R20634 GND.n9901 GND.n9816 99.6594
R20635 GND.n9899 GND.n9815 99.6594
R20636 GND.n9891 GND.n9814 99.6594
R20637 GND.n9889 GND.n9813 99.6594
R20638 GND.n9812 GND.n414 99.6594
R20639 GND.n1439 GND.n1352 99.6594
R20640 GND.n1441 GND.n1353 99.6594
R20641 GND.n1445 GND.n1354 99.6594
R20642 GND.n1447 GND.n1355 99.6594
R20643 GND.n1451 GND.n1356 99.6594
R20644 GND.n1440 GND.n1352 99.6594
R20645 GND.n1444 GND.n1353 99.6594
R20646 GND.n1446 GND.n1354 99.6594
R20647 GND.n1450 GND.n1355 99.6594
R20648 GND.n8220 GND.n1356 99.6594
R20649 GND.n1701 GND.n1681 99.6594
R20650 GND.n3858 GND.n1702 99.6594
R20651 GND.n3862 GND.n1703 99.6594
R20652 GND.n3866 GND.n1704 99.6594
R20653 GND.n3870 GND.n1705 99.6594
R20654 GND.n3854 GND.n1705 99.6594
R20655 GND.n3869 GND.n1704 99.6594
R20656 GND.n3865 GND.n1703 99.6594
R20657 GND.n3861 GND.n1702 99.6594
R20658 GND.n3857 GND.n1701 99.6594
R20659 GND.n8222 GND.n8221 97.552
R20660 GND.n1739 GND.n1738 97.552
R20661 GND.n1760 GND.n1759 97.552
R20662 GND.n1777 GND.n1776 97.552
R20663 GND.n1798 GND.n1797 97.552
R20664 GND.n1818 GND.n1817 97.552
R20665 GND.n7109 GND.n7108 97.552
R20666 GND.n7123 GND.n7122 97.552
R20667 GND.n5459 GND.n5458 97.552
R20668 GND.n9860 GND.n9859 97.552
R20669 GND.n9870 GND.n9869 97.552
R20670 GND.n9878 GND.n9877 97.552
R20671 GND.n9809 GND.n9808 97.552
R20672 GND.n6360 GND.n6359 97.552
R20673 GND.n1376 GND.n1375 97.552
R20674 GND.n1390 GND.n1389 97.552
R20675 GND.n1406 GND.n1405 97.552
R20676 GND.n1420 GND.n1419 97.552
R20677 GND.n1436 GND.n1435 97.552
R20678 GND.n3853 GND.n3852 97.552
R20679 GND.n1920 GND.n1919 76.4039
R20680 GND.n8 GND.t192 73.1986
R20681 GND.n15 GND.t241 73.1986
R20682 GND.n23 GND.t209 73.1986
R20683 GND.n31 GND.t158 73.1986
R20684 GND.n39 GND.t205 73.1986
R20685 GND.n1 GND.t233 73.1986
R20686 GND.n56 GND.t184 73.1986
R20687 GND.n63 GND.t238 73.1986
R20688 GND.n71 GND.t235 73.1986
R20689 GND.n79 GND.t266 73.1986
R20690 GND.n87 GND.t239 73.1986
R20691 GND.n95 GND.t172 73.1986
R20692 GND.n1921 GND.n1913 72.8411
R20693 GND.n1930 GND.n1910 72.8411
R20694 GND.n4753 GND.n4752 72.8411
R20695 GND.n7244 GND.n4730 71.676
R20696 GND.n7240 GND.n4729 71.676
R20697 GND.n7236 GND.n4728 71.676
R20698 GND.n7232 GND.n4727 71.676
R20699 GND.n7228 GND.n4726 71.676
R20700 GND.n7224 GND.n4725 71.676
R20701 GND.n7220 GND.n4724 71.676
R20702 GND.n7216 GND.n4723 71.676
R20703 GND.n7212 GND.n4722 71.676
R20704 GND.n7208 GND.n4721 71.676
R20705 GND.n7204 GND.n4720 71.676
R20706 GND.n7200 GND.n4719 71.676
R20707 GND.n7195 GND.n4718 71.676
R20708 GND.n7191 GND.n4717 71.676
R20709 GND.n4831 GND.n4715 71.676
R20710 GND.n4827 GND.n4714 71.676
R20711 GND.n4823 GND.n4713 71.676
R20712 GND.n4819 GND.n4712 71.676
R20713 GND.n4815 GND.n4711 71.676
R20714 GND.n4811 GND.n4710 71.676
R20715 GND.n4807 GND.n4709 71.676
R20716 GND.n4803 GND.n4708 71.676
R20717 GND.n4799 GND.n4707 71.676
R20718 GND.n4795 GND.n4706 71.676
R20719 GND.n4791 GND.n4705 71.676
R20720 GND.n4787 GND.n4704 71.676
R20721 GND.n4783 GND.n4703 71.676
R20722 GND.n4779 GND.n4702 71.676
R20723 GND.n4775 GND.n4701 71.676
R20724 GND.n7971 GND.n7970 71.676
R20725 GND.n7965 GND.n1877 71.676
R20726 GND.n7962 GND.n1878 71.676
R20727 GND.n7958 GND.n1879 71.676
R20728 GND.n7954 GND.n1880 71.676
R20729 GND.n7950 GND.n1881 71.676
R20730 GND.n7946 GND.n1882 71.676
R20731 GND.n7942 GND.n1883 71.676
R20732 GND.n7938 GND.n1884 71.676
R20733 GND.n7934 GND.n1885 71.676
R20734 GND.n7930 GND.n1886 71.676
R20735 GND.n7926 GND.n1887 71.676
R20736 GND.n7922 GND.n1888 71.676
R20737 GND.n7973 GND.n1875 71.676
R20738 GND.n1889 GND.n1873 71.676
R20739 GND.n2125 GND.n1891 71.676
R20740 GND.n2129 GND.n1892 71.676
R20741 GND.n2133 GND.n1893 71.676
R20742 GND.n2137 GND.n1894 71.676
R20743 GND.n2141 GND.n1895 71.676
R20744 GND.n2145 GND.n1896 71.676
R20745 GND.n2149 GND.n1897 71.676
R20746 GND.n2153 GND.n1898 71.676
R20747 GND.n2157 GND.n1899 71.676
R20748 GND.n2161 GND.n1900 71.676
R20749 GND.n2165 GND.n1901 71.676
R20750 GND.n2169 GND.n1902 71.676
R20751 GND.n2173 GND.n1903 71.676
R20752 GND.n2177 GND.n1904 71.676
R20753 GND.n7971 GND.n1907 71.676
R20754 GND.n7963 GND.n1877 71.676
R20755 GND.n7959 GND.n1878 71.676
R20756 GND.n7955 GND.n1879 71.676
R20757 GND.n7951 GND.n1880 71.676
R20758 GND.n7947 GND.n1881 71.676
R20759 GND.n7943 GND.n1882 71.676
R20760 GND.n7939 GND.n1883 71.676
R20761 GND.n7935 GND.n1884 71.676
R20762 GND.n7931 GND.n1885 71.676
R20763 GND.n7927 GND.n1886 71.676
R20764 GND.n7923 GND.n1887 71.676
R20765 GND.n7918 GND.n1888 71.676
R20766 GND.n7974 GND.n7973 71.676
R20767 GND.n2124 GND.n1890 71.676
R20768 GND.n2128 GND.n1891 71.676
R20769 GND.n2132 GND.n1892 71.676
R20770 GND.n2136 GND.n1893 71.676
R20771 GND.n2140 GND.n1894 71.676
R20772 GND.n2144 GND.n1895 71.676
R20773 GND.n2148 GND.n1896 71.676
R20774 GND.n2152 GND.n1897 71.676
R20775 GND.n2156 GND.n1898 71.676
R20776 GND.n2160 GND.n1899 71.676
R20777 GND.n2164 GND.n1900 71.676
R20778 GND.n2168 GND.n1901 71.676
R20779 GND.n2172 GND.n1902 71.676
R20780 GND.n2176 GND.n1903 71.676
R20781 GND.n2180 GND.n1904 71.676
R20782 GND.n4778 GND.n4701 71.676
R20783 GND.n4782 GND.n4702 71.676
R20784 GND.n4786 GND.n4703 71.676
R20785 GND.n4790 GND.n4704 71.676
R20786 GND.n4794 GND.n4705 71.676
R20787 GND.n4798 GND.n4706 71.676
R20788 GND.n4802 GND.n4707 71.676
R20789 GND.n4806 GND.n4708 71.676
R20790 GND.n4810 GND.n4709 71.676
R20791 GND.n4814 GND.n4710 71.676
R20792 GND.n4818 GND.n4711 71.676
R20793 GND.n4822 GND.n4712 71.676
R20794 GND.n4826 GND.n4713 71.676
R20795 GND.n4830 GND.n4714 71.676
R20796 GND.n7190 GND.n4716 71.676
R20797 GND.n7194 GND.n4717 71.676
R20798 GND.n7199 GND.n4718 71.676
R20799 GND.n7203 GND.n4719 71.676
R20800 GND.n7207 GND.n4720 71.676
R20801 GND.n7211 GND.n4721 71.676
R20802 GND.n7215 GND.n4722 71.676
R20803 GND.n7219 GND.n4723 71.676
R20804 GND.n7223 GND.n4724 71.676
R20805 GND.n7227 GND.n4725 71.676
R20806 GND.n7231 GND.n4726 71.676
R20807 GND.n7235 GND.n4727 71.676
R20808 GND.n7239 GND.n4728 71.676
R20809 GND.n7243 GND.n4729 71.676
R20810 GND.n4732 GND.n4730 71.676
R20811 GND.n13 GND.t253 71.5636
R20812 GND.n20 GND.t203 71.5636
R20813 GND.n28 GND.t217 71.5636
R20814 GND.n36 GND.t225 71.5636
R20815 GND.n44 GND.t257 71.5636
R20816 GND.n6 GND.t188 71.5636
R20817 GND.n61 GND.t182 71.5636
R20818 GND.n68 GND.t231 71.5636
R20819 GND.n76 GND.t220 71.5636
R20820 GND.n84 GND.t256 71.5636
R20821 GND.n92 GND.t230 71.5636
R20822 GND.n100 GND.t265 71.5636
R20823 GND.n8499 GND.n8498 70.6492
R20824 GND.n8499 GND.n1182 70.6492
R20825 GND.n8507 GND.n1182 70.6492
R20826 GND.n8508 GND.n8507 70.6492
R20827 GND.n8509 GND.n8508 70.6492
R20828 GND.n8509 GND.n1176 70.6492
R20829 GND.n8517 GND.n1176 70.6492
R20830 GND.n8518 GND.n8517 70.6492
R20831 GND.n8519 GND.n8518 70.6492
R20832 GND.n8519 GND.n1170 70.6492
R20833 GND.n8527 GND.n1170 70.6492
R20834 GND.n8528 GND.n8527 70.6492
R20835 GND.n8529 GND.n8528 70.6492
R20836 GND.n8529 GND.n1164 70.6492
R20837 GND.n8537 GND.n1164 70.6492
R20838 GND.n8538 GND.n8537 70.6492
R20839 GND.n8539 GND.n8538 70.6492
R20840 GND.n8539 GND.n1158 70.6492
R20841 GND.n8547 GND.n1158 70.6492
R20842 GND.n8548 GND.n8547 70.6492
R20843 GND.n8549 GND.n8548 70.6492
R20844 GND.n8549 GND.n1152 70.6492
R20845 GND.n8557 GND.n1152 70.6492
R20846 GND.n8558 GND.n8557 70.6492
R20847 GND.n8559 GND.n8558 70.6492
R20848 GND.n8559 GND.n1146 70.6492
R20849 GND.n8567 GND.n1146 70.6492
R20850 GND.n8568 GND.n8567 70.6492
R20851 GND.n8569 GND.n8568 70.6492
R20852 GND.n8569 GND.n1140 70.6492
R20853 GND.n8577 GND.n1140 70.6492
R20854 GND.n8578 GND.n8577 70.6492
R20855 GND.n8579 GND.n8578 70.6492
R20856 GND.n8579 GND.n1134 70.6492
R20857 GND.n8587 GND.n1134 70.6492
R20858 GND.n8588 GND.n8587 70.6492
R20859 GND.n8589 GND.n8588 70.6492
R20860 GND.n8589 GND.n1128 70.6492
R20861 GND.n8597 GND.n1128 70.6492
R20862 GND.n8598 GND.n8597 70.6492
R20863 GND.n8599 GND.n8598 70.6492
R20864 GND.n8599 GND.n1122 70.6492
R20865 GND.n8607 GND.n1122 70.6492
R20866 GND.n8608 GND.n8607 70.6492
R20867 GND.n8609 GND.n8608 70.6492
R20868 GND.n8609 GND.n1116 70.6492
R20869 GND.n8617 GND.n1116 70.6492
R20870 GND.n8618 GND.n8617 70.6492
R20871 GND.n8619 GND.n8618 70.6492
R20872 GND.n8619 GND.n1110 70.6492
R20873 GND.n8627 GND.n1110 70.6492
R20874 GND.n8628 GND.n8627 70.6492
R20875 GND.n8629 GND.n8628 70.6492
R20876 GND.n8629 GND.n1104 70.6492
R20877 GND.n8637 GND.n1104 70.6492
R20878 GND.n8638 GND.n8637 70.6492
R20879 GND.n8639 GND.n8638 70.6492
R20880 GND.n8639 GND.n1098 70.6492
R20881 GND.n8647 GND.n1098 70.6492
R20882 GND.n8648 GND.n8647 70.6492
R20883 GND.n8649 GND.n8648 70.6492
R20884 GND.n8649 GND.n1092 70.6492
R20885 GND.n8657 GND.n1092 70.6492
R20886 GND.n8658 GND.n8657 70.6492
R20887 GND.n8659 GND.n8658 70.6492
R20888 GND.n8659 GND.n1086 70.6492
R20889 GND.n8667 GND.n1086 70.6492
R20890 GND.n8668 GND.n8667 70.6492
R20891 GND.n8669 GND.n8668 70.6492
R20892 GND.n8669 GND.n1080 70.6492
R20893 GND.n8677 GND.n1080 70.6492
R20894 GND.n8678 GND.n8677 70.6492
R20895 GND.n8679 GND.n8678 70.6492
R20896 GND.n8679 GND.n1074 70.6492
R20897 GND.n8687 GND.n1074 70.6492
R20898 GND.n8688 GND.n8687 70.6492
R20899 GND.n8689 GND.n8688 70.6492
R20900 GND.n8689 GND.n1068 70.6492
R20901 GND.n8697 GND.n1068 70.6492
R20902 GND.n8698 GND.n8697 70.6492
R20903 GND.n8699 GND.n8698 70.6492
R20904 GND.n8699 GND.n1062 70.6492
R20905 GND.n8707 GND.n1062 70.6492
R20906 GND.n8708 GND.n8707 70.6492
R20907 GND.n8709 GND.n8708 70.6492
R20908 GND.n8709 GND.n1056 70.6492
R20909 GND.n8717 GND.n1056 70.6492
R20910 GND.n8718 GND.n8717 70.6492
R20911 GND.n8719 GND.n8718 70.6492
R20912 GND.n8719 GND.n1050 70.6492
R20913 GND.n8727 GND.n1050 70.6492
R20914 GND.n8728 GND.n8727 70.6492
R20915 GND.n8729 GND.n8728 70.6492
R20916 GND.n8729 GND.n1044 70.6492
R20917 GND.n8737 GND.n1044 70.6492
R20918 GND.n8738 GND.n8737 70.6492
R20919 GND.n8739 GND.n8738 70.6492
R20920 GND.n8739 GND.n1038 70.6492
R20921 GND.n8747 GND.n1038 70.6492
R20922 GND.n8748 GND.n8747 70.6492
R20923 GND.n8749 GND.n8748 70.6492
R20924 GND.n8749 GND.n1032 70.6492
R20925 GND.n8757 GND.n1032 70.6492
R20926 GND.n8758 GND.n8757 70.6492
R20927 GND.n8759 GND.n8758 70.6492
R20928 GND.n8759 GND.n1026 70.6492
R20929 GND.n8767 GND.n1026 70.6492
R20930 GND.n8768 GND.n8767 70.6492
R20931 GND.n8769 GND.n8768 70.6492
R20932 GND.n8769 GND.n1020 70.6492
R20933 GND.n8777 GND.n1020 70.6492
R20934 GND.n8778 GND.n8777 70.6492
R20935 GND.n8779 GND.n8778 70.6492
R20936 GND.n8779 GND.n1014 70.6492
R20937 GND.n8787 GND.n1014 70.6492
R20938 GND.n8788 GND.n8787 70.6492
R20939 GND.n8789 GND.n8788 70.6492
R20940 GND.n8789 GND.n1008 70.6492
R20941 GND.n8797 GND.n1008 70.6492
R20942 GND.n8798 GND.n8797 70.6492
R20943 GND.n8799 GND.n8798 70.6492
R20944 GND.n8799 GND.n1002 70.6492
R20945 GND.n8807 GND.n1002 70.6492
R20946 GND.n8808 GND.n8807 70.6492
R20947 GND.n8809 GND.n8808 70.6492
R20948 GND.n8809 GND.n996 70.6492
R20949 GND.n8817 GND.n996 70.6492
R20950 GND.n8818 GND.n8817 70.6492
R20951 GND.n8819 GND.n8818 70.6492
R20952 GND.n8819 GND.n990 70.6492
R20953 GND.n8827 GND.n990 70.6492
R20954 GND.n8828 GND.n8827 70.6492
R20955 GND.n8829 GND.n8828 70.6492
R20956 GND.n8829 GND.n984 70.6492
R20957 GND.n8837 GND.n984 70.6492
R20958 GND.n8838 GND.n8837 70.6492
R20959 GND.n8839 GND.n8838 70.6492
R20960 GND.n8839 GND.n978 70.6492
R20961 GND.n8847 GND.n978 70.6492
R20962 GND.n8848 GND.n8847 70.6492
R20963 GND.n8849 GND.n8848 70.6492
R20964 GND.n8849 GND.n972 70.6492
R20965 GND.n8857 GND.n972 70.6492
R20966 GND.n8858 GND.n8857 70.6492
R20967 GND.n8859 GND.n8858 70.6492
R20968 GND.n8859 GND.n966 70.6492
R20969 GND.n8867 GND.n966 70.6492
R20970 GND.n8868 GND.n8867 70.6492
R20971 GND.n8869 GND.n8868 70.6492
R20972 GND.n8869 GND.n960 70.6492
R20973 GND.n8877 GND.n960 70.6492
R20974 GND.n8878 GND.n8877 70.6492
R20975 GND.n8879 GND.n8878 70.6492
R20976 GND.n8879 GND.n954 70.6492
R20977 GND.n8887 GND.n954 70.6492
R20978 GND.n8888 GND.n8887 70.6492
R20979 GND.n8889 GND.n8888 70.6492
R20980 GND.n8889 GND.n948 70.6492
R20981 GND.n8897 GND.n948 70.6492
R20982 GND.n8898 GND.n8897 70.6492
R20983 GND.n8899 GND.n8898 70.6492
R20984 GND.n8899 GND.n942 70.6492
R20985 GND.n8907 GND.n942 70.6492
R20986 GND.n8908 GND.n8907 70.6492
R20987 GND.n8909 GND.n8908 70.6492
R20988 GND.n8909 GND.n936 70.6492
R20989 GND.n8917 GND.n936 70.6492
R20990 GND.n8918 GND.n8917 70.6492
R20991 GND.n8919 GND.n8918 70.6492
R20992 GND.n8919 GND.n930 70.6492
R20993 GND.n8927 GND.n930 70.6492
R20994 GND.n8928 GND.n8927 70.6492
R20995 GND.n8929 GND.n8928 70.6492
R20996 GND.n8929 GND.n924 70.6492
R20997 GND.n8937 GND.n924 70.6492
R20998 GND.n8938 GND.n8937 70.6492
R20999 GND.n8939 GND.n8938 70.6492
R21000 GND.n8939 GND.n918 70.6492
R21001 GND.n8947 GND.n918 70.6492
R21002 GND.n8948 GND.n8947 70.6492
R21003 GND.n8949 GND.n8948 70.6492
R21004 GND.n8949 GND.n912 70.6492
R21005 GND.n8957 GND.n912 70.6492
R21006 GND.n8958 GND.n8957 70.6492
R21007 GND.n8959 GND.n8958 70.6492
R21008 GND.n8959 GND.n906 70.6492
R21009 GND.n8967 GND.n906 70.6492
R21010 GND.n8968 GND.n8967 70.6492
R21011 GND.n8969 GND.n8968 70.6492
R21012 GND.n8969 GND.n900 70.6492
R21013 GND.n8977 GND.n900 70.6492
R21014 GND.n8978 GND.n8977 70.6492
R21015 GND.n8979 GND.n8978 70.6492
R21016 GND.n8979 GND.n894 70.6492
R21017 GND.n8987 GND.n894 70.6492
R21018 GND.n8988 GND.n8987 70.6492
R21019 GND.n8989 GND.n8988 70.6492
R21020 GND.n8989 GND.n888 70.6492
R21021 GND.n8997 GND.n888 70.6492
R21022 GND.n8998 GND.n8997 70.6492
R21023 GND.n8999 GND.n8998 70.6492
R21024 GND.n8999 GND.n882 70.6492
R21025 GND.n9007 GND.n882 70.6492
R21026 GND.n9008 GND.n9007 70.6492
R21027 GND.n9009 GND.n9008 70.6492
R21028 GND.n9009 GND.n876 70.6492
R21029 GND.n9017 GND.n876 70.6492
R21030 GND.n9018 GND.n9017 70.6492
R21031 GND.n9019 GND.n9018 70.6492
R21032 GND.n9019 GND.n870 70.6492
R21033 GND.n9027 GND.n870 70.6492
R21034 GND.n9028 GND.n9027 70.6492
R21035 GND.n9029 GND.n9028 70.6492
R21036 GND.n9029 GND.n864 70.6492
R21037 GND.n9037 GND.n864 70.6492
R21038 GND.n9038 GND.n9037 70.6492
R21039 GND.n9039 GND.n9038 70.6492
R21040 GND.n9039 GND.n858 70.6492
R21041 GND.n9047 GND.n858 70.6492
R21042 GND.n9048 GND.n9047 70.6492
R21043 GND.n9049 GND.n9048 70.6492
R21044 GND.n9049 GND.n852 70.6492
R21045 GND.n9057 GND.n852 70.6492
R21046 GND.n9058 GND.n9057 70.6492
R21047 GND.n9059 GND.n9058 70.6492
R21048 GND.n9059 GND.n846 70.6492
R21049 GND.n9067 GND.n846 70.6492
R21050 GND.n9068 GND.n9067 70.6492
R21051 GND.n9069 GND.n9068 70.6492
R21052 GND.n9069 GND.n840 70.6492
R21053 GND.n9077 GND.n840 70.6492
R21054 GND.n9078 GND.n9077 70.6492
R21055 GND.n9079 GND.n9078 70.6492
R21056 GND.n9079 GND.n834 70.6492
R21057 GND.n9087 GND.n834 70.6492
R21058 GND.n9088 GND.n9087 70.6492
R21059 GND.n9089 GND.n9088 70.6492
R21060 GND.n9089 GND.n828 70.6492
R21061 GND.n9097 GND.n828 70.6492
R21062 GND.n9098 GND.n9097 70.6492
R21063 GND.n9099 GND.n9098 70.6492
R21064 GND.n9099 GND.n822 70.6492
R21065 GND.n9107 GND.n822 70.6492
R21066 GND.n9108 GND.n9107 70.6492
R21067 GND.n9109 GND.n9108 70.6492
R21068 GND.n9109 GND.n816 70.6492
R21069 GND.n9117 GND.n816 70.6492
R21070 GND.n9118 GND.n9117 70.6492
R21071 GND.n9119 GND.n9118 70.6492
R21072 GND.n9119 GND.n810 70.6492
R21073 GND.n9127 GND.n810 70.6492
R21074 GND.n9128 GND.n9127 70.6492
R21075 GND.n9129 GND.n9128 70.6492
R21076 GND.n9129 GND.n804 70.6492
R21077 GND.n9137 GND.n804 70.6492
R21078 GND.n9138 GND.n9137 70.6492
R21079 GND.n9139 GND.n9138 70.6492
R21080 GND.n9139 GND.n798 70.6492
R21081 GND.n9147 GND.n798 70.6492
R21082 GND.n9148 GND.n9147 70.6492
R21083 GND.n9149 GND.n9148 70.6492
R21084 GND.n9149 GND.n792 70.6492
R21085 GND.n9157 GND.n792 70.6492
R21086 GND.n9158 GND.n9157 70.6492
R21087 GND.n9159 GND.n9158 70.6492
R21088 GND.n9159 GND.n786 70.6492
R21089 GND.n9167 GND.n786 70.6492
R21090 GND.n9168 GND.n9167 70.6492
R21091 GND.n9169 GND.n9168 70.6492
R21092 GND.n9169 GND.n780 70.6492
R21093 GND.n9177 GND.n780 70.6492
R21094 GND.n9178 GND.n9177 70.6492
R21095 GND.n9179 GND.n9178 70.6492
R21096 GND.n9179 GND.n774 70.6492
R21097 GND.n9187 GND.n774 70.6492
R21098 GND.n9188 GND.n9187 70.6492
R21099 GND.n9189 GND.n9188 70.6492
R21100 GND.n9189 GND.n768 70.6492
R21101 GND.n9197 GND.n768 70.6492
R21102 GND.n9198 GND.n9197 70.6492
R21103 GND.n9199 GND.n9198 70.6492
R21104 GND.n9199 GND.n762 70.6492
R21105 GND.n9207 GND.n762 70.6492
R21106 GND.n9208 GND.n9207 70.6492
R21107 GND.n9209 GND.n9208 70.6492
R21108 GND.n9209 GND.n756 70.6492
R21109 GND.n9217 GND.n756 70.6492
R21110 GND.n9218 GND.n9217 70.6492
R21111 GND.n9219 GND.n9218 70.6492
R21112 GND.n9219 GND.n750 70.6492
R21113 GND.n9227 GND.n750 70.6492
R21114 GND.n9228 GND.n9227 70.6492
R21115 GND.n9229 GND.n9228 70.6492
R21116 GND.n9229 GND.n744 70.6492
R21117 GND.n9237 GND.n744 70.6492
R21118 GND.n9238 GND.n9237 70.6492
R21119 GND.n9239 GND.n9238 70.6492
R21120 GND.n9239 GND.n738 70.6492
R21121 GND.n9247 GND.n738 70.6492
R21122 GND.n9248 GND.n9247 70.6492
R21123 GND.n9249 GND.n9248 70.6492
R21124 GND.n9249 GND.n732 70.6492
R21125 GND.n9257 GND.n732 70.6492
R21126 GND.n9258 GND.n9257 70.6492
R21127 GND.n9259 GND.n9258 70.6492
R21128 GND.n9259 GND.n726 70.6492
R21129 GND.n9267 GND.n726 70.6492
R21130 GND.n9268 GND.n9267 70.6492
R21131 GND.n9269 GND.n9268 70.6492
R21132 GND.n9269 GND.n720 70.6492
R21133 GND.n9277 GND.n720 70.6492
R21134 GND.n9278 GND.n9277 70.6492
R21135 GND.n9279 GND.n9278 70.6492
R21136 GND.n9279 GND.n714 70.6492
R21137 GND.n9287 GND.n714 70.6492
R21138 GND.n9288 GND.n9287 70.6492
R21139 GND.n9289 GND.n9288 70.6492
R21140 GND.n9289 GND.n708 70.6492
R21141 GND.n9297 GND.n708 70.6492
R21142 GND.n9298 GND.n9297 70.6492
R21143 GND.n9299 GND.n9298 70.6492
R21144 GND.n9299 GND.n702 70.6492
R21145 GND.n9307 GND.n702 70.6492
R21146 GND.n9308 GND.n9307 70.6492
R21147 GND.n9309 GND.n9308 70.6492
R21148 GND.n9309 GND.n696 70.6492
R21149 GND.n9317 GND.n696 70.6492
R21150 GND.n9318 GND.n9317 70.6492
R21151 GND.n9319 GND.n9318 70.6492
R21152 GND.n9319 GND.n690 70.6492
R21153 GND.n9327 GND.n690 70.6492
R21154 GND.n9328 GND.n9327 70.6492
R21155 GND.n9329 GND.n9328 70.6492
R21156 GND.n9329 GND.n684 70.6492
R21157 GND.n9337 GND.n684 70.6492
R21158 GND.n9338 GND.n9337 70.6492
R21159 GND.n9339 GND.n9338 70.6492
R21160 GND.n9339 GND.n678 70.6492
R21161 GND.n9347 GND.n678 70.6492
R21162 GND.n9348 GND.n9347 70.6492
R21163 GND.n9349 GND.n9348 70.6492
R21164 GND.n9349 GND.n672 70.6492
R21165 GND.n9357 GND.n672 70.6492
R21166 GND.n9358 GND.n9357 70.6492
R21167 GND.n9359 GND.n9358 70.6492
R21168 GND.n9359 GND.n666 70.6492
R21169 GND.n9367 GND.n666 70.6492
R21170 GND.n9368 GND.n9367 70.6492
R21171 GND.n9369 GND.n9368 70.6492
R21172 GND.n9369 GND.n660 70.6492
R21173 GND.n9377 GND.n660 70.6492
R21174 GND.n9378 GND.n9377 70.6492
R21175 GND.n9379 GND.n9378 70.6492
R21176 GND.n9379 GND.n654 70.6492
R21177 GND.n9387 GND.n654 70.6492
R21178 GND.n9388 GND.n9387 70.6492
R21179 GND.n9389 GND.n9388 70.6492
R21180 GND.n9389 GND.n648 70.6492
R21181 GND.n9397 GND.n648 70.6492
R21182 GND.n9398 GND.n9397 70.6492
R21183 GND.n9399 GND.n9398 70.6492
R21184 GND.n9399 GND.n642 70.6492
R21185 GND.n9407 GND.n642 70.6492
R21186 GND.n9408 GND.n9407 70.6492
R21187 GND.n9409 GND.n9408 70.6492
R21188 GND.n9409 GND.n636 70.6492
R21189 GND.n9417 GND.n636 70.6492
R21190 GND.n9418 GND.n9417 70.6492
R21191 GND.n9419 GND.n9418 70.6492
R21192 GND.n9419 GND.n630 70.6492
R21193 GND.n9427 GND.n630 70.6492
R21194 GND.n9428 GND.n9427 70.6492
R21195 GND.n9429 GND.n9428 70.6492
R21196 GND.n9429 GND.n624 70.6492
R21197 GND.n9437 GND.n624 70.6492
R21198 GND.n9438 GND.n9437 70.6492
R21199 GND.n9439 GND.n9438 70.6492
R21200 GND.n9439 GND.n618 70.6492
R21201 GND.n9447 GND.n618 70.6492
R21202 GND.n9448 GND.n9447 70.6492
R21203 GND.n9449 GND.n9448 70.6492
R21204 GND.n9449 GND.n612 70.6492
R21205 GND.n9457 GND.n612 70.6492
R21206 GND.n9458 GND.n9457 70.6492
R21207 GND.n9459 GND.n9458 70.6492
R21208 GND.n9459 GND.n606 70.6492
R21209 GND.n9467 GND.n606 70.6492
R21210 GND.n9468 GND.n9467 70.6492
R21211 GND.n9469 GND.n9468 70.6492
R21212 GND.n9469 GND.n600 70.6492
R21213 GND.n9477 GND.n600 70.6492
R21214 GND.n9478 GND.n9477 70.6492
R21215 GND.n9479 GND.n9478 70.6492
R21216 GND.n9479 GND.n594 70.6492
R21217 GND.n9487 GND.n594 70.6492
R21218 GND.n9488 GND.n9487 70.6492
R21219 GND.n9489 GND.n9488 70.6492
R21220 GND.n9489 GND.n588 70.6492
R21221 GND.n9497 GND.n588 70.6492
R21222 GND.n9498 GND.n9497 70.6492
R21223 GND.n9499 GND.n9498 70.6492
R21224 GND.n9499 GND.n582 70.6492
R21225 GND.n9507 GND.n582 70.6492
R21226 GND.n9508 GND.n9507 70.6492
R21227 GND.n9509 GND.n9508 70.6492
R21228 GND.n9509 GND.n576 70.6492
R21229 GND.n9518 GND.n576 70.6492
R21230 GND.n9519 GND.n9518 70.6492
R21231 GND.n9520 GND.n9519 70.6492
R21232 GND.n9520 GND.n571 70.6492
R21233 GND.n8222 GND.t146 66.6983
R21234 GND.n1739 GND.t59 66.6983
R21235 GND.n1760 GND.t117 66.6983
R21236 GND.n1777 GND.t83 66.6983
R21237 GND.n1798 GND.t24 66.6983
R21238 GND.n1818 GND.t141 66.6983
R21239 GND.n7109 GND.t110 66.6983
R21240 GND.n7123 GND.t46 66.6983
R21241 GND.n5459 GND.t134 66.6983
R21242 GND.n9860 GND.t132 66.6983
R21243 GND.n9870 GND.t32 66.6983
R21244 GND.n9878 GND.t95 66.6983
R21245 GND.n9809 GND.t39 66.6983
R21246 GND.n6360 GND.t55 66.6983
R21247 GND.n1376 GND.t73 66.6983
R21248 GND.n1390 GND.t122 66.6983
R21249 GND.n1406 GND.t85 66.6983
R21250 GND.n1420 GND.t35 66.6983
R21251 GND.n1436 GND.t101 66.6983
R21252 GND.n3853 GND.t65 66.6983
R21253 GND.n51 GND.t2 64.0712
R21254 GND.n5392 GND.t137 63.4983
R21255 GND.n5425 GND.t76 63.4983
R21256 GND.n9844 GND.t120 63.4983
R21257 GND.n10000 GND.t68 63.4983
R21258 GND.n53 GND.t16 63.2146
R21259 GND.n52 GND.t19 63.2146
R21260 GND.n51 GND.t269 63.2146
R21261 GND.n7915 GND.n1933 62.0895
R21262 GND.n8 GND.n7 57.37
R21263 GND.n10 GND.n9 57.37
R21264 GND.n12 GND.n11 57.37
R21265 GND.n15 GND.n14 57.37
R21266 GND.n17 GND.n16 57.37
R21267 GND.n19 GND.n18 57.37
R21268 GND.n23 GND.n22 57.37
R21269 GND.n25 GND.n24 57.37
R21270 GND.n27 GND.n26 57.37
R21271 GND.n31 GND.n30 57.37
R21272 GND.n33 GND.n32 57.37
R21273 GND.n35 GND.n34 57.37
R21274 GND.n39 GND.n38 57.37
R21275 GND.n41 GND.n40 57.37
R21276 GND.n43 GND.n42 57.37
R21277 GND.n1 GND.n0 57.37
R21278 GND.n3 GND.n2 57.37
R21279 GND.n5 GND.n4 57.37
R21280 GND.n60 GND.n59 57.37
R21281 GND.n58 GND.n57 57.37
R21282 GND.n56 GND.n55 57.37
R21283 GND.n67 GND.n66 57.37
R21284 GND.n65 GND.n64 57.37
R21285 GND.n63 GND.n62 57.37
R21286 GND.n75 GND.n74 57.37
R21287 GND.n73 GND.n72 57.37
R21288 GND.n71 GND.n70 57.37
R21289 GND.n83 GND.n82 57.37
R21290 GND.n81 GND.n80 57.37
R21291 GND.n79 GND.n78 57.37
R21292 GND.n91 GND.n90 57.37
R21293 GND.n89 GND.n88 57.37
R21294 GND.n87 GND.n86 57.37
R21295 GND.n99 GND.n98 57.37
R21296 GND.n97 GND.n96 57.37
R21297 GND.n95 GND.n94 57.37
R21298 GND.n8362 GND.n1358 57.0798
R21299 GND.n3877 GND.t42 55.9928
R21300 GND.n6343 GND.t154 55.9928
R21301 GND.n1918 GND.n1917 54.358
R21302 GND.n4750 GND.n4749 54.358
R21303 GND.n2122 GND.t143 53.9608
R21304 GND.n4761 GND.t28 53.9608
R21305 GND.n7917 GND.t98 53.9552
R21306 GND.n4759 GND.t108 53.9552
R21307 GND.n7920 GND.n7917 53.1399
R21308 GND.n2123 GND.n2122 53.1399
R21309 GND.n4762 GND.n4761 53.1399
R21310 GND.n7197 GND.n4759 53.1399
R21311 GND.n4739 GND.n4738 52.9692
R21312 GND.n5393 GND.n5392 48.6793
R21313 GND.n5426 GND.n5425 48.6793
R21314 GND.n9845 GND.n9844 48.6793
R21315 GND.n10001 GND.n10000 48.6793
R21316 GND.n3877 GND.n3876 47.5157
R21317 GND.n6343 GND.n6342 47.5157
R21318 GND.n1930 GND.n1929 46.0096
R21319 GND.n1923 GND.n1913 46.0096
R21320 GND.n4737 GND.n4736 46.0096
R21321 GND.n4753 GND.n4734 46.0096
R21322 GND.n4757 GND.n4756 44.3322
R21323 GND.n8497 GND.n1188 42.4674
R21324 GND.n8491 GND.n1188 42.4674
R21325 GND.n8491 GND.n8490 42.4674
R21326 GND.n8490 GND.n8489 42.4674
R21327 GND.n8489 GND.n1195 42.4674
R21328 GND.n8483 GND.n1195 42.4674
R21329 GND.n8483 GND.n8482 42.4674
R21330 GND.n8482 GND.n8481 42.4674
R21331 GND.n8481 GND.n1203 42.4674
R21332 GND.n8475 GND.n1203 42.4674
R21333 GND.n8475 GND.n8474 42.4674
R21334 GND.n8474 GND.n8473 42.4674
R21335 GND.n8473 GND.n1211 42.4674
R21336 GND.n8467 GND.n1211 42.4674
R21337 GND.n8467 GND.n8466 42.4674
R21338 GND.n8466 GND.n8465 42.4674
R21339 GND.n8465 GND.n1219 42.4674
R21340 GND.n8459 GND.n1219 42.4674
R21341 GND.n8459 GND.n8458 42.4674
R21342 GND.n8458 GND.n8457 42.4674
R21343 GND.n8457 GND.n1227 42.4674
R21344 GND.n8451 GND.n1227 42.4674
R21345 GND.n8451 GND.n8450 42.4674
R21346 GND.n8450 GND.n8449 42.4674
R21347 GND.n8449 GND.n1235 42.4674
R21348 GND.n8443 GND.n1235 42.4674
R21349 GND.n8443 GND.n8442 42.4674
R21350 GND.n8442 GND.n8441 42.4674
R21351 GND.n8441 GND.n1243 42.4674
R21352 GND.n8435 GND.n1243 42.4674
R21353 GND.n8435 GND.n8434 42.4674
R21354 GND.n8434 GND.n8433 42.4674
R21355 GND.n8433 GND.n1251 42.4674
R21356 GND.n8427 GND.n1251 42.4674
R21357 GND.n8427 GND.n8426 42.4674
R21358 GND.n8426 GND.n8425 42.4674
R21359 GND.n8425 GND.n1259 42.4674
R21360 GND.n8419 GND.n1259 42.4674
R21361 GND.n8419 GND.n8418 42.4674
R21362 GND.n8418 GND.n8417 42.4674
R21363 GND.n8417 GND.n1267 42.4674
R21364 GND.n8411 GND.n1267 42.4674
R21365 GND.n8411 GND.n8410 42.4674
R21366 GND.n8410 GND.n8409 42.4674
R21367 GND.n8409 GND.n1275 42.4674
R21368 GND.n8403 GND.n1275 42.4674
R21369 GND.n8403 GND.n8402 42.4674
R21370 GND.n8402 GND.n8401 42.4674
R21371 GND.n8401 GND.n1283 42.4674
R21372 GND.n8395 GND.n1283 42.4674
R21373 GND.n8395 GND.n8394 42.4674
R21374 GND.n8394 GND.n8393 42.4674
R21375 GND.n8393 GND.n1291 42.4674
R21376 GND.n8387 GND.n1291 42.4674
R21377 GND.n8387 GND.n8386 42.4674
R21378 GND.n8386 GND.n8385 42.4674
R21379 GND.n8385 GND.n1299 42.4674
R21380 GND.n8379 GND.n1299 42.4674
R21381 GND.n8379 GND.n8378 42.4674
R21382 GND.n8378 GND.n8377 42.4674
R21383 GND.n8377 GND.n1307 42.4674
R21384 GND.n8371 GND.n1307 42.4674
R21385 GND.n8371 GND.n8370 42.4674
R21386 GND.n8370 GND.n8369 42.4674
R21387 GND.n8369 GND.n1315 42.4674
R21388 GND.n8363 GND.n1315 42.4674
R21389 GND.n1920 GND.n1918 41.6274
R21390 GND.n4751 GND.n4750 41.6274
R21391 GND.n1919 GND.n1913 38.2165
R21392 GND.n8223 GND.n8222 35.8793
R21393 GND.n8005 GND.n1739 35.8793
R21394 GND.n7986 GND.n1760 35.8793
R21395 GND.n1860 GND.n1777 35.8793
R21396 GND.n1841 GND.n1798 35.8793
R21397 GND.n1822 GND.n1818 35.8793
R21398 GND.n7163 GND.n7109 35.8793
R21399 GND.n7124 GND.n7123 35.8793
R21400 GND.n5460 GND.n5459 35.8793
R21401 GND.n9971 GND.n9860 35.8793
R21402 GND.n9940 GND.n9870 35.8793
R21403 GND.n9909 GND.n9878 35.8793
R21404 GND.n9810 GND.n9809 35.8793
R21405 GND.n7708 GND.n3877 35.8793
R21406 GND.n6344 GND.n6343 35.8793
R21407 GND.n6385 GND.n6360 35.8793
R21408 GND.n8342 GND.n1376 35.8793
R21409 GND.n1391 GND.n1390 35.8793
R21410 GND.n8292 GND.n1406 35.8793
R21411 GND.n8267 GND.n1420 35.8793
R21412 GND.n8242 GND.n1436 35.8793
R21413 GND.n3872 GND.n3853 35.8793
R21414 GND.n4776 GND.n4763 34.1859
R21415 GND.n2182 GND.n2179 34.1859
R21416 GND.n9694 GND.n417 33.8941
R21417 GND.n2924 GND.n1358 32.6173
R21418 GND.n2944 GND.n2924 32.6173
R21419 GND.n2944 GND.n2912 32.6173
R21420 GND.n2953 GND.n2912 32.6173
R21421 GND.n2953 GND.n2904 32.6173
R21422 GND.n2961 GND.n2904 32.6173
R21423 GND.n2970 GND.n2892 32.6173
R21424 GND.n2970 GND.n2884 32.6173
R21425 GND.n2978 GND.n2884 32.6173
R21426 GND.n2978 GND.n2873 32.6173
R21427 GND.n2994 GND.n2873 32.6173
R21428 GND.n2994 GND.n2875 32.6173
R21429 GND.n1683 GND.n1679 32.6173
R21430 GND.n3436 GND.n1707 32.6173
R21431 GND.n3436 GND.n3435 32.6173
R21432 GND.n3435 GND.n1876 32.6173
R21433 GND.n7251 GND.n7250 32.6173
R21434 GND.n6401 GND.n6400 32.6173
R21435 GND.n6402 GND.n6401 32.6173
R21436 GND.n6402 GND.n4839 32.6173
R21437 GND.n6414 GND.n4869 32.6173
R21438 GND.n10171 GND.n358 32.6173
R21439 GND.n10171 GND.n361 32.6173
R21440 GND.n10165 GND.n361 32.6173
R21441 GND.n10165 GND.n370 32.6173
R21442 GND.n10159 GND.n370 32.6173
R21443 GND.n10159 GND.n380 32.6173
R21444 GND.n10153 GND.n389 32.6173
R21445 GND.n10147 GND.n389 32.6173
R21446 GND.n10147 GND.n399 32.6173
R21447 GND.n10141 GND.n399 32.6173
R21448 GND.n10141 GND.n408 32.6173
R21449 GND.n10135 GND.n408 32.6173
R21450 GND.n10135 GND.n417 32.6173
R21451 GND.n7977 GND.n7976 30.5925
R21452 GND.n7189 GND.n7187 30.5925
R21453 GND.n1931 GND.n1930 29.9429
R21454 GND.n4754 GND.n4753 29.9429
R21455 GND.n7972 GND.n1876 29.6817
R21456 GND.t79 GND.n1905 29.3556
R21457 GND.n8023 GND.n1707 28.3771
R21458 GND.n7183 GND.n4839 28.3771
R21459 GND.n6400 GND.t104 24.7892
R21460 GND.n10074 GND.n417 24.4631
R21461 GND.n1925 GND.n1911 24.1005
R21462 GND.n1925 GND.n1924 24.1005
R21463 GND.n4742 GND.n4741 24.1005
R21464 GND.n4743 GND.n4742 24.1005
R21465 GND.n7911 GND.n1936 22.1799
R21466 GND.n2190 GND.n1947 22.1799
R21467 GND.n7897 GND.n1955 22.1799
R21468 GND.n7890 GND.n1965 22.1799
R21469 GND.n2214 GND.n1973 22.1799
R21470 GND.n7876 GND.n1983 22.1799
R21471 GND.n2227 GND.n1991 22.1799
R21472 GND.n7862 GND.n2001 22.1799
R21473 GND.n2240 GND.n2009 22.1799
R21474 GND.n7848 GND.n2019 22.1799
R21475 GND.n2252 GND.n2027 22.1799
R21476 GND.n2252 GND.n2035 22.1799
R21477 GND.n7828 GND.n2043 22.1799
R21478 GND.n2265 GND.n2053 22.1799
R21479 GND.n7814 GND.n2061 22.1799
R21480 GND.n2278 GND.n2071 22.1799
R21481 GND.n7800 GND.n2079 22.1799
R21482 GND.n2291 GND.n2089 22.1799
R21483 GND.n7786 GND.n2097 22.1799
R21484 GND.n7779 GND.n2108 22.1799
R21485 GND.n7779 GND.n2110 22.1799
R21486 GND.n7767 GND.n2314 22.1799
R21487 GND.n5703 GND.n2327 22.1799
R21488 GND.n5712 GND.n3885 22.1799
R21489 GND.n5721 GND.n3894 22.1799
R21490 GND.n5730 GND.n3903 22.1799
R21491 GND.n5745 GND.n3913 22.1799
R21492 GND.n5758 GND.n3923 22.1799
R21493 GND.n7668 GND.n3933 22.1799
R21494 GND.n7668 GND.n3936 22.1799
R21495 GND.n7656 GND.n3950 22.1799
R21496 GND.n5807 GND.n3964 22.1799
R21497 GND.n5816 GND.n3987 22.1799
R21498 GND.n5825 GND.n3997 22.1799
R21499 GND.n5834 GND.n4007 22.1799
R21500 GND.n5849 GND.n4017 22.1799
R21501 GND.n7613 GND.n4037 22.1799
R21502 GND.n7613 GND.n4040 22.1799
R21503 GND.n7601 GND.n4054 22.1799
R21504 GND.n5910 GND.n4069 22.1799
R21505 GND.n5919 GND.n4092 22.1799
R21506 GND.n5928 GND.n4102 22.1799
R21507 GND.n5937 GND.n4112 22.1799
R21508 GND.n5965 GND.n4132 22.1799
R21509 GND.n7558 GND.n4142 22.1799
R21510 GND.n7558 GND.n4145 22.1799
R21511 GND.n7546 GND.n4159 22.1799
R21512 GND.n6022 GND.n4197 22.1799
R21513 GND.n6031 GND.n4206 22.1799
R21514 GND.n6040 GND.n4216 22.1799
R21515 GND.n6055 GND.n4226 22.1799
R21516 GND.n6068 GND.n4235 22.1799
R21517 GND.n7503 GND.n4245 22.1799
R21518 GND.n7503 GND.n4248 22.1799
R21519 GND.n6116 GND.n4277 22.1799
R21520 GND.n6125 GND.n4299 22.1799
R21521 GND.n6134 GND.n4309 22.1799
R21522 GND.n6143 GND.n4319 22.1799
R21523 GND.n6158 GND.n4329 22.1799
R21524 GND.n6171 GND.n4339 22.1799
R21525 GND.n7448 GND.n4349 22.1799
R21526 GND.n7448 GND.n4352 22.1799
R21527 GND.n7436 GND.n4366 22.1799
R21528 GND.n6209 GND.n4381 22.1799
R21529 GND.n6220 GND.n4404 22.1799
R21530 GND.n6228 GND.n5509 22.1799
R21531 GND.n6311 GND.n5499 22.1799
R21532 GND.n6303 GND.n4436 22.1799
R21533 GND.n7400 GND.n4449 22.1799
R21534 GND.n6291 GND.n4457 22.1799
R21535 GND.n6291 GND.n4465 22.1799
R21536 GND.n7380 GND.n4473 22.1799
R21537 GND.n6279 GND.n4483 22.1799
R21538 GND.n7366 GND.n4491 22.1799
R21539 GND.n6266 GND.n4501 22.1799
R21540 GND.n7352 GND.n4509 22.1799
R21541 GND.n6253 GND.n4519 22.1799
R21542 GND.n7338 GND.n4527 22.1799
R21543 GND.n7331 GND.n4538 22.1799
R21544 GND.n7331 GND.n4540 22.1799
R21545 GND.n7319 GND.n4556 22.1799
R21546 GND.n4635 GND.n4569 22.1799
R21547 GND.n7305 GND.n4577 22.1799
R21548 GND.n4648 GND.n4587 22.1799
R21549 GND.n7291 GND.n4595 22.1799
R21550 GND.n4661 GND.n4605 22.1799
R21551 GND.n7270 GND.n4623 22.1799
R21552 GND.n7258 GND.n4687 22.1799
R21553 GND.n4666 GND.t49 21.5276
R21554 GND.n7842 GND.n2025 20.8752
R21555 GND.n7834 GND.n2037 20.8752
R21556 GND.n7785 GND.n2099 20.8752
R21557 GND.n7773 GND.n2305 20.8752
R21558 GND.n7674 GND.n3925 20.8752
R21559 GND.n7662 GND.n3944 20.8752
R21560 GND.n7619 GND.n4029 20.8752
R21561 GND.n7607 GND.n4048 20.8752
R21562 GND.n7564 GND.n4134 20.8752
R21563 GND.n7552 GND.n4153 20.8752
R21564 GND.n7509 GND.n4237 20.8752
R21565 GND.n7497 GND.n4256 20.8752
R21566 GND.n7454 GND.n4341 20.8752
R21567 GND.n7442 GND.n4360 20.8752
R21568 GND.n7394 GND.n4455 20.8752
R21569 GND.n7386 GND.n4467 20.8752
R21570 GND.n7337 GND.n4529 20.8752
R21571 GND.n7325 GND.n4547 20.8752
R21572 GND.n7276 GND.n4614 20.8752
R21573 GND.n7264 GND.n4676 20.8752
R21574 GND.n7915 GND.n7914 20.7615
R21575 GND.n4769 GND.n4757 20.7615
R21576 GND.n2875 GND.n2863 20.2229
R21577 GND.n3005 GND.n3004 20.2229
R21578 GND.n3017 GND.n2862 20.2229
R21579 GND.n3018 GND.n2848 20.2229
R21580 GND.n3027 GND.n2850 20.2229
R21581 GND.n3036 GND.n2840 20.2229
R21582 GND.n3035 GND.n2834 20.2229
R21583 GND.n3045 GND.n3044 20.2229
R21584 GND.n3060 GND.n2825 20.2229
R21585 GND.n3071 GND.n2813 20.2229
R21586 GND.n3070 GND.n2816 20.2229
R21587 GND.n3081 GND.n2806 20.2229
R21588 GND.n3082 GND.n2795 20.2229
R21589 GND.n3097 GND.n2797 20.2229
R21590 GND.n3108 GND.n2785 20.2229
R21591 GND.n3107 GND.n2787 20.2229
R21592 GND.n3118 GND.n2777 20.2229
R21593 GND.n3119 GND.n2765 20.2229
R21594 GND.n3135 GND.n2768 20.2229
R21595 GND.n3145 GND.n2757 20.2229
R21596 GND.n3156 GND.n2749 20.2229
R21597 GND.n3158 GND.n2738 20.2229
R21598 GND.n3173 GND.n2740 20.2229
R21599 GND.n3184 GND.n2728 20.2229
R21600 GND.n3183 GND.n2730 20.2229
R21601 GND.n3194 GND.n2721 20.2229
R21602 GND.n3195 GND.n2709 20.2229
R21603 GND.n3210 GND.n2711 20.2229
R21604 GND.n3221 GND.n2698 20.2229
R21605 GND.n3231 GND.n2691 20.2229
R21606 GND.n3232 GND.n2680 20.2229
R21607 GND.n3247 GND.n2682 20.2229
R21608 GND.n3258 GND.n2670 20.2229
R21609 GND.n3257 GND.n2672 20.2229
R21610 GND.n3268 GND.n2662 20.2229
R21611 GND.n3269 GND.n2650 20.2229
R21612 GND.n3284 GND.n2653 20.2229
R21613 GND.n3296 GND.n2640 20.2229
R21614 GND.n3295 GND.n2642 20.2229
R21615 GND.n3306 GND.n2633 20.2229
R21616 GND.n3308 GND.n2622 20.2229
R21617 GND.n3320 GND.n2624 20.2229
R21618 GND.n3328 GND.n2615 20.2229
R21619 GND.n3327 GND.n2618 20.2229
R21620 GND.n3541 GND.n2610 20.2229
R21621 GND.n3542 GND.n1533 20.2229
R21622 GND.n8123 GND.n1535 20.2229
R21623 GND.n2600 GND.n2599 20.2229
R21624 GND.n3556 GND.n2596 20.2229
R21625 GND.n3559 GND.n1552 20.2229
R21626 GND.n8116 GND.n1555 20.2229
R21627 GND.n3570 GND.n2583 20.2229
R21628 GND.n3575 GND.n2586 20.2229
R21629 GND.n3572 GND.n2572 20.2229
R21630 GND.n3585 GND.n2573 20.2229
R21631 GND.n2577 GND.n2565 20.2229
R21632 GND.n3595 GND.n2561 20.2229
R21633 GND.n3601 GND.n2563 20.2229
R21634 GND.n3598 GND.n2550 20.2229
R21635 GND.n3611 GND.n2551 20.2229
R21636 GND.n2555 GND.n2544 20.2229
R21637 GND.n3627 GND.n2542 20.2229
R21638 GND.n3623 GND.n2529 20.2229
R21639 GND.n3637 GND.n2531 20.2229
R21640 GND.n2534 GND.n2523 20.2229
R21641 GND.n3647 GND.n2518 20.2229
R21642 GND.n3653 GND.n2520 20.2229
R21643 GND.n3650 GND.n2508 20.2229
R21644 GND.n3663 GND.n2509 20.2229
R21645 GND.n2512 GND.n2502 20.2229
R21646 GND.n3673 GND.n2496 20.2229
R21647 GND.n3678 GND.n2499 20.2229
R21648 GND.n3675 GND.n2485 20.2229
R21649 GND.n3688 GND.n2486 20.2229
R21650 GND.n2490 GND.n2478 20.2229
R21651 GND.n3698 GND.n2474 20.2229
R21652 GND.n3704 GND.n2476 20.2229
R21653 GND.n3701 GND.n2463 20.2229
R21654 GND.n3714 GND.n2464 20.2229
R21655 GND.n2468 GND.n2457 20.2229
R21656 GND.n3724 GND.n2453 20.2229
R21657 GND.n3730 GND.n2455 20.2229
R21658 GND.n3726 GND.n2444 20.2229
R21659 GND.n3473 GND.n2438 20.2229
R21660 GND.n3750 GND.n2433 20.2229
R21661 GND.n3756 GND.n2435 20.2229
R21662 GND.n3753 GND.n2423 20.2229
R21663 GND.n3766 GND.n2424 20.2229
R21664 GND.n2427 GND.n2417 20.2229
R21665 GND.n3776 GND.n2411 20.2229
R21666 GND.n3781 GND.n2414 20.2229
R21667 GND.n3778 GND.n2400 20.2229
R21668 GND.n3791 GND.n2401 20.2229
R21669 GND.n2405 GND.n2393 20.2229
R21670 GND.n3801 GND.n2389 20.2229
R21671 GND.n3807 GND.n2391 20.2229
R21672 GND.n3817 GND.n2379 20.2229
R21673 GND.n2383 GND.n2372 20.2229
R21674 GND.n3828 GND.n2368 20.2229
R21675 GND.n3834 GND.n2370 20.2229
R21676 GND.n3830 GND.n2362 20.2229
R21677 GND.n3843 GND.n1676 20.2229
R21678 GND.n8026 GND.n1679 20.2229
R21679 GND.n6416 GND.n6414 20.2229
R21680 GND.n7091 GND.n4882 20.2229
R21681 GND.n7084 GND.n4885 20.2229
R21682 GND.n7083 GND.n4896 20.2229
R21683 GND.n4906 GND.n4905 20.2229
R21684 GND.n7077 GND.n7076 20.2229
R21685 GND.n6473 GND.n4909 20.2229
R21686 GND.n6479 GND.n4926 20.2229
R21687 GND.n7064 GND.n4935 20.2229
R21688 GND.n6487 GND.n4938 20.2229
R21689 GND.n7058 GND.n4946 20.2229
R21690 GND.n6493 GND.n4949 20.2229
R21691 GND.n7052 GND.n4956 20.2229
R21692 GND.n6501 GND.n4959 20.2229
R21693 GND.n7046 GND.n4967 20.2229
R21694 GND.n6507 GND.n4970 20.2229
R21695 GND.n7040 GND.n4977 20.2229
R21696 GND.n6516 GND.n4980 20.2229
R21697 GND.n7034 GND.n4988 20.2229
R21698 GND.n6675 GND.n4991 20.2229
R21699 GND.n6669 GND.n5000 20.2229
R21700 GND.n7022 GND.n5008 20.2229
R21701 GND.n6663 GND.n5011 20.2229
R21702 GND.n7016 GND.n5018 20.2229
R21703 GND.n6657 GND.n5021 20.2229
R21704 GND.n7010 GND.n5029 20.2229
R21705 GND.n6651 GND.n5032 20.2229
R21706 GND.n7004 GND.n5039 20.2229
R21707 GND.n6645 GND.n5042 20.2229
R21708 GND.n6998 GND.n5050 20.2229
R21709 GND.n6639 GND.n5053 20.2229
R21710 GND.n6992 GND.n5060 20.2229
R21711 GND.n6633 GND.n5063 20.2229
R21712 GND.n6986 GND.n5071 20.2229
R21713 GND.n6627 GND.n5074 20.2229
R21714 GND.n6980 GND.n5081 20.2229
R21715 GND.n6621 GND.n5084 20.2229
R21716 GND.n6974 GND.n5092 20.2229
R21717 GND.n6615 GND.n5095 20.2229
R21718 GND.n6968 GND.n5102 20.2229
R21719 GND.n6609 GND.n5105 20.2229
R21720 GND.n6962 GND.n5113 20.2229
R21721 GND.n6956 GND.n5123 20.2229
R21722 GND.n6597 GND.n5126 20.2229
R21723 GND.n6950 GND.n5134 20.2229
R21724 GND.n6591 GND.n5137 20.2229
R21725 GND.n6944 GND.n5144 20.2229
R21726 GND.n6585 GND.n5147 20.2229
R21727 GND.n6938 GND.n5155 20.2229
R21728 GND.n6579 GND.n5158 20.2229
R21729 GND.n6932 GND.n5165 20.2229
R21730 GND.n6754 GND.n5168 20.2229
R21731 GND.n6769 GND.n5177 20.2229
R21732 GND.n6920 GND.n5184 20.2229
R21733 GND.n6916 GND.n5187 20.2229
R21734 GND.n6915 GND.n5192 20.2229
R21735 GND.n6779 GND.n5286 20.2229
R21736 GND.n10310 GND.n108 20.2229
R21737 GND.n6788 GND.n110 20.2229
R21738 GND.n6787 GND.n5269 20.2229
R21739 GND.n6902 GND.n6901 20.2229
R21740 GND.n10303 GND.n127 20.2229
R21741 GND.n6895 GND.n130 20.2229
R21742 GND.n10297 GND.n139 20.2229
R21743 GND.n6889 GND.n142 20.2229
R21744 GND.n10291 GND.n149 20.2229
R21745 GND.n6883 GND.n152 20.2229
R21746 GND.n10285 GND.n159 20.2229
R21747 GND.n6877 GND.n162 20.2229
R21748 GND.n10279 GND.n170 20.2229
R21749 GND.n6871 GND.n173 20.2229
R21750 GND.n10273 GND.n180 20.2229
R21751 GND.n6865 GND.n183 20.2229
R21752 GND.n10267 GND.n191 20.2229
R21753 GND.n10261 GND.n201 20.2229
R21754 GND.n6853 GND.n204 20.2229
R21755 GND.n10255 GND.n212 20.2229
R21756 GND.n6847 GND.n215 20.2229
R21757 GND.n10249 GND.n222 20.2229
R21758 GND.n6841 GND.n225 20.2229
R21759 GND.n10243 GND.n233 20.2229
R21760 GND.n6835 GND.n236 20.2229
R21761 GND.n10237 GND.n243 20.2229
R21762 GND.n9727 GND.n246 20.2229
R21763 GND.n9735 GND.n256 20.2229
R21764 GND.n10225 GND.n263 20.2229
R21765 GND.n9742 GND.n266 20.2229
R21766 GND.n10219 GND.n274 20.2229
R21767 GND.n9750 GND.n277 20.2229
R21768 GND.n10213 GND.n284 20.2229
R21769 GND.n9757 GND.n287 20.2229
R21770 GND.n10207 GND.n295 20.2229
R21771 GND.n9765 GND.n298 20.2229
R21772 GND.n10201 GND.n305 20.2229
R21773 GND.n9772 GND.n308 20.2229
R21774 GND.n10195 GND.n316 20.2229
R21775 GND.n9780 GND.n319 20.2229
R21776 GND.n10189 GND.n326 20.2229
R21777 GND.n9787 GND.n329 20.2229
R21778 GND.n10183 GND.n337 20.2229
R21779 GND.n10104 GND.n340 20.2229
R21780 GND.n10177 GND.n347 20.2229
R21781 GND.n358 GND.n350 20.2229
R21782 GND.n1916 GND.t89 19.8005
R21783 GND.n1916 GND.t114 19.8005
R21784 GND.n1915 GND.t80 19.8005
R21785 GND.n1915 GND.t129 19.8005
R21786 GND.n1914 GND.t53 19.8005
R21787 GND.n1914 GND.t92 19.8005
R21788 GND.n4748 GND.t62 19.8005
R21789 GND.n4748 GND.t126 19.8005
R21790 GND.n4747 GND.t50 19.8005
R21791 GND.n4747 GND.t150 19.8005
R21792 GND.n4746 GND.t71 19.8005
R21793 GND.n4746 GND.t105 19.8005
R21794 GND.n2237 GND.n2017 19.5706
R21795 GND.n2262 GND.n2045 19.5706
R21796 GND.n5694 GND.n2316 19.5706
R21797 GND.n7680 GND.n3915 19.5706
R21798 GND.n5798 GND.n5797 19.5706
R21799 GND.n7625 GND.n4019 19.5706
R21800 GND.n7570 GND.n4124 19.5706
R21801 GND.n6004 GND.n4162 19.5706
R21802 GND.n6107 GND.n4265 19.5706
R21803 GND.n7460 GND.n4331 19.5706
R21804 GND.n6203 GND.n4369 19.5706
R21805 GND.n6302 GND.n4447 19.5706
R21806 GND.n7345 GND.n7344 19.5706
R21807 GND.n4632 GND.n4558 19.5706
R21808 GND.n4768 GND.n4689 19.5706
R21809 GND.n1910 GND.n1909 19.5087
R21810 GND.n1928 GND.n1910 19.5087
R21811 GND.n1922 GND.n1921 19.5087
R21812 GND.n4752 GND.n4745 19.5087
R21813 GND.n8216 GND.n8215 19.3944
R21814 GND.n8215 GND.n8214 19.3944
R21815 GND.n8214 GND.n1457 19.3944
R21816 GND.n8210 GND.n1457 19.3944
R21817 GND.n8210 GND.n8209 19.3944
R21818 GND.n8209 GND.n8208 19.3944
R21819 GND.n8208 GND.n1462 19.3944
R21820 GND.n8204 GND.n1462 19.3944
R21821 GND.n8204 GND.n8203 19.3944
R21822 GND.n8203 GND.n8202 19.3944
R21823 GND.n8202 GND.n1467 19.3944
R21824 GND.n8198 GND.n1467 19.3944
R21825 GND.n8198 GND.n8197 19.3944
R21826 GND.n8197 GND.n8196 19.3944
R21827 GND.n8196 GND.n1472 19.3944
R21828 GND.n8192 GND.n1472 19.3944
R21829 GND.n8192 GND.n8191 19.3944
R21830 GND.n8191 GND.n8190 19.3944
R21831 GND.n8190 GND.n1477 19.3944
R21832 GND.n8186 GND.n1477 19.3944
R21833 GND.n8186 GND.n8185 19.3944
R21834 GND.n8185 GND.n8184 19.3944
R21835 GND.n8184 GND.n1482 19.3944
R21836 GND.n8180 GND.n1482 19.3944
R21837 GND.n8180 GND.n8179 19.3944
R21838 GND.n8179 GND.n8178 19.3944
R21839 GND.n8178 GND.n1487 19.3944
R21840 GND.n8174 GND.n1487 19.3944
R21841 GND.n8174 GND.n8173 19.3944
R21842 GND.n8173 GND.n8172 19.3944
R21843 GND.n8172 GND.n1492 19.3944
R21844 GND.n8168 GND.n1492 19.3944
R21845 GND.n8168 GND.n8167 19.3944
R21846 GND.n8167 GND.n8166 19.3944
R21847 GND.n8166 GND.n1497 19.3944
R21848 GND.n8162 GND.n1497 19.3944
R21849 GND.n8162 GND.n8161 19.3944
R21850 GND.n8161 GND.n8160 19.3944
R21851 GND.n8160 GND.n1502 19.3944
R21852 GND.n8156 GND.n1502 19.3944
R21853 GND.n8156 GND.n8155 19.3944
R21854 GND.n8155 GND.n8154 19.3944
R21855 GND.n8154 GND.n1507 19.3944
R21856 GND.n8150 GND.n1507 19.3944
R21857 GND.n8150 GND.n8149 19.3944
R21858 GND.n8149 GND.n8148 19.3944
R21859 GND.n8148 GND.n1512 19.3944
R21860 GND.n8144 GND.n1512 19.3944
R21861 GND.n8144 GND.n8143 19.3944
R21862 GND.n8143 GND.n8142 19.3944
R21863 GND.n8142 GND.n1517 19.3944
R21864 GND.n8138 GND.n1517 19.3944
R21865 GND.n8138 GND.n8137 19.3944
R21866 GND.n8137 GND.n8136 19.3944
R21867 GND.n8136 GND.n1522 19.3944
R21868 GND.n8132 GND.n1522 19.3944
R21869 GND.n8132 GND.n8131 19.3944
R21870 GND.n8131 GND.n8130 19.3944
R21871 GND.n8130 GND.n1527 19.3944
R21872 GND.n8126 GND.n1527 19.3944
R21873 GND.n8126 GND.n8125 19.3944
R21874 GND.n8125 GND.n1531 19.3944
R21875 GND.n2594 GND.n1531 19.3944
R21876 GND.n3561 GND.n2594 19.3944
R21877 GND.n3562 GND.n3561 19.3944
R21878 GND.n3562 GND.n2590 19.3944
R21879 GND.n3568 GND.n2590 19.3944
R21880 GND.n3568 GND.n3567 19.3944
R21881 GND.n3567 GND.n2570 19.3944
R21882 GND.n3587 GND.n2570 19.3944
R21883 GND.n3587 GND.n2568 19.3944
R21884 GND.n3593 GND.n2568 19.3944
R21885 GND.n3593 GND.n3592 19.3944
R21886 GND.n3592 GND.n2548 19.3944
R21887 GND.n3613 GND.n2548 19.3944
R21888 GND.n3613 GND.n2546 19.3944
R21889 GND.n3619 GND.n2546 19.3944
R21890 GND.n3619 GND.n3618 19.3944
R21891 GND.n3618 GND.n2527 19.3944
R21892 GND.n3639 GND.n2527 19.3944
R21893 GND.n3639 GND.n2525 19.3944
R21894 GND.n3645 GND.n2525 19.3944
R21895 GND.n3645 GND.n3644 19.3944
R21896 GND.n3644 GND.n2506 19.3944
R21897 GND.n3665 GND.n2506 19.3944
R21898 GND.n3665 GND.n2504 19.3944
R21899 GND.n3671 GND.n2504 19.3944
R21900 GND.n3671 GND.n3670 19.3944
R21901 GND.n3670 GND.n2483 19.3944
R21902 GND.n3690 GND.n2483 19.3944
R21903 GND.n3690 GND.n2481 19.3944
R21904 GND.n3696 GND.n2481 19.3944
R21905 GND.n3696 GND.n3695 19.3944
R21906 GND.n3695 GND.n2461 19.3944
R21907 GND.n3716 GND.n2461 19.3944
R21908 GND.n3716 GND.n2459 19.3944
R21909 GND.n3722 GND.n2459 19.3944
R21910 GND.n3722 GND.n3721 19.3944
R21911 GND.n3721 GND.n2442 19.3944
R21912 GND.n3742 GND.n2442 19.3944
R21913 GND.n3742 GND.n2440 19.3944
R21914 GND.n3748 GND.n2440 19.3944
R21915 GND.n3748 GND.n3747 19.3944
R21916 GND.n3747 GND.n2421 19.3944
R21917 GND.n3768 GND.n2421 19.3944
R21918 GND.n3768 GND.n2419 19.3944
R21919 GND.n3774 GND.n2419 19.3944
R21920 GND.n3774 GND.n3773 19.3944
R21921 GND.n3773 GND.n2398 19.3944
R21922 GND.n3793 GND.n2398 19.3944
R21923 GND.n3793 GND.n2396 19.3944
R21924 GND.n3799 GND.n2396 19.3944
R21925 GND.n3799 GND.n3798 19.3944
R21926 GND.n3798 GND.n2376 19.3944
R21927 GND.n3819 GND.n2376 19.3944
R21928 GND.n3819 GND.n2374 19.3944
R21929 GND.n3826 GND.n2374 19.3944
R21930 GND.n3826 GND.n3825 19.3944
R21931 GND.n3825 GND.n2360 19.3944
R21932 GND.n3845 GND.n2360 19.3944
R21933 GND.n3846 GND.n3845 19.3944
R21934 GND.n8237 GND.n8236 19.3944
R21935 GND.n8236 GND.n8235 19.3944
R21936 GND.n8235 GND.n1442 19.3944
R21937 GND.n8231 GND.n1442 19.3944
R21938 GND.n8231 GND.n8230 19.3944
R21939 GND.n8230 GND.n8229 19.3944
R21940 GND.n8229 GND.n1448 19.3944
R21941 GND.n8225 GND.n1448 19.3944
R21942 GND.n8225 GND.n8224 19.3944
R21943 GND.n2931 GND.n2930 19.3944
R21944 GND.n2931 GND.n2922 19.3944
R21945 GND.n2947 GND.n2922 19.3944
R21946 GND.n2949 GND.n2947 19.3944
R21947 GND.n2949 GND.n2948 19.3944
R21948 GND.n2948 GND.n2902 19.3944
R21949 GND.n2964 GND.n2902 19.3944
R21950 GND.n2966 GND.n2964 19.3944
R21951 GND.n2966 GND.n2965 19.3944
R21952 GND.n2965 GND.n2882 19.3944
R21953 GND.n2981 GND.n2882 19.3944
R21954 GND.n2990 GND.n2981 19.3944
R21955 GND.n2990 GND.n2989 19.3944
R21956 GND.n2989 GND.n2988 19.3944
R21957 GND.n2988 GND.n2859 19.3944
R21958 GND.n3020 GND.n2859 19.3944
R21959 GND.n3023 GND.n3020 19.3944
R21960 GND.n3023 GND.n3022 19.3944
R21961 GND.n3022 GND.n2832 19.3944
R21962 GND.n3047 GND.n2832 19.3944
R21963 GND.n3056 GND.n3047 19.3944
R21964 GND.n3056 GND.n3055 19.3944
R21965 GND.n3055 GND.n3054 19.3944
R21966 GND.n3054 GND.n2804 19.3944
R21967 GND.n3084 GND.n2804 19.3944
R21968 GND.n3093 GND.n3084 19.3944
R21969 GND.n3093 GND.n3092 19.3944
R21970 GND.n3092 GND.n3091 19.3944
R21971 GND.n3091 GND.n2775 19.3944
R21972 GND.n3121 GND.n2775 19.3944
R21973 GND.n3131 GND.n3121 19.3944
R21974 GND.n3131 GND.n3130 19.3944
R21975 GND.n3130 GND.n3129 19.3944
R21976 GND.n3129 GND.n2747 19.3944
R21977 GND.n3160 GND.n2747 19.3944
R21978 GND.n3169 GND.n3160 19.3944
R21979 GND.n3169 GND.n3168 19.3944
R21980 GND.n3168 GND.n3167 19.3944
R21981 GND.n3167 GND.n2718 19.3944
R21982 GND.n3197 GND.n2718 19.3944
R21983 GND.n3206 GND.n3197 19.3944
R21984 GND.n3206 GND.n3205 19.3944
R21985 GND.n3205 GND.n3204 19.3944
R21986 GND.n3204 GND.n2689 19.3944
R21987 GND.n3234 GND.n2689 19.3944
R21988 GND.n3243 GND.n3234 19.3944
R21989 GND.n3243 GND.n3242 19.3944
R21990 GND.n3242 GND.n3241 19.3944
R21991 GND.n3241 GND.n2660 19.3944
R21992 GND.n3271 GND.n2660 19.3944
R21993 GND.n3280 GND.n3271 19.3944
R21994 GND.n3280 GND.n3279 19.3944
R21995 GND.n3279 GND.n3278 19.3944
R21996 GND.n3278 GND.n2631 19.3944
R21997 GND.n3310 GND.n2631 19.3944
R21998 GND.n3316 GND.n3310 19.3944
R21999 GND.n3316 GND.n3315 19.3944
R22000 GND.n3315 GND.n3314 19.3944
R22001 GND.n3314 GND.n2604 19.3944
R22002 GND.n3547 GND.n2604 19.3944
R22003 GND.n3548 GND.n3547 19.3944
R22004 GND.n3549 GND.n3548 19.3944
R22005 GND.n3549 GND.n2598 19.3944
R22006 GND.n2598 GND.n1562 19.3944
R22007 GND.n8112 GND.n1562 19.3944
R22008 GND.n8112 GND.n8111 19.3944
R22009 GND.n8111 GND.n8110 19.3944
R22010 GND.n8110 GND.n1565 19.3944
R22011 GND.n8106 GND.n1565 19.3944
R22012 GND.n8106 GND.n8105 19.3944
R22013 GND.n8105 GND.n8104 19.3944
R22014 GND.n8104 GND.n1573 19.3944
R22015 GND.n8100 GND.n1573 19.3944
R22016 GND.n8100 GND.n8099 19.3944
R22017 GND.n8099 GND.n8098 19.3944
R22018 GND.n8098 GND.n1581 19.3944
R22019 GND.n8094 GND.n1581 19.3944
R22020 GND.n8094 GND.n8093 19.3944
R22021 GND.n8093 GND.n8092 19.3944
R22022 GND.n8092 GND.n1589 19.3944
R22023 GND.n8088 GND.n1589 19.3944
R22024 GND.n8088 GND.n8087 19.3944
R22025 GND.n8087 GND.n8086 19.3944
R22026 GND.n8086 GND.n1597 19.3944
R22027 GND.n8082 GND.n1597 19.3944
R22028 GND.n8082 GND.n8081 19.3944
R22029 GND.n8081 GND.n8080 19.3944
R22030 GND.n8080 GND.n1605 19.3944
R22031 GND.n8076 GND.n1605 19.3944
R22032 GND.n8076 GND.n8075 19.3944
R22033 GND.n8075 GND.n8074 19.3944
R22034 GND.n8074 GND.n1613 19.3944
R22035 GND.n8070 GND.n1613 19.3944
R22036 GND.n8070 GND.n8069 19.3944
R22037 GND.n8069 GND.n8068 19.3944
R22038 GND.n8068 GND.n1621 19.3944
R22039 GND.n8064 GND.n1621 19.3944
R22040 GND.n8064 GND.n8063 19.3944
R22041 GND.n8063 GND.n8062 19.3944
R22042 GND.n8062 GND.n1629 19.3944
R22043 GND.n8058 GND.n1629 19.3944
R22044 GND.n8058 GND.n8057 19.3944
R22045 GND.n8057 GND.n8056 19.3944
R22046 GND.n8056 GND.n1637 19.3944
R22047 GND.n8052 GND.n1637 19.3944
R22048 GND.n8052 GND.n8051 19.3944
R22049 GND.n8051 GND.n8050 19.3944
R22050 GND.n8050 GND.n1645 19.3944
R22051 GND.n8046 GND.n1645 19.3944
R22052 GND.n8046 GND.n8045 19.3944
R22053 GND.n8045 GND.n8044 19.3944
R22054 GND.n8044 GND.n1653 19.3944
R22055 GND.n8040 GND.n1653 19.3944
R22056 GND.n8040 GND.n8039 19.3944
R22057 GND.n8039 GND.n8038 19.3944
R22058 GND.n8038 GND.n1661 19.3944
R22059 GND.n8034 GND.n1661 19.3944
R22060 GND.n8034 GND.n8033 19.3944
R22061 GND.n8033 GND.n8032 19.3944
R22062 GND.n8032 GND.n1669 19.3944
R22063 GND.n8028 GND.n1669 19.3944
R22064 GND.n8021 GND.n1723 19.3944
R22065 GND.n8017 GND.n1723 19.3944
R22066 GND.n8017 GND.n8016 19.3944
R22067 GND.n8016 GND.n8015 19.3944
R22068 GND.n8015 GND.n1730 19.3944
R22069 GND.n8011 GND.n1730 19.3944
R22070 GND.n8011 GND.n8010 19.3944
R22071 GND.n8010 GND.n8009 19.3944
R22072 GND.n8009 GND.n1736 19.3944
R22073 GND.n8004 GND.n8003 19.3944
R22074 GND.n8003 GND.n1744 19.3944
R22075 GND.n7999 GND.n1744 19.3944
R22076 GND.n7999 GND.n7998 19.3944
R22077 GND.n7998 GND.n7997 19.3944
R22078 GND.n7997 GND.n1750 19.3944
R22079 GND.n7993 GND.n1750 19.3944
R22080 GND.n7993 GND.n7992 19.3944
R22081 GND.n7992 GND.n7991 19.3944
R22082 GND.n7991 GND.n1756 19.3944
R22083 GND.n7987 GND.n1756 19.3944
R22084 GND.n7985 GND.n7984 19.3944
R22085 GND.n7984 GND.n1764 19.3944
R22086 GND.n7980 GND.n1764 19.3944
R22087 GND.n7980 GND.n7979 19.3944
R22088 GND.n1866 GND.n1768 19.3944
R22089 GND.n1866 GND.n1865 19.3944
R22090 GND.n1865 GND.n1864 19.3944
R22091 GND.n1864 GND.n1774 19.3944
R22092 GND.n1859 GND.n1858 19.3944
R22093 GND.n1858 GND.n1782 19.3944
R22094 GND.n1854 GND.n1782 19.3944
R22095 GND.n1854 GND.n1853 19.3944
R22096 GND.n1853 GND.n1852 19.3944
R22097 GND.n1852 GND.n1788 19.3944
R22098 GND.n1848 GND.n1788 19.3944
R22099 GND.n1848 GND.n1847 19.3944
R22100 GND.n1847 GND.n1846 19.3944
R22101 GND.n1846 GND.n1794 19.3944
R22102 GND.n1842 GND.n1794 19.3944
R22103 GND.n1840 GND.n1839 19.3944
R22104 GND.n1839 GND.n1802 19.3944
R22105 GND.n1835 GND.n1802 19.3944
R22106 GND.n1835 GND.n1834 19.3944
R22107 GND.n1834 GND.n1833 19.3944
R22108 GND.n1833 GND.n1808 19.3944
R22109 GND.n1829 GND.n1808 19.3944
R22110 GND.n1829 GND.n1828 19.3944
R22111 GND.n1828 GND.n1827 19.3944
R22112 GND.n1827 GND.n1814 19.3944
R22113 GND.n1823 GND.n1814 19.3944
R22114 GND.n9526 GND.n569 19.3944
R22115 GND.n9532 GND.n569 19.3944
R22116 GND.n9532 GND.n567 19.3944
R22117 GND.n9536 GND.n567 19.3944
R22118 GND.n9536 GND.n563 19.3944
R22119 GND.n9542 GND.n563 19.3944
R22120 GND.n9542 GND.n561 19.3944
R22121 GND.n9546 GND.n561 19.3944
R22122 GND.n9546 GND.n557 19.3944
R22123 GND.n9552 GND.n557 19.3944
R22124 GND.n9552 GND.n555 19.3944
R22125 GND.n9556 GND.n555 19.3944
R22126 GND.n9556 GND.n551 19.3944
R22127 GND.n9562 GND.n551 19.3944
R22128 GND.n9562 GND.n549 19.3944
R22129 GND.n9566 GND.n549 19.3944
R22130 GND.n9566 GND.n545 19.3944
R22131 GND.n9572 GND.n545 19.3944
R22132 GND.n9572 GND.n543 19.3944
R22133 GND.n9576 GND.n543 19.3944
R22134 GND.n9576 GND.n539 19.3944
R22135 GND.n9582 GND.n539 19.3944
R22136 GND.n9582 GND.n537 19.3944
R22137 GND.n9586 GND.n537 19.3944
R22138 GND.n9586 GND.n533 19.3944
R22139 GND.n9592 GND.n533 19.3944
R22140 GND.n9592 GND.n531 19.3944
R22141 GND.n9596 GND.n531 19.3944
R22142 GND.n9596 GND.n527 19.3944
R22143 GND.n9602 GND.n527 19.3944
R22144 GND.n9602 GND.n525 19.3944
R22145 GND.n9606 GND.n525 19.3944
R22146 GND.n9606 GND.n521 19.3944
R22147 GND.n9612 GND.n521 19.3944
R22148 GND.n9612 GND.n519 19.3944
R22149 GND.n9616 GND.n519 19.3944
R22150 GND.n9616 GND.n515 19.3944
R22151 GND.n9622 GND.n515 19.3944
R22152 GND.n9622 GND.n513 19.3944
R22153 GND.n9626 GND.n513 19.3944
R22154 GND.n9626 GND.n509 19.3944
R22155 GND.n9632 GND.n509 19.3944
R22156 GND.n9632 GND.n507 19.3944
R22157 GND.n9636 GND.n507 19.3944
R22158 GND.n9636 GND.n503 19.3944
R22159 GND.n9642 GND.n503 19.3944
R22160 GND.n9642 GND.n501 19.3944
R22161 GND.n9646 GND.n501 19.3944
R22162 GND.n9646 GND.n497 19.3944
R22163 GND.n9652 GND.n497 19.3944
R22164 GND.n9652 GND.n495 19.3944
R22165 GND.n9656 GND.n495 19.3944
R22166 GND.n9656 GND.n491 19.3944
R22167 GND.n9662 GND.n491 19.3944
R22168 GND.n9662 GND.n489 19.3944
R22169 GND.n9666 GND.n489 19.3944
R22170 GND.n9666 GND.n485 19.3944
R22171 GND.n9672 GND.n485 19.3944
R22172 GND.n9672 GND.n483 19.3944
R22173 GND.n9676 GND.n483 19.3944
R22174 GND.n9676 GND.n479 19.3944
R22175 GND.n9682 GND.n479 19.3944
R22176 GND.n9682 GND.n477 19.3944
R22177 GND.n9690 GND.n477 19.3944
R22178 GND.n9690 GND.n9689 19.3944
R22179 GND.n9689 GND.n474 19.3944
R22180 GND.n8501 GND.n1186 19.3944
R22181 GND.n8501 GND.n1184 19.3944
R22182 GND.n8505 GND.n1184 19.3944
R22183 GND.n8505 GND.n1180 19.3944
R22184 GND.n8511 GND.n1180 19.3944
R22185 GND.n8511 GND.n1178 19.3944
R22186 GND.n8515 GND.n1178 19.3944
R22187 GND.n8515 GND.n1174 19.3944
R22188 GND.n8521 GND.n1174 19.3944
R22189 GND.n8521 GND.n1172 19.3944
R22190 GND.n8525 GND.n1172 19.3944
R22191 GND.n8525 GND.n1168 19.3944
R22192 GND.n8531 GND.n1168 19.3944
R22193 GND.n8531 GND.n1166 19.3944
R22194 GND.n8535 GND.n1166 19.3944
R22195 GND.n8535 GND.n1162 19.3944
R22196 GND.n8541 GND.n1162 19.3944
R22197 GND.n8541 GND.n1160 19.3944
R22198 GND.n8545 GND.n1160 19.3944
R22199 GND.n8545 GND.n1156 19.3944
R22200 GND.n8551 GND.n1156 19.3944
R22201 GND.n8551 GND.n1154 19.3944
R22202 GND.n8555 GND.n1154 19.3944
R22203 GND.n8555 GND.n1150 19.3944
R22204 GND.n8561 GND.n1150 19.3944
R22205 GND.n8561 GND.n1148 19.3944
R22206 GND.n8565 GND.n1148 19.3944
R22207 GND.n8565 GND.n1144 19.3944
R22208 GND.n8571 GND.n1144 19.3944
R22209 GND.n8571 GND.n1142 19.3944
R22210 GND.n8575 GND.n1142 19.3944
R22211 GND.n8575 GND.n1138 19.3944
R22212 GND.n8581 GND.n1138 19.3944
R22213 GND.n8581 GND.n1136 19.3944
R22214 GND.n8585 GND.n1136 19.3944
R22215 GND.n8585 GND.n1132 19.3944
R22216 GND.n8591 GND.n1132 19.3944
R22217 GND.n8591 GND.n1130 19.3944
R22218 GND.n8595 GND.n1130 19.3944
R22219 GND.n8595 GND.n1126 19.3944
R22220 GND.n8601 GND.n1126 19.3944
R22221 GND.n8601 GND.n1124 19.3944
R22222 GND.n8605 GND.n1124 19.3944
R22223 GND.n8605 GND.n1120 19.3944
R22224 GND.n8611 GND.n1120 19.3944
R22225 GND.n8611 GND.n1118 19.3944
R22226 GND.n8615 GND.n1118 19.3944
R22227 GND.n8615 GND.n1114 19.3944
R22228 GND.n8621 GND.n1114 19.3944
R22229 GND.n8621 GND.n1112 19.3944
R22230 GND.n8625 GND.n1112 19.3944
R22231 GND.n8625 GND.n1108 19.3944
R22232 GND.n8631 GND.n1108 19.3944
R22233 GND.n8631 GND.n1106 19.3944
R22234 GND.n8635 GND.n1106 19.3944
R22235 GND.n8635 GND.n1102 19.3944
R22236 GND.n8641 GND.n1102 19.3944
R22237 GND.n8641 GND.n1100 19.3944
R22238 GND.n8645 GND.n1100 19.3944
R22239 GND.n8645 GND.n1096 19.3944
R22240 GND.n8651 GND.n1096 19.3944
R22241 GND.n8651 GND.n1094 19.3944
R22242 GND.n8655 GND.n1094 19.3944
R22243 GND.n8655 GND.n1090 19.3944
R22244 GND.n8661 GND.n1090 19.3944
R22245 GND.n8661 GND.n1088 19.3944
R22246 GND.n8665 GND.n1088 19.3944
R22247 GND.n8665 GND.n1084 19.3944
R22248 GND.n8671 GND.n1084 19.3944
R22249 GND.n8671 GND.n1082 19.3944
R22250 GND.n8675 GND.n1082 19.3944
R22251 GND.n8675 GND.n1078 19.3944
R22252 GND.n8681 GND.n1078 19.3944
R22253 GND.n8681 GND.n1076 19.3944
R22254 GND.n8685 GND.n1076 19.3944
R22255 GND.n8685 GND.n1072 19.3944
R22256 GND.n8691 GND.n1072 19.3944
R22257 GND.n8691 GND.n1070 19.3944
R22258 GND.n8695 GND.n1070 19.3944
R22259 GND.n8695 GND.n1066 19.3944
R22260 GND.n8701 GND.n1066 19.3944
R22261 GND.n8701 GND.n1064 19.3944
R22262 GND.n8705 GND.n1064 19.3944
R22263 GND.n8705 GND.n1060 19.3944
R22264 GND.n8711 GND.n1060 19.3944
R22265 GND.n8711 GND.n1058 19.3944
R22266 GND.n8715 GND.n1058 19.3944
R22267 GND.n8715 GND.n1054 19.3944
R22268 GND.n8721 GND.n1054 19.3944
R22269 GND.n8721 GND.n1052 19.3944
R22270 GND.n8725 GND.n1052 19.3944
R22271 GND.n8725 GND.n1048 19.3944
R22272 GND.n8731 GND.n1048 19.3944
R22273 GND.n8731 GND.n1046 19.3944
R22274 GND.n8735 GND.n1046 19.3944
R22275 GND.n8735 GND.n1042 19.3944
R22276 GND.n8741 GND.n1042 19.3944
R22277 GND.n8741 GND.n1040 19.3944
R22278 GND.n8745 GND.n1040 19.3944
R22279 GND.n8745 GND.n1036 19.3944
R22280 GND.n8751 GND.n1036 19.3944
R22281 GND.n8751 GND.n1034 19.3944
R22282 GND.n8755 GND.n1034 19.3944
R22283 GND.n8755 GND.n1030 19.3944
R22284 GND.n8761 GND.n1030 19.3944
R22285 GND.n8761 GND.n1028 19.3944
R22286 GND.n8765 GND.n1028 19.3944
R22287 GND.n8765 GND.n1024 19.3944
R22288 GND.n8771 GND.n1024 19.3944
R22289 GND.n8771 GND.n1022 19.3944
R22290 GND.n8775 GND.n1022 19.3944
R22291 GND.n8775 GND.n1018 19.3944
R22292 GND.n8781 GND.n1018 19.3944
R22293 GND.n8781 GND.n1016 19.3944
R22294 GND.n8785 GND.n1016 19.3944
R22295 GND.n8785 GND.n1012 19.3944
R22296 GND.n8791 GND.n1012 19.3944
R22297 GND.n8791 GND.n1010 19.3944
R22298 GND.n8795 GND.n1010 19.3944
R22299 GND.n8795 GND.n1006 19.3944
R22300 GND.n8801 GND.n1006 19.3944
R22301 GND.n8801 GND.n1004 19.3944
R22302 GND.n8805 GND.n1004 19.3944
R22303 GND.n8805 GND.n1000 19.3944
R22304 GND.n8811 GND.n1000 19.3944
R22305 GND.n8811 GND.n998 19.3944
R22306 GND.n8815 GND.n998 19.3944
R22307 GND.n8815 GND.n994 19.3944
R22308 GND.n8821 GND.n994 19.3944
R22309 GND.n8821 GND.n992 19.3944
R22310 GND.n8825 GND.n992 19.3944
R22311 GND.n8825 GND.n988 19.3944
R22312 GND.n8831 GND.n988 19.3944
R22313 GND.n8831 GND.n986 19.3944
R22314 GND.n8835 GND.n986 19.3944
R22315 GND.n8835 GND.n982 19.3944
R22316 GND.n8841 GND.n982 19.3944
R22317 GND.n8841 GND.n980 19.3944
R22318 GND.n8845 GND.n980 19.3944
R22319 GND.n8845 GND.n976 19.3944
R22320 GND.n8851 GND.n976 19.3944
R22321 GND.n8851 GND.n974 19.3944
R22322 GND.n8855 GND.n974 19.3944
R22323 GND.n8855 GND.n970 19.3944
R22324 GND.n8861 GND.n970 19.3944
R22325 GND.n8861 GND.n968 19.3944
R22326 GND.n8865 GND.n968 19.3944
R22327 GND.n8865 GND.n964 19.3944
R22328 GND.n8871 GND.n964 19.3944
R22329 GND.n8871 GND.n962 19.3944
R22330 GND.n8875 GND.n962 19.3944
R22331 GND.n8875 GND.n958 19.3944
R22332 GND.n8881 GND.n958 19.3944
R22333 GND.n8881 GND.n956 19.3944
R22334 GND.n8885 GND.n956 19.3944
R22335 GND.n8885 GND.n952 19.3944
R22336 GND.n8891 GND.n952 19.3944
R22337 GND.n8891 GND.n950 19.3944
R22338 GND.n8895 GND.n950 19.3944
R22339 GND.n8895 GND.n946 19.3944
R22340 GND.n8901 GND.n946 19.3944
R22341 GND.n8901 GND.n944 19.3944
R22342 GND.n8905 GND.n944 19.3944
R22343 GND.n8905 GND.n940 19.3944
R22344 GND.n8911 GND.n940 19.3944
R22345 GND.n8911 GND.n938 19.3944
R22346 GND.n8915 GND.n938 19.3944
R22347 GND.n8915 GND.n934 19.3944
R22348 GND.n8921 GND.n934 19.3944
R22349 GND.n8921 GND.n932 19.3944
R22350 GND.n8925 GND.n932 19.3944
R22351 GND.n8925 GND.n928 19.3944
R22352 GND.n8931 GND.n928 19.3944
R22353 GND.n8931 GND.n926 19.3944
R22354 GND.n8935 GND.n926 19.3944
R22355 GND.n8935 GND.n922 19.3944
R22356 GND.n8941 GND.n922 19.3944
R22357 GND.n8941 GND.n920 19.3944
R22358 GND.n8945 GND.n920 19.3944
R22359 GND.n8945 GND.n916 19.3944
R22360 GND.n8951 GND.n916 19.3944
R22361 GND.n8951 GND.n914 19.3944
R22362 GND.n8955 GND.n914 19.3944
R22363 GND.n8955 GND.n910 19.3944
R22364 GND.n8961 GND.n910 19.3944
R22365 GND.n8961 GND.n908 19.3944
R22366 GND.n8965 GND.n908 19.3944
R22367 GND.n8965 GND.n904 19.3944
R22368 GND.n8971 GND.n904 19.3944
R22369 GND.n8971 GND.n902 19.3944
R22370 GND.n8975 GND.n902 19.3944
R22371 GND.n8975 GND.n898 19.3944
R22372 GND.n8981 GND.n898 19.3944
R22373 GND.n8981 GND.n896 19.3944
R22374 GND.n8985 GND.n896 19.3944
R22375 GND.n8985 GND.n892 19.3944
R22376 GND.n8991 GND.n892 19.3944
R22377 GND.n8991 GND.n890 19.3944
R22378 GND.n8995 GND.n890 19.3944
R22379 GND.n8995 GND.n886 19.3944
R22380 GND.n9001 GND.n886 19.3944
R22381 GND.n9001 GND.n884 19.3944
R22382 GND.n9005 GND.n884 19.3944
R22383 GND.n9005 GND.n880 19.3944
R22384 GND.n9011 GND.n880 19.3944
R22385 GND.n9011 GND.n878 19.3944
R22386 GND.n9015 GND.n878 19.3944
R22387 GND.n9015 GND.n874 19.3944
R22388 GND.n9021 GND.n874 19.3944
R22389 GND.n9021 GND.n872 19.3944
R22390 GND.n9025 GND.n872 19.3944
R22391 GND.n9025 GND.n868 19.3944
R22392 GND.n9031 GND.n868 19.3944
R22393 GND.n9031 GND.n866 19.3944
R22394 GND.n9035 GND.n866 19.3944
R22395 GND.n9035 GND.n862 19.3944
R22396 GND.n9041 GND.n862 19.3944
R22397 GND.n9041 GND.n860 19.3944
R22398 GND.n9045 GND.n860 19.3944
R22399 GND.n9045 GND.n856 19.3944
R22400 GND.n9051 GND.n856 19.3944
R22401 GND.n9051 GND.n854 19.3944
R22402 GND.n9055 GND.n854 19.3944
R22403 GND.n9055 GND.n850 19.3944
R22404 GND.n9061 GND.n850 19.3944
R22405 GND.n9061 GND.n848 19.3944
R22406 GND.n9065 GND.n848 19.3944
R22407 GND.n9065 GND.n844 19.3944
R22408 GND.n9071 GND.n844 19.3944
R22409 GND.n9071 GND.n842 19.3944
R22410 GND.n9075 GND.n842 19.3944
R22411 GND.n9075 GND.n838 19.3944
R22412 GND.n9081 GND.n838 19.3944
R22413 GND.n9081 GND.n836 19.3944
R22414 GND.n9085 GND.n836 19.3944
R22415 GND.n9085 GND.n832 19.3944
R22416 GND.n9091 GND.n832 19.3944
R22417 GND.n9091 GND.n830 19.3944
R22418 GND.n9095 GND.n830 19.3944
R22419 GND.n9095 GND.n826 19.3944
R22420 GND.n9101 GND.n826 19.3944
R22421 GND.n9101 GND.n824 19.3944
R22422 GND.n9105 GND.n824 19.3944
R22423 GND.n9105 GND.n820 19.3944
R22424 GND.n9111 GND.n820 19.3944
R22425 GND.n9111 GND.n818 19.3944
R22426 GND.n9115 GND.n818 19.3944
R22427 GND.n9115 GND.n814 19.3944
R22428 GND.n9121 GND.n814 19.3944
R22429 GND.n9121 GND.n812 19.3944
R22430 GND.n9125 GND.n812 19.3944
R22431 GND.n9125 GND.n808 19.3944
R22432 GND.n9131 GND.n808 19.3944
R22433 GND.n9131 GND.n806 19.3944
R22434 GND.n9135 GND.n806 19.3944
R22435 GND.n9135 GND.n802 19.3944
R22436 GND.n9141 GND.n802 19.3944
R22437 GND.n9141 GND.n800 19.3944
R22438 GND.n9145 GND.n800 19.3944
R22439 GND.n9145 GND.n796 19.3944
R22440 GND.n9151 GND.n796 19.3944
R22441 GND.n9151 GND.n794 19.3944
R22442 GND.n9155 GND.n794 19.3944
R22443 GND.n9155 GND.n790 19.3944
R22444 GND.n9161 GND.n790 19.3944
R22445 GND.n9161 GND.n788 19.3944
R22446 GND.n9165 GND.n788 19.3944
R22447 GND.n9165 GND.n784 19.3944
R22448 GND.n9171 GND.n784 19.3944
R22449 GND.n9171 GND.n782 19.3944
R22450 GND.n9175 GND.n782 19.3944
R22451 GND.n9175 GND.n778 19.3944
R22452 GND.n9181 GND.n778 19.3944
R22453 GND.n9181 GND.n776 19.3944
R22454 GND.n9185 GND.n776 19.3944
R22455 GND.n9185 GND.n772 19.3944
R22456 GND.n9191 GND.n772 19.3944
R22457 GND.n9191 GND.n770 19.3944
R22458 GND.n9195 GND.n770 19.3944
R22459 GND.n9195 GND.n766 19.3944
R22460 GND.n9201 GND.n766 19.3944
R22461 GND.n9201 GND.n764 19.3944
R22462 GND.n9205 GND.n764 19.3944
R22463 GND.n9205 GND.n760 19.3944
R22464 GND.n9211 GND.n760 19.3944
R22465 GND.n9211 GND.n758 19.3944
R22466 GND.n9215 GND.n758 19.3944
R22467 GND.n9215 GND.n754 19.3944
R22468 GND.n9221 GND.n754 19.3944
R22469 GND.n9221 GND.n752 19.3944
R22470 GND.n9225 GND.n752 19.3944
R22471 GND.n9225 GND.n748 19.3944
R22472 GND.n9231 GND.n748 19.3944
R22473 GND.n9231 GND.n746 19.3944
R22474 GND.n9235 GND.n746 19.3944
R22475 GND.n9235 GND.n742 19.3944
R22476 GND.n9241 GND.n742 19.3944
R22477 GND.n9241 GND.n740 19.3944
R22478 GND.n9245 GND.n740 19.3944
R22479 GND.n9245 GND.n736 19.3944
R22480 GND.n9251 GND.n736 19.3944
R22481 GND.n9251 GND.n734 19.3944
R22482 GND.n9255 GND.n734 19.3944
R22483 GND.n9255 GND.n730 19.3944
R22484 GND.n9261 GND.n730 19.3944
R22485 GND.n9261 GND.n728 19.3944
R22486 GND.n9265 GND.n728 19.3944
R22487 GND.n9265 GND.n724 19.3944
R22488 GND.n9271 GND.n724 19.3944
R22489 GND.n9271 GND.n722 19.3944
R22490 GND.n9275 GND.n722 19.3944
R22491 GND.n9275 GND.n718 19.3944
R22492 GND.n9281 GND.n718 19.3944
R22493 GND.n9281 GND.n716 19.3944
R22494 GND.n9285 GND.n716 19.3944
R22495 GND.n9285 GND.n712 19.3944
R22496 GND.n9291 GND.n712 19.3944
R22497 GND.n9291 GND.n710 19.3944
R22498 GND.n9295 GND.n710 19.3944
R22499 GND.n9295 GND.n706 19.3944
R22500 GND.n9301 GND.n706 19.3944
R22501 GND.n9301 GND.n704 19.3944
R22502 GND.n9305 GND.n704 19.3944
R22503 GND.n9305 GND.n700 19.3944
R22504 GND.n9311 GND.n700 19.3944
R22505 GND.n9311 GND.n698 19.3944
R22506 GND.n9315 GND.n698 19.3944
R22507 GND.n9315 GND.n694 19.3944
R22508 GND.n9321 GND.n694 19.3944
R22509 GND.n9321 GND.n692 19.3944
R22510 GND.n9325 GND.n692 19.3944
R22511 GND.n9325 GND.n688 19.3944
R22512 GND.n9331 GND.n688 19.3944
R22513 GND.n9331 GND.n686 19.3944
R22514 GND.n9335 GND.n686 19.3944
R22515 GND.n9335 GND.n682 19.3944
R22516 GND.n9341 GND.n682 19.3944
R22517 GND.n9341 GND.n680 19.3944
R22518 GND.n9345 GND.n680 19.3944
R22519 GND.n9345 GND.n676 19.3944
R22520 GND.n9351 GND.n676 19.3944
R22521 GND.n9351 GND.n674 19.3944
R22522 GND.n9355 GND.n674 19.3944
R22523 GND.n9355 GND.n670 19.3944
R22524 GND.n9361 GND.n670 19.3944
R22525 GND.n9361 GND.n668 19.3944
R22526 GND.n9365 GND.n668 19.3944
R22527 GND.n9365 GND.n664 19.3944
R22528 GND.n9371 GND.n664 19.3944
R22529 GND.n9371 GND.n662 19.3944
R22530 GND.n9375 GND.n662 19.3944
R22531 GND.n9375 GND.n658 19.3944
R22532 GND.n9381 GND.n658 19.3944
R22533 GND.n9381 GND.n656 19.3944
R22534 GND.n9385 GND.n656 19.3944
R22535 GND.n9385 GND.n652 19.3944
R22536 GND.n9391 GND.n652 19.3944
R22537 GND.n9391 GND.n650 19.3944
R22538 GND.n9395 GND.n650 19.3944
R22539 GND.n9395 GND.n646 19.3944
R22540 GND.n9401 GND.n646 19.3944
R22541 GND.n9401 GND.n644 19.3944
R22542 GND.n9405 GND.n644 19.3944
R22543 GND.n9405 GND.n640 19.3944
R22544 GND.n9411 GND.n640 19.3944
R22545 GND.n9411 GND.n638 19.3944
R22546 GND.n9415 GND.n638 19.3944
R22547 GND.n9415 GND.n634 19.3944
R22548 GND.n9421 GND.n634 19.3944
R22549 GND.n9421 GND.n632 19.3944
R22550 GND.n9425 GND.n632 19.3944
R22551 GND.n9425 GND.n628 19.3944
R22552 GND.n9431 GND.n628 19.3944
R22553 GND.n9431 GND.n626 19.3944
R22554 GND.n9435 GND.n626 19.3944
R22555 GND.n9435 GND.n622 19.3944
R22556 GND.n9441 GND.n622 19.3944
R22557 GND.n9441 GND.n620 19.3944
R22558 GND.n9445 GND.n620 19.3944
R22559 GND.n9445 GND.n616 19.3944
R22560 GND.n9451 GND.n616 19.3944
R22561 GND.n9451 GND.n614 19.3944
R22562 GND.n9455 GND.n614 19.3944
R22563 GND.n9455 GND.n610 19.3944
R22564 GND.n9461 GND.n610 19.3944
R22565 GND.n9461 GND.n608 19.3944
R22566 GND.n9465 GND.n608 19.3944
R22567 GND.n9465 GND.n604 19.3944
R22568 GND.n9471 GND.n604 19.3944
R22569 GND.n9471 GND.n602 19.3944
R22570 GND.n9475 GND.n602 19.3944
R22571 GND.n9475 GND.n598 19.3944
R22572 GND.n9481 GND.n598 19.3944
R22573 GND.n9481 GND.n596 19.3944
R22574 GND.n9485 GND.n596 19.3944
R22575 GND.n9485 GND.n592 19.3944
R22576 GND.n9491 GND.n592 19.3944
R22577 GND.n9491 GND.n590 19.3944
R22578 GND.n9495 GND.n590 19.3944
R22579 GND.n9495 GND.n586 19.3944
R22580 GND.n9501 GND.n586 19.3944
R22581 GND.n9501 GND.n584 19.3944
R22582 GND.n9505 GND.n584 19.3944
R22583 GND.n9505 GND.n580 19.3944
R22584 GND.n9511 GND.n580 19.3944
R22585 GND.n9511 GND.n578 19.3944
R22586 GND.n9516 GND.n578 19.3944
R22587 GND.n9516 GND.n574 19.3944
R22588 GND.n9522 GND.n574 19.3944
R22589 GND.n9523 GND.n9522 19.3944
R22590 GND.n7180 GND.n7179 19.3944
R22591 GND.n7179 GND.n7178 19.3944
R22592 GND.n7178 GND.n7177 19.3944
R22593 GND.n7177 GND.n7175 19.3944
R22594 GND.n7175 GND.n7172 19.3944
R22595 GND.n7172 GND.n7171 19.3944
R22596 GND.n7171 GND.n7168 19.3944
R22597 GND.n7168 GND.n7167 19.3944
R22598 GND.n7167 GND.n7164 19.3944
R22599 GND.n7162 GND.n7160 19.3944
R22600 GND.n7160 GND.n7157 19.3944
R22601 GND.n7157 GND.n7156 19.3944
R22602 GND.n7156 GND.n7153 19.3944
R22603 GND.n7153 GND.n7152 19.3944
R22604 GND.n7152 GND.n7149 19.3944
R22605 GND.n7149 GND.n7148 19.3944
R22606 GND.n7148 GND.n7145 19.3944
R22607 GND.n7145 GND.n7144 19.3944
R22608 GND.n7144 GND.n7141 19.3944
R22609 GND.n7141 GND.n7140 19.3944
R22610 GND.n7137 GND.n7136 19.3944
R22611 GND.n7136 GND.n7133 19.3944
R22612 GND.n7133 GND.n7132 19.3944
R22613 GND.n7132 GND.n4833 19.3944
R22614 GND.n7186 GND.n4837 19.3944
R22615 GND.n5384 GND.n4837 19.3944
R22616 GND.n5387 GND.n5384 19.3944
R22617 GND.n5387 GND.n5379 19.3944
R22618 GND.n5397 GND.n5394 19.3944
R22619 GND.n5397 GND.n5377 19.3944
R22620 GND.n5403 GND.n5377 19.3944
R22621 GND.n5404 GND.n5403 19.3944
R22622 GND.n5407 GND.n5404 19.3944
R22623 GND.n5407 GND.n5375 19.3944
R22624 GND.n5413 GND.n5375 19.3944
R22625 GND.n5414 GND.n5413 19.3944
R22626 GND.n5417 GND.n5414 19.3944
R22627 GND.n5417 GND.n5373 19.3944
R22628 GND.n5423 GND.n5373 19.3944
R22629 GND.n5430 GND.n5427 19.3944
R22630 GND.n5430 GND.n5371 19.3944
R22631 GND.n5436 GND.n5371 19.3944
R22632 GND.n5437 GND.n5436 19.3944
R22633 GND.n5440 GND.n5437 19.3944
R22634 GND.n5440 GND.n5369 19.3944
R22635 GND.n5446 GND.n5369 19.3944
R22636 GND.n5447 GND.n5446 19.3944
R22637 GND.n5450 GND.n5447 19.3944
R22638 GND.n5450 GND.n5367 19.3944
R22639 GND.n5456 GND.n5367 19.3944
R22640 GND.n7087 GND.n4892 19.3944
R22641 GND.n7087 GND.n7086 19.3944
R22642 GND.n7086 GND.n4893 19.3944
R22643 GND.n5353 GND.n4893 19.3944
R22644 GND.n5353 GND.n5351 19.3944
R22645 GND.n6475 GND.n5351 19.3944
R22646 GND.n6476 GND.n6475 19.3944
R22647 GND.n6477 GND.n6476 19.3944
R22648 GND.n6477 GND.n5346 19.3944
R22649 GND.n6489 GND.n5346 19.3944
R22650 GND.n6490 GND.n6489 19.3944
R22651 GND.n6491 GND.n6490 19.3944
R22652 GND.n6491 GND.n5341 19.3944
R22653 GND.n6503 GND.n5341 19.3944
R22654 GND.n6504 GND.n6503 19.3944
R22655 GND.n6505 GND.n6504 19.3944
R22656 GND.n6505 GND.n5336 19.3944
R22657 GND.n6518 GND.n5336 19.3944
R22658 GND.n6519 GND.n6518 19.3944
R22659 GND.n6520 GND.n6519 19.3944
R22660 GND.n6521 GND.n6520 19.3944
R22661 GND.n6667 GND.n6521 19.3944
R22662 GND.n6667 GND.n6666 19.3944
R22663 GND.n6666 GND.n6665 19.3944
R22664 GND.n6665 GND.n6523 19.3944
R22665 GND.n6655 GND.n6523 19.3944
R22666 GND.n6655 GND.n6654 19.3944
R22667 GND.n6654 GND.n6653 19.3944
R22668 GND.n6653 GND.n6530 19.3944
R22669 GND.n6643 GND.n6530 19.3944
R22670 GND.n6643 GND.n6642 19.3944
R22671 GND.n6642 GND.n6641 19.3944
R22672 GND.n6641 GND.n6537 19.3944
R22673 GND.n6631 GND.n6537 19.3944
R22674 GND.n6631 GND.n6630 19.3944
R22675 GND.n6630 GND.n6629 19.3944
R22676 GND.n6629 GND.n6544 19.3944
R22677 GND.n6619 GND.n6544 19.3944
R22678 GND.n6619 GND.n6618 19.3944
R22679 GND.n6618 GND.n6617 19.3944
R22680 GND.n6617 GND.n6551 19.3944
R22681 GND.n6607 GND.n6551 19.3944
R22682 GND.n6607 GND.n6606 19.3944
R22683 GND.n6606 GND.n6605 19.3944
R22684 GND.n6605 GND.n6558 19.3944
R22685 GND.n6595 GND.n6558 19.3944
R22686 GND.n6595 GND.n6594 19.3944
R22687 GND.n6594 GND.n6593 19.3944
R22688 GND.n6593 GND.n6565 19.3944
R22689 GND.n6583 GND.n6565 19.3944
R22690 GND.n6583 GND.n6582 19.3944
R22691 GND.n6582 GND.n6581 19.3944
R22692 GND.n6581 GND.n6574 19.3944
R22693 GND.n6574 GND.n6573 19.3944
R22694 GND.n6573 GND.n5287 19.3944
R22695 GND.n6771 GND.n5287 19.3944
R22696 GND.n6772 GND.n6771 19.3944
R22697 GND.n6773 GND.n6772 19.3944
R22698 GND.n6776 GND.n6773 19.3944
R22699 GND.n6776 GND.n5282 19.3944
R22700 GND.n6784 GND.n5282 19.3944
R22701 GND.n6785 GND.n6784 19.3944
R22702 GND.n6785 GND.n5278 19.3944
R22703 GND.n6794 GND.n5278 19.3944
R22704 GND.n6795 GND.n6794 19.3944
R22705 GND.n6893 GND.n6795 19.3944
R22706 GND.n6893 GND.n6892 19.3944
R22707 GND.n6892 GND.n6891 19.3944
R22708 GND.n6891 GND.n6797 19.3944
R22709 GND.n6881 GND.n6797 19.3944
R22710 GND.n6881 GND.n6880 19.3944
R22711 GND.n6880 GND.n6879 19.3944
R22712 GND.n6879 GND.n6804 19.3944
R22713 GND.n6869 GND.n6804 19.3944
R22714 GND.n6869 GND.n6868 19.3944
R22715 GND.n6868 GND.n6867 19.3944
R22716 GND.n6867 GND.n6811 19.3944
R22717 GND.n6857 GND.n6811 19.3944
R22718 GND.n6857 GND.n6856 19.3944
R22719 GND.n6856 GND.n6855 19.3944
R22720 GND.n6855 GND.n6818 19.3944
R22721 GND.n6845 GND.n6818 19.3944
R22722 GND.n6845 GND.n6844 19.3944
R22723 GND.n6844 GND.n6843 19.3944
R22724 GND.n6843 GND.n6825 19.3944
R22725 GND.n6833 GND.n6825 19.3944
R22726 GND.n6833 GND.n6832 19.3944
R22727 GND.n6832 GND.n6831 19.3944
R22728 GND.n6831 GND.n437 19.3944
R22729 GND.n9737 GND.n437 19.3944
R22730 GND.n9738 GND.n9737 19.3944
R22731 GND.n9740 GND.n9738 19.3944
R22732 GND.n9740 GND.n433 19.3944
R22733 GND.n9752 GND.n433 19.3944
R22734 GND.n9753 GND.n9752 19.3944
R22735 GND.n9755 GND.n9753 19.3944
R22736 GND.n9755 GND.n429 19.3944
R22737 GND.n9767 GND.n429 19.3944
R22738 GND.n9768 GND.n9767 19.3944
R22739 GND.n9770 GND.n9768 19.3944
R22740 GND.n9770 GND.n425 19.3944
R22741 GND.n9782 GND.n425 19.3944
R22742 GND.n9783 GND.n9782 19.3944
R22743 GND.n9785 GND.n9783 19.3944
R22744 GND.n9785 GND.n421 19.3944
R22745 GND.n10106 GND.n421 19.3944
R22746 GND.n10107 GND.n10106 19.3944
R22747 GND.n10110 GND.n10107 19.3944
R22748 GND.n10111 GND.n10110 19.3944
R22749 GND.n10113 GND.n10111 19.3944
R22750 GND.n10114 GND.n10113 19.3944
R22751 GND.n10117 GND.n10114 19.3944
R22752 GND.n10118 GND.n10117 19.3944
R22753 GND.n10120 GND.n10118 19.3944
R22754 GND.n10121 GND.n10120 19.3944
R22755 GND.n10124 GND.n10121 19.3944
R22756 GND.n10125 GND.n10124 19.3944
R22757 GND.n10127 GND.n10125 19.3944
R22758 GND.n10128 GND.n10127 19.3944
R22759 GND.n10130 GND.n10128 19.3944
R22760 GND.n10131 GND.n10130 19.3944
R22761 GND.n7089 GND.n4888 19.3944
R22762 GND.n7089 GND.n4889 19.3944
R22763 GND.n5356 GND.n4889 19.3944
R22764 GND.n5359 GND.n5356 19.3944
R22765 GND.n5360 GND.n5359 19.3944
R22766 GND.n5360 GND.n4929 19.3944
R22767 GND.n7068 GND.n4929 19.3944
R22768 GND.n7068 GND.n7067 19.3944
R22769 GND.n7067 GND.n7066 19.3944
R22770 GND.n7066 GND.n4933 19.3944
R22771 GND.n7056 GND.n4933 19.3944
R22772 GND.n7056 GND.n7055 19.3944
R22773 GND.n7055 GND.n7054 19.3944
R22774 GND.n7054 GND.n4954 19.3944
R22775 GND.n7044 GND.n4954 19.3944
R22776 GND.n7044 GND.n7043 19.3944
R22777 GND.n7043 GND.n7042 19.3944
R22778 GND.n7042 GND.n4975 19.3944
R22779 GND.n7032 GND.n4975 19.3944
R22780 GND.n7032 GND.n7031 19.3944
R22781 GND.n7031 GND.n7030 19.3944
R22782 GND.n7030 GND.n4996 19.3944
R22783 GND.n7020 GND.n4996 19.3944
R22784 GND.n7020 GND.n7019 19.3944
R22785 GND.n7019 GND.n7018 19.3944
R22786 GND.n7018 GND.n5016 19.3944
R22787 GND.n7008 GND.n5016 19.3944
R22788 GND.n7008 GND.n7007 19.3944
R22789 GND.n7007 GND.n7006 19.3944
R22790 GND.n7006 GND.n5037 19.3944
R22791 GND.n6996 GND.n5037 19.3944
R22792 GND.n6996 GND.n6995 19.3944
R22793 GND.n6995 GND.n6994 19.3944
R22794 GND.n6994 GND.n5058 19.3944
R22795 GND.n6984 GND.n5058 19.3944
R22796 GND.n6984 GND.n6983 19.3944
R22797 GND.n6983 GND.n6982 19.3944
R22798 GND.n6982 GND.n5079 19.3944
R22799 GND.n6972 GND.n5079 19.3944
R22800 GND.n6972 GND.n6971 19.3944
R22801 GND.n6971 GND.n6970 19.3944
R22802 GND.n6970 GND.n5100 19.3944
R22803 GND.n6960 GND.n5100 19.3944
R22804 GND.n6960 GND.n6959 19.3944
R22805 GND.n6959 GND.n6958 19.3944
R22806 GND.n6958 GND.n5121 19.3944
R22807 GND.n6948 GND.n5121 19.3944
R22808 GND.n6948 GND.n6947 19.3944
R22809 GND.n6947 GND.n6946 19.3944
R22810 GND.n6946 GND.n5142 19.3944
R22811 GND.n6936 GND.n5142 19.3944
R22812 GND.n6936 GND.n6935 19.3944
R22813 GND.n6935 GND.n6934 19.3944
R22814 GND.n6934 GND.n5163 19.3944
R22815 GND.n6924 GND.n5163 19.3944
R22816 GND.n6924 GND.n6923 19.3944
R22817 GND.n6923 GND.n6922 19.3944
R22818 GND.n6922 GND.n5182 19.3944
R22819 GND.n5284 GND.n5182 19.3944
R22820 GND.n6781 GND.n5284 19.3944
R22821 GND.n6782 GND.n6781 19.3944
R22822 GND.n6782 GND.n5280 19.3944
R22823 GND.n6791 GND.n5280 19.3944
R22824 GND.n6791 GND.n133 19.3944
R22825 GND.n10301 GND.n133 19.3944
R22826 GND.n10301 GND.n10300 19.3944
R22827 GND.n10300 GND.n10299 19.3944
R22828 GND.n10299 GND.n137 19.3944
R22829 GND.n10289 GND.n137 19.3944
R22830 GND.n10289 GND.n10288 19.3944
R22831 GND.n10288 GND.n10287 19.3944
R22832 GND.n10287 GND.n157 19.3944
R22833 GND.n10277 GND.n157 19.3944
R22834 GND.n10277 GND.n10276 19.3944
R22835 GND.n10276 GND.n10275 19.3944
R22836 GND.n10275 GND.n178 19.3944
R22837 GND.n10265 GND.n178 19.3944
R22838 GND.n10265 GND.n10264 19.3944
R22839 GND.n10264 GND.n10263 19.3944
R22840 GND.n10263 GND.n199 19.3944
R22841 GND.n10253 GND.n199 19.3944
R22842 GND.n10253 GND.n10252 19.3944
R22843 GND.n10252 GND.n10251 19.3944
R22844 GND.n10251 GND.n220 19.3944
R22845 GND.n10241 GND.n220 19.3944
R22846 GND.n10241 GND.n10240 19.3944
R22847 GND.n10240 GND.n10239 19.3944
R22848 GND.n10239 GND.n241 19.3944
R22849 GND.n10229 GND.n241 19.3944
R22850 GND.n10229 GND.n10228 19.3944
R22851 GND.n10228 GND.n10227 19.3944
R22852 GND.n10227 GND.n261 19.3944
R22853 GND.n10217 GND.n261 19.3944
R22854 GND.n10217 GND.n10216 19.3944
R22855 GND.n10216 GND.n10215 19.3944
R22856 GND.n10215 GND.n282 19.3944
R22857 GND.n10205 GND.n282 19.3944
R22858 GND.n10205 GND.n10204 19.3944
R22859 GND.n10204 GND.n10203 19.3944
R22860 GND.n10203 GND.n303 19.3944
R22861 GND.n10193 GND.n303 19.3944
R22862 GND.n10193 GND.n10192 19.3944
R22863 GND.n10192 GND.n10191 19.3944
R22864 GND.n10191 GND.n324 19.3944
R22865 GND.n10181 GND.n324 19.3944
R22866 GND.n10181 GND.n10180 19.3944
R22867 GND.n10180 GND.n10179 19.3944
R22868 GND.n10179 GND.n345 19.3944
R22869 GND.n10169 GND.n345 19.3944
R22870 GND.n10169 GND.n10168 19.3944
R22871 GND.n10168 GND.n10167 19.3944
R22872 GND.n10167 GND.n366 19.3944
R22873 GND.n10157 GND.n366 19.3944
R22874 GND.n10157 GND.n10156 19.3944
R22875 GND.n10156 GND.n10155 19.3944
R22876 GND.n10155 GND.n385 19.3944
R22877 GND.n10145 GND.n385 19.3944
R22878 GND.n10145 GND.n10144 19.3944
R22879 GND.n10144 GND.n10143 19.3944
R22880 GND.n10143 GND.n404 19.3944
R22881 GND.n10133 GND.n404 19.3944
R22882 GND.n10008 GND.n9851 19.3944
R22883 GND.n10011 GND.n10008 19.3944
R22884 GND.n10014 GND.n10011 19.3944
R22885 GND.n10014 GND.n9849 19.3944
R22886 GND.n10018 GND.n9849 19.3944
R22887 GND.n10021 GND.n10018 19.3944
R22888 GND.n10024 GND.n10021 19.3944
R22889 GND.n10024 GND.n9847 19.3944
R22890 GND.n10028 GND.n9847 19.3944
R22891 GND.n10031 GND.n10028 19.3944
R22892 GND.n10033 GND.n10031 19.3944
R22893 GND.n9975 GND.n9857 19.3944
R22894 GND.n9978 GND.n9975 19.3944
R22895 GND.n9981 GND.n9978 19.3944
R22896 GND.n9981 GND.n9855 19.3944
R22897 GND.n9985 GND.n9855 19.3944
R22898 GND.n9988 GND.n9985 19.3944
R22899 GND.n9991 GND.n9988 19.3944
R22900 GND.n9991 GND.n9853 19.3944
R22901 GND.n9995 GND.n9853 19.3944
R22902 GND.n9998 GND.n9995 19.3944
R22903 GND.n10004 GND.n9998 19.3944
R22904 GND.n9943 GND.n9867 19.3944
R22905 GND.n9947 GND.n9867 19.3944
R22906 GND.n9950 GND.n9947 19.3944
R22907 GND.n9953 GND.n9950 19.3944
R22908 GND.n9953 GND.n9865 19.3944
R22909 GND.n9957 GND.n9865 19.3944
R22910 GND.n9960 GND.n9957 19.3944
R22911 GND.n9963 GND.n9960 19.3944
R22912 GND.n9963 GND.n9863 19.3944
R22913 GND.n9967 GND.n9863 19.3944
R22914 GND.n9970 GND.n9967 19.3944
R22915 GND.n9912 GND.n9875 19.3944
R22916 GND.n9916 GND.n9875 19.3944
R22917 GND.n9919 GND.n9916 19.3944
R22918 GND.n9922 GND.n9919 19.3944
R22919 GND.n9922 GND.n9873 19.3944
R22920 GND.n9926 GND.n9873 19.3944
R22921 GND.n9929 GND.n9926 19.3944
R22922 GND.n9932 GND.n9929 19.3944
R22923 GND.n9932 GND.n9871 19.3944
R22924 GND.n9936 GND.n9871 19.3944
R22925 GND.n9939 GND.n9936 19.3944
R22926 GND.n9887 GND.n9884 19.3944
R22927 GND.n9890 GND.n9887 19.3944
R22928 GND.n9893 GND.n9890 19.3944
R22929 GND.n9893 GND.n9882 19.3944
R22930 GND.n9897 GND.n9882 19.3944
R22931 GND.n9900 GND.n9897 19.3944
R22932 GND.n9903 GND.n9900 19.3944
R22933 GND.n9903 GND.n9880 19.3944
R22934 GND.n9908 GND.n9880 19.3944
R22935 GND.n10052 GND.n10049 19.3944
R22936 GND.n10055 GND.n10052 19.3944
R22937 GND.n10058 GND.n10055 19.3944
R22938 GND.n10058 GND.n10047 19.3944
R22939 GND.n10062 GND.n10047 19.3944
R22940 GND.n10065 GND.n10062 19.3944
R22941 GND.n10067 GND.n10065 19.3944
R22942 GND.n10067 GND.n10045 19.3944
R22943 GND.n10071 GND.n10045 19.3944
R22944 GND.n6418 GND.n5365 19.3944
R22945 GND.n6422 GND.n5365 19.3944
R22946 GND.n6423 GND.n6422 19.3944
R22947 GND.n6426 GND.n6423 19.3944
R22948 GND.n6426 GND.n5363 19.3944
R22949 GND.n6430 GND.n5363 19.3944
R22950 GND.n6430 GND.n5350 19.3944
R22951 GND.n6481 GND.n5350 19.3944
R22952 GND.n6481 GND.n5348 19.3944
R22953 GND.n6485 GND.n5348 19.3944
R22954 GND.n6485 GND.n5345 19.3944
R22955 GND.n6495 GND.n5345 19.3944
R22956 GND.n6495 GND.n5343 19.3944
R22957 GND.n6499 GND.n5343 19.3944
R22958 GND.n6499 GND.n5340 19.3944
R22959 GND.n6509 GND.n5340 19.3944
R22960 GND.n6509 GND.n5338 19.3944
R22961 GND.n6514 GND.n5338 19.3944
R22962 GND.n6514 GND.n5331 19.3944
R22963 GND.n6673 GND.n5331 19.3944
R22964 GND.n6673 GND.n6672 19.3944
R22965 GND.n6672 GND.n6671 19.3944
R22966 GND.n6671 GND.n5335 19.3944
R22967 GND.n6661 GND.n5335 19.3944
R22968 GND.n6661 GND.n6660 19.3944
R22969 GND.n6660 GND.n6659 19.3944
R22970 GND.n6659 GND.n6528 19.3944
R22971 GND.n6649 GND.n6528 19.3944
R22972 GND.n6649 GND.n6648 19.3944
R22973 GND.n6648 GND.n6647 19.3944
R22974 GND.n6647 GND.n6535 19.3944
R22975 GND.n6637 GND.n6535 19.3944
R22976 GND.n6637 GND.n6636 19.3944
R22977 GND.n6636 GND.n6635 19.3944
R22978 GND.n6635 GND.n6542 19.3944
R22979 GND.n6625 GND.n6542 19.3944
R22980 GND.n6625 GND.n6624 19.3944
R22981 GND.n6624 GND.n6623 19.3944
R22982 GND.n6623 GND.n6549 19.3944
R22983 GND.n6613 GND.n6549 19.3944
R22984 GND.n6613 GND.n6612 19.3944
R22985 GND.n6612 GND.n6611 19.3944
R22986 GND.n6611 GND.n6556 19.3944
R22987 GND.n6601 GND.n6556 19.3944
R22988 GND.n6601 GND.n6600 19.3944
R22989 GND.n6600 GND.n6599 19.3944
R22990 GND.n6599 GND.n6563 19.3944
R22991 GND.n6589 GND.n6563 19.3944
R22992 GND.n6589 GND.n6588 19.3944
R22993 GND.n6588 GND.n6587 19.3944
R22994 GND.n6587 GND.n6570 19.3944
R22995 GND.n6577 GND.n6570 19.3944
R22996 GND.n6577 GND.n5290 19.3944
R22997 GND.n6756 GND.n5290 19.3944
R22998 GND.n6756 GND.n5288 19.3944
R22999 GND.n6767 GND.n5288 19.3944
R23000 GND.n6767 GND.n6766 19.3944
R23001 GND.n6766 GND.n6765 19.3944
R23002 GND.n6765 GND.n6764 19.3944
R23003 GND.n6764 GND.n104 19.3944
R23004 GND.n10312 GND.n104 19.3944
R23005 GND.n10312 GND.n105 19.3944
R23006 GND.n5272 GND.n105 19.3944
R23007 GND.n6899 GND.n5272 19.3944
R23008 GND.n6899 GND.n6898 19.3944
R23009 GND.n6898 GND.n6897 19.3944
R23010 GND.n6897 GND.n5277 19.3944
R23011 GND.n6887 GND.n5277 19.3944
R23012 GND.n6887 GND.n6886 19.3944
R23013 GND.n6886 GND.n6885 19.3944
R23014 GND.n6885 GND.n6802 19.3944
R23015 GND.n6875 GND.n6802 19.3944
R23016 GND.n6875 GND.n6874 19.3944
R23017 GND.n6874 GND.n6873 19.3944
R23018 GND.n6873 GND.n6809 19.3944
R23019 GND.n6863 GND.n6809 19.3944
R23020 GND.n6863 GND.n6862 19.3944
R23021 GND.n6862 GND.n6861 19.3944
R23022 GND.n6861 GND.n6816 19.3944
R23023 GND.n6851 GND.n6816 19.3944
R23024 GND.n6851 GND.n6850 19.3944
R23025 GND.n6850 GND.n6849 19.3944
R23026 GND.n6849 GND.n6823 19.3944
R23027 GND.n6839 GND.n6823 19.3944
R23028 GND.n6839 GND.n6838 19.3944
R23029 GND.n6838 GND.n6837 19.3944
R23030 GND.n6837 GND.n440 19.3944
R23031 GND.n9729 GND.n440 19.3944
R23032 GND.n9729 GND.n438 19.3944
R23033 GND.n9733 GND.n438 19.3944
R23034 GND.n9733 GND.n436 19.3944
R23035 GND.n9744 GND.n436 19.3944
R23036 GND.n9744 GND.n434 19.3944
R23037 GND.n9748 GND.n434 19.3944
R23038 GND.n9748 GND.n432 19.3944
R23039 GND.n9759 GND.n432 19.3944
R23040 GND.n9759 GND.n430 19.3944
R23041 GND.n9763 GND.n430 19.3944
R23042 GND.n9763 GND.n428 19.3944
R23043 GND.n9774 GND.n428 19.3944
R23044 GND.n9774 GND.n426 19.3944
R23045 GND.n9778 GND.n426 19.3944
R23046 GND.n9778 GND.n424 19.3944
R23047 GND.n9789 GND.n424 19.3944
R23048 GND.n9789 GND.n422 19.3944
R23049 GND.n10102 GND.n422 19.3944
R23050 GND.n10102 GND.n10101 19.3944
R23051 GND.n10101 GND.n10100 19.3944
R23052 GND.n10100 GND.n10098 19.3944
R23053 GND.n10098 GND.n10097 19.3944
R23054 GND.n10097 GND.n10095 19.3944
R23055 GND.n10095 GND.n10094 19.3944
R23056 GND.n10094 GND.n10092 19.3944
R23057 GND.n10092 GND.n10091 19.3944
R23058 GND.n10091 GND.n10089 19.3944
R23059 GND.n10089 GND.n10088 19.3944
R23060 GND.n10088 GND.n10086 19.3944
R23061 GND.n10086 GND.n10085 19.3944
R23062 GND.n10085 GND.n10083 19.3944
R23063 GND.n10083 GND.n10082 19.3944
R23064 GND.n10082 GND.n10080 19.3944
R23065 GND.n7699 GND.n3883 19.3944
R23066 GND.n7689 GND.n3883 19.3944
R23067 GND.n7689 GND.n7688 19.3944
R23068 GND.n7688 GND.n7687 19.3944
R23069 GND.n7687 GND.n3901 19.3944
R23070 GND.n7678 GND.n3901 19.3944
R23071 GND.n7678 GND.n7677 19.3944
R23072 GND.n7677 GND.n7676 19.3944
R23073 GND.n7676 GND.n3921 19.3944
R23074 GND.n3971 GND.n3921 19.3944
R23075 GND.n3975 GND.n3971 19.3944
R23076 GND.n3978 GND.n3975 19.3944
R23077 GND.n3979 GND.n3978 19.3944
R23078 GND.n3979 GND.n3969 19.3944
R23079 GND.n7647 GND.n3969 19.3944
R23080 GND.n7647 GND.n7646 19.3944
R23081 GND.n7646 GND.n7645 19.3944
R23082 GND.n7645 GND.n3985 19.3944
R23083 GND.n7635 GND.n3985 19.3944
R23084 GND.n7635 GND.n7634 19.3944
R23085 GND.n7634 GND.n7633 19.3944
R23086 GND.n7633 GND.n4005 19.3944
R23087 GND.n7623 GND.n4005 19.3944
R23088 GND.n7623 GND.n7622 19.3944
R23089 GND.n7622 GND.n7621 19.3944
R23090 GND.n7621 GND.n4025 19.3944
R23091 GND.n4076 GND.n4025 19.3944
R23092 GND.n4080 GND.n4076 19.3944
R23093 GND.n4083 GND.n4080 19.3944
R23094 GND.n4084 GND.n4083 19.3944
R23095 GND.n4084 GND.n4074 19.3944
R23096 GND.n7592 GND.n4074 19.3944
R23097 GND.n7592 GND.n7591 19.3944
R23098 GND.n7591 GND.n7590 19.3944
R23099 GND.n7590 GND.n4090 19.3944
R23100 GND.n7580 GND.n4090 19.3944
R23101 GND.n7580 GND.n7579 19.3944
R23102 GND.n7579 GND.n7578 19.3944
R23103 GND.n7578 GND.n4110 19.3944
R23104 GND.n7568 GND.n4110 19.3944
R23105 GND.n7568 GND.n7567 19.3944
R23106 GND.n7567 GND.n7566 19.3944
R23107 GND.n7566 GND.n4130 19.3944
R23108 GND.n4181 GND.n4130 19.3944
R23109 GND.n4185 GND.n4181 19.3944
R23110 GND.n4188 GND.n4185 19.3944
R23111 GND.n4189 GND.n4188 19.3944
R23112 GND.n4189 GND.n4179 19.3944
R23113 GND.n7537 GND.n4179 19.3944
R23114 GND.n7537 GND.n7536 19.3944
R23115 GND.n7536 GND.n7535 19.3944
R23116 GND.n7535 GND.n4195 19.3944
R23117 GND.n7525 GND.n4195 19.3944
R23118 GND.n7525 GND.n7524 19.3944
R23119 GND.n7524 GND.n7523 19.3944
R23120 GND.n7523 GND.n4214 19.3944
R23121 GND.n7513 GND.n4214 19.3944
R23122 GND.n7513 GND.n7512 19.3944
R23123 GND.n7512 GND.n7511 19.3944
R23124 GND.n7511 GND.n4233 19.3944
R23125 GND.n4283 GND.n4233 19.3944
R23126 GND.n4287 GND.n4283 19.3944
R23127 GND.n4290 GND.n4287 19.3944
R23128 GND.n4291 GND.n4290 19.3944
R23129 GND.n4291 GND.n4281 19.3944
R23130 GND.n7482 GND.n4281 19.3944
R23131 GND.n7482 GND.n7481 19.3944
R23132 GND.n7481 GND.n7480 19.3944
R23133 GND.n7480 GND.n4297 19.3944
R23134 GND.n7470 GND.n4297 19.3944
R23135 GND.n7470 GND.n7469 19.3944
R23136 GND.n7469 GND.n7468 19.3944
R23137 GND.n7468 GND.n4317 19.3944
R23138 GND.n7458 GND.n4317 19.3944
R23139 GND.n7458 GND.n7457 19.3944
R23140 GND.n7457 GND.n7456 19.3944
R23141 GND.n7456 GND.n4337 19.3944
R23142 GND.n4388 GND.n4337 19.3944
R23143 GND.n4392 GND.n4388 19.3944
R23144 GND.n4395 GND.n4392 19.3944
R23145 GND.n4396 GND.n4395 19.3944
R23146 GND.n4396 GND.n4386 19.3944
R23147 GND.n7427 GND.n4386 19.3944
R23148 GND.n7427 GND.n7426 19.3944
R23149 GND.n7426 GND.n7425 19.3944
R23150 GND.n7425 GND.n4402 19.3944
R23151 GND.n7415 GND.n4402 19.3944
R23152 GND.n7415 GND.n7414 19.3944
R23153 GND.n5683 GND.n5669 19.3944
R23154 GND.n5683 GND.n5670 19.3944
R23155 GND.n5679 GND.n5670 19.3944
R23156 GND.n5679 GND.n5677 19.3944
R23157 GND.n5677 GND.n5676 19.3944
R23158 GND.n5676 GND.n5653 19.3944
R23159 GND.n5761 GND.n5653 19.3944
R23160 GND.n5762 GND.n5761 19.3944
R23161 GND.n5762 GND.n5651 19.3944
R23162 GND.n5766 GND.n5651 19.3944
R23163 GND.n5767 GND.n5766 19.3944
R23164 GND.n5770 GND.n5767 19.3944
R23165 GND.n5770 GND.n5647 19.3944
R23166 GND.n5795 GND.n5647 19.3944
R23167 GND.n5795 GND.n5794 19.3944
R23168 GND.n5794 GND.n5793 19.3944
R23169 GND.n5793 GND.n5791 19.3944
R23170 GND.n5791 GND.n5790 19.3944
R23171 GND.n5790 GND.n5788 19.3944
R23172 GND.n5788 GND.n5787 19.3944
R23173 GND.n5787 GND.n5785 19.3944
R23174 GND.n5785 GND.n5784 19.3944
R23175 GND.n5784 GND.n5622 19.3944
R23176 GND.n5865 GND.n5622 19.3944
R23177 GND.n5866 GND.n5865 19.3944
R23178 GND.n5866 GND.n5620 19.3944
R23179 GND.n5870 GND.n5620 19.3944
R23180 GND.n5871 GND.n5870 19.3944
R23181 GND.n5874 GND.n5871 19.3944
R23182 GND.n5874 GND.n5616 19.3944
R23183 GND.n5899 GND.n5616 19.3944
R23184 GND.n5899 GND.n5898 19.3944
R23185 GND.n5898 GND.n5897 19.3944
R23186 GND.n5897 GND.n5895 19.3944
R23187 GND.n5895 GND.n5894 19.3944
R23188 GND.n5894 GND.n5892 19.3944
R23189 GND.n5892 GND.n5891 19.3944
R23190 GND.n5891 GND.n5889 19.3944
R23191 GND.n5889 GND.n5888 19.3944
R23192 GND.n5888 GND.n5591 19.3944
R23193 GND.n5968 GND.n5591 19.3944
R23194 GND.n5969 GND.n5968 19.3944
R23195 GND.n5969 GND.n5589 19.3944
R23196 GND.n5973 GND.n5589 19.3944
R23197 GND.n5974 GND.n5973 19.3944
R23198 GND.n5977 GND.n5974 19.3944
R23199 GND.n5977 GND.n5585 19.3944
R23200 GND.n6002 GND.n5585 19.3944
R23201 GND.n6002 GND.n6001 19.3944
R23202 GND.n6001 GND.n6000 19.3944
R23203 GND.n6000 GND.n5998 19.3944
R23204 GND.n5998 GND.n5997 19.3944
R23205 GND.n5997 GND.n5995 19.3944
R23206 GND.n5995 GND.n5994 19.3944
R23207 GND.n5994 GND.n5992 19.3944
R23208 GND.n5992 GND.n5991 19.3944
R23209 GND.n5991 GND.n5558 19.3944
R23210 GND.n6071 GND.n5558 19.3944
R23211 GND.n6072 GND.n6071 19.3944
R23212 GND.n6072 GND.n5556 19.3944
R23213 GND.n6076 GND.n5556 19.3944
R23214 GND.n6077 GND.n6076 19.3944
R23215 GND.n6080 GND.n6077 19.3944
R23216 GND.n6080 GND.n5552 19.3944
R23217 GND.n6105 GND.n5552 19.3944
R23218 GND.n6105 GND.n6104 19.3944
R23219 GND.n6104 GND.n6103 19.3944
R23220 GND.n6103 GND.n6101 19.3944
R23221 GND.n6101 GND.n6100 19.3944
R23222 GND.n6100 GND.n6098 19.3944
R23223 GND.n6098 GND.n6097 19.3944
R23224 GND.n6097 GND.n6095 19.3944
R23225 GND.n6095 GND.n6094 19.3944
R23226 GND.n6094 GND.n5526 19.3944
R23227 GND.n6174 GND.n5526 19.3944
R23228 GND.n6175 GND.n6174 19.3944
R23229 GND.n6175 GND.n5524 19.3944
R23230 GND.n6179 GND.n5524 19.3944
R23231 GND.n6180 GND.n6179 19.3944
R23232 GND.n6183 GND.n6180 19.3944
R23233 GND.n6183 GND.n5520 19.3944
R23234 GND.n6201 GND.n5520 19.3944
R23235 GND.n6201 GND.n6200 19.3944
R23236 GND.n6200 GND.n6199 19.3944
R23237 GND.n6199 GND.n6197 19.3944
R23238 GND.n6197 GND.n6196 19.3944
R23239 GND.n6196 GND.n6193 19.3944
R23240 GND.n6193 GND.n5496 19.3944
R23241 GND.n7756 GND.n7755 19.3944
R23242 GND.n7755 GND.n7754 19.3944
R23243 GND.n7754 GND.n7753 19.3944
R23244 GND.n7753 GND.n7751 19.3944
R23245 GND.n7751 GND.n7748 19.3944
R23246 GND.n7748 GND.n7747 19.3944
R23247 GND.n7747 GND.n7744 19.3944
R23248 GND.n7744 GND.n7743 19.3944
R23249 GND.n7743 GND.n7740 19.3944
R23250 GND.n7740 GND.n7739 19.3944
R23251 GND.n7739 GND.n2357 19.3944
R23252 GND.n7736 GND.n7735 19.3944
R23253 GND.n7731 GND.n7730 19.3944
R23254 GND.n7726 GND.n7725 19.3944
R23255 GND.n7721 GND.n7720 19.3944
R23256 GND.n7716 GND.n7715 19.3944
R23257 GND.n7711 GND.n7710 19.3944
R23258 GND.n7707 GND.n7704 19.3944
R23259 GND.n7704 GND.n7703 19.3944
R23260 GND.n7703 GND.n3881 19.3944
R23261 GND.n6349 GND.n6348 19.3944
R23262 GND.n6348 GND.n4420 19.3944
R23263 GND.n7411 GND.n4420 19.3944
R23264 GND.n6316 GND.n6315 19.3944
R23265 GND.n6319 GND.n6316 19.3944
R23266 GND.n6319 GND.n5493 19.3944
R23267 GND.n6325 GND.n5493 19.3944
R23268 GND.n6326 GND.n6325 19.3944
R23269 GND.n6329 GND.n6326 19.3944
R23270 GND.n6329 GND.n5491 19.3944
R23271 GND.n6335 GND.n5491 19.3944
R23272 GND.n6336 GND.n6335 19.3944
R23273 GND.n6339 GND.n6336 19.3944
R23274 GND.n5490 GND.n5487 19.3944
R23275 GND.n5485 GND.n5482 19.3944
R23276 GND.n5480 GND.n5477 19.3944
R23277 GND.n5475 GND.n5472 19.3944
R23278 GND.n5470 GND.n5467 19.3944
R23279 GND.n6355 GND.n6341 19.3944
R23280 GND.n6355 GND.n6352 19.3944
R23281 GND.n6366 GND.n6363 19.3944
R23282 GND.n6371 GND.n6368 19.3944
R23283 GND.n6376 GND.n6373 19.3944
R23284 GND.n6381 GND.n6378 19.3944
R23285 GND.n7094 GND.n7093 19.3944
R23286 GND.n7093 GND.n4880 19.3944
R23287 GND.n4916 GND.n4880 19.3944
R23288 GND.n4916 GND.n4913 19.3944
R23289 GND.n7074 GND.n4913 19.3944
R23290 GND.n7074 GND.n7073 19.3944
R23291 GND.n7073 GND.n7072 19.3944
R23292 GND.n7072 GND.n4922 19.3944
R23293 GND.n7062 GND.n4922 19.3944
R23294 GND.n7062 GND.n7061 19.3944
R23295 GND.n7061 GND.n7060 19.3944
R23296 GND.n7060 GND.n4944 19.3944
R23297 GND.n7050 GND.n4944 19.3944
R23298 GND.n7050 GND.n7049 19.3944
R23299 GND.n7049 GND.n7048 19.3944
R23300 GND.n7048 GND.n4965 19.3944
R23301 GND.n7038 GND.n4965 19.3944
R23302 GND.n7038 GND.n7037 19.3944
R23303 GND.n7037 GND.n7036 19.3944
R23304 GND.n7036 GND.n4986 19.3944
R23305 GND.n7026 GND.n4986 19.3944
R23306 GND.n7026 GND.n7025 19.3944
R23307 GND.n7025 GND.n7024 19.3944
R23308 GND.n7024 GND.n5006 19.3944
R23309 GND.n7014 GND.n5006 19.3944
R23310 GND.n7014 GND.n7013 19.3944
R23311 GND.n7013 GND.n7012 19.3944
R23312 GND.n7012 GND.n5027 19.3944
R23313 GND.n7002 GND.n5027 19.3944
R23314 GND.n7002 GND.n7001 19.3944
R23315 GND.n7001 GND.n7000 19.3944
R23316 GND.n7000 GND.n5048 19.3944
R23317 GND.n6990 GND.n5048 19.3944
R23318 GND.n6990 GND.n6989 19.3944
R23319 GND.n6989 GND.n6988 19.3944
R23320 GND.n6988 GND.n5069 19.3944
R23321 GND.n6978 GND.n5069 19.3944
R23322 GND.n6978 GND.n6977 19.3944
R23323 GND.n6977 GND.n6976 19.3944
R23324 GND.n6976 GND.n5090 19.3944
R23325 GND.n6966 GND.n5090 19.3944
R23326 GND.n6966 GND.n6965 19.3944
R23327 GND.n6965 GND.n6964 19.3944
R23328 GND.n6964 GND.n5111 19.3944
R23329 GND.n6954 GND.n5111 19.3944
R23330 GND.n6954 GND.n6953 19.3944
R23331 GND.n6953 GND.n6952 19.3944
R23332 GND.n6952 GND.n5132 19.3944
R23333 GND.n6942 GND.n5132 19.3944
R23334 GND.n6942 GND.n6941 19.3944
R23335 GND.n6941 GND.n6940 19.3944
R23336 GND.n6940 GND.n5153 19.3944
R23337 GND.n6930 GND.n5153 19.3944
R23338 GND.n6930 GND.n6929 19.3944
R23339 GND.n6929 GND.n6928 19.3944
R23340 GND.n6928 GND.n5173 19.3944
R23341 GND.n6918 GND.n121 19.3944
R23342 GND.n5188 GND.n121 19.3944
R23343 GND.n10308 GND.n114 19.3944
R23344 GND.n5267 GND.n115 19.3944
R23345 GND.n10305 GND.n123 19.3944
R23346 GND.n10305 GND.n124 19.3944
R23347 GND.n10295 GND.n124 19.3944
R23348 GND.n10295 GND.n10294 19.3944
R23349 GND.n10294 GND.n10293 19.3944
R23350 GND.n10293 GND.n147 19.3944
R23351 GND.n10283 GND.n147 19.3944
R23352 GND.n10283 GND.n10282 19.3944
R23353 GND.n10282 GND.n10281 19.3944
R23354 GND.n10281 GND.n168 19.3944
R23355 GND.n10271 GND.n168 19.3944
R23356 GND.n10271 GND.n10270 19.3944
R23357 GND.n10270 GND.n10269 19.3944
R23358 GND.n10269 GND.n189 19.3944
R23359 GND.n10259 GND.n189 19.3944
R23360 GND.n10259 GND.n10258 19.3944
R23361 GND.n10258 GND.n10257 19.3944
R23362 GND.n10257 GND.n210 19.3944
R23363 GND.n10247 GND.n210 19.3944
R23364 GND.n10247 GND.n10246 19.3944
R23365 GND.n10246 GND.n10245 19.3944
R23366 GND.n10245 GND.n231 19.3944
R23367 GND.n10235 GND.n231 19.3944
R23368 GND.n10235 GND.n10234 19.3944
R23369 GND.n10234 GND.n10233 19.3944
R23370 GND.n10233 GND.n252 19.3944
R23371 GND.n10223 GND.n252 19.3944
R23372 GND.n10223 GND.n10222 19.3944
R23373 GND.n10222 GND.n10221 19.3944
R23374 GND.n10221 GND.n272 19.3944
R23375 GND.n10211 GND.n272 19.3944
R23376 GND.n10211 GND.n10210 19.3944
R23377 GND.n10210 GND.n10209 19.3944
R23378 GND.n10209 GND.n293 19.3944
R23379 GND.n10199 GND.n293 19.3944
R23380 GND.n10199 GND.n10198 19.3944
R23381 GND.n10198 GND.n10197 19.3944
R23382 GND.n10197 GND.n314 19.3944
R23383 GND.n10187 GND.n314 19.3944
R23384 GND.n10187 GND.n10186 19.3944
R23385 GND.n10186 GND.n10185 19.3944
R23386 GND.n10185 GND.n335 19.3944
R23387 GND.n10175 GND.n335 19.3944
R23388 GND.n10175 GND.n10174 19.3944
R23389 GND.n10174 GND.n10173 19.3944
R23390 GND.n10173 GND.n356 19.3944
R23391 GND.n10163 GND.n356 19.3944
R23392 GND.n10163 GND.n10162 19.3944
R23393 GND.n10162 GND.n10161 19.3944
R23394 GND.n10161 GND.n376 19.3944
R23395 GND.n10151 GND.n376 19.3944
R23396 GND.n10151 GND.n10150 19.3944
R23397 GND.n10150 GND.n10149 19.3944
R23398 GND.n10149 GND.n395 19.3944
R23399 GND.n10139 GND.n395 19.3944
R23400 GND.n10139 GND.n10138 19.3944
R23401 GND.n10138 GND.n10137 19.3944
R23402 GND.n3009 GND.n3008 19.3944
R23403 GND.n3015 GND.n3008 19.3944
R23404 GND.n3015 GND.n3014 19.3944
R23405 GND.n3014 GND.n2838 19.3944
R23406 GND.n3038 GND.n2838 19.3944
R23407 GND.n3038 GND.n2836 19.3944
R23408 GND.n3042 GND.n2836 19.3944
R23409 GND.n3042 GND.n2811 19.3944
R23410 GND.n3073 GND.n2811 19.3944
R23411 GND.n3073 GND.n2809 19.3944
R23412 GND.n3079 GND.n2809 19.3944
R23413 GND.n3079 GND.n3078 19.3944
R23414 GND.n3078 GND.n2782 19.3944
R23415 GND.n3110 GND.n2782 19.3944
R23416 GND.n3110 GND.n2780 19.3944
R23417 GND.n3116 GND.n2780 19.3944
R23418 GND.n3116 GND.n3115 19.3944
R23419 GND.n3115 GND.n2754 19.3944
R23420 GND.n3148 GND.n2754 19.3944
R23421 GND.n3148 GND.n2752 19.3944
R23422 GND.n3154 GND.n2752 19.3944
R23423 GND.n3154 GND.n3153 19.3944
R23424 GND.n3153 GND.n2726 19.3944
R23425 GND.n3186 GND.n2726 19.3944
R23426 GND.n3186 GND.n2724 19.3944
R23427 GND.n3192 GND.n2724 19.3944
R23428 GND.n3192 GND.n3191 19.3944
R23429 GND.n3191 GND.n2696 19.3944
R23430 GND.n3223 GND.n2696 19.3944
R23431 GND.n3223 GND.n2694 19.3944
R23432 GND.n3229 GND.n2694 19.3944
R23433 GND.n3229 GND.n3228 19.3944
R23434 GND.n3228 GND.n2667 19.3944
R23435 GND.n3260 GND.n2667 19.3944
R23436 GND.n3260 GND.n2665 19.3944
R23437 GND.n3266 GND.n2665 19.3944
R23438 GND.n3266 GND.n3265 19.3944
R23439 GND.n3265 GND.n2638 19.3944
R23440 GND.n3298 GND.n2638 19.3944
R23441 GND.n3298 GND.n2636 19.3944
R23442 GND.n3304 GND.n2636 19.3944
R23443 GND.n3304 GND.n3303 19.3944
R23444 GND.n3330 GND.n2613 19.3944
R23445 GND.n3539 GND.n3332 19.3944
R23446 GND.n3537 GND.n3536 19.3944
R23447 GND.n3533 GND.n3532 19.3944
R23448 GND.n3530 GND.n3335 19.3944
R23449 GND.n3526 GND.n3335 19.3944
R23450 GND.n3526 GND.n3525 19.3944
R23451 GND.n3525 GND.n3524 19.3944
R23452 GND.n3524 GND.n3341 19.3944
R23453 GND.n3520 GND.n3341 19.3944
R23454 GND.n3520 GND.n3519 19.3944
R23455 GND.n3519 GND.n3518 19.3944
R23456 GND.n3518 GND.n3347 19.3944
R23457 GND.n3514 GND.n3347 19.3944
R23458 GND.n3514 GND.n3513 19.3944
R23459 GND.n3513 GND.n3512 19.3944
R23460 GND.n3512 GND.n3353 19.3944
R23461 GND.n3508 GND.n3353 19.3944
R23462 GND.n3508 GND.n3507 19.3944
R23463 GND.n3507 GND.n3506 19.3944
R23464 GND.n3506 GND.n3359 19.3944
R23465 GND.n3502 GND.n3359 19.3944
R23466 GND.n3502 GND.n3501 19.3944
R23467 GND.n3501 GND.n3500 19.3944
R23468 GND.n3500 GND.n3365 19.3944
R23469 GND.n3496 GND.n3365 19.3944
R23470 GND.n3496 GND.n3495 19.3944
R23471 GND.n3495 GND.n3494 19.3944
R23472 GND.n3494 GND.n3371 19.3944
R23473 GND.n3490 GND.n3371 19.3944
R23474 GND.n3490 GND.n3489 19.3944
R23475 GND.n3489 GND.n3488 19.3944
R23476 GND.n3488 GND.n3377 19.3944
R23477 GND.n3484 GND.n3377 19.3944
R23478 GND.n3484 GND.n3483 19.3944
R23479 GND.n3483 GND.n3482 19.3944
R23480 GND.n3482 GND.n3383 19.3944
R23481 GND.n3478 GND.n3383 19.3944
R23482 GND.n3478 GND.n3477 19.3944
R23483 GND.n3477 GND.n3476 19.3944
R23484 GND.n3476 GND.n3389 19.3944
R23485 GND.n3470 GND.n3389 19.3944
R23486 GND.n3470 GND.n3469 19.3944
R23487 GND.n3469 GND.n3468 19.3944
R23488 GND.n3468 GND.n3395 19.3944
R23489 GND.n3464 GND.n3395 19.3944
R23490 GND.n3464 GND.n3463 19.3944
R23491 GND.n3463 GND.n3462 19.3944
R23492 GND.n3462 GND.n3401 19.3944
R23493 GND.n3458 GND.n3401 19.3944
R23494 GND.n3458 GND.n3457 19.3944
R23495 GND.n3457 GND.n3456 19.3944
R23496 GND.n3456 GND.n3407 19.3944
R23497 GND.n3452 GND.n3407 19.3944
R23498 GND.n3452 GND.n3451 19.3944
R23499 GND.n3451 GND.n3450 19.3944
R23500 GND.n3450 GND.n3413 19.3944
R23501 GND.n3446 GND.n3413 19.3944
R23502 GND.n3446 GND.n3445 19.3944
R23503 GND.n3445 GND.n3444 19.3944
R23504 GND.n3444 GND.n3419 19.3944
R23505 GND.n3440 GND.n3419 19.3944
R23506 GND.n3440 GND.n3439 19.3944
R23507 GND.n3439 GND.n3438 19.3944
R23508 GND.n3438 GND.n3425 19.3944
R23509 GND.n3432 GND.n3425 19.3944
R23510 GND.n3432 GND.n3431 19.3944
R23511 GND.n3431 GND.n1941 19.3944
R23512 GND.n7908 GND.n1941 19.3944
R23513 GND.n7908 GND.n7907 19.3944
R23514 GND.n7907 GND.n7906 19.3944
R23515 GND.n7906 GND.n1945 19.3944
R23516 GND.n7895 GND.n1945 19.3944
R23517 GND.n7895 GND.n7894 19.3944
R23518 GND.n7894 GND.n7893 19.3944
R23519 GND.n7893 GND.n1962 19.3944
R23520 GND.n7881 GND.n1962 19.3944
R23521 GND.n7881 GND.n7880 19.3944
R23522 GND.n7880 GND.n7879 19.3944
R23523 GND.n7879 GND.n1979 19.3944
R23524 GND.n7867 GND.n1979 19.3944
R23525 GND.n7867 GND.n7866 19.3944
R23526 GND.n7866 GND.n7865 19.3944
R23527 GND.n7865 GND.n1997 19.3944
R23528 GND.n7853 GND.n1997 19.3944
R23529 GND.n7853 GND.n7852 19.3944
R23530 GND.n7852 GND.n7851 19.3944
R23531 GND.n7851 GND.n2015 19.3944
R23532 GND.n7839 GND.n2015 19.3944
R23533 GND.n7839 GND.n7838 19.3944
R23534 GND.n7838 GND.n7837 19.3944
R23535 GND.n7837 GND.n2033 19.3944
R23536 GND.n7825 GND.n2033 19.3944
R23537 GND.n7825 GND.n7824 19.3944
R23538 GND.n7824 GND.n7823 19.3944
R23539 GND.n7823 GND.n2051 19.3944
R23540 GND.n7811 GND.n2051 19.3944
R23541 GND.n7811 GND.n7810 19.3944
R23542 GND.n7810 GND.n7809 19.3944
R23543 GND.n7809 GND.n2069 19.3944
R23544 GND.n7797 GND.n2069 19.3944
R23545 GND.n7797 GND.n7796 19.3944
R23546 GND.n7796 GND.n7795 19.3944
R23547 GND.n7795 GND.n2087 19.3944
R23548 GND.n7783 GND.n2087 19.3944
R23549 GND.n7783 GND.n7782 19.3944
R23550 GND.n7782 GND.n7781 19.3944
R23551 GND.n7781 GND.n2105 19.3944
R23552 GND.n2319 GND.n2105 19.3944
R23553 GND.n7764 GND.n2319 19.3944
R23554 GND.n7764 GND.n7763 19.3944
R23555 GND.n7763 GND.n7762 19.3944
R23556 GND.n7762 GND.n2325 19.3944
R23557 GND.n7695 GND.n2325 19.3944
R23558 GND.n7695 GND.n7694 19.3944
R23559 GND.n7694 GND.n7693 19.3944
R23560 GND.n7693 GND.n3892 19.3944
R23561 GND.n7684 GND.n3892 19.3944
R23562 GND.n7684 GND.n7683 19.3944
R23563 GND.n7683 GND.n7682 19.3944
R23564 GND.n7682 GND.n3911 19.3944
R23565 GND.n7672 GND.n3911 19.3944
R23566 GND.n7672 GND.n7671 19.3944
R23567 GND.n7671 GND.n7670 19.3944
R23568 GND.n7670 GND.n3931 19.3944
R23569 GND.n3956 GND.n3931 19.3944
R23570 GND.n7653 GND.n3956 19.3944
R23571 GND.n7653 GND.n7652 19.3944
R23572 GND.n7652 GND.n7651 19.3944
R23573 GND.n7651 GND.n3962 19.3944
R23574 GND.n7641 GND.n3962 19.3944
R23575 GND.n7641 GND.n7640 19.3944
R23576 GND.n7640 GND.n7639 19.3944
R23577 GND.n7639 GND.n3995 19.3944
R23578 GND.n7629 GND.n3995 19.3944
R23579 GND.n7629 GND.n7628 19.3944
R23580 GND.n7628 GND.n7627 19.3944
R23581 GND.n7627 GND.n4015 19.3944
R23582 GND.n7617 GND.n4015 19.3944
R23583 GND.n7617 GND.n7616 19.3944
R23584 GND.n7616 GND.n7615 19.3944
R23585 GND.n7615 GND.n4035 19.3944
R23586 GND.n4061 GND.n4035 19.3944
R23587 GND.n7598 GND.n4061 19.3944
R23588 GND.n7598 GND.n7597 19.3944
R23589 GND.n7597 GND.n7596 19.3944
R23590 GND.n7596 GND.n4067 19.3944
R23591 GND.n7586 GND.n4067 19.3944
R23592 GND.n7586 GND.n7585 19.3944
R23593 GND.n7585 GND.n7584 19.3944
R23594 GND.n7584 GND.n4100 19.3944
R23595 GND.n7574 GND.n4100 19.3944
R23596 GND.n7574 GND.n7573 19.3944
R23597 GND.n7573 GND.n7572 19.3944
R23598 GND.n7572 GND.n4120 19.3944
R23599 GND.n7562 GND.n4120 19.3944
R23600 GND.n7562 GND.n7561 19.3944
R23601 GND.n7561 GND.n7560 19.3944
R23602 GND.n7560 GND.n4140 19.3944
R23603 GND.n4166 GND.n4140 19.3944
R23604 GND.n7543 GND.n4166 19.3944
R23605 GND.n7543 GND.n7542 19.3944
R23606 GND.n7542 GND.n7541 19.3944
R23607 GND.n7541 GND.n4172 19.3944
R23608 GND.n7531 GND.n4172 19.3944
R23609 GND.n7531 GND.n7530 19.3944
R23610 GND.n7530 GND.n7529 19.3944
R23611 GND.n7529 GND.n4204 19.3944
R23612 GND.n7519 GND.n4204 19.3944
R23613 GND.n7519 GND.n7518 19.3944
R23614 GND.n7518 GND.n7517 19.3944
R23615 GND.n7517 GND.n4224 19.3944
R23616 GND.n7507 GND.n4224 19.3944
R23617 GND.n7507 GND.n7506 19.3944
R23618 GND.n7506 GND.n7505 19.3944
R23619 GND.n7505 GND.n4243 19.3944
R23620 GND.n4269 GND.n4243 19.3944
R23621 GND.n7488 GND.n4269 19.3944
R23622 GND.n7488 GND.n7487 19.3944
R23623 GND.n7487 GND.n7486 19.3944
R23624 GND.n7486 GND.n4275 19.3944
R23625 GND.n7476 GND.n4275 19.3944
R23626 GND.n7476 GND.n7475 19.3944
R23627 GND.n7475 GND.n7474 19.3944
R23628 GND.n7474 GND.n4307 19.3944
R23629 GND.n7464 GND.n4307 19.3944
R23630 GND.n7464 GND.n7463 19.3944
R23631 GND.n7463 GND.n7462 19.3944
R23632 GND.n7462 GND.n4327 19.3944
R23633 GND.n7452 GND.n4327 19.3944
R23634 GND.n7452 GND.n7451 19.3944
R23635 GND.n7451 GND.n7450 19.3944
R23636 GND.n7450 GND.n4347 19.3944
R23637 GND.n4373 GND.n4347 19.3944
R23638 GND.n7433 GND.n4373 19.3944
R23639 GND.n7433 GND.n7432 19.3944
R23640 GND.n7432 GND.n7431 19.3944
R23641 GND.n7431 GND.n4379 19.3944
R23642 GND.n7421 GND.n4379 19.3944
R23643 GND.n7421 GND.n7420 19.3944
R23644 GND.n7420 GND.n7419 19.3944
R23645 GND.n7419 GND.n4412 19.3944
R23646 GND.n4439 GND.n4412 19.3944
R23647 GND.n7405 GND.n4439 19.3944
R23648 GND.n7405 GND.n7404 19.3944
R23649 GND.n7404 GND.n7403 19.3944
R23650 GND.n7403 GND.n4445 19.3944
R23651 GND.n7391 GND.n4445 19.3944
R23652 GND.n7391 GND.n7390 19.3944
R23653 GND.n7390 GND.n7389 19.3944
R23654 GND.n7389 GND.n4463 19.3944
R23655 GND.n7377 GND.n4463 19.3944
R23656 GND.n7377 GND.n7376 19.3944
R23657 GND.n7376 GND.n7375 19.3944
R23658 GND.n7375 GND.n4481 19.3944
R23659 GND.n7363 GND.n4481 19.3944
R23660 GND.n7363 GND.n7362 19.3944
R23661 GND.n7362 GND.n7361 19.3944
R23662 GND.n7361 GND.n4499 19.3944
R23663 GND.n7349 GND.n4499 19.3944
R23664 GND.n7349 GND.n7348 19.3944
R23665 GND.n7348 GND.n7347 19.3944
R23666 GND.n7347 GND.n4517 19.3944
R23667 GND.n7335 GND.n4517 19.3944
R23668 GND.n7335 GND.n7334 19.3944
R23669 GND.n7334 GND.n7333 19.3944
R23670 GND.n7333 GND.n4535 19.3944
R23671 GND.n4561 GND.n4535 19.3944
R23672 GND.n7316 GND.n4561 19.3944
R23673 GND.n7316 GND.n7315 19.3944
R23674 GND.n7315 GND.n7314 19.3944
R23675 GND.n7314 GND.n4567 19.3944
R23676 GND.n7302 GND.n4567 19.3944
R23677 GND.n7302 GND.n7301 19.3944
R23678 GND.n7301 GND.n7300 19.3944
R23679 GND.n7300 GND.n4585 19.3944
R23680 GND.n7288 GND.n4585 19.3944
R23681 GND.n7288 GND.n7287 19.3944
R23682 GND.n7287 GND.n7286 19.3944
R23683 GND.n7286 GND.n4603 19.3944
R23684 GND.n7274 GND.n4603 19.3944
R23685 GND.n7274 GND.n7273 19.3944
R23686 GND.n7273 GND.n7272 19.3944
R23687 GND.n7272 GND.n4620 19.3944
R23688 GND.n4692 GND.n4620 19.3944
R23689 GND.n7255 GND.n4692 19.3944
R23690 GND.n7255 GND.n7254 19.3944
R23691 GND.n7254 GND.n7253 19.3944
R23692 GND.n7253 GND.n4698 19.3944
R23693 GND.n6398 GND.n4698 19.3944
R23694 GND.n6398 GND.n6397 19.3944
R23695 GND.n6397 GND.n6392 19.3944
R23696 GND.n6405 GND.n6392 19.3944
R23697 GND.n6405 GND.n6390 19.3944
R23698 GND.n6412 GND.n6390 19.3944
R23699 GND.n6412 GND.n6411 19.3944
R23700 GND.n6411 GND.n4899 19.3944
R23701 GND.n7081 GND.n4899 19.3944
R23702 GND.n7081 GND.n7080 19.3944
R23703 GND.n7080 GND.n7079 19.3944
R23704 GND.n7079 GND.n4903 19.3944
R23705 GND.n6470 GND.n4903 19.3944
R23706 GND.n6470 GND.n6469 19.3944
R23707 GND.n6469 GND.n6468 19.3944
R23708 GND.n6468 GND.n6437 19.3944
R23709 GND.n6464 GND.n6437 19.3944
R23710 GND.n6464 GND.n6463 19.3944
R23711 GND.n6463 GND.n6462 19.3944
R23712 GND.n6462 GND.n6443 19.3944
R23713 GND.n6458 GND.n6443 19.3944
R23714 GND.n6458 GND.n6457 19.3944
R23715 GND.n6457 GND.n6456 19.3944
R23716 GND.n6456 GND.n6449 19.3944
R23717 GND.n6452 GND.n6449 19.3944
R23718 GND.n6452 GND.n5328 19.3944
R23719 GND.n6678 GND.n5328 19.3944
R23720 GND.n6678 GND.n5326 19.3944
R23721 GND.n6682 GND.n5326 19.3944
R23722 GND.n6682 GND.n5324 19.3944
R23723 GND.n6686 GND.n5324 19.3944
R23724 GND.n6686 GND.n5322 19.3944
R23725 GND.n6690 GND.n5322 19.3944
R23726 GND.n6690 GND.n5320 19.3944
R23727 GND.n6694 GND.n5320 19.3944
R23728 GND.n6694 GND.n5318 19.3944
R23729 GND.n6698 GND.n5318 19.3944
R23730 GND.n6698 GND.n5316 19.3944
R23731 GND.n6702 GND.n5316 19.3944
R23732 GND.n6702 GND.n5314 19.3944
R23733 GND.n6706 GND.n5314 19.3944
R23734 GND.n6706 GND.n5312 19.3944
R23735 GND.n6710 GND.n5312 19.3944
R23736 GND.n6710 GND.n5310 19.3944
R23737 GND.n6714 GND.n5310 19.3944
R23738 GND.n6714 GND.n5308 19.3944
R23739 GND.n6718 GND.n5308 19.3944
R23740 GND.n6718 GND.n5306 19.3944
R23741 GND.n6722 GND.n5306 19.3944
R23742 GND.n6722 GND.n5304 19.3944
R23743 GND.n6726 GND.n5304 19.3944
R23744 GND.n6726 GND.n5302 19.3944
R23745 GND.n6730 GND.n5302 19.3944
R23746 GND.n6730 GND.n5300 19.3944
R23747 GND.n6734 GND.n5300 19.3944
R23748 GND.n6734 GND.n5298 19.3944
R23749 GND.n6738 GND.n5298 19.3944
R23750 GND.n6738 GND.n5296 19.3944
R23751 GND.n6742 GND.n5296 19.3944
R23752 GND.n6742 GND.n5294 19.3944
R23753 GND.n6751 GND.n5294 19.3944
R23754 GND.n6751 GND.n6750 19.3944
R23755 GND.n6750 GND.n6749 19.3944
R23756 GND.n6913 GND.n5195 19.3944
R23757 GND.n6911 GND.n6910 19.3944
R23758 GND.n6907 GND.n6906 19.3944
R23759 GND.n6904 GND.n5198 19.3944
R23760 GND.n5264 GND.n5263 19.3944
R23761 GND.n5263 GND.n5262 19.3944
R23762 GND.n5262 GND.n5203 19.3944
R23763 GND.n5258 GND.n5203 19.3944
R23764 GND.n5258 GND.n5257 19.3944
R23765 GND.n5257 GND.n5256 19.3944
R23766 GND.n5256 GND.n5209 19.3944
R23767 GND.n5252 GND.n5209 19.3944
R23768 GND.n5252 GND.n5251 19.3944
R23769 GND.n5251 GND.n5250 19.3944
R23770 GND.n5250 GND.n5215 19.3944
R23771 GND.n5246 GND.n5215 19.3944
R23772 GND.n5246 GND.n5245 19.3944
R23773 GND.n5245 GND.n5244 19.3944
R23774 GND.n5244 GND.n5221 19.3944
R23775 GND.n5240 GND.n5221 19.3944
R23776 GND.n5240 GND.n5239 19.3944
R23777 GND.n5239 GND.n5238 19.3944
R23778 GND.n5238 GND.n5227 19.3944
R23779 GND.n5234 GND.n5227 19.3944
R23780 GND.n5234 GND.n5233 19.3944
R23781 GND.n5233 GND.n444 19.3944
R23782 GND.n9724 GND.n444 19.3944
R23783 GND.n9724 GND.n9723 19.3944
R23784 GND.n9723 GND.n9722 19.3944
R23785 GND.n9722 GND.n448 19.3944
R23786 GND.n9718 GND.n448 19.3944
R23787 GND.n9718 GND.n9717 19.3944
R23788 GND.n9717 GND.n9716 19.3944
R23789 GND.n9716 GND.n454 19.3944
R23790 GND.n9712 GND.n454 19.3944
R23791 GND.n9712 GND.n9711 19.3944
R23792 GND.n9711 GND.n9710 19.3944
R23793 GND.n9710 GND.n460 19.3944
R23794 GND.n9706 GND.n460 19.3944
R23795 GND.n9706 GND.n9705 19.3944
R23796 GND.n9705 GND.n9704 19.3944
R23797 GND.n9704 GND.n466 19.3944
R23798 GND.n9700 GND.n466 19.3944
R23799 GND.n9700 GND.n9699 19.3944
R23800 GND.n9699 GND.n9698 19.3944
R23801 GND.n9698 GND.n472 19.3944
R23802 GND.n8359 GND.n8358 19.3944
R23803 GND.n8358 GND.n8357 19.3944
R23804 GND.n8357 GND.n8356 19.3944
R23805 GND.n8356 GND.n8354 19.3944
R23806 GND.n8354 GND.n8351 19.3944
R23807 GND.n8351 GND.n8350 19.3944
R23808 GND.n8350 GND.n8347 19.3944
R23809 GND.n8347 GND.n8346 19.3944
R23810 GND.n8346 GND.n8343 19.3944
R23811 GND.n8341 GND.n8339 19.3944
R23812 GND.n8339 GND.n8336 19.3944
R23813 GND.n8336 GND.n8335 19.3944
R23814 GND.n8335 GND.n8332 19.3944
R23815 GND.n8332 GND.n8331 19.3944
R23816 GND.n8331 GND.n8328 19.3944
R23817 GND.n8328 GND.n8327 19.3944
R23818 GND.n8327 GND.n8324 19.3944
R23819 GND.n8324 GND.n8323 19.3944
R23820 GND.n8323 GND.n8320 19.3944
R23821 GND.n8320 GND.n8319 19.3944
R23822 GND.n8316 GND.n8315 19.3944
R23823 GND.n8315 GND.n8312 19.3944
R23824 GND.n8312 GND.n8311 19.3944
R23825 GND.n8311 GND.n8308 19.3944
R23826 GND.n8308 GND.n8307 19.3944
R23827 GND.n8307 GND.n8304 19.3944
R23828 GND.n8304 GND.n8303 19.3944
R23829 GND.n8303 GND.n8300 19.3944
R23830 GND.n8300 GND.n8299 19.3944
R23831 GND.n8299 GND.n8296 19.3944
R23832 GND.n8296 GND.n8295 19.3944
R23833 GND.n8291 GND.n8288 19.3944
R23834 GND.n8288 GND.n8287 19.3944
R23835 GND.n8287 GND.n8284 19.3944
R23836 GND.n8284 GND.n8283 19.3944
R23837 GND.n8283 GND.n8280 19.3944
R23838 GND.n8280 GND.n8279 19.3944
R23839 GND.n8279 GND.n8276 19.3944
R23840 GND.n8276 GND.n8275 19.3944
R23841 GND.n8275 GND.n8272 19.3944
R23842 GND.n8272 GND.n8271 19.3944
R23843 GND.n8271 GND.n8268 19.3944
R23844 GND.n8266 GND.n8263 19.3944
R23845 GND.n8263 GND.n8262 19.3944
R23846 GND.n8262 GND.n8259 19.3944
R23847 GND.n8259 GND.n8258 19.3944
R23848 GND.n8258 GND.n8255 19.3944
R23849 GND.n8255 GND.n8254 19.3944
R23850 GND.n8254 GND.n8251 19.3944
R23851 GND.n8251 GND.n8250 19.3944
R23852 GND.n8250 GND.n8247 19.3944
R23853 GND.n8247 GND.n8246 19.3944
R23854 GND.n8246 GND.n8243 19.3944
R23855 GND.n2938 GND.n2937 19.3944
R23856 GND.n2942 GND.n2937 19.3944
R23857 GND.n2942 GND.n2909 19.3944
R23858 GND.n2955 GND.n2909 19.3944
R23859 GND.n2955 GND.n2907 19.3944
R23860 GND.n2959 GND.n2907 19.3944
R23861 GND.n2959 GND.n2889 19.3944
R23862 GND.n2972 GND.n2889 19.3944
R23863 GND.n2972 GND.n2887 19.3944
R23864 GND.n2976 GND.n2887 19.3944
R23865 GND.n2976 GND.n2870 19.3944
R23866 GND.n2996 GND.n2870 19.3944
R23867 GND.n2996 GND.n2868 19.3944
R23868 GND.n3002 GND.n2868 19.3944
R23869 GND.n3002 GND.n3001 19.3944
R23870 GND.n3001 GND.n2846 19.3944
R23871 GND.n3029 GND.n2846 19.3944
R23872 GND.n3029 GND.n2844 19.3944
R23873 GND.n3033 GND.n2844 19.3944
R23874 GND.n3033 GND.n2822 19.3944
R23875 GND.n3062 GND.n2822 19.3944
R23876 GND.n3062 GND.n2820 19.3944
R23877 GND.n3068 GND.n2820 19.3944
R23878 GND.n3068 GND.n3067 19.3944
R23879 GND.n3067 GND.n2793 19.3944
R23880 GND.n3099 GND.n2793 19.3944
R23881 GND.n3099 GND.n2791 19.3944
R23882 GND.n3105 GND.n2791 19.3944
R23883 GND.n3105 GND.n3104 19.3944
R23884 GND.n3104 GND.n2763 19.3944
R23885 GND.n3137 GND.n2763 19.3944
R23886 GND.n3137 GND.n2761 19.3944
R23887 GND.n3143 GND.n2761 19.3944
R23888 GND.n3143 GND.n3142 19.3944
R23889 GND.n3142 GND.n2736 19.3944
R23890 GND.n3175 GND.n2736 19.3944
R23891 GND.n3175 GND.n2734 19.3944
R23892 GND.n3181 GND.n2734 19.3944
R23893 GND.n3181 GND.n3180 19.3944
R23894 GND.n3180 GND.n2707 19.3944
R23895 GND.n3212 GND.n2707 19.3944
R23896 GND.n3212 GND.n2705 19.3944
R23897 GND.n3218 GND.n2705 19.3944
R23898 GND.n3218 GND.n3217 19.3944
R23899 GND.n3217 GND.n2678 19.3944
R23900 GND.n3249 GND.n2678 19.3944
R23901 GND.n3249 GND.n2676 19.3944
R23902 GND.n3255 GND.n2676 19.3944
R23903 GND.n3255 GND.n3254 19.3944
R23904 GND.n3254 GND.n2648 19.3944
R23905 GND.n3286 GND.n2648 19.3944
R23906 GND.n3286 GND.n2646 19.3944
R23907 GND.n3293 GND.n2646 19.3944
R23908 GND.n3293 GND.n3292 19.3944
R23909 GND.n3292 GND.n3291 19.3944
R23910 GND.n3291 GND.n2621 19.3944
R23911 GND.n3322 GND.n1546 19.3944
R23912 GND.n3324 GND.n1546 19.3944
R23913 GND.n8121 GND.n1539 19.3944
R23914 GND.n3554 GND.n1540 19.3944
R23915 GND.n8118 GND.n1548 19.3944
R23916 GND.n8118 GND.n1549 19.3944
R23917 GND.n2581 GND.n1549 19.3944
R23918 GND.n3577 GND.n2581 19.3944
R23919 GND.n3577 GND.n2579 19.3944
R23920 GND.n3583 GND.n2579 19.3944
R23921 GND.n3583 GND.n3582 19.3944
R23922 GND.n3582 GND.n2559 19.3944
R23923 GND.n3603 GND.n2559 19.3944
R23924 GND.n3603 GND.n2557 19.3944
R23925 GND.n3609 GND.n2557 19.3944
R23926 GND.n3609 GND.n3608 19.3944
R23927 GND.n3608 GND.n2538 19.3944
R23928 GND.n3629 GND.n2538 19.3944
R23929 GND.n3629 GND.n2536 19.3944
R23930 GND.n3635 GND.n2536 19.3944
R23931 GND.n3635 GND.n3634 19.3944
R23932 GND.n3634 GND.n2516 19.3944
R23933 GND.n3655 GND.n2516 19.3944
R23934 GND.n3655 GND.n2514 19.3944
R23935 GND.n3661 GND.n2514 19.3944
R23936 GND.n3661 GND.n3660 19.3944
R23937 GND.n3660 GND.n2494 19.3944
R23938 GND.n3680 GND.n2494 19.3944
R23939 GND.n3680 GND.n2492 19.3944
R23940 GND.n3686 GND.n2492 19.3944
R23941 GND.n3686 GND.n3685 19.3944
R23942 GND.n3685 GND.n2472 19.3944
R23943 GND.n3706 GND.n2472 19.3944
R23944 GND.n3706 GND.n2470 19.3944
R23945 GND.n3712 GND.n2470 19.3944
R23946 GND.n3712 GND.n3711 19.3944
R23947 GND.n3711 GND.n2451 19.3944
R23948 GND.n3732 GND.n2451 19.3944
R23949 GND.n3732 GND.n2449 19.3944
R23950 GND.n3738 GND.n2449 19.3944
R23951 GND.n3738 GND.n3737 19.3944
R23952 GND.n3737 GND.n2431 19.3944
R23953 GND.n3758 GND.n2431 19.3944
R23954 GND.n3758 GND.n2429 19.3944
R23955 GND.n3764 GND.n2429 19.3944
R23956 GND.n3764 GND.n3763 19.3944
R23957 GND.n3763 GND.n2409 19.3944
R23958 GND.n3783 GND.n2409 19.3944
R23959 GND.n3783 GND.n2407 19.3944
R23960 GND.n3789 GND.n2407 19.3944
R23961 GND.n3789 GND.n3788 19.3944
R23962 GND.n3788 GND.n2387 19.3944
R23963 GND.n3809 GND.n2387 19.3944
R23964 GND.n3809 GND.n2385 19.3944
R23965 GND.n3815 GND.n2385 19.3944
R23966 GND.n3815 GND.n3814 19.3944
R23967 GND.n3814 GND.n2366 19.3944
R23968 GND.n3836 GND.n2366 19.3944
R23969 GND.n3836 GND.n2364 19.3944
R23970 GND.n3841 GND.n2364 19.3944
R23971 GND.n3841 GND.n3840 19.3944
R23972 GND.n8495 GND.n8494 19.3944
R23973 GND.n8494 GND.n8493 19.3944
R23974 GND.n8493 GND.n1193 19.3944
R23975 GND.n8487 GND.n1193 19.3944
R23976 GND.n8487 GND.n8486 19.3944
R23977 GND.n8486 GND.n8485 19.3944
R23978 GND.n8485 GND.n1201 19.3944
R23979 GND.n8479 GND.n1201 19.3944
R23980 GND.n8479 GND.n8478 19.3944
R23981 GND.n8478 GND.n8477 19.3944
R23982 GND.n8477 GND.n1209 19.3944
R23983 GND.n8471 GND.n1209 19.3944
R23984 GND.n8471 GND.n8470 19.3944
R23985 GND.n8470 GND.n8469 19.3944
R23986 GND.n8469 GND.n1217 19.3944
R23987 GND.n8463 GND.n1217 19.3944
R23988 GND.n8463 GND.n8462 19.3944
R23989 GND.n8462 GND.n8461 19.3944
R23990 GND.n8461 GND.n1225 19.3944
R23991 GND.n8455 GND.n1225 19.3944
R23992 GND.n8455 GND.n8454 19.3944
R23993 GND.n8454 GND.n8453 19.3944
R23994 GND.n8453 GND.n1233 19.3944
R23995 GND.n8447 GND.n1233 19.3944
R23996 GND.n8447 GND.n8446 19.3944
R23997 GND.n8446 GND.n8445 19.3944
R23998 GND.n8445 GND.n1241 19.3944
R23999 GND.n8439 GND.n1241 19.3944
R24000 GND.n8439 GND.n8438 19.3944
R24001 GND.n8438 GND.n8437 19.3944
R24002 GND.n8437 GND.n1249 19.3944
R24003 GND.n8431 GND.n1249 19.3944
R24004 GND.n8431 GND.n8430 19.3944
R24005 GND.n8430 GND.n8429 19.3944
R24006 GND.n8429 GND.n1257 19.3944
R24007 GND.n8423 GND.n1257 19.3944
R24008 GND.n8423 GND.n8422 19.3944
R24009 GND.n8422 GND.n8421 19.3944
R24010 GND.n8421 GND.n1265 19.3944
R24011 GND.n8415 GND.n1265 19.3944
R24012 GND.n8415 GND.n8414 19.3944
R24013 GND.n8414 GND.n8413 19.3944
R24014 GND.n8413 GND.n1273 19.3944
R24015 GND.n8407 GND.n1273 19.3944
R24016 GND.n8407 GND.n8406 19.3944
R24017 GND.n8406 GND.n8405 19.3944
R24018 GND.n8405 GND.n1281 19.3944
R24019 GND.n8399 GND.n1281 19.3944
R24020 GND.n8399 GND.n8398 19.3944
R24021 GND.n8398 GND.n8397 19.3944
R24022 GND.n8397 GND.n1289 19.3944
R24023 GND.n8391 GND.n1289 19.3944
R24024 GND.n8391 GND.n8390 19.3944
R24025 GND.n8390 GND.n8389 19.3944
R24026 GND.n8389 GND.n1297 19.3944
R24027 GND.n8383 GND.n1297 19.3944
R24028 GND.n8383 GND.n8382 19.3944
R24029 GND.n8382 GND.n8381 19.3944
R24030 GND.n8381 GND.n1305 19.3944
R24031 GND.n8375 GND.n1305 19.3944
R24032 GND.n8375 GND.n8374 19.3944
R24033 GND.n8374 GND.n8373 19.3944
R24034 GND.n8373 GND.n1313 19.3944
R24035 GND.n8367 GND.n1313 19.3944
R24036 GND.n8367 GND.n8366 19.3944
R24037 GND.n8366 GND.n8365 19.3944
R24038 GND.n2928 GND.n2927 19.3944
R24039 GND.n2934 GND.n2928 19.3944
R24040 GND.n2934 GND.n2916 19.3944
R24041 GND.n2951 GND.n2916 19.3944
R24042 GND.n2951 GND.n2917 19.3944
R24043 GND.n2919 GND.n2917 19.3944
R24044 GND.n2919 GND.n2896 19.3944
R24045 GND.n2968 GND.n2896 19.3944
R24046 GND.n2968 GND.n2897 19.3944
R24047 GND.n2899 GND.n2897 19.3944
R24048 GND.n2899 GND.n2878 19.3944
R24049 GND.n2992 GND.n2878 19.3944
R24050 GND.n2992 GND.n2879 19.3944
R24051 GND.n2983 GND.n2879 19.3944
R24052 GND.n2985 GND.n2983 19.3944
R24053 GND.n2985 GND.n2853 19.3944
R24054 GND.n3025 GND.n2853 19.3944
R24055 GND.n3025 GND.n2854 19.3944
R24056 GND.n2856 GND.n2854 19.3944
R24057 GND.n2856 GND.n2828 19.3944
R24058 GND.n3058 GND.n2828 19.3944
R24059 GND.n3058 GND.n2829 19.3944
R24060 GND.n3049 GND.n2829 19.3944
R24061 GND.n3051 GND.n3049 19.3944
R24062 GND.n3051 GND.n2800 19.3944
R24063 GND.n3095 GND.n2800 19.3944
R24064 GND.n3095 GND.n2801 19.3944
R24065 GND.n3086 GND.n2801 19.3944
R24066 GND.n3088 GND.n3086 19.3944
R24067 GND.n3088 GND.n2771 19.3944
R24068 GND.n3133 GND.n2771 19.3944
R24069 GND.n3133 GND.n2772 19.3944
R24070 GND.n3124 GND.n2772 19.3944
R24071 GND.n3126 GND.n3124 19.3944
R24072 GND.n3126 GND.n2743 19.3944
R24073 GND.n3171 GND.n2743 19.3944
R24074 GND.n3171 GND.n2744 19.3944
R24075 GND.n3162 GND.n2744 19.3944
R24076 GND.n3164 GND.n3162 19.3944
R24077 GND.n3164 GND.n2714 19.3944
R24078 GND.n3208 GND.n2714 19.3944
R24079 GND.n3208 GND.n2715 19.3944
R24080 GND.n3199 GND.n2715 19.3944
R24081 GND.n3201 GND.n3199 19.3944
R24082 GND.n3201 GND.n2685 19.3944
R24083 GND.n3245 GND.n2685 19.3944
R24084 GND.n3245 GND.n2686 19.3944
R24085 GND.n3236 GND.n2686 19.3944
R24086 GND.n3238 GND.n3236 19.3944
R24087 GND.n3238 GND.n2656 19.3944
R24088 GND.n3282 GND.n2656 19.3944
R24089 GND.n3282 GND.n2657 19.3944
R24090 GND.n3273 GND.n2657 19.3944
R24091 GND.n3275 GND.n3273 19.3944
R24092 GND.n3275 GND.n2627 19.3944
R24093 GND.n3318 GND.n2627 19.3944
R24094 GND.n3318 GND.n2628 19.3944
R24095 GND.n3312 GND.n2628 19.3944
R24096 GND.n3312 GND.n2607 19.3944
R24097 GND.n3545 GND.n2607 19.3944
R24098 GND.n3545 GND.n3544 19.3944
R24099 GND.n3544 GND.n2602 19.3944
R24100 GND.n3552 GND.n2602 19.3944
R24101 GND.n3552 GND.n1558 19.3944
R24102 GND.n8114 GND.n1558 19.3944
R24103 GND.n8114 GND.n1559 19.3944
R24104 GND.n1566 GND.n1559 19.3944
R24105 GND.n1567 GND.n1566 19.3944
R24106 GND.n1568 GND.n1567 19.3944
R24107 GND.n2574 GND.n1568 19.3944
R24108 GND.n2574 GND.n1574 19.3944
R24109 GND.n1575 GND.n1574 19.3944
R24110 GND.n1576 GND.n1575 19.3944
R24111 GND.n3597 GND.n1576 19.3944
R24112 GND.n3597 GND.n1582 19.3944
R24113 GND.n1583 GND.n1582 19.3944
R24114 GND.n1584 GND.n1583 19.3944
R24115 GND.n3625 GND.n1584 19.3944
R24116 GND.n3625 GND.n1590 19.3944
R24117 GND.n1591 GND.n1590 19.3944
R24118 GND.n1592 GND.n1591 19.3944
R24119 GND.n2522 GND.n1592 19.3944
R24120 GND.n2522 GND.n1598 19.3944
R24121 GND.n1599 GND.n1598 19.3944
R24122 GND.n1600 GND.n1599 19.3944
R24123 GND.n2500 GND.n1600 19.3944
R24124 GND.n2500 GND.n1606 19.3944
R24125 GND.n1607 GND.n1606 19.3944
R24126 GND.n1608 GND.n1607 19.3944
R24127 GND.n2487 GND.n1608 19.3944
R24128 GND.n2487 GND.n1614 19.3944
R24129 GND.n1615 GND.n1614 19.3944
R24130 GND.n1616 GND.n1615 19.3944
R24131 GND.n3700 GND.n1616 19.3944
R24132 GND.n3700 GND.n1622 19.3944
R24133 GND.n1623 GND.n1622 19.3944
R24134 GND.n1624 GND.n1623 19.3944
R24135 GND.n3728 GND.n1624 19.3944
R24136 GND.n3728 GND.n1630 19.3944
R24137 GND.n1631 GND.n1630 19.3944
R24138 GND.n1632 GND.n1631 19.3944
R24139 GND.n2437 GND.n1632 19.3944
R24140 GND.n2437 GND.n1638 19.3944
R24141 GND.n1639 GND.n1638 19.3944
R24142 GND.n1640 GND.n1639 19.3944
R24143 GND.n2415 GND.n1640 19.3944
R24144 GND.n2415 GND.n1646 19.3944
R24145 GND.n1647 GND.n1646 19.3944
R24146 GND.n1648 GND.n1647 19.3944
R24147 GND.n2402 GND.n1648 19.3944
R24148 GND.n2402 GND.n1654 19.3944
R24149 GND.n1655 GND.n1654 19.3944
R24150 GND.n1656 GND.n1655 19.3944
R24151 GND.n3803 GND.n1656 19.3944
R24152 GND.n3803 GND.n1662 19.3944
R24153 GND.n1663 GND.n1662 19.3944
R24154 GND.n1664 GND.n1663 19.3944
R24155 GND.n3832 GND.n1664 19.3944
R24156 GND.n3832 GND.n1670 19.3944
R24157 GND.n1671 GND.n1670 19.3944
R24158 GND.n1672 GND.n1671 19.3944
R24159 GND.n3856 GND.n3855 19.3944
R24160 GND.n3860 GND.n3859 19.3944
R24161 GND.n3864 GND.n3863 19.3944
R24162 GND.n3868 GND.n3867 19.3944
R24163 GND.n3146 GND.t194 18.592
R24164 GND.n3621 GND.t167 18.592
R24165 GND.n6603 GND.t177 18.592
R24166 GND.n9726 GND.t161 18.592
R24167 GND.n7910 GND.t128 18.2659
R24168 GND.n2195 GND.t113 18.2659
R24169 GND.n7877 GND.n1981 18.2659
R24170 GND.n7856 GND.n2007 18.2659
R24171 GND.n7820 GND.n2055 18.2659
R24172 GND.n7799 GND.n2081 18.2659
R24173 GND.n5690 GND.n2341 18.2659
R24174 GND.t41 GND.n3905 18.2659
R24175 GND.n5643 GND.n3966 18.2659
R24176 GND.n7631 GND.n4009 18.2659
R24177 GND.n5612 GND.n4071 18.2659
R24178 GND.n7576 GND.n4114 18.2659
R24179 GND.n5581 GND.n4176 18.2659
R24180 GND.n7521 GND.n4218 18.2659
R24181 GND.n5548 GND.n5547 18.2659
R24182 GND.n7466 GND.n4321 18.2659
R24183 GND.t152 GND.n4383 18.2659
R24184 GND.n5498 GND.n4422 18.2659
R24185 GND.n7372 GND.n4485 18.2659
R24186 GND.n7351 GND.n4511 18.2659
R24187 GND.n7311 GND.n4571 18.2659
R24188 GND.n7290 GND.n4597 18.2659
R24189 GND.n1932 GND.n1931 18.2581
R24190 GND.n4755 GND.n4754 18.2581
R24191 GND.n1921 GND.n1920 17.9571
R24192 GND.n4752 GND.n4751 17.9571
R24193 GND.t34 GND.n2892 17.9397
R24194 GND.n3804 GND.t22 17.9397
R24195 GND.n7070 GND.t45 17.9397
R24196 GND.t30 GND.n380 17.9397
R24197 GND.n7870 GND.n7869 16.9612
R24198 GND.n2224 GND.n1999 16.9612
R24199 GND.n2275 GND.n2063 16.9612
R24200 GND.n7807 GND.n7806 16.9612
R24201 GND.n5685 GND.n3886 16.9612
R24202 GND.n7691 GND.n3896 16.9612
R24203 GND.n5638 GND.n3989 16.9612
R24204 GND.n7637 GND.n3999 16.9612
R24205 GND.n5607 GND.n4094 16.9612
R24206 GND.n7582 GND.n4104 16.9612
R24207 GND.n5576 GND.n5575 16.9612
R24208 GND.n7527 GND.n4208 16.9612
R24209 GND.n5542 GND.n4301 16.9612
R24210 GND.n7472 GND.n4311 16.9612
R24211 GND.n6194 GND.n4406 16.9612
R24212 GND.n7417 GND.n4415 16.9612
R24213 GND.n6263 GND.n4493 16.9612
R24214 GND.n7359 GND.n7358 16.9612
R24215 GND.n4645 GND.n4579 16.9612
R24216 GND.n7298 GND.n7297 16.9612
R24217 GND.n5862 GND.t267 16.635
R24218 GND.n7491 GND.t9 16.635
R24219 GND.n8005 GND.n1736 16.4853
R24220 GND.n7164 GND.n7163 16.4853
R24221 GND.n9909 GND.n9908 16.4853
R24222 GND.n8343 GND.n8342 16.4853
R24223 GND.n4772 GND.t70 16.3089
R24224 GND.n8224 GND.n8223 15.7096
R24225 GND.n10071 GND.n9810 15.7096
R24226 GND.n6385 GND.n6384 15.7096
R24227 GND.n3872 GND.n3871 15.7096
R24228 GND.n7870 GND.n1989 15.6565
R24229 GND.n7863 GND.n1999 15.6565
R24230 GND.n7813 GND.n2063 15.6565
R24231 GND.n7806 GND.n2073 15.6565
R24232 GND.n7697 GND.n3886 15.6565
R24233 GND.n5664 GND.n3896 15.6565
R24234 GND.n7643 GND.n3989 15.6565
R24235 GND.n5633 GND.n3999 15.6565
R24236 GND.n7588 GND.n4094 15.6565
R24237 GND.n5570 GND.n4208 15.6565
R24238 GND.n7478 GND.n4301 15.6565
R24239 GND.n5537 GND.n4311 15.6565
R24240 GND.n7423 GND.n4406 15.6565
R24241 GND.n6312 GND.n4415 15.6565
R24242 GND.n7365 GND.n4493 15.6565
R24243 GND.n7358 GND.n4503 15.6565
R24244 GND.n7304 GND.n4579 15.6565
R24245 GND.n7297 GND.n4589 15.6565
R24246 GND.n7891 GND.t52 15.0042
R24247 GND.n2961 GND.t34 14.678
R24248 GND.n10153 GND.t30 14.678
R24249 GND.n2211 GND.n1981 14.3519
R24250 GND.n7856 GND.n7855 14.3519
R24251 GND.n7821 GND.n7820 14.3519
R24252 GND.n2288 GND.n2081 14.3519
R24253 GND.n5659 GND.n3905 14.3519
R24254 GND.n7649 GND.n3966 14.3519
R24255 GND.n7594 GND.n4071 14.3519
R24256 GND.n5597 GND.n4114 14.3519
R24257 GND.n7539 GND.n4176 14.3519
R24258 GND.n5565 GND.n4218 14.3519
R24259 GND.n5532 GND.n4321 14.3519
R24260 GND.n7429 GND.n4383 14.3519
R24261 GND.n7373 GND.n7372 14.3519
R24262 GND.n6250 GND.n4511 14.3519
R24263 GND.n7312 GND.n7311 14.3519
R24264 GND.n4658 GND.n4597 14.3519
R24265 GND.n7 GND.t222 14.194
R24266 GND.n7 GND.t198 14.194
R24267 GND.n9 GND.t254 14.194
R24268 GND.n9 GND.t226 14.194
R24269 GND.n11 GND.t251 14.194
R24270 GND.n11 GND.t249 14.194
R24271 GND.n14 GND.t168 14.194
R24272 GND.n14 GND.t244 14.194
R24273 GND.n16 GND.t208 14.194
R24274 GND.n16 GND.t170 14.194
R24275 GND.n18 GND.t195 14.194
R24276 GND.n18 GND.t191 14.194
R24277 GND.n22 GND.t261 14.194
R24278 GND.n22 GND.t196 14.194
R24279 GND.n24 GND.t242 14.194
R24280 GND.n24 GND.t255 14.194
R24281 GND.n26 GND.t228 14.194
R24282 GND.n26 GND.t236 14.194
R24283 GND.n30 GND.t204 14.194
R24284 GND.n30 GND.t166 14.194
R24285 GND.n32 GND.t229 14.194
R24286 GND.n32 GND.t206 14.194
R24287 GND.n34 GND.t221 14.194
R24288 GND.n34 GND.t219 14.194
R24289 GND.n38 GND.t263 14.194
R24290 GND.n38 GND.t250 14.194
R24291 GND.n40 GND.t234 14.194
R24292 GND.n40 GND.t213 14.194
R24293 GND.n42 GND.t212 14.194
R24294 GND.n42 GND.t260 14.194
R24295 GND.n0 GND.t202 14.194
R24296 GND.n0 GND.t179 14.194
R24297 GND.n2 GND.t160 14.194
R24298 GND.n2 GND.t248 14.194
R24299 GND.n4 GND.t245 14.194
R24300 GND.n4 GND.t197 14.194
R24301 GND.n59 GND.t240 14.194
R24302 GND.n59 GND.t162 14.194
R24303 GND.n57 GND.t247 14.194
R24304 GND.n57 GND.t252 14.194
R24305 GND.n55 GND.t211 14.194
R24306 GND.n55 GND.t246 14.194
R24307 GND.n66 GND.t183 14.194
R24308 GND.n66 GND.t216 14.194
R24309 GND.n64 GND.t193 14.194
R24310 GND.n64 GND.t200 14.194
R24311 GND.n62 GND.t156 14.194
R24312 GND.n62 GND.t189 14.194
R24313 GND.n74 GND.t174 14.194
R24314 GND.n74 GND.t264 14.194
R24315 GND.n72 GND.t185 14.194
R24316 GND.n72 GND.t180 14.194
R24317 GND.n70 GND.t232 14.194
R24318 GND.n70 GND.t199 14.194
R24319 GND.n82 GND.t215 14.194
R24320 GND.n82 GND.t243 14.194
R24321 GND.n80 GND.t164 14.194
R24322 GND.n80 GND.t223 14.194
R24323 GND.n78 GND.t186 14.194
R24324 GND.n78 GND.t218 14.194
R24325 GND.n90 GND.t207 14.194
R24326 GND.n90 GND.t224 14.194
R24327 GND.n88 GND.t227 14.194
R24328 GND.n88 GND.t176 14.194
R24329 GND.n86 GND.t262 14.194
R24330 GND.n86 GND.t178 14.194
R24331 GND.n98 GND.t237 14.194
R24332 GND.n98 GND.t258 14.194
R24333 GND.n96 GND.t259 14.194
R24334 GND.n96 GND.t210 14.194
R24335 GND.n94 GND.t201 14.194
R24336 GND.n94 GND.t214 14.194
R24337 GND.n1860 GND.n1774 14.1581
R24338 GND.n1822 GND.n1821 14.1581
R24339 GND.n5393 GND.n5379 14.1581
R24340 GND.n5461 GND.n5460 14.1581
R24341 GND.n10037 GND.n9845 14.1581
R24342 GND.n9971 GND.n9970 14.1581
R24343 GND.n8295 GND.n8292 14.1581
R24344 GND.n8242 GND.n1433 14.1581
R24345 GND.n3220 GND.t190 14.0257
R24346 GND.t169 GND.n2587 14.0257
R24347 GND.n6753 GND.t163 14.0257
R24348 GND.n6859 GND.t173 14.0257
R24349 GND.t88 GND.n7903 13.6995
R24350 GND.n4738 GND.n4737 13.5524
R24351 GND.n7969 GND.n7915 13.4249
R24352 GND.n7247 GND.n4757 13.4249
R24353 GND.n1933 GND.n1909 13.1884
R24354 GND.n1928 GND.n1927 13.1884
R24355 GND.n1927 GND.n1926 13.1884
R24356 GND.n1926 GND.n1912 13.1884
R24357 GND.n1922 GND.n1912 13.1884
R24358 GND.n4740 GND.n4739 13.1884
R24359 GND.n4740 GND.n4735 13.1884
R24360 GND.n4744 GND.n4735 13.1884
R24361 GND.n4745 GND.n4744 13.1884
R24362 GND.n2187 GND.n2186 13.0472
R24363 GND.n7849 GND.n2017 13.0472
R24364 GND.n7827 GND.n2045 13.0472
R24365 GND.n7792 GND.n2091 13.0472
R24366 GND.n7766 GND.n2316 13.0472
R24367 GND.n5759 GND.n3915 13.0472
R24368 GND.n5863 GND.n4019 13.0472
R24369 GND.n7600 GND.n4057 13.0472
R24370 GND.n5966 GND.n4124 13.0472
R24371 GND.n7545 GND.n4162 13.0472
R24372 GND.n6069 GND.n5559 13.0472
R24373 GND.n7490 GND.n4265 13.0472
R24374 GND.n7435 GND.n4369 13.0472
R24375 GND.n7401 GND.n4447 13.0472
R24376 GND.n7379 GND.n4475 13.0472
R24377 GND.n7344 GND.n4521 13.0472
R24378 GND.n7318 GND.n4558 13.0472
R24379 GND.n7283 GND.n4607 13.0472
R24380 GND.n7270 GND.t149 13.0472
R24381 GND.n7257 GND.n4689 13.0472
R24382 GND.t3 GND.n7792 12.721
R24383 GND.t5 GND.n4475 12.721
R24384 GND.n3004 GND.n2863 12.3949
R24385 GND.n3005 GND.n2862 12.3949
R24386 GND.n3018 GND.n3017 12.3949
R24387 GND.n3027 GND.n2848 12.3949
R24388 GND.n2850 GND.n2840 12.3949
R24389 GND.n3036 GND.n3035 12.3949
R24390 GND.n3045 GND.n2834 12.3949
R24391 GND.n2825 GND.n2813 12.3949
R24392 GND.n3071 GND.n3070 12.3949
R24393 GND.n2816 GND.n2806 12.3949
R24394 GND.n3082 GND.n3081 12.3949
R24395 GND.n3097 GND.n2795 12.3949
R24396 GND.n2797 GND.n2785 12.3949
R24397 GND.n3108 GND.n3107 12.3949
R24398 GND.n2787 GND.n2777 12.3949
R24399 GND.n3119 GND.n3118 12.3949
R24400 GND.n3135 GND.n2765 12.3949
R24401 GND.n3122 GND.n2768 12.3949
R24402 GND.n3146 GND.n3145 12.3949
R24403 GND.n2757 GND.n2749 12.3949
R24404 GND.n3158 GND.n3156 12.3949
R24405 GND.n3173 GND.n2738 12.3949
R24406 GND.n2740 GND.n2728 12.3949
R24407 GND.n3184 GND.n3183 12.3949
R24408 GND.n2730 GND.n2721 12.3949
R24409 GND.n3195 GND.n3194 12.3949
R24410 GND.n3210 GND.n2709 12.3949
R24411 GND.n2711 GND.n2698 12.3949
R24412 GND.n3221 GND.n3220 12.3949
R24413 GND.n2701 GND.n2691 12.3949
R24414 GND.n3232 GND.n3231 12.3949
R24415 GND.n3247 GND.n2680 12.3949
R24416 GND.n2682 GND.n2670 12.3949
R24417 GND.n3258 GND.n3257 12.3949
R24418 GND.n2672 GND.n2662 12.3949
R24419 GND.n3269 GND.n3268 12.3949
R24420 GND.n3284 GND.n2650 12.3949
R24421 GND.n2653 GND.n2640 12.3949
R24422 GND.n3296 GND.n3295 12.3949
R24423 GND.n2642 GND.n2633 12.3949
R24424 GND.n3320 GND.n2622 12.3949
R24425 GND.n2624 GND.n2615 12.3949
R24426 GND.n3328 GND.n3327 12.3949
R24427 GND.n2618 GND.n2610 12.3949
R24428 GND.n3542 GND.n3541 12.3949
R24429 GND.n8123 GND.n1533 12.3949
R24430 GND.n2600 GND.n1535 12.3949
R24431 GND.n3556 GND.n2599 12.3949
R24432 GND.n3559 GND.n2596 12.3949
R24433 GND.n8116 GND.n1552 12.3949
R24434 GND.n2588 GND.n1555 12.3949
R24435 GND.n3570 GND.n2587 12.3949
R24436 GND.n3575 GND.n2583 12.3949
R24437 GND.n3572 GND.n2586 12.3949
R24438 GND.n3585 GND.n2572 12.3949
R24439 GND.n2577 GND.n2573 12.3949
R24440 GND.n3595 GND.n2565 12.3949
R24441 GND.n3601 GND.n2561 12.3949
R24442 GND.n3598 GND.n2563 12.3949
R24443 GND.n3611 GND.n2550 12.3949
R24444 GND.n2555 GND.n2551 12.3949
R24445 GND.n3621 GND.n2544 12.3949
R24446 GND.n3627 GND.n2540 12.3949
R24447 GND.n3623 GND.n2542 12.3949
R24448 GND.n3637 GND.n2529 12.3949
R24449 GND.n2534 GND.n2531 12.3949
R24450 GND.n3647 GND.n2523 12.3949
R24451 GND.n3653 GND.n2518 12.3949
R24452 GND.n3650 GND.n2520 12.3949
R24453 GND.n3663 GND.n2508 12.3949
R24454 GND.n2512 GND.n2509 12.3949
R24455 GND.n3673 GND.n2502 12.3949
R24456 GND.n3678 GND.n2496 12.3949
R24457 GND.n3688 GND.n2485 12.3949
R24458 GND.n2490 GND.n2486 12.3949
R24459 GND.n3698 GND.n2478 12.3949
R24460 GND.n3704 GND.n2474 12.3949
R24461 GND.n3701 GND.n2476 12.3949
R24462 GND.n3714 GND.n2463 12.3949
R24463 GND.n2468 GND.n2464 12.3949
R24464 GND.n3724 GND.n2457 12.3949
R24465 GND.n3730 GND.n2453 12.3949
R24466 GND.n3726 GND.n2455 12.3949
R24467 GND.n3740 GND.n2444 12.3949
R24468 GND.n3474 GND.n3473 12.3949
R24469 GND.n3750 GND.n2438 12.3949
R24470 GND.n3756 GND.n2433 12.3949
R24471 GND.n3753 GND.n2435 12.3949
R24472 GND.n3766 GND.n2423 12.3949
R24473 GND.n2427 GND.n2424 12.3949
R24474 GND.n3776 GND.n2417 12.3949
R24475 GND.n3781 GND.n2411 12.3949
R24476 GND.n3778 GND.n2414 12.3949
R24477 GND.n3791 GND.n2400 12.3949
R24478 GND.n2405 GND.n2401 12.3949
R24479 GND.n3801 GND.n2393 12.3949
R24480 GND.n3807 GND.n2389 12.3949
R24481 GND.n3804 GND.n2391 12.3949
R24482 GND.n3817 GND.n2378 12.3949
R24483 GND.n2383 GND.n2379 12.3949
R24484 GND.n3828 GND.n2372 12.3949
R24485 GND.n3834 GND.n2368 12.3949
R24486 GND.n3830 GND.n2370 12.3949
R24487 GND.n3843 GND.n2362 12.3949
R24488 GND.n8026 GND.n1676 12.3949
R24489 GND.n7760 GND.n7759 12.3949
R24490 GND.n7408 GND.n7407 12.3949
R24491 GND.n6416 GND.n4882 12.3949
R24492 GND.n7091 GND.n4885 12.3949
R24493 GND.n7084 GND.n7083 12.3949
R24494 GND.n4905 GND.n4896 12.3949
R24495 GND.n7077 GND.n4906 12.3949
R24496 GND.n7076 GND.n4909 12.3949
R24497 GND.n6473 GND.n6472 12.3949
R24498 GND.n7070 GND.n4926 12.3949
R24499 GND.n6479 GND.n4935 12.3949
R24500 GND.n7064 GND.n4938 12.3949
R24501 GND.n6487 GND.n4946 12.3949
R24502 GND.n7058 GND.n4949 12.3949
R24503 GND.n6493 GND.n4956 12.3949
R24504 GND.n7052 GND.n4959 12.3949
R24505 GND.n6501 GND.n4967 12.3949
R24506 GND.n7046 GND.n4970 12.3949
R24507 GND.n6507 GND.n4977 12.3949
R24508 GND.n7040 GND.n4980 12.3949
R24509 GND.n6516 GND.n4988 12.3949
R24510 GND.n7034 GND.n4991 12.3949
R24511 GND.n6676 GND.n6675 12.3949
R24512 GND.n7028 GND.n5000 12.3949
R24513 GND.n6669 GND.n5008 12.3949
R24514 GND.n7022 GND.n5011 12.3949
R24515 GND.n6663 GND.n5018 12.3949
R24516 GND.n7016 GND.n5021 12.3949
R24517 GND.n6657 GND.n5029 12.3949
R24518 GND.n7010 GND.n5032 12.3949
R24519 GND.n6651 GND.n5039 12.3949
R24520 GND.n7004 GND.n5042 12.3949
R24521 GND.n6645 GND.n5050 12.3949
R24522 GND.n6998 GND.n5053 12.3949
R24523 GND.n6992 GND.n5063 12.3949
R24524 GND.n6633 GND.n5071 12.3949
R24525 GND.n6986 GND.n5074 12.3949
R24526 GND.n6627 GND.n5081 12.3949
R24527 GND.n6980 GND.n5084 12.3949
R24528 GND.n6621 GND.n5092 12.3949
R24529 GND.n6974 GND.n5095 12.3949
R24530 GND.n6615 GND.n5102 12.3949
R24531 GND.n6968 GND.n5105 12.3949
R24532 GND.n6609 GND.n5113 12.3949
R24533 GND.n6962 GND.n5116 12.3949
R24534 GND.n6603 GND.n5123 12.3949
R24535 GND.n6956 GND.n5126 12.3949
R24536 GND.n6597 GND.n5134 12.3949
R24537 GND.n6950 GND.n5137 12.3949
R24538 GND.n6591 GND.n5144 12.3949
R24539 GND.n6944 GND.n5147 12.3949
R24540 GND.n6585 GND.n5155 12.3949
R24541 GND.n6938 GND.n5158 12.3949
R24542 GND.n6579 GND.n5165 12.3949
R24543 GND.n6932 GND.n5168 12.3949
R24544 GND.n6754 GND.n6753 12.3949
R24545 GND.n6926 GND.n5177 12.3949
R24546 GND.n6769 GND.n5184 12.3949
R24547 GND.n6920 GND.n5187 12.3949
R24548 GND.n6916 GND.n6915 12.3949
R24549 GND.n5286 GND.n5192 12.3949
R24550 GND.n6779 GND.n108 12.3949
R24551 GND.n10310 GND.n110 12.3949
R24552 GND.n6788 GND.n6787 12.3949
R24553 GND.n6902 GND.n5269 12.3949
R24554 GND.n6901 GND.n127 12.3949
R24555 GND.n10303 GND.n130 12.3949
R24556 GND.n10297 GND.n142 12.3949
R24557 GND.n6889 GND.n149 12.3949
R24558 GND.n10291 GND.n152 12.3949
R24559 GND.n6883 GND.n159 12.3949
R24560 GND.n10285 GND.n162 12.3949
R24561 GND.n6877 GND.n170 12.3949
R24562 GND.n10279 GND.n173 12.3949
R24563 GND.n6871 GND.n180 12.3949
R24564 GND.n10273 GND.n183 12.3949
R24565 GND.n6865 GND.n191 12.3949
R24566 GND.n10267 GND.n194 12.3949
R24567 GND.n6859 GND.n201 12.3949
R24568 GND.n10261 GND.n204 12.3949
R24569 GND.n6853 GND.n212 12.3949
R24570 GND.n10255 GND.n215 12.3949
R24571 GND.n6847 GND.n222 12.3949
R24572 GND.n10249 GND.n225 12.3949
R24573 GND.n6841 GND.n233 12.3949
R24574 GND.n10243 GND.n236 12.3949
R24575 GND.n6835 GND.n243 12.3949
R24576 GND.n10237 GND.n246 12.3949
R24577 GND.n9727 GND.n9726 12.3949
R24578 GND.n10231 GND.n256 12.3949
R24579 GND.n9735 GND.n263 12.3949
R24580 GND.n10225 GND.n266 12.3949
R24581 GND.n9742 GND.n274 12.3949
R24582 GND.n10219 GND.n277 12.3949
R24583 GND.n9750 GND.n284 12.3949
R24584 GND.n10213 GND.n287 12.3949
R24585 GND.n9757 GND.n295 12.3949
R24586 GND.n10207 GND.n298 12.3949
R24587 GND.n9765 GND.n305 12.3949
R24588 GND.n10201 GND.n308 12.3949
R24589 GND.n10195 GND.n319 12.3949
R24590 GND.n9780 GND.n326 12.3949
R24591 GND.n10189 GND.n329 12.3949
R24592 GND.n9787 GND.n337 12.3949
R24593 GND.n10183 GND.n340 12.3949
R24594 GND.n10104 GND.n347 12.3949
R24595 GND.n10177 GND.n350 12.3949
R24596 GND.n1860 GND.n1859 11.8308
R24597 GND.n1823 GND.n1822 11.8308
R24598 GND.n5394 GND.n5393 11.8308
R24599 GND.n5460 GND.n5456 11.8308
R24600 GND.n10033 GND.n9845 11.8308
R24601 GND.n9971 GND.n9857 11.8308
R24602 GND.n8292 GND.n8291 11.8308
R24603 GND.n8243 GND.n8242 11.8308
R24604 GND.n7903 GND.n1949 11.7425
R24605 GND.n2202 GND.n2201 11.7425
R24606 GND.n7842 GND.n7841 11.7425
R24607 GND.n2107 GND.n2099 11.7425
R24608 GND.n7773 GND.n2304 11.7425
R24609 GND.n5649 GND.n3925 11.7425
R24610 GND.n7662 GND.n3943 11.7425
R24611 GND.n5618 GND.n4029 11.7425
R24612 GND.n7607 GND.n4047 11.7425
R24613 GND.n5587 GND.n4134 11.7425
R24614 GND.n7552 GND.n4152 11.7425
R24615 GND.n5554 GND.n4237 11.7425
R24616 GND.n7497 GND.n4255 11.7425
R24617 GND.n5522 GND.n4341 11.7425
R24618 GND.n7442 GND.n4359 11.7425
R24619 GND.n7394 GND.n7393 11.7425
R24620 GND.n7387 GND.n7386 11.7425
R24621 GND.n7325 GND.n4546 11.7425
R24622 GND.n4679 GND.n4614 11.7425
R24623 GND.n4756 GND.n4733 11.6369
R24624 GND.t97 GND.n7883 11.4164
R24625 GND.n7835 GND.t17 11.4164
R24626 GND.n5602 GND.t4 11.4164
R24627 GND.n7533 GND.t10 11.4164
R24628 GND.n4537 GND.t6 11.4164
R24629 GND.n7284 GND.t26 11.4164
R24630 GND.n5798 GND.t270 11.0902
R24631 GND.t1 GND.n4009 11.0902
R24632 GND.t13 GND.n4057 11.0902
R24633 GND.n5952 GND.t268 11.0902
R24634 GND.t268 GND.n4122 11.0902
R24635 GND.n6013 GND.t11 11.0902
R24636 GND.t11 GND.n4174 11.0902
R24637 GND.n5559 GND.t18 11.0902
R24638 GND.n5548 GND.t272 11.0902
R24639 GND.t15 GND.n4331 11.0902
R24640 GND.n3060 GND.t187 10.764
R24641 GND.t165 GND.n2499 10.764
R24642 GND.n3740 GND.t157 10.764
R24643 GND.n7028 GND.t171 10.764
R24644 GND.t155 GND.n5060 10.764
R24645 GND.n9772 GND.t181 10.764
R24646 GND.n7977 GND.n1768 10.6672
R24647 GND.n7187 GND.n7186 10.6672
R24648 GND.n4832 GND.n4829 10.6151
R24649 GND.n4829 GND.n4828 10.6151
R24650 GND.n4825 GND.n4824 10.6151
R24651 GND.n4824 GND.n4821 10.6151
R24652 GND.n4821 GND.n4820 10.6151
R24653 GND.n4820 GND.n4817 10.6151
R24654 GND.n4817 GND.n4816 10.6151
R24655 GND.n4816 GND.n4813 10.6151
R24656 GND.n4813 GND.n4812 10.6151
R24657 GND.n4812 GND.n4809 10.6151
R24658 GND.n4809 GND.n4808 10.6151
R24659 GND.n4808 GND.n4805 10.6151
R24660 GND.n4805 GND.n4804 10.6151
R24661 GND.n4804 GND.n4801 10.6151
R24662 GND.n4801 GND.n4800 10.6151
R24663 GND.n4800 GND.n4797 10.6151
R24664 GND.n4797 GND.n4796 10.6151
R24665 GND.n4796 GND.n4793 10.6151
R24666 GND.n4793 GND.n4792 10.6151
R24667 GND.n4792 GND.n4789 10.6151
R24668 GND.n4789 GND.n4788 10.6151
R24669 GND.n4788 GND.n4785 10.6151
R24670 GND.n4785 GND.n4784 10.6151
R24671 GND.n4784 GND.n4781 10.6151
R24672 GND.n4781 GND.n4780 10.6151
R24673 GND.n4780 GND.n4777 10.6151
R24674 GND.n4777 GND.n4776 10.6151
R24675 GND.n2183 GND.n2182 10.6151
R24676 GND.n2184 GND.n2183 10.6151
R24677 GND.n2184 GND.n2120 10.6151
R24678 GND.n2193 GND.n2120 10.6151
R24679 GND.n2194 GND.n2193 10.6151
R24680 GND.n2197 GND.n2194 10.6151
R24681 GND.n2198 GND.n2197 10.6151
R24682 GND.n2199 GND.n2198 10.6151
R24683 GND.n2204 GND.n2199 10.6151
R24684 GND.n2205 GND.n2204 10.6151
R24685 GND.n2207 GND.n2205 10.6151
R24686 GND.n2208 GND.n2207 10.6151
R24687 GND.n2209 GND.n2208 10.6151
R24688 GND.n2209 GND.n2119 10.6151
R24689 GND.n2217 GND.n2119 10.6151
R24690 GND.n2218 GND.n2217 10.6151
R24691 GND.n2220 GND.n2218 10.6151
R24692 GND.n2221 GND.n2220 10.6151
R24693 GND.n2222 GND.n2221 10.6151
R24694 GND.n2222 GND.n2118 10.6151
R24695 GND.n2230 GND.n2118 10.6151
R24696 GND.n2231 GND.n2230 10.6151
R24697 GND.n2233 GND.n2231 10.6151
R24698 GND.n2234 GND.n2233 10.6151
R24699 GND.n2235 GND.n2234 10.6151
R24700 GND.n2235 GND.n2117 10.6151
R24701 GND.n2243 GND.n2117 10.6151
R24702 GND.n2244 GND.n2243 10.6151
R24703 GND.n2246 GND.n2244 10.6151
R24704 GND.n2247 GND.n2246 10.6151
R24705 GND.n2248 GND.n2247 10.6151
R24706 GND.n2248 GND.n2116 10.6151
R24707 GND.n2255 GND.n2116 10.6151
R24708 GND.n2256 GND.n2255 10.6151
R24709 GND.n2258 GND.n2256 10.6151
R24710 GND.n2259 GND.n2258 10.6151
R24711 GND.n2260 GND.n2259 10.6151
R24712 GND.n2260 GND.n2115 10.6151
R24713 GND.n2268 GND.n2115 10.6151
R24714 GND.n2269 GND.n2268 10.6151
R24715 GND.n2271 GND.n2269 10.6151
R24716 GND.n2272 GND.n2271 10.6151
R24717 GND.n2273 GND.n2272 10.6151
R24718 GND.n2273 GND.n2114 10.6151
R24719 GND.n2281 GND.n2114 10.6151
R24720 GND.n2282 GND.n2281 10.6151
R24721 GND.n2284 GND.n2282 10.6151
R24722 GND.n2285 GND.n2284 10.6151
R24723 GND.n2286 GND.n2285 10.6151
R24724 GND.n2286 GND.n2113 10.6151
R24725 GND.n2294 GND.n2113 10.6151
R24726 GND.n2295 GND.n2294 10.6151
R24727 GND.n2297 GND.n2295 10.6151
R24728 GND.n2298 GND.n2297 10.6151
R24729 GND.n2300 GND.n2298 10.6151
R24730 GND.n2301 GND.n2300 10.6151
R24731 GND.n7777 GND.n2301 10.6151
R24732 GND.n7777 GND.n7776 10.6151
R24733 GND.n7776 GND.n7775 10.6151
R24734 GND.n7775 GND.n2302 10.6151
R24735 GND.n5697 GND.n2302 10.6151
R24736 GND.n5698 GND.n5697 10.6151
R24737 GND.n5701 GND.n5698 10.6151
R24738 GND.n5701 GND.n5700 10.6151
R24739 GND.n5700 GND.n5699 10.6151
R24740 GND.n5699 GND.n5688 10.6151
R24741 GND.n5715 GND.n5688 10.6151
R24742 GND.n5716 GND.n5715 10.6151
R24743 GND.n5719 GND.n5716 10.6151
R24744 GND.n5719 GND.n5718 10.6151
R24745 GND.n5718 GND.n5717 10.6151
R24746 GND.n5717 GND.n5662 10.6151
R24747 GND.n5733 GND.n5662 10.6151
R24748 GND.n5734 GND.n5733 10.6151
R24749 GND.n5743 GND.n5734 10.6151
R24750 GND.n5743 GND.n5742 10.6151
R24751 GND.n5742 GND.n5741 10.6151
R24752 GND.n5741 GND.n5739 10.6151
R24753 GND.n5739 GND.n5738 10.6151
R24754 GND.n5738 GND.n5735 10.6151
R24755 GND.n5735 GND.n3940 10.6151
R24756 GND.n7666 GND.n3940 10.6151
R24757 GND.n7666 GND.n7665 10.6151
R24758 GND.n7665 GND.n7664 10.6151
R24759 GND.n7664 GND.n3941 10.6151
R24760 GND.n5801 GND.n3941 10.6151
R24761 GND.n5802 GND.n5801 10.6151
R24762 GND.n5805 GND.n5802 10.6151
R24763 GND.n5805 GND.n5804 10.6151
R24764 GND.n5804 GND.n5803 10.6151
R24765 GND.n5803 GND.n5641 10.6151
R24766 GND.n5819 GND.n5641 10.6151
R24767 GND.n5820 GND.n5819 10.6151
R24768 GND.n5823 GND.n5820 10.6151
R24769 GND.n5823 GND.n5822 10.6151
R24770 GND.n5822 GND.n5821 10.6151
R24771 GND.n5821 GND.n5631 10.6151
R24772 GND.n5837 GND.n5631 10.6151
R24773 GND.n5838 GND.n5837 10.6151
R24774 GND.n5847 GND.n5838 10.6151
R24775 GND.n5847 GND.n5846 10.6151
R24776 GND.n5846 GND.n5845 10.6151
R24777 GND.n5845 GND.n5843 10.6151
R24778 GND.n5843 GND.n5842 10.6151
R24779 GND.n5842 GND.n5839 10.6151
R24780 GND.n5839 GND.n4044 10.6151
R24781 GND.n7611 GND.n4044 10.6151
R24782 GND.n7611 GND.n7610 10.6151
R24783 GND.n7610 GND.n7609 10.6151
R24784 GND.n7609 GND.n4045 10.6151
R24785 GND.n5904 GND.n4045 10.6151
R24786 GND.n5905 GND.n5904 10.6151
R24787 GND.n5908 GND.n5905 10.6151
R24788 GND.n5908 GND.n5907 10.6151
R24789 GND.n5907 GND.n5906 10.6151
R24790 GND.n5906 GND.n5610 10.6151
R24791 GND.n5922 GND.n5610 10.6151
R24792 GND.n5923 GND.n5922 10.6151
R24793 GND.n5926 GND.n5923 10.6151
R24794 GND.n5926 GND.n5925 10.6151
R24795 GND.n5925 GND.n5924 10.6151
R24796 GND.n5924 GND.n5600 10.6151
R24797 GND.n5940 GND.n5600 10.6151
R24798 GND.n5941 GND.n5940 10.6151
R24799 GND.n5950 GND.n5941 10.6151
R24800 GND.n5950 GND.n5949 10.6151
R24801 GND.n5949 GND.n5948 10.6151
R24802 GND.n5948 GND.n5946 10.6151
R24803 GND.n5946 GND.n5945 10.6151
R24804 GND.n5945 GND.n5942 10.6151
R24805 GND.n5942 GND.n4149 10.6151
R24806 GND.n7556 GND.n4149 10.6151
R24807 GND.n7556 GND.n7555 10.6151
R24808 GND.n7555 GND.n7554 10.6151
R24809 GND.n7554 GND.n4150 10.6151
R24810 GND.n6007 GND.n4150 10.6151
R24811 GND.n6008 GND.n6007 10.6151
R24812 GND.n6011 GND.n6008 10.6151
R24813 GND.n6011 GND.n6010 10.6151
R24814 GND.n6010 GND.n6009 10.6151
R24815 GND.n6009 GND.n5579 10.6151
R24816 GND.n6025 GND.n5579 10.6151
R24817 GND.n6026 GND.n6025 10.6151
R24818 GND.n6029 GND.n6026 10.6151
R24819 GND.n6029 GND.n6028 10.6151
R24820 GND.n6028 GND.n6027 10.6151
R24821 GND.n6027 GND.n5568 10.6151
R24822 GND.n6043 GND.n5568 10.6151
R24823 GND.n6044 GND.n6043 10.6151
R24824 GND.n6053 GND.n6044 10.6151
R24825 GND.n6053 GND.n6052 10.6151
R24826 GND.n6052 GND.n6051 10.6151
R24827 GND.n6051 GND.n6049 10.6151
R24828 GND.n6049 GND.n6048 10.6151
R24829 GND.n6048 GND.n6045 10.6151
R24830 GND.n6045 GND.n4252 10.6151
R24831 GND.n7501 GND.n4252 10.6151
R24832 GND.n7501 GND.n7500 10.6151
R24833 GND.n7500 GND.n7499 10.6151
R24834 GND.n7499 GND.n4253 10.6151
R24835 GND.n6110 GND.n4253 10.6151
R24836 GND.n6111 GND.n6110 10.6151
R24837 GND.n6114 GND.n6111 10.6151
R24838 GND.n6114 GND.n6113 10.6151
R24839 GND.n6113 GND.n6112 10.6151
R24840 GND.n6112 GND.n5545 10.6151
R24841 GND.n6128 GND.n5545 10.6151
R24842 GND.n6129 GND.n6128 10.6151
R24843 GND.n6132 GND.n6129 10.6151
R24844 GND.n6132 GND.n6131 10.6151
R24845 GND.n6131 GND.n6130 10.6151
R24846 GND.n6130 GND.n5535 10.6151
R24847 GND.n6146 GND.n5535 10.6151
R24848 GND.n6147 GND.n6146 10.6151
R24849 GND.n6156 GND.n6147 10.6151
R24850 GND.n6156 GND.n6155 10.6151
R24851 GND.n6155 GND.n6154 10.6151
R24852 GND.n6154 GND.n6152 10.6151
R24853 GND.n6152 GND.n6151 10.6151
R24854 GND.n6151 GND.n6148 10.6151
R24855 GND.n6148 GND.n4356 10.6151
R24856 GND.n7446 GND.n4356 10.6151
R24857 GND.n7446 GND.n7445 10.6151
R24858 GND.n7445 GND.n7444 10.6151
R24859 GND.n7444 GND.n4357 10.6151
R24860 GND.n5517 GND.n4357 10.6151
R24861 GND.n5518 GND.n5517 10.6151
R24862 GND.n5518 GND.n5516 10.6151
R24863 GND.n6212 GND.n5516 10.6151
R24864 GND.n6213 GND.n6212 10.6151
R24865 GND.n6218 GND.n6213 10.6151
R24866 GND.n6218 GND.n6217 10.6151
R24867 GND.n6217 GND.n6216 10.6151
R24868 GND.n6216 GND.n6214 10.6151
R24869 GND.n6214 GND.n5507 10.6151
R24870 GND.n6231 GND.n5507 10.6151
R24871 GND.n6232 GND.n6231 10.6151
R24872 GND.n6233 GND.n6232 10.6151
R24873 GND.n6236 GND.n6233 10.6151
R24874 GND.n6237 GND.n6236 10.6151
R24875 GND.n6300 GND.n6237 10.6151
R24876 GND.n6300 GND.n6299 10.6151
R24877 GND.n6299 GND.n6298 10.6151
R24878 GND.n6298 GND.n6297 10.6151
R24879 GND.n6297 GND.n6295 10.6151
R24880 GND.n6295 GND.n6294 10.6151
R24881 GND.n6294 GND.n6238 10.6151
R24882 GND.n6287 GND.n6238 10.6151
R24883 GND.n6287 GND.n6286 10.6151
R24884 GND.n6286 GND.n6285 10.6151
R24885 GND.n6285 GND.n6283 10.6151
R24886 GND.n6283 GND.n6282 10.6151
R24887 GND.n6282 GND.n6239 10.6151
R24888 GND.n6274 GND.n6239 10.6151
R24889 GND.n6274 GND.n6273 10.6151
R24890 GND.n6273 GND.n6272 10.6151
R24891 GND.n6272 GND.n6270 10.6151
R24892 GND.n6270 GND.n6269 10.6151
R24893 GND.n6269 GND.n6240 10.6151
R24894 GND.n6261 GND.n6240 10.6151
R24895 GND.n6261 GND.n6260 10.6151
R24896 GND.n6260 GND.n6259 10.6151
R24897 GND.n6259 GND.n6257 10.6151
R24898 GND.n6257 GND.n6256 10.6151
R24899 GND.n6256 GND.n6241 10.6151
R24900 GND.n6248 GND.n6241 10.6151
R24901 GND.n6248 GND.n6247 10.6151
R24902 GND.n6247 GND.n6246 10.6151
R24903 GND.n6246 GND.n6244 10.6151
R24904 GND.n6244 GND.n6243 10.6151
R24905 GND.n6243 GND.n4543 10.6151
R24906 GND.n7329 GND.n4543 10.6151
R24907 GND.n7329 GND.n7328 10.6151
R24908 GND.n7328 GND.n7327 10.6151
R24909 GND.n7327 GND.n4544 10.6151
R24910 GND.n4629 GND.n4544 10.6151
R24911 GND.n4630 GND.n4629 10.6151
R24912 GND.n4630 GND.n4628 10.6151
R24913 GND.n4638 GND.n4628 10.6151
R24914 GND.n4639 GND.n4638 10.6151
R24915 GND.n4641 GND.n4639 10.6151
R24916 GND.n4642 GND.n4641 10.6151
R24917 GND.n4643 GND.n4642 10.6151
R24918 GND.n4643 GND.n4627 10.6151
R24919 GND.n4651 GND.n4627 10.6151
R24920 GND.n4652 GND.n4651 10.6151
R24921 GND.n4654 GND.n4652 10.6151
R24922 GND.n4655 GND.n4654 10.6151
R24923 GND.n4656 GND.n4655 10.6151
R24924 GND.n4656 GND.n4626 10.6151
R24925 GND.n4664 GND.n4626 10.6151
R24926 GND.n4665 GND.n4664 10.6151
R24927 GND.n4668 GND.n4665 10.6151
R24928 GND.n4669 GND.n4668 10.6151
R24929 GND.n4671 GND.n4669 10.6151
R24930 GND.n4672 GND.n4671 10.6151
R24931 GND.n7268 GND.n4672 10.6151
R24932 GND.n7268 GND.n7267 10.6151
R24933 GND.n7267 GND.n7266 10.6151
R24934 GND.n7266 GND.n4673 10.6151
R24935 GND.n4765 GND.n4673 10.6151
R24936 GND.n4766 GND.n4765 10.6151
R24937 GND.n4767 GND.n4766 10.6151
R24938 GND.n4767 GND.n4763 10.6151
R24939 GND.n2126 GND.n1871 10.6151
R24940 GND.n2127 GND.n2126 10.6151
R24941 GND.n2131 GND.n2130 10.6151
R24942 GND.n2134 GND.n2131 10.6151
R24943 GND.n2135 GND.n2134 10.6151
R24944 GND.n2138 GND.n2135 10.6151
R24945 GND.n2139 GND.n2138 10.6151
R24946 GND.n2142 GND.n2139 10.6151
R24947 GND.n2143 GND.n2142 10.6151
R24948 GND.n2146 GND.n2143 10.6151
R24949 GND.n2147 GND.n2146 10.6151
R24950 GND.n2150 GND.n2147 10.6151
R24951 GND.n2151 GND.n2150 10.6151
R24952 GND.n2154 GND.n2151 10.6151
R24953 GND.n2155 GND.n2154 10.6151
R24954 GND.n2158 GND.n2155 10.6151
R24955 GND.n2159 GND.n2158 10.6151
R24956 GND.n2162 GND.n2159 10.6151
R24957 GND.n2163 GND.n2162 10.6151
R24958 GND.n2166 GND.n2163 10.6151
R24959 GND.n2167 GND.n2166 10.6151
R24960 GND.n2170 GND.n2167 10.6151
R24961 GND.n2171 GND.n2170 10.6151
R24962 GND.n2174 GND.n2171 10.6151
R24963 GND.n2175 GND.n2174 10.6151
R24964 GND.n2178 GND.n2175 10.6151
R24965 GND.n2179 GND.n2178 10.6151
R24966 GND.n7969 GND.n7968 10.6151
R24967 GND.n7968 GND.n7967 10.6151
R24968 GND.n7967 GND.n7966 10.6151
R24969 GND.n7966 GND.n7964 10.6151
R24970 GND.n7964 GND.n7961 10.6151
R24971 GND.n7961 GND.n7960 10.6151
R24972 GND.n7960 GND.n7957 10.6151
R24973 GND.n7957 GND.n7956 10.6151
R24974 GND.n7956 GND.n7953 10.6151
R24975 GND.n7953 GND.n7952 10.6151
R24976 GND.n7952 GND.n7949 10.6151
R24977 GND.n7949 GND.n7948 10.6151
R24978 GND.n7948 GND.n7945 10.6151
R24979 GND.n7945 GND.n7944 10.6151
R24980 GND.n7944 GND.n7941 10.6151
R24981 GND.n7941 GND.n7940 10.6151
R24982 GND.n7940 GND.n7937 10.6151
R24983 GND.n7937 GND.n7936 10.6151
R24984 GND.n7936 GND.n7933 10.6151
R24985 GND.n7933 GND.n7932 10.6151
R24986 GND.n7932 GND.n7929 10.6151
R24987 GND.n7929 GND.n7928 10.6151
R24988 GND.n7928 GND.n7925 10.6151
R24989 GND.n7925 GND.n7924 10.6151
R24990 GND.n7924 GND.n7921 10.6151
R24991 GND.n7919 GND.n1874 10.6151
R24992 GND.n7975 GND.n1874 10.6151
R24993 GND.n7247 GND.n7246 10.6151
R24994 GND.n7246 GND.n7245 10.6151
R24995 GND.n7245 GND.n7242 10.6151
R24996 GND.n7242 GND.n7241 10.6151
R24997 GND.n7241 GND.n7238 10.6151
R24998 GND.n7238 GND.n7237 10.6151
R24999 GND.n7237 GND.n7234 10.6151
R25000 GND.n7234 GND.n7233 10.6151
R25001 GND.n7233 GND.n7230 10.6151
R25002 GND.n7230 GND.n7229 10.6151
R25003 GND.n7229 GND.n7226 10.6151
R25004 GND.n7226 GND.n7225 10.6151
R25005 GND.n7225 GND.n7222 10.6151
R25006 GND.n7222 GND.n7221 10.6151
R25007 GND.n7221 GND.n7218 10.6151
R25008 GND.n7218 GND.n7217 10.6151
R25009 GND.n7217 GND.n7214 10.6151
R25010 GND.n7214 GND.n7213 10.6151
R25011 GND.n7213 GND.n7210 10.6151
R25012 GND.n7210 GND.n7209 10.6151
R25013 GND.n7209 GND.n7206 10.6151
R25014 GND.n7206 GND.n7205 10.6151
R25015 GND.n7205 GND.n7202 10.6151
R25016 GND.n7202 GND.n7201 10.6151
R25017 GND.n7201 GND.n7198 10.6151
R25018 GND.n7196 GND.n7193 10.6151
R25019 GND.n7193 GND.n7192 10.6151
R25020 GND.n7914 GND.n7913 10.6151
R25021 GND.n7913 GND.n1934 10.6151
R25022 GND.n2188 GND.n1934 10.6151
R25023 GND.n2188 GND.n1952 10.6151
R25024 GND.n7901 GND.n1952 10.6151
R25025 GND.n7901 GND.n7900 10.6151
R25026 GND.n7900 GND.n7899 10.6151
R25027 GND.n7899 GND.n1953 10.6151
R25028 GND.n1968 GND.n1953 10.6151
R25029 GND.n7888 GND.n1968 10.6151
R25030 GND.n7888 GND.n7887 10.6151
R25031 GND.n7887 GND.n7886 10.6151
R25032 GND.n7886 GND.n1969 10.6151
R25033 GND.n2212 GND.n1969 10.6151
R25034 GND.n2212 GND.n1986 10.6151
R25035 GND.n7874 GND.n1986 10.6151
R25036 GND.n7874 GND.n7873 10.6151
R25037 GND.n7873 GND.n7872 10.6151
R25038 GND.n7872 GND.n1987 10.6151
R25039 GND.n2225 GND.n1987 10.6151
R25040 GND.n2225 GND.n2004 10.6151
R25041 GND.n7860 GND.n2004 10.6151
R25042 GND.n7860 GND.n7859 10.6151
R25043 GND.n7859 GND.n7858 10.6151
R25044 GND.n7858 GND.n2005 10.6151
R25045 GND.n2238 GND.n2005 10.6151
R25046 GND.n2238 GND.n2022 10.6151
R25047 GND.n7846 GND.n2022 10.6151
R25048 GND.n7846 GND.n7845 10.6151
R25049 GND.n7845 GND.n7844 10.6151
R25050 GND.n7844 GND.n2023 10.6151
R25051 GND.n2250 GND.n2023 10.6151
R25052 GND.n2250 GND.n2040 10.6151
R25053 GND.n7832 GND.n2040 10.6151
R25054 GND.n7832 GND.n7831 10.6151
R25055 GND.n7831 GND.n7830 10.6151
R25056 GND.n7830 GND.n2041 10.6151
R25057 GND.n2263 GND.n2041 10.6151
R25058 GND.n2263 GND.n2058 10.6151
R25059 GND.n7818 GND.n2058 10.6151
R25060 GND.n7818 GND.n7817 10.6151
R25061 GND.n7817 GND.n7816 10.6151
R25062 GND.n7816 GND.n2059 10.6151
R25063 GND.n2276 GND.n2059 10.6151
R25064 GND.n2276 GND.n2076 10.6151
R25065 GND.n7804 GND.n2076 10.6151
R25066 GND.n7804 GND.n7803 10.6151
R25067 GND.n7803 GND.n7802 10.6151
R25068 GND.n7802 GND.n2077 10.6151
R25069 GND.n2289 GND.n2077 10.6151
R25070 GND.n2289 GND.n2094 10.6151
R25071 GND.n7790 GND.n2094 10.6151
R25072 GND.n7790 GND.n7789 10.6151
R25073 GND.n7789 GND.n7788 10.6151
R25074 GND.n7788 GND.n2095 10.6151
R25075 GND.n2309 GND.n2095 10.6151
R25076 GND.n2310 GND.n2309 10.6151
R25077 GND.n2311 GND.n2310 10.6151
R25078 GND.n7771 GND.n2311 10.6151
R25079 GND.n7771 GND.n7770 10.6151
R25080 GND.n7770 GND.n7769 10.6151
R25081 GND.n7769 GND.n2312 10.6151
R25082 GND.n5693 GND.n2312 10.6151
R25083 GND.n5706 GND.n5693 10.6151
R25084 GND.n5707 GND.n5706 10.6151
R25085 GND.n5710 GND.n5707 10.6151
R25086 GND.n5710 GND.n5709 10.6151
R25087 GND.n5709 GND.n5708 10.6151
R25088 GND.n5708 GND.n5667 10.6151
R25089 GND.n5724 GND.n5667 10.6151
R25090 GND.n5725 GND.n5724 10.6151
R25091 GND.n5728 GND.n5725 10.6151
R25092 GND.n5728 GND.n5727 10.6151
R25093 GND.n5727 GND.n5726 10.6151
R25094 GND.n5726 GND.n5657 10.6151
R25095 GND.n5748 GND.n5657 10.6151
R25096 GND.n5749 GND.n5748 10.6151
R25097 GND.n5756 GND.n5749 10.6151
R25098 GND.n5756 GND.n5755 10.6151
R25099 GND.n5755 GND.n5754 10.6151
R25100 GND.n5754 GND.n5751 10.6151
R25101 GND.n5751 GND.n5750 10.6151
R25102 GND.n5750 GND.n3947 10.6151
R25103 GND.n7660 GND.n3947 10.6151
R25104 GND.n7660 GND.n7659 10.6151
R25105 GND.n7659 GND.n7658 10.6151
R25106 GND.n7658 GND.n3948 10.6151
R25107 GND.n5646 GND.n3948 10.6151
R25108 GND.n5810 GND.n5646 10.6151
R25109 GND.n5811 GND.n5810 10.6151
R25110 GND.n5814 GND.n5811 10.6151
R25111 GND.n5814 GND.n5813 10.6151
R25112 GND.n5813 GND.n5812 10.6151
R25113 GND.n5812 GND.n5636 10.6151
R25114 GND.n5828 GND.n5636 10.6151
R25115 GND.n5829 GND.n5828 10.6151
R25116 GND.n5832 GND.n5829 10.6151
R25117 GND.n5832 GND.n5831 10.6151
R25118 GND.n5831 GND.n5830 10.6151
R25119 GND.n5830 GND.n5626 10.6151
R25120 GND.n5852 GND.n5626 10.6151
R25121 GND.n5853 GND.n5852 10.6151
R25122 GND.n5860 GND.n5853 10.6151
R25123 GND.n5860 GND.n5859 10.6151
R25124 GND.n5859 GND.n5858 10.6151
R25125 GND.n5858 GND.n5855 10.6151
R25126 GND.n5855 GND.n5854 10.6151
R25127 GND.n5854 GND.n4051 10.6151
R25128 GND.n7605 GND.n4051 10.6151
R25129 GND.n7605 GND.n7604 10.6151
R25130 GND.n7604 GND.n7603 10.6151
R25131 GND.n7603 GND.n4052 10.6151
R25132 GND.n5615 GND.n4052 10.6151
R25133 GND.n5913 GND.n5615 10.6151
R25134 GND.n5914 GND.n5913 10.6151
R25135 GND.n5917 GND.n5914 10.6151
R25136 GND.n5917 GND.n5916 10.6151
R25137 GND.n5916 GND.n5915 10.6151
R25138 GND.n5915 GND.n5605 10.6151
R25139 GND.n5931 GND.n5605 10.6151
R25140 GND.n5932 GND.n5931 10.6151
R25141 GND.n5935 GND.n5932 10.6151
R25142 GND.n5935 GND.n5934 10.6151
R25143 GND.n5934 GND.n5933 10.6151
R25144 GND.n5933 GND.n5595 10.6151
R25145 GND.n5955 GND.n5595 10.6151
R25146 GND.n5956 GND.n5955 10.6151
R25147 GND.n5963 GND.n5956 10.6151
R25148 GND.n5963 GND.n5962 10.6151
R25149 GND.n5962 GND.n5961 10.6151
R25150 GND.n5961 GND.n5958 10.6151
R25151 GND.n5958 GND.n5957 10.6151
R25152 GND.n5957 GND.n4156 10.6151
R25153 GND.n7550 GND.n4156 10.6151
R25154 GND.n7550 GND.n7549 10.6151
R25155 GND.n7549 GND.n7548 10.6151
R25156 GND.n7548 GND.n4157 10.6151
R25157 GND.n5584 GND.n4157 10.6151
R25158 GND.n6016 GND.n5584 10.6151
R25159 GND.n6017 GND.n6016 10.6151
R25160 GND.n6020 GND.n6017 10.6151
R25161 GND.n6020 GND.n6019 10.6151
R25162 GND.n6019 GND.n6018 10.6151
R25163 GND.n6018 GND.n5573 10.6151
R25164 GND.n6034 GND.n5573 10.6151
R25165 GND.n6035 GND.n6034 10.6151
R25166 GND.n6038 GND.n6035 10.6151
R25167 GND.n6038 GND.n6037 10.6151
R25168 GND.n6037 GND.n6036 10.6151
R25169 GND.n6036 GND.n5563 10.6151
R25170 GND.n6058 GND.n5563 10.6151
R25171 GND.n6059 GND.n6058 10.6151
R25172 GND.n6066 GND.n6059 10.6151
R25173 GND.n6066 GND.n6065 10.6151
R25174 GND.n6065 GND.n6064 10.6151
R25175 GND.n6064 GND.n6061 10.6151
R25176 GND.n6061 GND.n6060 10.6151
R25177 GND.n6060 GND.n4259 10.6151
R25178 GND.n7495 GND.n4259 10.6151
R25179 GND.n7495 GND.n7494 10.6151
R25180 GND.n7494 GND.n7493 10.6151
R25181 GND.n7493 GND.n4260 10.6151
R25182 GND.n5551 GND.n4260 10.6151
R25183 GND.n6119 GND.n5551 10.6151
R25184 GND.n6120 GND.n6119 10.6151
R25185 GND.n6123 GND.n6120 10.6151
R25186 GND.n6123 GND.n6122 10.6151
R25187 GND.n6122 GND.n6121 10.6151
R25188 GND.n6121 GND.n5540 10.6151
R25189 GND.n6137 GND.n5540 10.6151
R25190 GND.n6138 GND.n6137 10.6151
R25191 GND.n6141 GND.n6138 10.6151
R25192 GND.n6141 GND.n6140 10.6151
R25193 GND.n6140 GND.n6139 10.6151
R25194 GND.n6139 GND.n5530 10.6151
R25195 GND.n6161 GND.n5530 10.6151
R25196 GND.n6162 GND.n6161 10.6151
R25197 GND.n6169 GND.n6162 10.6151
R25198 GND.n6169 GND.n6168 10.6151
R25199 GND.n6168 GND.n6167 10.6151
R25200 GND.n6167 GND.n6164 10.6151
R25201 GND.n6164 GND.n6163 10.6151
R25202 GND.n6163 GND.n4363 10.6151
R25203 GND.n7440 GND.n4363 10.6151
R25204 GND.n7440 GND.n7439 10.6151
R25205 GND.n7439 GND.n7438 10.6151
R25206 GND.n7438 GND.n4364 10.6151
R25207 GND.n6207 GND.n4364 10.6151
R25208 GND.n6207 GND.n6206 10.6151
R25209 GND.n6206 GND.n6205 10.6151
R25210 GND.n6205 GND.n5513 10.6151
R25211 GND.n5513 GND.n5511 10.6151
R25212 GND.n6224 GND.n5511 10.6151
R25213 GND.n6225 GND.n6224 10.6151
R25214 GND.n6226 GND.n6225 10.6151
R25215 GND.n6226 GND.n5502 10.6151
R25216 GND.n6309 GND.n5502 10.6151
R25217 GND.n6309 GND.n6308 10.6151
R25218 GND.n6308 GND.n6307 10.6151
R25219 GND.n6307 GND.n5503 10.6151
R25220 GND.n5504 GND.n5503 10.6151
R25221 GND.n5504 GND.n4452 10.6151
R25222 GND.n7398 GND.n4452 10.6151
R25223 GND.n7398 GND.n7397 10.6151
R25224 GND.n7397 GND.n7396 10.6151
R25225 GND.n7396 GND.n4453 10.6151
R25226 GND.n6289 GND.n4453 10.6151
R25227 GND.n6289 GND.n4470 10.6151
R25228 GND.n7384 GND.n4470 10.6151
R25229 GND.n7384 GND.n7383 10.6151
R25230 GND.n7383 GND.n7382 10.6151
R25231 GND.n7382 GND.n4471 10.6151
R25232 GND.n6277 GND.n4471 10.6151
R25233 GND.n6277 GND.n4488 10.6151
R25234 GND.n7370 GND.n4488 10.6151
R25235 GND.n7370 GND.n7369 10.6151
R25236 GND.n7369 GND.n7368 10.6151
R25237 GND.n7368 GND.n4489 10.6151
R25238 GND.n6264 GND.n4489 10.6151
R25239 GND.n6264 GND.n4506 10.6151
R25240 GND.n7356 GND.n4506 10.6151
R25241 GND.n7356 GND.n7355 10.6151
R25242 GND.n7355 GND.n7354 10.6151
R25243 GND.n7354 GND.n4507 10.6151
R25244 GND.n6251 GND.n4507 10.6151
R25245 GND.n6251 GND.n4524 10.6151
R25246 GND.n7342 GND.n4524 10.6151
R25247 GND.n7342 GND.n7341 10.6151
R25248 GND.n7341 GND.n7340 10.6151
R25249 GND.n7340 GND.n4525 10.6151
R25250 GND.n4551 GND.n4525 10.6151
R25251 GND.n4552 GND.n4551 10.6151
R25252 GND.n4553 GND.n4552 10.6151
R25253 GND.n7323 GND.n4553 10.6151
R25254 GND.n7323 GND.n7322 10.6151
R25255 GND.n7322 GND.n7321 10.6151
R25256 GND.n7321 GND.n4554 10.6151
R25257 GND.n4633 GND.n4554 10.6151
R25258 GND.n4633 GND.n4574 10.6151
R25259 GND.n7309 GND.n4574 10.6151
R25260 GND.n7309 GND.n7308 10.6151
R25261 GND.n7308 GND.n7307 10.6151
R25262 GND.n7307 GND.n4575 10.6151
R25263 GND.n4646 GND.n4575 10.6151
R25264 GND.n4646 GND.n4592 10.6151
R25265 GND.n7295 GND.n4592 10.6151
R25266 GND.n7295 GND.n7294 10.6151
R25267 GND.n7294 GND.n7293 10.6151
R25268 GND.n7293 GND.n4593 10.6151
R25269 GND.n4659 GND.n4593 10.6151
R25270 GND.n4659 GND.n4610 10.6151
R25271 GND.n7281 GND.n4610 10.6151
R25272 GND.n7281 GND.n7280 10.6151
R25273 GND.n7280 GND.n7279 10.6151
R25274 GND.n7279 GND.n4611 10.6151
R25275 GND.n4682 GND.n4611 10.6151
R25276 GND.n4683 GND.n4682 10.6151
R25277 GND.n4684 GND.n4683 10.6151
R25278 GND.n7262 GND.n4684 10.6151
R25279 GND.n7262 GND.n7261 10.6151
R25280 GND.n7261 GND.n7260 10.6151
R25281 GND.n7260 GND.n4685 10.6151
R25282 GND.n4770 GND.n4685 10.6151
R25283 GND.n4770 GND.n4769 10.6151
R25284 GND.n2195 GND.n1949 10.4379
R25285 GND.n2201 GND.n1955 10.4379
R25286 GND.n7841 GND.n2027 10.4379
R25287 GND.n7835 GND.n2035 10.4379
R25288 GND.n2108 GND.n2107 10.4379
R25289 GND.n2304 GND.n2110 10.4379
R25290 GND.n5649 GND.n3933 10.4379
R25291 GND.n3943 GND.n3936 10.4379
R25292 GND.n5618 GND.n4037 10.4379
R25293 GND.n4047 GND.n4040 10.4379
R25294 GND.n5587 GND.n4142 10.4379
R25295 GND.n4152 GND.n4145 10.4379
R25296 GND.n5554 GND.n4245 10.4379
R25297 GND.n4255 GND.n4248 10.4379
R25298 GND.n5522 GND.n4349 10.4379
R25299 GND.n4359 GND.n4352 10.4379
R25300 GND.n7393 GND.n4457 10.4379
R25301 GND.n7387 GND.n4465 10.4379
R25302 GND.n4538 GND.n4537 10.4379
R25303 GND.n4546 GND.n4540 10.4379
R25304 GND.n4680 GND.n4679 10.4379
R25305 GND.n4675 GND.n4623 10.4379
R25306 GND.n8223 GND.n1452 10.2793
R25307 GND.n10077 GND.n9810 10.2793
R25308 GND.n8005 GND.n8004 9.50353
R25309 GND.n7163 GND.n7162 9.50353
R25310 GND.n9912 GND.n9909 9.50353
R25311 GND.n8342 GND.n8341 9.50353
R25312 GND.n3474 GND.t157 9.45936
R25313 GND.n6676 GND.t171 9.45936
R25314 GND.n8125 GND.n1530 9.3005
R25315 GND.n2592 GND.n1531 9.3005
R25316 GND.n2594 GND.n2593 9.3005
R25317 GND.n3561 GND.n2591 9.3005
R25318 GND.n3563 GND.n3562 9.3005
R25319 GND.n3564 GND.n2590 9.3005
R25320 GND.n3568 GND.n3565 9.3005
R25321 GND.n3567 GND.n3566 9.3005
R25322 GND.n2570 GND.n2569 9.3005
R25323 GND.n3588 GND.n3587 9.3005
R25324 GND.n3589 GND.n2568 9.3005
R25325 GND.n3593 GND.n3590 9.3005
R25326 GND.n3592 GND.n3591 9.3005
R25327 GND.n2548 GND.n2547 9.3005
R25328 GND.n3614 GND.n3613 9.3005
R25329 GND.n3615 GND.n2546 9.3005
R25330 GND.n3619 GND.n3616 9.3005
R25331 GND.n3618 GND.n3617 9.3005
R25332 GND.n2527 GND.n2526 9.3005
R25333 GND.n3640 GND.n3639 9.3005
R25334 GND.n3641 GND.n2525 9.3005
R25335 GND.n3645 GND.n3642 9.3005
R25336 GND.n3644 GND.n3643 9.3005
R25337 GND.n2506 GND.n2505 9.3005
R25338 GND.n3666 GND.n3665 9.3005
R25339 GND.n3667 GND.n2504 9.3005
R25340 GND.n3671 GND.n3668 9.3005
R25341 GND.n3670 GND.n3669 9.3005
R25342 GND.n2483 GND.n2482 9.3005
R25343 GND.n3691 GND.n3690 9.3005
R25344 GND.n3692 GND.n2481 9.3005
R25345 GND.n3696 GND.n3693 9.3005
R25346 GND.n3695 GND.n3694 9.3005
R25347 GND.n2461 GND.n2460 9.3005
R25348 GND.n3717 GND.n3716 9.3005
R25349 GND.n3718 GND.n2459 9.3005
R25350 GND.n3722 GND.n3719 9.3005
R25351 GND.n3721 GND.n3720 9.3005
R25352 GND.n2442 GND.n2441 9.3005
R25353 GND.n3743 GND.n3742 9.3005
R25354 GND.n3744 GND.n2440 9.3005
R25355 GND.n3748 GND.n3745 9.3005
R25356 GND.n3747 GND.n3746 9.3005
R25357 GND.n2421 GND.n2420 9.3005
R25358 GND.n3769 GND.n3768 9.3005
R25359 GND.n3770 GND.n2419 9.3005
R25360 GND.n3774 GND.n3771 9.3005
R25361 GND.n3773 GND.n3772 9.3005
R25362 GND.n2398 GND.n2397 9.3005
R25363 GND.n3794 GND.n3793 9.3005
R25364 GND.n3795 GND.n2396 9.3005
R25365 GND.n3799 GND.n3796 9.3005
R25366 GND.n3798 GND.n3797 9.3005
R25367 GND.n2376 GND.n2375 9.3005
R25368 GND.n3820 GND.n3819 9.3005
R25369 GND.n3821 GND.n2374 9.3005
R25370 GND.n3826 GND.n3822 9.3005
R25371 GND.n3825 GND.n3824 9.3005
R25372 GND.n3823 GND.n2360 9.3005
R25373 GND.n3845 GND.n2359 9.3005
R25374 GND.n3847 GND.n3846 9.3005
R25375 GND.n1186 GND.n1185 9.3005
R25376 GND.n8502 GND.n8501 9.3005
R25377 GND.n8503 GND.n1184 9.3005
R25378 GND.n8505 GND.n8504 9.3005
R25379 GND.n1180 GND.n1179 9.3005
R25380 GND.n8512 GND.n8511 9.3005
R25381 GND.n8513 GND.n1178 9.3005
R25382 GND.n8515 GND.n8514 9.3005
R25383 GND.n1174 GND.n1173 9.3005
R25384 GND.n8522 GND.n8521 9.3005
R25385 GND.n8523 GND.n1172 9.3005
R25386 GND.n8525 GND.n8524 9.3005
R25387 GND.n1168 GND.n1167 9.3005
R25388 GND.n8532 GND.n8531 9.3005
R25389 GND.n8533 GND.n1166 9.3005
R25390 GND.n8535 GND.n8534 9.3005
R25391 GND.n1162 GND.n1161 9.3005
R25392 GND.n8542 GND.n8541 9.3005
R25393 GND.n8543 GND.n1160 9.3005
R25394 GND.n8545 GND.n8544 9.3005
R25395 GND.n1156 GND.n1155 9.3005
R25396 GND.n8552 GND.n8551 9.3005
R25397 GND.n8553 GND.n1154 9.3005
R25398 GND.n8555 GND.n8554 9.3005
R25399 GND.n1150 GND.n1149 9.3005
R25400 GND.n8562 GND.n8561 9.3005
R25401 GND.n8563 GND.n1148 9.3005
R25402 GND.n8565 GND.n8564 9.3005
R25403 GND.n1144 GND.n1143 9.3005
R25404 GND.n8572 GND.n8571 9.3005
R25405 GND.n8573 GND.n1142 9.3005
R25406 GND.n8575 GND.n8574 9.3005
R25407 GND.n1138 GND.n1137 9.3005
R25408 GND.n8582 GND.n8581 9.3005
R25409 GND.n8583 GND.n1136 9.3005
R25410 GND.n8585 GND.n8584 9.3005
R25411 GND.n1132 GND.n1131 9.3005
R25412 GND.n8592 GND.n8591 9.3005
R25413 GND.n8593 GND.n1130 9.3005
R25414 GND.n8595 GND.n8594 9.3005
R25415 GND.n1126 GND.n1125 9.3005
R25416 GND.n8602 GND.n8601 9.3005
R25417 GND.n8603 GND.n1124 9.3005
R25418 GND.n8605 GND.n8604 9.3005
R25419 GND.n1120 GND.n1119 9.3005
R25420 GND.n8612 GND.n8611 9.3005
R25421 GND.n8613 GND.n1118 9.3005
R25422 GND.n8615 GND.n8614 9.3005
R25423 GND.n1114 GND.n1113 9.3005
R25424 GND.n8622 GND.n8621 9.3005
R25425 GND.n8623 GND.n1112 9.3005
R25426 GND.n8625 GND.n8624 9.3005
R25427 GND.n1108 GND.n1107 9.3005
R25428 GND.n8632 GND.n8631 9.3005
R25429 GND.n8633 GND.n1106 9.3005
R25430 GND.n8635 GND.n8634 9.3005
R25431 GND.n1102 GND.n1101 9.3005
R25432 GND.n8642 GND.n8641 9.3005
R25433 GND.n8643 GND.n1100 9.3005
R25434 GND.n8645 GND.n8644 9.3005
R25435 GND.n1096 GND.n1095 9.3005
R25436 GND.n8652 GND.n8651 9.3005
R25437 GND.n8653 GND.n1094 9.3005
R25438 GND.n8655 GND.n8654 9.3005
R25439 GND.n1090 GND.n1089 9.3005
R25440 GND.n8662 GND.n8661 9.3005
R25441 GND.n8663 GND.n1088 9.3005
R25442 GND.n8665 GND.n8664 9.3005
R25443 GND.n1084 GND.n1083 9.3005
R25444 GND.n8672 GND.n8671 9.3005
R25445 GND.n8673 GND.n1082 9.3005
R25446 GND.n8675 GND.n8674 9.3005
R25447 GND.n1078 GND.n1077 9.3005
R25448 GND.n8682 GND.n8681 9.3005
R25449 GND.n8683 GND.n1076 9.3005
R25450 GND.n8685 GND.n8684 9.3005
R25451 GND.n1072 GND.n1071 9.3005
R25452 GND.n8692 GND.n8691 9.3005
R25453 GND.n8693 GND.n1070 9.3005
R25454 GND.n8695 GND.n8694 9.3005
R25455 GND.n1066 GND.n1065 9.3005
R25456 GND.n8702 GND.n8701 9.3005
R25457 GND.n8703 GND.n1064 9.3005
R25458 GND.n8705 GND.n8704 9.3005
R25459 GND.n1060 GND.n1059 9.3005
R25460 GND.n8712 GND.n8711 9.3005
R25461 GND.n8713 GND.n1058 9.3005
R25462 GND.n8715 GND.n8714 9.3005
R25463 GND.n1054 GND.n1053 9.3005
R25464 GND.n8722 GND.n8721 9.3005
R25465 GND.n8723 GND.n1052 9.3005
R25466 GND.n8725 GND.n8724 9.3005
R25467 GND.n1048 GND.n1047 9.3005
R25468 GND.n8732 GND.n8731 9.3005
R25469 GND.n8733 GND.n1046 9.3005
R25470 GND.n8735 GND.n8734 9.3005
R25471 GND.n1042 GND.n1041 9.3005
R25472 GND.n8742 GND.n8741 9.3005
R25473 GND.n8743 GND.n1040 9.3005
R25474 GND.n8745 GND.n8744 9.3005
R25475 GND.n1036 GND.n1035 9.3005
R25476 GND.n8752 GND.n8751 9.3005
R25477 GND.n8753 GND.n1034 9.3005
R25478 GND.n8755 GND.n8754 9.3005
R25479 GND.n1030 GND.n1029 9.3005
R25480 GND.n8762 GND.n8761 9.3005
R25481 GND.n8763 GND.n1028 9.3005
R25482 GND.n8765 GND.n8764 9.3005
R25483 GND.n1024 GND.n1023 9.3005
R25484 GND.n8772 GND.n8771 9.3005
R25485 GND.n8773 GND.n1022 9.3005
R25486 GND.n8775 GND.n8774 9.3005
R25487 GND.n1018 GND.n1017 9.3005
R25488 GND.n8782 GND.n8781 9.3005
R25489 GND.n8783 GND.n1016 9.3005
R25490 GND.n8785 GND.n8784 9.3005
R25491 GND.n1012 GND.n1011 9.3005
R25492 GND.n8792 GND.n8791 9.3005
R25493 GND.n8793 GND.n1010 9.3005
R25494 GND.n8795 GND.n8794 9.3005
R25495 GND.n1006 GND.n1005 9.3005
R25496 GND.n8802 GND.n8801 9.3005
R25497 GND.n8803 GND.n1004 9.3005
R25498 GND.n8805 GND.n8804 9.3005
R25499 GND.n1000 GND.n999 9.3005
R25500 GND.n8812 GND.n8811 9.3005
R25501 GND.n8813 GND.n998 9.3005
R25502 GND.n8815 GND.n8814 9.3005
R25503 GND.n994 GND.n993 9.3005
R25504 GND.n8822 GND.n8821 9.3005
R25505 GND.n8823 GND.n992 9.3005
R25506 GND.n8825 GND.n8824 9.3005
R25507 GND.n988 GND.n987 9.3005
R25508 GND.n8832 GND.n8831 9.3005
R25509 GND.n8833 GND.n986 9.3005
R25510 GND.n8835 GND.n8834 9.3005
R25511 GND.n982 GND.n981 9.3005
R25512 GND.n8842 GND.n8841 9.3005
R25513 GND.n8843 GND.n980 9.3005
R25514 GND.n8845 GND.n8844 9.3005
R25515 GND.n976 GND.n975 9.3005
R25516 GND.n8852 GND.n8851 9.3005
R25517 GND.n8853 GND.n974 9.3005
R25518 GND.n8855 GND.n8854 9.3005
R25519 GND.n970 GND.n969 9.3005
R25520 GND.n8862 GND.n8861 9.3005
R25521 GND.n8863 GND.n968 9.3005
R25522 GND.n8865 GND.n8864 9.3005
R25523 GND.n964 GND.n963 9.3005
R25524 GND.n8872 GND.n8871 9.3005
R25525 GND.n8873 GND.n962 9.3005
R25526 GND.n8875 GND.n8874 9.3005
R25527 GND.n958 GND.n957 9.3005
R25528 GND.n8882 GND.n8881 9.3005
R25529 GND.n8883 GND.n956 9.3005
R25530 GND.n8885 GND.n8884 9.3005
R25531 GND.n952 GND.n951 9.3005
R25532 GND.n8892 GND.n8891 9.3005
R25533 GND.n8893 GND.n950 9.3005
R25534 GND.n8895 GND.n8894 9.3005
R25535 GND.n946 GND.n945 9.3005
R25536 GND.n8902 GND.n8901 9.3005
R25537 GND.n8903 GND.n944 9.3005
R25538 GND.n8905 GND.n8904 9.3005
R25539 GND.n940 GND.n939 9.3005
R25540 GND.n8912 GND.n8911 9.3005
R25541 GND.n8913 GND.n938 9.3005
R25542 GND.n8915 GND.n8914 9.3005
R25543 GND.n934 GND.n933 9.3005
R25544 GND.n8922 GND.n8921 9.3005
R25545 GND.n8923 GND.n932 9.3005
R25546 GND.n8925 GND.n8924 9.3005
R25547 GND.n928 GND.n927 9.3005
R25548 GND.n8932 GND.n8931 9.3005
R25549 GND.n8933 GND.n926 9.3005
R25550 GND.n8935 GND.n8934 9.3005
R25551 GND.n922 GND.n921 9.3005
R25552 GND.n8942 GND.n8941 9.3005
R25553 GND.n8943 GND.n920 9.3005
R25554 GND.n8945 GND.n8944 9.3005
R25555 GND.n916 GND.n915 9.3005
R25556 GND.n8952 GND.n8951 9.3005
R25557 GND.n8953 GND.n914 9.3005
R25558 GND.n8955 GND.n8954 9.3005
R25559 GND.n910 GND.n909 9.3005
R25560 GND.n8962 GND.n8961 9.3005
R25561 GND.n8963 GND.n908 9.3005
R25562 GND.n8965 GND.n8964 9.3005
R25563 GND.n904 GND.n903 9.3005
R25564 GND.n8972 GND.n8971 9.3005
R25565 GND.n8973 GND.n902 9.3005
R25566 GND.n8975 GND.n8974 9.3005
R25567 GND.n898 GND.n897 9.3005
R25568 GND.n8982 GND.n8981 9.3005
R25569 GND.n8983 GND.n896 9.3005
R25570 GND.n8985 GND.n8984 9.3005
R25571 GND.n892 GND.n891 9.3005
R25572 GND.n8992 GND.n8991 9.3005
R25573 GND.n8993 GND.n890 9.3005
R25574 GND.n8995 GND.n8994 9.3005
R25575 GND.n886 GND.n885 9.3005
R25576 GND.n9002 GND.n9001 9.3005
R25577 GND.n9003 GND.n884 9.3005
R25578 GND.n9005 GND.n9004 9.3005
R25579 GND.n880 GND.n879 9.3005
R25580 GND.n9012 GND.n9011 9.3005
R25581 GND.n9013 GND.n878 9.3005
R25582 GND.n9015 GND.n9014 9.3005
R25583 GND.n874 GND.n873 9.3005
R25584 GND.n9022 GND.n9021 9.3005
R25585 GND.n9023 GND.n872 9.3005
R25586 GND.n9025 GND.n9024 9.3005
R25587 GND.n868 GND.n867 9.3005
R25588 GND.n9032 GND.n9031 9.3005
R25589 GND.n9033 GND.n866 9.3005
R25590 GND.n9035 GND.n9034 9.3005
R25591 GND.n862 GND.n861 9.3005
R25592 GND.n9042 GND.n9041 9.3005
R25593 GND.n9043 GND.n860 9.3005
R25594 GND.n9045 GND.n9044 9.3005
R25595 GND.n856 GND.n855 9.3005
R25596 GND.n9052 GND.n9051 9.3005
R25597 GND.n9053 GND.n854 9.3005
R25598 GND.n9055 GND.n9054 9.3005
R25599 GND.n850 GND.n849 9.3005
R25600 GND.n9062 GND.n9061 9.3005
R25601 GND.n9063 GND.n848 9.3005
R25602 GND.n9065 GND.n9064 9.3005
R25603 GND.n844 GND.n843 9.3005
R25604 GND.n9072 GND.n9071 9.3005
R25605 GND.n9073 GND.n842 9.3005
R25606 GND.n9075 GND.n9074 9.3005
R25607 GND.n838 GND.n837 9.3005
R25608 GND.n9082 GND.n9081 9.3005
R25609 GND.n9083 GND.n836 9.3005
R25610 GND.n9085 GND.n9084 9.3005
R25611 GND.n832 GND.n831 9.3005
R25612 GND.n9092 GND.n9091 9.3005
R25613 GND.n9093 GND.n830 9.3005
R25614 GND.n9095 GND.n9094 9.3005
R25615 GND.n826 GND.n825 9.3005
R25616 GND.n9102 GND.n9101 9.3005
R25617 GND.n9103 GND.n824 9.3005
R25618 GND.n9105 GND.n9104 9.3005
R25619 GND.n820 GND.n819 9.3005
R25620 GND.n9112 GND.n9111 9.3005
R25621 GND.n9113 GND.n818 9.3005
R25622 GND.n9115 GND.n9114 9.3005
R25623 GND.n814 GND.n813 9.3005
R25624 GND.n9122 GND.n9121 9.3005
R25625 GND.n9123 GND.n812 9.3005
R25626 GND.n9125 GND.n9124 9.3005
R25627 GND.n808 GND.n807 9.3005
R25628 GND.n9132 GND.n9131 9.3005
R25629 GND.n9133 GND.n806 9.3005
R25630 GND.n9135 GND.n9134 9.3005
R25631 GND.n802 GND.n801 9.3005
R25632 GND.n9142 GND.n9141 9.3005
R25633 GND.n9143 GND.n800 9.3005
R25634 GND.n9145 GND.n9144 9.3005
R25635 GND.n796 GND.n795 9.3005
R25636 GND.n9152 GND.n9151 9.3005
R25637 GND.n9153 GND.n794 9.3005
R25638 GND.n9155 GND.n9154 9.3005
R25639 GND.n790 GND.n789 9.3005
R25640 GND.n9162 GND.n9161 9.3005
R25641 GND.n9163 GND.n788 9.3005
R25642 GND.n9165 GND.n9164 9.3005
R25643 GND.n784 GND.n783 9.3005
R25644 GND.n9172 GND.n9171 9.3005
R25645 GND.n9173 GND.n782 9.3005
R25646 GND.n9175 GND.n9174 9.3005
R25647 GND.n778 GND.n777 9.3005
R25648 GND.n9182 GND.n9181 9.3005
R25649 GND.n9183 GND.n776 9.3005
R25650 GND.n9185 GND.n9184 9.3005
R25651 GND.n772 GND.n771 9.3005
R25652 GND.n9192 GND.n9191 9.3005
R25653 GND.n9193 GND.n770 9.3005
R25654 GND.n9195 GND.n9194 9.3005
R25655 GND.n766 GND.n765 9.3005
R25656 GND.n9202 GND.n9201 9.3005
R25657 GND.n9203 GND.n764 9.3005
R25658 GND.n9205 GND.n9204 9.3005
R25659 GND.n760 GND.n759 9.3005
R25660 GND.n9212 GND.n9211 9.3005
R25661 GND.n9213 GND.n758 9.3005
R25662 GND.n9215 GND.n9214 9.3005
R25663 GND.n754 GND.n753 9.3005
R25664 GND.n9222 GND.n9221 9.3005
R25665 GND.n9223 GND.n752 9.3005
R25666 GND.n9225 GND.n9224 9.3005
R25667 GND.n748 GND.n747 9.3005
R25668 GND.n9232 GND.n9231 9.3005
R25669 GND.n9233 GND.n746 9.3005
R25670 GND.n9235 GND.n9234 9.3005
R25671 GND.n742 GND.n741 9.3005
R25672 GND.n9242 GND.n9241 9.3005
R25673 GND.n9243 GND.n740 9.3005
R25674 GND.n9245 GND.n9244 9.3005
R25675 GND.n736 GND.n735 9.3005
R25676 GND.n9252 GND.n9251 9.3005
R25677 GND.n9253 GND.n734 9.3005
R25678 GND.n9255 GND.n9254 9.3005
R25679 GND.n730 GND.n729 9.3005
R25680 GND.n9262 GND.n9261 9.3005
R25681 GND.n9263 GND.n728 9.3005
R25682 GND.n9265 GND.n9264 9.3005
R25683 GND.n724 GND.n723 9.3005
R25684 GND.n9272 GND.n9271 9.3005
R25685 GND.n9273 GND.n722 9.3005
R25686 GND.n9275 GND.n9274 9.3005
R25687 GND.n718 GND.n717 9.3005
R25688 GND.n9282 GND.n9281 9.3005
R25689 GND.n9283 GND.n716 9.3005
R25690 GND.n9285 GND.n9284 9.3005
R25691 GND.n712 GND.n711 9.3005
R25692 GND.n9292 GND.n9291 9.3005
R25693 GND.n9293 GND.n710 9.3005
R25694 GND.n9295 GND.n9294 9.3005
R25695 GND.n706 GND.n705 9.3005
R25696 GND.n9302 GND.n9301 9.3005
R25697 GND.n9303 GND.n704 9.3005
R25698 GND.n9305 GND.n9304 9.3005
R25699 GND.n700 GND.n699 9.3005
R25700 GND.n9312 GND.n9311 9.3005
R25701 GND.n9313 GND.n698 9.3005
R25702 GND.n9315 GND.n9314 9.3005
R25703 GND.n694 GND.n693 9.3005
R25704 GND.n9322 GND.n9321 9.3005
R25705 GND.n9323 GND.n692 9.3005
R25706 GND.n9325 GND.n9324 9.3005
R25707 GND.n688 GND.n687 9.3005
R25708 GND.n9332 GND.n9331 9.3005
R25709 GND.n9333 GND.n686 9.3005
R25710 GND.n9335 GND.n9334 9.3005
R25711 GND.n682 GND.n681 9.3005
R25712 GND.n9342 GND.n9341 9.3005
R25713 GND.n9343 GND.n680 9.3005
R25714 GND.n9345 GND.n9344 9.3005
R25715 GND.n676 GND.n675 9.3005
R25716 GND.n9352 GND.n9351 9.3005
R25717 GND.n9353 GND.n674 9.3005
R25718 GND.n9355 GND.n9354 9.3005
R25719 GND.n670 GND.n669 9.3005
R25720 GND.n9362 GND.n9361 9.3005
R25721 GND.n9363 GND.n668 9.3005
R25722 GND.n9365 GND.n9364 9.3005
R25723 GND.n664 GND.n663 9.3005
R25724 GND.n9372 GND.n9371 9.3005
R25725 GND.n9373 GND.n662 9.3005
R25726 GND.n9375 GND.n9374 9.3005
R25727 GND.n658 GND.n657 9.3005
R25728 GND.n9382 GND.n9381 9.3005
R25729 GND.n9383 GND.n656 9.3005
R25730 GND.n9385 GND.n9384 9.3005
R25731 GND.n652 GND.n651 9.3005
R25732 GND.n9392 GND.n9391 9.3005
R25733 GND.n9393 GND.n650 9.3005
R25734 GND.n9395 GND.n9394 9.3005
R25735 GND.n646 GND.n645 9.3005
R25736 GND.n9402 GND.n9401 9.3005
R25737 GND.n9403 GND.n644 9.3005
R25738 GND.n9405 GND.n9404 9.3005
R25739 GND.n640 GND.n639 9.3005
R25740 GND.n9412 GND.n9411 9.3005
R25741 GND.n9413 GND.n638 9.3005
R25742 GND.n9415 GND.n9414 9.3005
R25743 GND.n634 GND.n633 9.3005
R25744 GND.n9422 GND.n9421 9.3005
R25745 GND.n9423 GND.n632 9.3005
R25746 GND.n9425 GND.n9424 9.3005
R25747 GND.n628 GND.n627 9.3005
R25748 GND.n9432 GND.n9431 9.3005
R25749 GND.n9433 GND.n626 9.3005
R25750 GND.n9435 GND.n9434 9.3005
R25751 GND.n622 GND.n621 9.3005
R25752 GND.n9442 GND.n9441 9.3005
R25753 GND.n9443 GND.n620 9.3005
R25754 GND.n9445 GND.n9444 9.3005
R25755 GND.n616 GND.n615 9.3005
R25756 GND.n9452 GND.n9451 9.3005
R25757 GND.n9453 GND.n614 9.3005
R25758 GND.n9455 GND.n9454 9.3005
R25759 GND.n610 GND.n609 9.3005
R25760 GND.n9462 GND.n9461 9.3005
R25761 GND.n9463 GND.n608 9.3005
R25762 GND.n9465 GND.n9464 9.3005
R25763 GND.n604 GND.n603 9.3005
R25764 GND.n9472 GND.n9471 9.3005
R25765 GND.n9473 GND.n602 9.3005
R25766 GND.n9475 GND.n9474 9.3005
R25767 GND.n598 GND.n597 9.3005
R25768 GND.n9482 GND.n9481 9.3005
R25769 GND.n9483 GND.n596 9.3005
R25770 GND.n9485 GND.n9484 9.3005
R25771 GND.n592 GND.n591 9.3005
R25772 GND.n9492 GND.n9491 9.3005
R25773 GND.n9493 GND.n590 9.3005
R25774 GND.n9495 GND.n9494 9.3005
R25775 GND.n586 GND.n585 9.3005
R25776 GND.n9502 GND.n9501 9.3005
R25777 GND.n9503 GND.n584 9.3005
R25778 GND.n9505 GND.n9504 9.3005
R25779 GND.n580 GND.n579 9.3005
R25780 GND.n9512 GND.n9511 9.3005
R25781 GND.n9513 GND.n578 9.3005
R25782 GND.n9516 GND.n9515 9.3005
R25783 GND.n9514 GND.n574 9.3005
R25784 GND.n9522 GND.n573 9.3005
R25785 GND.n9524 GND.n9523 9.3005
R25786 GND.n569 GND.n568 9.3005
R25787 GND.n9533 GND.n9532 9.3005
R25788 GND.n9534 GND.n567 9.3005
R25789 GND.n9536 GND.n9535 9.3005
R25790 GND.n563 GND.n562 9.3005
R25791 GND.n9543 GND.n9542 9.3005
R25792 GND.n9544 GND.n561 9.3005
R25793 GND.n9546 GND.n9545 9.3005
R25794 GND.n557 GND.n556 9.3005
R25795 GND.n9553 GND.n9552 9.3005
R25796 GND.n9554 GND.n555 9.3005
R25797 GND.n9556 GND.n9555 9.3005
R25798 GND.n551 GND.n550 9.3005
R25799 GND.n9563 GND.n9562 9.3005
R25800 GND.n9564 GND.n549 9.3005
R25801 GND.n9566 GND.n9565 9.3005
R25802 GND.n545 GND.n544 9.3005
R25803 GND.n9573 GND.n9572 9.3005
R25804 GND.n9574 GND.n543 9.3005
R25805 GND.n9576 GND.n9575 9.3005
R25806 GND.n539 GND.n538 9.3005
R25807 GND.n9583 GND.n9582 9.3005
R25808 GND.n9584 GND.n537 9.3005
R25809 GND.n9586 GND.n9585 9.3005
R25810 GND.n533 GND.n532 9.3005
R25811 GND.n9593 GND.n9592 9.3005
R25812 GND.n9594 GND.n531 9.3005
R25813 GND.n9596 GND.n9595 9.3005
R25814 GND.n527 GND.n526 9.3005
R25815 GND.n9603 GND.n9602 9.3005
R25816 GND.n9604 GND.n525 9.3005
R25817 GND.n9606 GND.n9605 9.3005
R25818 GND.n521 GND.n520 9.3005
R25819 GND.n9613 GND.n9612 9.3005
R25820 GND.n9614 GND.n519 9.3005
R25821 GND.n9616 GND.n9615 9.3005
R25822 GND.n515 GND.n514 9.3005
R25823 GND.n9623 GND.n9622 9.3005
R25824 GND.n9624 GND.n513 9.3005
R25825 GND.n9626 GND.n9625 9.3005
R25826 GND.n509 GND.n508 9.3005
R25827 GND.n9633 GND.n9632 9.3005
R25828 GND.n9634 GND.n507 9.3005
R25829 GND.n9636 GND.n9635 9.3005
R25830 GND.n503 GND.n502 9.3005
R25831 GND.n9643 GND.n9642 9.3005
R25832 GND.n9644 GND.n501 9.3005
R25833 GND.n9646 GND.n9645 9.3005
R25834 GND.n497 GND.n496 9.3005
R25835 GND.n9653 GND.n9652 9.3005
R25836 GND.n9654 GND.n495 9.3005
R25837 GND.n9656 GND.n9655 9.3005
R25838 GND.n491 GND.n490 9.3005
R25839 GND.n9663 GND.n9662 9.3005
R25840 GND.n9664 GND.n489 9.3005
R25841 GND.n9666 GND.n9665 9.3005
R25842 GND.n485 GND.n484 9.3005
R25843 GND.n9673 GND.n9672 9.3005
R25844 GND.n9674 GND.n483 9.3005
R25845 GND.n9676 GND.n9675 9.3005
R25846 GND.n479 GND.n478 9.3005
R25847 GND.n9683 GND.n9682 9.3005
R25848 GND.n9684 GND.n477 9.3005
R25849 GND.n9690 GND.n9685 9.3005
R25850 GND.n9689 GND.n9688 9.3005
R25851 GND.n9687 GND.n474 9.3005
R25852 GND.n9526 GND.n9525 9.3005
R25853 GND.n5683 GND.n5682 9.3005
R25854 GND.n5681 GND.n5670 9.3005
R25855 GND.n5680 GND.n5679 9.3005
R25856 GND.n5677 GND.n5672 9.3005
R25857 GND.n5676 GND.n5674 9.3005
R25858 GND.n5673 GND.n5653 9.3005
R25859 GND.n5761 GND.n5652 9.3005
R25860 GND.n5763 GND.n5762 9.3005
R25861 GND.n5764 GND.n5651 9.3005
R25862 GND.n5766 GND.n5765 9.3005
R25863 GND.n5767 GND.n5648 9.3005
R25864 GND.n5771 GND.n5770 9.3005
R25865 GND.n5772 GND.n5647 9.3005
R25866 GND.n5795 GND.n5773 9.3005
R25867 GND.n5794 GND.n5774 9.3005
R25868 GND.n5793 GND.n5775 9.3005
R25869 GND.n5791 GND.n5776 9.3005
R25870 GND.n5790 GND.n5777 9.3005
R25871 GND.n5788 GND.n5778 9.3005
R25872 GND.n5787 GND.n5779 9.3005
R25873 GND.n5785 GND.n5780 9.3005
R25874 GND.n5784 GND.n5782 9.3005
R25875 GND.n5781 GND.n5622 9.3005
R25876 GND.n5865 GND.n5621 9.3005
R25877 GND.n5867 GND.n5866 9.3005
R25878 GND.n5868 GND.n5620 9.3005
R25879 GND.n5870 GND.n5869 9.3005
R25880 GND.n5871 GND.n5617 9.3005
R25881 GND.n5875 GND.n5874 9.3005
R25882 GND.n5876 GND.n5616 9.3005
R25883 GND.n5899 GND.n5877 9.3005
R25884 GND.n5898 GND.n5878 9.3005
R25885 GND.n5897 GND.n5879 9.3005
R25886 GND.n5895 GND.n5880 9.3005
R25887 GND.n5894 GND.n5881 9.3005
R25888 GND.n5892 GND.n5882 9.3005
R25889 GND.n5891 GND.n5883 9.3005
R25890 GND.n5889 GND.n5884 9.3005
R25891 GND.n5888 GND.n5886 9.3005
R25892 GND.n5885 GND.n5591 9.3005
R25893 GND.n5968 GND.n5590 9.3005
R25894 GND.n5970 GND.n5969 9.3005
R25895 GND.n5971 GND.n5589 9.3005
R25896 GND.n5973 GND.n5972 9.3005
R25897 GND.n5974 GND.n5586 9.3005
R25898 GND.n5978 GND.n5977 9.3005
R25899 GND.n5979 GND.n5585 9.3005
R25900 GND.n6002 GND.n5980 9.3005
R25901 GND.n6001 GND.n5981 9.3005
R25902 GND.n6000 GND.n5982 9.3005
R25903 GND.n5998 GND.n5983 9.3005
R25904 GND.n5997 GND.n5984 9.3005
R25905 GND.n5995 GND.n5985 9.3005
R25906 GND.n5994 GND.n5986 9.3005
R25907 GND.n5992 GND.n5987 9.3005
R25908 GND.n5991 GND.n5989 9.3005
R25909 GND.n5988 GND.n5558 9.3005
R25910 GND.n6071 GND.n5557 9.3005
R25911 GND.n6073 GND.n6072 9.3005
R25912 GND.n6074 GND.n5556 9.3005
R25913 GND.n6076 GND.n6075 9.3005
R25914 GND.n6077 GND.n5553 9.3005
R25915 GND.n6081 GND.n6080 9.3005
R25916 GND.n6082 GND.n5552 9.3005
R25917 GND.n6105 GND.n6083 9.3005
R25918 GND.n6104 GND.n6084 9.3005
R25919 GND.n6103 GND.n6085 9.3005
R25920 GND.n6101 GND.n6086 9.3005
R25921 GND.n6100 GND.n6087 9.3005
R25922 GND.n6098 GND.n6088 9.3005
R25923 GND.n6097 GND.n6089 9.3005
R25924 GND.n6095 GND.n6090 9.3005
R25925 GND.n6094 GND.n6092 9.3005
R25926 GND.n6091 GND.n5526 9.3005
R25927 GND.n6174 GND.n5525 9.3005
R25928 GND.n6176 GND.n6175 9.3005
R25929 GND.n6177 GND.n5524 9.3005
R25930 GND.n6179 GND.n6178 9.3005
R25931 GND.n6180 GND.n5521 9.3005
R25932 GND.n6184 GND.n6183 9.3005
R25933 GND.n6185 GND.n5520 9.3005
R25934 GND.n6201 GND.n6186 9.3005
R25935 GND.n6200 GND.n6187 9.3005
R25936 GND.n6199 GND.n6188 9.3005
R25937 GND.n6197 GND.n6189 9.3005
R25938 GND.n6196 GND.n6190 9.3005
R25939 GND.n6193 GND.n6192 9.3005
R25940 GND.n6191 GND.n5496 9.3005
R25941 GND.n5671 GND.n5669 9.3005
R25942 GND.n7740 GND.n2354 9.3005
R25943 GND.n7743 GND.n2353 9.3005
R25944 GND.n7744 GND.n2352 9.3005
R25945 GND.n7747 GND.n2351 9.3005
R25946 GND.n7748 GND.n2350 9.3005
R25947 GND.n7751 GND.n2349 9.3005
R25948 GND.n7753 GND.n2348 9.3005
R25949 GND.n7754 GND.n2347 9.3005
R25950 GND.n7755 GND.n2346 9.3005
R25951 GND.n7756 GND.n2345 9.3005
R25952 GND.n7703 GND.n7702 9.3005
R25953 GND.n7704 GND.n3879 9.3005
R25954 GND.n7707 GND.n3878 9.3005
R25955 GND.n7710 GND.n2358 9.3005
R25956 GND.n7701 GND.n3881 9.3005
R25957 GND.n3883 GND.n3882 9.3005
R25958 GND.n7689 GND.n3898 9.3005
R25959 GND.n7688 GND.n3899 9.3005
R25960 GND.n7687 GND.n3900 9.3005
R25961 GND.n3917 GND.n3901 9.3005
R25962 GND.n7678 GND.n3918 9.3005
R25963 GND.n7677 GND.n3919 9.3005
R25964 GND.n7676 GND.n3920 9.3005
R25965 GND.n3972 GND.n3921 9.3005
R25966 GND.n3973 GND.n3971 9.3005
R25967 GND.n3975 GND.n3974 9.3005
R25968 GND.n3978 GND.n3970 9.3005
R25969 GND.n3980 GND.n3979 9.3005
R25970 GND.n3981 GND.n3969 9.3005
R25971 GND.n7647 GND.n3982 9.3005
R25972 GND.n7646 GND.n3983 9.3005
R25973 GND.n7645 GND.n3984 9.3005
R25974 GND.n4001 GND.n3985 9.3005
R25975 GND.n7635 GND.n4002 9.3005
R25976 GND.n7634 GND.n4003 9.3005
R25977 GND.n7633 GND.n4004 9.3005
R25978 GND.n4021 GND.n4005 9.3005
R25979 GND.n7623 GND.n4022 9.3005
R25980 GND.n7622 GND.n4023 9.3005
R25981 GND.n7621 GND.n4024 9.3005
R25982 GND.n4077 GND.n4025 9.3005
R25983 GND.n4078 GND.n4076 9.3005
R25984 GND.n4080 GND.n4079 9.3005
R25985 GND.n4083 GND.n4075 9.3005
R25986 GND.n4085 GND.n4084 9.3005
R25987 GND.n4086 GND.n4074 9.3005
R25988 GND.n7592 GND.n4087 9.3005
R25989 GND.n7591 GND.n4088 9.3005
R25990 GND.n7590 GND.n4089 9.3005
R25991 GND.n4106 GND.n4090 9.3005
R25992 GND.n7580 GND.n4107 9.3005
R25993 GND.n7579 GND.n4108 9.3005
R25994 GND.n7578 GND.n4109 9.3005
R25995 GND.n4126 GND.n4110 9.3005
R25996 GND.n7568 GND.n4127 9.3005
R25997 GND.n7567 GND.n4128 9.3005
R25998 GND.n7566 GND.n4129 9.3005
R25999 GND.n4182 GND.n4130 9.3005
R26000 GND.n4183 GND.n4181 9.3005
R26001 GND.n4185 GND.n4184 9.3005
R26002 GND.n4188 GND.n4180 9.3005
R26003 GND.n4190 GND.n4189 9.3005
R26004 GND.n4191 GND.n4179 9.3005
R26005 GND.n7537 GND.n4192 9.3005
R26006 GND.n7536 GND.n4193 9.3005
R26007 GND.n7535 GND.n4194 9.3005
R26008 GND.n4210 GND.n4195 9.3005
R26009 GND.n7525 GND.n4211 9.3005
R26010 GND.n7524 GND.n4212 9.3005
R26011 GND.n7523 GND.n4213 9.3005
R26012 GND.n4229 GND.n4214 9.3005
R26013 GND.n7513 GND.n4230 9.3005
R26014 GND.n7512 GND.n4231 9.3005
R26015 GND.n7511 GND.n4232 9.3005
R26016 GND.n4284 GND.n4233 9.3005
R26017 GND.n4285 GND.n4283 9.3005
R26018 GND.n4287 GND.n4286 9.3005
R26019 GND.n4290 GND.n4282 9.3005
R26020 GND.n4292 GND.n4291 9.3005
R26021 GND.n4293 GND.n4281 9.3005
R26022 GND.n7482 GND.n4294 9.3005
R26023 GND.n7481 GND.n4295 9.3005
R26024 GND.n7480 GND.n4296 9.3005
R26025 GND.n4313 GND.n4297 9.3005
R26026 GND.n7470 GND.n4314 9.3005
R26027 GND.n7469 GND.n4315 9.3005
R26028 GND.n7468 GND.n4316 9.3005
R26029 GND.n4333 GND.n4317 9.3005
R26030 GND.n7458 GND.n4334 9.3005
R26031 GND.n7457 GND.n4335 9.3005
R26032 GND.n7456 GND.n4336 9.3005
R26033 GND.n4389 GND.n4337 9.3005
R26034 GND.n4390 GND.n4388 9.3005
R26035 GND.n4392 GND.n4391 9.3005
R26036 GND.n4395 GND.n4387 9.3005
R26037 GND.n4397 GND.n4396 9.3005
R26038 GND.n4398 GND.n4386 9.3005
R26039 GND.n7427 GND.n4399 9.3005
R26040 GND.n7426 GND.n4400 9.3005
R26041 GND.n7425 GND.n4401 9.3005
R26042 GND.n4417 GND.n4402 9.3005
R26043 GND.n7415 GND.n4418 9.3005
R26044 GND.n7414 GND.n7413 9.3005
R26045 GND.n7700 GND.n7699 9.3005
R26046 GND.n6349 GND.n6345 9.3005
R26047 GND.n6348 GND.n6346 9.3005
R26048 GND.n4420 GND.n4419 9.3005
R26049 GND.n7412 GND.n7411 9.3005
R26050 GND.n6316 GND.n5494 9.3005
R26051 GND.n6320 GND.n6319 9.3005
R26052 GND.n6321 GND.n5493 9.3005
R26053 GND.n6325 GND.n6322 9.3005
R26054 GND.n6326 GND.n5492 9.3005
R26055 GND.n6330 GND.n6329 9.3005
R26056 GND.n6331 GND.n5491 9.3005
R26057 GND.n6335 GND.n6332 9.3005
R26058 GND.n6336 GND.n5464 9.3005
R26059 GND.n6352 GND.n5465 9.3005
R26060 GND.n6315 GND.n5495 9.3005
R26061 GND.n6356 GND.n6355 9.3005
R26062 GND.n6420 GND.n5365 9.3005
R26063 GND.n6422 GND.n6421 9.3005
R26064 GND.n6423 GND.n5364 9.3005
R26065 GND.n6427 GND.n6426 9.3005
R26066 GND.n6428 GND.n5363 9.3005
R26067 GND.n6430 GND.n6429 9.3005
R26068 GND.n5350 GND.n5349 9.3005
R26069 GND.n6482 GND.n6481 9.3005
R26070 GND.n6483 GND.n5348 9.3005
R26071 GND.n6485 GND.n6484 9.3005
R26072 GND.n5345 GND.n5344 9.3005
R26073 GND.n6496 GND.n6495 9.3005
R26074 GND.n6497 GND.n5343 9.3005
R26075 GND.n6499 GND.n6498 9.3005
R26076 GND.n5340 GND.n5339 9.3005
R26077 GND.n6510 GND.n6509 9.3005
R26078 GND.n6511 GND.n5338 9.3005
R26079 GND.n6514 GND.n6513 9.3005
R26080 GND.n6512 GND.n5331 9.3005
R26081 GND.n6673 GND.n5332 9.3005
R26082 GND.n6672 GND.n5333 9.3005
R26083 GND.n6671 GND.n5334 9.3005
R26084 GND.n6524 GND.n5335 9.3005
R26085 GND.n6661 GND.n6525 9.3005
R26086 GND.n6660 GND.n6526 9.3005
R26087 GND.n6659 GND.n6527 9.3005
R26088 GND.n6531 GND.n6528 9.3005
R26089 GND.n6649 GND.n6532 9.3005
R26090 GND.n6648 GND.n6533 9.3005
R26091 GND.n6647 GND.n6534 9.3005
R26092 GND.n6538 GND.n6535 9.3005
R26093 GND.n6637 GND.n6539 9.3005
R26094 GND.n6636 GND.n6540 9.3005
R26095 GND.n6635 GND.n6541 9.3005
R26096 GND.n6545 GND.n6542 9.3005
R26097 GND.n6625 GND.n6546 9.3005
R26098 GND.n6624 GND.n6547 9.3005
R26099 GND.n6623 GND.n6548 9.3005
R26100 GND.n6552 GND.n6549 9.3005
R26101 GND.n6613 GND.n6553 9.3005
R26102 GND.n6612 GND.n6554 9.3005
R26103 GND.n6611 GND.n6555 9.3005
R26104 GND.n6559 GND.n6556 9.3005
R26105 GND.n6601 GND.n6560 9.3005
R26106 GND.n6600 GND.n6561 9.3005
R26107 GND.n6599 GND.n6562 9.3005
R26108 GND.n6566 GND.n6563 9.3005
R26109 GND.n6589 GND.n6567 9.3005
R26110 GND.n6588 GND.n6568 9.3005
R26111 GND.n6587 GND.n6569 9.3005
R26112 GND.n6575 GND.n6570 9.3005
R26113 GND.n6577 GND.n6576 9.3005
R26114 GND.n5290 GND.n5289 9.3005
R26115 GND.n6757 GND.n6756 9.3005
R26116 GND.n6758 GND.n5288 9.3005
R26117 GND.n6767 GND.n6759 9.3005
R26118 GND.n6766 GND.n6760 9.3005
R26119 GND.n6765 GND.n6761 9.3005
R26120 GND.n6764 GND.n6762 9.3005
R26121 GND.n104 GND.n102 9.3005
R26122 GND.n6419 GND.n6418 9.3005
R26123 GND.n10313 GND.n10312 9.3005
R26124 GND.n105 GND.n103 9.3005
R26125 GND.n5273 GND.n5272 9.3005
R26126 GND.n6899 GND.n5274 9.3005
R26127 GND.n6898 GND.n5275 9.3005
R26128 GND.n6897 GND.n5276 9.3005
R26129 GND.n6798 GND.n5277 9.3005
R26130 GND.n6887 GND.n6799 9.3005
R26131 GND.n6886 GND.n6800 9.3005
R26132 GND.n6885 GND.n6801 9.3005
R26133 GND.n6805 GND.n6802 9.3005
R26134 GND.n6875 GND.n6806 9.3005
R26135 GND.n6874 GND.n6807 9.3005
R26136 GND.n6873 GND.n6808 9.3005
R26137 GND.n6812 GND.n6809 9.3005
R26138 GND.n6863 GND.n6813 9.3005
R26139 GND.n6862 GND.n6814 9.3005
R26140 GND.n6861 GND.n6815 9.3005
R26141 GND.n6819 GND.n6816 9.3005
R26142 GND.n6851 GND.n6820 9.3005
R26143 GND.n6850 GND.n6821 9.3005
R26144 GND.n6849 GND.n6822 9.3005
R26145 GND.n6826 GND.n6823 9.3005
R26146 GND.n6839 GND.n6827 9.3005
R26147 GND.n6838 GND.n6828 9.3005
R26148 GND.n6837 GND.n6829 9.3005
R26149 GND.n440 GND.n439 9.3005
R26150 GND.n9730 GND.n9729 9.3005
R26151 GND.n9731 GND.n438 9.3005
R26152 GND.n9733 GND.n9732 9.3005
R26153 GND.n436 GND.n435 9.3005
R26154 GND.n9745 GND.n9744 9.3005
R26155 GND.n9746 GND.n434 9.3005
R26156 GND.n9748 GND.n9747 9.3005
R26157 GND.n432 GND.n431 9.3005
R26158 GND.n9760 GND.n9759 9.3005
R26159 GND.n9761 GND.n430 9.3005
R26160 GND.n9763 GND.n9762 9.3005
R26161 GND.n428 GND.n427 9.3005
R26162 GND.n9775 GND.n9774 9.3005
R26163 GND.n9776 GND.n426 9.3005
R26164 GND.n9778 GND.n9777 9.3005
R26165 GND.n424 GND.n423 9.3005
R26166 GND.n9790 GND.n9789 9.3005
R26167 GND.n9791 GND.n422 9.3005
R26168 GND.n10102 GND.n9792 9.3005
R26169 GND.n10101 GND.n9793 9.3005
R26170 GND.n10100 GND.n9794 9.3005
R26171 GND.n10098 GND.n9795 9.3005
R26172 GND.n10097 GND.n9796 9.3005
R26173 GND.n10095 GND.n9797 9.3005
R26174 GND.n10094 GND.n9798 9.3005
R26175 GND.n10092 GND.n9799 9.3005
R26176 GND.n10091 GND.n9800 9.3005
R26177 GND.n10089 GND.n9801 9.3005
R26178 GND.n10088 GND.n9802 9.3005
R26179 GND.n10086 GND.n9803 9.3005
R26180 GND.n10085 GND.n9804 9.3005
R26181 GND.n10083 GND.n9805 9.3005
R26182 GND.n10082 GND.n9806 9.3005
R26183 GND.n10080 GND.n10079 9.3005
R26184 GND.n10052 GND.n10051 9.3005
R26185 GND.n10055 GND.n10048 9.3005
R26186 GND.n10059 GND.n10058 9.3005
R26187 GND.n10060 GND.n10047 9.3005
R26188 GND.n10062 GND.n10061 9.3005
R26189 GND.n10065 GND.n10046 9.3005
R26190 GND.n10068 GND.n10067 9.3005
R26191 GND.n10069 GND.n10045 9.3005
R26192 GND.n10071 GND.n10070 9.3005
R26193 GND.n9810 GND.n9807 9.3005
R26194 GND.n10078 GND.n10077 9.3005
R26195 GND.n10050 GND.n10049 9.3005
R26196 GND.n9887 GND.n9886 9.3005
R26197 GND.n9890 GND.n9883 9.3005
R26198 GND.n9894 GND.n9893 9.3005
R26199 GND.n9895 GND.n9882 9.3005
R26200 GND.n9897 GND.n9896 9.3005
R26201 GND.n9900 GND.n9881 9.3005
R26202 GND.n9904 GND.n9903 9.3005
R26203 GND.n9905 GND.n9880 9.3005
R26204 GND.n9908 GND.n9906 9.3005
R26205 GND.n9909 GND.n9876 9.3005
R26206 GND.n9913 GND.n9912 9.3005
R26207 GND.n9914 GND.n9875 9.3005
R26208 GND.n9916 GND.n9915 9.3005
R26209 GND.n9919 GND.n9874 9.3005
R26210 GND.n9923 GND.n9922 9.3005
R26211 GND.n9924 GND.n9873 9.3005
R26212 GND.n9926 GND.n9925 9.3005
R26213 GND.n9929 GND.n9872 9.3005
R26214 GND.n9933 GND.n9932 9.3005
R26215 GND.n9934 GND.n9871 9.3005
R26216 GND.n9936 GND.n9935 9.3005
R26217 GND.n9939 GND.n9868 9.3005
R26218 GND.n9944 GND.n9943 9.3005
R26219 GND.n9945 GND.n9867 9.3005
R26220 GND.n9947 GND.n9946 9.3005
R26221 GND.n9950 GND.n9866 9.3005
R26222 GND.n9954 GND.n9953 9.3005
R26223 GND.n9955 GND.n9865 9.3005
R26224 GND.n9957 GND.n9956 9.3005
R26225 GND.n9960 GND.n9864 9.3005
R26226 GND.n9964 GND.n9963 9.3005
R26227 GND.n9965 GND.n9863 9.3005
R26228 GND.n9967 GND.n9966 9.3005
R26229 GND.n9970 GND.n9858 9.3005
R26230 GND.n9972 GND.n9971 9.3005
R26231 GND.n9973 GND.n9857 9.3005
R26232 GND.n9975 GND.n9974 9.3005
R26233 GND.n9978 GND.n9856 9.3005
R26234 GND.n9982 GND.n9981 9.3005
R26235 GND.n9983 GND.n9855 9.3005
R26236 GND.n9985 GND.n9984 9.3005
R26237 GND.n9988 GND.n9854 9.3005
R26238 GND.n9992 GND.n9991 9.3005
R26239 GND.n9993 GND.n9853 9.3005
R26240 GND.n9995 GND.n9994 9.3005
R26241 GND.n9998 GND.n9852 9.3005
R26242 GND.n10005 GND.n10004 9.3005
R26243 GND.n10006 GND.n9851 9.3005
R26244 GND.n10008 GND.n10007 9.3005
R26245 GND.n10011 GND.n9850 9.3005
R26246 GND.n10015 GND.n10014 9.3005
R26247 GND.n10016 GND.n9849 9.3005
R26248 GND.n10018 GND.n10017 9.3005
R26249 GND.n10021 GND.n9848 9.3005
R26250 GND.n10025 GND.n10024 9.3005
R26251 GND.n10026 GND.n9847 9.3005
R26252 GND.n10028 GND.n10027 9.3005
R26253 GND.n10031 GND.n9846 9.3005
R26254 GND.n10034 GND.n10033 9.3005
R26255 GND.n10035 GND.n9845 9.3005
R26256 GND.n10037 GND.n10036 9.3005
R26257 GND.n9885 GND.n9884 9.3005
R26258 GND.n7089 GND.n7088 9.3005
R26259 GND.n4891 GND.n4889 9.3005
R26260 GND.n5356 GND.n5355 9.3005
R26261 GND.n5359 GND.n5354 9.3005
R26262 GND.n5361 GND.n5360 9.3005
R26263 GND.n5362 GND.n4929 9.3005
R26264 GND.n7068 GND.n4930 9.3005
R26265 GND.n7067 GND.n4931 9.3005
R26266 GND.n7066 GND.n4932 9.3005
R26267 GND.n5347 GND.n4933 9.3005
R26268 GND.n7056 GND.n4951 9.3005
R26269 GND.n7055 GND.n4952 9.3005
R26270 GND.n7054 GND.n4953 9.3005
R26271 GND.n5342 GND.n4954 9.3005
R26272 GND.n7044 GND.n4972 9.3005
R26273 GND.n7043 GND.n4973 9.3005
R26274 GND.n7042 GND.n4974 9.3005
R26275 GND.n5337 GND.n4975 9.3005
R26276 GND.n7032 GND.n4993 9.3005
R26277 GND.n7031 GND.n4994 9.3005
R26278 GND.n7030 GND.n4995 9.3005
R26279 GND.n6522 GND.n4996 9.3005
R26280 GND.n7020 GND.n5013 9.3005
R26281 GND.n7019 GND.n5014 9.3005
R26282 GND.n7018 GND.n5015 9.3005
R26283 GND.n6529 GND.n5016 9.3005
R26284 GND.n7008 GND.n5034 9.3005
R26285 GND.n7007 GND.n5035 9.3005
R26286 GND.n7006 GND.n5036 9.3005
R26287 GND.n6536 GND.n5037 9.3005
R26288 GND.n6996 GND.n5055 9.3005
R26289 GND.n6995 GND.n5056 9.3005
R26290 GND.n6994 GND.n5057 9.3005
R26291 GND.n6543 GND.n5058 9.3005
R26292 GND.n6984 GND.n5076 9.3005
R26293 GND.n6983 GND.n5077 9.3005
R26294 GND.n6982 GND.n5078 9.3005
R26295 GND.n6550 GND.n5079 9.3005
R26296 GND.n6972 GND.n5097 9.3005
R26297 GND.n6971 GND.n5098 9.3005
R26298 GND.n6970 GND.n5099 9.3005
R26299 GND.n6557 GND.n5100 9.3005
R26300 GND.n6960 GND.n5118 9.3005
R26301 GND.n6959 GND.n5119 9.3005
R26302 GND.n6958 GND.n5120 9.3005
R26303 GND.n6564 GND.n5121 9.3005
R26304 GND.n6948 GND.n5139 9.3005
R26305 GND.n6947 GND.n5140 9.3005
R26306 GND.n6946 GND.n5141 9.3005
R26307 GND.n6571 GND.n5142 9.3005
R26308 GND.n6936 GND.n5160 9.3005
R26309 GND.n6935 GND.n5161 9.3005
R26310 GND.n6934 GND.n5162 9.3005
R26311 GND.n6572 GND.n5163 9.3005
R26312 GND.n6924 GND.n5179 9.3005
R26313 GND.n6923 GND.n5180 9.3005
R26314 GND.n6922 GND.n5181 9.3005
R26315 GND.n6774 GND.n5182 9.3005
R26316 GND.n6775 GND.n5284 9.3005
R26317 GND.n6781 GND.n5283 9.3005
R26318 GND.n6783 GND.n6782 9.3005
R26319 GND.n5280 GND.n5279 9.3005
R26320 GND.n6792 GND.n6791 9.3005
R26321 GND.n6793 GND.n133 9.3005
R26322 GND.n10301 GND.n134 9.3005
R26323 GND.n10300 GND.n135 9.3005
R26324 GND.n10299 GND.n136 9.3005
R26325 GND.n6796 GND.n137 9.3005
R26326 GND.n10289 GND.n154 9.3005
R26327 GND.n10288 GND.n155 9.3005
R26328 GND.n10287 GND.n156 9.3005
R26329 GND.n6803 GND.n157 9.3005
R26330 GND.n10277 GND.n175 9.3005
R26331 GND.n10276 GND.n176 9.3005
R26332 GND.n10275 GND.n177 9.3005
R26333 GND.n6810 GND.n178 9.3005
R26334 GND.n10265 GND.n196 9.3005
R26335 GND.n10264 GND.n197 9.3005
R26336 GND.n10263 GND.n198 9.3005
R26337 GND.n6817 GND.n199 9.3005
R26338 GND.n10253 GND.n217 9.3005
R26339 GND.n10252 GND.n218 9.3005
R26340 GND.n10251 GND.n219 9.3005
R26341 GND.n6824 GND.n220 9.3005
R26342 GND.n10241 GND.n238 9.3005
R26343 GND.n10240 GND.n239 9.3005
R26344 GND.n10239 GND.n240 9.3005
R26345 GND.n6830 GND.n241 9.3005
R26346 GND.n10229 GND.n258 9.3005
R26347 GND.n10228 GND.n259 9.3005
R26348 GND.n10227 GND.n260 9.3005
R26349 GND.n9739 GND.n261 9.3005
R26350 GND.n10217 GND.n279 9.3005
R26351 GND.n10216 GND.n280 9.3005
R26352 GND.n10215 GND.n281 9.3005
R26353 GND.n9754 GND.n282 9.3005
R26354 GND.n10205 GND.n300 9.3005
R26355 GND.n10204 GND.n301 9.3005
R26356 GND.n10203 GND.n302 9.3005
R26357 GND.n9769 GND.n303 9.3005
R26358 GND.n10193 GND.n321 9.3005
R26359 GND.n10192 GND.n322 9.3005
R26360 GND.n10191 GND.n323 9.3005
R26361 GND.n9784 GND.n324 9.3005
R26362 GND.n10181 GND.n342 9.3005
R26363 GND.n10180 GND.n343 9.3005
R26364 GND.n10179 GND.n344 9.3005
R26365 GND.n10108 GND.n345 9.3005
R26366 GND.n10169 GND.n363 9.3005
R26367 GND.n10168 GND.n364 9.3005
R26368 GND.n10167 GND.n365 9.3005
R26369 GND.n10115 GND.n366 9.3005
R26370 GND.n10157 GND.n382 9.3005
R26371 GND.n10156 GND.n383 9.3005
R26372 GND.n10155 GND.n384 9.3005
R26373 GND.n10122 GND.n385 9.3005
R26374 GND.n10145 GND.n401 9.3005
R26375 GND.n10144 GND.n402 9.3005
R26376 GND.n10143 GND.n403 9.3005
R26377 GND.n419 GND.n404 9.3005
R26378 GND.n10133 GND.n10132 9.3005
R26379 GND.n4890 GND.n4888 9.3005
R26380 GND.n7088 GND.n7087 9.3005
R26381 GND.n7086 GND.n4891 9.3005
R26382 GND.n5355 GND.n4893 9.3005
R26383 GND.n5354 GND.n5353 9.3005
R26384 GND.n5361 GND.n5351 9.3005
R26385 GND.n6475 GND.n5362 9.3005
R26386 GND.n6476 GND.n4930 9.3005
R26387 GND.n6477 GND.n4931 9.3005
R26388 GND.n5346 GND.n4932 9.3005
R26389 GND.n6489 GND.n5347 9.3005
R26390 GND.n6490 GND.n4951 9.3005
R26391 GND.n6491 GND.n4952 9.3005
R26392 GND.n5341 GND.n4953 9.3005
R26393 GND.n6503 GND.n5342 9.3005
R26394 GND.n6504 GND.n4972 9.3005
R26395 GND.n6505 GND.n4973 9.3005
R26396 GND.n5336 GND.n4974 9.3005
R26397 GND.n6518 GND.n5337 9.3005
R26398 GND.n6519 GND.n4993 9.3005
R26399 GND.n6520 GND.n4994 9.3005
R26400 GND.n6521 GND.n4995 9.3005
R26401 GND.n6667 GND.n6522 9.3005
R26402 GND.n6666 GND.n5013 9.3005
R26403 GND.n6665 GND.n5014 9.3005
R26404 GND.n6523 GND.n5015 9.3005
R26405 GND.n6655 GND.n6529 9.3005
R26406 GND.n6654 GND.n5034 9.3005
R26407 GND.n6653 GND.n5035 9.3005
R26408 GND.n6530 GND.n5036 9.3005
R26409 GND.n6643 GND.n6536 9.3005
R26410 GND.n6642 GND.n5055 9.3005
R26411 GND.n6641 GND.n5056 9.3005
R26412 GND.n6537 GND.n5057 9.3005
R26413 GND.n6631 GND.n6543 9.3005
R26414 GND.n6630 GND.n5076 9.3005
R26415 GND.n6629 GND.n5077 9.3005
R26416 GND.n6544 GND.n5078 9.3005
R26417 GND.n6619 GND.n6550 9.3005
R26418 GND.n6618 GND.n5097 9.3005
R26419 GND.n6617 GND.n5098 9.3005
R26420 GND.n6551 GND.n5099 9.3005
R26421 GND.n6607 GND.n6557 9.3005
R26422 GND.n6606 GND.n5118 9.3005
R26423 GND.n6605 GND.n5119 9.3005
R26424 GND.n6558 GND.n5120 9.3005
R26425 GND.n6595 GND.n6564 9.3005
R26426 GND.n6594 GND.n5139 9.3005
R26427 GND.n6593 GND.n5140 9.3005
R26428 GND.n6565 GND.n5141 9.3005
R26429 GND.n6583 GND.n6571 9.3005
R26430 GND.n6582 GND.n5160 9.3005
R26431 GND.n6581 GND.n5161 9.3005
R26432 GND.n6574 GND.n5162 9.3005
R26433 GND.n6573 GND.n6572 9.3005
R26434 GND.n5287 GND.n5179 9.3005
R26435 GND.n6771 GND.n5180 9.3005
R26436 GND.n6772 GND.n5181 9.3005
R26437 GND.n6774 GND.n6773 9.3005
R26438 GND.n6776 GND.n6775 9.3005
R26439 GND.n5283 GND.n5282 9.3005
R26440 GND.n6784 GND.n6783 9.3005
R26441 GND.n6785 GND.n5279 9.3005
R26442 GND.n6792 GND.n5278 9.3005
R26443 GND.n6794 GND.n6793 9.3005
R26444 GND.n6795 GND.n134 9.3005
R26445 GND.n6893 GND.n135 9.3005
R26446 GND.n6892 GND.n136 9.3005
R26447 GND.n6891 GND.n6796 9.3005
R26448 GND.n6797 GND.n154 9.3005
R26449 GND.n6881 GND.n155 9.3005
R26450 GND.n6880 GND.n156 9.3005
R26451 GND.n6879 GND.n6803 9.3005
R26452 GND.n6804 GND.n175 9.3005
R26453 GND.n6869 GND.n176 9.3005
R26454 GND.n6868 GND.n177 9.3005
R26455 GND.n6867 GND.n6810 9.3005
R26456 GND.n6811 GND.n196 9.3005
R26457 GND.n6857 GND.n197 9.3005
R26458 GND.n6856 GND.n198 9.3005
R26459 GND.n6855 GND.n6817 9.3005
R26460 GND.n6818 GND.n217 9.3005
R26461 GND.n6845 GND.n218 9.3005
R26462 GND.n6844 GND.n219 9.3005
R26463 GND.n6843 GND.n6824 9.3005
R26464 GND.n6825 GND.n238 9.3005
R26465 GND.n6833 GND.n239 9.3005
R26466 GND.n6832 GND.n240 9.3005
R26467 GND.n6831 GND.n6830 9.3005
R26468 GND.n437 GND.n258 9.3005
R26469 GND.n9737 GND.n259 9.3005
R26470 GND.n9738 GND.n260 9.3005
R26471 GND.n9740 GND.n9739 9.3005
R26472 GND.n433 GND.n279 9.3005
R26473 GND.n9752 GND.n280 9.3005
R26474 GND.n9753 GND.n281 9.3005
R26475 GND.n9755 GND.n9754 9.3005
R26476 GND.n429 GND.n300 9.3005
R26477 GND.n9767 GND.n301 9.3005
R26478 GND.n9768 GND.n302 9.3005
R26479 GND.n9770 GND.n9769 9.3005
R26480 GND.n425 GND.n321 9.3005
R26481 GND.n9782 GND.n322 9.3005
R26482 GND.n9783 GND.n323 9.3005
R26483 GND.n9785 GND.n9784 9.3005
R26484 GND.n421 GND.n342 9.3005
R26485 GND.n10106 GND.n343 9.3005
R26486 GND.n10107 GND.n344 9.3005
R26487 GND.n10110 GND.n10108 9.3005
R26488 GND.n10111 GND.n363 9.3005
R26489 GND.n10113 GND.n364 9.3005
R26490 GND.n10114 GND.n365 9.3005
R26491 GND.n10117 GND.n10115 9.3005
R26492 GND.n10118 GND.n382 9.3005
R26493 GND.n10120 GND.n383 9.3005
R26494 GND.n10121 GND.n384 9.3005
R26495 GND.n10124 GND.n10122 9.3005
R26496 GND.n10125 GND.n401 9.3005
R26497 GND.n10127 GND.n402 9.3005
R26498 GND.n10128 GND.n403 9.3005
R26499 GND.n10130 GND.n419 9.3005
R26500 GND.n10132 GND.n10131 9.3005
R26501 GND.n4892 GND.n4890 9.3005
R26502 GND.n5460 GND.n5366 9.3005
R26503 GND.n5456 GND.n5453 9.3005
R26504 GND.n5452 GND.n5367 9.3005
R26505 GND.n5451 GND.n5450 9.3005
R26506 GND.n5447 GND.n5368 9.3005
R26507 GND.n5446 GND.n5443 9.3005
R26508 GND.n5442 GND.n5369 9.3005
R26509 GND.n5441 GND.n5440 9.3005
R26510 GND.n5437 GND.n5370 9.3005
R26511 GND.n5436 GND.n5433 9.3005
R26512 GND.n5432 GND.n5371 9.3005
R26513 GND.n5431 GND.n5430 9.3005
R26514 GND.n5427 GND.n5372 9.3005
R26515 GND.n5423 GND.n5420 9.3005
R26516 GND.n5419 GND.n5373 9.3005
R26517 GND.n5418 GND.n5417 9.3005
R26518 GND.n5414 GND.n5374 9.3005
R26519 GND.n5413 GND.n5410 9.3005
R26520 GND.n5409 GND.n5375 9.3005
R26521 GND.n5408 GND.n5407 9.3005
R26522 GND.n5404 GND.n5376 9.3005
R26523 GND.n5403 GND.n5400 9.3005
R26524 GND.n5399 GND.n5377 9.3005
R26525 GND.n5398 GND.n5397 9.3005
R26526 GND.n5394 GND.n5378 9.3005
R26527 GND.n5389 GND.n5379 9.3005
R26528 GND.n5388 GND.n5387 9.3005
R26529 GND.n5384 GND.n5383 9.3005
R26530 GND.n5382 GND.n4837 9.3005
R26531 GND.n7186 GND.n4836 9.3005
R26532 GND.n7128 GND.n4833 9.3005
R26533 GND.n7132 GND.n7129 9.3005
R26534 GND.n7133 GND.n7127 9.3005
R26535 GND.n7136 GND.n7126 9.3005
R26536 GND.n7137 GND.n7125 9.3005
R26537 GND.n7140 GND.n7121 9.3005
R26538 GND.n7141 GND.n7120 9.3005
R26539 GND.n7144 GND.n7119 9.3005
R26540 GND.n7145 GND.n7118 9.3005
R26541 GND.n7148 GND.n7117 9.3005
R26542 GND.n7149 GND.n7116 9.3005
R26543 GND.n7152 GND.n7115 9.3005
R26544 GND.n7153 GND.n7114 9.3005
R26545 GND.n7156 GND.n7113 9.3005
R26546 GND.n7157 GND.n7112 9.3005
R26547 GND.n7160 GND.n7111 9.3005
R26548 GND.n7162 GND.n7110 9.3005
R26549 GND.n7164 GND.n7105 9.3005
R26550 GND.n7167 GND.n7104 9.3005
R26551 GND.n7168 GND.n7103 9.3005
R26552 GND.n7171 GND.n7102 9.3005
R26553 GND.n7172 GND.n7101 9.3005
R26554 GND.n7175 GND.n7100 9.3005
R26555 GND.n7177 GND.n7099 9.3005
R26556 GND.n7178 GND.n7098 9.3005
R26557 GND.n7179 GND.n7097 9.3005
R26558 GND.n7180 GND.n7096 9.3005
R26559 GND.n7163 GND.n7107 9.3005
R26560 GND.n5393 GND.n5390 9.3005
R26561 GND.n5462 GND.n5461 9.3005
R26562 GND.n7093 GND.n4879 9.3005
R26563 GND.n4914 GND.n4880 9.3005
R26564 GND.n4917 GND.n4916 9.3005
R26565 GND.n4918 GND.n4913 9.3005
R26566 GND.n7074 GND.n4919 9.3005
R26567 GND.n7073 GND.n4920 9.3005
R26568 GND.n7072 GND.n4921 9.3005
R26569 GND.n4940 GND.n4922 9.3005
R26570 GND.n7062 GND.n4941 9.3005
R26571 GND.n7061 GND.n4942 9.3005
R26572 GND.n7060 GND.n4943 9.3005
R26573 GND.n4961 GND.n4944 9.3005
R26574 GND.n7050 GND.n4962 9.3005
R26575 GND.n7049 GND.n4963 9.3005
R26576 GND.n7048 GND.n4964 9.3005
R26577 GND.n4982 GND.n4965 9.3005
R26578 GND.n7038 GND.n4983 9.3005
R26579 GND.n7037 GND.n4984 9.3005
R26580 GND.n7036 GND.n4985 9.3005
R26581 GND.n5002 GND.n4986 9.3005
R26582 GND.n7026 GND.n5003 9.3005
R26583 GND.n7025 GND.n5004 9.3005
R26584 GND.n7024 GND.n5005 9.3005
R26585 GND.n5023 GND.n5006 9.3005
R26586 GND.n7014 GND.n5024 9.3005
R26587 GND.n7013 GND.n5025 9.3005
R26588 GND.n7012 GND.n5026 9.3005
R26589 GND.n5044 GND.n5027 9.3005
R26590 GND.n7002 GND.n5045 9.3005
R26591 GND.n7001 GND.n5046 9.3005
R26592 GND.n7000 GND.n5047 9.3005
R26593 GND.n5065 GND.n5048 9.3005
R26594 GND.n6990 GND.n5066 9.3005
R26595 GND.n6989 GND.n5067 9.3005
R26596 GND.n6988 GND.n5068 9.3005
R26597 GND.n5086 GND.n5069 9.3005
R26598 GND.n6978 GND.n5087 9.3005
R26599 GND.n6977 GND.n5088 9.3005
R26600 GND.n6976 GND.n5089 9.3005
R26601 GND.n5107 GND.n5090 9.3005
R26602 GND.n6966 GND.n5108 9.3005
R26603 GND.n6965 GND.n5109 9.3005
R26604 GND.n6964 GND.n5110 9.3005
R26605 GND.n5128 GND.n5111 9.3005
R26606 GND.n6954 GND.n5129 9.3005
R26607 GND.n6953 GND.n5130 9.3005
R26608 GND.n6952 GND.n5131 9.3005
R26609 GND.n5149 GND.n5132 9.3005
R26610 GND.n6942 GND.n5150 9.3005
R26611 GND.n6941 GND.n5151 9.3005
R26612 GND.n6940 GND.n5152 9.3005
R26613 GND.n5170 GND.n5153 9.3005
R26614 GND.n6930 GND.n5171 9.3005
R26615 GND.n6929 GND.n5172 9.3005
R26616 GND.n6928 GND.n117 9.3005
R26617 GND.n124 GND.n116 9.3005
R26618 GND.n10295 GND.n144 9.3005
R26619 GND.n10294 GND.n145 9.3005
R26620 GND.n10293 GND.n146 9.3005
R26621 GND.n164 GND.n147 9.3005
R26622 GND.n10283 GND.n165 9.3005
R26623 GND.n10282 GND.n166 9.3005
R26624 GND.n10281 GND.n167 9.3005
R26625 GND.n185 GND.n168 9.3005
R26626 GND.n10271 GND.n186 9.3005
R26627 GND.n10270 GND.n187 9.3005
R26628 GND.n10269 GND.n188 9.3005
R26629 GND.n206 GND.n189 9.3005
R26630 GND.n10259 GND.n207 9.3005
R26631 GND.n10258 GND.n208 9.3005
R26632 GND.n10257 GND.n209 9.3005
R26633 GND.n227 GND.n210 9.3005
R26634 GND.n10247 GND.n228 9.3005
R26635 GND.n10246 GND.n229 9.3005
R26636 GND.n10245 GND.n230 9.3005
R26637 GND.n248 GND.n231 9.3005
R26638 GND.n10235 GND.n249 9.3005
R26639 GND.n10234 GND.n250 9.3005
R26640 GND.n10233 GND.n251 9.3005
R26641 GND.n268 GND.n252 9.3005
R26642 GND.n10223 GND.n269 9.3005
R26643 GND.n10222 GND.n270 9.3005
R26644 GND.n10221 GND.n271 9.3005
R26645 GND.n289 GND.n272 9.3005
R26646 GND.n10211 GND.n290 9.3005
R26647 GND.n10210 GND.n291 9.3005
R26648 GND.n10209 GND.n292 9.3005
R26649 GND.n310 GND.n293 9.3005
R26650 GND.n10199 GND.n311 9.3005
R26651 GND.n10198 GND.n312 9.3005
R26652 GND.n10197 GND.n313 9.3005
R26653 GND.n331 GND.n314 9.3005
R26654 GND.n10187 GND.n332 9.3005
R26655 GND.n10186 GND.n333 9.3005
R26656 GND.n10185 GND.n334 9.3005
R26657 GND.n352 GND.n335 9.3005
R26658 GND.n10175 GND.n353 9.3005
R26659 GND.n10174 GND.n354 9.3005
R26660 GND.n10173 GND.n355 9.3005
R26661 GND.n372 GND.n356 9.3005
R26662 GND.n10163 GND.n373 9.3005
R26663 GND.n10162 GND.n374 9.3005
R26664 GND.n10161 GND.n375 9.3005
R26665 GND.n391 GND.n376 9.3005
R26666 GND.n10151 GND.n392 9.3005
R26667 GND.n10150 GND.n393 9.3005
R26668 GND.n10149 GND.n394 9.3005
R26669 GND.n410 GND.n395 9.3005
R26670 GND.n10139 GND.n411 9.3005
R26671 GND.n10138 GND.n412 9.3005
R26672 GND.n10137 GND.n413 9.3005
R26673 GND.n7095 GND.n7094 9.3005
R26674 GND.n10306 GND.n121 9.3005
R26675 GND.n10306 GND.n10305 9.3005
R26676 GND.n3337 GND.n3335 9.3005
R26677 GND.n3526 GND.n3338 9.3005
R26678 GND.n3525 GND.n3339 9.3005
R26679 GND.n3524 GND.n3340 9.3005
R26680 GND.n3343 GND.n3341 9.3005
R26681 GND.n3520 GND.n3344 9.3005
R26682 GND.n3519 GND.n3345 9.3005
R26683 GND.n3518 GND.n3346 9.3005
R26684 GND.n3349 GND.n3347 9.3005
R26685 GND.n3514 GND.n3350 9.3005
R26686 GND.n3513 GND.n3351 9.3005
R26687 GND.n3512 GND.n3352 9.3005
R26688 GND.n3355 GND.n3353 9.3005
R26689 GND.n3508 GND.n3356 9.3005
R26690 GND.n3507 GND.n3357 9.3005
R26691 GND.n3506 GND.n3358 9.3005
R26692 GND.n3361 GND.n3359 9.3005
R26693 GND.n3502 GND.n3362 9.3005
R26694 GND.n3501 GND.n3363 9.3005
R26695 GND.n3500 GND.n3364 9.3005
R26696 GND.n3367 GND.n3365 9.3005
R26697 GND.n3496 GND.n3368 9.3005
R26698 GND.n3495 GND.n3369 9.3005
R26699 GND.n3494 GND.n3370 9.3005
R26700 GND.n3373 GND.n3371 9.3005
R26701 GND.n3490 GND.n3374 9.3005
R26702 GND.n3489 GND.n3375 9.3005
R26703 GND.n3488 GND.n3376 9.3005
R26704 GND.n3379 GND.n3377 9.3005
R26705 GND.n3484 GND.n3380 9.3005
R26706 GND.n3483 GND.n3381 9.3005
R26707 GND.n3482 GND.n3382 9.3005
R26708 GND.n3385 GND.n3383 9.3005
R26709 GND.n3478 GND.n3386 9.3005
R26710 GND.n3477 GND.n3387 9.3005
R26711 GND.n3476 GND.n3388 9.3005
R26712 GND.n3391 GND.n3389 9.3005
R26713 GND.n3470 GND.n3392 9.3005
R26714 GND.n3469 GND.n3393 9.3005
R26715 GND.n3468 GND.n3394 9.3005
R26716 GND.n3397 GND.n3395 9.3005
R26717 GND.n3464 GND.n3398 9.3005
R26718 GND.n3463 GND.n3399 9.3005
R26719 GND.n3462 GND.n3400 9.3005
R26720 GND.n3403 GND.n3401 9.3005
R26721 GND.n3458 GND.n3404 9.3005
R26722 GND.n3457 GND.n3405 9.3005
R26723 GND.n3456 GND.n3406 9.3005
R26724 GND.n3409 GND.n3407 9.3005
R26725 GND.n3452 GND.n3410 9.3005
R26726 GND.n3451 GND.n3411 9.3005
R26727 GND.n3450 GND.n3412 9.3005
R26728 GND.n3415 GND.n3413 9.3005
R26729 GND.n3446 GND.n3416 9.3005
R26730 GND.n3445 GND.n3417 9.3005
R26731 GND.n3444 GND.n3418 9.3005
R26732 GND.n3421 GND.n3419 9.3005
R26733 GND.n3440 GND.n3422 9.3005
R26734 GND.n3439 GND.n3423 9.3005
R26735 GND.n3438 GND.n3424 9.3005
R26736 GND.n3427 GND.n3425 9.3005
R26737 GND.n3432 GND.n3428 9.3005
R26738 GND.n3431 GND.n3430 9.3005
R26739 GND.n3429 GND.n1941 9.3005
R26740 GND.n7908 GND.n1942 9.3005
R26741 GND.n7907 GND.n1943 9.3005
R26742 GND.n7906 GND.n1944 9.3005
R26743 GND.n1958 GND.n1945 9.3005
R26744 GND.n7895 GND.n1959 9.3005
R26745 GND.n7894 GND.n1960 9.3005
R26746 GND.n7893 GND.n1961 9.3005
R26747 GND.n1975 GND.n1962 9.3005
R26748 GND.n7881 GND.n1976 9.3005
R26749 GND.n7880 GND.n1977 9.3005
R26750 GND.n7879 GND.n1978 9.3005
R26751 GND.n1993 GND.n1979 9.3005
R26752 GND.n7867 GND.n1994 9.3005
R26753 GND.n7866 GND.n1995 9.3005
R26754 GND.n7865 GND.n1996 9.3005
R26755 GND.n2011 GND.n1997 9.3005
R26756 GND.n7853 GND.n2012 9.3005
R26757 GND.n7852 GND.n2013 9.3005
R26758 GND.n7851 GND.n2014 9.3005
R26759 GND.n2029 GND.n2015 9.3005
R26760 GND.n7839 GND.n2030 9.3005
R26761 GND.n7838 GND.n2031 9.3005
R26762 GND.n7837 GND.n2032 9.3005
R26763 GND.n2047 GND.n2033 9.3005
R26764 GND.n7825 GND.n2048 9.3005
R26765 GND.n7824 GND.n2049 9.3005
R26766 GND.n7823 GND.n2050 9.3005
R26767 GND.n2065 GND.n2051 9.3005
R26768 GND.n7811 GND.n2066 9.3005
R26769 GND.n7810 GND.n2067 9.3005
R26770 GND.n7809 GND.n2068 9.3005
R26771 GND.n2083 GND.n2069 9.3005
R26772 GND.n7797 GND.n2084 9.3005
R26773 GND.n7796 GND.n2085 9.3005
R26774 GND.n7795 GND.n2086 9.3005
R26775 GND.n2101 GND.n2087 9.3005
R26776 GND.n7783 GND.n2102 9.3005
R26777 GND.n7782 GND.n2103 9.3005
R26778 GND.n7781 GND.n2104 9.3005
R26779 GND.n2320 GND.n2105 9.3005
R26780 GND.n2321 GND.n2319 9.3005
R26781 GND.n7764 GND.n2322 9.3005
R26782 GND.n7763 GND.n2323 9.3005
R26783 GND.n7762 GND.n2324 9.3005
R26784 GND.n3888 GND.n2325 9.3005
R26785 GND.n7695 GND.n3889 9.3005
R26786 GND.n7694 GND.n3890 9.3005
R26787 GND.n7693 GND.n3891 9.3005
R26788 GND.n3907 GND.n3892 9.3005
R26789 GND.n7684 GND.n3908 9.3005
R26790 GND.n7683 GND.n3909 9.3005
R26791 GND.n7682 GND.n3910 9.3005
R26792 GND.n3927 GND.n3911 9.3005
R26793 GND.n7672 GND.n3928 9.3005
R26794 GND.n7671 GND.n3929 9.3005
R26795 GND.n7670 GND.n3930 9.3005
R26796 GND.n3957 GND.n3931 9.3005
R26797 GND.n3958 GND.n3956 9.3005
R26798 GND.n7653 GND.n3959 9.3005
R26799 GND.n7652 GND.n3960 9.3005
R26800 GND.n7651 GND.n3961 9.3005
R26801 GND.n3991 GND.n3962 9.3005
R26802 GND.n7641 GND.n3992 9.3005
R26803 GND.n7640 GND.n3993 9.3005
R26804 GND.n7639 GND.n3994 9.3005
R26805 GND.n4011 GND.n3995 9.3005
R26806 GND.n7629 GND.n4012 9.3005
R26807 GND.n7628 GND.n4013 9.3005
R26808 GND.n7627 GND.n4014 9.3005
R26809 GND.n4031 GND.n4015 9.3005
R26810 GND.n7617 GND.n4032 9.3005
R26811 GND.n7616 GND.n4033 9.3005
R26812 GND.n7615 GND.n4034 9.3005
R26813 GND.n4062 GND.n4035 9.3005
R26814 GND.n4063 GND.n4061 9.3005
R26815 GND.n7598 GND.n4064 9.3005
R26816 GND.n7597 GND.n4065 9.3005
R26817 GND.n7596 GND.n4066 9.3005
R26818 GND.n4096 GND.n4067 9.3005
R26819 GND.n7586 GND.n4097 9.3005
R26820 GND.n7585 GND.n4098 9.3005
R26821 GND.n7584 GND.n4099 9.3005
R26822 GND.n4116 GND.n4100 9.3005
R26823 GND.n7574 GND.n4117 9.3005
R26824 GND.n7573 GND.n4118 9.3005
R26825 GND.n7572 GND.n4119 9.3005
R26826 GND.n4136 GND.n4120 9.3005
R26827 GND.n7562 GND.n4137 9.3005
R26828 GND.n7561 GND.n4138 9.3005
R26829 GND.n7560 GND.n4139 9.3005
R26830 GND.n4167 GND.n4140 9.3005
R26831 GND.n4168 GND.n4166 9.3005
R26832 GND.n7543 GND.n4169 9.3005
R26833 GND.n7542 GND.n4170 9.3005
R26834 GND.n7541 GND.n4171 9.3005
R26835 GND.n4200 GND.n4172 9.3005
R26836 GND.n7531 GND.n4201 9.3005
R26837 GND.n7530 GND.n4202 9.3005
R26838 GND.n7529 GND.n4203 9.3005
R26839 GND.n4220 GND.n4204 9.3005
R26840 GND.n7519 GND.n4221 9.3005
R26841 GND.n7518 GND.n4222 9.3005
R26842 GND.n7517 GND.n4223 9.3005
R26843 GND.n4239 GND.n4224 9.3005
R26844 GND.n7507 GND.n4240 9.3005
R26845 GND.n7506 GND.n4241 9.3005
R26846 GND.n7505 GND.n4242 9.3005
R26847 GND.n4270 GND.n4243 9.3005
R26848 GND.n4271 GND.n4269 9.3005
R26849 GND.n7488 GND.n4272 9.3005
R26850 GND.n7487 GND.n4273 9.3005
R26851 GND.n7486 GND.n4274 9.3005
R26852 GND.n4303 GND.n4275 9.3005
R26853 GND.n7476 GND.n4304 9.3005
R26854 GND.n7475 GND.n4305 9.3005
R26855 GND.n7474 GND.n4306 9.3005
R26856 GND.n4323 GND.n4307 9.3005
R26857 GND.n7464 GND.n4324 9.3005
R26858 GND.n7463 GND.n4325 9.3005
R26859 GND.n7462 GND.n4326 9.3005
R26860 GND.n4343 GND.n4327 9.3005
R26861 GND.n7452 GND.n4344 9.3005
R26862 GND.n7451 GND.n4345 9.3005
R26863 GND.n7450 GND.n4346 9.3005
R26864 GND.n4374 GND.n4347 9.3005
R26865 GND.n4375 GND.n4373 9.3005
R26866 GND.n7433 GND.n4376 9.3005
R26867 GND.n7432 GND.n4377 9.3005
R26868 GND.n7431 GND.n4378 9.3005
R26869 GND.n4408 GND.n4379 9.3005
R26870 GND.n7421 GND.n4409 9.3005
R26871 GND.n7420 GND.n4410 9.3005
R26872 GND.n7419 GND.n4411 9.3005
R26873 GND.n4440 GND.n4412 9.3005
R26874 GND.n4441 GND.n4439 9.3005
R26875 GND.n7405 GND.n4442 9.3005
R26876 GND.n7404 GND.n4443 9.3005
R26877 GND.n7403 GND.n4444 9.3005
R26878 GND.n4459 GND.n4445 9.3005
R26879 GND.n7391 GND.n4460 9.3005
R26880 GND.n7390 GND.n4461 9.3005
R26881 GND.n7389 GND.n4462 9.3005
R26882 GND.n4477 GND.n4463 9.3005
R26883 GND.n7377 GND.n4478 9.3005
R26884 GND.n7376 GND.n4479 9.3005
R26885 GND.n7375 GND.n4480 9.3005
R26886 GND.n4495 GND.n4481 9.3005
R26887 GND.n7363 GND.n4496 9.3005
R26888 GND.n7362 GND.n4497 9.3005
R26889 GND.n7361 GND.n4498 9.3005
R26890 GND.n4513 GND.n4499 9.3005
R26891 GND.n7349 GND.n4514 9.3005
R26892 GND.n7348 GND.n4515 9.3005
R26893 GND.n7347 GND.n4516 9.3005
R26894 GND.n4531 GND.n4517 9.3005
R26895 GND.n7335 GND.n4532 9.3005
R26896 GND.n7334 GND.n4533 9.3005
R26897 GND.n7333 GND.n4534 9.3005
R26898 GND.n4562 GND.n4535 9.3005
R26899 GND.n4563 GND.n4561 9.3005
R26900 GND.n7316 GND.n4564 9.3005
R26901 GND.n7315 GND.n4565 9.3005
R26902 GND.n7314 GND.n4566 9.3005
R26903 GND.n4581 GND.n4567 9.3005
R26904 GND.n7302 GND.n4582 9.3005
R26905 GND.n7301 GND.n4583 9.3005
R26906 GND.n7300 GND.n4584 9.3005
R26907 GND.n4599 GND.n4585 9.3005
R26908 GND.n7288 GND.n4600 9.3005
R26909 GND.n7287 GND.n4601 9.3005
R26910 GND.n7286 GND.n4602 9.3005
R26911 GND.n4616 GND.n4603 9.3005
R26912 GND.n7274 GND.n4617 9.3005
R26913 GND.n7273 GND.n4618 9.3005
R26914 GND.n7272 GND.n4619 9.3005
R26915 GND.n4693 GND.n4620 9.3005
R26916 GND.n4694 GND.n4692 9.3005
R26917 GND.n7255 GND.n4695 9.3005
R26918 GND.n7254 GND.n4696 9.3005
R26919 GND.n7253 GND.n4697 9.3005
R26920 GND.n6394 GND.n4698 9.3005
R26921 GND.n6398 GND.n6395 9.3005
R26922 GND.n6397 GND.n6396 9.3005
R26923 GND.n6392 GND.n6391 9.3005
R26924 GND.n6406 GND.n6405 9.3005
R26925 GND.n6407 GND.n6390 9.3005
R26926 GND.n6412 GND.n6408 9.3005
R26927 GND.n6411 GND.n6410 9.3005
R26928 GND.n6409 GND.n4899 9.3005
R26929 GND.n7081 GND.n4900 9.3005
R26930 GND.n7080 GND.n4901 9.3005
R26931 GND.n7079 GND.n4902 9.3005
R26932 GND.n6433 GND.n4903 9.3005
R26933 GND.n6470 GND.n6434 9.3005
R26934 GND.n6469 GND.n6435 9.3005
R26935 GND.n6468 GND.n6436 9.3005
R26936 GND.n6439 GND.n6437 9.3005
R26937 GND.n6464 GND.n6440 9.3005
R26938 GND.n6463 GND.n6441 9.3005
R26939 GND.n6462 GND.n6442 9.3005
R26940 GND.n6445 GND.n6443 9.3005
R26941 GND.n6458 GND.n6446 9.3005
R26942 GND.n6457 GND.n6447 9.3005
R26943 GND.n6456 GND.n6448 9.3005
R26944 GND.n6450 GND.n6449 9.3005
R26945 GND.n6452 GND.n6451 9.3005
R26946 GND.n5328 GND.n5327 9.3005
R26947 GND.n6679 GND.n6678 9.3005
R26948 GND.n6680 GND.n5326 9.3005
R26949 GND.n6682 GND.n6681 9.3005
R26950 GND.n5324 GND.n5323 9.3005
R26951 GND.n6687 GND.n6686 9.3005
R26952 GND.n6688 GND.n5322 9.3005
R26953 GND.n6690 GND.n6689 9.3005
R26954 GND.n5320 GND.n5319 9.3005
R26955 GND.n6695 GND.n6694 9.3005
R26956 GND.n6696 GND.n5318 9.3005
R26957 GND.n6698 GND.n6697 9.3005
R26958 GND.n5316 GND.n5315 9.3005
R26959 GND.n6703 GND.n6702 9.3005
R26960 GND.n6704 GND.n5314 9.3005
R26961 GND.n6706 GND.n6705 9.3005
R26962 GND.n5312 GND.n5311 9.3005
R26963 GND.n6711 GND.n6710 9.3005
R26964 GND.n6712 GND.n5310 9.3005
R26965 GND.n6714 GND.n6713 9.3005
R26966 GND.n5308 GND.n5307 9.3005
R26967 GND.n6719 GND.n6718 9.3005
R26968 GND.n6720 GND.n5306 9.3005
R26969 GND.n6722 GND.n6721 9.3005
R26970 GND.n5304 GND.n5303 9.3005
R26971 GND.n6727 GND.n6726 9.3005
R26972 GND.n6728 GND.n5302 9.3005
R26973 GND.n6730 GND.n6729 9.3005
R26974 GND.n5300 GND.n5299 9.3005
R26975 GND.n6735 GND.n6734 9.3005
R26976 GND.n6736 GND.n5298 9.3005
R26977 GND.n6738 GND.n6737 9.3005
R26978 GND.n5296 GND.n5295 9.3005
R26979 GND.n6743 GND.n6742 9.3005
R26980 GND.n6744 GND.n5294 9.3005
R26981 GND.n6751 GND.n6745 9.3005
R26982 GND.n6750 GND.n6746 9.3005
R26983 GND.n5263 GND.n5201 9.3005
R26984 GND.n5262 GND.n5202 9.3005
R26985 GND.n5205 GND.n5203 9.3005
R26986 GND.n5258 GND.n5206 9.3005
R26987 GND.n5257 GND.n5207 9.3005
R26988 GND.n5256 GND.n5208 9.3005
R26989 GND.n5211 GND.n5209 9.3005
R26990 GND.n5252 GND.n5212 9.3005
R26991 GND.n5251 GND.n5213 9.3005
R26992 GND.n5250 GND.n5214 9.3005
R26993 GND.n5217 GND.n5215 9.3005
R26994 GND.n5246 GND.n5218 9.3005
R26995 GND.n5245 GND.n5219 9.3005
R26996 GND.n5244 GND.n5220 9.3005
R26997 GND.n5223 GND.n5221 9.3005
R26998 GND.n5240 GND.n5224 9.3005
R26999 GND.n5239 GND.n5225 9.3005
R27000 GND.n5238 GND.n5226 9.3005
R27001 GND.n5229 GND.n5227 9.3005
R27002 GND.n5234 GND.n5230 9.3005
R27003 GND.n5233 GND.n5232 9.3005
R27004 GND.n5231 GND.n444 9.3005
R27005 GND.n9724 GND.n445 9.3005
R27006 GND.n9723 GND.n446 9.3005
R27007 GND.n9722 GND.n447 9.3005
R27008 GND.n450 GND.n448 9.3005
R27009 GND.n9718 GND.n451 9.3005
R27010 GND.n9717 GND.n452 9.3005
R27011 GND.n9716 GND.n453 9.3005
R27012 GND.n456 GND.n454 9.3005
R27013 GND.n9712 GND.n457 9.3005
R27014 GND.n9711 GND.n458 9.3005
R27015 GND.n9710 GND.n459 9.3005
R27016 GND.n462 GND.n460 9.3005
R27017 GND.n9706 GND.n463 9.3005
R27018 GND.n9705 GND.n464 9.3005
R27019 GND.n9704 GND.n465 9.3005
R27020 GND.n468 GND.n466 9.3005
R27021 GND.n9700 GND.n469 9.3005
R27022 GND.n9699 GND.n470 9.3005
R27023 GND.n9698 GND.n471 9.3005
R27024 GND.n9686 GND.n472 9.3005
R27025 GND.n8242 GND.n8241 9.3005
R27026 GND.n8243 GND.n1432 9.3005
R27027 GND.n8246 GND.n1431 9.3005
R27028 GND.n8247 GND.n1430 9.3005
R27029 GND.n8250 GND.n1429 9.3005
R27030 GND.n8251 GND.n1428 9.3005
R27031 GND.n8254 GND.n1427 9.3005
R27032 GND.n8255 GND.n1426 9.3005
R27033 GND.n8258 GND.n1425 9.3005
R27034 GND.n8259 GND.n1424 9.3005
R27035 GND.n8262 GND.n1423 9.3005
R27036 GND.n8263 GND.n1422 9.3005
R27037 GND.n8266 GND.n1421 9.3005
R27038 GND.n8268 GND.n1418 9.3005
R27039 GND.n8271 GND.n1417 9.3005
R27040 GND.n8272 GND.n1416 9.3005
R27041 GND.n8275 GND.n1415 9.3005
R27042 GND.n8276 GND.n1414 9.3005
R27043 GND.n8279 GND.n1413 9.3005
R27044 GND.n8280 GND.n1412 9.3005
R27045 GND.n8283 GND.n1411 9.3005
R27046 GND.n8284 GND.n1410 9.3005
R27047 GND.n8287 GND.n1409 9.3005
R27048 GND.n8288 GND.n1408 9.3005
R27049 GND.n8291 GND.n1407 9.3005
R27050 GND.n8295 GND.n1403 9.3005
R27051 GND.n8296 GND.n1402 9.3005
R27052 GND.n8299 GND.n1401 9.3005
R27053 GND.n8300 GND.n1400 9.3005
R27054 GND.n8303 GND.n1399 9.3005
R27055 GND.n8304 GND.n1398 9.3005
R27056 GND.n8307 GND.n1397 9.3005
R27057 GND.n8308 GND.n1396 9.3005
R27058 GND.n8311 GND.n1395 9.3005
R27059 GND.n8312 GND.n1394 9.3005
R27060 GND.n8315 GND.n1393 9.3005
R27061 GND.n8316 GND.n1392 9.3005
R27062 GND.n8319 GND.n1388 9.3005
R27063 GND.n8320 GND.n1387 9.3005
R27064 GND.n8323 GND.n1386 9.3005
R27065 GND.n8324 GND.n1385 9.3005
R27066 GND.n8327 GND.n1384 9.3005
R27067 GND.n8328 GND.n1383 9.3005
R27068 GND.n8331 GND.n1382 9.3005
R27069 GND.n8332 GND.n1381 9.3005
R27070 GND.n8335 GND.n1380 9.3005
R27071 GND.n8336 GND.n1379 9.3005
R27072 GND.n8339 GND.n1378 9.3005
R27073 GND.n8341 GND.n1377 9.3005
R27074 GND.n8343 GND.n1372 9.3005
R27075 GND.n8346 GND.n1371 9.3005
R27076 GND.n8347 GND.n1370 9.3005
R27077 GND.n8350 GND.n1369 9.3005
R27078 GND.n8351 GND.n1368 9.3005
R27079 GND.n8354 GND.n1367 9.3005
R27080 GND.n8356 GND.n1366 9.3005
R27081 GND.n8357 GND.n1365 9.3005
R27082 GND.n8358 GND.n1364 9.3005
R27083 GND.n8359 GND.n1363 9.3005
R27084 GND.n8342 GND.n1374 9.3005
R27085 GND.n8292 GND.n1404 9.3005
R27086 GND.n8240 GND.n1433 9.3005
R27087 GND.n2940 GND.n2937 9.3005
R27088 GND.n2942 GND.n2941 9.3005
R27089 GND.n2909 GND.n2908 9.3005
R27090 GND.n2956 GND.n2955 9.3005
R27091 GND.n2957 GND.n2907 9.3005
R27092 GND.n2959 GND.n2958 9.3005
R27093 GND.n2889 GND.n2888 9.3005
R27094 GND.n2973 GND.n2972 9.3005
R27095 GND.n2974 GND.n2887 9.3005
R27096 GND.n2976 GND.n2975 9.3005
R27097 GND.n2870 GND.n2869 9.3005
R27098 GND.n2997 GND.n2996 9.3005
R27099 GND.n2998 GND.n2868 9.3005
R27100 GND.n3002 GND.n2999 9.3005
R27101 GND.n3001 GND.n3000 9.3005
R27102 GND.n2846 GND.n2845 9.3005
R27103 GND.n3030 GND.n3029 9.3005
R27104 GND.n3031 GND.n2844 9.3005
R27105 GND.n3033 GND.n3032 9.3005
R27106 GND.n2822 GND.n2821 9.3005
R27107 GND.n3063 GND.n3062 9.3005
R27108 GND.n3064 GND.n2820 9.3005
R27109 GND.n3068 GND.n3065 9.3005
R27110 GND.n3067 GND.n3066 9.3005
R27111 GND.n2793 GND.n2792 9.3005
R27112 GND.n3100 GND.n3099 9.3005
R27113 GND.n3101 GND.n2791 9.3005
R27114 GND.n3105 GND.n3102 9.3005
R27115 GND.n3104 GND.n3103 9.3005
R27116 GND.n2763 GND.n2762 9.3005
R27117 GND.n3138 GND.n3137 9.3005
R27118 GND.n3139 GND.n2761 9.3005
R27119 GND.n3143 GND.n3140 9.3005
R27120 GND.n3142 GND.n3141 9.3005
R27121 GND.n2736 GND.n2735 9.3005
R27122 GND.n3176 GND.n3175 9.3005
R27123 GND.n3177 GND.n2734 9.3005
R27124 GND.n3181 GND.n3178 9.3005
R27125 GND.n3180 GND.n3179 9.3005
R27126 GND.n2707 GND.n2706 9.3005
R27127 GND.n3213 GND.n3212 9.3005
R27128 GND.n3214 GND.n2705 9.3005
R27129 GND.n3218 GND.n3215 9.3005
R27130 GND.n3217 GND.n3216 9.3005
R27131 GND.n2678 GND.n2677 9.3005
R27132 GND.n3250 GND.n3249 9.3005
R27133 GND.n3251 GND.n2676 9.3005
R27134 GND.n3255 GND.n3252 9.3005
R27135 GND.n3254 GND.n3253 9.3005
R27136 GND.n2648 GND.n2647 9.3005
R27137 GND.n3287 GND.n3286 9.3005
R27138 GND.n3288 GND.n2646 9.3005
R27139 GND.n3293 GND.n3289 9.3005
R27140 GND.n3292 GND.n3290 9.3005
R27141 GND.n3291 GND.n1542 9.3005
R27142 GND.n1549 GND.n1541 9.3005
R27143 GND.n2581 GND.n2580 9.3005
R27144 GND.n3578 GND.n3577 9.3005
R27145 GND.n3579 GND.n2579 9.3005
R27146 GND.n3583 GND.n3580 9.3005
R27147 GND.n3582 GND.n3581 9.3005
R27148 GND.n2559 GND.n2558 9.3005
R27149 GND.n3604 GND.n3603 9.3005
R27150 GND.n3605 GND.n2557 9.3005
R27151 GND.n3609 GND.n3606 9.3005
R27152 GND.n3608 GND.n3607 9.3005
R27153 GND.n2538 GND.n2537 9.3005
R27154 GND.n3630 GND.n3629 9.3005
R27155 GND.n3631 GND.n2536 9.3005
R27156 GND.n3635 GND.n3632 9.3005
R27157 GND.n3634 GND.n3633 9.3005
R27158 GND.n2516 GND.n2515 9.3005
R27159 GND.n3656 GND.n3655 9.3005
R27160 GND.n3657 GND.n2514 9.3005
R27161 GND.n3661 GND.n3658 9.3005
R27162 GND.n3660 GND.n3659 9.3005
R27163 GND.n2494 GND.n2493 9.3005
R27164 GND.n3681 GND.n3680 9.3005
R27165 GND.n3682 GND.n2492 9.3005
R27166 GND.n3686 GND.n3683 9.3005
R27167 GND.n3685 GND.n3684 9.3005
R27168 GND.n2472 GND.n2471 9.3005
R27169 GND.n3707 GND.n3706 9.3005
R27170 GND.n3708 GND.n2470 9.3005
R27171 GND.n3712 GND.n3709 9.3005
R27172 GND.n3711 GND.n3710 9.3005
R27173 GND.n2451 GND.n2450 9.3005
R27174 GND.n3733 GND.n3732 9.3005
R27175 GND.n3734 GND.n2449 9.3005
R27176 GND.n3738 GND.n3735 9.3005
R27177 GND.n3737 GND.n3736 9.3005
R27178 GND.n2431 GND.n2430 9.3005
R27179 GND.n3759 GND.n3758 9.3005
R27180 GND.n3760 GND.n2429 9.3005
R27181 GND.n3764 GND.n3761 9.3005
R27182 GND.n3763 GND.n3762 9.3005
R27183 GND.n2409 GND.n2408 9.3005
R27184 GND.n3784 GND.n3783 9.3005
R27185 GND.n3785 GND.n2407 9.3005
R27186 GND.n3789 GND.n3786 9.3005
R27187 GND.n3788 GND.n3787 9.3005
R27188 GND.n2387 GND.n2386 9.3005
R27189 GND.n3810 GND.n3809 9.3005
R27190 GND.n3811 GND.n2385 9.3005
R27191 GND.n3815 GND.n3812 9.3005
R27192 GND.n3814 GND.n3813 9.3005
R27193 GND.n2366 GND.n2365 9.3005
R27194 GND.n3837 GND.n3836 9.3005
R27195 GND.n3838 GND.n2364 9.3005
R27196 GND.n3841 GND.n3839 9.3005
R27197 GND.n3840 GND.n1724 9.3005
R27198 GND.n2939 GND.n2938 9.3005
R27199 GND.n8119 GND.n1546 9.3005
R27200 GND.n8119 GND.n8118 9.3005
R27201 GND.n3011 GND.n3008 9.3005
R27202 GND.n3015 GND.n3012 9.3005
R27203 GND.n3014 GND.n3013 9.3005
R27204 GND.n2838 GND.n2837 9.3005
R27205 GND.n3039 GND.n3038 9.3005
R27206 GND.n3040 GND.n2836 9.3005
R27207 GND.n3042 GND.n3041 9.3005
R27208 GND.n2811 GND.n2810 9.3005
R27209 GND.n3074 GND.n3073 9.3005
R27210 GND.n3075 GND.n2809 9.3005
R27211 GND.n3079 GND.n3076 9.3005
R27212 GND.n3078 GND.n3077 9.3005
R27213 GND.n2782 GND.n2781 9.3005
R27214 GND.n3111 GND.n3110 9.3005
R27215 GND.n3112 GND.n2780 9.3005
R27216 GND.n3116 GND.n3113 9.3005
R27217 GND.n3115 GND.n3114 9.3005
R27218 GND.n2754 GND.n2753 9.3005
R27219 GND.n3149 GND.n3148 9.3005
R27220 GND.n3150 GND.n2752 9.3005
R27221 GND.n3154 GND.n3151 9.3005
R27222 GND.n3153 GND.n3152 9.3005
R27223 GND.n2726 GND.n2725 9.3005
R27224 GND.n3187 GND.n3186 9.3005
R27225 GND.n3188 GND.n2724 9.3005
R27226 GND.n3192 GND.n3189 9.3005
R27227 GND.n3191 GND.n3190 9.3005
R27228 GND.n2696 GND.n2695 9.3005
R27229 GND.n3224 GND.n3223 9.3005
R27230 GND.n3225 GND.n2694 9.3005
R27231 GND.n3229 GND.n3226 9.3005
R27232 GND.n3228 GND.n3227 9.3005
R27233 GND.n2667 GND.n2666 9.3005
R27234 GND.n3261 GND.n3260 9.3005
R27235 GND.n3262 GND.n2665 9.3005
R27236 GND.n3266 GND.n3263 9.3005
R27237 GND.n3265 GND.n3264 9.3005
R27238 GND.n2638 GND.n2637 9.3005
R27239 GND.n3299 GND.n3298 9.3005
R27240 GND.n3300 GND.n2636 9.3005
R27241 GND.n3304 GND.n3301 9.3005
R27242 GND.n3010 GND.n3009 9.3005
R27243 GND.n8366 GND.n1319 9.3005
R27244 GND.n8367 GND.n1318 9.3005
R27245 GND.n1317 GND.n1313 9.3005
R27246 GND.n8373 GND.n1312 9.3005
R27247 GND.n8374 GND.n1311 9.3005
R27248 GND.n8375 GND.n1310 9.3005
R27249 GND.n1309 GND.n1305 9.3005
R27250 GND.n8381 GND.n1304 9.3005
R27251 GND.n8382 GND.n1303 9.3005
R27252 GND.n8383 GND.n1302 9.3005
R27253 GND.n1301 GND.n1297 9.3005
R27254 GND.n8389 GND.n1296 9.3005
R27255 GND.n8390 GND.n1295 9.3005
R27256 GND.n8391 GND.n1294 9.3005
R27257 GND.n1293 GND.n1289 9.3005
R27258 GND.n8397 GND.n1288 9.3005
R27259 GND.n8398 GND.n1287 9.3005
R27260 GND.n8399 GND.n1286 9.3005
R27261 GND.n1285 GND.n1281 9.3005
R27262 GND.n8405 GND.n1280 9.3005
R27263 GND.n8406 GND.n1279 9.3005
R27264 GND.n8407 GND.n1278 9.3005
R27265 GND.n1277 GND.n1273 9.3005
R27266 GND.n8413 GND.n1272 9.3005
R27267 GND.n8414 GND.n1271 9.3005
R27268 GND.n8415 GND.n1270 9.3005
R27269 GND.n1269 GND.n1265 9.3005
R27270 GND.n8421 GND.n1264 9.3005
R27271 GND.n8422 GND.n1263 9.3005
R27272 GND.n8423 GND.n1262 9.3005
R27273 GND.n1261 GND.n1257 9.3005
R27274 GND.n8429 GND.n1256 9.3005
R27275 GND.n8430 GND.n1255 9.3005
R27276 GND.n8431 GND.n1254 9.3005
R27277 GND.n1253 GND.n1249 9.3005
R27278 GND.n8437 GND.n1248 9.3005
R27279 GND.n8438 GND.n1247 9.3005
R27280 GND.n8439 GND.n1246 9.3005
R27281 GND.n1245 GND.n1241 9.3005
R27282 GND.n8445 GND.n1240 9.3005
R27283 GND.n8446 GND.n1239 9.3005
R27284 GND.n8447 GND.n1238 9.3005
R27285 GND.n1237 GND.n1233 9.3005
R27286 GND.n8453 GND.n1232 9.3005
R27287 GND.n8454 GND.n1231 9.3005
R27288 GND.n8455 GND.n1230 9.3005
R27289 GND.n1229 GND.n1225 9.3005
R27290 GND.n8461 GND.n1224 9.3005
R27291 GND.n8462 GND.n1223 9.3005
R27292 GND.n8463 GND.n1222 9.3005
R27293 GND.n1221 GND.n1217 9.3005
R27294 GND.n8469 GND.n1216 9.3005
R27295 GND.n8470 GND.n1215 9.3005
R27296 GND.n8471 GND.n1214 9.3005
R27297 GND.n1213 GND.n1209 9.3005
R27298 GND.n8477 GND.n1208 9.3005
R27299 GND.n8478 GND.n1207 9.3005
R27300 GND.n8479 GND.n1206 9.3005
R27301 GND.n1205 GND.n1201 9.3005
R27302 GND.n8485 GND.n1200 9.3005
R27303 GND.n8486 GND.n1199 9.3005
R27304 GND.n8487 GND.n1198 9.3005
R27305 GND.n1197 GND.n1193 9.3005
R27306 GND.n8493 GND.n1192 9.3005
R27307 GND.n8494 GND.n1191 9.3005
R27308 GND.n8495 GND.n1190 9.3005
R27309 GND.n8365 GND.n1320 9.3005
R27310 GND.n7739 GND.n7738 9.3005
R27311 GND.n7979 GND.n1765 9.3005
R27312 GND.n7981 GND.n7980 9.3005
R27313 GND.n7982 GND.n1764 9.3005
R27314 GND.n7984 GND.n7983 9.3005
R27315 GND.n7985 GND.n1757 9.3005
R27316 GND.n7988 GND.n7987 9.3005
R27317 GND.n7989 GND.n1756 9.3005
R27318 GND.n7991 GND.n7990 9.3005
R27319 GND.n7992 GND.n1751 9.3005
R27320 GND.n7994 GND.n7993 9.3005
R27321 GND.n7995 GND.n1750 9.3005
R27322 GND.n7997 GND.n7996 9.3005
R27323 GND.n7998 GND.n1745 9.3005
R27324 GND.n8000 GND.n7999 9.3005
R27325 GND.n8001 GND.n1744 9.3005
R27326 GND.n8003 GND.n8002 9.3005
R27327 GND.n8004 GND.n1737 9.3005
R27328 GND.n8006 GND.n8005 9.3005
R27329 GND.n8007 GND.n1736 9.3005
R27330 GND.n8009 GND.n8008 9.3005
R27331 GND.n8010 GND.n1731 9.3005
R27332 GND.n8012 GND.n8011 9.3005
R27333 GND.n8013 GND.n1730 9.3005
R27334 GND.n8015 GND.n8014 9.3005
R27335 GND.n8016 GND.n1725 9.3005
R27336 GND.n8018 GND.n8017 9.3005
R27337 GND.n8019 GND.n1723 9.3005
R27338 GND.n8021 GND.n8020 9.3005
R27339 GND.n1868 GND.n1768 9.3005
R27340 GND.n1867 GND.n1866 9.3005
R27341 GND.n1865 GND.n1769 9.3005
R27342 GND.n1864 GND.n1863 9.3005
R27343 GND.n1862 GND.n1774 9.3005
R27344 GND.n1861 GND.n1860 9.3005
R27345 GND.n1859 GND.n1775 9.3005
R27346 GND.n1858 GND.n1857 9.3005
R27347 GND.n1856 GND.n1782 9.3005
R27348 GND.n1855 GND.n1854 9.3005
R27349 GND.n1853 GND.n1783 9.3005
R27350 GND.n1852 GND.n1851 9.3005
R27351 GND.n1850 GND.n1788 9.3005
R27352 GND.n1849 GND.n1848 9.3005
R27353 GND.n1847 GND.n1789 9.3005
R27354 GND.n1846 GND.n1845 9.3005
R27355 GND.n1844 GND.n1794 9.3005
R27356 GND.n1843 GND.n1842 9.3005
R27357 GND.n1840 GND.n1795 9.3005
R27358 GND.n1839 GND.n1838 9.3005
R27359 GND.n1837 GND.n1802 9.3005
R27360 GND.n1836 GND.n1835 9.3005
R27361 GND.n1834 GND.n1803 9.3005
R27362 GND.n1833 GND.n1832 9.3005
R27363 GND.n1831 GND.n1808 9.3005
R27364 GND.n1830 GND.n1829 9.3005
R27365 GND.n1828 GND.n1809 9.3005
R27366 GND.n1827 GND.n1826 9.3005
R27367 GND.n1825 GND.n1814 9.3005
R27368 GND.n1824 GND.n1823 9.3005
R27369 GND.n1822 GND.n1815 9.3005
R27370 GND.n1821 GND.n1820 9.3005
R27371 GND.n2932 GND.n2928 9.3005
R27372 GND.n2934 GND.n2933 9.3005
R27373 GND.n2918 GND.n2916 9.3005
R27374 GND.n2951 GND.n2950 9.3005
R27375 GND.n2921 GND.n2917 9.3005
R27376 GND.n2920 GND.n2919 9.3005
R27377 GND.n2898 GND.n2896 9.3005
R27378 GND.n2968 GND.n2967 9.3005
R27379 GND.n2901 GND.n2897 9.3005
R27380 GND.n2900 GND.n2899 9.3005
R27381 GND.n2880 GND.n2878 9.3005
R27382 GND.n2992 GND.n2991 9.3005
R27383 GND.n2881 GND.n2879 9.3005
R27384 GND.n2987 GND.n2983 9.3005
R27385 GND.n2986 GND.n2985 9.3005
R27386 GND.n2855 GND.n2853 9.3005
R27387 GND.n3025 GND.n3024 9.3005
R27388 GND.n2858 GND.n2854 9.3005
R27389 GND.n2857 GND.n2856 9.3005
R27390 GND.n2830 GND.n2828 9.3005
R27391 GND.n3058 GND.n3057 9.3005
R27392 GND.n2831 GND.n2829 9.3005
R27393 GND.n3053 GND.n3049 9.3005
R27394 GND.n3052 GND.n3051 9.3005
R27395 GND.n2802 GND.n2800 9.3005
R27396 GND.n3095 GND.n3094 9.3005
R27397 GND.n2803 GND.n2801 9.3005
R27398 GND.n3090 GND.n3086 9.3005
R27399 GND.n3089 GND.n3088 9.3005
R27400 GND.n2773 GND.n2771 9.3005
R27401 GND.n3133 GND.n3132 9.3005
R27402 GND.n2774 GND.n2772 9.3005
R27403 GND.n3128 GND.n3124 9.3005
R27404 GND.n3127 GND.n3126 9.3005
R27405 GND.n2745 GND.n2743 9.3005
R27406 GND.n3171 GND.n3170 9.3005
R27407 GND.n2746 GND.n2744 9.3005
R27408 GND.n3166 GND.n3162 9.3005
R27409 GND.n3165 GND.n3164 9.3005
R27410 GND.n2716 GND.n2714 9.3005
R27411 GND.n3208 GND.n3207 9.3005
R27412 GND.n2717 GND.n2715 9.3005
R27413 GND.n3203 GND.n3199 9.3005
R27414 GND.n3202 GND.n3201 9.3005
R27415 GND.n2687 GND.n2685 9.3005
R27416 GND.n3245 GND.n3244 9.3005
R27417 GND.n2688 GND.n2686 9.3005
R27418 GND.n3240 GND.n3236 9.3005
R27419 GND.n3239 GND.n3238 9.3005
R27420 GND.n2658 GND.n2656 9.3005
R27421 GND.n3282 GND.n3281 9.3005
R27422 GND.n2659 GND.n2657 9.3005
R27423 GND.n3277 GND.n3273 9.3005
R27424 GND.n3276 GND.n3275 9.3005
R27425 GND.n2629 GND.n2627 9.3005
R27426 GND.n3318 GND.n3317 9.3005
R27427 GND.n2630 GND.n2628 9.3005
R27428 GND.n3313 GND.n3312 9.3005
R27429 GND.n2607 GND.n2606 9.3005
R27430 GND.n3546 GND.n3545 9.3005
R27431 GND.n3544 GND.n2603 9.3005
R27432 GND.n3550 GND.n2602 9.3005
R27433 GND.n3552 GND.n3551 9.3005
R27434 GND.n1560 GND.n1558 9.3005
R27435 GND.n8114 GND.n8113 9.3005
R27436 GND.n1561 GND.n1559 9.3005
R27437 GND.n8109 GND.n1566 9.3005
R27438 GND.n8108 GND.n1567 9.3005
R27439 GND.n8107 GND.n1568 9.3005
R27440 GND.n2574 GND.n1569 9.3005
R27441 GND.n8103 GND.n1574 9.3005
R27442 GND.n8102 GND.n1575 9.3005
R27443 GND.n8101 GND.n1576 9.3005
R27444 GND.n3597 GND.n1577 9.3005
R27445 GND.n8097 GND.n1582 9.3005
R27446 GND.n8096 GND.n1583 9.3005
R27447 GND.n8095 GND.n1584 9.3005
R27448 GND.n3625 GND.n1585 9.3005
R27449 GND.n8091 GND.n1590 9.3005
R27450 GND.n8090 GND.n1591 9.3005
R27451 GND.n8089 GND.n1592 9.3005
R27452 GND.n2522 GND.n1593 9.3005
R27453 GND.n8085 GND.n1598 9.3005
R27454 GND.n8084 GND.n1599 9.3005
R27455 GND.n8083 GND.n1600 9.3005
R27456 GND.n2500 GND.n1601 9.3005
R27457 GND.n8079 GND.n1606 9.3005
R27458 GND.n8078 GND.n1607 9.3005
R27459 GND.n8077 GND.n1608 9.3005
R27460 GND.n2487 GND.n1609 9.3005
R27461 GND.n8073 GND.n1614 9.3005
R27462 GND.n8072 GND.n1615 9.3005
R27463 GND.n8071 GND.n1616 9.3005
R27464 GND.n3700 GND.n1617 9.3005
R27465 GND.n8067 GND.n1622 9.3005
R27466 GND.n8066 GND.n1623 9.3005
R27467 GND.n8065 GND.n1624 9.3005
R27468 GND.n3728 GND.n1625 9.3005
R27469 GND.n8061 GND.n1630 9.3005
R27470 GND.n8060 GND.n1631 9.3005
R27471 GND.n8059 GND.n1632 9.3005
R27472 GND.n2437 GND.n1633 9.3005
R27473 GND.n8055 GND.n1638 9.3005
R27474 GND.n8054 GND.n1639 9.3005
R27475 GND.n8053 GND.n1640 9.3005
R27476 GND.n2415 GND.n1641 9.3005
R27477 GND.n8049 GND.n1646 9.3005
R27478 GND.n8048 GND.n1647 9.3005
R27479 GND.n8047 GND.n1648 9.3005
R27480 GND.n2402 GND.n1649 9.3005
R27481 GND.n8043 GND.n1654 9.3005
R27482 GND.n8042 GND.n1655 9.3005
R27483 GND.n8041 GND.n1656 9.3005
R27484 GND.n3803 GND.n1657 9.3005
R27485 GND.n8037 GND.n1662 9.3005
R27486 GND.n8036 GND.n1663 9.3005
R27487 GND.n8035 GND.n1664 9.3005
R27488 GND.n3832 GND.n1665 9.3005
R27489 GND.n8031 GND.n1670 9.3005
R27490 GND.n8030 GND.n1671 9.3005
R27491 GND.n8029 GND.n1672 9.3005
R27492 GND.n2927 GND.n1437 9.3005
R27493 GND.n2932 GND.n2931 9.3005
R27494 GND.n2933 GND.n2922 9.3005
R27495 GND.n2947 GND.n2918 9.3005
R27496 GND.n2950 GND.n2949 9.3005
R27497 GND.n2948 GND.n2921 9.3005
R27498 GND.n2920 GND.n2902 9.3005
R27499 GND.n2964 GND.n2898 9.3005
R27500 GND.n2967 GND.n2966 9.3005
R27501 GND.n2965 GND.n2901 9.3005
R27502 GND.n2900 GND.n2882 9.3005
R27503 GND.n2981 GND.n2880 9.3005
R27504 GND.n2991 GND.n2990 9.3005
R27505 GND.n2989 GND.n2881 9.3005
R27506 GND.n2988 GND.n2987 9.3005
R27507 GND.n2986 GND.n2859 9.3005
R27508 GND.n3020 GND.n2855 9.3005
R27509 GND.n3024 GND.n3023 9.3005
R27510 GND.n3022 GND.n2858 9.3005
R27511 GND.n2857 GND.n2832 9.3005
R27512 GND.n3047 GND.n2830 9.3005
R27513 GND.n3057 GND.n3056 9.3005
R27514 GND.n3055 GND.n2831 9.3005
R27515 GND.n3054 GND.n3053 9.3005
R27516 GND.n3052 GND.n2804 9.3005
R27517 GND.n3084 GND.n2802 9.3005
R27518 GND.n3094 GND.n3093 9.3005
R27519 GND.n3092 GND.n2803 9.3005
R27520 GND.n3091 GND.n3090 9.3005
R27521 GND.n3089 GND.n2775 9.3005
R27522 GND.n3121 GND.n2773 9.3005
R27523 GND.n3132 GND.n3131 9.3005
R27524 GND.n3130 GND.n2774 9.3005
R27525 GND.n3129 GND.n3128 9.3005
R27526 GND.n3127 GND.n2747 9.3005
R27527 GND.n3160 GND.n2745 9.3005
R27528 GND.n3170 GND.n3169 9.3005
R27529 GND.n3168 GND.n2746 9.3005
R27530 GND.n3167 GND.n3166 9.3005
R27531 GND.n3165 GND.n2718 9.3005
R27532 GND.n3197 GND.n2716 9.3005
R27533 GND.n3207 GND.n3206 9.3005
R27534 GND.n3205 GND.n2717 9.3005
R27535 GND.n3204 GND.n3203 9.3005
R27536 GND.n3202 GND.n2689 9.3005
R27537 GND.n3234 GND.n2687 9.3005
R27538 GND.n3244 GND.n3243 9.3005
R27539 GND.n3242 GND.n2688 9.3005
R27540 GND.n3241 GND.n3240 9.3005
R27541 GND.n3239 GND.n2660 9.3005
R27542 GND.n3271 GND.n2658 9.3005
R27543 GND.n3281 GND.n3280 9.3005
R27544 GND.n3279 GND.n2659 9.3005
R27545 GND.n3278 GND.n3277 9.3005
R27546 GND.n3276 GND.n2631 9.3005
R27547 GND.n3310 GND.n2629 9.3005
R27548 GND.n3317 GND.n3316 9.3005
R27549 GND.n3315 GND.n2630 9.3005
R27550 GND.n3314 GND.n3313 9.3005
R27551 GND.n2606 GND.n2604 9.3005
R27552 GND.n3547 GND.n3546 9.3005
R27553 GND.n3548 GND.n2603 9.3005
R27554 GND.n3550 GND.n3549 9.3005
R27555 GND.n3551 GND.n2598 9.3005
R27556 GND.n1562 GND.n1560 9.3005
R27557 GND.n8113 GND.n8112 9.3005
R27558 GND.n8111 GND.n1561 9.3005
R27559 GND.n8110 GND.n8109 9.3005
R27560 GND.n8108 GND.n1565 9.3005
R27561 GND.n8107 GND.n8106 9.3005
R27562 GND.n8105 GND.n1569 9.3005
R27563 GND.n8104 GND.n8103 9.3005
R27564 GND.n8102 GND.n1573 9.3005
R27565 GND.n8101 GND.n8100 9.3005
R27566 GND.n8099 GND.n1577 9.3005
R27567 GND.n8098 GND.n8097 9.3005
R27568 GND.n8096 GND.n1581 9.3005
R27569 GND.n8095 GND.n8094 9.3005
R27570 GND.n8093 GND.n1585 9.3005
R27571 GND.n8092 GND.n8091 9.3005
R27572 GND.n8090 GND.n1589 9.3005
R27573 GND.n8089 GND.n8088 9.3005
R27574 GND.n8087 GND.n1593 9.3005
R27575 GND.n8086 GND.n8085 9.3005
R27576 GND.n8084 GND.n1597 9.3005
R27577 GND.n8083 GND.n8082 9.3005
R27578 GND.n8081 GND.n1601 9.3005
R27579 GND.n8080 GND.n8079 9.3005
R27580 GND.n8078 GND.n1605 9.3005
R27581 GND.n8077 GND.n8076 9.3005
R27582 GND.n8075 GND.n1609 9.3005
R27583 GND.n8074 GND.n8073 9.3005
R27584 GND.n8072 GND.n1613 9.3005
R27585 GND.n8071 GND.n8070 9.3005
R27586 GND.n8069 GND.n1617 9.3005
R27587 GND.n8068 GND.n8067 9.3005
R27588 GND.n8066 GND.n1621 9.3005
R27589 GND.n8065 GND.n8064 9.3005
R27590 GND.n8063 GND.n1625 9.3005
R27591 GND.n8062 GND.n8061 9.3005
R27592 GND.n8060 GND.n1629 9.3005
R27593 GND.n8059 GND.n8058 9.3005
R27594 GND.n8057 GND.n1633 9.3005
R27595 GND.n8056 GND.n8055 9.3005
R27596 GND.n8054 GND.n1637 9.3005
R27597 GND.n8053 GND.n8052 9.3005
R27598 GND.n8051 GND.n1641 9.3005
R27599 GND.n8050 GND.n8049 9.3005
R27600 GND.n8048 GND.n1645 9.3005
R27601 GND.n8047 GND.n8046 9.3005
R27602 GND.n8045 GND.n1649 9.3005
R27603 GND.n8044 GND.n8043 9.3005
R27604 GND.n8042 GND.n1653 9.3005
R27605 GND.n8041 GND.n8040 9.3005
R27606 GND.n8039 GND.n1657 9.3005
R27607 GND.n8038 GND.n8037 9.3005
R27608 GND.n8036 GND.n1661 9.3005
R27609 GND.n8035 GND.n8034 9.3005
R27610 GND.n8033 GND.n1665 9.3005
R27611 GND.n8032 GND.n8031 9.3005
R27612 GND.n8030 GND.n1669 9.3005
R27613 GND.n8029 GND.n8028 9.3005
R27614 GND.n2930 GND.n1437 9.3005
R27615 GND.n8224 GND.n1449 9.3005
R27616 GND.n8226 GND.n8225 9.3005
R27617 GND.n8227 GND.n1448 9.3005
R27618 GND.n8229 GND.n8228 9.3005
R27619 GND.n8230 GND.n1443 9.3005
R27620 GND.n8232 GND.n8231 9.3005
R27621 GND.n8233 GND.n1442 9.3005
R27622 GND.n8235 GND.n8234 9.3005
R27623 GND.n8236 GND.n1438 9.3005
R27624 GND.n8238 GND.n8237 9.3005
R27625 GND.n8223 GND.n8219 9.3005
R27626 GND.n8218 GND.n1452 9.3005
R27627 GND.n8215 GND.n1453 9.3005
R27628 GND.n8214 GND.n8213 9.3005
R27629 GND.n8212 GND.n1457 9.3005
R27630 GND.n8211 GND.n8210 9.3005
R27631 GND.n8209 GND.n1458 9.3005
R27632 GND.n8208 GND.n8207 9.3005
R27633 GND.n8206 GND.n1462 9.3005
R27634 GND.n8205 GND.n8204 9.3005
R27635 GND.n8203 GND.n1463 9.3005
R27636 GND.n8202 GND.n8201 9.3005
R27637 GND.n8200 GND.n1467 9.3005
R27638 GND.n8199 GND.n8198 9.3005
R27639 GND.n8197 GND.n1468 9.3005
R27640 GND.n8196 GND.n8195 9.3005
R27641 GND.n8194 GND.n1472 9.3005
R27642 GND.n8193 GND.n8192 9.3005
R27643 GND.n8191 GND.n1473 9.3005
R27644 GND.n8190 GND.n8189 9.3005
R27645 GND.n8188 GND.n1477 9.3005
R27646 GND.n8187 GND.n8186 9.3005
R27647 GND.n8185 GND.n1478 9.3005
R27648 GND.n8184 GND.n8183 9.3005
R27649 GND.n8182 GND.n1482 9.3005
R27650 GND.n8181 GND.n8180 9.3005
R27651 GND.n8179 GND.n1483 9.3005
R27652 GND.n8178 GND.n8177 9.3005
R27653 GND.n8176 GND.n1487 9.3005
R27654 GND.n8175 GND.n8174 9.3005
R27655 GND.n8173 GND.n1488 9.3005
R27656 GND.n8172 GND.n8171 9.3005
R27657 GND.n8170 GND.n1492 9.3005
R27658 GND.n8169 GND.n8168 9.3005
R27659 GND.n8167 GND.n1493 9.3005
R27660 GND.n8166 GND.n8165 9.3005
R27661 GND.n8164 GND.n1497 9.3005
R27662 GND.n8163 GND.n8162 9.3005
R27663 GND.n8161 GND.n1498 9.3005
R27664 GND.n8160 GND.n8159 9.3005
R27665 GND.n8158 GND.n1502 9.3005
R27666 GND.n8157 GND.n8156 9.3005
R27667 GND.n8155 GND.n1503 9.3005
R27668 GND.n8154 GND.n8153 9.3005
R27669 GND.n8152 GND.n1507 9.3005
R27670 GND.n8151 GND.n8150 9.3005
R27671 GND.n8149 GND.n1508 9.3005
R27672 GND.n8148 GND.n8147 9.3005
R27673 GND.n8146 GND.n1512 9.3005
R27674 GND.n8145 GND.n8144 9.3005
R27675 GND.n8143 GND.n1513 9.3005
R27676 GND.n8142 GND.n8141 9.3005
R27677 GND.n8140 GND.n1517 9.3005
R27678 GND.n8139 GND.n8138 9.3005
R27679 GND.n8137 GND.n1518 9.3005
R27680 GND.n8136 GND.n8135 9.3005
R27681 GND.n8134 GND.n1522 9.3005
R27682 GND.n8133 GND.n8132 9.3005
R27683 GND.n8131 GND.n1523 9.3005
R27684 GND.n8130 GND.n8129 9.3005
R27685 GND.n8128 GND.n1527 9.3005
R27686 GND.n8127 GND.n8126 9.3005
R27687 GND.n8217 GND.n8216 9.3005
R27688 GND.n2190 GND.n2187 9.13319
R27689 GND.n1971 GND.n1965 9.13319
R27690 GND.n7849 GND.n7848 9.13319
R27691 GND.n7828 GND.n7827 9.13319
R27692 GND.n2097 GND.n2091 9.13319
R27693 GND.n7767 GND.n7766 9.13319
R27694 GND.n5759 GND.n5758 9.13319
R27695 GND.n5863 GND.n5862 9.13319
R27696 GND.n7601 GND.n7600 9.13319
R27697 GND.n5966 GND.n5965 9.13319
R27698 GND.n7546 GND.n7545 9.13319
R27699 GND.n6069 GND.n6068 9.13319
R27700 GND.n7491 GND.n7490 9.13319
R27701 GND.n7436 GND.n7435 9.13319
R27702 GND.n7401 GND.n7400 9.13319
R27703 GND.n7380 GND.n7379 9.13319
R27704 GND.n4527 GND.n4521 9.13319
R27705 GND.n7319 GND.n7318 9.13319
R27706 GND.n4666 GND.n4607 9.13319
R27707 GND.n4680 GND.t149 9.13319
R27708 GND.n7979 GND.n7977 8.72777
R27709 GND.n7187 GND.n4833 8.72777
R27710 GND.n5901 GND.t13 8.48086
R27711 GND.n7515 GND.t18 8.48086
R27712 GND.t61 GND.n4675 8.48086
R27713 GND.n10315 GND.n10314 8.23019
R27714 GND.n1528 GND.n47 8.23019
R27715 GND.n7884 GND.t97 8.15469
R27716 GND.t26 GND.n7283 8.15469
R27717 GND.n1938 GND.n1936 7.82852
R27718 GND.n2214 GND.n2211 7.82852
R27719 GND.n7855 GND.n2009 7.82852
R27720 GND.n7821 GND.n2053 7.82852
R27721 GND.n2291 GND.n2288 7.82852
R27722 GND.n7760 GND.n2327 7.82852
R27723 GND.n5745 GND.n5659 7.82852
R27724 GND.n7649 GND.n3964 7.82852
R27725 GND.n5849 GND.n5628 7.82852
R27726 GND.n7594 GND.n4069 7.82852
R27727 GND.n5952 GND.n5597 7.82852
R27728 GND.n7539 GND.n4174 7.82852
R27729 GND.n6055 GND.n5565 7.82852
R27730 GND.n7484 GND.n4277 7.82852
R27731 GND.n6158 GND.n5532 7.82852
R27732 GND.n7429 GND.n4381 7.82852
R27733 GND.n7407 GND.n4436 7.82852
R27734 GND.n7373 GND.n4483 7.82852
R27735 GND.n6253 GND.n6250 7.82852
R27736 GND.n7312 GND.n4569 7.82852
R27737 GND.n4661 GND.n4658 7.82852
R27738 GND.n7251 GND.n4700 7.82852
R27739 GND.n7904 GND.t88 7.17619
R27740 GND.n7793 GND.t3 6.85002
R27741 GND.n7656 GND.t20 6.85002
R27742 GND.t7 GND.n6171 6.85002
R27743 GND.n6276 GND.t5 6.85002
R27744 GND.n4828 GND.n4762 6.5566
R27745 GND.n2127 GND.n2123 6.5566
R27746 GND.n7920 GND.n7919 6.5566
R27747 GND.n7197 GND.n7196 6.5566
R27748 GND.t91 GND.n1971 6.52385
R27749 GND.n7884 GND.t91 6.52385
R27750 GND.n1989 GND.n1983 6.52385
R27751 GND.n7863 GND.n7862 6.52385
R27752 GND.n7814 GND.n7813 6.52385
R27753 GND.n2079 GND.n2073 6.52385
R27754 GND.n7697 GND.n3885 6.52385
R27755 GND.n5730 GND.n5664 6.52385
R27756 GND.n7643 GND.n3987 6.52385
R27757 GND.n5834 GND.n5633 6.52385
R27758 GND.n7588 GND.n4092 6.52385
R27759 GND.n5937 GND.n5602 6.52385
R27760 GND.n7533 GND.n4197 6.52385
R27761 GND.n6040 GND.n5570 6.52385
R27762 GND.n7478 GND.n4299 6.52385
R27763 GND.n6143 GND.n5537 6.52385
R27764 GND.n7423 GND.n4404 6.52385
R27765 GND.n6312 GND.n6311 6.52385
R27766 GND.n7366 GND.n7365 6.52385
R27767 GND.n4509 GND.n4503 6.52385
R27768 GND.n7305 GND.n7304 6.52385
R27769 GND.n4595 GND.n4589 6.52385
R27770 GND.n7258 GND.t125 6.52385
R27771 GND.t190 GND.n2701 6.19768
R27772 GND.t159 GND.n3306 6.19768
R27773 GND.n3308 GND.t159 6.19768
R27774 GND.n2588 GND.t169 6.19768
R27775 GND.n6926 GND.t163 6.19768
R27776 GND.n6895 GND.t175 6.19768
R27777 GND.t175 GND.n139 6.19768
R27778 GND.t173 GND.n194 6.19768
R27779 GND.n2202 GND.t52 5.87152
R27780 GND.t70 GND.n4700 5.87152
R27781 GND.n7987 GND.n7986 5.62474
R27782 GND.n7140 GND.n7124 5.62474
R27783 GND.n9940 GND.n9939 5.62474
R27784 GND.n8319 GND.n1391 5.62474
R27785 GND.n7189 GND.n4832 5.62001
R27786 GND.n7976 GND.n1871 5.62001
R27787 GND.n7976 GND.n7975 5.62001
R27788 GND.n7192 GND.n7189 5.62001
R27789 GND.t267 GND.n4027 5.54535
R27790 GND.t9 GND.n4262 5.54535
R27791 GND.n21 GND.n13 5.53211
R27792 GND.n69 GND.n61 5.53211
R27793 GND.n47 GND.n46 5.44637
R27794 GND.n10315 GND.n101 5.44637
R27795 GND.n7869 GND.n1991 5.21918
R27796 GND.n2227 GND.n2224 5.21918
R27797 GND.n2278 GND.n2275 5.21918
R27798 GND.n7807 GND.n2071 5.21918
R27799 GND.n7691 GND.n3894 5.21918
R27800 GND.n5825 GND.n5638 5.21918
R27801 GND.n7637 GND.n3997 5.21918
R27802 GND.n5928 GND.n5607 5.21918
R27803 GND.n7582 GND.n4102 5.21918
R27804 GND.n6031 GND.n5575 5.21918
R27805 GND.n7527 GND.n4206 5.21918
R27806 GND.n6134 GND.n5542 5.21918
R27807 GND.n7472 GND.n4309 5.21918
R27808 GND.n6194 GND.n5509 5.21918
R27809 GND.n6266 GND.n6263 5.21918
R27810 GND.n7359 GND.n4501 5.21918
R27811 GND.n4648 GND.n4645 5.21918
R27812 GND.n7298 GND.n4587 5.21918
R27813 GND.n7249 GND.t104 4.89301
R27814 GND.n7737 GND.n7736 4.74817
R27815 GND.n7732 GND.n7731 4.74817
R27816 GND.n7727 GND.n7726 4.74817
R27817 GND.n7722 GND.n7721 4.74817
R27818 GND.n7717 GND.n7716 4.74817
R27819 GND.n7712 GND.n7711 4.74817
R27820 GND.n6340 GND.n6339 4.74817
R27821 GND.n5486 GND.n5485 4.74817
R27822 GND.n5481 GND.n5480 4.74817
R27823 GND.n5476 GND.n5475 4.74817
R27824 GND.n5471 GND.n5470 4.74817
R27825 GND.n6341 GND.n5466 4.74817
R27826 GND.n6367 GND.n6366 4.74817
R27827 GND.n6372 GND.n6371 4.74817
R27828 GND.n6377 GND.n6376 4.74817
R27829 GND.n6384 GND.n6382 4.74817
R27830 GND.n6382 GND.n6381 4.74817
R27831 GND.n6378 GND.n6377 4.74817
R27832 GND.n6373 GND.n6372 4.74817
R27833 GND.n6368 GND.n6367 4.74817
R27834 GND.n6363 GND.n6362 4.74817
R27835 GND.n6340 GND.n5490 4.74817
R27836 GND.n5487 GND.n5486 4.74817
R27837 GND.n5482 GND.n5481 4.74817
R27838 GND.n5477 GND.n5476 4.74817
R27839 GND.n5472 GND.n5471 4.74817
R27840 GND.n5467 GND.n5466 4.74817
R27841 GND.n5173 GND.n122 4.74817
R27842 GND.n120 GND.n114 4.74817
R27843 GND.n10307 GND.n115 4.74817
R27844 GND.n123 GND.n119 4.74817
R27845 GND.n6918 GND.n122 4.74817
R27846 GND.n5188 GND.n120 4.74817
R27847 GND.n10308 GND.n10307 4.74817
R27848 GND.n5267 GND.n119 4.74817
R27849 GND.n3303 GND.n3302 4.74817
R27850 GND.n3332 GND.n3331 4.74817
R27851 GND.n3538 GND.n3537 4.74817
R27852 GND.n3533 GND.n3333 4.74817
R27853 GND.n3531 GND.n3530 4.74817
R27854 GND.n6747 GND.n5195 4.74817
R27855 GND.n6912 GND.n6911 4.74817
R27856 GND.n6907 GND.n5196 4.74817
R27857 GND.n6905 GND.n6904 4.74817
R27858 GND.n5264 GND.n5200 4.74817
R27859 GND.n6749 GND.n6747 4.74817
R27860 GND.n6913 GND.n6912 4.74817
R27861 GND.n6910 GND.n5196 4.74817
R27862 GND.n6906 GND.n6905 4.74817
R27863 GND.n5200 GND.n5198 4.74817
R27864 GND.n2621 GND.n1547 4.74817
R27865 GND.n1545 GND.n1539 4.74817
R27866 GND.n8120 GND.n1540 4.74817
R27867 GND.n1548 GND.n1544 4.74817
R27868 GND.n3322 GND.n1547 4.74817
R27869 GND.n3324 GND.n1545 4.74817
R27870 GND.n8121 GND.n8120 4.74817
R27871 GND.n3554 GND.n1544 4.74817
R27872 GND.n3302 GND.n2613 4.74817
R27873 GND.n3331 GND.n3330 4.74817
R27874 GND.n3539 GND.n3538 4.74817
R27875 GND.n3536 GND.n3333 4.74817
R27876 GND.n3532 GND.n3531 4.74817
R27877 GND.n3855 GND.n1682 4.74817
R27878 GND.n3856 GND.n3851 4.74817
R27879 GND.n3860 GND.n3850 4.74817
R27880 GND.n3864 GND.n3849 4.74817
R27881 GND.n3868 GND.n3848 4.74817
R27882 GND.n3859 GND.n3851 4.74817
R27883 GND.n3863 GND.n3850 4.74817
R27884 GND.n3867 GND.n3849 4.74817
R27885 GND.n3871 GND.n3848 4.74817
R27886 GND.n7715 GND.n7712 4.74817
R27887 GND.n7720 GND.n7717 4.74817
R27888 GND.n7725 GND.n7722 4.74817
R27889 GND.n7730 GND.n7727 4.74817
R27890 GND.n7735 GND.n7732 4.74817
R27891 GND.n7737 GND.n2357 4.74817
R27892 GND.n46 GND.n6 4.70093
R27893 GND.n101 GND.n100 4.70093
R27894 GND.n21 GND.n20 4.63843
R27895 GND.n29 GND.n28 4.63843
R27896 GND.n37 GND.n36 4.63843
R27897 GND.n45 GND.n44 4.63843
R27898 GND.n69 GND.n68 4.63843
R27899 GND.n77 GND.n76 4.63843
R27900 GND.n85 GND.n84 4.63843
R27901 GND.n93 GND.n92 4.63843
R27902 GND.n7187 GND.n4835 4.6132
R27903 GND.n7977 GND.n1869 4.6132
R27904 GND.n8023 GND.n1683 4.24068
R27905 GND.t4 GND.n4104 4.24068
R27906 GND.n5576 GND.t10 4.24068
R27907 GND.n7183 GND.n4869 4.24068
R27908 GND.n7708 GND.n7707 4.07323
R27909 GND.n6349 GND.n6344 4.07323
R27910 GND.n54 GND.n50 4.06868
R27911 GND.n4825 GND.n4762 4.05904
R27912 GND.n2130 GND.n2123 4.05904
R27913 GND.n7921 GND.n7920 4.05904
R27914 GND.n7198 GND.n7197 4.05904
R27915 GND.n7897 GND.t113 3.91451
R27916 GND.n7877 GND.n7876 3.91451
R27917 GND.n2007 GND.n2001 3.91451
R27918 GND.n2061 GND.n2055 3.91451
R27919 GND.n7800 GND.n7799 3.91451
R27920 GND.n5712 GND.n5690 3.91451
R27921 GND.t41 GND.n3903 3.91451
R27922 GND.n5816 GND.n5643 3.91451
R27923 GND.n7631 GND.n4007 3.91451
R27924 GND.n5919 GND.n5612 3.91451
R27925 GND.n7576 GND.n4112 3.91451
R27926 GND.n6022 GND.n5581 3.91451
R27927 GND.n7521 GND.n4216 3.91451
R27928 GND.n6125 GND.n5547 3.91451
R27929 GND.n7466 GND.n4319 3.91451
R27930 GND.n6220 GND.t152 3.91451
R27931 GND.n5499 GND.n5498 3.91451
R27932 GND.n4491 GND.n4485 3.91451
R27933 GND.n7352 GND.n7351 3.91451
R27934 GND.n4577 GND.n4571 3.91451
R27935 GND.n7291 GND.n7290 3.91451
R27936 GND.n54 GND.n53 3.53792
R27937 GND.n6386 GND.n6385 3.31114
R27938 GND.n3873 GND.n3872 3.31114
R27939 GND.n1842 GND.n1841 3.29747
R27940 GND.n1841 GND.n1840 3.29747
R27941 GND.n5426 GND.n5423 3.29747
R27942 GND.n5427 GND.n5426 3.29747
R27943 GND.n10001 GND.n9851 3.29747
R27944 GND.n10004 GND.n10001 3.29747
R27945 GND.n8268 GND.n8267 3.29747
R27946 GND.n8267 GND.n8266 3.29747
R27947 GND.n1938 GND.t79 3.26218
R27948 GND.n5628 GND.t1 3.26218
R27949 GND.n7484 GND.t272 3.26218
R27950 GND.n7264 GND.t61 3.26218
R27951 GND.n6386 GND.n6357 2.99593
R27952 GND.n3874 GND.n3873 2.99593
R27953 GND.n7972 GND.n1905 2.93601
R27954 GND.n5721 GND.t8 2.93601
R27955 GND.n6228 GND.t0 2.93601
R27956 GND.n7250 GND.n7249 2.93601
R27957 GND.n7911 GND.n7910 2.60984
R27958 GND.n7883 GND.n1973 2.60984
R27959 GND.n2240 GND.n2237 2.60984
R27960 GND.n2265 GND.n2262 2.60984
R27961 GND.n7793 GND.n2089 2.60984
R27962 GND.n5703 GND.n5694 2.60984
R27963 GND.n7680 GND.n3913 2.60984
R27964 GND.n5807 GND.n5797 2.60984
R27965 GND.n7625 GND.n4017 2.60984
R27966 GND.n5910 GND.n5901 2.60984
R27967 GND.n7570 GND.n4122 2.60984
R27968 GND.n6013 GND.n6004 2.60984
R27969 GND.n7515 GND.n4226 2.60984
R27970 GND.n6116 GND.n6107 2.60984
R27971 GND.n7460 GND.n4329 2.60984
R27972 GND.n6209 GND.n6203 2.60984
R27973 GND.n6303 GND.n6302 2.60984
R27974 GND.n6279 GND.n6276 2.60984
R27975 GND.n7345 GND.n4519 2.60984
R27976 GND.n4635 GND.n4632 2.60984
R27977 GND.n7284 GND.n4605 2.60984
R27978 GND.t125 GND.n7257 2.60984
R27979 GND.n4772 GND.n4768 2.60984
R27980 GND.n7710 GND.n7708 2.52171
R27981 GND.n6352 GND.n6344 2.52171
R27982 GND GND.n47 2.45421
R27983 GND.t22 GND.n2378 2.28367
R27984 GND.t8 GND.n5685 2.28367
R27985 GND.t20 GND.n7655 2.28367
R27986 GND.n6172 GND.t7 2.28367
R27987 GND.n7417 GND.t0 2.28367
R27988 GND.n6472 GND.t45 2.28367
R27989 GND.n6382 GND.n6357 2.27742
R27990 GND.n6377 GND.n6357 2.27742
R27991 GND.n6372 GND.n6357 2.27742
R27992 GND.n6367 GND.n6357 2.27742
R27993 GND.n6362 GND.n6357 2.27742
R27994 GND.n6356 GND.n6340 2.27742
R27995 GND.n6356 GND.n5486 2.27742
R27996 GND.n6356 GND.n5481 2.27742
R27997 GND.n6356 GND.n5476 2.27742
R27998 GND.n6356 GND.n5471 2.27742
R27999 GND.n6356 GND.n5466 2.27742
R28000 GND.n10306 GND.n122 2.27742
R28001 GND.n10306 GND.n120 2.27742
R28002 GND.n10307 GND.n10306 2.27742
R28003 GND.n10306 GND.n119 2.27742
R28004 GND.n6747 GND.n118 2.27742
R28005 GND.n6912 GND.n118 2.27742
R28006 GND.n5196 GND.n118 2.27742
R28007 GND.n6905 GND.n118 2.27742
R28008 GND.n5200 GND.n118 2.27742
R28009 GND.n8119 GND.n1547 2.27742
R28010 GND.n8119 GND.n1545 2.27742
R28011 GND.n8120 GND.n8119 2.27742
R28012 GND.n8119 GND.n1544 2.27742
R28013 GND.n3302 GND.n1543 2.27742
R28014 GND.n3331 GND.n1543 2.27742
R28015 GND.n3538 GND.n1543 2.27742
R28016 GND.n3333 GND.n1543 2.27742
R28017 GND.n3531 GND.n1543 2.27742
R28018 GND.n3874 GND.n1682 2.27742
R28019 GND.n3874 GND.n3851 2.27742
R28020 GND.n3874 GND.n3850 2.27742
R28021 GND.n3874 GND.n3849 2.27742
R28022 GND.n3874 GND.n3848 2.27742
R28023 GND.n7738 GND.n7712 2.27742
R28024 GND.n7738 GND.n7717 2.27742
R28025 GND.n7738 GND.n7722 2.27742
R28026 GND.n7738 GND.n7727 2.27742
R28027 GND.n7738 GND.n7732 2.27742
R28028 GND.n7738 GND.n7737 2.27742
R28029 GND.n1929 GND.n1911 2.19141
R28030 GND.n1924 GND.n1923 2.19141
R28031 GND.n4741 GND.n4736 2.19141
R28032 GND.n4743 GND.n4734 2.19141
R28033 GND.n7759 GND.n2341 1.95751
R28034 GND.n7655 GND.t270 1.95751
R28035 GND.n6172 GND.t15 1.95751
R28036 GND.n7408 GND.n4422 1.95751
R28037 GND.n10316 GND.n10315 1.89914
R28038 GND.n13 GND.n12 1.63556
R28039 GND.n12 GND.n10 1.63556
R28040 GND.n10 GND.n8 1.63556
R28041 GND.n20 GND.n19 1.63556
R28042 GND.n19 GND.n17 1.63556
R28043 GND.n17 GND.n15 1.63556
R28044 GND.n28 GND.n27 1.63556
R28045 GND.n27 GND.n25 1.63556
R28046 GND.n25 GND.n23 1.63556
R28047 GND.n36 GND.n35 1.63556
R28048 GND.n35 GND.n33 1.63556
R28049 GND.n33 GND.n31 1.63556
R28050 GND.n44 GND.n43 1.63556
R28051 GND.n43 GND.n41 1.63556
R28052 GND.n41 GND.n39 1.63556
R28053 GND.n6 GND.n5 1.63556
R28054 GND.n5 GND.n3 1.63556
R28055 GND.n3 GND.n1 1.63556
R28056 GND.n58 GND.n56 1.63556
R28057 GND.n60 GND.n58 1.63556
R28058 GND.n61 GND.n60 1.63556
R28059 GND.n65 GND.n63 1.63556
R28060 GND.n67 GND.n65 1.63556
R28061 GND.n68 GND.n67 1.63556
R28062 GND.n73 GND.n71 1.63556
R28063 GND.n75 GND.n73 1.63556
R28064 GND.n76 GND.n75 1.63556
R28065 GND.n81 GND.n79 1.63556
R28066 GND.n83 GND.n81 1.63556
R28067 GND.n84 GND.n83 1.63556
R28068 GND.n89 GND.n87 1.63556
R28069 GND.n91 GND.n89 1.63556
R28070 GND.n92 GND.n91 1.63556
R28071 GND.n97 GND.n95 1.63556
R28072 GND.n99 GND.n97 1.63556
R28073 GND.n100 GND.n99 1.63556
R28074 GND.n3044 GND.t187 1.63134
R28075 GND.n3122 GND.t194 1.63134
R28076 GND.t167 GND.n2540 1.63134
R28077 GND.n3675 GND.t165 1.63134
R28078 GND.n6639 GND.t155 1.63134
R28079 GND.t177 GND.n5116 1.63134
R28080 GND.n10231 GND.t161 1.63134
R28081 GND.t181 GND.n316 1.63134
R28082 GND.n4751 GND.n4733 1.55202
R28083 GND.n2186 GND.t128 1.30517
R28084 GND.n7904 GND.n1947 1.30517
R28085 GND.n7891 GND.n7890 1.30517
R28086 GND.n2025 GND.n2019 1.30517
R28087 GND.n2043 GND.n2037 1.30517
R28088 GND.n7786 GND.n7785 1.30517
R28089 GND.n2314 GND.n2305 1.30517
R28090 GND.n7674 GND.n3923 1.30517
R28091 GND.n3950 GND.n3944 1.30517
R28092 GND.n7619 GND.n4027 1.30517
R28093 GND.n4054 GND.n4048 1.30517
R28094 GND.n7564 GND.n4132 1.30517
R28095 GND.n4159 GND.n4153 1.30517
R28096 GND.n7509 GND.n4235 1.30517
R28097 GND.n4262 GND.n4256 1.30517
R28098 GND.n7454 GND.n4339 1.30517
R28099 GND.n4366 GND.n4360 1.30517
R28100 GND.n4455 GND.n4449 1.30517
R28101 GND.n4473 GND.n4467 1.30517
R28102 GND.n7338 GND.n7337 1.30517
R28103 GND.n4556 GND.n4547 1.30517
R28104 GND.n7277 GND.n7276 1.30517
R28105 GND.n4687 GND.n4676 1.30517
R28106 GND.n46 GND.n45 1.23398
R28107 GND.n101 GND.n93 1.23398
R28108 GND.n7986 GND.n7985 0.970197
R28109 GND.n7137 GND.n7124 0.970197
R28110 GND.n9943 GND.n9940 0.970197
R28111 GND.n8316 GND.n1391 0.970197
R28112 GND.n29 GND.n21 0.894178
R28113 GND.n37 GND.n29 0.894178
R28114 GND.n45 GND.n37 0.894178
R28115 GND.n77 GND.n69 0.894178
R28116 GND.n85 GND.n77 0.894178
R28117 GND.n93 GND.n85 0.894178
R28118 GND.n49 GND.n48 0.857089
R28119 GND.n50 GND.n49 0.857089
R28120 GND.n52 GND.n51 0.857089
R28121 GND.n53 GND.n52 0.857089
R28122 GND.n7277 GND.t49 0.652835
R28123 GND.n10079 GND.n10078 0.479159
R28124 GND.n8218 GND.n8217 0.479158
R28125 GND.n9885 GND.n413 0.471537
R28126 GND.n7096 GND.n7095 0.471537
R28127 GND.n8020 GND.n1724 0.471537
R28128 GND.n2939 GND.n1363 0.471537
R28129 GND.n1190 GND.n1185 0.459341
R28130 GND.n9525 GND.n9524 0.459341
R28131 GND.n9687 GND.n9686 0.459341
R28132 GND.n3010 GND.n1320 0.459341
R28133 GND.n6357 GND.n6356 0.456324
R28134 GND.n7738 GND.n3874 0.456324
R28135 GND.n6191 GND.n5495 0.436476
R28136 GND.n5671 GND.n2345 0.436476
R28137 GND.n7701 GND.n7700 0.436476
R28138 GND.n7413 GND.n7412 0.436476
R28139 GND.n10306 GND.n118 0.394875
R28140 GND.n8119 GND.n1543 0.394875
R28141 GND.t17 GND.n7834 0.326668
R28142 GND.t6 GND.n4529 0.326668
R28143 GND.n10316 GND.n54 0.305843
R28144 GND GND.n10316 0.279993
R28145 GND.n10050 GND.n420 0.27489
R28146 GND.n8239 GND.n8238 0.27489
R28147 GND.n3874 GND.n3847 0.267268
R28148 GND.n6419 GND.n6357 0.267268
R28149 GND.n10036 GND.n420 0.267268
R28150 GND.n5463 GND.n5462 0.267268
R28151 GND.n8240 GND.n8239 0.267268
R28152 GND.n1820 GND.n1673 0.267268
R28153 GND.n7128 GND.n4835 0.229039
R28154 GND.n4836 GND.n4835 0.229039
R28155 GND.n1869 GND.n1765 0.229039
R28156 GND.n1869 GND.n1868 0.229039
R28157 GND.n2592 GND.n1530 0.152939
R28158 GND.n2593 GND.n2592 0.152939
R28159 GND.n2593 GND.n2591 0.152939
R28160 GND.n3563 GND.n2591 0.152939
R28161 GND.n3564 GND.n3563 0.152939
R28162 GND.n3565 GND.n3564 0.152939
R28163 GND.n3566 GND.n3565 0.152939
R28164 GND.n3566 GND.n2569 0.152939
R28165 GND.n3588 GND.n2569 0.152939
R28166 GND.n3589 GND.n3588 0.152939
R28167 GND.n3590 GND.n3589 0.152939
R28168 GND.n3591 GND.n3590 0.152939
R28169 GND.n3591 GND.n2547 0.152939
R28170 GND.n3614 GND.n2547 0.152939
R28171 GND.n3615 GND.n3614 0.152939
R28172 GND.n3616 GND.n3615 0.152939
R28173 GND.n3617 GND.n3616 0.152939
R28174 GND.n3617 GND.n2526 0.152939
R28175 GND.n3640 GND.n2526 0.152939
R28176 GND.n3641 GND.n3640 0.152939
R28177 GND.n3642 GND.n3641 0.152939
R28178 GND.n3643 GND.n3642 0.152939
R28179 GND.n3643 GND.n2505 0.152939
R28180 GND.n3666 GND.n2505 0.152939
R28181 GND.n3667 GND.n3666 0.152939
R28182 GND.n3668 GND.n3667 0.152939
R28183 GND.n3669 GND.n3668 0.152939
R28184 GND.n3669 GND.n2482 0.152939
R28185 GND.n3691 GND.n2482 0.152939
R28186 GND.n3692 GND.n3691 0.152939
R28187 GND.n3693 GND.n3692 0.152939
R28188 GND.n3694 GND.n3693 0.152939
R28189 GND.n3694 GND.n2460 0.152939
R28190 GND.n3717 GND.n2460 0.152939
R28191 GND.n3718 GND.n3717 0.152939
R28192 GND.n3719 GND.n3718 0.152939
R28193 GND.n3720 GND.n3719 0.152939
R28194 GND.n3720 GND.n2441 0.152939
R28195 GND.n3743 GND.n2441 0.152939
R28196 GND.n3744 GND.n3743 0.152939
R28197 GND.n3745 GND.n3744 0.152939
R28198 GND.n3746 GND.n3745 0.152939
R28199 GND.n3746 GND.n2420 0.152939
R28200 GND.n3769 GND.n2420 0.152939
R28201 GND.n3770 GND.n3769 0.152939
R28202 GND.n3771 GND.n3770 0.152939
R28203 GND.n3772 GND.n3771 0.152939
R28204 GND.n3772 GND.n2397 0.152939
R28205 GND.n3794 GND.n2397 0.152939
R28206 GND.n3795 GND.n3794 0.152939
R28207 GND.n3796 GND.n3795 0.152939
R28208 GND.n3797 GND.n3796 0.152939
R28209 GND.n3797 GND.n2375 0.152939
R28210 GND.n3820 GND.n2375 0.152939
R28211 GND.n3821 GND.n3820 0.152939
R28212 GND.n3822 GND.n3821 0.152939
R28213 GND.n3824 GND.n3822 0.152939
R28214 GND.n3824 GND.n3823 0.152939
R28215 GND.n3823 GND.n2359 0.152939
R28216 GND.n3847 GND.n2359 0.152939
R28217 GND.n8502 GND.n1185 0.152939
R28218 GND.n8503 GND.n8502 0.152939
R28219 GND.n8504 GND.n8503 0.152939
R28220 GND.n8504 GND.n1179 0.152939
R28221 GND.n8512 GND.n1179 0.152939
R28222 GND.n8513 GND.n8512 0.152939
R28223 GND.n8514 GND.n8513 0.152939
R28224 GND.n8514 GND.n1173 0.152939
R28225 GND.n8522 GND.n1173 0.152939
R28226 GND.n8523 GND.n8522 0.152939
R28227 GND.n8524 GND.n8523 0.152939
R28228 GND.n8524 GND.n1167 0.152939
R28229 GND.n8532 GND.n1167 0.152939
R28230 GND.n8533 GND.n8532 0.152939
R28231 GND.n8534 GND.n8533 0.152939
R28232 GND.n8534 GND.n1161 0.152939
R28233 GND.n8542 GND.n1161 0.152939
R28234 GND.n8543 GND.n8542 0.152939
R28235 GND.n8544 GND.n8543 0.152939
R28236 GND.n8544 GND.n1155 0.152939
R28237 GND.n8552 GND.n1155 0.152939
R28238 GND.n8553 GND.n8552 0.152939
R28239 GND.n8554 GND.n8553 0.152939
R28240 GND.n8554 GND.n1149 0.152939
R28241 GND.n8562 GND.n1149 0.152939
R28242 GND.n8563 GND.n8562 0.152939
R28243 GND.n8564 GND.n8563 0.152939
R28244 GND.n8564 GND.n1143 0.152939
R28245 GND.n8572 GND.n1143 0.152939
R28246 GND.n8573 GND.n8572 0.152939
R28247 GND.n8574 GND.n8573 0.152939
R28248 GND.n8574 GND.n1137 0.152939
R28249 GND.n8582 GND.n1137 0.152939
R28250 GND.n8583 GND.n8582 0.152939
R28251 GND.n8584 GND.n8583 0.152939
R28252 GND.n8584 GND.n1131 0.152939
R28253 GND.n8592 GND.n1131 0.152939
R28254 GND.n8593 GND.n8592 0.152939
R28255 GND.n8594 GND.n8593 0.152939
R28256 GND.n8594 GND.n1125 0.152939
R28257 GND.n8602 GND.n1125 0.152939
R28258 GND.n8603 GND.n8602 0.152939
R28259 GND.n8604 GND.n8603 0.152939
R28260 GND.n8604 GND.n1119 0.152939
R28261 GND.n8612 GND.n1119 0.152939
R28262 GND.n8613 GND.n8612 0.152939
R28263 GND.n8614 GND.n8613 0.152939
R28264 GND.n8614 GND.n1113 0.152939
R28265 GND.n8622 GND.n1113 0.152939
R28266 GND.n8623 GND.n8622 0.152939
R28267 GND.n8624 GND.n8623 0.152939
R28268 GND.n8624 GND.n1107 0.152939
R28269 GND.n8632 GND.n1107 0.152939
R28270 GND.n8633 GND.n8632 0.152939
R28271 GND.n8634 GND.n8633 0.152939
R28272 GND.n8634 GND.n1101 0.152939
R28273 GND.n8642 GND.n1101 0.152939
R28274 GND.n8643 GND.n8642 0.152939
R28275 GND.n8644 GND.n8643 0.152939
R28276 GND.n8644 GND.n1095 0.152939
R28277 GND.n8652 GND.n1095 0.152939
R28278 GND.n8653 GND.n8652 0.152939
R28279 GND.n8654 GND.n8653 0.152939
R28280 GND.n8654 GND.n1089 0.152939
R28281 GND.n8662 GND.n1089 0.152939
R28282 GND.n8663 GND.n8662 0.152939
R28283 GND.n8664 GND.n8663 0.152939
R28284 GND.n8664 GND.n1083 0.152939
R28285 GND.n8672 GND.n1083 0.152939
R28286 GND.n8673 GND.n8672 0.152939
R28287 GND.n8674 GND.n8673 0.152939
R28288 GND.n8674 GND.n1077 0.152939
R28289 GND.n8682 GND.n1077 0.152939
R28290 GND.n8683 GND.n8682 0.152939
R28291 GND.n8684 GND.n8683 0.152939
R28292 GND.n8684 GND.n1071 0.152939
R28293 GND.n8692 GND.n1071 0.152939
R28294 GND.n8693 GND.n8692 0.152939
R28295 GND.n8694 GND.n8693 0.152939
R28296 GND.n8694 GND.n1065 0.152939
R28297 GND.n8702 GND.n1065 0.152939
R28298 GND.n8703 GND.n8702 0.152939
R28299 GND.n8704 GND.n8703 0.152939
R28300 GND.n8704 GND.n1059 0.152939
R28301 GND.n8712 GND.n1059 0.152939
R28302 GND.n8713 GND.n8712 0.152939
R28303 GND.n8714 GND.n8713 0.152939
R28304 GND.n8714 GND.n1053 0.152939
R28305 GND.n8722 GND.n1053 0.152939
R28306 GND.n8723 GND.n8722 0.152939
R28307 GND.n8724 GND.n8723 0.152939
R28308 GND.n8724 GND.n1047 0.152939
R28309 GND.n8732 GND.n1047 0.152939
R28310 GND.n8733 GND.n8732 0.152939
R28311 GND.n8734 GND.n8733 0.152939
R28312 GND.n8734 GND.n1041 0.152939
R28313 GND.n8742 GND.n1041 0.152939
R28314 GND.n8743 GND.n8742 0.152939
R28315 GND.n8744 GND.n8743 0.152939
R28316 GND.n8744 GND.n1035 0.152939
R28317 GND.n8752 GND.n1035 0.152939
R28318 GND.n8753 GND.n8752 0.152939
R28319 GND.n8754 GND.n8753 0.152939
R28320 GND.n8754 GND.n1029 0.152939
R28321 GND.n8762 GND.n1029 0.152939
R28322 GND.n8763 GND.n8762 0.152939
R28323 GND.n8764 GND.n8763 0.152939
R28324 GND.n8764 GND.n1023 0.152939
R28325 GND.n8772 GND.n1023 0.152939
R28326 GND.n8773 GND.n8772 0.152939
R28327 GND.n8774 GND.n8773 0.152939
R28328 GND.n8774 GND.n1017 0.152939
R28329 GND.n8782 GND.n1017 0.152939
R28330 GND.n8783 GND.n8782 0.152939
R28331 GND.n8784 GND.n8783 0.152939
R28332 GND.n8784 GND.n1011 0.152939
R28333 GND.n8792 GND.n1011 0.152939
R28334 GND.n8793 GND.n8792 0.152939
R28335 GND.n8794 GND.n8793 0.152939
R28336 GND.n8794 GND.n1005 0.152939
R28337 GND.n8802 GND.n1005 0.152939
R28338 GND.n8803 GND.n8802 0.152939
R28339 GND.n8804 GND.n8803 0.152939
R28340 GND.n8804 GND.n999 0.152939
R28341 GND.n8812 GND.n999 0.152939
R28342 GND.n8813 GND.n8812 0.152939
R28343 GND.n8814 GND.n8813 0.152939
R28344 GND.n8814 GND.n993 0.152939
R28345 GND.n8822 GND.n993 0.152939
R28346 GND.n8823 GND.n8822 0.152939
R28347 GND.n8824 GND.n8823 0.152939
R28348 GND.n8824 GND.n987 0.152939
R28349 GND.n8832 GND.n987 0.152939
R28350 GND.n8833 GND.n8832 0.152939
R28351 GND.n8834 GND.n8833 0.152939
R28352 GND.n8834 GND.n981 0.152939
R28353 GND.n8842 GND.n981 0.152939
R28354 GND.n8843 GND.n8842 0.152939
R28355 GND.n8844 GND.n8843 0.152939
R28356 GND.n8844 GND.n975 0.152939
R28357 GND.n8852 GND.n975 0.152939
R28358 GND.n8853 GND.n8852 0.152939
R28359 GND.n8854 GND.n8853 0.152939
R28360 GND.n8854 GND.n969 0.152939
R28361 GND.n8862 GND.n969 0.152939
R28362 GND.n8863 GND.n8862 0.152939
R28363 GND.n8864 GND.n8863 0.152939
R28364 GND.n8864 GND.n963 0.152939
R28365 GND.n8872 GND.n963 0.152939
R28366 GND.n8873 GND.n8872 0.152939
R28367 GND.n8874 GND.n8873 0.152939
R28368 GND.n8874 GND.n957 0.152939
R28369 GND.n8882 GND.n957 0.152939
R28370 GND.n8883 GND.n8882 0.152939
R28371 GND.n8884 GND.n8883 0.152939
R28372 GND.n8884 GND.n951 0.152939
R28373 GND.n8892 GND.n951 0.152939
R28374 GND.n8893 GND.n8892 0.152939
R28375 GND.n8894 GND.n8893 0.152939
R28376 GND.n8894 GND.n945 0.152939
R28377 GND.n8902 GND.n945 0.152939
R28378 GND.n8903 GND.n8902 0.152939
R28379 GND.n8904 GND.n8903 0.152939
R28380 GND.n8904 GND.n939 0.152939
R28381 GND.n8912 GND.n939 0.152939
R28382 GND.n8913 GND.n8912 0.152939
R28383 GND.n8914 GND.n8913 0.152939
R28384 GND.n8914 GND.n933 0.152939
R28385 GND.n8922 GND.n933 0.152939
R28386 GND.n8923 GND.n8922 0.152939
R28387 GND.n8924 GND.n8923 0.152939
R28388 GND.n8924 GND.n927 0.152939
R28389 GND.n8932 GND.n927 0.152939
R28390 GND.n8933 GND.n8932 0.152939
R28391 GND.n8934 GND.n8933 0.152939
R28392 GND.n8934 GND.n921 0.152939
R28393 GND.n8942 GND.n921 0.152939
R28394 GND.n8943 GND.n8942 0.152939
R28395 GND.n8944 GND.n8943 0.152939
R28396 GND.n8944 GND.n915 0.152939
R28397 GND.n8952 GND.n915 0.152939
R28398 GND.n8953 GND.n8952 0.152939
R28399 GND.n8954 GND.n8953 0.152939
R28400 GND.n8954 GND.n909 0.152939
R28401 GND.n8962 GND.n909 0.152939
R28402 GND.n8963 GND.n8962 0.152939
R28403 GND.n8964 GND.n8963 0.152939
R28404 GND.n8964 GND.n903 0.152939
R28405 GND.n8972 GND.n903 0.152939
R28406 GND.n8973 GND.n8972 0.152939
R28407 GND.n8974 GND.n8973 0.152939
R28408 GND.n8974 GND.n897 0.152939
R28409 GND.n8982 GND.n897 0.152939
R28410 GND.n8983 GND.n8982 0.152939
R28411 GND.n8984 GND.n8983 0.152939
R28412 GND.n8984 GND.n891 0.152939
R28413 GND.n8992 GND.n891 0.152939
R28414 GND.n8993 GND.n8992 0.152939
R28415 GND.n8994 GND.n8993 0.152939
R28416 GND.n8994 GND.n885 0.152939
R28417 GND.n9002 GND.n885 0.152939
R28418 GND.n9003 GND.n9002 0.152939
R28419 GND.n9004 GND.n9003 0.152939
R28420 GND.n9004 GND.n879 0.152939
R28421 GND.n9012 GND.n879 0.152939
R28422 GND.n9013 GND.n9012 0.152939
R28423 GND.n9014 GND.n9013 0.152939
R28424 GND.n9014 GND.n873 0.152939
R28425 GND.n9022 GND.n873 0.152939
R28426 GND.n9023 GND.n9022 0.152939
R28427 GND.n9024 GND.n9023 0.152939
R28428 GND.n9024 GND.n867 0.152939
R28429 GND.n9032 GND.n867 0.152939
R28430 GND.n9033 GND.n9032 0.152939
R28431 GND.n9034 GND.n9033 0.152939
R28432 GND.n9034 GND.n861 0.152939
R28433 GND.n9042 GND.n861 0.152939
R28434 GND.n9043 GND.n9042 0.152939
R28435 GND.n9044 GND.n9043 0.152939
R28436 GND.n9044 GND.n855 0.152939
R28437 GND.n9052 GND.n855 0.152939
R28438 GND.n9053 GND.n9052 0.152939
R28439 GND.n9054 GND.n9053 0.152939
R28440 GND.n9054 GND.n849 0.152939
R28441 GND.n9062 GND.n849 0.152939
R28442 GND.n9063 GND.n9062 0.152939
R28443 GND.n9064 GND.n9063 0.152939
R28444 GND.n9064 GND.n843 0.152939
R28445 GND.n9072 GND.n843 0.152939
R28446 GND.n9073 GND.n9072 0.152939
R28447 GND.n9074 GND.n9073 0.152939
R28448 GND.n9074 GND.n837 0.152939
R28449 GND.n9082 GND.n837 0.152939
R28450 GND.n9083 GND.n9082 0.152939
R28451 GND.n9084 GND.n9083 0.152939
R28452 GND.n9084 GND.n831 0.152939
R28453 GND.n9092 GND.n831 0.152939
R28454 GND.n9093 GND.n9092 0.152939
R28455 GND.n9094 GND.n9093 0.152939
R28456 GND.n9094 GND.n825 0.152939
R28457 GND.n9102 GND.n825 0.152939
R28458 GND.n9103 GND.n9102 0.152939
R28459 GND.n9104 GND.n9103 0.152939
R28460 GND.n9104 GND.n819 0.152939
R28461 GND.n9112 GND.n819 0.152939
R28462 GND.n9113 GND.n9112 0.152939
R28463 GND.n9114 GND.n9113 0.152939
R28464 GND.n9114 GND.n813 0.152939
R28465 GND.n9122 GND.n813 0.152939
R28466 GND.n9123 GND.n9122 0.152939
R28467 GND.n9124 GND.n9123 0.152939
R28468 GND.n9124 GND.n807 0.152939
R28469 GND.n9132 GND.n807 0.152939
R28470 GND.n9133 GND.n9132 0.152939
R28471 GND.n9134 GND.n9133 0.152939
R28472 GND.n9134 GND.n801 0.152939
R28473 GND.n9142 GND.n801 0.152939
R28474 GND.n9143 GND.n9142 0.152939
R28475 GND.n9144 GND.n9143 0.152939
R28476 GND.n9144 GND.n795 0.152939
R28477 GND.n9152 GND.n795 0.152939
R28478 GND.n9153 GND.n9152 0.152939
R28479 GND.n9154 GND.n9153 0.152939
R28480 GND.n9154 GND.n789 0.152939
R28481 GND.n9162 GND.n789 0.152939
R28482 GND.n9163 GND.n9162 0.152939
R28483 GND.n9164 GND.n9163 0.152939
R28484 GND.n9164 GND.n783 0.152939
R28485 GND.n9172 GND.n783 0.152939
R28486 GND.n9173 GND.n9172 0.152939
R28487 GND.n9174 GND.n9173 0.152939
R28488 GND.n9174 GND.n777 0.152939
R28489 GND.n9182 GND.n777 0.152939
R28490 GND.n9183 GND.n9182 0.152939
R28491 GND.n9184 GND.n9183 0.152939
R28492 GND.n9184 GND.n771 0.152939
R28493 GND.n9192 GND.n771 0.152939
R28494 GND.n9193 GND.n9192 0.152939
R28495 GND.n9194 GND.n9193 0.152939
R28496 GND.n9194 GND.n765 0.152939
R28497 GND.n9202 GND.n765 0.152939
R28498 GND.n9203 GND.n9202 0.152939
R28499 GND.n9204 GND.n9203 0.152939
R28500 GND.n9204 GND.n759 0.152939
R28501 GND.n9212 GND.n759 0.152939
R28502 GND.n9213 GND.n9212 0.152939
R28503 GND.n9214 GND.n9213 0.152939
R28504 GND.n9214 GND.n753 0.152939
R28505 GND.n9222 GND.n753 0.152939
R28506 GND.n9223 GND.n9222 0.152939
R28507 GND.n9224 GND.n9223 0.152939
R28508 GND.n9224 GND.n747 0.152939
R28509 GND.n9232 GND.n747 0.152939
R28510 GND.n9233 GND.n9232 0.152939
R28511 GND.n9234 GND.n9233 0.152939
R28512 GND.n9234 GND.n741 0.152939
R28513 GND.n9242 GND.n741 0.152939
R28514 GND.n9243 GND.n9242 0.152939
R28515 GND.n9244 GND.n9243 0.152939
R28516 GND.n9244 GND.n735 0.152939
R28517 GND.n9252 GND.n735 0.152939
R28518 GND.n9253 GND.n9252 0.152939
R28519 GND.n9254 GND.n9253 0.152939
R28520 GND.n9254 GND.n729 0.152939
R28521 GND.n9262 GND.n729 0.152939
R28522 GND.n9263 GND.n9262 0.152939
R28523 GND.n9264 GND.n9263 0.152939
R28524 GND.n9264 GND.n723 0.152939
R28525 GND.n9272 GND.n723 0.152939
R28526 GND.n9273 GND.n9272 0.152939
R28527 GND.n9274 GND.n9273 0.152939
R28528 GND.n9274 GND.n717 0.152939
R28529 GND.n9282 GND.n717 0.152939
R28530 GND.n9283 GND.n9282 0.152939
R28531 GND.n9284 GND.n9283 0.152939
R28532 GND.n9284 GND.n711 0.152939
R28533 GND.n9292 GND.n711 0.152939
R28534 GND.n9293 GND.n9292 0.152939
R28535 GND.n9294 GND.n9293 0.152939
R28536 GND.n9294 GND.n705 0.152939
R28537 GND.n9302 GND.n705 0.152939
R28538 GND.n9303 GND.n9302 0.152939
R28539 GND.n9304 GND.n9303 0.152939
R28540 GND.n9304 GND.n699 0.152939
R28541 GND.n9312 GND.n699 0.152939
R28542 GND.n9313 GND.n9312 0.152939
R28543 GND.n9314 GND.n9313 0.152939
R28544 GND.n9314 GND.n693 0.152939
R28545 GND.n9322 GND.n693 0.152939
R28546 GND.n9323 GND.n9322 0.152939
R28547 GND.n9324 GND.n9323 0.152939
R28548 GND.n9324 GND.n687 0.152939
R28549 GND.n9332 GND.n687 0.152939
R28550 GND.n9333 GND.n9332 0.152939
R28551 GND.n9334 GND.n9333 0.152939
R28552 GND.n9334 GND.n681 0.152939
R28553 GND.n9342 GND.n681 0.152939
R28554 GND.n9343 GND.n9342 0.152939
R28555 GND.n9344 GND.n9343 0.152939
R28556 GND.n9344 GND.n675 0.152939
R28557 GND.n9352 GND.n675 0.152939
R28558 GND.n9353 GND.n9352 0.152939
R28559 GND.n9354 GND.n9353 0.152939
R28560 GND.n9354 GND.n669 0.152939
R28561 GND.n9362 GND.n669 0.152939
R28562 GND.n9363 GND.n9362 0.152939
R28563 GND.n9364 GND.n9363 0.152939
R28564 GND.n9364 GND.n663 0.152939
R28565 GND.n9372 GND.n663 0.152939
R28566 GND.n9373 GND.n9372 0.152939
R28567 GND.n9374 GND.n9373 0.152939
R28568 GND.n9374 GND.n657 0.152939
R28569 GND.n9382 GND.n657 0.152939
R28570 GND.n9383 GND.n9382 0.152939
R28571 GND.n9384 GND.n9383 0.152939
R28572 GND.n9384 GND.n651 0.152939
R28573 GND.n9392 GND.n651 0.152939
R28574 GND.n9393 GND.n9392 0.152939
R28575 GND.n9394 GND.n9393 0.152939
R28576 GND.n9394 GND.n645 0.152939
R28577 GND.n9402 GND.n645 0.152939
R28578 GND.n9403 GND.n9402 0.152939
R28579 GND.n9404 GND.n9403 0.152939
R28580 GND.n9404 GND.n639 0.152939
R28581 GND.n9412 GND.n639 0.152939
R28582 GND.n9413 GND.n9412 0.152939
R28583 GND.n9414 GND.n9413 0.152939
R28584 GND.n9414 GND.n633 0.152939
R28585 GND.n9422 GND.n633 0.152939
R28586 GND.n9423 GND.n9422 0.152939
R28587 GND.n9424 GND.n9423 0.152939
R28588 GND.n9424 GND.n627 0.152939
R28589 GND.n9432 GND.n627 0.152939
R28590 GND.n9433 GND.n9432 0.152939
R28591 GND.n9434 GND.n9433 0.152939
R28592 GND.n9434 GND.n621 0.152939
R28593 GND.n9442 GND.n621 0.152939
R28594 GND.n9443 GND.n9442 0.152939
R28595 GND.n9444 GND.n9443 0.152939
R28596 GND.n9444 GND.n615 0.152939
R28597 GND.n9452 GND.n615 0.152939
R28598 GND.n9453 GND.n9452 0.152939
R28599 GND.n9454 GND.n9453 0.152939
R28600 GND.n9454 GND.n609 0.152939
R28601 GND.n9462 GND.n609 0.152939
R28602 GND.n9463 GND.n9462 0.152939
R28603 GND.n9464 GND.n9463 0.152939
R28604 GND.n9464 GND.n603 0.152939
R28605 GND.n9472 GND.n603 0.152939
R28606 GND.n9473 GND.n9472 0.152939
R28607 GND.n9474 GND.n9473 0.152939
R28608 GND.n9474 GND.n597 0.152939
R28609 GND.n9482 GND.n597 0.152939
R28610 GND.n9483 GND.n9482 0.152939
R28611 GND.n9484 GND.n9483 0.152939
R28612 GND.n9484 GND.n591 0.152939
R28613 GND.n9492 GND.n591 0.152939
R28614 GND.n9493 GND.n9492 0.152939
R28615 GND.n9494 GND.n9493 0.152939
R28616 GND.n9494 GND.n585 0.152939
R28617 GND.n9502 GND.n585 0.152939
R28618 GND.n9503 GND.n9502 0.152939
R28619 GND.n9504 GND.n9503 0.152939
R28620 GND.n9504 GND.n579 0.152939
R28621 GND.n9512 GND.n579 0.152939
R28622 GND.n9513 GND.n9512 0.152939
R28623 GND.n9515 GND.n9513 0.152939
R28624 GND.n9515 GND.n9514 0.152939
R28625 GND.n9514 GND.n573 0.152939
R28626 GND.n9524 GND.n573 0.152939
R28627 GND.n9525 GND.n568 0.152939
R28628 GND.n9533 GND.n568 0.152939
R28629 GND.n9534 GND.n9533 0.152939
R28630 GND.n9535 GND.n9534 0.152939
R28631 GND.n9535 GND.n562 0.152939
R28632 GND.n9543 GND.n562 0.152939
R28633 GND.n9544 GND.n9543 0.152939
R28634 GND.n9545 GND.n9544 0.152939
R28635 GND.n9545 GND.n556 0.152939
R28636 GND.n9553 GND.n556 0.152939
R28637 GND.n9554 GND.n9553 0.152939
R28638 GND.n9555 GND.n9554 0.152939
R28639 GND.n9555 GND.n550 0.152939
R28640 GND.n9563 GND.n550 0.152939
R28641 GND.n9564 GND.n9563 0.152939
R28642 GND.n9565 GND.n9564 0.152939
R28643 GND.n9565 GND.n544 0.152939
R28644 GND.n9573 GND.n544 0.152939
R28645 GND.n9574 GND.n9573 0.152939
R28646 GND.n9575 GND.n9574 0.152939
R28647 GND.n9575 GND.n538 0.152939
R28648 GND.n9583 GND.n538 0.152939
R28649 GND.n9584 GND.n9583 0.152939
R28650 GND.n9585 GND.n9584 0.152939
R28651 GND.n9585 GND.n532 0.152939
R28652 GND.n9593 GND.n532 0.152939
R28653 GND.n9594 GND.n9593 0.152939
R28654 GND.n9595 GND.n9594 0.152939
R28655 GND.n9595 GND.n526 0.152939
R28656 GND.n9603 GND.n526 0.152939
R28657 GND.n9604 GND.n9603 0.152939
R28658 GND.n9605 GND.n9604 0.152939
R28659 GND.n9605 GND.n520 0.152939
R28660 GND.n9613 GND.n520 0.152939
R28661 GND.n9614 GND.n9613 0.152939
R28662 GND.n9615 GND.n9614 0.152939
R28663 GND.n9615 GND.n514 0.152939
R28664 GND.n9623 GND.n514 0.152939
R28665 GND.n9624 GND.n9623 0.152939
R28666 GND.n9625 GND.n9624 0.152939
R28667 GND.n9625 GND.n508 0.152939
R28668 GND.n9633 GND.n508 0.152939
R28669 GND.n9634 GND.n9633 0.152939
R28670 GND.n9635 GND.n9634 0.152939
R28671 GND.n9635 GND.n502 0.152939
R28672 GND.n9643 GND.n502 0.152939
R28673 GND.n9644 GND.n9643 0.152939
R28674 GND.n9645 GND.n9644 0.152939
R28675 GND.n9645 GND.n496 0.152939
R28676 GND.n9653 GND.n496 0.152939
R28677 GND.n9654 GND.n9653 0.152939
R28678 GND.n9655 GND.n9654 0.152939
R28679 GND.n9655 GND.n490 0.152939
R28680 GND.n9663 GND.n490 0.152939
R28681 GND.n9664 GND.n9663 0.152939
R28682 GND.n9665 GND.n9664 0.152939
R28683 GND.n9665 GND.n484 0.152939
R28684 GND.n9673 GND.n484 0.152939
R28685 GND.n9674 GND.n9673 0.152939
R28686 GND.n9675 GND.n9674 0.152939
R28687 GND.n9675 GND.n478 0.152939
R28688 GND.n9683 GND.n478 0.152939
R28689 GND.n9684 GND.n9683 0.152939
R28690 GND.n9685 GND.n9684 0.152939
R28691 GND.n9688 GND.n9685 0.152939
R28692 GND.n9688 GND.n9687 0.152939
R28693 GND.n5202 GND.n5201 0.152939
R28694 GND.n5205 GND.n5202 0.152939
R28695 GND.n5206 GND.n5205 0.152939
R28696 GND.n5207 GND.n5206 0.152939
R28697 GND.n5208 GND.n5207 0.152939
R28698 GND.n5211 GND.n5208 0.152939
R28699 GND.n5212 GND.n5211 0.152939
R28700 GND.n5213 GND.n5212 0.152939
R28701 GND.n5214 GND.n5213 0.152939
R28702 GND.n5217 GND.n5214 0.152939
R28703 GND.n5218 GND.n5217 0.152939
R28704 GND.n5219 GND.n5218 0.152939
R28705 GND.n5220 GND.n5219 0.152939
R28706 GND.n5223 GND.n5220 0.152939
R28707 GND.n5224 GND.n5223 0.152939
R28708 GND.n5225 GND.n5224 0.152939
R28709 GND.n5226 GND.n5225 0.152939
R28710 GND.n5229 GND.n5226 0.152939
R28711 GND.n5230 GND.n5229 0.152939
R28712 GND.n5232 GND.n5230 0.152939
R28713 GND.n5232 GND.n5231 0.152939
R28714 GND.n5231 GND.n445 0.152939
R28715 GND.n446 GND.n445 0.152939
R28716 GND.n447 GND.n446 0.152939
R28717 GND.n450 GND.n447 0.152939
R28718 GND.n451 GND.n450 0.152939
R28719 GND.n452 GND.n451 0.152939
R28720 GND.n453 GND.n452 0.152939
R28721 GND.n456 GND.n453 0.152939
R28722 GND.n457 GND.n456 0.152939
R28723 GND.n458 GND.n457 0.152939
R28724 GND.n459 GND.n458 0.152939
R28725 GND.n462 GND.n459 0.152939
R28726 GND.n463 GND.n462 0.152939
R28727 GND.n464 GND.n463 0.152939
R28728 GND.n465 GND.n464 0.152939
R28729 GND.n468 GND.n465 0.152939
R28730 GND.n469 GND.n468 0.152939
R28731 GND.n470 GND.n469 0.152939
R28732 GND.n471 GND.n470 0.152939
R28733 GND.n9686 GND.n471 0.152939
R28734 GND.n144 GND.n116 0.152939
R28735 GND.n145 GND.n144 0.152939
R28736 GND.n146 GND.n145 0.152939
R28737 GND.n164 GND.n146 0.152939
R28738 GND.n165 GND.n164 0.152939
R28739 GND.n166 GND.n165 0.152939
R28740 GND.n167 GND.n166 0.152939
R28741 GND.n185 GND.n167 0.152939
R28742 GND.n186 GND.n185 0.152939
R28743 GND.n187 GND.n186 0.152939
R28744 GND.n188 GND.n187 0.152939
R28745 GND.n206 GND.n188 0.152939
R28746 GND.n207 GND.n206 0.152939
R28747 GND.n208 GND.n207 0.152939
R28748 GND.n209 GND.n208 0.152939
R28749 GND.n227 GND.n209 0.152939
R28750 GND.n228 GND.n227 0.152939
R28751 GND.n229 GND.n228 0.152939
R28752 GND.n230 GND.n229 0.152939
R28753 GND.n248 GND.n230 0.152939
R28754 GND.n249 GND.n248 0.152939
R28755 GND.n250 GND.n249 0.152939
R28756 GND.n251 GND.n250 0.152939
R28757 GND.n268 GND.n251 0.152939
R28758 GND.n269 GND.n268 0.152939
R28759 GND.n270 GND.n269 0.152939
R28760 GND.n271 GND.n270 0.152939
R28761 GND.n289 GND.n271 0.152939
R28762 GND.n290 GND.n289 0.152939
R28763 GND.n291 GND.n290 0.152939
R28764 GND.n292 GND.n291 0.152939
R28765 GND.n310 GND.n292 0.152939
R28766 GND.n311 GND.n310 0.152939
R28767 GND.n312 GND.n311 0.152939
R28768 GND.n313 GND.n312 0.152939
R28769 GND.n331 GND.n313 0.152939
R28770 GND.n332 GND.n331 0.152939
R28771 GND.n333 GND.n332 0.152939
R28772 GND.n334 GND.n333 0.152939
R28773 GND.n352 GND.n334 0.152939
R28774 GND.n353 GND.n352 0.152939
R28775 GND.n354 GND.n353 0.152939
R28776 GND.n355 GND.n354 0.152939
R28777 GND.n372 GND.n355 0.152939
R28778 GND.n373 GND.n372 0.152939
R28779 GND.n374 GND.n373 0.152939
R28780 GND.n375 GND.n374 0.152939
R28781 GND.n391 GND.n375 0.152939
R28782 GND.n392 GND.n391 0.152939
R28783 GND.n393 GND.n392 0.152939
R28784 GND.n394 GND.n393 0.152939
R28785 GND.n410 GND.n394 0.152939
R28786 GND.n411 GND.n410 0.152939
R28787 GND.n412 GND.n411 0.152939
R28788 GND.n413 GND.n412 0.152939
R28789 GND.n5495 GND.n5494 0.152939
R28790 GND.n6320 GND.n5494 0.152939
R28791 GND.n6321 GND.n6320 0.152939
R28792 GND.n6322 GND.n6321 0.152939
R28793 GND.n6322 GND.n5492 0.152939
R28794 GND.n6330 GND.n5492 0.152939
R28795 GND.n6331 GND.n6330 0.152939
R28796 GND.n6332 GND.n6331 0.152939
R28797 GND.n6332 GND.n5464 0.152939
R28798 GND.n5682 GND.n5671 0.152939
R28799 GND.n5682 GND.n5681 0.152939
R28800 GND.n5681 GND.n5680 0.152939
R28801 GND.n5680 GND.n5672 0.152939
R28802 GND.n5674 GND.n5672 0.152939
R28803 GND.n5674 GND.n5673 0.152939
R28804 GND.n5673 GND.n5652 0.152939
R28805 GND.n5763 GND.n5652 0.152939
R28806 GND.n5764 GND.n5763 0.152939
R28807 GND.n5765 GND.n5764 0.152939
R28808 GND.n5765 GND.n5648 0.152939
R28809 GND.n5771 GND.n5648 0.152939
R28810 GND.n5772 GND.n5771 0.152939
R28811 GND.n5773 GND.n5772 0.152939
R28812 GND.n5774 GND.n5773 0.152939
R28813 GND.n5775 GND.n5774 0.152939
R28814 GND.n5776 GND.n5775 0.152939
R28815 GND.n5777 GND.n5776 0.152939
R28816 GND.n5778 GND.n5777 0.152939
R28817 GND.n5779 GND.n5778 0.152939
R28818 GND.n5780 GND.n5779 0.152939
R28819 GND.n5782 GND.n5780 0.152939
R28820 GND.n5782 GND.n5781 0.152939
R28821 GND.n5781 GND.n5621 0.152939
R28822 GND.n5867 GND.n5621 0.152939
R28823 GND.n5868 GND.n5867 0.152939
R28824 GND.n5869 GND.n5868 0.152939
R28825 GND.n5869 GND.n5617 0.152939
R28826 GND.n5875 GND.n5617 0.152939
R28827 GND.n5876 GND.n5875 0.152939
R28828 GND.n5877 GND.n5876 0.152939
R28829 GND.n5878 GND.n5877 0.152939
R28830 GND.n5879 GND.n5878 0.152939
R28831 GND.n5880 GND.n5879 0.152939
R28832 GND.n5881 GND.n5880 0.152939
R28833 GND.n5882 GND.n5881 0.152939
R28834 GND.n5883 GND.n5882 0.152939
R28835 GND.n5884 GND.n5883 0.152939
R28836 GND.n5886 GND.n5884 0.152939
R28837 GND.n5886 GND.n5885 0.152939
R28838 GND.n5885 GND.n5590 0.152939
R28839 GND.n5970 GND.n5590 0.152939
R28840 GND.n5971 GND.n5970 0.152939
R28841 GND.n5972 GND.n5971 0.152939
R28842 GND.n5972 GND.n5586 0.152939
R28843 GND.n5978 GND.n5586 0.152939
R28844 GND.n5979 GND.n5978 0.152939
R28845 GND.n5980 GND.n5979 0.152939
R28846 GND.n5981 GND.n5980 0.152939
R28847 GND.n5982 GND.n5981 0.152939
R28848 GND.n5983 GND.n5982 0.152939
R28849 GND.n5984 GND.n5983 0.152939
R28850 GND.n5985 GND.n5984 0.152939
R28851 GND.n5986 GND.n5985 0.152939
R28852 GND.n5987 GND.n5986 0.152939
R28853 GND.n5989 GND.n5987 0.152939
R28854 GND.n5989 GND.n5988 0.152939
R28855 GND.n5988 GND.n5557 0.152939
R28856 GND.n6073 GND.n5557 0.152939
R28857 GND.n6074 GND.n6073 0.152939
R28858 GND.n6075 GND.n6074 0.152939
R28859 GND.n6075 GND.n5553 0.152939
R28860 GND.n6081 GND.n5553 0.152939
R28861 GND.n6082 GND.n6081 0.152939
R28862 GND.n6083 GND.n6082 0.152939
R28863 GND.n6084 GND.n6083 0.152939
R28864 GND.n6085 GND.n6084 0.152939
R28865 GND.n6086 GND.n6085 0.152939
R28866 GND.n6087 GND.n6086 0.152939
R28867 GND.n6088 GND.n6087 0.152939
R28868 GND.n6089 GND.n6088 0.152939
R28869 GND.n6090 GND.n6089 0.152939
R28870 GND.n6092 GND.n6090 0.152939
R28871 GND.n6092 GND.n6091 0.152939
R28872 GND.n6091 GND.n5525 0.152939
R28873 GND.n6176 GND.n5525 0.152939
R28874 GND.n6177 GND.n6176 0.152939
R28875 GND.n6178 GND.n6177 0.152939
R28876 GND.n6178 GND.n5521 0.152939
R28877 GND.n6184 GND.n5521 0.152939
R28878 GND.n6185 GND.n6184 0.152939
R28879 GND.n6186 GND.n6185 0.152939
R28880 GND.n6187 GND.n6186 0.152939
R28881 GND.n6188 GND.n6187 0.152939
R28882 GND.n6189 GND.n6188 0.152939
R28883 GND.n6190 GND.n6189 0.152939
R28884 GND.n6192 GND.n6190 0.152939
R28885 GND.n6192 GND.n6191 0.152939
R28886 GND.n2346 GND.n2345 0.152939
R28887 GND.n2347 GND.n2346 0.152939
R28888 GND.n2348 GND.n2347 0.152939
R28889 GND.n2349 GND.n2348 0.152939
R28890 GND.n2350 GND.n2349 0.152939
R28891 GND.n2351 GND.n2350 0.152939
R28892 GND.n2352 GND.n2351 0.152939
R28893 GND.n2353 GND.n2352 0.152939
R28894 GND.n2354 GND.n2353 0.152939
R28895 GND.n3878 GND.n2358 0.152939
R28896 GND.n3879 GND.n3878 0.152939
R28897 GND.n7702 GND.n3879 0.152939
R28898 GND.n7702 GND.n7701 0.152939
R28899 GND.n7700 GND.n3882 0.152939
R28900 GND.n3898 GND.n3882 0.152939
R28901 GND.n3899 GND.n3898 0.152939
R28902 GND.n3900 GND.n3899 0.152939
R28903 GND.n3917 GND.n3900 0.152939
R28904 GND.n3918 GND.n3917 0.152939
R28905 GND.n3919 GND.n3918 0.152939
R28906 GND.n3920 GND.n3919 0.152939
R28907 GND.n3972 GND.n3920 0.152939
R28908 GND.n3973 GND.n3972 0.152939
R28909 GND.n3974 GND.n3973 0.152939
R28910 GND.n3974 GND.n3970 0.152939
R28911 GND.n3980 GND.n3970 0.152939
R28912 GND.n3981 GND.n3980 0.152939
R28913 GND.n3982 GND.n3981 0.152939
R28914 GND.n3983 GND.n3982 0.152939
R28915 GND.n3984 GND.n3983 0.152939
R28916 GND.n4001 GND.n3984 0.152939
R28917 GND.n4002 GND.n4001 0.152939
R28918 GND.n4003 GND.n4002 0.152939
R28919 GND.n4004 GND.n4003 0.152939
R28920 GND.n4021 GND.n4004 0.152939
R28921 GND.n4022 GND.n4021 0.152939
R28922 GND.n4023 GND.n4022 0.152939
R28923 GND.n4024 GND.n4023 0.152939
R28924 GND.n4077 GND.n4024 0.152939
R28925 GND.n4078 GND.n4077 0.152939
R28926 GND.n4079 GND.n4078 0.152939
R28927 GND.n4079 GND.n4075 0.152939
R28928 GND.n4085 GND.n4075 0.152939
R28929 GND.n4086 GND.n4085 0.152939
R28930 GND.n4087 GND.n4086 0.152939
R28931 GND.n4088 GND.n4087 0.152939
R28932 GND.n4089 GND.n4088 0.152939
R28933 GND.n4106 GND.n4089 0.152939
R28934 GND.n4107 GND.n4106 0.152939
R28935 GND.n4108 GND.n4107 0.152939
R28936 GND.n4109 GND.n4108 0.152939
R28937 GND.n4126 GND.n4109 0.152939
R28938 GND.n4127 GND.n4126 0.152939
R28939 GND.n4128 GND.n4127 0.152939
R28940 GND.n4129 GND.n4128 0.152939
R28941 GND.n4182 GND.n4129 0.152939
R28942 GND.n4183 GND.n4182 0.152939
R28943 GND.n4184 GND.n4183 0.152939
R28944 GND.n4184 GND.n4180 0.152939
R28945 GND.n4190 GND.n4180 0.152939
R28946 GND.n4191 GND.n4190 0.152939
R28947 GND.n4192 GND.n4191 0.152939
R28948 GND.n4193 GND.n4192 0.152939
R28949 GND.n4194 GND.n4193 0.152939
R28950 GND.n4210 GND.n4194 0.152939
R28951 GND.n4211 GND.n4210 0.152939
R28952 GND.n4212 GND.n4211 0.152939
R28953 GND.n4213 GND.n4212 0.152939
R28954 GND.n4229 GND.n4213 0.152939
R28955 GND.n4230 GND.n4229 0.152939
R28956 GND.n4231 GND.n4230 0.152939
R28957 GND.n4232 GND.n4231 0.152939
R28958 GND.n4284 GND.n4232 0.152939
R28959 GND.n4285 GND.n4284 0.152939
R28960 GND.n4286 GND.n4285 0.152939
R28961 GND.n4286 GND.n4282 0.152939
R28962 GND.n4292 GND.n4282 0.152939
R28963 GND.n4293 GND.n4292 0.152939
R28964 GND.n4294 GND.n4293 0.152939
R28965 GND.n4295 GND.n4294 0.152939
R28966 GND.n4296 GND.n4295 0.152939
R28967 GND.n4313 GND.n4296 0.152939
R28968 GND.n4314 GND.n4313 0.152939
R28969 GND.n4315 GND.n4314 0.152939
R28970 GND.n4316 GND.n4315 0.152939
R28971 GND.n4333 GND.n4316 0.152939
R28972 GND.n4334 GND.n4333 0.152939
R28973 GND.n4335 GND.n4334 0.152939
R28974 GND.n4336 GND.n4335 0.152939
R28975 GND.n4389 GND.n4336 0.152939
R28976 GND.n4390 GND.n4389 0.152939
R28977 GND.n4391 GND.n4390 0.152939
R28978 GND.n4391 GND.n4387 0.152939
R28979 GND.n4397 GND.n4387 0.152939
R28980 GND.n4398 GND.n4397 0.152939
R28981 GND.n4399 GND.n4398 0.152939
R28982 GND.n4400 GND.n4399 0.152939
R28983 GND.n4401 GND.n4400 0.152939
R28984 GND.n4417 GND.n4401 0.152939
R28985 GND.n4418 GND.n4417 0.152939
R28986 GND.n7413 GND.n4418 0.152939
R28987 GND.n6345 GND.n5465 0.152939
R28988 GND.n6346 GND.n6345 0.152939
R28989 GND.n6346 GND.n4419 0.152939
R28990 GND.n7412 GND.n4419 0.152939
R28991 GND.n6420 GND.n6419 0.152939
R28992 GND.n6421 GND.n6420 0.152939
R28993 GND.n6421 GND.n5364 0.152939
R28994 GND.n6427 GND.n5364 0.152939
R28995 GND.n6428 GND.n6427 0.152939
R28996 GND.n6429 GND.n6428 0.152939
R28997 GND.n6429 GND.n5349 0.152939
R28998 GND.n6482 GND.n5349 0.152939
R28999 GND.n6483 GND.n6482 0.152939
R29000 GND.n6484 GND.n6483 0.152939
R29001 GND.n6484 GND.n5344 0.152939
R29002 GND.n6496 GND.n5344 0.152939
R29003 GND.n6497 GND.n6496 0.152939
R29004 GND.n6498 GND.n6497 0.152939
R29005 GND.n6498 GND.n5339 0.152939
R29006 GND.n6510 GND.n5339 0.152939
R29007 GND.n6511 GND.n6510 0.152939
R29008 GND.n6513 GND.n6511 0.152939
R29009 GND.n6513 GND.n6512 0.152939
R29010 GND.n6512 GND.n5332 0.152939
R29011 GND.n5333 GND.n5332 0.152939
R29012 GND.n5334 GND.n5333 0.152939
R29013 GND.n6524 GND.n5334 0.152939
R29014 GND.n6525 GND.n6524 0.152939
R29015 GND.n6526 GND.n6525 0.152939
R29016 GND.n6527 GND.n6526 0.152939
R29017 GND.n6531 GND.n6527 0.152939
R29018 GND.n6532 GND.n6531 0.152939
R29019 GND.n6533 GND.n6532 0.152939
R29020 GND.n6534 GND.n6533 0.152939
R29021 GND.n6538 GND.n6534 0.152939
R29022 GND.n6539 GND.n6538 0.152939
R29023 GND.n6540 GND.n6539 0.152939
R29024 GND.n6541 GND.n6540 0.152939
R29025 GND.n6545 GND.n6541 0.152939
R29026 GND.n6546 GND.n6545 0.152939
R29027 GND.n6547 GND.n6546 0.152939
R29028 GND.n6548 GND.n6547 0.152939
R29029 GND.n6552 GND.n6548 0.152939
R29030 GND.n6553 GND.n6552 0.152939
R29031 GND.n6554 GND.n6553 0.152939
R29032 GND.n6555 GND.n6554 0.152939
R29033 GND.n6559 GND.n6555 0.152939
R29034 GND.n6560 GND.n6559 0.152939
R29035 GND.n6561 GND.n6560 0.152939
R29036 GND.n6562 GND.n6561 0.152939
R29037 GND.n6566 GND.n6562 0.152939
R29038 GND.n6567 GND.n6566 0.152939
R29039 GND.n6568 GND.n6567 0.152939
R29040 GND.n6569 GND.n6568 0.152939
R29041 GND.n6575 GND.n6569 0.152939
R29042 GND.n6576 GND.n6575 0.152939
R29043 GND.n6576 GND.n5289 0.152939
R29044 GND.n6757 GND.n5289 0.152939
R29045 GND.n6758 GND.n6757 0.152939
R29046 GND.n6759 GND.n6758 0.152939
R29047 GND.n6760 GND.n6759 0.152939
R29048 GND.n6761 GND.n6760 0.152939
R29049 GND.n6762 GND.n6761 0.152939
R29050 GND.n6762 GND.n102 0.152939
R29051 GND.n10313 GND.n103 0.152939
R29052 GND.n5273 GND.n103 0.152939
R29053 GND.n5274 GND.n5273 0.152939
R29054 GND.n5275 GND.n5274 0.152939
R29055 GND.n5276 GND.n5275 0.152939
R29056 GND.n6798 GND.n5276 0.152939
R29057 GND.n6799 GND.n6798 0.152939
R29058 GND.n6800 GND.n6799 0.152939
R29059 GND.n6801 GND.n6800 0.152939
R29060 GND.n6805 GND.n6801 0.152939
R29061 GND.n6806 GND.n6805 0.152939
R29062 GND.n6807 GND.n6806 0.152939
R29063 GND.n6808 GND.n6807 0.152939
R29064 GND.n6812 GND.n6808 0.152939
R29065 GND.n6813 GND.n6812 0.152939
R29066 GND.n6814 GND.n6813 0.152939
R29067 GND.n6815 GND.n6814 0.152939
R29068 GND.n6819 GND.n6815 0.152939
R29069 GND.n6820 GND.n6819 0.152939
R29070 GND.n6821 GND.n6820 0.152939
R29071 GND.n6822 GND.n6821 0.152939
R29072 GND.n6826 GND.n6822 0.152939
R29073 GND.n6827 GND.n6826 0.152939
R29074 GND.n6828 GND.n6827 0.152939
R29075 GND.n6829 GND.n6828 0.152939
R29076 GND.n6829 GND.n439 0.152939
R29077 GND.n9730 GND.n439 0.152939
R29078 GND.n9731 GND.n9730 0.152939
R29079 GND.n9732 GND.n9731 0.152939
R29080 GND.n9732 GND.n435 0.152939
R29081 GND.n9745 GND.n435 0.152939
R29082 GND.n9746 GND.n9745 0.152939
R29083 GND.n9747 GND.n9746 0.152939
R29084 GND.n9747 GND.n431 0.152939
R29085 GND.n9760 GND.n431 0.152939
R29086 GND.n9761 GND.n9760 0.152939
R29087 GND.n9762 GND.n9761 0.152939
R29088 GND.n9762 GND.n427 0.152939
R29089 GND.n9775 GND.n427 0.152939
R29090 GND.n9776 GND.n9775 0.152939
R29091 GND.n9777 GND.n9776 0.152939
R29092 GND.n9777 GND.n423 0.152939
R29093 GND.n9790 GND.n423 0.152939
R29094 GND.n9791 GND.n9790 0.152939
R29095 GND.n9792 GND.n9791 0.152939
R29096 GND.n9793 GND.n9792 0.152939
R29097 GND.n9794 GND.n9793 0.152939
R29098 GND.n9795 GND.n9794 0.152939
R29099 GND.n9796 GND.n9795 0.152939
R29100 GND.n9797 GND.n9796 0.152939
R29101 GND.n9798 GND.n9797 0.152939
R29102 GND.n9799 GND.n9798 0.152939
R29103 GND.n9800 GND.n9799 0.152939
R29104 GND.n9801 GND.n9800 0.152939
R29105 GND.n9802 GND.n9801 0.152939
R29106 GND.n9803 GND.n9802 0.152939
R29107 GND.n9804 GND.n9803 0.152939
R29108 GND.n9805 GND.n9804 0.152939
R29109 GND.n9806 GND.n9805 0.152939
R29110 GND.n10079 GND.n9806 0.152939
R29111 GND.n10051 GND.n10050 0.152939
R29112 GND.n10051 GND.n10048 0.152939
R29113 GND.n10059 GND.n10048 0.152939
R29114 GND.n10060 GND.n10059 0.152939
R29115 GND.n10061 GND.n10060 0.152939
R29116 GND.n10061 GND.n10046 0.152939
R29117 GND.n10068 GND.n10046 0.152939
R29118 GND.n10069 GND.n10068 0.152939
R29119 GND.n10070 GND.n10069 0.152939
R29120 GND.n10070 GND.n9807 0.152939
R29121 GND.n10078 GND.n9807 0.152939
R29122 GND.n9886 GND.n9885 0.152939
R29123 GND.n9886 GND.n9883 0.152939
R29124 GND.n9894 GND.n9883 0.152939
R29125 GND.n9895 GND.n9894 0.152939
R29126 GND.n9896 GND.n9895 0.152939
R29127 GND.n9896 GND.n9881 0.152939
R29128 GND.n9904 GND.n9881 0.152939
R29129 GND.n9905 GND.n9904 0.152939
R29130 GND.n9906 GND.n9905 0.152939
R29131 GND.n9906 GND.n9876 0.152939
R29132 GND.n9913 GND.n9876 0.152939
R29133 GND.n9914 GND.n9913 0.152939
R29134 GND.n9915 GND.n9914 0.152939
R29135 GND.n9915 GND.n9874 0.152939
R29136 GND.n9923 GND.n9874 0.152939
R29137 GND.n9924 GND.n9923 0.152939
R29138 GND.n9925 GND.n9924 0.152939
R29139 GND.n9925 GND.n9872 0.152939
R29140 GND.n9933 GND.n9872 0.152939
R29141 GND.n9934 GND.n9933 0.152939
R29142 GND.n9935 GND.n9934 0.152939
R29143 GND.n9935 GND.n9868 0.152939
R29144 GND.n9944 GND.n9868 0.152939
R29145 GND.n9945 GND.n9944 0.152939
R29146 GND.n9946 GND.n9945 0.152939
R29147 GND.n9946 GND.n9866 0.152939
R29148 GND.n9954 GND.n9866 0.152939
R29149 GND.n9955 GND.n9954 0.152939
R29150 GND.n9956 GND.n9955 0.152939
R29151 GND.n9956 GND.n9864 0.152939
R29152 GND.n9964 GND.n9864 0.152939
R29153 GND.n9965 GND.n9964 0.152939
R29154 GND.n9966 GND.n9965 0.152939
R29155 GND.n9966 GND.n9858 0.152939
R29156 GND.n9972 GND.n9858 0.152939
R29157 GND.n9973 GND.n9972 0.152939
R29158 GND.n9974 GND.n9973 0.152939
R29159 GND.n9974 GND.n9856 0.152939
R29160 GND.n9982 GND.n9856 0.152939
R29161 GND.n9983 GND.n9982 0.152939
R29162 GND.n9984 GND.n9983 0.152939
R29163 GND.n9984 GND.n9854 0.152939
R29164 GND.n9992 GND.n9854 0.152939
R29165 GND.n9993 GND.n9992 0.152939
R29166 GND.n9994 GND.n9993 0.152939
R29167 GND.n9994 GND.n9852 0.152939
R29168 GND.n10005 GND.n9852 0.152939
R29169 GND.n10006 GND.n10005 0.152939
R29170 GND.n10007 GND.n10006 0.152939
R29171 GND.n10007 GND.n9850 0.152939
R29172 GND.n10015 GND.n9850 0.152939
R29173 GND.n10016 GND.n10015 0.152939
R29174 GND.n10017 GND.n10016 0.152939
R29175 GND.n10017 GND.n9848 0.152939
R29176 GND.n10025 GND.n9848 0.152939
R29177 GND.n10026 GND.n10025 0.152939
R29178 GND.n10027 GND.n10026 0.152939
R29179 GND.n10027 GND.n9846 0.152939
R29180 GND.n10034 GND.n9846 0.152939
R29181 GND.n10035 GND.n10034 0.152939
R29182 GND.n10036 GND.n10035 0.152939
R29183 GND.n7097 GND.n7096 0.152939
R29184 GND.n7098 GND.n7097 0.152939
R29185 GND.n7099 GND.n7098 0.152939
R29186 GND.n7100 GND.n7099 0.152939
R29187 GND.n7101 GND.n7100 0.152939
R29188 GND.n7102 GND.n7101 0.152939
R29189 GND.n7103 GND.n7102 0.152939
R29190 GND.n7104 GND.n7103 0.152939
R29191 GND.n7105 GND.n7104 0.152939
R29192 GND.n7107 GND.n7105 0.152939
R29193 GND.n7110 GND.n7107 0.152939
R29194 GND.n7111 GND.n7110 0.152939
R29195 GND.n7112 GND.n7111 0.152939
R29196 GND.n7113 GND.n7112 0.152939
R29197 GND.n7114 GND.n7113 0.152939
R29198 GND.n7115 GND.n7114 0.152939
R29199 GND.n7116 GND.n7115 0.152939
R29200 GND.n7117 GND.n7116 0.152939
R29201 GND.n7118 GND.n7117 0.152939
R29202 GND.n7119 GND.n7118 0.152939
R29203 GND.n7120 GND.n7119 0.152939
R29204 GND.n7121 GND.n7120 0.152939
R29205 GND.n7125 GND.n7121 0.152939
R29206 GND.n7126 GND.n7125 0.152939
R29207 GND.n7127 GND.n7126 0.152939
R29208 GND.n7129 GND.n7127 0.152939
R29209 GND.n7129 GND.n7128 0.152939
R29210 GND.n5382 GND.n4836 0.152939
R29211 GND.n5383 GND.n5382 0.152939
R29212 GND.n5388 GND.n5383 0.152939
R29213 GND.n5389 GND.n5388 0.152939
R29214 GND.n5390 GND.n5389 0.152939
R29215 GND.n5390 GND.n5378 0.152939
R29216 GND.n5398 GND.n5378 0.152939
R29217 GND.n5399 GND.n5398 0.152939
R29218 GND.n5400 GND.n5399 0.152939
R29219 GND.n5400 GND.n5376 0.152939
R29220 GND.n5408 GND.n5376 0.152939
R29221 GND.n5409 GND.n5408 0.152939
R29222 GND.n5410 GND.n5409 0.152939
R29223 GND.n5410 GND.n5374 0.152939
R29224 GND.n5418 GND.n5374 0.152939
R29225 GND.n5419 GND.n5418 0.152939
R29226 GND.n5420 GND.n5419 0.152939
R29227 GND.n5420 GND.n5372 0.152939
R29228 GND.n5431 GND.n5372 0.152939
R29229 GND.n5432 GND.n5431 0.152939
R29230 GND.n5433 GND.n5432 0.152939
R29231 GND.n5433 GND.n5370 0.152939
R29232 GND.n5441 GND.n5370 0.152939
R29233 GND.n5442 GND.n5441 0.152939
R29234 GND.n5443 GND.n5442 0.152939
R29235 GND.n5443 GND.n5368 0.152939
R29236 GND.n5451 GND.n5368 0.152939
R29237 GND.n5452 GND.n5451 0.152939
R29238 GND.n5453 GND.n5452 0.152939
R29239 GND.n5453 GND.n5366 0.152939
R29240 GND.n5462 GND.n5366 0.152939
R29241 GND.n7095 GND.n4879 0.152939
R29242 GND.n4914 GND.n4879 0.152939
R29243 GND.n4917 GND.n4914 0.152939
R29244 GND.n4918 GND.n4917 0.152939
R29245 GND.n4919 GND.n4918 0.152939
R29246 GND.n4920 GND.n4919 0.152939
R29247 GND.n4921 GND.n4920 0.152939
R29248 GND.n4940 GND.n4921 0.152939
R29249 GND.n4941 GND.n4940 0.152939
R29250 GND.n4942 GND.n4941 0.152939
R29251 GND.n4943 GND.n4942 0.152939
R29252 GND.n4961 GND.n4943 0.152939
R29253 GND.n4962 GND.n4961 0.152939
R29254 GND.n4963 GND.n4962 0.152939
R29255 GND.n4964 GND.n4963 0.152939
R29256 GND.n4982 GND.n4964 0.152939
R29257 GND.n4983 GND.n4982 0.152939
R29258 GND.n4984 GND.n4983 0.152939
R29259 GND.n4985 GND.n4984 0.152939
R29260 GND.n5002 GND.n4985 0.152939
R29261 GND.n5003 GND.n5002 0.152939
R29262 GND.n5004 GND.n5003 0.152939
R29263 GND.n5005 GND.n5004 0.152939
R29264 GND.n5023 GND.n5005 0.152939
R29265 GND.n5024 GND.n5023 0.152939
R29266 GND.n5025 GND.n5024 0.152939
R29267 GND.n5026 GND.n5025 0.152939
R29268 GND.n5044 GND.n5026 0.152939
R29269 GND.n5045 GND.n5044 0.152939
R29270 GND.n5046 GND.n5045 0.152939
R29271 GND.n5047 GND.n5046 0.152939
R29272 GND.n5065 GND.n5047 0.152939
R29273 GND.n5066 GND.n5065 0.152939
R29274 GND.n5067 GND.n5066 0.152939
R29275 GND.n5068 GND.n5067 0.152939
R29276 GND.n5086 GND.n5068 0.152939
R29277 GND.n5087 GND.n5086 0.152939
R29278 GND.n5088 GND.n5087 0.152939
R29279 GND.n5089 GND.n5088 0.152939
R29280 GND.n5107 GND.n5089 0.152939
R29281 GND.n5108 GND.n5107 0.152939
R29282 GND.n5109 GND.n5108 0.152939
R29283 GND.n5110 GND.n5109 0.152939
R29284 GND.n5128 GND.n5110 0.152939
R29285 GND.n5129 GND.n5128 0.152939
R29286 GND.n5130 GND.n5129 0.152939
R29287 GND.n5131 GND.n5130 0.152939
R29288 GND.n5149 GND.n5131 0.152939
R29289 GND.n5150 GND.n5149 0.152939
R29290 GND.n5151 GND.n5150 0.152939
R29291 GND.n5152 GND.n5151 0.152939
R29292 GND.n5170 GND.n5152 0.152939
R29293 GND.n5171 GND.n5170 0.152939
R29294 GND.n5172 GND.n5171 0.152939
R29295 GND.n5172 GND.n117 0.152939
R29296 GND.n3338 GND.n3337 0.152939
R29297 GND.n3339 GND.n3338 0.152939
R29298 GND.n3340 GND.n3339 0.152939
R29299 GND.n3343 GND.n3340 0.152939
R29300 GND.n3344 GND.n3343 0.152939
R29301 GND.n3345 GND.n3344 0.152939
R29302 GND.n3346 GND.n3345 0.152939
R29303 GND.n3349 GND.n3346 0.152939
R29304 GND.n3350 GND.n3349 0.152939
R29305 GND.n3351 GND.n3350 0.152939
R29306 GND.n3352 GND.n3351 0.152939
R29307 GND.n3355 GND.n3352 0.152939
R29308 GND.n3356 GND.n3355 0.152939
R29309 GND.n3357 GND.n3356 0.152939
R29310 GND.n3358 GND.n3357 0.152939
R29311 GND.n3361 GND.n3358 0.152939
R29312 GND.n3362 GND.n3361 0.152939
R29313 GND.n3363 GND.n3362 0.152939
R29314 GND.n3364 GND.n3363 0.152939
R29315 GND.n3367 GND.n3364 0.152939
R29316 GND.n3368 GND.n3367 0.152939
R29317 GND.n3369 GND.n3368 0.152939
R29318 GND.n3370 GND.n3369 0.152939
R29319 GND.n3373 GND.n3370 0.152939
R29320 GND.n3374 GND.n3373 0.152939
R29321 GND.n3375 GND.n3374 0.152939
R29322 GND.n3376 GND.n3375 0.152939
R29323 GND.n3379 GND.n3376 0.152939
R29324 GND.n3380 GND.n3379 0.152939
R29325 GND.n3381 GND.n3380 0.152939
R29326 GND.n3382 GND.n3381 0.152939
R29327 GND.n3385 GND.n3382 0.152939
R29328 GND.n3386 GND.n3385 0.152939
R29329 GND.n3387 GND.n3386 0.152939
R29330 GND.n3388 GND.n3387 0.152939
R29331 GND.n3391 GND.n3388 0.152939
R29332 GND.n3392 GND.n3391 0.152939
R29333 GND.n3393 GND.n3392 0.152939
R29334 GND.n3394 GND.n3393 0.152939
R29335 GND.n3397 GND.n3394 0.152939
R29336 GND.n3398 GND.n3397 0.152939
R29337 GND.n3399 GND.n3398 0.152939
R29338 GND.n3400 GND.n3399 0.152939
R29339 GND.n3403 GND.n3400 0.152939
R29340 GND.n3404 GND.n3403 0.152939
R29341 GND.n3405 GND.n3404 0.152939
R29342 GND.n3406 GND.n3405 0.152939
R29343 GND.n3409 GND.n3406 0.152939
R29344 GND.n3410 GND.n3409 0.152939
R29345 GND.n3411 GND.n3410 0.152939
R29346 GND.n3412 GND.n3411 0.152939
R29347 GND.n3415 GND.n3412 0.152939
R29348 GND.n3416 GND.n3415 0.152939
R29349 GND.n3417 GND.n3416 0.152939
R29350 GND.n3418 GND.n3417 0.152939
R29351 GND.n3421 GND.n3418 0.152939
R29352 GND.n3422 GND.n3421 0.152939
R29353 GND.n3423 GND.n3422 0.152939
R29354 GND.n3424 GND.n3423 0.152939
R29355 GND.n3427 GND.n3424 0.152939
R29356 GND.n3428 GND.n3427 0.152939
R29357 GND.n3430 GND.n3428 0.152939
R29358 GND.n3430 GND.n3429 0.152939
R29359 GND.n3429 GND.n1942 0.152939
R29360 GND.n1943 GND.n1942 0.152939
R29361 GND.n1944 GND.n1943 0.152939
R29362 GND.n1958 GND.n1944 0.152939
R29363 GND.n1959 GND.n1958 0.152939
R29364 GND.n1960 GND.n1959 0.152939
R29365 GND.n1961 GND.n1960 0.152939
R29366 GND.n1975 GND.n1961 0.152939
R29367 GND.n1976 GND.n1975 0.152939
R29368 GND.n1977 GND.n1976 0.152939
R29369 GND.n1978 GND.n1977 0.152939
R29370 GND.n1993 GND.n1978 0.152939
R29371 GND.n1994 GND.n1993 0.152939
R29372 GND.n1995 GND.n1994 0.152939
R29373 GND.n1996 GND.n1995 0.152939
R29374 GND.n2011 GND.n1996 0.152939
R29375 GND.n2012 GND.n2011 0.152939
R29376 GND.n2013 GND.n2012 0.152939
R29377 GND.n2014 GND.n2013 0.152939
R29378 GND.n2029 GND.n2014 0.152939
R29379 GND.n2030 GND.n2029 0.152939
R29380 GND.n2031 GND.n2030 0.152939
R29381 GND.n2032 GND.n2031 0.152939
R29382 GND.n2047 GND.n2032 0.152939
R29383 GND.n2048 GND.n2047 0.152939
R29384 GND.n2049 GND.n2048 0.152939
R29385 GND.n2050 GND.n2049 0.152939
R29386 GND.n2065 GND.n2050 0.152939
R29387 GND.n2066 GND.n2065 0.152939
R29388 GND.n2067 GND.n2066 0.152939
R29389 GND.n2068 GND.n2067 0.152939
R29390 GND.n2083 GND.n2068 0.152939
R29391 GND.n2084 GND.n2083 0.152939
R29392 GND.n2085 GND.n2084 0.152939
R29393 GND.n2086 GND.n2085 0.152939
R29394 GND.n2101 GND.n2086 0.152939
R29395 GND.n2102 GND.n2101 0.152939
R29396 GND.n2103 GND.n2102 0.152939
R29397 GND.n2104 GND.n2103 0.152939
R29398 GND.n2320 GND.n2104 0.152939
R29399 GND.n2321 GND.n2320 0.152939
R29400 GND.n2322 GND.n2321 0.152939
R29401 GND.n2323 GND.n2322 0.152939
R29402 GND.n2324 GND.n2323 0.152939
R29403 GND.n3888 GND.n2324 0.152939
R29404 GND.n3889 GND.n3888 0.152939
R29405 GND.n3890 GND.n3889 0.152939
R29406 GND.n3891 GND.n3890 0.152939
R29407 GND.n3907 GND.n3891 0.152939
R29408 GND.n3908 GND.n3907 0.152939
R29409 GND.n3909 GND.n3908 0.152939
R29410 GND.n3910 GND.n3909 0.152939
R29411 GND.n3927 GND.n3910 0.152939
R29412 GND.n3928 GND.n3927 0.152939
R29413 GND.n3929 GND.n3928 0.152939
R29414 GND.n3930 GND.n3929 0.152939
R29415 GND.n3957 GND.n3930 0.152939
R29416 GND.n3958 GND.n3957 0.152939
R29417 GND.n3959 GND.n3958 0.152939
R29418 GND.n3960 GND.n3959 0.152939
R29419 GND.n3961 GND.n3960 0.152939
R29420 GND.n3991 GND.n3961 0.152939
R29421 GND.n3992 GND.n3991 0.152939
R29422 GND.n3993 GND.n3992 0.152939
R29423 GND.n3994 GND.n3993 0.152939
R29424 GND.n4011 GND.n3994 0.152939
R29425 GND.n4012 GND.n4011 0.152939
R29426 GND.n4013 GND.n4012 0.152939
R29427 GND.n4014 GND.n4013 0.152939
R29428 GND.n4031 GND.n4014 0.152939
R29429 GND.n4032 GND.n4031 0.152939
R29430 GND.n4033 GND.n4032 0.152939
R29431 GND.n4034 GND.n4033 0.152939
R29432 GND.n4062 GND.n4034 0.152939
R29433 GND.n4063 GND.n4062 0.152939
R29434 GND.n4064 GND.n4063 0.152939
R29435 GND.n4065 GND.n4064 0.152939
R29436 GND.n4066 GND.n4065 0.152939
R29437 GND.n4096 GND.n4066 0.152939
R29438 GND.n4097 GND.n4096 0.152939
R29439 GND.n4098 GND.n4097 0.152939
R29440 GND.n4099 GND.n4098 0.152939
R29441 GND.n4116 GND.n4099 0.152939
R29442 GND.n4117 GND.n4116 0.152939
R29443 GND.n4118 GND.n4117 0.152939
R29444 GND.n4119 GND.n4118 0.152939
R29445 GND.n4136 GND.n4119 0.152939
R29446 GND.n4137 GND.n4136 0.152939
R29447 GND.n4138 GND.n4137 0.152939
R29448 GND.n4139 GND.n4138 0.152939
R29449 GND.n4167 GND.n4139 0.152939
R29450 GND.n4168 GND.n4167 0.152939
R29451 GND.n4169 GND.n4168 0.152939
R29452 GND.n4170 GND.n4169 0.152939
R29453 GND.n4171 GND.n4170 0.152939
R29454 GND.n4200 GND.n4171 0.152939
R29455 GND.n4201 GND.n4200 0.152939
R29456 GND.n4202 GND.n4201 0.152939
R29457 GND.n4203 GND.n4202 0.152939
R29458 GND.n4220 GND.n4203 0.152939
R29459 GND.n4221 GND.n4220 0.152939
R29460 GND.n4222 GND.n4221 0.152939
R29461 GND.n4223 GND.n4222 0.152939
R29462 GND.n4239 GND.n4223 0.152939
R29463 GND.n4240 GND.n4239 0.152939
R29464 GND.n4241 GND.n4240 0.152939
R29465 GND.n4242 GND.n4241 0.152939
R29466 GND.n4270 GND.n4242 0.152939
R29467 GND.n4271 GND.n4270 0.152939
R29468 GND.n4272 GND.n4271 0.152939
R29469 GND.n4273 GND.n4272 0.152939
R29470 GND.n4274 GND.n4273 0.152939
R29471 GND.n4303 GND.n4274 0.152939
R29472 GND.n4304 GND.n4303 0.152939
R29473 GND.n4305 GND.n4304 0.152939
R29474 GND.n4306 GND.n4305 0.152939
R29475 GND.n4323 GND.n4306 0.152939
R29476 GND.n4324 GND.n4323 0.152939
R29477 GND.n4325 GND.n4324 0.152939
R29478 GND.n4326 GND.n4325 0.152939
R29479 GND.n4343 GND.n4326 0.152939
R29480 GND.n4344 GND.n4343 0.152939
R29481 GND.n4345 GND.n4344 0.152939
R29482 GND.n4346 GND.n4345 0.152939
R29483 GND.n4374 GND.n4346 0.152939
R29484 GND.n4375 GND.n4374 0.152939
R29485 GND.n4376 GND.n4375 0.152939
R29486 GND.n4377 GND.n4376 0.152939
R29487 GND.n4378 GND.n4377 0.152939
R29488 GND.n4408 GND.n4378 0.152939
R29489 GND.n4409 GND.n4408 0.152939
R29490 GND.n4410 GND.n4409 0.152939
R29491 GND.n4411 GND.n4410 0.152939
R29492 GND.n4440 GND.n4411 0.152939
R29493 GND.n4441 GND.n4440 0.152939
R29494 GND.n4442 GND.n4441 0.152939
R29495 GND.n4443 GND.n4442 0.152939
R29496 GND.n4444 GND.n4443 0.152939
R29497 GND.n4459 GND.n4444 0.152939
R29498 GND.n4460 GND.n4459 0.152939
R29499 GND.n4461 GND.n4460 0.152939
R29500 GND.n4462 GND.n4461 0.152939
R29501 GND.n4477 GND.n4462 0.152939
R29502 GND.n4478 GND.n4477 0.152939
R29503 GND.n4479 GND.n4478 0.152939
R29504 GND.n4480 GND.n4479 0.152939
R29505 GND.n4495 GND.n4480 0.152939
R29506 GND.n4496 GND.n4495 0.152939
R29507 GND.n4497 GND.n4496 0.152939
R29508 GND.n4498 GND.n4497 0.152939
R29509 GND.n4513 GND.n4498 0.152939
R29510 GND.n4514 GND.n4513 0.152939
R29511 GND.n4515 GND.n4514 0.152939
R29512 GND.n4516 GND.n4515 0.152939
R29513 GND.n4531 GND.n4516 0.152939
R29514 GND.n4532 GND.n4531 0.152939
R29515 GND.n4533 GND.n4532 0.152939
R29516 GND.n4534 GND.n4533 0.152939
R29517 GND.n4562 GND.n4534 0.152939
R29518 GND.n4563 GND.n4562 0.152939
R29519 GND.n4564 GND.n4563 0.152939
R29520 GND.n4565 GND.n4564 0.152939
R29521 GND.n4566 GND.n4565 0.152939
R29522 GND.n4581 GND.n4566 0.152939
R29523 GND.n4582 GND.n4581 0.152939
R29524 GND.n4583 GND.n4582 0.152939
R29525 GND.n4584 GND.n4583 0.152939
R29526 GND.n4599 GND.n4584 0.152939
R29527 GND.n4600 GND.n4599 0.152939
R29528 GND.n4601 GND.n4600 0.152939
R29529 GND.n4602 GND.n4601 0.152939
R29530 GND.n4616 GND.n4602 0.152939
R29531 GND.n4617 GND.n4616 0.152939
R29532 GND.n4618 GND.n4617 0.152939
R29533 GND.n4619 GND.n4618 0.152939
R29534 GND.n4693 GND.n4619 0.152939
R29535 GND.n4694 GND.n4693 0.152939
R29536 GND.n4695 GND.n4694 0.152939
R29537 GND.n4696 GND.n4695 0.152939
R29538 GND.n4697 GND.n4696 0.152939
R29539 GND.n6394 GND.n4697 0.152939
R29540 GND.n6395 GND.n6394 0.152939
R29541 GND.n6396 GND.n6395 0.152939
R29542 GND.n6396 GND.n6391 0.152939
R29543 GND.n6406 GND.n6391 0.152939
R29544 GND.n6407 GND.n6406 0.152939
R29545 GND.n6408 GND.n6407 0.152939
R29546 GND.n6410 GND.n6408 0.152939
R29547 GND.n6410 GND.n6409 0.152939
R29548 GND.n6409 GND.n4900 0.152939
R29549 GND.n4901 GND.n4900 0.152939
R29550 GND.n4902 GND.n4901 0.152939
R29551 GND.n6433 GND.n4902 0.152939
R29552 GND.n6434 GND.n6433 0.152939
R29553 GND.n6435 GND.n6434 0.152939
R29554 GND.n6436 GND.n6435 0.152939
R29555 GND.n6439 GND.n6436 0.152939
R29556 GND.n6440 GND.n6439 0.152939
R29557 GND.n6441 GND.n6440 0.152939
R29558 GND.n6442 GND.n6441 0.152939
R29559 GND.n6445 GND.n6442 0.152939
R29560 GND.n6446 GND.n6445 0.152939
R29561 GND.n6447 GND.n6446 0.152939
R29562 GND.n6448 GND.n6447 0.152939
R29563 GND.n6450 GND.n6448 0.152939
R29564 GND.n6451 GND.n6450 0.152939
R29565 GND.n6451 GND.n5327 0.152939
R29566 GND.n6679 GND.n5327 0.152939
R29567 GND.n6680 GND.n6679 0.152939
R29568 GND.n6681 GND.n6680 0.152939
R29569 GND.n6681 GND.n5323 0.152939
R29570 GND.n6687 GND.n5323 0.152939
R29571 GND.n6688 GND.n6687 0.152939
R29572 GND.n6689 GND.n6688 0.152939
R29573 GND.n6689 GND.n5319 0.152939
R29574 GND.n6695 GND.n5319 0.152939
R29575 GND.n6696 GND.n6695 0.152939
R29576 GND.n6697 GND.n6696 0.152939
R29577 GND.n6697 GND.n5315 0.152939
R29578 GND.n6703 GND.n5315 0.152939
R29579 GND.n6704 GND.n6703 0.152939
R29580 GND.n6705 GND.n6704 0.152939
R29581 GND.n6705 GND.n5311 0.152939
R29582 GND.n6711 GND.n5311 0.152939
R29583 GND.n6712 GND.n6711 0.152939
R29584 GND.n6713 GND.n6712 0.152939
R29585 GND.n6713 GND.n5307 0.152939
R29586 GND.n6719 GND.n5307 0.152939
R29587 GND.n6720 GND.n6719 0.152939
R29588 GND.n6721 GND.n6720 0.152939
R29589 GND.n6721 GND.n5303 0.152939
R29590 GND.n6727 GND.n5303 0.152939
R29591 GND.n6728 GND.n6727 0.152939
R29592 GND.n6729 GND.n6728 0.152939
R29593 GND.n6729 GND.n5299 0.152939
R29594 GND.n6735 GND.n5299 0.152939
R29595 GND.n6736 GND.n6735 0.152939
R29596 GND.n6737 GND.n6736 0.152939
R29597 GND.n6737 GND.n5295 0.152939
R29598 GND.n6743 GND.n5295 0.152939
R29599 GND.n6744 GND.n6743 0.152939
R29600 GND.n6745 GND.n6744 0.152939
R29601 GND.n6746 GND.n6745 0.152939
R29602 GND.n2580 GND.n1541 0.152939
R29603 GND.n3578 GND.n2580 0.152939
R29604 GND.n3579 GND.n3578 0.152939
R29605 GND.n3580 GND.n3579 0.152939
R29606 GND.n3581 GND.n3580 0.152939
R29607 GND.n3581 GND.n2558 0.152939
R29608 GND.n3604 GND.n2558 0.152939
R29609 GND.n3605 GND.n3604 0.152939
R29610 GND.n3606 GND.n3605 0.152939
R29611 GND.n3607 GND.n3606 0.152939
R29612 GND.n3607 GND.n2537 0.152939
R29613 GND.n3630 GND.n2537 0.152939
R29614 GND.n3631 GND.n3630 0.152939
R29615 GND.n3632 GND.n3631 0.152939
R29616 GND.n3633 GND.n3632 0.152939
R29617 GND.n3633 GND.n2515 0.152939
R29618 GND.n3656 GND.n2515 0.152939
R29619 GND.n3657 GND.n3656 0.152939
R29620 GND.n3658 GND.n3657 0.152939
R29621 GND.n3659 GND.n3658 0.152939
R29622 GND.n3659 GND.n2493 0.152939
R29623 GND.n3681 GND.n2493 0.152939
R29624 GND.n3682 GND.n3681 0.152939
R29625 GND.n3683 GND.n3682 0.152939
R29626 GND.n3684 GND.n3683 0.152939
R29627 GND.n3684 GND.n2471 0.152939
R29628 GND.n3707 GND.n2471 0.152939
R29629 GND.n3708 GND.n3707 0.152939
R29630 GND.n3709 GND.n3708 0.152939
R29631 GND.n3710 GND.n3709 0.152939
R29632 GND.n3710 GND.n2450 0.152939
R29633 GND.n3733 GND.n2450 0.152939
R29634 GND.n3734 GND.n3733 0.152939
R29635 GND.n3735 GND.n3734 0.152939
R29636 GND.n3736 GND.n3735 0.152939
R29637 GND.n3736 GND.n2430 0.152939
R29638 GND.n3759 GND.n2430 0.152939
R29639 GND.n3760 GND.n3759 0.152939
R29640 GND.n3761 GND.n3760 0.152939
R29641 GND.n3762 GND.n3761 0.152939
R29642 GND.n3762 GND.n2408 0.152939
R29643 GND.n3784 GND.n2408 0.152939
R29644 GND.n3785 GND.n3784 0.152939
R29645 GND.n3786 GND.n3785 0.152939
R29646 GND.n3787 GND.n3786 0.152939
R29647 GND.n3787 GND.n2386 0.152939
R29648 GND.n3810 GND.n2386 0.152939
R29649 GND.n3811 GND.n3810 0.152939
R29650 GND.n3812 GND.n3811 0.152939
R29651 GND.n3813 GND.n3812 0.152939
R29652 GND.n3813 GND.n2365 0.152939
R29653 GND.n3837 GND.n2365 0.152939
R29654 GND.n3838 GND.n3837 0.152939
R29655 GND.n3839 GND.n3838 0.152939
R29656 GND.n3839 GND.n1724 0.152939
R29657 GND.n1364 GND.n1363 0.152939
R29658 GND.n1365 GND.n1364 0.152939
R29659 GND.n1366 GND.n1365 0.152939
R29660 GND.n1367 GND.n1366 0.152939
R29661 GND.n1368 GND.n1367 0.152939
R29662 GND.n1369 GND.n1368 0.152939
R29663 GND.n1370 GND.n1369 0.152939
R29664 GND.n1371 GND.n1370 0.152939
R29665 GND.n1372 GND.n1371 0.152939
R29666 GND.n1374 GND.n1372 0.152939
R29667 GND.n1377 GND.n1374 0.152939
R29668 GND.n1378 GND.n1377 0.152939
R29669 GND.n1379 GND.n1378 0.152939
R29670 GND.n1380 GND.n1379 0.152939
R29671 GND.n1381 GND.n1380 0.152939
R29672 GND.n1382 GND.n1381 0.152939
R29673 GND.n1383 GND.n1382 0.152939
R29674 GND.n1384 GND.n1383 0.152939
R29675 GND.n1385 GND.n1384 0.152939
R29676 GND.n1386 GND.n1385 0.152939
R29677 GND.n1387 GND.n1386 0.152939
R29678 GND.n1388 GND.n1387 0.152939
R29679 GND.n1392 GND.n1388 0.152939
R29680 GND.n1393 GND.n1392 0.152939
R29681 GND.n1394 GND.n1393 0.152939
R29682 GND.n1395 GND.n1394 0.152939
R29683 GND.n1396 GND.n1395 0.152939
R29684 GND.n1397 GND.n1396 0.152939
R29685 GND.n1398 GND.n1397 0.152939
R29686 GND.n1399 GND.n1398 0.152939
R29687 GND.n1400 GND.n1399 0.152939
R29688 GND.n1401 GND.n1400 0.152939
R29689 GND.n1402 GND.n1401 0.152939
R29690 GND.n1403 GND.n1402 0.152939
R29691 GND.n1404 GND.n1403 0.152939
R29692 GND.n1407 GND.n1404 0.152939
R29693 GND.n1408 GND.n1407 0.152939
R29694 GND.n1409 GND.n1408 0.152939
R29695 GND.n1410 GND.n1409 0.152939
R29696 GND.n1411 GND.n1410 0.152939
R29697 GND.n1412 GND.n1411 0.152939
R29698 GND.n1413 GND.n1412 0.152939
R29699 GND.n1414 GND.n1413 0.152939
R29700 GND.n1415 GND.n1414 0.152939
R29701 GND.n1416 GND.n1415 0.152939
R29702 GND.n1417 GND.n1416 0.152939
R29703 GND.n1418 GND.n1417 0.152939
R29704 GND.n1421 GND.n1418 0.152939
R29705 GND.n1422 GND.n1421 0.152939
R29706 GND.n1423 GND.n1422 0.152939
R29707 GND.n1424 GND.n1423 0.152939
R29708 GND.n1425 GND.n1424 0.152939
R29709 GND.n1426 GND.n1425 0.152939
R29710 GND.n1427 GND.n1426 0.152939
R29711 GND.n1428 GND.n1427 0.152939
R29712 GND.n1429 GND.n1428 0.152939
R29713 GND.n1430 GND.n1429 0.152939
R29714 GND.n1431 GND.n1430 0.152939
R29715 GND.n1432 GND.n1431 0.152939
R29716 GND.n8241 GND.n1432 0.152939
R29717 GND.n8241 GND.n8240 0.152939
R29718 GND.n2940 GND.n2939 0.152939
R29719 GND.n2941 GND.n2940 0.152939
R29720 GND.n2941 GND.n2908 0.152939
R29721 GND.n2956 GND.n2908 0.152939
R29722 GND.n2957 GND.n2956 0.152939
R29723 GND.n2958 GND.n2957 0.152939
R29724 GND.n2958 GND.n2888 0.152939
R29725 GND.n2973 GND.n2888 0.152939
R29726 GND.n2974 GND.n2973 0.152939
R29727 GND.n2975 GND.n2974 0.152939
R29728 GND.n2975 GND.n2869 0.152939
R29729 GND.n2997 GND.n2869 0.152939
R29730 GND.n2998 GND.n2997 0.152939
R29731 GND.n2999 GND.n2998 0.152939
R29732 GND.n3000 GND.n2999 0.152939
R29733 GND.n3000 GND.n2845 0.152939
R29734 GND.n3030 GND.n2845 0.152939
R29735 GND.n3031 GND.n3030 0.152939
R29736 GND.n3032 GND.n3031 0.152939
R29737 GND.n3032 GND.n2821 0.152939
R29738 GND.n3063 GND.n2821 0.152939
R29739 GND.n3064 GND.n3063 0.152939
R29740 GND.n3065 GND.n3064 0.152939
R29741 GND.n3066 GND.n3065 0.152939
R29742 GND.n3066 GND.n2792 0.152939
R29743 GND.n3100 GND.n2792 0.152939
R29744 GND.n3101 GND.n3100 0.152939
R29745 GND.n3102 GND.n3101 0.152939
R29746 GND.n3103 GND.n3102 0.152939
R29747 GND.n3103 GND.n2762 0.152939
R29748 GND.n3138 GND.n2762 0.152939
R29749 GND.n3139 GND.n3138 0.152939
R29750 GND.n3140 GND.n3139 0.152939
R29751 GND.n3141 GND.n3140 0.152939
R29752 GND.n3141 GND.n2735 0.152939
R29753 GND.n3176 GND.n2735 0.152939
R29754 GND.n3177 GND.n3176 0.152939
R29755 GND.n3178 GND.n3177 0.152939
R29756 GND.n3179 GND.n3178 0.152939
R29757 GND.n3179 GND.n2706 0.152939
R29758 GND.n3213 GND.n2706 0.152939
R29759 GND.n3214 GND.n3213 0.152939
R29760 GND.n3215 GND.n3214 0.152939
R29761 GND.n3216 GND.n3215 0.152939
R29762 GND.n3216 GND.n2677 0.152939
R29763 GND.n3250 GND.n2677 0.152939
R29764 GND.n3251 GND.n3250 0.152939
R29765 GND.n3252 GND.n3251 0.152939
R29766 GND.n3253 GND.n3252 0.152939
R29767 GND.n3253 GND.n2647 0.152939
R29768 GND.n3287 GND.n2647 0.152939
R29769 GND.n3288 GND.n3287 0.152939
R29770 GND.n3289 GND.n3288 0.152939
R29771 GND.n3290 GND.n3289 0.152939
R29772 GND.n3290 GND.n1542 0.152939
R29773 GND.n3011 GND.n3010 0.152939
R29774 GND.n3012 GND.n3011 0.152939
R29775 GND.n3013 GND.n3012 0.152939
R29776 GND.n3013 GND.n2837 0.152939
R29777 GND.n3039 GND.n2837 0.152939
R29778 GND.n3040 GND.n3039 0.152939
R29779 GND.n3041 GND.n3040 0.152939
R29780 GND.n3041 GND.n2810 0.152939
R29781 GND.n3074 GND.n2810 0.152939
R29782 GND.n3075 GND.n3074 0.152939
R29783 GND.n3076 GND.n3075 0.152939
R29784 GND.n3077 GND.n3076 0.152939
R29785 GND.n3077 GND.n2781 0.152939
R29786 GND.n3111 GND.n2781 0.152939
R29787 GND.n3112 GND.n3111 0.152939
R29788 GND.n3113 GND.n3112 0.152939
R29789 GND.n3114 GND.n3113 0.152939
R29790 GND.n3114 GND.n2753 0.152939
R29791 GND.n3149 GND.n2753 0.152939
R29792 GND.n3150 GND.n3149 0.152939
R29793 GND.n3151 GND.n3150 0.152939
R29794 GND.n3152 GND.n3151 0.152939
R29795 GND.n3152 GND.n2725 0.152939
R29796 GND.n3187 GND.n2725 0.152939
R29797 GND.n3188 GND.n3187 0.152939
R29798 GND.n3189 GND.n3188 0.152939
R29799 GND.n3190 GND.n3189 0.152939
R29800 GND.n3190 GND.n2695 0.152939
R29801 GND.n3224 GND.n2695 0.152939
R29802 GND.n3225 GND.n3224 0.152939
R29803 GND.n3226 GND.n3225 0.152939
R29804 GND.n3227 GND.n3226 0.152939
R29805 GND.n3227 GND.n2666 0.152939
R29806 GND.n3261 GND.n2666 0.152939
R29807 GND.n3262 GND.n3261 0.152939
R29808 GND.n3263 GND.n3262 0.152939
R29809 GND.n3264 GND.n3263 0.152939
R29810 GND.n3264 GND.n2637 0.152939
R29811 GND.n3299 GND.n2637 0.152939
R29812 GND.n3300 GND.n3299 0.152939
R29813 GND.n3301 GND.n3300 0.152939
R29814 GND.n1191 GND.n1190 0.152939
R29815 GND.n1192 GND.n1191 0.152939
R29816 GND.n1197 GND.n1192 0.152939
R29817 GND.n1198 GND.n1197 0.152939
R29818 GND.n1199 GND.n1198 0.152939
R29819 GND.n1200 GND.n1199 0.152939
R29820 GND.n1205 GND.n1200 0.152939
R29821 GND.n1206 GND.n1205 0.152939
R29822 GND.n1207 GND.n1206 0.152939
R29823 GND.n1208 GND.n1207 0.152939
R29824 GND.n1213 GND.n1208 0.152939
R29825 GND.n1214 GND.n1213 0.152939
R29826 GND.n1215 GND.n1214 0.152939
R29827 GND.n1216 GND.n1215 0.152939
R29828 GND.n1221 GND.n1216 0.152939
R29829 GND.n1222 GND.n1221 0.152939
R29830 GND.n1223 GND.n1222 0.152939
R29831 GND.n1224 GND.n1223 0.152939
R29832 GND.n1229 GND.n1224 0.152939
R29833 GND.n1230 GND.n1229 0.152939
R29834 GND.n1231 GND.n1230 0.152939
R29835 GND.n1232 GND.n1231 0.152939
R29836 GND.n1237 GND.n1232 0.152939
R29837 GND.n1238 GND.n1237 0.152939
R29838 GND.n1239 GND.n1238 0.152939
R29839 GND.n1240 GND.n1239 0.152939
R29840 GND.n1245 GND.n1240 0.152939
R29841 GND.n1246 GND.n1245 0.152939
R29842 GND.n1247 GND.n1246 0.152939
R29843 GND.n1248 GND.n1247 0.152939
R29844 GND.n1253 GND.n1248 0.152939
R29845 GND.n1254 GND.n1253 0.152939
R29846 GND.n1255 GND.n1254 0.152939
R29847 GND.n1256 GND.n1255 0.152939
R29848 GND.n1261 GND.n1256 0.152939
R29849 GND.n1262 GND.n1261 0.152939
R29850 GND.n1263 GND.n1262 0.152939
R29851 GND.n1264 GND.n1263 0.152939
R29852 GND.n1269 GND.n1264 0.152939
R29853 GND.n1270 GND.n1269 0.152939
R29854 GND.n1271 GND.n1270 0.152939
R29855 GND.n1272 GND.n1271 0.152939
R29856 GND.n1277 GND.n1272 0.152939
R29857 GND.n1278 GND.n1277 0.152939
R29858 GND.n1279 GND.n1278 0.152939
R29859 GND.n1280 GND.n1279 0.152939
R29860 GND.n1285 GND.n1280 0.152939
R29861 GND.n1286 GND.n1285 0.152939
R29862 GND.n1287 GND.n1286 0.152939
R29863 GND.n1288 GND.n1287 0.152939
R29864 GND.n1293 GND.n1288 0.152939
R29865 GND.n1294 GND.n1293 0.152939
R29866 GND.n1295 GND.n1294 0.152939
R29867 GND.n1296 GND.n1295 0.152939
R29868 GND.n1301 GND.n1296 0.152939
R29869 GND.n1302 GND.n1301 0.152939
R29870 GND.n1303 GND.n1302 0.152939
R29871 GND.n1304 GND.n1303 0.152939
R29872 GND.n1309 GND.n1304 0.152939
R29873 GND.n1310 GND.n1309 0.152939
R29874 GND.n1311 GND.n1310 0.152939
R29875 GND.n1312 GND.n1311 0.152939
R29876 GND.n1317 GND.n1312 0.152939
R29877 GND.n1318 GND.n1317 0.152939
R29878 GND.n1319 GND.n1318 0.152939
R29879 GND.n1320 GND.n1319 0.152939
R29880 GND.n8020 GND.n8019 0.152939
R29881 GND.n8019 GND.n8018 0.152939
R29882 GND.n8018 GND.n1725 0.152939
R29883 GND.n8014 GND.n1725 0.152939
R29884 GND.n8014 GND.n8013 0.152939
R29885 GND.n8013 GND.n8012 0.152939
R29886 GND.n8012 GND.n1731 0.152939
R29887 GND.n8008 GND.n1731 0.152939
R29888 GND.n8008 GND.n8007 0.152939
R29889 GND.n8007 GND.n8006 0.152939
R29890 GND.n8006 GND.n1737 0.152939
R29891 GND.n8002 GND.n1737 0.152939
R29892 GND.n8002 GND.n8001 0.152939
R29893 GND.n8001 GND.n8000 0.152939
R29894 GND.n8000 GND.n1745 0.152939
R29895 GND.n7996 GND.n1745 0.152939
R29896 GND.n7996 GND.n7995 0.152939
R29897 GND.n7995 GND.n7994 0.152939
R29898 GND.n7994 GND.n1751 0.152939
R29899 GND.n7990 GND.n1751 0.152939
R29900 GND.n7990 GND.n7989 0.152939
R29901 GND.n7989 GND.n7988 0.152939
R29902 GND.n7988 GND.n1757 0.152939
R29903 GND.n7983 GND.n1757 0.152939
R29904 GND.n7983 GND.n7982 0.152939
R29905 GND.n7982 GND.n7981 0.152939
R29906 GND.n7981 GND.n1765 0.152939
R29907 GND.n1868 GND.n1867 0.152939
R29908 GND.n1867 GND.n1769 0.152939
R29909 GND.n1863 GND.n1769 0.152939
R29910 GND.n1863 GND.n1862 0.152939
R29911 GND.n1862 GND.n1861 0.152939
R29912 GND.n1861 GND.n1775 0.152939
R29913 GND.n1857 GND.n1775 0.152939
R29914 GND.n1857 GND.n1856 0.152939
R29915 GND.n1856 GND.n1855 0.152939
R29916 GND.n1855 GND.n1783 0.152939
R29917 GND.n1851 GND.n1783 0.152939
R29918 GND.n1851 GND.n1850 0.152939
R29919 GND.n1850 GND.n1849 0.152939
R29920 GND.n1849 GND.n1789 0.152939
R29921 GND.n1845 GND.n1789 0.152939
R29922 GND.n1845 GND.n1844 0.152939
R29923 GND.n1844 GND.n1843 0.152939
R29924 GND.n1843 GND.n1795 0.152939
R29925 GND.n1838 GND.n1795 0.152939
R29926 GND.n1838 GND.n1837 0.152939
R29927 GND.n1837 GND.n1836 0.152939
R29928 GND.n1836 GND.n1803 0.152939
R29929 GND.n1832 GND.n1803 0.152939
R29930 GND.n1832 GND.n1831 0.152939
R29931 GND.n1831 GND.n1830 0.152939
R29932 GND.n1830 GND.n1809 0.152939
R29933 GND.n1826 GND.n1809 0.152939
R29934 GND.n1826 GND.n1825 0.152939
R29935 GND.n1825 GND.n1824 0.152939
R29936 GND.n1824 GND.n1815 0.152939
R29937 GND.n1820 GND.n1815 0.152939
R29938 GND.n8238 GND.n1438 0.152939
R29939 GND.n8234 GND.n1438 0.152939
R29940 GND.n8234 GND.n8233 0.152939
R29941 GND.n8233 GND.n8232 0.152939
R29942 GND.n8232 GND.n1443 0.152939
R29943 GND.n8228 GND.n1443 0.152939
R29944 GND.n8228 GND.n8227 0.152939
R29945 GND.n8227 GND.n8226 0.152939
R29946 GND.n8226 GND.n1449 0.152939
R29947 GND.n8219 GND.n1449 0.152939
R29948 GND.n8219 GND.n8218 0.152939
R29949 GND.n8217 GND.n1453 0.152939
R29950 GND.n8213 GND.n1453 0.152939
R29951 GND.n8213 GND.n8212 0.152939
R29952 GND.n8212 GND.n8211 0.152939
R29953 GND.n8211 GND.n1458 0.152939
R29954 GND.n8207 GND.n1458 0.152939
R29955 GND.n8207 GND.n8206 0.152939
R29956 GND.n8206 GND.n8205 0.152939
R29957 GND.n8205 GND.n1463 0.152939
R29958 GND.n8201 GND.n1463 0.152939
R29959 GND.n8201 GND.n8200 0.152939
R29960 GND.n8200 GND.n8199 0.152939
R29961 GND.n8199 GND.n1468 0.152939
R29962 GND.n8195 GND.n1468 0.152939
R29963 GND.n8195 GND.n8194 0.152939
R29964 GND.n8194 GND.n8193 0.152939
R29965 GND.n8193 GND.n1473 0.152939
R29966 GND.n8189 GND.n1473 0.152939
R29967 GND.n8189 GND.n8188 0.152939
R29968 GND.n8188 GND.n8187 0.152939
R29969 GND.n8187 GND.n1478 0.152939
R29970 GND.n8183 GND.n1478 0.152939
R29971 GND.n8183 GND.n8182 0.152939
R29972 GND.n8182 GND.n8181 0.152939
R29973 GND.n8181 GND.n1483 0.152939
R29974 GND.n8177 GND.n1483 0.152939
R29975 GND.n8177 GND.n8176 0.152939
R29976 GND.n8176 GND.n8175 0.152939
R29977 GND.n8175 GND.n1488 0.152939
R29978 GND.n8171 GND.n1488 0.152939
R29979 GND.n8171 GND.n8170 0.152939
R29980 GND.n8170 GND.n8169 0.152939
R29981 GND.n8169 GND.n1493 0.152939
R29982 GND.n8165 GND.n1493 0.152939
R29983 GND.n8165 GND.n8164 0.152939
R29984 GND.n8164 GND.n8163 0.152939
R29985 GND.n8163 GND.n1498 0.152939
R29986 GND.n8159 GND.n1498 0.152939
R29987 GND.n8159 GND.n8158 0.152939
R29988 GND.n8158 GND.n8157 0.152939
R29989 GND.n8157 GND.n1503 0.152939
R29990 GND.n8153 GND.n1503 0.152939
R29991 GND.n8153 GND.n8152 0.152939
R29992 GND.n8152 GND.n8151 0.152939
R29993 GND.n8151 GND.n1508 0.152939
R29994 GND.n8147 GND.n1508 0.152939
R29995 GND.n8147 GND.n8146 0.152939
R29996 GND.n8146 GND.n8145 0.152939
R29997 GND.n8145 GND.n1513 0.152939
R29998 GND.n8141 GND.n1513 0.152939
R29999 GND.n8141 GND.n8140 0.152939
R30000 GND.n8140 GND.n8139 0.152939
R30001 GND.n8139 GND.n1518 0.152939
R30002 GND.n8135 GND.n1518 0.152939
R30003 GND.n8135 GND.n8134 0.152939
R30004 GND.n8134 GND.n8133 0.152939
R30005 GND.n8133 GND.n1523 0.152939
R30006 GND.n8129 GND.n1523 0.152939
R30007 GND.n8129 GND.n8128 0.152939
R30008 GND.n8128 GND.n8127 0.152939
R30009 GND.n5201 GND.n118 0.134646
R30010 GND.n3301 GND.n1543 0.134646
R30011 GND.n10306 GND.n116 0.0767195
R30012 GND.n10306 GND.n117 0.0767195
R30013 GND.n8119 GND.n1541 0.0767195
R30014 GND.n8119 GND.n1542 0.0767195
R30015 GND.n1530 GND.n1528 0.0695946
R30016 GND.n10314 GND.n102 0.0695946
R30017 GND.n10314 GND.n10313 0.0695946
R30018 GND.n8127 GND.n1528 0.0695946
R30019 GND.n6357 GND.n5463 0.063
R30020 GND.n3874 GND.n1673 0.063
R30021 GND.n5463 GND.n4890 0.0460163
R30022 GND.n10132 GND.n420 0.0460163
R30023 GND.n8239 GND.n1437 0.0460163
R30024 GND.n8029 GND.n1673 0.0460163
R30025 GND.n7088 GND.n4890 0.0344674
R30026 GND.n7088 GND.n4891 0.0344674
R30027 GND.n5355 GND.n4891 0.0344674
R30028 GND.n5355 GND.n5354 0.0344674
R30029 GND.n5361 GND.n5354 0.0344674
R30030 GND.n5362 GND.n5361 0.0344674
R30031 GND.n5362 GND.n4930 0.0344674
R30032 GND.n4931 GND.n4930 0.0344674
R30033 GND.n4932 GND.n4931 0.0344674
R30034 GND.n5347 GND.n4932 0.0344674
R30035 GND.n5347 GND.n4951 0.0344674
R30036 GND.n4952 GND.n4951 0.0344674
R30037 GND.n4953 GND.n4952 0.0344674
R30038 GND.n5342 GND.n4953 0.0344674
R30039 GND.n5342 GND.n4972 0.0344674
R30040 GND.n4973 GND.n4972 0.0344674
R30041 GND.n4974 GND.n4973 0.0344674
R30042 GND.n5337 GND.n4974 0.0344674
R30043 GND.n5337 GND.n4993 0.0344674
R30044 GND.n4994 GND.n4993 0.0344674
R30045 GND.n4995 GND.n4994 0.0344674
R30046 GND.n6522 GND.n4995 0.0344674
R30047 GND.n6522 GND.n5013 0.0344674
R30048 GND.n5014 GND.n5013 0.0344674
R30049 GND.n5015 GND.n5014 0.0344674
R30050 GND.n6529 GND.n5015 0.0344674
R30051 GND.n6529 GND.n5034 0.0344674
R30052 GND.n5035 GND.n5034 0.0344674
R30053 GND.n5036 GND.n5035 0.0344674
R30054 GND.n6536 GND.n5036 0.0344674
R30055 GND.n6536 GND.n5055 0.0344674
R30056 GND.n5056 GND.n5055 0.0344674
R30057 GND.n5057 GND.n5056 0.0344674
R30058 GND.n6543 GND.n5057 0.0344674
R30059 GND.n6543 GND.n5076 0.0344674
R30060 GND.n5077 GND.n5076 0.0344674
R30061 GND.n5078 GND.n5077 0.0344674
R30062 GND.n6550 GND.n5078 0.0344674
R30063 GND.n6550 GND.n5097 0.0344674
R30064 GND.n5098 GND.n5097 0.0344674
R30065 GND.n5099 GND.n5098 0.0344674
R30066 GND.n6557 GND.n5099 0.0344674
R30067 GND.n6557 GND.n5118 0.0344674
R30068 GND.n5119 GND.n5118 0.0344674
R30069 GND.n5120 GND.n5119 0.0344674
R30070 GND.n6564 GND.n5120 0.0344674
R30071 GND.n6564 GND.n5139 0.0344674
R30072 GND.n5140 GND.n5139 0.0344674
R30073 GND.n5141 GND.n5140 0.0344674
R30074 GND.n6571 GND.n5141 0.0344674
R30075 GND.n6571 GND.n5160 0.0344674
R30076 GND.n5161 GND.n5160 0.0344674
R30077 GND.n5162 GND.n5161 0.0344674
R30078 GND.n6572 GND.n5162 0.0344674
R30079 GND.n6572 GND.n5179 0.0344674
R30080 GND.n5180 GND.n5179 0.0344674
R30081 GND.n5181 GND.n5180 0.0344674
R30082 GND.n6774 GND.n5181 0.0344674
R30083 GND.n6775 GND.n6774 0.0344674
R30084 GND.n6775 GND.n5283 0.0344674
R30085 GND.n6783 GND.n5283 0.0344674
R30086 GND.n6783 GND.n5279 0.0344674
R30087 GND.n6792 GND.n5279 0.0344674
R30088 GND.n6793 GND.n6792 0.0344674
R30089 GND.n6793 GND.n134 0.0344674
R30090 GND.n135 GND.n134 0.0344674
R30091 GND.n136 GND.n135 0.0344674
R30092 GND.n6796 GND.n136 0.0344674
R30093 GND.n6796 GND.n154 0.0344674
R30094 GND.n155 GND.n154 0.0344674
R30095 GND.n156 GND.n155 0.0344674
R30096 GND.n6803 GND.n156 0.0344674
R30097 GND.n6803 GND.n175 0.0344674
R30098 GND.n176 GND.n175 0.0344674
R30099 GND.n177 GND.n176 0.0344674
R30100 GND.n6810 GND.n177 0.0344674
R30101 GND.n6810 GND.n196 0.0344674
R30102 GND.n197 GND.n196 0.0344674
R30103 GND.n198 GND.n197 0.0344674
R30104 GND.n6817 GND.n198 0.0344674
R30105 GND.n6817 GND.n217 0.0344674
R30106 GND.n218 GND.n217 0.0344674
R30107 GND.n219 GND.n218 0.0344674
R30108 GND.n6824 GND.n219 0.0344674
R30109 GND.n6824 GND.n238 0.0344674
R30110 GND.n239 GND.n238 0.0344674
R30111 GND.n240 GND.n239 0.0344674
R30112 GND.n6830 GND.n240 0.0344674
R30113 GND.n6830 GND.n258 0.0344674
R30114 GND.n259 GND.n258 0.0344674
R30115 GND.n260 GND.n259 0.0344674
R30116 GND.n9739 GND.n260 0.0344674
R30117 GND.n9739 GND.n279 0.0344674
R30118 GND.n280 GND.n279 0.0344674
R30119 GND.n281 GND.n280 0.0344674
R30120 GND.n9754 GND.n281 0.0344674
R30121 GND.n9754 GND.n300 0.0344674
R30122 GND.n301 GND.n300 0.0344674
R30123 GND.n302 GND.n301 0.0344674
R30124 GND.n9769 GND.n302 0.0344674
R30125 GND.n9769 GND.n321 0.0344674
R30126 GND.n322 GND.n321 0.0344674
R30127 GND.n323 GND.n322 0.0344674
R30128 GND.n9784 GND.n323 0.0344674
R30129 GND.n9784 GND.n342 0.0344674
R30130 GND.n343 GND.n342 0.0344674
R30131 GND.n344 GND.n343 0.0344674
R30132 GND.n10108 GND.n344 0.0344674
R30133 GND.n10108 GND.n363 0.0344674
R30134 GND.n364 GND.n363 0.0344674
R30135 GND.n365 GND.n364 0.0344674
R30136 GND.n10115 GND.n365 0.0344674
R30137 GND.n10115 GND.n382 0.0344674
R30138 GND.n383 GND.n382 0.0344674
R30139 GND.n384 GND.n383 0.0344674
R30140 GND.n10122 GND.n384 0.0344674
R30141 GND.n10122 GND.n401 0.0344674
R30142 GND.n402 GND.n401 0.0344674
R30143 GND.n403 GND.n402 0.0344674
R30144 GND.n419 GND.n403 0.0344674
R30145 GND.n10132 GND.n419 0.0344674
R30146 GND.n2932 GND.n1437 0.0344674
R30147 GND.n2933 GND.n2932 0.0344674
R30148 GND.n2933 GND.n2918 0.0344674
R30149 GND.n2950 GND.n2918 0.0344674
R30150 GND.n2950 GND.n2921 0.0344674
R30151 GND.n2921 GND.n2920 0.0344674
R30152 GND.n2920 GND.n2898 0.0344674
R30153 GND.n2967 GND.n2898 0.0344674
R30154 GND.n2967 GND.n2901 0.0344674
R30155 GND.n2901 GND.n2900 0.0344674
R30156 GND.n2900 GND.n2880 0.0344674
R30157 GND.n2991 GND.n2880 0.0344674
R30158 GND.n2991 GND.n2881 0.0344674
R30159 GND.n2987 GND.n2881 0.0344674
R30160 GND.n2987 GND.n2986 0.0344674
R30161 GND.n2986 GND.n2855 0.0344674
R30162 GND.n3024 GND.n2855 0.0344674
R30163 GND.n3024 GND.n2858 0.0344674
R30164 GND.n2858 GND.n2857 0.0344674
R30165 GND.n2857 GND.n2830 0.0344674
R30166 GND.n3057 GND.n2830 0.0344674
R30167 GND.n3057 GND.n2831 0.0344674
R30168 GND.n3053 GND.n2831 0.0344674
R30169 GND.n3053 GND.n3052 0.0344674
R30170 GND.n3052 GND.n2802 0.0344674
R30171 GND.n3094 GND.n2802 0.0344674
R30172 GND.n3094 GND.n2803 0.0344674
R30173 GND.n3090 GND.n2803 0.0344674
R30174 GND.n3090 GND.n3089 0.0344674
R30175 GND.n3089 GND.n2773 0.0344674
R30176 GND.n3132 GND.n2773 0.0344674
R30177 GND.n3132 GND.n2774 0.0344674
R30178 GND.n3128 GND.n2774 0.0344674
R30179 GND.n3128 GND.n3127 0.0344674
R30180 GND.n3127 GND.n2745 0.0344674
R30181 GND.n3170 GND.n2745 0.0344674
R30182 GND.n3170 GND.n2746 0.0344674
R30183 GND.n3166 GND.n2746 0.0344674
R30184 GND.n3166 GND.n3165 0.0344674
R30185 GND.n3165 GND.n2716 0.0344674
R30186 GND.n3207 GND.n2716 0.0344674
R30187 GND.n3207 GND.n2717 0.0344674
R30188 GND.n3203 GND.n2717 0.0344674
R30189 GND.n3203 GND.n3202 0.0344674
R30190 GND.n3202 GND.n2687 0.0344674
R30191 GND.n3244 GND.n2687 0.0344674
R30192 GND.n3244 GND.n2688 0.0344674
R30193 GND.n3240 GND.n2688 0.0344674
R30194 GND.n3240 GND.n3239 0.0344674
R30195 GND.n3239 GND.n2658 0.0344674
R30196 GND.n3281 GND.n2658 0.0344674
R30197 GND.n3281 GND.n2659 0.0344674
R30198 GND.n3277 GND.n2659 0.0344674
R30199 GND.n3277 GND.n3276 0.0344674
R30200 GND.n3276 GND.n2629 0.0344674
R30201 GND.n3317 GND.n2629 0.0344674
R30202 GND.n3317 GND.n2630 0.0344674
R30203 GND.n3313 GND.n2630 0.0344674
R30204 GND.n3313 GND.n2606 0.0344674
R30205 GND.n3546 GND.n2606 0.0344674
R30206 GND.n3546 GND.n2603 0.0344674
R30207 GND.n3550 GND.n2603 0.0344674
R30208 GND.n3551 GND.n3550 0.0344674
R30209 GND.n3551 GND.n1560 0.0344674
R30210 GND.n8113 GND.n1560 0.0344674
R30211 GND.n8113 GND.n1561 0.0344674
R30212 GND.n8109 GND.n1561 0.0344674
R30213 GND.n8109 GND.n8108 0.0344674
R30214 GND.n8108 GND.n8107 0.0344674
R30215 GND.n8107 GND.n1569 0.0344674
R30216 GND.n8103 GND.n1569 0.0344674
R30217 GND.n8103 GND.n8102 0.0344674
R30218 GND.n8102 GND.n8101 0.0344674
R30219 GND.n8101 GND.n1577 0.0344674
R30220 GND.n8097 GND.n1577 0.0344674
R30221 GND.n8097 GND.n8096 0.0344674
R30222 GND.n8096 GND.n8095 0.0344674
R30223 GND.n8095 GND.n1585 0.0344674
R30224 GND.n8091 GND.n1585 0.0344674
R30225 GND.n8091 GND.n8090 0.0344674
R30226 GND.n8090 GND.n8089 0.0344674
R30227 GND.n8089 GND.n1593 0.0344674
R30228 GND.n8085 GND.n1593 0.0344674
R30229 GND.n8085 GND.n8084 0.0344674
R30230 GND.n8084 GND.n8083 0.0344674
R30231 GND.n8083 GND.n1601 0.0344674
R30232 GND.n8079 GND.n1601 0.0344674
R30233 GND.n8079 GND.n8078 0.0344674
R30234 GND.n8078 GND.n8077 0.0344674
R30235 GND.n8077 GND.n1609 0.0344674
R30236 GND.n8073 GND.n1609 0.0344674
R30237 GND.n8073 GND.n8072 0.0344674
R30238 GND.n8072 GND.n8071 0.0344674
R30239 GND.n8071 GND.n1617 0.0344674
R30240 GND.n8067 GND.n1617 0.0344674
R30241 GND.n8067 GND.n8066 0.0344674
R30242 GND.n8066 GND.n8065 0.0344674
R30243 GND.n8065 GND.n1625 0.0344674
R30244 GND.n8061 GND.n1625 0.0344674
R30245 GND.n8061 GND.n8060 0.0344674
R30246 GND.n8060 GND.n8059 0.0344674
R30247 GND.n8059 GND.n1633 0.0344674
R30248 GND.n8055 GND.n1633 0.0344674
R30249 GND.n8055 GND.n8054 0.0344674
R30250 GND.n8054 GND.n8053 0.0344674
R30251 GND.n8053 GND.n1641 0.0344674
R30252 GND.n8049 GND.n1641 0.0344674
R30253 GND.n8049 GND.n8048 0.0344674
R30254 GND.n8048 GND.n8047 0.0344674
R30255 GND.n8047 GND.n1649 0.0344674
R30256 GND.n8043 GND.n1649 0.0344674
R30257 GND.n8043 GND.n8042 0.0344674
R30258 GND.n8042 GND.n8041 0.0344674
R30259 GND.n8041 GND.n1657 0.0344674
R30260 GND.n8037 GND.n1657 0.0344674
R30261 GND.n8037 GND.n8036 0.0344674
R30262 GND.n8036 GND.n8035 0.0344674
R30263 GND.n8035 GND.n1665 0.0344674
R30264 GND.n8031 GND.n1665 0.0344674
R30265 GND.n8031 GND.n8030 0.0344674
R30266 GND.n8030 GND.n8029 0.0344674
R30267 GND.n6356 GND.n5464 0.0248902
R30268 GND.n7738 GND.n2354 0.0248902
R30269 GND.n3337 GND.n1543 0.0187927
R30270 GND.n6746 GND.n118 0.0187927
R30271 GND.n7738 GND.n2358 0.00964634
R30272 GND.n6356 GND.n5465 0.00964634
R30273 VP.n204 VP.t0 243.97
R30274 VP.n207 VP.t3 243.255
R30275 VP.n206 VP.n205 223.454
R30276 VP.n204 VP.n203 223.454
R30277 VP.n130 VP.n127 161.3
R30278 VP.n132 VP.n131 161.3
R30279 VP.n133 VP.n126 161.3
R30280 VP.n135 VP.n134 161.3
R30281 VP.n136 VP.n125 161.3
R30282 VP.n138 VP.n137 161.3
R30283 VP.n139 VP.n124 161.3
R30284 VP.n141 VP.n140 161.3
R30285 VP.n142 VP.n123 161.3
R30286 VP.n144 VP.n143 161.3
R30287 VP.n145 VP.n122 161.3
R30288 VP.n147 VP.n146 161.3
R30289 VP.n149 VP.n148 161.3
R30290 VP.n150 VP.n120 161.3
R30291 VP.n152 VP.n151 161.3
R30292 VP.n153 VP.n119 161.3
R30293 VP.n155 VP.n154 161.3
R30294 VP.n156 VP.n118 161.3
R30295 VP.n158 VP.n157 161.3
R30296 VP.n159 VP.n117 161.3
R30297 VP.n161 VP.n160 161.3
R30298 VP.n162 VP.n115 161.3
R30299 VP.n164 VP.n163 161.3
R30300 VP.n165 VP.n114 161.3
R30301 VP.n167 VP.n166 161.3
R30302 VP.n168 VP.n113 161.3
R30303 VP.n170 VP.n169 161.3
R30304 VP.n171 VP.n112 161.3
R30305 VP.n173 VP.n172 161.3
R30306 VP.n174 VP.n111 161.3
R30307 VP.n176 VP.n175 161.3
R30308 VP.n177 VP.n110 161.3
R30309 VP.n179 VP.n178 161.3
R30310 VP.n180 VP.n108 161.3
R30311 VP.n182 VP.n181 161.3
R30312 VP.n183 VP.n107 161.3
R30313 VP.n185 VP.n184 161.3
R30314 VP.n186 VP.n106 161.3
R30315 VP.n188 VP.n187 161.3
R30316 VP.n189 VP.n105 161.3
R30317 VP.n191 VP.n190 161.3
R30318 VP.n192 VP.n104 161.3
R30319 VP.n194 VP.n193 161.3
R30320 VP.n195 VP.n103 161.3
R30321 VP.n197 VP.n196 161.3
R30322 VP.n198 VP.n102 161.3
R30323 VP.n200 VP.n199 161.3
R30324 VP.n99 VP.n98 161.3
R30325 VP.n97 VP.n1 161.3
R30326 VP.n96 VP.n95 161.3
R30327 VP.n94 VP.n2 161.3
R30328 VP.n93 VP.n92 161.3
R30329 VP.n91 VP.n3 161.3
R30330 VP.n90 VP.n89 161.3
R30331 VP.n88 VP.n4 161.3
R30332 VP.n87 VP.n86 161.3
R30333 VP.n85 VP.n5 161.3
R30334 VP.n84 VP.n83 161.3
R30335 VP.n82 VP.n6 161.3
R30336 VP.n81 VP.n80 161.3
R30337 VP.n78 VP.n7 161.3
R30338 VP.n77 VP.n76 161.3
R30339 VP.n75 VP.n8 161.3
R30340 VP.n74 VP.n73 161.3
R30341 VP.n72 VP.n9 161.3
R30342 VP.n71 VP.n70 161.3
R30343 VP.n69 VP.n10 161.3
R30344 VP.n68 VP.n67 161.3
R30345 VP.n66 VP.n11 161.3
R30346 VP.n65 VP.n64 161.3
R30347 VP.n63 VP.n12 161.3
R30348 VP.n62 VP.n61 161.3
R30349 VP.n59 VP.n13 161.3
R30350 VP.n58 VP.n57 161.3
R30351 VP.n56 VP.n14 161.3
R30352 VP.n55 VP.n54 161.3
R30353 VP.n53 VP.n15 161.3
R30354 VP.n52 VP.n51 161.3
R30355 VP.n50 VP.n16 161.3
R30356 VP.n49 VP.n48 161.3
R30357 VP.n47 VP.n17 161.3
R30358 VP.n46 VP.n45 161.3
R30359 VP.n44 VP.n43 161.3
R30360 VP.n42 VP.n19 161.3
R30361 VP.n41 VP.n40 161.3
R30362 VP.n39 VP.n20 161.3
R30363 VP.n38 VP.n37 161.3
R30364 VP.n36 VP.n21 161.3
R30365 VP.n35 VP.n34 161.3
R30366 VP.n33 VP.n22 161.3
R30367 VP.n32 VP.n31 161.3
R30368 VP.n30 VP.n23 161.3
R30369 VP.n29 VP.n28 161.3
R30370 VP.n27 VP.n24 161.3
R30371 VP.n192 VP.n191 70.1245
R30372 VP.n91 VP.n90 70.1245
R30373 VP.n174 VP.n173 63.3431
R30374 VP.n139 VP.n138 63.3431
R30375 VP.n36 VP.n35 63.3431
R30376 VP.n72 VP.n71 63.3431
R30377 VP.n201 VP.n101 63.0449
R30378 VP.n100 VP.n0 63.0449
R30379 VP.n26 VP.t14 58.8464
R30380 VP.n129 VP.t13 58.8463
R30381 VP.n202 VP.n201 57.3936
R30382 VP.n129 VP.n128 56.805
R30383 VP.n26 VP.n25 56.805
R30384 VP.n157 VP.n156 56.5617
R30385 VP.n156 VP.n155 56.5617
R30386 VP.n53 VP.n52 56.5617
R30387 VP.n54 VP.n53 56.5617
R30388 VP.n175 VP.n174 49.7803
R30389 VP.n138 VP.n125 49.7803
R30390 VP.n35 VP.n22 49.7803
R30391 VP.n73 VP.n72 49.7803
R30392 VP.n193 VP.n192 42.999
R30393 VP.n92 VP.n91 42.999
R30394 VP.n101 VP.t17 24.8779
R30395 VP.n109 VP.t6 24.8779
R30396 VP.n116 VP.t9 24.8779
R30397 VP.n121 VP.t16 24.8779
R30398 VP.n128 VP.t7 24.8779
R30399 VP.n25 VP.t8 24.8779
R30400 VP.n18 VP.t15 24.8779
R30401 VP.n60 VP.t10 24.8779
R30402 VP.n79 VP.t12 24.8779
R30403 VP.n0 VP.t11 24.8779
R30404 VP.n199 VP.n198 24.5923
R30405 VP.n198 VP.n197 24.5923
R30406 VP.n197 VP.n103 24.5923
R30407 VP.n193 VP.n103 24.5923
R30408 VP.n191 VP.n105 24.5923
R30409 VP.n187 VP.n105 24.5923
R30410 VP.n187 VP.n186 24.5923
R30411 VP.n186 VP.n185 24.5923
R30412 VP.n185 VP.n107 24.5923
R30413 VP.n181 VP.n180 24.5923
R30414 VP.n180 VP.n179 24.5923
R30415 VP.n179 VP.n110 24.5923
R30416 VP.n175 VP.n110 24.5923
R30417 VP.n173 VP.n112 24.5923
R30418 VP.n169 VP.n112 24.5923
R30419 VP.n169 VP.n168 24.5923
R30420 VP.n168 VP.n167 24.5923
R30421 VP.n167 VP.n114 24.5923
R30422 VP.n163 VP.n162 24.5923
R30423 VP.n162 VP.n161 24.5923
R30424 VP.n161 VP.n117 24.5923
R30425 VP.n157 VP.n117 24.5923
R30426 VP.n155 VP.n119 24.5923
R30427 VP.n151 VP.n119 24.5923
R30428 VP.n151 VP.n150 24.5923
R30429 VP.n150 VP.n149 24.5923
R30430 VP.n146 VP.n145 24.5923
R30431 VP.n145 VP.n144 24.5923
R30432 VP.n144 VP.n123 24.5923
R30433 VP.n140 VP.n123 24.5923
R30434 VP.n140 VP.n139 24.5923
R30435 VP.n134 VP.n125 24.5923
R30436 VP.n134 VP.n133 24.5923
R30437 VP.n133 VP.n132 24.5923
R30438 VP.n132 VP.n127 24.5923
R30439 VP.n29 VP.n24 24.5923
R30440 VP.n30 VP.n29 24.5923
R30441 VP.n31 VP.n30 24.5923
R30442 VP.n31 VP.n22 24.5923
R30443 VP.n37 VP.n36 24.5923
R30444 VP.n37 VP.n20 24.5923
R30445 VP.n41 VP.n20 24.5923
R30446 VP.n42 VP.n41 24.5923
R30447 VP.n43 VP.n42 24.5923
R30448 VP.n47 VP.n46 24.5923
R30449 VP.n48 VP.n47 24.5923
R30450 VP.n48 VP.n16 24.5923
R30451 VP.n52 VP.n16 24.5923
R30452 VP.n54 VP.n14 24.5923
R30453 VP.n58 VP.n14 24.5923
R30454 VP.n59 VP.n58 24.5923
R30455 VP.n61 VP.n59 24.5923
R30456 VP.n65 VP.n12 24.5923
R30457 VP.n66 VP.n65 24.5923
R30458 VP.n67 VP.n66 24.5923
R30459 VP.n67 VP.n10 24.5923
R30460 VP.n71 VP.n10 24.5923
R30461 VP.n73 VP.n8 24.5923
R30462 VP.n77 VP.n8 24.5923
R30463 VP.n78 VP.n77 24.5923
R30464 VP.n80 VP.n78 24.5923
R30465 VP.n84 VP.n6 24.5923
R30466 VP.n85 VP.n84 24.5923
R30467 VP.n86 VP.n85 24.5923
R30468 VP.n86 VP.n4 24.5923
R30469 VP.n90 VP.n4 24.5923
R30470 VP.n92 VP.n2 24.5923
R30471 VP.n96 VP.n2 24.5923
R30472 VP.n97 VP.n96 24.5923
R30473 VP.n98 VP.n97 24.5923
R30474 VP.n163 VP.n116 22.8709
R30475 VP.n149 VP.n121 22.8709
R30476 VP.n46 VP.n18 22.8709
R30477 VP.n61 VP.n60 22.8709
R30478 VP.n205 VP.t4 19.8005
R30479 VP.n205 VP.t2 19.8005
R30480 VP.n203 VP.t5 19.8005
R30481 VP.n203 VP.t1 19.8005
R30482 VP.n181 VP.n109 19.4281
R30483 VP.n128 VP.n127 19.4281
R30484 VP.n25 VP.n24 19.4281
R30485 VP.n80 VP.n79 19.4281
R30486 VP.n199 VP.n101 15.9852
R30487 VP.n98 VP.n0 15.9852
R30488 VP.n202 VP.n100 14.2914
R30489 VP VP.n208 13.3464
R30490 VP.n109 VP.n107 5.16479
R30491 VP.n79 VP.n6 5.16479
R30492 VP.n208 VP.n207 4.80222
R30493 VP.n116 VP.n114 1.72193
R30494 VP.n146 VP.n121 1.72193
R30495 VP.n43 VP.n18 1.72193
R30496 VP.n60 VP.n12 1.72193
R30497 VP.n208 VP.n202 0.972091
R30498 VP.n27 VP.n26 0.940476
R30499 VP.n130 VP.n129 0.940474
R30500 VP.n206 VP.n204 0.716017
R30501 VP.n207 VP.n206 0.716017
R30502 VP.n201 VP.n200 0.46582
R30503 VP.n100 VP.n99 0.46582
R30504 VP.n200 VP.n102 0.189894
R30505 VP.n196 VP.n102 0.189894
R30506 VP.n196 VP.n195 0.189894
R30507 VP.n195 VP.n194 0.189894
R30508 VP.n194 VP.n104 0.189894
R30509 VP.n190 VP.n104 0.189894
R30510 VP.n190 VP.n189 0.189894
R30511 VP.n189 VP.n188 0.189894
R30512 VP.n188 VP.n106 0.189894
R30513 VP.n184 VP.n106 0.189894
R30514 VP.n184 VP.n183 0.189894
R30515 VP.n183 VP.n182 0.189894
R30516 VP.n182 VP.n108 0.189894
R30517 VP.n178 VP.n108 0.189894
R30518 VP.n178 VP.n177 0.189894
R30519 VP.n177 VP.n176 0.189894
R30520 VP.n176 VP.n111 0.189894
R30521 VP.n172 VP.n111 0.189894
R30522 VP.n172 VP.n171 0.189894
R30523 VP.n171 VP.n170 0.189894
R30524 VP.n170 VP.n113 0.189894
R30525 VP.n166 VP.n113 0.189894
R30526 VP.n166 VP.n165 0.189894
R30527 VP.n165 VP.n164 0.189894
R30528 VP.n164 VP.n115 0.189894
R30529 VP.n160 VP.n115 0.189894
R30530 VP.n160 VP.n159 0.189894
R30531 VP.n159 VP.n158 0.189894
R30532 VP.n158 VP.n118 0.189894
R30533 VP.n154 VP.n118 0.189894
R30534 VP.n154 VP.n153 0.189894
R30535 VP.n153 VP.n152 0.189894
R30536 VP.n152 VP.n120 0.189894
R30537 VP.n148 VP.n120 0.189894
R30538 VP.n148 VP.n147 0.189894
R30539 VP.n147 VP.n122 0.189894
R30540 VP.n143 VP.n122 0.189894
R30541 VP.n143 VP.n142 0.189894
R30542 VP.n142 VP.n141 0.189894
R30543 VP.n141 VP.n124 0.189894
R30544 VP.n137 VP.n124 0.189894
R30545 VP.n137 VP.n136 0.189894
R30546 VP.n136 VP.n135 0.189894
R30547 VP.n135 VP.n126 0.189894
R30548 VP.n131 VP.n126 0.189894
R30549 VP.n131 VP.n130 0.189894
R30550 VP.n28 VP.n27 0.189894
R30551 VP.n28 VP.n23 0.189894
R30552 VP.n32 VP.n23 0.189894
R30553 VP.n33 VP.n32 0.189894
R30554 VP.n34 VP.n33 0.189894
R30555 VP.n34 VP.n21 0.189894
R30556 VP.n38 VP.n21 0.189894
R30557 VP.n39 VP.n38 0.189894
R30558 VP.n40 VP.n39 0.189894
R30559 VP.n40 VP.n19 0.189894
R30560 VP.n44 VP.n19 0.189894
R30561 VP.n45 VP.n44 0.189894
R30562 VP.n45 VP.n17 0.189894
R30563 VP.n49 VP.n17 0.189894
R30564 VP.n50 VP.n49 0.189894
R30565 VP.n51 VP.n50 0.189894
R30566 VP.n51 VP.n15 0.189894
R30567 VP.n55 VP.n15 0.189894
R30568 VP.n56 VP.n55 0.189894
R30569 VP.n57 VP.n56 0.189894
R30570 VP.n57 VP.n13 0.189894
R30571 VP.n62 VP.n13 0.189894
R30572 VP.n63 VP.n62 0.189894
R30573 VP.n64 VP.n63 0.189894
R30574 VP.n64 VP.n11 0.189894
R30575 VP.n68 VP.n11 0.189894
R30576 VP.n69 VP.n68 0.189894
R30577 VP.n70 VP.n69 0.189894
R30578 VP.n70 VP.n9 0.189894
R30579 VP.n74 VP.n9 0.189894
R30580 VP.n75 VP.n74 0.189894
R30581 VP.n76 VP.n75 0.189894
R30582 VP.n76 VP.n7 0.189894
R30583 VP.n81 VP.n7 0.189894
R30584 VP.n82 VP.n81 0.189894
R30585 VP.n83 VP.n82 0.189894
R30586 VP.n83 VP.n5 0.189894
R30587 VP.n87 VP.n5 0.189894
R30588 VP.n88 VP.n87 0.189894
R30589 VP.n89 VP.n88 0.189894
R30590 VP.n89 VP.n3 0.189894
R30591 VP.n93 VP.n3 0.189894
R30592 VP.n94 VP.n93 0.189894
R30593 VP.n95 VP.n94 0.189894
R30594 VP.n95 VP.n1 0.189894
R30595 VP.n99 VP.n1 0.189894
R30596 a_n7336_n129.n3 a_n7336_n129.t27 161.155
R30597 a_n7336_n129.n4 a_n7336_n129.t7 161.155
R30598 a_n7336_n129.n5 a_n7336_n129.t8 161.155
R30599 a_n7336_n129.n6 a_n7336_n129.t26 161.155
R30600 a_n7336_n129.n1 a_n7336_n129.t23 52.3106
R30601 a_n7336_n129.n1 a_n7336_n129.t13 52.3106
R30602 a_n7336_n129.n2 a_n7336_n129.t9 52.3106
R30603 a_n7336_n129.n19 a_n7336_n129.t5 52.3097
R30604 a_n7336_n129.n17 a_n7336_n129.t15 52.3096
R30605 a_n7336_n129.n0 a_n7336_n129.t12 52.3096
R30606 a_n7336_n129.n0 a_n7336_n129.t2 52.3096
R30607 a_n7336_n129.n8 a_n7336_n129.t22 52.3096
R30608 a_n7336_n129.n21 a_n7336_n129.n20 45.0312
R30609 a_n7336_n129.n23 a_n7336_n129.n22 45.0312
R30610 a_n7336_n129.n25 a_n7336_n129.n24 45.0312
R30611 a_n7336_n129.n27 a_n7336_n129.n26 45.0312
R30612 a_n7336_n129.n16 a_n7336_n129.n15 45.0311
R30613 a_n7336_n129.n14 a_n7336_n129.n13 45.0311
R30614 a_n7336_n129.n12 a_n7336_n129.n11 45.0311
R30615 a_n7336_n129.n10 a_n7336_n129.n9 45.0311
R30616 a_n7336_n129.n7 a_n7336_n129.n2 11.5857
R30617 a_n7336_n129.n19 a_n7336_n129.n18 11.5857
R30618 a_n7336_n129.n20 a_n7336_n129.t0 7.27991
R30619 a_n7336_n129.n20 a_n7336_n129.t3 7.27991
R30620 a_n7336_n129.n22 a_n7336_n129.t25 7.27991
R30621 a_n7336_n129.n22 a_n7336_n129.t4 7.27991
R30622 a_n7336_n129.n24 a_n7336_n129.t10 7.27991
R30623 a_n7336_n129.n24 a_n7336_n129.t19 7.27991
R30624 a_n7336_n129.n15 a_n7336_n129.t16 7.27991
R30625 a_n7336_n129.n15 a_n7336_n129.t14 7.27991
R30626 a_n7336_n129.n13 a_n7336_n129.t18 7.27991
R30627 a_n7336_n129.n13 a_n7336_n129.t11 7.27991
R30628 a_n7336_n129.n11 a_n7336_n129.t21 7.27991
R30629 a_n7336_n129.n11 a_n7336_n129.t24 7.27991
R30630 a_n7336_n129.n9 a_n7336_n129.t1 7.27991
R30631 a_n7336_n129.n9 a_n7336_n129.t6 7.27991
R30632 a_n7336_n129.t20 a_n7336_n129.n27 7.27991
R30633 a_n7336_n129.n27 a_n7336_n129.t17 7.27991
R30634 a_n7336_n129.n18 a_n7336_n129.n3 5.79551
R30635 a_n7336_n129.n8 a_n7336_n129.n7 5.688
R30636 a_n7336_n129.n18 a_n7336_n129.n17 5.688
R30637 a_n7336_n129.n7 a_n7336_n129.n6 5.06586
R30638 a_n7336_n129.n25 a_n7336_n129.n1 1.90855
R30639 a_n7336_n129.n14 a_n7336_n129.n0 1.90855
R30640 a_n7336_n129.n10 a_n7336_n129.n8 1.70452
R30641 a_n7336_n129.n12 a_n7336_n129.n10 1.70452
R30642 a_n7336_n129.n0 a_n7336_n129.n12 1.70452
R30643 a_n7336_n129.n16 a_n7336_n129.n14 1.70452
R30644 a_n7336_n129.n17 a_n7336_n129.n16 1.70452
R30645 a_n7336_n129.n26 a_n7336_n129.n2 1.70452
R30646 a_n7336_n129.n26 a_n7336_n129.n25 1.70452
R30647 a_n7336_n129.n1 a_n7336_n129.n23 1.70452
R30648 a_n7336_n129.n23 a_n7336_n129.n21 1.70452
R30649 a_n7336_n129.n21 a_n7336_n129.n19 1.70452
R30650 a_n7336_n129.n6 a_n7336_n129.n5 0.857089
R30651 a_n7336_n129.n5 a_n7336_n129.n4 0.857089
R30652 a_n7336_n129.n4 a_n7336_n129.n3 0.857089
R30653 VN.n204 VN.t3 243.97
R30654 VN.n207 VN.t1 243.255
R30655 VN.n204 VN.n203 223.454
R30656 VN.n206 VN.n205 223.454
R30657 VN.n200 VN.n199 161.3
R30658 VN.n198 VN.n102 161.3
R30659 VN.n197 VN.n196 161.3
R30660 VN.n195 VN.n103 161.3
R30661 VN.n194 VN.n193 161.3
R30662 VN.n192 VN.n104 161.3
R30663 VN.n191 VN.n190 161.3
R30664 VN.n189 VN.n105 161.3
R30665 VN.n188 VN.n187 161.3
R30666 VN.n186 VN.n106 161.3
R30667 VN.n185 VN.n184 161.3
R30668 VN.n183 VN.n107 161.3
R30669 VN.n182 VN.n181 161.3
R30670 VN.n179 VN.n108 161.3
R30671 VN.n178 VN.n177 161.3
R30672 VN.n176 VN.n109 161.3
R30673 VN.n175 VN.n174 161.3
R30674 VN.n173 VN.n110 161.3
R30675 VN.n172 VN.n171 161.3
R30676 VN.n170 VN.n111 161.3
R30677 VN.n169 VN.n168 161.3
R30678 VN.n167 VN.n112 161.3
R30679 VN.n166 VN.n165 161.3
R30680 VN.n164 VN.n113 161.3
R30681 VN.n163 VN.n162 161.3
R30682 VN.n160 VN.n114 161.3
R30683 VN.n159 VN.n158 161.3
R30684 VN.n157 VN.n115 161.3
R30685 VN.n156 VN.n155 161.3
R30686 VN.n154 VN.n116 161.3
R30687 VN.n153 VN.n152 161.3
R30688 VN.n151 VN.n117 161.3
R30689 VN.n150 VN.n149 161.3
R30690 VN.n148 VN.n118 161.3
R30691 VN.n147 VN.n146 161.3
R30692 VN.n145 VN.n144 161.3
R30693 VN.n143 VN.n120 161.3
R30694 VN.n142 VN.n141 161.3
R30695 VN.n140 VN.n121 161.3
R30696 VN.n139 VN.n138 161.3
R30697 VN.n137 VN.n122 161.3
R30698 VN.n136 VN.n135 161.3
R30699 VN.n134 VN.n123 161.3
R30700 VN.n133 VN.n132 161.3
R30701 VN.n131 VN.n124 161.3
R30702 VN.n130 VN.n129 161.3
R30703 VN.n128 VN.n125 161.3
R30704 VN.n29 VN.n26 161.3
R30705 VN.n31 VN.n30 161.3
R30706 VN.n32 VN.n25 161.3
R30707 VN.n34 VN.n33 161.3
R30708 VN.n35 VN.n24 161.3
R30709 VN.n37 VN.n36 161.3
R30710 VN.n38 VN.n23 161.3
R30711 VN.n40 VN.n39 161.3
R30712 VN.n41 VN.n22 161.3
R30713 VN.n43 VN.n42 161.3
R30714 VN.n44 VN.n21 161.3
R30715 VN.n46 VN.n45 161.3
R30716 VN.n48 VN.n47 161.3
R30717 VN.n49 VN.n19 161.3
R30718 VN.n51 VN.n50 161.3
R30719 VN.n52 VN.n18 161.3
R30720 VN.n54 VN.n53 161.3
R30721 VN.n55 VN.n17 161.3
R30722 VN.n57 VN.n56 161.3
R30723 VN.n58 VN.n16 161.3
R30724 VN.n60 VN.n59 161.3
R30725 VN.n61 VN.n14 161.3
R30726 VN.n63 VN.n62 161.3
R30727 VN.n64 VN.n13 161.3
R30728 VN.n66 VN.n65 161.3
R30729 VN.n67 VN.n12 161.3
R30730 VN.n69 VN.n68 161.3
R30731 VN.n70 VN.n11 161.3
R30732 VN.n72 VN.n71 161.3
R30733 VN.n73 VN.n10 161.3
R30734 VN.n75 VN.n74 161.3
R30735 VN.n76 VN.n9 161.3
R30736 VN.n78 VN.n77 161.3
R30737 VN.n79 VN.n7 161.3
R30738 VN.n81 VN.n80 161.3
R30739 VN.n82 VN.n6 161.3
R30740 VN.n84 VN.n83 161.3
R30741 VN.n85 VN.n5 161.3
R30742 VN.n87 VN.n86 161.3
R30743 VN.n88 VN.n4 161.3
R30744 VN.n90 VN.n89 161.3
R30745 VN.n91 VN.n3 161.3
R30746 VN.n93 VN.n92 161.3
R30747 VN.n94 VN.n2 161.3
R30748 VN.n96 VN.n95 161.3
R30749 VN.n97 VN.n1 161.3
R30750 VN.n99 VN.n98 161.3
R30751 VN.n192 VN.n191 70.1245
R30752 VN.n91 VN.n90 70.1245
R30753 VN.n137 VN.n136 63.3431
R30754 VN.n173 VN.n172 63.3431
R30755 VN.n73 VN.n72 63.3431
R30756 VN.n38 VN.n37 63.3431
R30757 VN.n201 VN.n101 63.0449
R30758 VN.n100 VN.n0 63.0449
R30759 VN.n127 VN.t17 58.8464
R30760 VN.n28 VN.t6 58.8463
R30761 VN.n202 VN.n201 57.1777
R30762 VN.n28 VN.n27 56.805
R30763 VN.n127 VN.n126 56.805
R30764 VN.n154 VN.n153 56.5617
R30765 VN.n155 VN.n154 56.5617
R30766 VN.n56 VN.n55 56.5617
R30767 VN.n55 VN.n54 56.5617
R30768 VN.n136 VN.n123 49.7803
R30769 VN.n174 VN.n173 49.7803
R30770 VN.n74 VN.n73 49.7803
R30771 VN.n37 VN.n24 49.7803
R30772 VN.n193 VN.n192 42.999
R30773 VN.n92 VN.n91 42.999
R30774 VN.n126 VN.t9 24.8779
R30775 VN.n119 VN.t7 24.8779
R30776 VN.n161 VN.t12 24.8779
R30777 VN.n180 VN.t15 24.8779
R30778 VN.n101 VN.t14 24.8779
R30779 VN.n0 VN.t10 24.8779
R30780 VN.n8 VN.t11 24.8779
R30781 VN.n15 VN.t16 24.8779
R30782 VN.n20 VN.t8 24.8779
R30783 VN.n27 VN.t13 24.8779
R30784 VN.n130 VN.n125 24.5923
R30785 VN.n131 VN.n130 24.5923
R30786 VN.n132 VN.n131 24.5923
R30787 VN.n132 VN.n123 24.5923
R30788 VN.n138 VN.n137 24.5923
R30789 VN.n138 VN.n121 24.5923
R30790 VN.n142 VN.n121 24.5923
R30791 VN.n143 VN.n142 24.5923
R30792 VN.n144 VN.n143 24.5923
R30793 VN.n148 VN.n147 24.5923
R30794 VN.n149 VN.n148 24.5923
R30795 VN.n149 VN.n117 24.5923
R30796 VN.n153 VN.n117 24.5923
R30797 VN.n155 VN.n115 24.5923
R30798 VN.n159 VN.n115 24.5923
R30799 VN.n160 VN.n159 24.5923
R30800 VN.n162 VN.n160 24.5923
R30801 VN.n166 VN.n113 24.5923
R30802 VN.n167 VN.n166 24.5923
R30803 VN.n168 VN.n167 24.5923
R30804 VN.n168 VN.n111 24.5923
R30805 VN.n172 VN.n111 24.5923
R30806 VN.n174 VN.n109 24.5923
R30807 VN.n178 VN.n109 24.5923
R30808 VN.n179 VN.n178 24.5923
R30809 VN.n181 VN.n179 24.5923
R30810 VN.n185 VN.n107 24.5923
R30811 VN.n186 VN.n185 24.5923
R30812 VN.n187 VN.n186 24.5923
R30813 VN.n187 VN.n105 24.5923
R30814 VN.n191 VN.n105 24.5923
R30815 VN.n193 VN.n103 24.5923
R30816 VN.n197 VN.n103 24.5923
R30817 VN.n198 VN.n197 24.5923
R30818 VN.n199 VN.n198 24.5923
R30819 VN.n98 VN.n97 24.5923
R30820 VN.n97 VN.n96 24.5923
R30821 VN.n96 VN.n2 24.5923
R30822 VN.n92 VN.n2 24.5923
R30823 VN.n90 VN.n4 24.5923
R30824 VN.n86 VN.n4 24.5923
R30825 VN.n86 VN.n85 24.5923
R30826 VN.n85 VN.n84 24.5923
R30827 VN.n84 VN.n6 24.5923
R30828 VN.n80 VN.n79 24.5923
R30829 VN.n79 VN.n78 24.5923
R30830 VN.n78 VN.n9 24.5923
R30831 VN.n74 VN.n9 24.5923
R30832 VN.n72 VN.n11 24.5923
R30833 VN.n68 VN.n11 24.5923
R30834 VN.n68 VN.n67 24.5923
R30835 VN.n67 VN.n66 24.5923
R30836 VN.n66 VN.n13 24.5923
R30837 VN.n62 VN.n61 24.5923
R30838 VN.n61 VN.n60 24.5923
R30839 VN.n60 VN.n16 24.5923
R30840 VN.n56 VN.n16 24.5923
R30841 VN.n54 VN.n18 24.5923
R30842 VN.n50 VN.n18 24.5923
R30843 VN.n50 VN.n49 24.5923
R30844 VN.n49 VN.n48 24.5923
R30845 VN.n45 VN.n44 24.5923
R30846 VN.n44 VN.n43 24.5923
R30847 VN.n43 VN.n22 24.5923
R30848 VN.n39 VN.n22 24.5923
R30849 VN.n39 VN.n38 24.5923
R30850 VN.n33 VN.n24 24.5923
R30851 VN.n33 VN.n32 24.5923
R30852 VN.n32 VN.n31 24.5923
R30853 VN.n31 VN.n26 24.5923
R30854 VN.n147 VN.n119 22.8709
R30855 VN.n162 VN.n161 22.8709
R30856 VN.n62 VN.n15 22.8709
R30857 VN.n48 VN.n20 22.8709
R30858 VN VN.n208 20.1061
R30859 VN.n203 VN.t4 19.8005
R30860 VN.n203 VN.t0 19.8005
R30861 VN.n205 VN.t5 19.8005
R30862 VN.n205 VN.t2 19.8005
R30863 VN.n126 VN.n125 19.4281
R30864 VN.n181 VN.n180 19.4281
R30865 VN.n80 VN.n8 19.4281
R30866 VN.n27 VN.n26 19.4281
R30867 VN.n199 VN.n101 15.9852
R30868 VN.n98 VN.n0 15.9852
R30869 VN.n202 VN.n100 14.0755
R30870 VN.n180 VN.n107 5.16479
R30871 VN.n8 VN.n6 5.16479
R30872 VN.n208 VN.n207 5.04791
R30873 VN.n144 VN.n119 1.72193
R30874 VN.n161 VN.n113 1.72193
R30875 VN.n15 VN.n13 1.72193
R30876 VN.n45 VN.n20 1.72193
R30877 VN.n208 VN.n202 1.188
R30878 VN.n128 VN.n127 0.940476
R30879 VN.n29 VN.n28 0.940474
R30880 VN.n207 VN.n206 0.716017
R30881 VN.n206 VN.n204 0.716017
R30882 VN.n201 VN.n200 0.46582
R30883 VN.n100 VN.n99 0.46582
R30884 VN.n129 VN.n128 0.189894
R30885 VN.n129 VN.n124 0.189894
R30886 VN.n133 VN.n124 0.189894
R30887 VN.n134 VN.n133 0.189894
R30888 VN.n135 VN.n134 0.189894
R30889 VN.n135 VN.n122 0.189894
R30890 VN.n139 VN.n122 0.189894
R30891 VN.n140 VN.n139 0.189894
R30892 VN.n141 VN.n140 0.189894
R30893 VN.n141 VN.n120 0.189894
R30894 VN.n145 VN.n120 0.189894
R30895 VN.n146 VN.n145 0.189894
R30896 VN.n146 VN.n118 0.189894
R30897 VN.n150 VN.n118 0.189894
R30898 VN.n151 VN.n150 0.189894
R30899 VN.n152 VN.n151 0.189894
R30900 VN.n152 VN.n116 0.189894
R30901 VN.n156 VN.n116 0.189894
R30902 VN.n157 VN.n156 0.189894
R30903 VN.n158 VN.n157 0.189894
R30904 VN.n158 VN.n114 0.189894
R30905 VN.n163 VN.n114 0.189894
R30906 VN.n164 VN.n163 0.189894
R30907 VN.n165 VN.n164 0.189894
R30908 VN.n165 VN.n112 0.189894
R30909 VN.n169 VN.n112 0.189894
R30910 VN.n170 VN.n169 0.189894
R30911 VN.n171 VN.n170 0.189894
R30912 VN.n171 VN.n110 0.189894
R30913 VN.n175 VN.n110 0.189894
R30914 VN.n176 VN.n175 0.189894
R30915 VN.n177 VN.n176 0.189894
R30916 VN.n177 VN.n108 0.189894
R30917 VN.n182 VN.n108 0.189894
R30918 VN.n183 VN.n182 0.189894
R30919 VN.n184 VN.n183 0.189894
R30920 VN.n184 VN.n106 0.189894
R30921 VN.n188 VN.n106 0.189894
R30922 VN.n189 VN.n188 0.189894
R30923 VN.n190 VN.n189 0.189894
R30924 VN.n190 VN.n104 0.189894
R30925 VN.n194 VN.n104 0.189894
R30926 VN.n195 VN.n194 0.189894
R30927 VN.n196 VN.n195 0.189894
R30928 VN.n196 VN.n102 0.189894
R30929 VN.n200 VN.n102 0.189894
R30930 VN.n99 VN.n1 0.189894
R30931 VN.n95 VN.n1 0.189894
R30932 VN.n95 VN.n94 0.189894
R30933 VN.n94 VN.n93 0.189894
R30934 VN.n93 VN.n3 0.189894
R30935 VN.n89 VN.n3 0.189894
R30936 VN.n89 VN.n88 0.189894
R30937 VN.n88 VN.n87 0.189894
R30938 VN.n87 VN.n5 0.189894
R30939 VN.n83 VN.n5 0.189894
R30940 VN.n83 VN.n82 0.189894
R30941 VN.n82 VN.n81 0.189894
R30942 VN.n81 VN.n7 0.189894
R30943 VN.n77 VN.n7 0.189894
R30944 VN.n77 VN.n76 0.189894
R30945 VN.n76 VN.n75 0.189894
R30946 VN.n75 VN.n10 0.189894
R30947 VN.n71 VN.n10 0.189894
R30948 VN.n71 VN.n70 0.189894
R30949 VN.n70 VN.n69 0.189894
R30950 VN.n69 VN.n12 0.189894
R30951 VN.n65 VN.n12 0.189894
R30952 VN.n65 VN.n64 0.189894
R30953 VN.n64 VN.n63 0.189894
R30954 VN.n63 VN.n14 0.189894
R30955 VN.n59 VN.n14 0.189894
R30956 VN.n59 VN.n58 0.189894
R30957 VN.n58 VN.n57 0.189894
R30958 VN.n57 VN.n17 0.189894
R30959 VN.n53 VN.n17 0.189894
R30960 VN.n53 VN.n52 0.189894
R30961 VN.n52 VN.n51 0.189894
R30962 VN.n51 VN.n19 0.189894
R30963 VN.n47 VN.n19 0.189894
R30964 VN.n47 VN.n46 0.189894
R30965 VN.n46 VN.n21 0.189894
R30966 VN.n42 VN.n21 0.189894
R30967 VN.n42 VN.n41 0.189894
R30968 VN.n41 VN.n40 0.189894
R30969 VN.n40 VN.n23 0.189894
R30970 VN.n36 VN.n23 0.189894
R30971 VN.n36 VN.n35 0.189894
R30972 VN.n35 VN.n34 0.189894
R30973 VN.n34 VN.n25 0.189894
R30974 VN.n30 VN.n25 0.189894
R30975 VN.n30 VN.n29 0.189894
R30976 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t10 146
R30977 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.t8 143.429
R30978 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.t11 143.429
R30979 DIFFPAIR_BIAS.n0 DIFFPAIR_BIAS.t9 143.429
R30980 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t2 108.409
R30981 DIFFPAIR_BIAS.n4 DIFFPAIR_BIAS.t6 105.838
R30982 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.t0 105.838
R30983 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.t4 105.838
R30984 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t3 94.5196
R30985 DIFFPAIR_BIAS.n1 DIFFPAIR_BIAS.t7 93.6631
R30986 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.t1 93.6631
R30987 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.t5 93.6631
R30988 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n6 5.59755
R30989 DIFFPAIR_BIAS.n8 DIFFPAIR_BIAS.n7 4.34994
R30990 DIFFPAIR_BIAS.n7 DIFFPAIR_BIAS.n3 4.25114
R30991 DIFFPAIR_BIAS.n6 DIFFPAIR_BIAS.n5 2.57195
R30992 DIFFPAIR_BIAS.n5 DIFFPAIR_BIAS.n4 2.57195
R30993 DIFFPAIR_BIAS.n9 DIFFPAIR_BIAS.n8 2.57192
R30994 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n9 1.78314
R30995 DIFFPAIR_BIAS.n3 DIFFPAIR_BIAS.n2 0.857089
R30996 DIFFPAIR_BIAS.n2 DIFFPAIR_BIAS.n1 0.857089
R30997 DIFFPAIR_BIAS DIFFPAIR_BIAS.n10 0.68425
R30998 DIFFPAIR_BIAS.n10 DIFFPAIR_BIAS.n0 0.498588
R30999 a_n7981_10383.n3 a_n7981_10383.n1 96.0321
R31000 a_n7981_10383.n6 a_n7981_10383.n4 95.3226
R31001 a_n7981_10383.n6 a_n7981_10383.n5 94.7763
R31002 a_n7981_10383.n3 a_n7981_10383.n2 94.7752
R31003 a_n7981_10383.n11 a_n7981_10383.t4 89.0675
R31004 a_n7981_10383.n8 a_n7981_10383.t5 87.8118
R31005 a_n7981_10383.n0 a_n7981_10383.t0 87.8118
R31006 a_n7981_10383.n0 a_n7981_10383.t1 87.8118
R31007 a_n7981_10383.n10 a_n7981_10383.n9 75.1885
R31008 a_n7981_10383.n12 a_n7981_10383.n11 75.1885
R31009 a_n7981_10383.n7 a_n7981_10383.n6 15.9535
R31010 a_n7981_10383.n7 a_n7981_10383.n3 12.7231
R31011 a_n7981_10383.n9 a_n7981_10383.t6 12.6238
R31012 a_n7981_10383.n9 a_n7981_10383.t3 12.6238
R31013 a_n7981_10383.n2 a_n7981_10383.t13 12.6238
R31014 a_n7981_10383.n2 a_n7981_10383.t12 12.6238
R31015 a_n7981_10383.n1 a_n7981_10383.t11 12.6238
R31016 a_n7981_10383.n1 a_n7981_10383.t8 12.6238
R31017 a_n7981_10383.n5 a_n7981_10383.t10 12.6238
R31018 a_n7981_10383.n5 a_n7981_10383.t14 12.6238
R31019 a_n7981_10383.n4 a_n7981_10383.t15 12.6238
R31020 a_n7981_10383.n4 a_n7981_10383.t9 12.6238
R31021 a_n7981_10383.n12 a_n7981_10383.t2 12.6238
R31022 a_n7981_10383.t7 a_n7981_10383.n12 12.6238
R31023 a_n7981_10383.n8 a_n7981_10383.n7 5.53642
R31024 a_n7981_10383.n11 a_n7981_10383.n0 1.55438
R31025 a_n7981_10383.n0 a_n7981_10383.n10 1.25625
R31026 a_n7981_10383.n10 a_n7981_10383.n8 1.25625
C0 VP DIFFPAIR_BIAS 1.8e-19
C1 VN CS_BIAS 0.358004f
C2 VN DIFFPAIR_BIAS 9.49e-20
C3 a_8109_10383# VDD 1.56827f
C4 VDD VOUT 62.338398f
C5 VDD VN 0.212967f
C6 VOUT VP 4.24797f
C7 a_n9139_10383# VDD 1.56831f
C8 VOUT VN 1.31691f
C9 VP VN 18.5785f
C10 VOUT CS_BIAS 62.7803f
C11 VP CS_BIAS 0.446266f
C12 DIFFPAIR_BIAS GND 37.021748f
C13 CS_BIAS GND 0.322645p
C14 VN GND 66.9698f
C15 VP GND 52.80977f
C16 VOUT GND 0.159031p
C17 VDD GND 0.828995p
C18 a_8109_10383# GND 0.484863f
C19 a_n9139_10383# GND 0.484697f
C20 a_n7981_10383.n0 GND 3.10977f
C21 a_n7981_10383.t2 GND 0.154859f
C22 a_n7981_10383.t4 GND 0.969734f
C23 a_n7981_10383.t11 GND 0.154859f
C24 a_n7981_10383.t8 GND 0.154859f
C25 a_n7981_10383.n1 GND 0.881751f
C26 a_n7981_10383.t13 GND 0.154859f
C27 a_n7981_10383.t12 GND 0.154859f
C28 a_n7981_10383.n2 GND 0.856179f
C29 a_n7981_10383.n3 GND 6.72004f
C30 a_n7981_10383.t15 GND 0.154859f
C31 a_n7981_10383.t9 GND 0.154859f
C32 a_n7981_10383.n4 GND 0.877872f
C33 a_n7981_10383.t10 GND 0.154859f
C34 a_n7981_10383.t14 GND 0.154859f
C35 a_n7981_10383.n5 GND 0.856182f
C36 a_n7981_10383.n6 GND 14.027901f
C37 a_n7981_10383.n7 GND 4.11102f
C38 a_n7981_10383.t5 GND 0.949807f
C39 a_n7981_10383.n8 GND 2.45428f
C40 a_n7981_10383.t6 GND 0.154859f
C41 a_n7981_10383.t3 GND 0.154859f
C42 a_n7981_10383.n9 GND 0.717241f
C43 a_n7981_10383.n10 GND 1.94979f
C44 a_n7981_10383.t0 GND 0.949807f
C45 a_n7981_10383.t1 GND 0.949807f
C46 a_n7981_10383.n11 GND 3.34324f
C47 a_n7981_10383.n12 GND 0.717241f
C48 a_n7981_10383.t7 GND 0.154859f
C49 DIFFPAIR_BIAS.t9 GND 0.095723f
C50 DIFFPAIR_BIAS.t10 GND 0.096863f
C51 DIFFPAIR_BIAS.n0 GND 0.112211f
C52 DIFFPAIR_BIAS.t3 GND 0.05722f
C53 DIFFPAIR_BIAS.t7 GND 0.056272f
C54 DIFFPAIR_BIAS.n1 GND 0.219023f
C55 DIFFPAIR_BIAS.t1 GND 0.056272f
C56 DIFFPAIR_BIAS.n2 GND 0.115359f
C57 DIFFPAIR_BIAS.t5 GND 0.056272f
C58 DIFFPAIR_BIAS.n3 GND 0.135895f
C59 DIFFPAIR_BIAS.t4 GND 0.091422f
C60 DIFFPAIR_BIAS.t0 GND 0.091422f
C61 DIFFPAIR_BIAS.t6 GND 0.091422f
C62 DIFFPAIR_BIAS.t2 GND 0.092641f
C63 DIFFPAIR_BIAS.n4 GND 0.111526f
C64 DIFFPAIR_BIAS.n5 GND 0.061371f
C65 DIFFPAIR_BIAS.n6 GND 0.066549f
C66 DIFFPAIR_BIAS.n7 GND 0.125951f
C67 DIFFPAIR_BIAS.t11 GND 0.095723f
C68 DIFFPAIR_BIAS.n8 GND 0.056034f
C69 DIFFPAIR_BIAS.t8 GND 0.095723f
C70 DIFFPAIR_BIAS.n9 GND 0.056343f
C71 DIFFPAIR_BIAS.n10 GND 0.035819f
C72 VN.t10 GND 0.924272f
C73 VN.n0 GND 0.393886f
C74 VN.n1 GND 0.012255f
C75 VN.n2 GND 0.022726f
C76 VN.n3 GND 0.012255f
C77 VN.n4 GND 0.022726f
C78 VN.n5 GND 0.012255f
C79 VN.n6 GND 0.013863f
C80 VN.n7 GND 0.012255f
C81 VN.t11 GND 0.924272f
C82 VN.n8 GND 0.33942f
C83 VN.n9 GND 0.022726f
C84 VN.n10 GND 0.012255f
C85 VN.n11 GND 0.022726f
C86 VN.n12 GND 0.012255f
C87 VN.n13 GND 0.012292f
C88 VN.n14 GND 0.012255f
C89 VN.t16 GND 0.924272f
C90 VN.n15 GND 0.33942f
C91 VN.n16 GND 0.022726f
C92 VN.n17 GND 0.012255f
C93 VN.n18 GND 0.022726f
C94 VN.n19 GND 0.012255f
C95 VN.t8 GND 0.924272f
C96 VN.n20 GND 0.33942f
C97 VN.n21 GND 0.012255f
C98 VN.n22 GND 0.022726f
C99 VN.n23 GND 0.012255f
C100 VN.n24 GND 0.022499f
C101 VN.n25 GND 0.012255f
C102 VN.n26 GND 0.02037f
C103 VN.t6 GND 1.18563f
C104 VN.t13 GND 0.924272f
C105 VN.n27 GND 0.391406f
C106 VN.n28 GND 0.469716f
C107 VN.n29 GND 0.136158f
C108 VN.n30 GND 0.012255f
C109 VN.n31 GND 0.022726f
C110 VN.n32 GND 0.022726f
C111 VN.n33 GND 0.022726f
C112 VN.n34 GND 0.012255f
C113 VN.n35 GND 0.012255f
C114 VN.n36 GND 0.012255f
C115 VN.n37 GND 0.007426f
C116 VN.n38 GND 0.018608f
C117 VN.n39 GND 0.022726f
C118 VN.n40 GND 0.012255f
C119 VN.n41 GND 0.012255f
C120 VN.n42 GND 0.012255f
C121 VN.n43 GND 0.022726f
C122 VN.n44 GND 0.022726f
C123 VN.n45 GND 0.012292f
C124 VN.n46 GND 0.012255f
C125 VN.n47 GND 0.012255f
C126 VN.n48 GND 0.02194f
C127 VN.n49 GND 0.022726f
C128 VN.n50 GND 0.022726f
C129 VN.n51 GND 0.012255f
C130 VN.n52 GND 0.012255f
C131 VN.n53 GND 0.012255f
C132 VN.n54 GND 0.020696f
C133 VN.n55 GND 0.007139f
C134 VN.n56 GND 0.020696f
C135 VN.n57 GND 0.012255f
C136 VN.n58 GND 0.012255f
C137 VN.n59 GND 0.012255f
C138 VN.n60 GND 0.022726f
C139 VN.n61 GND 0.022726f
C140 VN.n62 GND 0.02194f
C141 VN.n63 GND 0.012255f
C142 VN.n64 GND 0.012255f
C143 VN.n65 GND 0.012255f
C144 VN.n66 GND 0.022726f
C145 VN.n67 GND 0.022726f
C146 VN.n68 GND 0.022726f
C147 VN.n69 GND 0.012255f
C148 VN.n70 GND 0.012255f
C149 VN.n71 GND 0.012255f
C150 VN.n72 GND 0.018608f
C151 VN.n73 GND 0.007426f
C152 VN.n74 GND 0.022499f
C153 VN.n75 GND 0.012255f
C154 VN.n76 GND 0.012255f
C155 VN.n77 GND 0.012255f
C156 VN.n78 GND 0.022726f
C157 VN.n79 GND 0.022726f
C158 VN.n80 GND 0.02037f
C159 VN.n81 GND 0.012255f
C160 VN.n82 GND 0.012255f
C161 VN.n83 GND 0.012255f
C162 VN.n84 GND 0.022726f
C163 VN.n85 GND 0.022726f
C164 VN.n86 GND 0.022726f
C165 VN.n87 GND 0.012255f
C166 VN.n88 GND 0.012255f
C167 VN.n89 GND 0.012255f
C168 VN.n90 GND 0.016315f
C169 VN.n91 GND 0.008339f
C170 VN.n92 GND 0.023878f
C171 VN.n93 GND 0.012255f
C172 VN.n94 GND 0.012255f
C173 VN.n95 GND 0.012255f
C174 VN.n96 GND 0.022726f
C175 VN.n97 GND 0.022726f
C176 VN.n98 GND 0.018799f
C177 VN.n99 GND 0.02592f
C178 VN.n100 GND 0.279693f
C179 VN.t14 GND 0.924272f
C180 VN.n101 GND 0.393886f
C181 VN.n102 GND 0.012255f
C182 VN.n103 GND 0.022726f
C183 VN.n104 GND 0.012255f
C184 VN.n105 GND 0.022726f
C185 VN.n106 GND 0.012255f
C186 VN.n107 GND 0.013863f
C187 VN.n108 GND 0.012255f
C188 VN.n109 GND 0.022726f
C189 VN.n110 GND 0.012255f
C190 VN.n111 GND 0.022726f
C191 VN.n112 GND 0.012255f
C192 VN.n113 GND 0.012292f
C193 VN.n114 GND 0.012255f
C194 VN.n115 GND 0.022726f
C195 VN.n116 GND 0.012255f
C196 VN.n117 GND 0.022726f
C197 VN.n118 GND 0.012255f
C198 VN.t7 GND 0.924272f
C199 VN.n119 GND 0.33942f
C200 VN.n120 GND 0.012255f
C201 VN.n121 GND 0.022726f
C202 VN.n122 GND 0.012255f
C203 VN.n123 GND 0.022499f
C204 VN.n124 GND 0.012255f
C205 VN.n125 GND 0.02037f
C206 VN.t9 GND 0.924272f
C207 VN.n126 GND 0.391406f
C208 VN.t17 GND 1.18563f
C209 VN.n127 GND 0.469715f
C210 VN.n128 GND 0.136158f
C211 VN.n129 GND 0.012255f
C212 VN.n130 GND 0.022726f
C213 VN.n131 GND 0.022726f
C214 VN.n132 GND 0.022726f
C215 VN.n133 GND 0.012255f
C216 VN.n134 GND 0.012255f
C217 VN.n135 GND 0.012255f
C218 VN.n136 GND 0.007426f
C219 VN.n137 GND 0.018608f
C220 VN.n138 GND 0.022726f
C221 VN.n139 GND 0.012255f
C222 VN.n140 GND 0.012255f
C223 VN.n141 GND 0.012255f
C224 VN.n142 GND 0.022726f
C225 VN.n143 GND 0.022726f
C226 VN.n144 GND 0.012292f
C227 VN.n145 GND 0.012255f
C228 VN.n146 GND 0.012255f
C229 VN.n147 GND 0.02194f
C230 VN.n148 GND 0.022726f
C231 VN.n149 GND 0.022726f
C232 VN.n150 GND 0.012255f
C233 VN.n151 GND 0.012255f
C234 VN.n152 GND 0.012255f
C235 VN.n153 GND 0.020696f
C236 VN.n154 GND 0.007139f
C237 VN.n155 GND 0.020696f
C238 VN.n156 GND 0.012255f
C239 VN.n157 GND 0.012255f
C240 VN.n158 GND 0.012255f
C241 VN.n159 GND 0.022726f
C242 VN.n160 GND 0.022726f
C243 VN.t12 GND 0.924272f
C244 VN.n161 GND 0.33942f
C245 VN.n162 GND 0.02194f
C246 VN.n163 GND 0.012255f
C247 VN.n164 GND 0.012255f
C248 VN.n165 GND 0.012255f
C249 VN.n166 GND 0.022726f
C250 VN.n167 GND 0.022726f
C251 VN.n168 GND 0.022726f
C252 VN.n169 GND 0.012255f
C253 VN.n170 GND 0.012255f
C254 VN.n171 GND 0.012255f
C255 VN.n172 GND 0.018608f
C256 VN.n173 GND 0.007426f
C257 VN.n174 GND 0.022499f
C258 VN.n175 GND 0.012255f
C259 VN.n176 GND 0.012255f
C260 VN.n177 GND 0.012255f
C261 VN.n178 GND 0.022726f
C262 VN.n179 GND 0.022726f
C263 VN.t15 GND 0.924272f
C264 VN.n180 GND 0.33942f
C265 VN.n181 GND 0.02037f
C266 VN.n182 GND 0.012255f
C267 VN.n183 GND 0.012255f
C268 VN.n184 GND 0.012255f
C269 VN.n185 GND 0.022726f
C270 VN.n186 GND 0.022726f
C271 VN.n187 GND 0.022726f
C272 VN.n188 GND 0.012255f
C273 VN.n189 GND 0.012255f
C274 VN.n190 GND 0.012255f
C275 VN.n191 GND 0.016315f
C276 VN.n192 GND 0.008339f
C277 VN.n193 GND 0.023878f
C278 VN.n194 GND 0.012255f
C279 VN.n195 GND 0.012255f
C280 VN.n196 GND 0.012255f
C281 VN.n197 GND 0.022726f
C282 VN.n198 GND 0.022726f
C283 VN.n199 GND 0.018799f
C284 VN.n200 GND 0.02592f
C285 VN.n201 GND 0.943104f
C286 VN.n202 GND 1.12834f
C287 VN.t3 GND 0.021156f
C288 VN.t4 GND 0.003778f
C289 VN.t0 GND 0.003778f
C290 VN.n203 GND 0.012252f
C291 VN.n204 GND 0.095115f
C292 VN.t5 GND 0.003778f
C293 VN.t2 GND 0.003778f
C294 VN.n205 GND 0.012252f
C295 VN.n206 GND 0.051406f
C296 VN.t1 GND 0.021027f
C297 VN.n207 GND 0.063709f
C298 VN.n208 GND 4.03065f
C299 a_n7336_n129.n0 GND 1.69787f
C300 a_n7336_n129.n1 GND 1.69787f
C301 a_n7336_n129.t17 GND 0.089858f
C302 a_n7336_n129.t9 GND 0.682781f
C303 a_n7336_n129.n2 GND 1.62055f
C304 a_n7336_n129.t27 GND 0.905428f
C305 a_n7336_n129.n3 GND 4.1434f
C306 a_n7336_n129.t7 GND 0.905428f
C307 a_n7336_n129.n4 GND 1.46162f
C308 a_n7336_n129.t8 GND 0.905428f
C309 a_n7336_n129.n5 GND 1.46162f
C310 a_n7336_n129.t26 GND 0.905428f
C311 a_n7336_n129.n6 GND 3.56946f
C312 a_n7336_n129.n7 GND 1.611f
C313 a_n7336_n129.t22 GND 0.68278f
C314 a_n7336_n129.n8 GND 1.4466f
C315 a_n7336_n129.t1 GND 0.089858f
C316 a_n7336_n129.t6 GND 0.089858f
C317 a_n7336_n129.n9 GND 0.566236f
C318 a_n7336_n129.n10 GND 1.20772f
C319 a_n7336_n129.t21 GND 0.089858f
C320 a_n7336_n129.t24 GND 0.089858f
C321 a_n7336_n129.n11 GND 0.566236f
C322 a_n7336_n129.n12 GND 1.20772f
C323 a_n7336_n129.t2 GND 0.68278f
C324 a_n7336_n129.t12 GND 0.68278f
C325 a_n7336_n129.t18 GND 0.089858f
C326 a_n7336_n129.t11 GND 0.089858f
C327 a_n7336_n129.n13 GND 0.566236f
C328 a_n7336_n129.n14 GND 1.20772f
C329 a_n7336_n129.t16 GND 0.089858f
C330 a_n7336_n129.t14 GND 0.089858f
C331 a_n7336_n129.n15 GND 0.566236f
C332 a_n7336_n129.n16 GND 1.20772f
C333 a_n7336_n129.t15 GND 0.68278f
C334 a_n7336_n129.n17 GND 1.4466f
C335 a_n7336_n129.n18 GND 2.00949f
C336 a_n7336_n129.t5 GND 0.682777f
C337 a_n7336_n129.n19 GND 1.62055f
C338 a_n7336_n129.t0 GND 0.089858f
C339 a_n7336_n129.t3 GND 0.089858f
C340 a_n7336_n129.n20 GND 0.566238f
C341 a_n7336_n129.n21 GND 1.20772f
C342 a_n7336_n129.t25 GND 0.089858f
C343 a_n7336_n129.t4 GND 0.089858f
C344 a_n7336_n129.n22 GND 0.566238f
C345 a_n7336_n129.n23 GND 1.20772f
C346 a_n7336_n129.t23 GND 0.682781f
C347 a_n7336_n129.t13 GND 0.682781f
C348 a_n7336_n129.t10 GND 0.089858f
C349 a_n7336_n129.t19 GND 0.089858f
C350 a_n7336_n129.n24 GND 0.566238f
C351 a_n7336_n129.n25 GND 1.20772f
C352 a_n7336_n129.n26 GND 1.20772f
C353 a_n7336_n129.n27 GND 0.566238f
C354 a_n7336_n129.t20 GND 0.089858f
C355 VP.t11 GND 1.27568f
C356 VP.n0 GND 0.54364f
C357 VP.n1 GND 0.016914f
C358 VP.n2 GND 0.031366f
C359 VP.n3 GND 0.016914f
C360 VP.n4 GND 0.031366f
C361 VP.n5 GND 0.016914f
C362 VP.n6 GND 0.019133f
C363 VP.n7 GND 0.016914f
C364 VP.n8 GND 0.031366f
C365 VP.n9 GND 0.016914f
C366 VP.n10 GND 0.031366f
C367 VP.n11 GND 0.016914f
C368 VP.n12 GND 0.016965f
C369 VP.n13 GND 0.016914f
C370 VP.n14 GND 0.031366f
C371 VP.n15 GND 0.016914f
C372 VP.n16 GND 0.031366f
C373 VP.n17 GND 0.016914f
C374 VP.t15 GND 1.27568f
C375 VP.n18 GND 0.468466f
C376 VP.n19 GND 0.016914f
C377 VP.n20 GND 0.031366f
C378 VP.n21 GND 0.016914f
C379 VP.n22 GND 0.031052f
C380 VP.n23 GND 0.016914f
C381 VP.n24 GND 0.028114f
C382 VP.t8 GND 1.27568f
C383 VP.n25 GND 0.540218f
C384 VP.t14 GND 1.6364f
C385 VP.n26 GND 0.648299f
C386 VP.n27 GND 0.187925f
C387 VP.n28 GND 0.016914f
C388 VP.n29 GND 0.031366f
C389 VP.n30 GND 0.031366f
C390 VP.n31 GND 0.031366f
C391 VP.n32 GND 0.016914f
C392 VP.n33 GND 0.016914f
C393 VP.n34 GND 0.016914f
C394 VP.n35 GND 0.010249f
C395 VP.n36 GND 0.025682f
C396 VP.n37 GND 0.031366f
C397 VP.n38 GND 0.016914f
C398 VP.n39 GND 0.016914f
C399 VP.n40 GND 0.016914f
C400 VP.n41 GND 0.031366f
C401 VP.n42 GND 0.031366f
C402 VP.n43 GND 0.016965f
C403 VP.n44 GND 0.016914f
C404 VP.n45 GND 0.016914f
C405 VP.n46 GND 0.030282f
C406 VP.n47 GND 0.031366f
C407 VP.n48 GND 0.031366f
C408 VP.n49 GND 0.016914f
C409 VP.n50 GND 0.016914f
C410 VP.n51 GND 0.016914f
C411 VP.n52 GND 0.028565f
C412 VP.n53 GND 0.009853f
C413 VP.n54 GND 0.028565f
C414 VP.n55 GND 0.016914f
C415 VP.n56 GND 0.016914f
C416 VP.n57 GND 0.016914f
C417 VP.n58 GND 0.031366f
C418 VP.n59 GND 0.031366f
C419 VP.t10 GND 1.27568f
C420 VP.n60 GND 0.468466f
C421 VP.n61 GND 0.030282f
C422 VP.n62 GND 0.016914f
C423 VP.n63 GND 0.016914f
C424 VP.n64 GND 0.016914f
C425 VP.n65 GND 0.031366f
C426 VP.n66 GND 0.031366f
C427 VP.n67 GND 0.031366f
C428 VP.n68 GND 0.016914f
C429 VP.n69 GND 0.016914f
C430 VP.n70 GND 0.016914f
C431 VP.n71 GND 0.025682f
C432 VP.n72 GND 0.010249f
C433 VP.n73 GND 0.031052f
C434 VP.n74 GND 0.016914f
C435 VP.n75 GND 0.016914f
C436 VP.n76 GND 0.016914f
C437 VP.n77 GND 0.031366f
C438 VP.n78 GND 0.031366f
C439 VP.t12 GND 1.27568f
C440 VP.n79 GND 0.468466f
C441 VP.n80 GND 0.028114f
C442 VP.n81 GND 0.016914f
C443 VP.n82 GND 0.016914f
C444 VP.n83 GND 0.016914f
C445 VP.n84 GND 0.031366f
C446 VP.n85 GND 0.031366f
C447 VP.n86 GND 0.031366f
C448 VP.n87 GND 0.016914f
C449 VP.n88 GND 0.016914f
C450 VP.n89 GND 0.016914f
C451 VP.n90 GND 0.022518f
C452 VP.n91 GND 0.011509f
C453 VP.n92 GND 0.032957f
C454 VP.n93 GND 0.016914f
C455 VP.n94 GND 0.016914f
C456 VP.n95 GND 0.016914f
C457 VP.n96 GND 0.031366f
C458 VP.n97 GND 0.031366f
C459 VP.n98 GND 0.025946f
C460 VP.n99 GND 0.035775f
C461 VP.n100 GND 0.39022f
C462 VP.t17 GND 1.27568f
C463 VP.n101 GND 0.54364f
C464 VP.n102 GND 0.016914f
C465 VP.n103 GND 0.031366f
C466 VP.n104 GND 0.016914f
C467 VP.n105 GND 0.031366f
C468 VP.n106 GND 0.016914f
C469 VP.n107 GND 0.019133f
C470 VP.n108 GND 0.016914f
C471 VP.t6 GND 1.27568f
C472 VP.n109 GND 0.468466f
C473 VP.n110 GND 0.031366f
C474 VP.n111 GND 0.016914f
C475 VP.n112 GND 0.031366f
C476 VP.n113 GND 0.016914f
C477 VP.n114 GND 0.016965f
C478 VP.n115 GND 0.016914f
C479 VP.t9 GND 1.27568f
C480 VP.n116 GND 0.468466f
C481 VP.n117 GND 0.031366f
C482 VP.n118 GND 0.016914f
C483 VP.n119 GND 0.031366f
C484 VP.n120 GND 0.016914f
C485 VP.t16 GND 1.27568f
C486 VP.n121 GND 0.468466f
C487 VP.n122 GND 0.016914f
C488 VP.n123 GND 0.031366f
C489 VP.n124 GND 0.016914f
C490 VP.n125 GND 0.031052f
C491 VP.n126 GND 0.016914f
C492 VP.n127 GND 0.028114f
C493 VP.t13 GND 1.6364f
C494 VP.t7 GND 1.27568f
C495 VP.n128 GND 0.540218f
C496 VP.n129 GND 0.6483f
C497 VP.n130 GND 0.187925f
C498 VP.n131 GND 0.016914f
C499 VP.n132 GND 0.031366f
C500 VP.n133 GND 0.031366f
C501 VP.n134 GND 0.031366f
C502 VP.n135 GND 0.016914f
C503 VP.n136 GND 0.016914f
C504 VP.n137 GND 0.016914f
C505 VP.n138 GND 0.010249f
C506 VP.n139 GND 0.025682f
C507 VP.n140 GND 0.031366f
C508 VP.n141 GND 0.016914f
C509 VP.n142 GND 0.016914f
C510 VP.n143 GND 0.016914f
C511 VP.n144 GND 0.031366f
C512 VP.n145 GND 0.031366f
C513 VP.n146 GND 0.016965f
C514 VP.n147 GND 0.016914f
C515 VP.n148 GND 0.016914f
C516 VP.n149 GND 0.030282f
C517 VP.n150 GND 0.031366f
C518 VP.n151 GND 0.031366f
C519 VP.n152 GND 0.016914f
C520 VP.n153 GND 0.016914f
C521 VP.n154 GND 0.016914f
C522 VP.n155 GND 0.028565f
C523 VP.n156 GND 0.009853f
C524 VP.n157 GND 0.028565f
C525 VP.n158 GND 0.016914f
C526 VP.n159 GND 0.016914f
C527 VP.n160 GND 0.016914f
C528 VP.n161 GND 0.031366f
C529 VP.n162 GND 0.031366f
C530 VP.n163 GND 0.030282f
C531 VP.n164 GND 0.016914f
C532 VP.n165 GND 0.016914f
C533 VP.n166 GND 0.016914f
C534 VP.n167 GND 0.031366f
C535 VP.n168 GND 0.031366f
C536 VP.n169 GND 0.031366f
C537 VP.n170 GND 0.016914f
C538 VP.n171 GND 0.016914f
C539 VP.n172 GND 0.016914f
C540 VP.n173 GND 0.025682f
C541 VP.n174 GND 0.010249f
C542 VP.n175 GND 0.031052f
C543 VP.n176 GND 0.016914f
C544 VP.n177 GND 0.016914f
C545 VP.n178 GND 0.016914f
C546 VP.n179 GND 0.031366f
C547 VP.n180 GND 0.031366f
C548 VP.n181 GND 0.028114f
C549 VP.n182 GND 0.016914f
C550 VP.n183 GND 0.016914f
C551 VP.n184 GND 0.016914f
C552 VP.n185 GND 0.031366f
C553 VP.n186 GND 0.031366f
C554 VP.n187 GND 0.031366f
C555 VP.n188 GND 0.016914f
C556 VP.n189 GND 0.016914f
C557 VP.n190 GND 0.016914f
C558 VP.n191 GND 0.022518f
C559 VP.n192 GND 0.011509f
C560 VP.n193 GND 0.032957f
C561 VP.n194 GND 0.016914f
C562 VP.n195 GND 0.016914f
C563 VP.n196 GND 0.016914f
C564 VP.n197 GND 0.031366f
C565 VP.n198 GND 0.031366f
C566 VP.n199 GND 0.025946f
C567 VP.n200 GND 0.035775f
C568 VP.n201 GND 1.3082f
C569 VP.n202 GND 1.56445f
C570 VP.t0 GND 0.029199f
C571 VP.t5 GND 0.005214f
C572 VP.t1 GND 0.005214f
C573 VP.n203 GND 0.01691f
C574 VP.n204 GND 0.131277f
C575 VP.t4 GND 0.005214f
C576 VP.t2 GND 0.005214f
C577 VP.n205 GND 0.01691f
C578 VP.n206 GND 0.07095f
C579 VP.t3 GND 0.029021f
C580 VP.n207 GND 0.078756f
C581 VP.n208 GND 1.84514f
C582 VOUT.t82 GND 0.045214f
C583 VOUT.t85 GND 0.045214f
C584 VOUT.n0 GND 0.256126f
C585 VOUT.t108 GND 0.045214f
C586 VOUT.t109 GND 0.045214f
C587 VOUT.n1 GND 0.242959f
C588 VOUT.n2 GND 1.49185f
C589 VOUT.t94 GND 0.045214f
C590 VOUT.t107 GND 0.045214f
C591 VOUT.n3 GND 0.242959f
C592 VOUT.n4 GND 0.867394f
C593 VOUT.t83 GND 0.045214f
C594 VOUT.t92 GND 0.045214f
C595 VOUT.n5 GND 0.256126f
C596 VOUT.t105 GND 0.045214f
C597 VOUT.t115 GND 0.045214f
C598 VOUT.n6 GND 0.242959f
C599 VOUT.n7 GND 1.49185f
C600 VOUT.t96 GND 0.045214f
C601 VOUT.t91 GND 0.045214f
C602 VOUT.n8 GND 0.242959f
C603 VOUT.n9 GND 0.822833f
C604 VOUT.n10 GND 0.660834f
C605 VOUT.t84 GND 0.045214f
C606 VOUT.t93 GND 0.045214f
C607 VOUT.n11 GND 0.256126f
C608 VOUT.t103 GND 0.045214f
C609 VOUT.t114 GND 0.045214f
C610 VOUT.n12 GND 0.242959f
C611 VOUT.n13 GND 1.49185f
C612 VOUT.t95 GND 0.045214f
C613 VOUT.t89 GND 0.045214f
C614 VOUT.n14 GND 0.242959f
C615 VOUT.n15 GND 0.822833f
C616 VOUT.n16 GND 0.734024f
C617 VOUT.n17 GND 10.3095f
C618 VOUT.n18 GND 4.82392f
C619 VOUT.n19 GND 3.8282f
C620 VOUT.n20 GND 3.8282f
C621 VOUT.t122 GND 12.836401f
C622 VOUT.t118 GND 11.7599f
C623 VOUT.t121 GND 11.7599f
C624 VOUT.t123 GND 13.0908f
C625 VOUT.n21 GND 9.19657f
C626 VOUT.n22 GND 4.54901f
C627 VOUT.n23 GND 3.8282f
C628 VOUT.n24 GND 3.8232f
C629 VOUT.n25 GND 4.3338f
C630 VOUT.n26 GND 3.8282f
C631 VOUT.n27 GND 4.29575f
C632 VOUT.n28 GND 9.74233f
C633 VOUT.t120 GND 12.836401f
C634 VOUT.n29 GND 11.5029f
C635 VOUT.n30 GND 4.11597f
C636 VOUT.t116 GND 11.7599f
C637 VOUT.n31 GND 4.3338f
C638 VOUT.n32 GND 3.8232f
C639 VOUT.t117 GND 11.7599f
C640 VOUT.n33 GND 4.3338f
C641 VOUT.n34 GND 3.8232f
C642 VOUT.t119 GND 11.7599f
C643 VOUT.n35 GND 5.7609f
C644 VOUT.n36 GND 1.9557f
C645 VOUT.t87 GND 0.045214f
C646 VOUT.t86 GND 0.045214f
C647 VOUT.n37 GND 0.256126f
C648 VOUT.t102 GND 0.045214f
C649 VOUT.t101 GND 0.045214f
C650 VOUT.n38 GND 0.242959f
C651 VOUT.n39 GND 1.49185f
C652 VOUT.t100 GND 0.045214f
C653 VOUT.t99 GND 0.045214f
C654 VOUT.n40 GND 0.242959f
C655 VOUT.n41 GND 0.867394f
C656 VOUT.t111 GND 0.045214f
C657 VOUT.t98 GND 0.045214f
C658 VOUT.n42 GND 0.256126f
C659 VOUT.t106 GND 0.045214f
C660 VOUT.t88 GND 0.045214f
C661 VOUT.n43 GND 0.242959f
C662 VOUT.n44 GND 1.49185f
C663 VOUT.t80 GND 0.045214f
C664 VOUT.t112 GND 0.045214f
C665 VOUT.n45 GND 0.242959f
C666 VOUT.n46 GND 0.822833f
C667 VOUT.n47 GND 0.660834f
C668 VOUT.t110 GND 0.045214f
C669 VOUT.t97 GND 0.045214f
C670 VOUT.n48 GND 0.256126f
C671 VOUT.t104 GND 0.045214f
C672 VOUT.t90 GND 0.045214f
C673 VOUT.n49 GND 0.242959f
C674 VOUT.n50 GND 1.49185f
C675 VOUT.t81 GND 0.045214f
C676 VOUT.t113 GND 0.045214f
C677 VOUT.n51 GND 0.242958f
C678 VOUT.n52 GND 0.822834f
C679 VOUT.n53 GND 0.734024f
C680 VOUT.n54 GND 12.4979f
C681 VOUT.t30 GND 0.025956f
C682 VOUT.t49 GND 0.025956f
C683 VOUT.n55 GND 0.182203f
C684 VOUT.t5 GND 0.025956f
C685 VOUT.t20 GND 0.025956f
C686 VOUT.n56 GND 0.16846f
C687 VOUT.n57 GND 1.30028f
C688 VOUT.t4 GND 0.025956f
C689 VOUT.t53 GND 0.025956f
C690 VOUT.n58 GND 0.16846f
C691 VOUT.n59 GND 0.653454f
C692 VOUT.t17 GND 0.025956f
C693 VOUT.t23 GND 0.025956f
C694 VOUT.n60 GND 0.16846f
C695 VOUT.n61 GND 0.757185f
C696 VOUT.t10 GND 0.025956f
C697 VOUT.t76 GND 0.025956f
C698 VOUT.n62 GND 0.182203f
C699 VOUT.t11 GND 0.025956f
C700 VOUT.t9 GND 0.025956f
C701 VOUT.n63 GND 0.16846f
C702 VOUT.n64 GND 1.30028f
C703 VOUT.t16 GND 0.025956f
C704 VOUT.t59 GND 0.025956f
C705 VOUT.n65 GND 0.16846f
C706 VOUT.n66 GND 0.653454f
C707 VOUT.t34 GND 0.025956f
C708 VOUT.t45 GND 0.025956f
C709 VOUT.n67 GND 0.16846f
C710 VOUT.n68 GND 0.729257f
C711 VOUT.n69 GND 0.521685f
C712 VOUT.t27 GND 0.025956f
C713 VOUT.t25 GND 0.025956f
C714 VOUT.n70 GND 0.182203f
C715 VOUT.t66 GND 0.025956f
C716 VOUT.t75 GND 0.025956f
C717 VOUT.n71 GND 0.16846f
C718 VOUT.n72 GND 1.30028f
C719 VOUT.t71 GND 0.025956f
C720 VOUT.t3 GND 0.025956f
C721 VOUT.n73 GND 0.16846f
C722 VOUT.n74 GND 0.653454f
C723 VOUT.t51 GND 0.025956f
C724 VOUT.t13 GND 0.025956f
C725 VOUT.n75 GND 0.16846f
C726 VOUT.n76 GND 0.729257f
C727 VOUT.n77 GND 0.345811f
C728 VOUT.t29 GND 0.025956f
C729 VOUT.t6 GND 0.025956f
C730 VOUT.n78 GND 0.182203f
C731 VOUT.t77 GND 0.025956f
C732 VOUT.t62 GND 0.025956f
C733 VOUT.n79 GND 0.16846f
C734 VOUT.n80 GND 1.30028f
C735 VOUT.t67 GND 0.025956f
C736 VOUT.t73 GND 0.025956f
C737 VOUT.n81 GND 0.16846f
C738 VOUT.n82 GND 0.653454f
C739 VOUT.t60 GND 0.025956f
C740 VOUT.t24 GND 0.025956f
C741 VOUT.n83 GND 0.16846f
C742 VOUT.n84 GND 0.729257f
C743 VOUT.n85 GND 0.345811f
C744 VOUT.t74 GND 0.025956f
C745 VOUT.t56 GND 0.025956f
C746 VOUT.n86 GND 0.182203f
C747 VOUT.t36 GND 0.025956f
C748 VOUT.t37 GND 0.025956f
C749 VOUT.n87 GND 0.16846f
C750 VOUT.n88 GND 1.30028f
C751 VOUT.t41 GND 0.025956f
C752 VOUT.t31 GND 0.025956f
C753 VOUT.n89 GND 0.16846f
C754 VOUT.n90 GND 0.653454f
C755 VOUT.t8 GND 0.025956f
C756 VOUT.t72 GND 0.025956f
C757 VOUT.n91 GND 0.16846f
C758 VOUT.n92 GND 0.729257f
C759 VOUT.n93 GND 0.536437f
C760 VOUT.n94 GND 12.665f
C761 VOUT.t39 GND 0.025956f
C762 VOUT.t70 GND 0.025956f
C763 VOUT.n95 GND 0.182203f
C764 VOUT.t58 GND 0.025956f
C765 VOUT.t50 GND 0.025956f
C766 VOUT.n96 GND 0.16846f
C767 VOUT.n97 GND 1.30028f
C768 VOUT.t47 GND 0.025956f
C769 VOUT.t26 GND 0.025956f
C770 VOUT.n98 GND 0.16846f
C771 VOUT.n99 GND 0.653454f
C772 VOUT.t46 GND 0.025956f
C773 VOUT.t57 GND 0.025956f
C774 VOUT.n100 GND 0.16846f
C775 VOUT.n101 GND 0.757185f
C776 VOUT.t0 GND 0.025956f
C777 VOUT.t7 GND 0.025956f
C778 VOUT.n102 GND 0.182203f
C779 VOUT.t52 GND 0.025956f
C780 VOUT.t69 GND 0.025956f
C781 VOUT.n103 GND 0.16846f
C782 VOUT.n104 GND 1.30028f
C783 VOUT.t12 GND 0.025956f
C784 VOUT.t22 GND 0.025956f
C785 VOUT.n105 GND 0.16846f
C786 VOUT.n106 GND 0.653454f
C787 VOUT.t18 GND 0.025956f
C788 VOUT.t14 GND 0.025956f
C789 VOUT.n107 GND 0.16846f
C790 VOUT.n108 GND 0.729257f
C791 VOUT.n109 GND 0.521685f
C792 VOUT.t64 GND 0.025956f
C793 VOUT.t55 GND 0.025956f
C794 VOUT.n110 GND 0.182203f
C795 VOUT.t44 GND 0.025956f
C796 VOUT.t48 GND 0.025956f
C797 VOUT.n111 GND 0.16846f
C798 VOUT.n112 GND 1.30028f
C799 VOUT.t28 GND 0.025956f
C800 VOUT.t33 GND 0.025956f
C801 VOUT.n113 GND 0.16846f
C802 VOUT.n114 GND 0.653454f
C803 VOUT.t61 GND 0.025956f
C804 VOUT.t21 GND 0.025956f
C805 VOUT.n115 GND 0.16846f
C806 VOUT.n116 GND 0.729257f
C807 VOUT.n117 GND 0.345811f
C808 VOUT.t35 GND 0.025956f
C809 VOUT.t32 GND 0.025956f
C810 VOUT.n118 GND 0.182203f
C811 VOUT.t2 GND 0.025956f
C812 VOUT.t1 GND 0.025956f
C813 VOUT.n119 GND 0.16846f
C814 VOUT.n120 GND 1.30028f
C815 VOUT.t78 GND 0.025956f
C816 VOUT.t54 GND 0.025956f
C817 VOUT.n121 GND 0.16846f
C818 VOUT.n122 GND 0.653454f
C819 VOUT.t68 GND 0.025956f
C820 VOUT.t63 GND 0.025956f
C821 VOUT.n123 GND 0.16846f
C822 VOUT.n124 GND 0.729257f
C823 VOUT.n125 GND 0.345811f
C824 VOUT.t65 GND 0.025956f
C825 VOUT.t79 GND 0.025956f
C826 VOUT.n126 GND 0.182203f
C827 VOUT.t19 GND 0.025956f
C828 VOUT.t15 GND 0.025956f
C829 VOUT.n127 GND 0.16846f
C830 VOUT.n128 GND 1.30028f
C831 VOUT.t38 GND 0.025956f
C832 VOUT.t43 GND 0.025956f
C833 VOUT.n129 GND 0.16846f
C834 VOUT.n130 GND 0.653454f
C835 VOUT.t42 GND 0.025956f
C836 VOUT.t40 GND 0.025956f
C837 VOUT.n131 GND 0.16846f
C838 VOUT.n132 GND 0.729257f
C839 VOUT.n133 GND 0.536437f
C840 VOUT.n134 GND 9.66788f
C841 VOUT.n135 GND 5.31068f
C842 CS_BIAS.t55 GND 0.226601f
C843 CS_BIAS.n0 GND 0.122067f
C844 CS_BIAS.n1 GND 0.006543f
C845 CS_BIAS.n2 GND 0.012195f
C846 CS_BIAS.n3 GND 0.006543f
C847 CS_BIAS.n4 GND 0.012195f
C848 CS_BIAS.n5 GND 0.006543f
C849 CS_BIAS.t35 GND 0.226601f
C850 CS_BIAS.n6 GND 0.091803f
C851 CS_BIAS.n7 GND 0.006543f
C852 CS_BIAS.n8 GND 0.012195f
C853 CS_BIAS.n9 GND 0.006543f
C854 CS_BIAS.n10 GND 0.012195f
C855 CS_BIAS.n11 GND 0.006543f
C856 CS_BIAS.t103 GND 0.226601f
C857 CS_BIAS.n12 GND 0.091803f
C858 CS_BIAS.n13 GND 0.006543f
C859 CS_BIAS.n14 GND 0.012195f
C860 CS_BIAS.n15 GND 0.006543f
C861 CS_BIAS.n16 GND 0.013142f
C862 CS_BIAS.n17 GND 0.006543f
C863 CS_BIAS.n18 GND 0.008041f
C864 CS_BIAS.n19 GND 0.006543f
C865 CS_BIAS.t64 GND 0.226601f
C866 CS_BIAS.n20 GND 0.091803f
C867 CS_BIAS.n21 GND 0.012195f
C868 CS_BIAS.t0 GND 0.226601f
C869 CS_BIAS.n22 GND 0.122067f
C870 CS_BIAS.n23 GND 0.006543f
C871 CS_BIAS.n24 GND 0.012195f
C872 CS_BIAS.n25 GND 0.006543f
C873 CS_BIAS.n26 GND 0.012195f
C874 CS_BIAS.n27 GND 0.006543f
C875 CS_BIAS.t26 GND 0.226601f
C876 CS_BIAS.n28 GND 0.091803f
C877 CS_BIAS.n29 GND 0.006543f
C878 CS_BIAS.n30 GND 0.012195f
C879 CS_BIAS.n31 GND 0.006543f
C880 CS_BIAS.n32 GND 0.012195f
C881 CS_BIAS.n33 GND 0.006543f
C882 CS_BIAS.t22 GND 0.226601f
C883 CS_BIAS.n34 GND 0.091803f
C884 CS_BIAS.n35 GND 0.006543f
C885 CS_BIAS.n36 GND 0.012195f
C886 CS_BIAS.n37 GND 0.006543f
C887 CS_BIAS.n38 GND 0.013142f
C888 CS_BIAS.n39 GND 0.006543f
C889 CS_BIAS.n40 GND 0.008041f
C890 CS_BIAS.n41 GND 0.006543f
C891 CS_BIAS.t16 GND 0.226601f
C892 CS_BIAS.n42 GND 0.091803f
C893 CS_BIAS.n43 GND 0.012195f
C894 CS_BIAS.n44 GND 0.006543f
C895 CS_BIAS.n45 GND 0.012195f
C896 CS_BIAS.n46 GND 0.006543f
C897 CS_BIAS.t20 GND 0.226601f
C898 CS_BIAS.n47 GND 0.091803f
C899 CS_BIAS.n48 GND 0.006543f
C900 CS_BIAS.n49 GND 0.012195f
C901 CS_BIAS.n50 GND 0.006543f
C902 CS_BIAS.n51 GND 0.012603f
C903 CS_BIAS.n52 GND 0.006543f
C904 CS_BIAS.n53 GND 0.006596f
C905 CS_BIAS.n54 GND 0.006543f
C906 CS_BIAS.t8 GND 0.226601f
C907 CS_BIAS.n55 GND 0.091803f
C908 CS_BIAS.n56 GND 0.012195f
C909 CS_BIAS.n57 GND 0.006543f
C910 CS_BIAS.n58 GND 0.012195f
C911 CS_BIAS.n59 GND 0.006543f
C912 CS_BIAS.t14 GND 0.226601f
C913 CS_BIAS.n60 GND 0.117336f
C914 CS_BIAS.t18 GND 0.334543f
C915 CS_BIAS.n61 GND 0.172166f
C916 CS_BIAS.n62 GND 0.079011f
C917 CS_BIAS.n63 GND 0.008884f
C918 CS_BIAS.n64 GND 0.012195f
C919 CS_BIAS.n65 GND 0.012195f
C920 CS_BIAS.n66 GND 0.006543f
C921 CS_BIAS.n67 GND 0.006543f
C922 CS_BIAS.n68 GND 0.006543f
C923 CS_BIAS.n69 GND 0.012633f
C924 CS_BIAS.n70 GND 0.004276f
C925 CS_BIAS.n71 GND 0.009107f
C926 CS_BIAS.n72 GND 0.006543f
C927 CS_BIAS.n73 GND 0.006543f
C928 CS_BIAS.n74 GND 0.006543f
C929 CS_BIAS.n75 GND 0.012195f
C930 CS_BIAS.n76 GND 0.012195f
C931 CS_BIAS.n77 GND 0.011774f
C932 CS_BIAS.n78 GND 0.006543f
C933 CS_BIAS.n79 GND 0.006543f
C934 CS_BIAS.n80 GND 0.006543f
C935 CS_BIAS.n81 GND 0.012195f
C936 CS_BIAS.n82 GND 0.012195f
C937 CS_BIAS.n83 GND 0.012195f
C938 CS_BIAS.n84 GND 0.006543f
C939 CS_BIAS.n85 GND 0.006543f
C940 CS_BIAS.n86 GND 0.006543f
C941 CS_BIAS.n87 GND 0.007464f
C942 CS_BIAS.n88 GND 0.005003f
C943 CS_BIAS.n89 GND 0.013142f
C944 CS_BIAS.n90 GND 0.006543f
C945 CS_BIAS.n91 GND 0.006543f
C946 CS_BIAS.n92 GND 0.006543f
C947 CS_BIAS.n93 GND 0.012195f
C948 CS_BIAS.n94 GND 0.012195f
C949 CS_BIAS.n95 GND 0.008041f
C950 CS_BIAS.n96 GND 0.006543f
C951 CS_BIAS.n97 GND 0.006543f
C952 CS_BIAS.n98 GND 0.010328f
C953 CS_BIAS.n99 GND 0.012195f
C954 CS_BIAS.n100 GND 0.012195f
C955 CS_BIAS.n101 GND 0.006543f
C956 CS_BIAS.n102 GND 0.006543f
C957 CS_BIAS.n103 GND 0.006543f
C958 CS_BIAS.n104 GND 0.011103f
C959 CS_BIAS.n105 GND 0.003811f
C960 CS_BIAS.n106 GND 0.011103f
C961 CS_BIAS.n107 GND 0.006543f
C962 CS_BIAS.n108 GND 0.006543f
C963 CS_BIAS.n109 GND 0.006543f
C964 CS_BIAS.n110 GND 0.012195f
C965 CS_BIAS.n111 GND 0.012195f
C966 CS_BIAS.n112 GND 0.010328f
C967 CS_BIAS.n113 GND 0.006543f
C968 CS_BIAS.n114 GND 0.006543f
C969 CS_BIAS.n115 GND 0.006543f
C970 CS_BIAS.n116 GND 0.012195f
C971 CS_BIAS.n117 GND 0.012195f
C972 CS_BIAS.n118 GND 0.012195f
C973 CS_BIAS.n119 GND 0.006543f
C974 CS_BIAS.n120 GND 0.006543f
C975 CS_BIAS.n121 GND 0.006543f
C976 CS_BIAS.n122 GND 0.005003f
C977 CS_BIAS.n123 GND 0.007464f
C978 CS_BIAS.n124 GND 0.012603f
C979 CS_BIAS.n125 GND 0.006543f
C980 CS_BIAS.n126 GND 0.006543f
C981 CS_BIAS.n127 GND 0.006543f
C982 CS_BIAS.n128 GND 0.012195f
C983 CS_BIAS.n129 GND 0.012195f
C984 CS_BIAS.n130 GND 0.006596f
C985 CS_BIAS.n131 GND 0.006543f
C986 CS_BIAS.n132 GND 0.006543f
C987 CS_BIAS.n133 GND 0.011774f
C988 CS_BIAS.n134 GND 0.012195f
C989 CS_BIAS.n135 GND 0.012195f
C990 CS_BIAS.n136 GND 0.006543f
C991 CS_BIAS.n137 GND 0.006543f
C992 CS_BIAS.n138 GND 0.006543f
C993 CS_BIAS.n139 GND 0.009107f
C994 CS_BIAS.n140 GND 0.004276f
C995 CS_BIAS.n141 GND 0.012633f
C996 CS_BIAS.n142 GND 0.006543f
C997 CS_BIAS.n143 GND 0.006543f
C998 CS_BIAS.n144 GND 0.006543f
C999 CS_BIAS.n145 GND 0.012195f
C1000 CS_BIAS.n146 GND 0.012195f
C1001 CS_BIAS.n147 GND 0.008884f
C1002 CS_BIAS.n148 GND 0.006543f
C1003 CS_BIAS.n149 GND 0.006543f
C1004 CS_BIAS.n150 GND 0.009486f
C1005 CS_BIAS.n151 GND 0.012195f
C1006 CS_BIAS.n152 GND 0.012195f
C1007 CS_BIAS.n153 GND 0.006543f
C1008 CS_BIAS.n154 GND 0.006543f
C1009 CS_BIAS.n155 GND 0.006543f
C1010 CS_BIAS.n156 GND 0.012073f
C1011 CS_BIAS.n157 GND 0.003964f
C1012 CS_BIAS.n158 GND 0.009979f
C1013 CS_BIAS.n159 GND 0.006543f
C1014 CS_BIAS.n160 GND 0.006543f
C1015 CS_BIAS.n161 GND 0.006543f
C1016 CS_BIAS.n162 GND 0.012195f
C1017 CS_BIAS.n163 GND 0.012195f
C1018 CS_BIAS.n164 GND 0.011172f
C1019 CS_BIAS.n165 GND 0.013846f
C1020 CS_BIAS.n166 GND 0.107996f
C1021 CS_BIAS.t1 GND 0.011256f
C1022 CS_BIAS.t27 GND 0.011256f
C1023 CS_BIAS.n167 GND 0.073052f
C1024 CS_BIAS.n168 GND 0.321859f
C1025 CS_BIAS.t23 GND 0.011256f
C1026 CS_BIAS.t17 GND 0.011256f
C1027 CS_BIAS.n169 GND 0.073052f
C1028 CS_BIAS.n170 GND 0.22285f
C1029 CS_BIAS.t15 GND 0.011256f
C1030 CS_BIAS.t19 GND 0.011256f
C1031 CS_BIAS.n171 GND 0.079012f
C1032 CS_BIAS.t21 GND 0.011256f
C1033 CS_BIAS.t9 GND 0.011256f
C1034 CS_BIAS.n172 GND 0.073052f
C1035 CS_BIAS.n173 GND 0.503344f
C1036 CS_BIAS.n174 GND 0.160155f
C1037 CS_BIAS.n175 GND 0.047301f
C1038 CS_BIAS.n176 GND 0.012195f
C1039 CS_BIAS.n177 GND 0.006543f
C1040 CS_BIAS.t105 GND 0.226601f
C1041 CS_BIAS.n178 GND 0.091803f
C1042 CS_BIAS.n179 GND 0.006543f
C1043 CS_BIAS.n180 GND 0.012195f
C1044 CS_BIAS.n181 GND 0.006543f
C1045 CS_BIAS.n182 GND 0.012603f
C1046 CS_BIAS.n183 GND 0.006543f
C1047 CS_BIAS.n184 GND 0.006596f
C1048 CS_BIAS.n185 GND 0.006543f
C1049 CS_BIAS.t83 GND 0.226601f
C1050 CS_BIAS.n186 GND 0.091803f
C1051 CS_BIAS.n187 GND 0.012195f
C1052 CS_BIAS.n188 GND 0.006543f
C1053 CS_BIAS.n189 GND 0.012195f
C1054 CS_BIAS.n190 GND 0.006543f
C1055 CS_BIAS.t67 GND 0.226601f
C1056 CS_BIAS.n191 GND 0.117336f
C1057 CS_BIAS.t61 GND 0.334543f
C1058 CS_BIAS.n192 GND 0.172166f
C1059 CS_BIAS.n193 GND 0.079011f
C1060 CS_BIAS.n194 GND 0.008884f
C1061 CS_BIAS.n195 GND 0.012195f
C1062 CS_BIAS.n196 GND 0.012195f
C1063 CS_BIAS.n197 GND 0.006543f
C1064 CS_BIAS.n198 GND 0.006543f
C1065 CS_BIAS.n199 GND 0.006543f
C1066 CS_BIAS.n200 GND 0.012633f
C1067 CS_BIAS.n201 GND 0.004276f
C1068 CS_BIAS.n202 GND 0.009107f
C1069 CS_BIAS.n203 GND 0.006543f
C1070 CS_BIAS.n204 GND 0.006543f
C1071 CS_BIAS.n205 GND 0.006543f
C1072 CS_BIAS.n206 GND 0.012195f
C1073 CS_BIAS.n207 GND 0.012195f
C1074 CS_BIAS.n208 GND 0.011774f
C1075 CS_BIAS.n209 GND 0.006543f
C1076 CS_BIAS.n210 GND 0.006543f
C1077 CS_BIAS.n211 GND 0.006543f
C1078 CS_BIAS.n212 GND 0.012195f
C1079 CS_BIAS.n213 GND 0.012195f
C1080 CS_BIAS.n214 GND 0.012195f
C1081 CS_BIAS.n215 GND 0.006543f
C1082 CS_BIAS.n216 GND 0.006543f
C1083 CS_BIAS.n217 GND 0.006543f
C1084 CS_BIAS.n218 GND 0.007464f
C1085 CS_BIAS.n219 GND 0.005003f
C1086 CS_BIAS.n220 GND 0.013142f
C1087 CS_BIAS.n221 GND 0.006543f
C1088 CS_BIAS.n222 GND 0.006543f
C1089 CS_BIAS.n223 GND 0.006543f
C1090 CS_BIAS.n224 GND 0.012195f
C1091 CS_BIAS.n225 GND 0.012195f
C1092 CS_BIAS.n226 GND 0.008041f
C1093 CS_BIAS.n227 GND 0.006543f
C1094 CS_BIAS.n228 GND 0.006543f
C1095 CS_BIAS.n229 GND 0.010328f
C1096 CS_BIAS.n230 GND 0.012195f
C1097 CS_BIAS.n231 GND 0.012195f
C1098 CS_BIAS.n232 GND 0.006543f
C1099 CS_BIAS.n233 GND 0.006543f
C1100 CS_BIAS.n234 GND 0.006512f
C1101 CS_BIAS.n235 GND 0.011103f
C1102 CS_BIAS.n236 GND 0.003811f
C1103 CS_BIAS.n237 GND 0.011103f
C1104 CS_BIAS.n238 GND 0.006512f
C1105 CS_BIAS.n239 GND 0.006543f
C1106 CS_BIAS.n240 GND 0.006543f
C1107 CS_BIAS.n241 GND 0.012195f
C1108 CS_BIAS.n242 GND 0.012195f
C1109 CS_BIAS.n243 GND 0.010328f
C1110 CS_BIAS.n244 GND 0.006543f
C1111 CS_BIAS.n245 GND 0.006543f
C1112 CS_BIAS.n246 GND 0.006543f
C1113 CS_BIAS.n247 GND 0.012195f
C1114 CS_BIAS.n248 GND 0.012195f
C1115 CS_BIAS.n249 GND 0.012195f
C1116 CS_BIAS.n250 GND 0.006543f
C1117 CS_BIAS.n251 GND 0.006543f
C1118 CS_BIAS.n252 GND 0.006543f
C1119 CS_BIAS.n253 GND 0.005003f
C1120 CS_BIAS.n254 GND 0.007464f
C1121 CS_BIAS.n255 GND 0.012603f
C1122 CS_BIAS.n256 GND 0.006543f
C1123 CS_BIAS.n257 GND 0.006543f
C1124 CS_BIAS.n258 GND 0.006543f
C1125 CS_BIAS.n259 GND 0.012195f
C1126 CS_BIAS.n260 GND 0.012195f
C1127 CS_BIAS.n261 GND 0.006596f
C1128 CS_BIAS.n262 GND 0.006543f
C1129 CS_BIAS.n263 GND 0.006543f
C1130 CS_BIAS.n264 GND 0.011774f
C1131 CS_BIAS.n265 GND 0.012195f
C1132 CS_BIAS.n266 GND 0.012195f
C1133 CS_BIAS.n267 GND 0.006543f
C1134 CS_BIAS.n268 GND 0.006543f
C1135 CS_BIAS.n269 GND 0.006543f
C1136 CS_BIAS.n270 GND 0.009107f
C1137 CS_BIAS.n271 GND 0.004276f
C1138 CS_BIAS.n272 GND 0.012633f
C1139 CS_BIAS.n273 GND 0.006543f
C1140 CS_BIAS.n274 GND 0.006543f
C1141 CS_BIAS.n275 GND 0.006543f
C1142 CS_BIAS.n276 GND 0.012195f
C1143 CS_BIAS.n277 GND 0.012195f
C1144 CS_BIAS.n278 GND 0.008884f
C1145 CS_BIAS.n279 GND 0.006543f
C1146 CS_BIAS.n280 GND 0.006543f
C1147 CS_BIAS.n281 GND 0.009486f
C1148 CS_BIAS.n282 GND 0.012195f
C1149 CS_BIAS.n283 GND 0.012195f
C1150 CS_BIAS.n284 GND 0.006543f
C1151 CS_BIAS.n285 GND 0.006543f
C1152 CS_BIAS.n286 GND 0.006543f
C1153 CS_BIAS.n287 GND 0.012073f
C1154 CS_BIAS.n288 GND 0.003964f
C1155 CS_BIAS.n289 GND 0.009979f
C1156 CS_BIAS.n290 GND 0.006543f
C1157 CS_BIAS.n291 GND 0.006543f
C1158 CS_BIAS.n292 GND 0.006543f
C1159 CS_BIAS.n293 GND 0.012195f
C1160 CS_BIAS.n294 GND 0.012195f
C1161 CS_BIAS.n295 GND 0.011172f
C1162 CS_BIAS.n296 GND 0.013846f
C1163 CS_BIAS.n297 GND 0.071671f
C1164 CS_BIAS.t32 GND 0.226601f
C1165 CS_BIAS.n298 GND 0.122067f
C1166 CS_BIAS.n299 GND 0.006543f
C1167 CS_BIAS.n300 GND 0.012195f
C1168 CS_BIAS.n301 GND 0.006543f
C1169 CS_BIAS.n302 GND 0.012195f
C1170 CS_BIAS.n303 GND 0.006543f
C1171 CS_BIAS.t97 GND 0.226601f
C1172 CS_BIAS.n304 GND 0.091803f
C1173 CS_BIAS.n305 GND 0.006543f
C1174 CS_BIAS.n306 GND 0.012195f
C1175 CS_BIAS.n307 GND 0.006543f
C1176 CS_BIAS.n308 GND 0.012195f
C1177 CS_BIAS.n309 GND 0.006543f
C1178 CS_BIAS.t74 GND 0.226601f
C1179 CS_BIAS.n310 GND 0.091803f
C1180 CS_BIAS.n311 GND 0.006543f
C1181 CS_BIAS.n312 GND 0.012195f
C1182 CS_BIAS.n313 GND 0.006543f
C1183 CS_BIAS.n314 GND 0.013142f
C1184 CS_BIAS.n315 GND 0.006543f
C1185 CS_BIAS.n316 GND 0.008041f
C1186 CS_BIAS.n317 GND 0.006543f
C1187 CS_BIAS.t72 GND 0.226601f
C1188 CS_BIAS.n318 GND 0.091803f
C1189 CS_BIAS.n319 GND 0.012195f
C1190 CS_BIAS.n320 GND 0.006543f
C1191 CS_BIAS.n321 GND 0.012195f
C1192 CS_BIAS.n322 GND 0.006543f
C1193 CS_BIAS.t68 GND 0.226601f
C1194 CS_BIAS.n323 GND 0.091803f
C1195 CS_BIAS.n324 GND 0.006543f
C1196 CS_BIAS.n325 GND 0.012195f
C1197 CS_BIAS.n326 GND 0.006543f
C1198 CS_BIAS.n327 GND 0.012603f
C1199 CS_BIAS.n328 GND 0.006543f
C1200 CS_BIAS.n329 GND 0.006596f
C1201 CS_BIAS.n330 GND 0.006543f
C1202 CS_BIAS.t78 GND 0.226601f
C1203 CS_BIAS.n331 GND 0.091803f
C1204 CS_BIAS.n332 GND 0.012195f
C1205 CS_BIAS.n333 GND 0.006543f
C1206 CS_BIAS.n334 GND 0.012195f
C1207 CS_BIAS.n335 GND 0.006543f
C1208 CS_BIAS.t51 GND 0.226601f
C1209 CS_BIAS.n336 GND 0.117336f
C1210 CS_BIAS.t39 GND 0.334543f
C1211 CS_BIAS.n337 GND 0.172166f
C1212 CS_BIAS.n338 GND 0.079011f
C1213 CS_BIAS.n339 GND 0.008884f
C1214 CS_BIAS.n340 GND 0.012195f
C1215 CS_BIAS.n341 GND 0.012195f
C1216 CS_BIAS.n342 GND 0.006543f
C1217 CS_BIAS.n343 GND 0.006543f
C1218 CS_BIAS.n344 GND 0.006543f
C1219 CS_BIAS.n345 GND 0.012633f
C1220 CS_BIAS.n346 GND 0.004276f
C1221 CS_BIAS.n347 GND 0.009107f
C1222 CS_BIAS.n348 GND 0.006543f
C1223 CS_BIAS.n349 GND 0.006543f
C1224 CS_BIAS.n350 GND 0.006543f
C1225 CS_BIAS.n351 GND 0.012195f
C1226 CS_BIAS.n352 GND 0.012195f
C1227 CS_BIAS.n353 GND 0.011774f
C1228 CS_BIAS.n354 GND 0.006543f
C1229 CS_BIAS.n355 GND 0.006543f
C1230 CS_BIAS.n356 GND 0.006543f
C1231 CS_BIAS.n357 GND 0.012195f
C1232 CS_BIAS.n358 GND 0.012195f
C1233 CS_BIAS.n359 GND 0.012195f
C1234 CS_BIAS.n360 GND 0.006543f
C1235 CS_BIAS.n361 GND 0.006543f
C1236 CS_BIAS.n362 GND 0.006543f
C1237 CS_BIAS.n363 GND 0.007464f
C1238 CS_BIAS.n364 GND 0.005003f
C1239 CS_BIAS.n365 GND 0.013142f
C1240 CS_BIAS.n366 GND 0.006543f
C1241 CS_BIAS.n367 GND 0.006543f
C1242 CS_BIAS.n368 GND 0.006543f
C1243 CS_BIAS.n369 GND 0.012195f
C1244 CS_BIAS.n370 GND 0.012195f
C1245 CS_BIAS.n371 GND 0.008041f
C1246 CS_BIAS.n372 GND 0.006543f
C1247 CS_BIAS.n373 GND 0.006543f
C1248 CS_BIAS.n374 GND 0.010328f
C1249 CS_BIAS.n375 GND 0.012195f
C1250 CS_BIAS.n376 GND 0.012195f
C1251 CS_BIAS.n377 GND 0.006543f
C1252 CS_BIAS.n378 GND 0.006543f
C1253 CS_BIAS.n379 GND 0.006543f
C1254 CS_BIAS.n380 GND 0.011103f
C1255 CS_BIAS.n381 GND 0.003811f
C1256 CS_BIAS.n382 GND 0.011103f
C1257 CS_BIAS.n383 GND 0.006543f
C1258 CS_BIAS.n384 GND 0.006543f
C1259 CS_BIAS.n385 GND 0.006543f
C1260 CS_BIAS.n386 GND 0.012195f
C1261 CS_BIAS.n387 GND 0.012195f
C1262 CS_BIAS.n388 GND 0.010328f
C1263 CS_BIAS.n389 GND 0.006543f
C1264 CS_BIAS.n390 GND 0.006543f
C1265 CS_BIAS.n391 GND 0.006543f
C1266 CS_BIAS.n392 GND 0.012195f
C1267 CS_BIAS.n393 GND 0.012195f
C1268 CS_BIAS.n394 GND 0.012195f
C1269 CS_BIAS.n395 GND 0.006543f
C1270 CS_BIAS.n396 GND 0.006543f
C1271 CS_BIAS.n397 GND 0.006543f
C1272 CS_BIAS.n398 GND 0.005003f
C1273 CS_BIAS.n399 GND 0.007464f
C1274 CS_BIAS.n400 GND 0.012603f
C1275 CS_BIAS.n401 GND 0.006543f
C1276 CS_BIAS.n402 GND 0.006543f
C1277 CS_BIAS.n403 GND 0.006543f
C1278 CS_BIAS.n404 GND 0.012195f
C1279 CS_BIAS.n405 GND 0.012195f
C1280 CS_BIAS.n406 GND 0.006596f
C1281 CS_BIAS.n407 GND 0.006543f
C1282 CS_BIAS.n408 GND 0.006543f
C1283 CS_BIAS.n409 GND 0.011774f
C1284 CS_BIAS.n410 GND 0.012195f
C1285 CS_BIAS.n411 GND 0.012195f
C1286 CS_BIAS.n412 GND 0.006543f
C1287 CS_BIAS.n413 GND 0.006543f
C1288 CS_BIAS.n414 GND 0.006543f
C1289 CS_BIAS.n415 GND 0.009107f
C1290 CS_BIAS.n416 GND 0.004276f
C1291 CS_BIAS.n417 GND 0.012633f
C1292 CS_BIAS.n418 GND 0.006543f
C1293 CS_BIAS.n419 GND 0.006543f
C1294 CS_BIAS.n420 GND 0.006543f
C1295 CS_BIAS.n421 GND 0.012195f
C1296 CS_BIAS.n422 GND 0.012195f
C1297 CS_BIAS.n423 GND 0.008884f
C1298 CS_BIAS.n424 GND 0.006543f
C1299 CS_BIAS.n425 GND 0.006543f
C1300 CS_BIAS.n426 GND 0.009486f
C1301 CS_BIAS.n427 GND 0.012195f
C1302 CS_BIAS.n428 GND 0.012195f
C1303 CS_BIAS.n429 GND 0.006543f
C1304 CS_BIAS.n430 GND 0.006543f
C1305 CS_BIAS.n431 GND 0.006543f
C1306 CS_BIAS.n432 GND 0.012073f
C1307 CS_BIAS.n433 GND 0.003964f
C1308 CS_BIAS.n434 GND 0.009979f
C1309 CS_BIAS.n435 GND 0.006543f
C1310 CS_BIAS.n436 GND 0.006543f
C1311 CS_BIAS.n437 GND 0.006543f
C1312 CS_BIAS.n438 GND 0.012195f
C1313 CS_BIAS.n439 GND 0.012195f
C1314 CS_BIAS.n440 GND 0.011172f
C1315 CS_BIAS.n441 GND 0.013846f
C1316 CS_BIAS.n442 GND 0.062082f
C1317 CS_BIAS.n443 GND 0.077922f
C1318 CS_BIAS.t50 GND 0.226601f
C1319 CS_BIAS.n444 GND 0.122067f
C1320 CS_BIAS.n445 GND 0.006543f
C1321 CS_BIAS.n446 GND 0.012195f
C1322 CS_BIAS.n447 GND 0.006543f
C1323 CS_BIAS.n448 GND 0.012195f
C1324 CS_BIAS.n449 GND 0.006543f
C1325 CS_BIAS.t59 GND 0.226601f
C1326 CS_BIAS.n450 GND 0.091803f
C1327 CS_BIAS.n451 GND 0.006543f
C1328 CS_BIAS.n452 GND 0.012195f
C1329 CS_BIAS.n453 GND 0.006543f
C1330 CS_BIAS.n454 GND 0.012195f
C1331 CS_BIAS.n455 GND 0.006543f
C1332 CS_BIAS.t86 GND 0.226601f
C1333 CS_BIAS.n456 GND 0.091803f
C1334 CS_BIAS.n457 GND 0.006543f
C1335 CS_BIAS.n458 GND 0.012195f
C1336 CS_BIAS.n459 GND 0.006543f
C1337 CS_BIAS.n460 GND 0.013142f
C1338 CS_BIAS.n461 GND 0.006543f
C1339 CS_BIAS.n462 GND 0.008041f
C1340 CS_BIAS.n463 GND 0.006543f
C1341 CS_BIAS.t98 GND 0.226601f
C1342 CS_BIAS.n464 GND 0.091803f
C1343 CS_BIAS.n465 GND 0.012195f
C1344 CS_BIAS.n466 GND 0.006543f
C1345 CS_BIAS.n467 GND 0.012195f
C1346 CS_BIAS.n468 GND 0.006543f
C1347 CS_BIAS.t102 GND 0.226601f
C1348 CS_BIAS.n469 GND 0.091803f
C1349 CS_BIAS.n470 GND 0.006543f
C1350 CS_BIAS.n471 GND 0.012195f
C1351 CS_BIAS.n472 GND 0.006543f
C1352 CS_BIAS.n473 GND 0.012603f
C1353 CS_BIAS.n474 GND 0.006543f
C1354 CS_BIAS.n475 GND 0.006596f
C1355 CS_BIAS.n476 GND 0.006543f
C1356 CS_BIAS.t104 GND 0.226601f
C1357 CS_BIAS.n477 GND 0.091803f
C1358 CS_BIAS.n478 GND 0.012195f
C1359 CS_BIAS.n479 GND 0.006543f
C1360 CS_BIAS.n480 GND 0.012195f
C1361 CS_BIAS.n481 GND 0.006543f
C1362 CS_BIAS.t33 GND 0.226601f
C1363 CS_BIAS.n482 GND 0.117336f
C1364 CS_BIAS.t71 GND 0.334543f
C1365 CS_BIAS.n483 GND 0.172166f
C1366 CS_BIAS.n484 GND 0.079011f
C1367 CS_BIAS.n485 GND 0.008884f
C1368 CS_BIAS.n486 GND 0.012195f
C1369 CS_BIAS.n487 GND 0.012195f
C1370 CS_BIAS.n488 GND 0.006543f
C1371 CS_BIAS.n489 GND 0.006543f
C1372 CS_BIAS.n490 GND 0.006543f
C1373 CS_BIAS.n491 GND 0.012633f
C1374 CS_BIAS.n492 GND 0.004276f
C1375 CS_BIAS.n493 GND 0.009107f
C1376 CS_BIAS.n494 GND 0.006543f
C1377 CS_BIAS.n495 GND 0.006543f
C1378 CS_BIAS.n496 GND 0.006543f
C1379 CS_BIAS.n497 GND 0.012195f
C1380 CS_BIAS.n498 GND 0.012195f
C1381 CS_BIAS.n499 GND 0.011774f
C1382 CS_BIAS.n500 GND 0.006543f
C1383 CS_BIAS.n501 GND 0.006543f
C1384 CS_BIAS.n502 GND 0.006543f
C1385 CS_BIAS.n503 GND 0.012195f
C1386 CS_BIAS.n504 GND 0.012195f
C1387 CS_BIAS.n505 GND 0.012195f
C1388 CS_BIAS.n506 GND 0.006543f
C1389 CS_BIAS.n507 GND 0.006543f
C1390 CS_BIAS.n508 GND 0.006543f
C1391 CS_BIAS.n509 GND 0.007464f
C1392 CS_BIAS.n510 GND 0.005003f
C1393 CS_BIAS.n511 GND 0.013142f
C1394 CS_BIAS.n512 GND 0.006543f
C1395 CS_BIAS.n513 GND 0.006543f
C1396 CS_BIAS.n514 GND 0.006543f
C1397 CS_BIAS.n515 GND 0.012195f
C1398 CS_BIAS.n516 GND 0.012195f
C1399 CS_BIAS.n517 GND 0.008041f
C1400 CS_BIAS.n518 GND 0.006543f
C1401 CS_BIAS.n519 GND 0.006543f
C1402 CS_BIAS.n520 GND 0.010328f
C1403 CS_BIAS.n521 GND 0.012195f
C1404 CS_BIAS.n522 GND 0.012195f
C1405 CS_BIAS.n523 GND 0.006543f
C1406 CS_BIAS.n524 GND 0.006543f
C1407 CS_BIAS.n525 GND 0.006543f
C1408 CS_BIAS.n526 GND 0.011103f
C1409 CS_BIAS.n527 GND 0.003811f
C1410 CS_BIAS.n528 GND 0.011103f
C1411 CS_BIAS.n529 GND 0.006543f
C1412 CS_BIAS.n530 GND 0.006543f
C1413 CS_BIAS.n531 GND 0.006543f
C1414 CS_BIAS.n532 GND 0.012195f
C1415 CS_BIAS.n533 GND 0.012195f
C1416 CS_BIAS.n534 GND 0.010328f
C1417 CS_BIAS.n535 GND 0.006543f
C1418 CS_BIAS.n536 GND 0.006543f
C1419 CS_BIAS.n537 GND 0.006543f
C1420 CS_BIAS.n538 GND 0.012195f
C1421 CS_BIAS.n539 GND 0.012195f
C1422 CS_BIAS.n540 GND 0.012195f
C1423 CS_BIAS.n541 GND 0.006543f
C1424 CS_BIAS.n542 GND 0.006543f
C1425 CS_BIAS.n543 GND 0.006543f
C1426 CS_BIAS.n544 GND 0.005003f
C1427 CS_BIAS.n545 GND 0.007464f
C1428 CS_BIAS.n546 GND 0.012603f
C1429 CS_BIAS.n547 GND 0.006543f
C1430 CS_BIAS.n548 GND 0.006543f
C1431 CS_BIAS.n549 GND 0.006543f
C1432 CS_BIAS.n550 GND 0.012195f
C1433 CS_BIAS.n551 GND 0.012195f
C1434 CS_BIAS.n552 GND 0.006596f
C1435 CS_BIAS.n553 GND 0.006543f
C1436 CS_BIAS.n554 GND 0.006543f
C1437 CS_BIAS.n555 GND 0.011774f
C1438 CS_BIAS.n556 GND 0.012195f
C1439 CS_BIAS.n557 GND 0.012195f
C1440 CS_BIAS.n558 GND 0.006543f
C1441 CS_BIAS.n559 GND 0.006543f
C1442 CS_BIAS.n560 GND 0.006543f
C1443 CS_BIAS.n561 GND 0.009107f
C1444 CS_BIAS.n562 GND 0.004276f
C1445 CS_BIAS.n563 GND 0.012633f
C1446 CS_BIAS.n564 GND 0.006543f
C1447 CS_BIAS.n565 GND 0.006543f
C1448 CS_BIAS.n566 GND 0.006543f
C1449 CS_BIAS.n567 GND 0.012195f
C1450 CS_BIAS.n568 GND 0.012195f
C1451 CS_BIAS.n569 GND 0.008884f
C1452 CS_BIAS.n570 GND 0.006543f
C1453 CS_BIAS.n571 GND 0.006543f
C1454 CS_BIAS.n572 GND 0.009486f
C1455 CS_BIAS.n573 GND 0.012195f
C1456 CS_BIAS.n574 GND 0.012195f
C1457 CS_BIAS.n575 GND 0.006543f
C1458 CS_BIAS.n576 GND 0.006543f
C1459 CS_BIAS.n577 GND 0.006543f
C1460 CS_BIAS.n578 GND 0.012073f
C1461 CS_BIAS.n579 GND 0.003964f
C1462 CS_BIAS.n580 GND 0.009979f
C1463 CS_BIAS.n581 GND 0.006543f
C1464 CS_BIAS.n582 GND 0.006543f
C1465 CS_BIAS.n583 GND 0.006543f
C1466 CS_BIAS.n584 GND 0.012195f
C1467 CS_BIAS.n585 GND 0.012195f
C1468 CS_BIAS.n586 GND 0.011172f
C1469 CS_BIAS.n587 GND 0.013846f
C1470 CS_BIAS.n588 GND 0.062082f
C1471 CS_BIAS.n589 GND 0.055435f
C1472 CS_BIAS.t56 GND 0.226601f
C1473 CS_BIAS.n590 GND 0.122067f
C1474 CS_BIAS.n591 GND 0.006543f
C1475 CS_BIAS.n592 GND 0.012195f
C1476 CS_BIAS.n593 GND 0.006543f
C1477 CS_BIAS.n594 GND 0.012195f
C1478 CS_BIAS.n595 GND 0.006543f
C1479 CS_BIAS.t111 GND 0.226601f
C1480 CS_BIAS.n596 GND 0.091803f
C1481 CS_BIAS.n597 GND 0.006543f
C1482 CS_BIAS.n598 GND 0.012195f
C1483 CS_BIAS.n599 GND 0.006543f
C1484 CS_BIAS.n600 GND 0.012195f
C1485 CS_BIAS.n601 GND 0.006543f
C1486 CS_BIAS.t96 GND 0.226601f
C1487 CS_BIAS.n602 GND 0.091803f
C1488 CS_BIAS.n603 GND 0.006543f
C1489 CS_BIAS.n604 GND 0.012195f
C1490 CS_BIAS.n605 GND 0.006543f
C1491 CS_BIAS.n606 GND 0.013142f
C1492 CS_BIAS.n607 GND 0.006543f
C1493 CS_BIAS.n608 GND 0.008041f
C1494 CS_BIAS.n609 GND 0.006543f
C1495 CS_BIAS.t93 GND 0.226601f
C1496 CS_BIAS.n610 GND 0.091803f
C1497 CS_BIAS.n611 GND 0.012195f
C1498 CS_BIAS.n612 GND 0.006543f
C1499 CS_BIAS.n613 GND 0.012195f
C1500 CS_BIAS.n614 GND 0.006543f
C1501 CS_BIAS.t89 GND 0.226601f
C1502 CS_BIAS.n615 GND 0.091803f
C1503 CS_BIAS.n616 GND 0.006543f
C1504 CS_BIAS.n617 GND 0.012195f
C1505 CS_BIAS.n618 GND 0.006543f
C1506 CS_BIAS.n619 GND 0.012603f
C1507 CS_BIAS.n620 GND 0.006543f
C1508 CS_BIAS.n621 GND 0.006596f
C1509 CS_BIAS.n622 GND 0.006543f
C1510 CS_BIAS.t100 GND 0.226601f
C1511 CS_BIAS.n623 GND 0.091803f
C1512 CS_BIAS.n624 GND 0.012195f
C1513 CS_BIAS.n625 GND 0.006543f
C1514 CS_BIAS.n626 GND 0.012195f
C1515 CS_BIAS.n627 GND 0.006543f
C1516 CS_BIAS.t77 GND 0.226601f
C1517 CS_BIAS.n628 GND 0.117336f
C1518 CS_BIAS.t60 GND 0.334543f
C1519 CS_BIAS.n629 GND 0.172166f
C1520 CS_BIAS.n630 GND 0.079011f
C1521 CS_BIAS.n631 GND 0.008884f
C1522 CS_BIAS.n632 GND 0.012195f
C1523 CS_BIAS.n633 GND 0.012195f
C1524 CS_BIAS.n634 GND 0.006543f
C1525 CS_BIAS.n635 GND 0.006543f
C1526 CS_BIAS.n636 GND 0.006543f
C1527 CS_BIAS.n637 GND 0.012633f
C1528 CS_BIAS.n638 GND 0.004276f
C1529 CS_BIAS.n639 GND 0.009107f
C1530 CS_BIAS.n640 GND 0.006543f
C1531 CS_BIAS.n641 GND 0.006543f
C1532 CS_BIAS.n642 GND 0.006543f
C1533 CS_BIAS.n643 GND 0.012195f
C1534 CS_BIAS.n644 GND 0.012195f
C1535 CS_BIAS.n645 GND 0.011774f
C1536 CS_BIAS.n646 GND 0.006543f
C1537 CS_BIAS.n647 GND 0.006543f
C1538 CS_BIAS.n648 GND 0.006543f
C1539 CS_BIAS.n649 GND 0.012195f
C1540 CS_BIAS.n650 GND 0.012195f
C1541 CS_BIAS.n651 GND 0.012195f
C1542 CS_BIAS.n652 GND 0.006543f
C1543 CS_BIAS.n653 GND 0.006543f
C1544 CS_BIAS.n654 GND 0.006543f
C1545 CS_BIAS.n655 GND 0.007464f
C1546 CS_BIAS.n656 GND 0.005003f
C1547 CS_BIAS.n657 GND 0.013142f
C1548 CS_BIAS.n658 GND 0.006543f
C1549 CS_BIAS.n659 GND 0.006543f
C1550 CS_BIAS.n660 GND 0.006543f
C1551 CS_BIAS.n661 GND 0.012195f
C1552 CS_BIAS.n662 GND 0.012195f
C1553 CS_BIAS.n663 GND 0.008041f
C1554 CS_BIAS.n664 GND 0.006543f
C1555 CS_BIAS.n665 GND 0.006543f
C1556 CS_BIAS.n666 GND 0.010328f
C1557 CS_BIAS.n667 GND 0.012195f
C1558 CS_BIAS.n668 GND 0.012195f
C1559 CS_BIAS.n669 GND 0.006543f
C1560 CS_BIAS.n670 GND 0.006543f
C1561 CS_BIAS.n671 GND 0.006543f
C1562 CS_BIAS.n672 GND 0.011103f
C1563 CS_BIAS.n673 GND 0.003811f
C1564 CS_BIAS.n674 GND 0.011103f
C1565 CS_BIAS.n675 GND 0.006543f
C1566 CS_BIAS.n676 GND 0.006543f
C1567 CS_BIAS.n677 GND 0.006543f
C1568 CS_BIAS.n678 GND 0.012195f
C1569 CS_BIAS.n679 GND 0.012195f
C1570 CS_BIAS.n680 GND 0.010328f
C1571 CS_BIAS.n681 GND 0.006543f
C1572 CS_BIAS.n682 GND 0.006543f
C1573 CS_BIAS.n683 GND 0.006543f
C1574 CS_BIAS.n684 GND 0.012195f
C1575 CS_BIAS.n685 GND 0.012195f
C1576 CS_BIAS.n686 GND 0.012195f
C1577 CS_BIAS.n687 GND 0.006543f
C1578 CS_BIAS.n688 GND 0.006543f
C1579 CS_BIAS.n689 GND 0.006543f
C1580 CS_BIAS.n690 GND 0.005003f
C1581 CS_BIAS.n691 GND 0.007464f
C1582 CS_BIAS.n692 GND 0.012603f
C1583 CS_BIAS.n693 GND 0.006543f
C1584 CS_BIAS.n694 GND 0.006543f
C1585 CS_BIAS.n695 GND 0.006543f
C1586 CS_BIAS.n696 GND 0.012195f
C1587 CS_BIAS.n697 GND 0.012195f
C1588 CS_BIAS.n698 GND 0.006596f
C1589 CS_BIAS.n699 GND 0.006543f
C1590 CS_BIAS.n700 GND 0.006543f
C1591 CS_BIAS.n701 GND 0.011774f
C1592 CS_BIAS.n702 GND 0.012195f
C1593 CS_BIAS.n703 GND 0.012195f
C1594 CS_BIAS.n704 GND 0.006543f
C1595 CS_BIAS.n705 GND 0.006543f
C1596 CS_BIAS.n706 GND 0.006543f
C1597 CS_BIAS.n707 GND 0.009107f
C1598 CS_BIAS.n708 GND 0.004276f
C1599 CS_BIAS.n709 GND 0.012633f
C1600 CS_BIAS.n710 GND 0.006543f
C1601 CS_BIAS.n711 GND 0.006543f
C1602 CS_BIAS.n712 GND 0.006543f
C1603 CS_BIAS.n713 GND 0.012195f
C1604 CS_BIAS.n714 GND 0.012195f
C1605 CS_BIAS.n715 GND 0.008884f
C1606 CS_BIAS.n716 GND 0.006543f
C1607 CS_BIAS.n717 GND 0.006543f
C1608 CS_BIAS.n718 GND 0.009486f
C1609 CS_BIAS.n719 GND 0.012195f
C1610 CS_BIAS.n720 GND 0.012195f
C1611 CS_BIAS.n721 GND 0.006543f
C1612 CS_BIAS.n722 GND 0.006543f
C1613 CS_BIAS.n723 GND 0.006543f
C1614 CS_BIAS.n724 GND 0.012073f
C1615 CS_BIAS.n725 GND 0.003964f
C1616 CS_BIAS.n726 GND 0.009979f
C1617 CS_BIAS.n727 GND 0.006543f
C1618 CS_BIAS.n728 GND 0.006543f
C1619 CS_BIAS.n729 GND 0.006543f
C1620 CS_BIAS.n730 GND 0.012195f
C1621 CS_BIAS.n731 GND 0.012195f
C1622 CS_BIAS.n732 GND 0.011172f
C1623 CS_BIAS.n733 GND 0.013846f
C1624 CS_BIAS.n734 GND 0.062082f
C1625 CS_BIAS.n735 GND 0.055435f
C1626 CS_BIAS.t99 GND 0.226601f
C1627 CS_BIAS.n736 GND 0.122067f
C1628 CS_BIAS.n737 GND 0.006543f
C1629 CS_BIAS.n738 GND 0.012195f
C1630 CS_BIAS.n739 GND 0.006543f
C1631 CS_BIAS.n740 GND 0.012195f
C1632 CS_BIAS.n741 GND 0.006543f
C1633 CS_BIAS.t76 GND 0.226601f
C1634 CS_BIAS.n742 GND 0.091803f
C1635 CS_BIAS.n743 GND 0.006543f
C1636 CS_BIAS.n744 GND 0.012195f
C1637 CS_BIAS.n745 GND 0.006543f
C1638 CS_BIAS.n746 GND 0.012195f
C1639 CS_BIAS.n747 GND 0.006543f
C1640 CS_BIAS.t48 GND 0.226601f
C1641 CS_BIAS.n748 GND 0.091803f
C1642 CS_BIAS.n749 GND 0.006543f
C1643 CS_BIAS.n750 GND 0.012195f
C1644 CS_BIAS.n751 GND 0.006543f
C1645 CS_BIAS.n752 GND 0.013142f
C1646 CS_BIAS.n753 GND 0.006543f
C1647 CS_BIAS.n754 GND 0.008041f
C1648 CS_BIAS.n755 GND 0.006543f
C1649 CS_BIAS.t46 GND 0.226601f
C1650 CS_BIAS.n756 GND 0.091803f
C1651 CS_BIAS.n757 GND 0.012195f
C1652 CS_BIAS.n758 GND 0.006543f
C1653 CS_BIAS.n759 GND 0.012195f
C1654 CS_BIAS.n760 GND 0.006543f
C1655 CS_BIAS.t43 GND 0.226601f
C1656 CS_BIAS.n761 GND 0.091803f
C1657 CS_BIAS.n762 GND 0.006543f
C1658 CS_BIAS.n763 GND 0.012195f
C1659 CS_BIAS.n764 GND 0.006543f
C1660 CS_BIAS.n765 GND 0.012603f
C1661 CS_BIAS.n766 GND 0.006543f
C1662 CS_BIAS.n767 GND 0.006596f
C1663 CS_BIAS.n768 GND 0.006543f
C1664 CS_BIAS.t54 GND 0.226601f
C1665 CS_BIAS.n769 GND 0.091803f
C1666 CS_BIAS.n770 GND 0.012195f
C1667 CS_BIAS.n771 GND 0.006543f
C1668 CS_BIAS.n772 GND 0.012195f
C1669 CS_BIAS.n773 GND 0.006543f
C1670 CS_BIAS.t109 GND 0.226601f
C1671 CS_BIAS.n774 GND 0.117336f
C1672 CS_BIAS.t101 GND 0.334543f
C1673 CS_BIAS.n775 GND 0.172165f
C1674 CS_BIAS.n776 GND 0.079011f
C1675 CS_BIAS.n777 GND 0.008884f
C1676 CS_BIAS.n778 GND 0.012195f
C1677 CS_BIAS.n779 GND 0.012195f
C1678 CS_BIAS.n780 GND 0.006543f
C1679 CS_BIAS.n781 GND 0.006543f
C1680 CS_BIAS.n782 GND 0.006543f
C1681 CS_BIAS.n783 GND 0.012633f
C1682 CS_BIAS.n784 GND 0.004276f
C1683 CS_BIAS.n785 GND 0.009107f
C1684 CS_BIAS.n786 GND 0.006543f
C1685 CS_BIAS.n787 GND 0.006543f
C1686 CS_BIAS.n788 GND 0.006543f
C1687 CS_BIAS.n789 GND 0.012195f
C1688 CS_BIAS.n790 GND 0.012195f
C1689 CS_BIAS.n791 GND 0.011774f
C1690 CS_BIAS.n792 GND 0.006543f
C1691 CS_BIAS.n793 GND 0.006543f
C1692 CS_BIAS.n794 GND 0.006543f
C1693 CS_BIAS.n795 GND 0.012195f
C1694 CS_BIAS.n796 GND 0.012195f
C1695 CS_BIAS.n797 GND 0.012195f
C1696 CS_BIAS.n798 GND 0.006543f
C1697 CS_BIAS.n799 GND 0.006543f
C1698 CS_BIAS.n800 GND 0.006543f
C1699 CS_BIAS.n801 GND 0.007464f
C1700 CS_BIAS.n802 GND 0.005003f
C1701 CS_BIAS.n803 GND 0.013142f
C1702 CS_BIAS.n804 GND 0.006543f
C1703 CS_BIAS.n805 GND 0.006543f
C1704 CS_BIAS.n806 GND 0.006543f
C1705 CS_BIAS.n807 GND 0.012195f
C1706 CS_BIAS.n808 GND 0.012195f
C1707 CS_BIAS.n809 GND 0.008041f
C1708 CS_BIAS.n810 GND 0.006543f
C1709 CS_BIAS.n811 GND 0.006543f
C1710 CS_BIAS.n812 GND 0.010328f
C1711 CS_BIAS.n813 GND 0.012195f
C1712 CS_BIAS.n814 GND 0.012195f
C1713 CS_BIAS.n815 GND 0.006543f
C1714 CS_BIAS.n816 GND 0.006543f
C1715 CS_BIAS.n817 GND 0.006543f
C1716 CS_BIAS.n818 GND 0.011103f
C1717 CS_BIAS.n819 GND 0.003811f
C1718 CS_BIAS.n820 GND 0.011103f
C1719 CS_BIAS.n821 GND 0.006543f
C1720 CS_BIAS.n822 GND 0.006543f
C1721 CS_BIAS.n823 GND 0.006543f
C1722 CS_BIAS.n824 GND 0.012195f
C1723 CS_BIAS.n825 GND 0.012195f
C1724 CS_BIAS.n826 GND 0.010328f
C1725 CS_BIAS.n827 GND 0.006543f
C1726 CS_BIAS.n828 GND 0.006543f
C1727 CS_BIAS.n829 GND 0.006543f
C1728 CS_BIAS.n830 GND 0.012195f
C1729 CS_BIAS.n831 GND 0.012195f
C1730 CS_BIAS.n832 GND 0.012195f
C1731 CS_BIAS.n833 GND 0.006543f
C1732 CS_BIAS.n834 GND 0.006543f
C1733 CS_BIAS.n835 GND 0.006543f
C1734 CS_BIAS.n836 GND 0.005003f
C1735 CS_BIAS.n837 GND 0.007464f
C1736 CS_BIAS.n838 GND 0.012603f
C1737 CS_BIAS.n839 GND 0.006543f
C1738 CS_BIAS.n840 GND 0.006543f
C1739 CS_BIAS.n841 GND 0.006543f
C1740 CS_BIAS.n842 GND 0.012195f
C1741 CS_BIAS.n843 GND 0.012195f
C1742 CS_BIAS.n844 GND 0.006596f
C1743 CS_BIAS.n845 GND 0.006543f
C1744 CS_BIAS.n846 GND 0.006543f
C1745 CS_BIAS.n847 GND 0.011774f
C1746 CS_BIAS.n848 GND 0.012195f
C1747 CS_BIAS.n849 GND 0.012195f
C1748 CS_BIAS.n850 GND 0.006543f
C1749 CS_BIAS.n851 GND 0.006543f
C1750 CS_BIAS.n852 GND 0.006543f
C1751 CS_BIAS.n853 GND 0.009107f
C1752 CS_BIAS.n854 GND 0.004276f
C1753 CS_BIAS.n855 GND 0.012633f
C1754 CS_BIAS.n856 GND 0.006543f
C1755 CS_BIAS.n857 GND 0.006543f
C1756 CS_BIAS.n858 GND 0.006543f
C1757 CS_BIAS.n859 GND 0.012195f
C1758 CS_BIAS.n860 GND 0.012195f
C1759 CS_BIAS.n861 GND 0.008884f
C1760 CS_BIAS.n862 GND 0.006543f
C1761 CS_BIAS.n863 GND 0.006543f
C1762 CS_BIAS.n864 GND 0.009486f
C1763 CS_BIAS.n865 GND 0.012195f
C1764 CS_BIAS.n866 GND 0.012195f
C1765 CS_BIAS.n867 GND 0.006543f
C1766 CS_BIAS.n868 GND 0.006543f
C1767 CS_BIAS.n869 GND 0.006543f
C1768 CS_BIAS.n870 GND 0.012073f
C1769 CS_BIAS.n871 GND 0.003964f
C1770 CS_BIAS.n872 GND 0.009979f
C1771 CS_BIAS.n873 GND 0.006543f
C1772 CS_BIAS.n874 GND 0.006543f
C1773 CS_BIAS.n875 GND 0.006543f
C1774 CS_BIAS.n876 GND 0.012195f
C1775 CS_BIAS.n877 GND 0.012195f
C1776 CS_BIAS.n878 GND 0.011172f
C1777 CS_BIAS.n879 GND 0.013846f
C1778 CS_BIAS.n880 GND 0.062082f
C1779 CS_BIAS.n881 GND 0.864455f
C1780 CS_BIAS.t85 GND 0.226601f
C1781 CS_BIAS.n882 GND 0.122067f
C1782 CS_BIAS.n883 GND 0.006543f
C1783 CS_BIAS.n884 GND 0.012195f
C1784 CS_BIAS.n885 GND 0.006543f
C1785 CS_BIAS.n886 GND 0.012195f
C1786 CS_BIAS.n887 GND 0.006543f
C1787 CS_BIAS.t45 GND 0.226601f
C1788 CS_BIAS.n888 GND 0.091803f
C1789 CS_BIAS.n889 GND 0.006543f
C1790 CS_BIAS.n890 GND 0.012195f
C1791 CS_BIAS.n891 GND 0.006543f
C1792 CS_BIAS.n892 GND 0.012195f
C1793 CS_BIAS.n893 GND 0.006543f
C1794 CS_BIAS.t34 GND 0.226601f
C1795 CS_BIAS.n894 GND 0.091803f
C1796 CS_BIAS.n895 GND 0.006543f
C1797 CS_BIAS.n896 GND 0.012195f
C1798 CS_BIAS.n897 GND 0.006543f
C1799 CS_BIAS.n898 GND 0.013142f
C1800 CS_BIAS.n899 GND 0.006543f
C1801 CS_BIAS.n900 GND 0.008041f
C1802 CS_BIAS.n901 GND 0.006543f
C1803 CS_BIAS.n902 GND 0.012195f
C1804 CS_BIAS.t31 GND 0.011256f
C1805 CS_BIAS.t11 GND 0.011256f
C1806 CS_BIAS.n903 GND 0.079012f
C1807 CS_BIAS.t25 GND 0.011256f
C1808 CS_BIAS.t5 GND 0.011256f
C1809 CS_BIAS.n904 GND 0.073052f
C1810 CS_BIAS.n905 GND 0.503344f
C1811 CS_BIAS.t6 GND 0.226601f
C1812 CS_BIAS.n906 GND 0.122067f
C1813 CS_BIAS.n907 GND 0.006543f
C1814 CS_BIAS.n908 GND 0.012195f
C1815 CS_BIAS.n909 GND 0.006543f
C1816 CS_BIAS.n910 GND 0.012195f
C1817 CS_BIAS.n911 GND 0.006543f
C1818 CS_BIAS.t2 GND 0.226601f
C1819 CS_BIAS.n912 GND 0.091803f
C1820 CS_BIAS.n913 GND 0.006543f
C1821 CS_BIAS.n914 GND 0.012195f
C1822 CS_BIAS.n915 GND 0.006543f
C1823 CS_BIAS.n916 GND 0.012195f
C1824 CS_BIAS.n917 GND 0.006543f
C1825 CS_BIAS.t28 GND 0.226601f
C1826 CS_BIAS.n918 GND 0.091803f
C1827 CS_BIAS.n919 GND 0.006543f
C1828 CS_BIAS.n920 GND 0.012195f
C1829 CS_BIAS.n921 GND 0.006543f
C1830 CS_BIAS.n922 GND 0.013142f
C1831 CS_BIAS.n923 GND 0.006543f
C1832 CS_BIAS.n924 GND 0.008041f
C1833 CS_BIAS.n925 GND 0.006543f
C1834 CS_BIAS.n926 GND 0.012195f
C1835 CS_BIAS.n927 GND 0.006543f
C1836 CS_BIAS.n928 GND 0.012195f
C1837 CS_BIAS.n929 GND 0.006543f
C1838 CS_BIAS.t4 GND 0.226601f
C1839 CS_BIAS.n930 GND 0.091803f
C1840 CS_BIAS.n931 GND 0.006543f
C1841 CS_BIAS.n932 GND 0.012195f
C1842 CS_BIAS.n933 GND 0.006543f
C1843 CS_BIAS.n934 GND 0.012603f
C1844 CS_BIAS.n935 GND 0.006543f
C1845 CS_BIAS.n936 GND 0.006596f
C1846 CS_BIAS.n937 GND 0.006543f
C1847 CS_BIAS.n938 GND 0.012195f
C1848 CS_BIAS.n939 GND 0.006543f
C1849 CS_BIAS.n940 GND 0.012195f
C1850 CS_BIAS.n941 GND 0.006543f
C1851 CS_BIAS.t10 GND 0.226601f
C1852 CS_BIAS.n942 GND 0.117336f
C1853 CS_BIAS.t30 GND 0.334543f
C1854 CS_BIAS.n943 GND 0.172165f
C1855 CS_BIAS.n944 GND 0.079011f
C1856 CS_BIAS.n945 GND 0.008884f
C1857 CS_BIAS.n946 GND 0.012195f
C1858 CS_BIAS.n947 GND 0.012195f
C1859 CS_BIAS.n948 GND 0.006543f
C1860 CS_BIAS.n949 GND 0.006543f
C1861 CS_BIAS.n950 GND 0.006543f
C1862 CS_BIAS.n951 GND 0.012633f
C1863 CS_BIAS.n952 GND 0.004276f
C1864 CS_BIAS.n953 GND 0.009107f
C1865 CS_BIAS.n954 GND 0.006543f
C1866 CS_BIAS.n955 GND 0.006543f
C1867 CS_BIAS.n956 GND 0.006543f
C1868 CS_BIAS.n957 GND 0.012195f
C1869 CS_BIAS.n958 GND 0.012195f
C1870 CS_BIAS.t24 GND 0.226601f
C1871 CS_BIAS.n959 GND 0.091803f
C1872 CS_BIAS.n960 GND 0.011774f
C1873 CS_BIAS.n961 GND 0.006543f
C1874 CS_BIAS.n962 GND 0.006543f
C1875 CS_BIAS.n963 GND 0.006543f
C1876 CS_BIAS.n964 GND 0.012195f
C1877 CS_BIAS.n965 GND 0.012195f
C1878 CS_BIAS.n966 GND 0.012195f
C1879 CS_BIAS.n967 GND 0.006543f
C1880 CS_BIAS.n968 GND 0.006543f
C1881 CS_BIAS.n969 GND 0.006543f
C1882 CS_BIAS.n970 GND 0.007464f
C1883 CS_BIAS.n971 GND 0.005003f
C1884 CS_BIAS.n972 GND 0.013142f
C1885 CS_BIAS.n973 GND 0.006543f
C1886 CS_BIAS.n974 GND 0.006543f
C1887 CS_BIAS.n975 GND 0.006543f
C1888 CS_BIAS.n976 GND 0.012195f
C1889 CS_BIAS.n977 GND 0.012195f
C1890 CS_BIAS.n978 GND 0.008041f
C1891 CS_BIAS.n979 GND 0.006543f
C1892 CS_BIAS.n980 GND 0.006543f
C1893 CS_BIAS.n981 GND 0.010328f
C1894 CS_BIAS.n982 GND 0.012195f
C1895 CS_BIAS.n983 GND 0.012195f
C1896 CS_BIAS.n984 GND 0.006543f
C1897 CS_BIAS.n985 GND 0.006543f
C1898 CS_BIAS.n986 GND 0.006543f
C1899 CS_BIAS.n987 GND 0.011103f
C1900 CS_BIAS.n988 GND 0.003811f
C1901 CS_BIAS.n989 GND 0.011103f
C1902 CS_BIAS.n990 GND 0.006543f
C1903 CS_BIAS.n991 GND 0.006543f
C1904 CS_BIAS.n992 GND 0.006543f
C1905 CS_BIAS.n993 GND 0.012195f
C1906 CS_BIAS.n994 GND 0.012195f
C1907 CS_BIAS.t12 GND 0.226601f
C1908 CS_BIAS.n995 GND 0.091803f
C1909 CS_BIAS.n996 GND 0.010328f
C1910 CS_BIAS.n997 GND 0.006543f
C1911 CS_BIAS.n998 GND 0.006543f
C1912 CS_BIAS.n999 GND 0.006543f
C1913 CS_BIAS.n1000 GND 0.012195f
C1914 CS_BIAS.n1001 GND 0.012195f
C1915 CS_BIAS.n1002 GND 0.012195f
C1916 CS_BIAS.n1003 GND 0.006543f
C1917 CS_BIAS.n1004 GND 0.006543f
C1918 CS_BIAS.n1005 GND 0.006543f
C1919 CS_BIAS.n1006 GND 0.005003f
C1920 CS_BIAS.n1007 GND 0.007464f
C1921 CS_BIAS.n1008 GND 0.012603f
C1922 CS_BIAS.n1009 GND 0.006543f
C1923 CS_BIAS.n1010 GND 0.006543f
C1924 CS_BIAS.n1011 GND 0.006543f
C1925 CS_BIAS.n1012 GND 0.012195f
C1926 CS_BIAS.n1013 GND 0.012195f
C1927 CS_BIAS.n1014 GND 0.006596f
C1928 CS_BIAS.n1015 GND 0.006543f
C1929 CS_BIAS.n1016 GND 0.006543f
C1930 CS_BIAS.n1017 GND 0.011774f
C1931 CS_BIAS.n1018 GND 0.012195f
C1932 CS_BIAS.n1019 GND 0.012195f
C1933 CS_BIAS.n1020 GND 0.006543f
C1934 CS_BIAS.n1021 GND 0.006543f
C1935 CS_BIAS.n1022 GND 0.006543f
C1936 CS_BIAS.n1023 GND 0.009107f
C1937 CS_BIAS.n1024 GND 0.004276f
C1938 CS_BIAS.n1025 GND 0.012633f
C1939 CS_BIAS.n1026 GND 0.006543f
C1940 CS_BIAS.n1027 GND 0.006543f
C1941 CS_BIAS.n1028 GND 0.006543f
C1942 CS_BIAS.n1029 GND 0.012195f
C1943 CS_BIAS.n1030 GND 0.012195f
C1944 CS_BIAS.n1031 GND 0.008884f
C1945 CS_BIAS.n1032 GND 0.006543f
C1946 CS_BIAS.n1033 GND 0.006543f
C1947 CS_BIAS.n1034 GND 0.009486f
C1948 CS_BIAS.n1035 GND 0.012195f
C1949 CS_BIAS.n1036 GND 0.012195f
C1950 CS_BIAS.n1037 GND 0.006543f
C1951 CS_BIAS.n1038 GND 0.006543f
C1952 CS_BIAS.n1039 GND 0.006543f
C1953 CS_BIAS.n1040 GND 0.012073f
C1954 CS_BIAS.n1041 GND 0.003964f
C1955 CS_BIAS.n1042 GND 0.009979f
C1956 CS_BIAS.n1043 GND 0.006543f
C1957 CS_BIAS.n1044 GND 0.006543f
C1958 CS_BIAS.n1045 GND 0.006543f
C1959 CS_BIAS.n1046 GND 0.012195f
C1960 CS_BIAS.n1047 GND 0.012195f
C1961 CS_BIAS.n1048 GND 0.011172f
C1962 CS_BIAS.n1049 GND 0.013846f
C1963 CS_BIAS.n1050 GND 0.107996f
C1964 CS_BIAS.t3 GND 0.011256f
C1965 CS_BIAS.t7 GND 0.011256f
C1966 CS_BIAS.n1051 GND 0.073052f
C1967 CS_BIAS.n1052 GND 0.321859f
C1968 CS_BIAS.t13 GND 0.011256f
C1969 CS_BIAS.t29 GND 0.011256f
C1970 CS_BIAS.n1053 GND 0.073052f
C1971 CS_BIAS.n1054 GND 0.22285f
C1972 CS_BIAS.n1055 GND 0.160155f
C1973 CS_BIAS.n1056 GND 0.047301f
C1974 CS_BIAS.n1057 GND 0.012195f
C1975 CS_BIAS.n1058 GND 0.006543f
C1976 CS_BIAS.t57 GND 0.226601f
C1977 CS_BIAS.n1059 GND 0.091803f
C1978 CS_BIAS.n1060 GND 0.006543f
C1979 CS_BIAS.n1061 GND 0.012195f
C1980 CS_BIAS.n1062 GND 0.006543f
C1981 CS_BIAS.n1063 GND 0.012603f
C1982 CS_BIAS.n1064 GND 0.006543f
C1983 CS_BIAS.n1065 GND 0.006596f
C1984 CS_BIAS.n1066 GND 0.006543f
C1985 CS_BIAS.n1067 GND 0.012195f
C1986 CS_BIAS.n1068 GND 0.006543f
C1987 CS_BIAS.n1069 GND 0.012195f
C1988 CS_BIAS.n1070 GND 0.006543f
C1989 CS_BIAS.t80 GND 0.226601f
C1990 CS_BIAS.n1071 GND 0.117336f
C1991 CS_BIAS.t38 GND 0.334543f
C1992 CS_BIAS.n1072 GND 0.172165f
C1993 CS_BIAS.n1073 GND 0.079011f
C1994 CS_BIAS.n1074 GND 0.008884f
C1995 CS_BIAS.n1075 GND 0.012195f
C1996 CS_BIAS.n1076 GND 0.012195f
C1997 CS_BIAS.n1077 GND 0.006543f
C1998 CS_BIAS.n1078 GND 0.006543f
C1999 CS_BIAS.n1079 GND 0.006543f
C2000 CS_BIAS.n1080 GND 0.012633f
C2001 CS_BIAS.n1081 GND 0.004276f
C2002 CS_BIAS.n1082 GND 0.009107f
C2003 CS_BIAS.n1083 GND 0.006543f
C2004 CS_BIAS.n1084 GND 0.006543f
C2005 CS_BIAS.n1085 GND 0.006543f
C2006 CS_BIAS.n1086 GND 0.012195f
C2007 CS_BIAS.n1087 GND 0.012195f
C2008 CS_BIAS.t37 GND 0.226601f
C2009 CS_BIAS.n1088 GND 0.091803f
C2010 CS_BIAS.n1089 GND 0.011774f
C2011 CS_BIAS.n1090 GND 0.006543f
C2012 CS_BIAS.n1091 GND 0.006543f
C2013 CS_BIAS.n1092 GND 0.006543f
C2014 CS_BIAS.n1093 GND 0.012195f
C2015 CS_BIAS.n1094 GND 0.012195f
C2016 CS_BIAS.n1095 GND 0.012195f
C2017 CS_BIAS.n1096 GND 0.006543f
C2018 CS_BIAS.n1097 GND 0.006543f
C2019 CS_BIAS.n1098 GND 0.006543f
C2020 CS_BIAS.n1099 GND 0.007464f
C2021 CS_BIAS.n1100 GND 0.005003f
C2022 CS_BIAS.n1101 GND 0.013142f
C2023 CS_BIAS.n1102 GND 0.006543f
C2024 CS_BIAS.n1103 GND 0.006543f
C2025 CS_BIAS.n1104 GND 0.006543f
C2026 CS_BIAS.n1105 GND 0.012195f
C2027 CS_BIAS.n1106 GND 0.012195f
C2028 CS_BIAS.n1107 GND 0.008041f
C2029 CS_BIAS.n1108 GND 0.006543f
C2030 CS_BIAS.n1109 GND 0.006543f
C2031 CS_BIAS.n1110 GND 0.010328f
C2032 CS_BIAS.n1111 GND 0.012195f
C2033 CS_BIAS.n1112 GND 0.012195f
C2034 CS_BIAS.n1113 GND 0.006543f
C2035 CS_BIAS.n1114 GND 0.006543f
C2036 CS_BIAS.n1115 GND 0.006512f
C2037 CS_BIAS.n1116 GND 0.011103f
C2038 CS_BIAS.n1117 GND 0.003811f
C2039 CS_BIAS.n1118 GND 0.011103f
C2040 CS_BIAS.n1119 GND 0.006512f
C2041 CS_BIAS.n1120 GND 0.006543f
C2042 CS_BIAS.n1121 GND 0.006543f
C2043 CS_BIAS.n1122 GND 0.012195f
C2044 CS_BIAS.n1123 GND 0.012195f
C2045 CS_BIAS.t79 GND 0.226601f
C2046 CS_BIAS.n1124 GND 0.091803f
C2047 CS_BIAS.n1125 GND 0.010328f
C2048 CS_BIAS.n1126 GND 0.006543f
C2049 CS_BIAS.n1127 GND 0.006543f
C2050 CS_BIAS.n1128 GND 0.006543f
C2051 CS_BIAS.n1129 GND 0.012195f
C2052 CS_BIAS.n1130 GND 0.012195f
C2053 CS_BIAS.n1131 GND 0.012195f
C2054 CS_BIAS.n1132 GND 0.006543f
C2055 CS_BIAS.n1133 GND 0.006543f
C2056 CS_BIAS.n1134 GND 0.006543f
C2057 CS_BIAS.n1135 GND 0.005003f
C2058 CS_BIAS.n1136 GND 0.007464f
C2059 CS_BIAS.n1137 GND 0.012603f
C2060 CS_BIAS.n1138 GND 0.006543f
C2061 CS_BIAS.n1139 GND 0.006543f
C2062 CS_BIAS.n1140 GND 0.006543f
C2063 CS_BIAS.n1141 GND 0.012195f
C2064 CS_BIAS.n1142 GND 0.012195f
C2065 CS_BIAS.n1143 GND 0.006596f
C2066 CS_BIAS.n1144 GND 0.006543f
C2067 CS_BIAS.n1145 GND 0.006543f
C2068 CS_BIAS.n1146 GND 0.011774f
C2069 CS_BIAS.n1147 GND 0.012195f
C2070 CS_BIAS.n1148 GND 0.012195f
C2071 CS_BIAS.n1149 GND 0.006543f
C2072 CS_BIAS.n1150 GND 0.006543f
C2073 CS_BIAS.n1151 GND 0.006543f
C2074 CS_BIAS.n1152 GND 0.009107f
C2075 CS_BIAS.n1153 GND 0.004276f
C2076 CS_BIAS.n1154 GND 0.012633f
C2077 CS_BIAS.n1155 GND 0.006543f
C2078 CS_BIAS.n1156 GND 0.006543f
C2079 CS_BIAS.n1157 GND 0.006543f
C2080 CS_BIAS.n1158 GND 0.012195f
C2081 CS_BIAS.n1159 GND 0.012195f
C2082 CS_BIAS.n1160 GND 0.008884f
C2083 CS_BIAS.n1161 GND 0.006543f
C2084 CS_BIAS.n1162 GND 0.006543f
C2085 CS_BIAS.n1163 GND 0.009486f
C2086 CS_BIAS.n1164 GND 0.012195f
C2087 CS_BIAS.n1165 GND 0.012195f
C2088 CS_BIAS.n1166 GND 0.006543f
C2089 CS_BIAS.n1167 GND 0.006543f
C2090 CS_BIAS.n1168 GND 0.006543f
C2091 CS_BIAS.n1169 GND 0.012073f
C2092 CS_BIAS.n1170 GND 0.003964f
C2093 CS_BIAS.n1171 GND 0.009979f
C2094 CS_BIAS.n1172 GND 0.006543f
C2095 CS_BIAS.n1173 GND 0.006543f
C2096 CS_BIAS.n1174 GND 0.006543f
C2097 CS_BIAS.n1175 GND 0.012195f
C2098 CS_BIAS.n1176 GND 0.012195f
C2099 CS_BIAS.n1177 GND 0.011172f
C2100 CS_BIAS.n1178 GND 0.013846f
C2101 CS_BIAS.n1179 GND 0.071671f
C2102 CS_BIAS.t110 GND 0.226601f
C2103 CS_BIAS.n1180 GND 0.122067f
C2104 CS_BIAS.n1181 GND 0.006543f
C2105 CS_BIAS.n1182 GND 0.012195f
C2106 CS_BIAS.n1183 GND 0.006543f
C2107 CS_BIAS.n1184 GND 0.012195f
C2108 CS_BIAS.n1185 GND 0.006543f
C2109 CS_BIAS.t108 GND 0.226601f
C2110 CS_BIAS.n1186 GND 0.091803f
C2111 CS_BIAS.n1187 GND 0.006543f
C2112 CS_BIAS.n1188 GND 0.012195f
C2113 CS_BIAS.n1189 GND 0.006543f
C2114 CS_BIAS.n1190 GND 0.012195f
C2115 CS_BIAS.n1191 GND 0.006543f
C2116 CS_BIAS.t87 GND 0.226601f
C2117 CS_BIAS.n1192 GND 0.091803f
C2118 CS_BIAS.n1193 GND 0.006543f
C2119 CS_BIAS.n1194 GND 0.012195f
C2120 CS_BIAS.n1195 GND 0.006543f
C2121 CS_BIAS.n1196 GND 0.013142f
C2122 CS_BIAS.n1197 GND 0.006543f
C2123 CS_BIAS.n1198 GND 0.008041f
C2124 CS_BIAS.n1199 GND 0.006543f
C2125 CS_BIAS.n1200 GND 0.012195f
C2126 CS_BIAS.n1201 GND 0.006543f
C2127 CS_BIAS.n1202 GND 0.012195f
C2128 CS_BIAS.n1203 GND 0.006543f
C2129 CS_BIAS.t62 GND 0.226601f
C2130 CS_BIAS.n1204 GND 0.091803f
C2131 CS_BIAS.n1205 GND 0.006543f
C2132 CS_BIAS.n1206 GND 0.012195f
C2133 CS_BIAS.n1207 GND 0.006543f
C2134 CS_BIAS.n1208 GND 0.012603f
C2135 CS_BIAS.n1209 GND 0.006543f
C2136 CS_BIAS.n1210 GND 0.006596f
C2137 CS_BIAS.n1211 GND 0.006543f
C2138 CS_BIAS.n1212 GND 0.012195f
C2139 CS_BIAS.n1213 GND 0.006543f
C2140 CS_BIAS.n1214 GND 0.012195f
C2141 CS_BIAS.n1215 GND 0.006543f
C2142 CS_BIAS.t70 GND 0.226601f
C2143 CS_BIAS.n1216 GND 0.117336f
C2144 CS_BIAS.t66 GND 0.334543f
C2145 CS_BIAS.n1217 GND 0.172165f
C2146 CS_BIAS.n1218 GND 0.079011f
C2147 CS_BIAS.n1219 GND 0.008884f
C2148 CS_BIAS.n1220 GND 0.012195f
C2149 CS_BIAS.n1221 GND 0.012195f
C2150 CS_BIAS.n1222 GND 0.006543f
C2151 CS_BIAS.n1223 GND 0.006543f
C2152 CS_BIAS.n1224 GND 0.006543f
C2153 CS_BIAS.n1225 GND 0.012633f
C2154 CS_BIAS.n1226 GND 0.004276f
C2155 CS_BIAS.n1227 GND 0.009107f
C2156 CS_BIAS.n1228 GND 0.006543f
C2157 CS_BIAS.n1229 GND 0.006543f
C2158 CS_BIAS.n1230 GND 0.006543f
C2159 CS_BIAS.n1231 GND 0.012195f
C2160 CS_BIAS.n1232 GND 0.012195f
C2161 CS_BIAS.t73 GND 0.226601f
C2162 CS_BIAS.n1233 GND 0.091803f
C2163 CS_BIAS.n1234 GND 0.011774f
C2164 CS_BIAS.n1235 GND 0.006543f
C2165 CS_BIAS.n1236 GND 0.006543f
C2166 CS_BIAS.n1237 GND 0.006543f
C2167 CS_BIAS.n1238 GND 0.012195f
C2168 CS_BIAS.n1239 GND 0.012195f
C2169 CS_BIAS.n1240 GND 0.012195f
C2170 CS_BIAS.n1241 GND 0.006543f
C2171 CS_BIAS.n1242 GND 0.006543f
C2172 CS_BIAS.n1243 GND 0.006543f
C2173 CS_BIAS.n1244 GND 0.007464f
C2174 CS_BIAS.n1245 GND 0.005003f
C2175 CS_BIAS.n1246 GND 0.013142f
C2176 CS_BIAS.n1247 GND 0.006543f
C2177 CS_BIAS.n1248 GND 0.006543f
C2178 CS_BIAS.n1249 GND 0.006543f
C2179 CS_BIAS.n1250 GND 0.012195f
C2180 CS_BIAS.n1251 GND 0.012195f
C2181 CS_BIAS.n1252 GND 0.008041f
C2182 CS_BIAS.n1253 GND 0.006543f
C2183 CS_BIAS.n1254 GND 0.006543f
C2184 CS_BIAS.n1255 GND 0.010328f
C2185 CS_BIAS.n1256 GND 0.012195f
C2186 CS_BIAS.n1257 GND 0.012195f
C2187 CS_BIAS.n1258 GND 0.006543f
C2188 CS_BIAS.n1259 GND 0.006543f
C2189 CS_BIAS.n1260 GND 0.006543f
C2190 CS_BIAS.n1261 GND 0.011103f
C2191 CS_BIAS.n1262 GND 0.003811f
C2192 CS_BIAS.n1263 GND 0.011103f
C2193 CS_BIAS.n1264 GND 0.006543f
C2194 CS_BIAS.n1265 GND 0.006543f
C2195 CS_BIAS.n1266 GND 0.006543f
C2196 CS_BIAS.n1267 GND 0.012195f
C2197 CS_BIAS.n1268 GND 0.012195f
C2198 CS_BIAS.t84 GND 0.226601f
C2199 CS_BIAS.n1269 GND 0.091803f
C2200 CS_BIAS.n1270 GND 0.010328f
C2201 CS_BIAS.n1271 GND 0.006543f
C2202 CS_BIAS.n1272 GND 0.006543f
C2203 CS_BIAS.n1273 GND 0.006543f
C2204 CS_BIAS.n1274 GND 0.012195f
C2205 CS_BIAS.n1275 GND 0.012195f
C2206 CS_BIAS.n1276 GND 0.012195f
C2207 CS_BIAS.n1277 GND 0.006543f
C2208 CS_BIAS.n1278 GND 0.006543f
C2209 CS_BIAS.n1279 GND 0.006543f
C2210 CS_BIAS.n1280 GND 0.005003f
C2211 CS_BIAS.n1281 GND 0.007464f
C2212 CS_BIAS.n1282 GND 0.012603f
C2213 CS_BIAS.n1283 GND 0.006543f
C2214 CS_BIAS.n1284 GND 0.006543f
C2215 CS_BIAS.n1285 GND 0.006543f
C2216 CS_BIAS.n1286 GND 0.012195f
C2217 CS_BIAS.n1287 GND 0.012195f
C2218 CS_BIAS.n1288 GND 0.006596f
C2219 CS_BIAS.n1289 GND 0.006543f
C2220 CS_BIAS.n1290 GND 0.006543f
C2221 CS_BIAS.n1291 GND 0.011774f
C2222 CS_BIAS.n1292 GND 0.012195f
C2223 CS_BIAS.n1293 GND 0.012195f
C2224 CS_BIAS.n1294 GND 0.006543f
C2225 CS_BIAS.n1295 GND 0.006543f
C2226 CS_BIAS.n1296 GND 0.006543f
C2227 CS_BIAS.n1297 GND 0.009107f
C2228 CS_BIAS.n1298 GND 0.004276f
C2229 CS_BIAS.n1299 GND 0.012633f
C2230 CS_BIAS.n1300 GND 0.006543f
C2231 CS_BIAS.n1301 GND 0.006543f
C2232 CS_BIAS.n1302 GND 0.006543f
C2233 CS_BIAS.n1303 GND 0.012195f
C2234 CS_BIAS.n1304 GND 0.012195f
C2235 CS_BIAS.n1305 GND 0.008884f
C2236 CS_BIAS.n1306 GND 0.006543f
C2237 CS_BIAS.n1307 GND 0.006543f
C2238 CS_BIAS.n1308 GND 0.009486f
C2239 CS_BIAS.n1309 GND 0.012195f
C2240 CS_BIAS.n1310 GND 0.012195f
C2241 CS_BIAS.n1311 GND 0.006543f
C2242 CS_BIAS.n1312 GND 0.006543f
C2243 CS_BIAS.n1313 GND 0.006543f
C2244 CS_BIAS.n1314 GND 0.012073f
C2245 CS_BIAS.n1315 GND 0.003964f
C2246 CS_BIAS.n1316 GND 0.009979f
C2247 CS_BIAS.n1317 GND 0.006543f
C2248 CS_BIAS.n1318 GND 0.006543f
C2249 CS_BIAS.n1319 GND 0.006543f
C2250 CS_BIAS.n1320 GND 0.012195f
C2251 CS_BIAS.n1321 GND 0.012195f
C2252 CS_BIAS.n1322 GND 0.011172f
C2253 CS_BIAS.n1323 GND 0.013846f
C2254 CS_BIAS.n1324 GND 0.062082f
C2255 CS_BIAS.n1325 GND 0.077922f
C2256 CS_BIAS.t81 GND 0.226601f
C2257 CS_BIAS.n1326 GND 0.122067f
C2258 CS_BIAS.n1327 GND 0.006543f
C2259 CS_BIAS.n1328 GND 0.012195f
C2260 CS_BIAS.n1329 GND 0.006543f
C2261 CS_BIAS.n1330 GND 0.012195f
C2262 CS_BIAS.n1331 GND 0.006543f
C2263 CS_BIAS.t91 GND 0.226601f
C2264 CS_BIAS.n1332 GND 0.091803f
C2265 CS_BIAS.n1333 GND 0.006543f
C2266 CS_BIAS.n1334 GND 0.012195f
C2267 CS_BIAS.n1335 GND 0.006543f
C2268 CS_BIAS.n1336 GND 0.012195f
C2269 CS_BIAS.n1337 GND 0.006543f
C2270 CS_BIAS.t36 GND 0.226601f
C2271 CS_BIAS.n1338 GND 0.091803f
C2272 CS_BIAS.n1339 GND 0.006543f
C2273 CS_BIAS.n1340 GND 0.012195f
C2274 CS_BIAS.n1341 GND 0.006543f
C2275 CS_BIAS.n1342 GND 0.013142f
C2276 CS_BIAS.n1343 GND 0.006543f
C2277 CS_BIAS.n1344 GND 0.008041f
C2278 CS_BIAS.n1345 GND 0.006543f
C2279 CS_BIAS.n1346 GND 0.012195f
C2280 CS_BIAS.n1347 GND 0.006543f
C2281 CS_BIAS.n1348 GND 0.012195f
C2282 CS_BIAS.n1349 GND 0.006543f
C2283 CS_BIAS.t52 GND 0.226601f
C2284 CS_BIAS.n1350 GND 0.091803f
C2285 CS_BIAS.n1351 GND 0.006543f
C2286 CS_BIAS.n1352 GND 0.012195f
C2287 CS_BIAS.n1353 GND 0.006543f
C2288 CS_BIAS.n1354 GND 0.012603f
C2289 CS_BIAS.n1355 GND 0.006543f
C2290 CS_BIAS.n1356 GND 0.006596f
C2291 CS_BIAS.n1357 GND 0.006543f
C2292 CS_BIAS.n1358 GND 0.012195f
C2293 CS_BIAS.n1359 GND 0.006543f
C2294 CS_BIAS.n1360 GND 0.012195f
C2295 CS_BIAS.n1361 GND 0.006543f
C2296 CS_BIAS.t63 GND 0.226601f
C2297 CS_BIAS.n1362 GND 0.117336f
C2298 CS_BIAS.t75 GND 0.334543f
C2299 CS_BIAS.n1363 GND 0.172165f
C2300 CS_BIAS.n1364 GND 0.079011f
C2301 CS_BIAS.n1365 GND 0.008884f
C2302 CS_BIAS.n1366 GND 0.012195f
C2303 CS_BIAS.n1367 GND 0.012195f
C2304 CS_BIAS.n1368 GND 0.006543f
C2305 CS_BIAS.n1369 GND 0.006543f
C2306 CS_BIAS.n1370 GND 0.006543f
C2307 CS_BIAS.n1371 GND 0.012633f
C2308 CS_BIAS.n1372 GND 0.004276f
C2309 CS_BIAS.n1373 GND 0.009107f
C2310 CS_BIAS.n1374 GND 0.006543f
C2311 CS_BIAS.n1375 GND 0.006543f
C2312 CS_BIAS.n1376 GND 0.006543f
C2313 CS_BIAS.n1377 GND 0.012195f
C2314 CS_BIAS.n1378 GND 0.012195f
C2315 CS_BIAS.t58 GND 0.226601f
C2316 CS_BIAS.n1379 GND 0.091803f
C2317 CS_BIAS.n1380 GND 0.011774f
C2318 CS_BIAS.n1381 GND 0.006543f
C2319 CS_BIAS.n1382 GND 0.006543f
C2320 CS_BIAS.n1383 GND 0.006543f
C2321 CS_BIAS.n1384 GND 0.012195f
C2322 CS_BIAS.n1385 GND 0.012195f
C2323 CS_BIAS.n1386 GND 0.012195f
C2324 CS_BIAS.n1387 GND 0.006543f
C2325 CS_BIAS.n1388 GND 0.006543f
C2326 CS_BIAS.n1389 GND 0.006543f
C2327 CS_BIAS.n1390 GND 0.007464f
C2328 CS_BIAS.n1391 GND 0.005003f
C2329 CS_BIAS.n1392 GND 0.013142f
C2330 CS_BIAS.n1393 GND 0.006543f
C2331 CS_BIAS.n1394 GND 0.006543f
C2332 CS_BIAS.n1395 GND 0.006543f
C2333 CS_BIAS.n1396 GND 0.012195f
C2334 CS_BIAS.n1397 GND 0.012195f
C2335 CS_BIAS.n1398 GND 0.008041f
C2336 CS_BIAS.n1399 GND 0.006543f
C2337 CS_BIAS.n1400 GND 0.006543f
C2338 CS_BIAS.n1401 GND 0.010328f
C2339 CS_BIAS.n1402 GND 0.012195f
C2340 CS_BIAS.n1403 GND 0.012195f
C2341 CS_BIAS.n1404 GND 0.006543f
C2342 CS_BIAS.n1405 GND 0.006543f
C2343 CS_BIAS.n1406 GND 0.006543f
C2344 CS_BIAS.n1407 GND 0.011103f
C2345 CS_BIAS.n1408 GND 0.003811f
C2346 CS_BIAS.n1409 GND 0.011103f
C2347 CS_BIAS.n1410 GND 0.006543f
C2348 CS_BIAS.n1411 GND 0.006543f
C2349 CS_BIAS.n1412 GND 0.006543f
C2350 CS_BIAS.n1413 GND 0.012195f
C2351 CS_BIAS.n1414 GND 0.012195f
C2352 CS_BIAS.t40 GND 0.226601f
C2353 CS_BIAS.n1415 GND 0.091803f
C2354 CS_BIAS.n1416 GND 0.010328f
C2355 CS_BIAS.n1417 GND 0.006543f
C2356 CS_BIAS.n1418 GND 0.006543f
C2357 CS_BIAS.n1419 GND 0.006543f
C2358 CS_BIAS.n1420 GND 0.012195f
C2359 CS_BIAS.n1421 GND 0.012195f
C2360 CS_BIAS.n1422 GND 0.012195f
C2361 CS_BIAS.n1423 GND 0.006543f
C2362 CS_BIAS.n1424 GND 0.006543f
C2363 CS_BIAS.n1425 GND 0.006543f
C2364 CS_BIAS.n1426 GND 0.005003f
C2365 CS_BIAS.n1427 GND 0.007464f
C2366 CS_BIAS.n1428 GND 0.012603f
C2367 CS_BIAS.n1429 GND 0.006543f
C2368 CS_BIAS.n1430 GND 0.006543f
C2369 CS_BIAS.n1431 GND 0.006543f
C2370 CS_BIAS.n1432 GND 0.012195f
C2371 CS_BIAS.n1433 GND 0.012195f
C2372 CS_BIAS.n1434 GND 0.006596f
C2373 CS_BIAS.n1435 GND 0.006543f
C2374 CS_BIAS.n1436 GND 0.006543f
C2375 CS_BIAS.n1437 GND 0.011774f
C2376 CS_BIAS.n1438 GND 0.012195f
C2377 CS_BIAS.n1439 GND 0.012195f
C2378 CS_BIAS.n1440 GND 0.006543f
C2379 CS_BIAS.n1441 GND 0.006543f
C2380 CS_BIAS.n1442 GND 0.006543f
C2381 CS_BIAS.n1443 GND 0.009107f
C2382 CS_BIAS.n1444 GND 0.004276f
C2383 CS_BIAS.n1445 GND 0.012633f
C2384 CS_BIAS.n1446 GND 0.006543f
C2385 CS_BIAS.n1447 GND 0.006543f
C2386 CS_BIAS.n1448 GND 0.006543f
C2387 CS_BIAS.n1449 GND 0.012195f
C2388 CS_BIAS.n1450 GND 0.012195f
C2389 CS_BIAS.n1451 GND 0.008884f
C2390 CS_BIAS.n1452 GND 0.006543f
C2391 CS_BIAS.n1453 GND 0.006543f
C2392 CS_BIAS.n1454 GND 0.009486f
C2393 CS_BIAS.n1455 GND 0.012195f
C2394 CS_BIAS.n1456 GND 0.012195f
C2395 CS_BIAS.n1457 GND 0.006543f
C2396 CS_BIAS.n1458 GND 0.006543f
C2397 CS_BIAS.n1459 GND 0.006543f
C2398 CS_BIAS.n1460 GND 0.012073f
C2399 CS_BIAS.n1461 GND 0.003964f
C2400 CS_BIAS.n1462 GND 0.009979f
C2401 CS_BIAS.n1463 GND 0.006543f
C2402 CS_BIAS.n1464 GND 0.006543f
C2403 CS_BIAS.n1465 GND 0.006543f
C2404 CS_BIAS.n1466 GND 0.012195f
C2405 CS_BIAS.n1467 GND 0.012195f
C2406 CS_BIAS.n1468 GND 0.011172f
C2407 CS_BIAS.n1469 GND 0.013846f
C2408 CS_BIAS.n1470 GND 0.062082f
C2409 CS_BIAS.n1471 GND 0.055435f
C2410 CS_BIAS.t53 GND 0.226601f
C2411 CS_BIAS.n1472 GND 0.122067f
C2412 CS_BIAS.n1473 GND 0.006543f
C2413 CS_BIAS.n1474 GND 0.012195f
C2414 CS_BIAS.n1475 GND 0.006543f
C2415 CS_BIAS.n1476 GND 0.012195f
C2416 CS_BIAS.n1477 GND 0.006543f
C2417 CS_BIAS.t49 GND 0.226601f
C2418 CS_BIAS.n1478 GND 0.091803f
C2419 CS_BIAS.n1479 GND 0.006543f
C2420 CS_BIAS.n1480 GND 0.012195f
C2421 CS_BIAS.n1481 GND 0.006543f
C2422 CS_BIAS.n1482 GND 0.012195f
C2423 CS_BIAS.n1483 GND 0.006543f
C2424 CS_BIAS.t107 GND 0.226601f
C2425 CS_BIAS.n1484 GND 0.091803f
C2426 CS_BIAS.n1485 GND 0.006543f
C2427 CS_BIAS.n1486 GND 0.012195f
C2428 CS_BIAS.n1487 GND 0.006543f
C2429 CS_BIAS.n1488 GND 0.013142f
C2430 CS_BIAS.n1489 GND 0.006543f
C2431 CS_BIAS.n1490 GND 0.008041f
C2432 CS_BIAS.n1491 GND 0.006543f
C2433 CS_BIAS.n1492 GND 0.012195f
C2434 CS_BIAS.n1493 GND 0.006543f
C2435 CS_BIAS.n1494 GND 0.012195f
C2436 CS_BIAS.n1495 GND 0.006543f
C2437 CS_BIAS.t82 GND 0.226601f
C2438 CS_BIAS.n1496 GND 0.091803f
C2439 CS_BIAS.n1497 GND 0.006543f
C2440 CS_BIAS.n1498 GND 0.012195f
C2441 CS_BIAS.n1499 GND 0.006543f
C2442 CS_BIAS.n1500 GND 0.012603f
C2443 CS_BIAS.n1501 GND 0.006543f
C2444 CS_BIAS.n1502 GND 0.006596f
C2445 CS_BIAS.n1503 GND 0.006543f
C2446 CS_BIAS.n1504 GND 0.012195f
C2447 CS_BIAS.n1505 GND 0.006543f
C2448 CS_BIAS.n1506 GND 0.012195f
C2449 CS_BIAS.n1507 GND 0.006543f
C2450 CS_BIAS.t92 GND 0.226601f
C2451 CS_BIAS.n1508 GND 0.117336f
C2452 CS_BIAS.t88 GND 0.334543f
C2453 CS_BIAS.n1509 GND 0.172165f
C2454 CS_BIAS.n1510 GND 0.079011f
C2455 CS_BIAS.n1511 GND 0.008884f
C2456 CS_BIAS.n1512 GND 0.012195f
C2457 CS_BIAS.n1513 GND 0.012195f
C2458 CS_BIAS.n1514 GND 0.006543f
C2459 CS_BIAS.n1515 GND 0.006543f
C2460 CS_BIAS.n1516 GND 0.006543f
C2461 CS_BIAS.n1517 GND 0.012633f
C2462 CS_BIAS.n1518 GND 0.004276f
C2463 CS_BIAS.n1519 GND 0.009107f
C2464 CS_BIAS.n1520 GND 0.006543f
C2465 CS_BIAS.n1521 GND 0.006543f
C2466 CS_BIAS.n1522 GND 0.006543f
C2467 CS_BIAS.n1523 GND 0.012195f
C2468 CS_BIAS.n1524 GND 0.012195f
C2469 CS_BIAS.t95 GND 0.226601f
C2470 CS_BIAS.n1525 GND 0.091803f
C2471 CS_BIAS.n1526 GND 0.011774f
C2472 CS_BIAS.n1527 GND 0.006543f
C2473 CS_BIAS.n1528 GND 0.006543f
C2474 CS_BIAS.n1529 GND 0.006543f
C2475 CS_BIAS.n1530 GND 0.012195f
C2476 CS_BIAS.n1531 GND 0.012195f
C2477 CS_BIAS.n1532 GND 0.012195f
C2478 CS_BIAS.n1533 GND 0.006543f
C2479 CS_BIAS.n1534 GND 0.006543f
C2480 CS_BIAS.n1535 GND 0.006543f
C2481 CS_BIAS.n1536 GND 0.007464f
C2482 CS_BIAS.n1537 GND 0.005003f
C2483 CS_BIAS.n1538 GND 0.013142f
C2484 CS_BIAS.n1539 GND 0.006543f
C2485 CS_BIAS.n1540 GND 0.006543f
C2486 CS_BIAS.n1541 GND 0.006543f
C2487 CS_BIAS.n1542 GND 0.012195f
C2488 CS_BIAS.n1543 GND 0.012195f
C2489 CS_BIAS.n1544 GND 0.008041f
C2490 CS_BIAS.n1545 GND 0.006543f
C2491 CS_BIAS.n1546 GND 0.006543f
C2492 CS_BIAS.n1547 GND 0.010328f
C2493 CS_BIAS.n1548 GND 0.012195f
C2494 CS_BIAS.n1549 GND 0.012195f
C2495 CS_BIAS.n1550 GND 0.006543f
C2496 CS_BIAS.n1551 GND 0.006543f
C2497 CS_BIAS.n1552 GND 0.006543f
C2498 CS_BIAS.n1553 GND 0.011103f
C2499 CS_BIAS.n1554 GND 0.003811f
C2500 CS_BIAS.n1555 GND 0.011103f
C2501 CS_BIAS.n1556 GND 0.006543f
C2502 CS_BIAS.n1557 GND 0.006543f
C2503 CS_BIAS.n1558 GND 0.006543f
C2504 CS_BIAS.n1559 GND 0.012195f
C2505 CS_BIAS.n1560 GND 0.012195f
C2506 CS_BIAS.t106 GND 0.226601f
C2507 CS_BIAS.n1561 GND 0.091803f
C2508 CS_BIAS.n1562 GND 0.010328f
C2509 CS_BIAS.n1563 GND 0.006543f
C2510 CS_BIAS.n1564 GND 0.006543f
C2511 CS_BIAS.n1565 GND 0.006543f
C2512 CS_BIAS.n1566 GND 0.012195f
C2513 CS_BIAS.n1567 GND 0.012195f
C2514 CS_BIAS.n1568 GND 0.012195f
C2515 CS_BIAS.n1569 GND 0.006543f
C2516 CS_BIAS.n1570 GND 0.006543f
C2517 CS_BIAS.n1571 GND 0.006543f
C2518 CS_BIAS.n1572 GND 0.005003f
C2519 CS_BIAS.n1573 GND 0.007464f
C2520 CS_BIAS.n1574 GND 0.012603f
C2521 CS_BIAS.n1575 GND 0.006543f
C2522 CS_BIAS.n1576 GND 0.006543f
C2523 CS_BIAS.n1577 GND 0.006543f
C2524 CS_BIAS.n1578 GND 0.012195f
C2525 CS_BIAS.n1579 GND 0.012195f
C2526 CS_BIAS.n1580 GND 0.006596f
C2527 CS_BIAS.n1581 GND 0.006543f
C2528 CS_BIAS.n1582 GND 0.006543f
C2529 CS_BIAS.n1583 GND 0.011774f
C2530 CS_BIAS.n1584 GND 0.012195f
C2531 CS_BIAS.n1585 GND 0.012195f
C2532 CS_BIAS.n1586 GND 0.006543f
C2533 CS_BIAS.n1587 GND 0.006543f
C2534 CS_BIAS.n1588 GND 0.006543f
C2535 CS_BIAS.n1589 GND 0.009107f
C2536 CS_BIAS.n1590 GND 0.004276f
C2537 CS_BIAS.n1591 GND 0.012633f
C2538 CS_BIAS.n1592 GND 0.006543f
C2539 CS_BIAS.n1593 GND 0.006543f
C2540 CS_BIAS.n1594 GND 0.006543f
C2541 CS_BIAS.n1595 GND 0.012195f
C2542 CS_BIAS.n1596 GND 0.012195f
C2543 CS_BIAS.n1597 GND 0.008884f
C2544 CS_BIAS.n1598 GND 0.006543f
C2545 CS_BIAS.n1599 GND 0.006543f
C2546 CS_BIAS.n1600 GND 0.009486f
C2547 CS_BIAS.n1601 GND 0.012195f
C2548 CS_BIAS.n1602 GND 0.012195f
C2549 CS_BIAS.n1603 GND 0.006543f
C2550 CS_BIAS.n1604 GND 0.006543f
C2551 CS_BIAS.n1605 GND 0.006543f
C2552 CS_BIAS.n1606 GND 0.012073f
C2553 CS_BIAS.n1607 GND 0.003964f
C2554 CS_BIAS.n1608 GND 0.009979f
C2555 CS_BIAS.n1609 GND 0.006543f
C2556 CS_BIAS.n1610 GND 0.006543f
C2557 CS_BIAS.n1611 GND 0.006543f
C2558 CS_BIAS.n1612 GND 0.012195f
C2559 CS_BIAS.n1613 GND 0.012195f
C2560 CS_BIAS.n1614 GND 0.011172f
C2561 CS_BIAS.n1615 GND 0.013846f
C2562 CS_BIAS.n1616 GND 0.062082f
C2563 CS_BIAS.n1617 GND 0.055435f
C2564 CS_BIAS.t94 GND 0.226601f
C2565 CS_BIAS.n1618 GND 0.122067f
C2566 CS_BIAS.n1619 GND 0.006543f
C2567 CS_BIAS.n1620 GND 0.012195f
C2568 CS_BIAS.n1621 GND 0.006543f
C2569 CS_BIAS.n1622 GND 0.012195f
C2570 CS_BIAS.n1623 GND 0.006543f
C2571 CS_BIAS.t90 GND 0.226601f
C2572 CS_BIAS.n1624 GND 0.091803f
C2573 CS_BIAS.n1625 GND 0.006543f
C2574 CS_BIAS.n1626 GND 0.012195f
C2575 CS_BIAS.n1627 GND 0.006543f
C2576 CS_BIAS.n1628 GND 0.012195f
C2577 CS_BIAS.n1629 GND 0.006543f
C2578 CS_BIAS.t69 GND 0.226601f
C2579 CS_BIAS.n1630 GND 0.091803f
C2580 CS_BIAS.n1631 GND 0.006543f
C2581 CS_BIAS.n1632 GND 0.012195f
C2582 CS_BIAS.n1633 GND 0.006543f
C2583 CS_BIAS.n1634 GND 0.013142f
C2584 CS_BIAS.n1635 GND 0.006543f
C2585 CS_BIAS.n1636 GND 0.008041f
C2586 CS_BIAS.n1637 GND 0.006543f
C2587 CS_BIAS.n1638 GND 0.012195f
C2588 CS_BIAS.n1639 GND 0.006543f
C2589 CS_BIAS.n1640 GND 0.012195f
C2590 CS_BIAS.n1641 GND 0.006543f
C2591 CS_BIAS.t41 GND 0.226601f
C2592 CS_BIAS.n1642 GND 0.091803f
C2593 CS_BIAS.n1643 GND 0.006543f
C2594 CS_BIAS.n1644 GND 0.012195f
C2595 CS_BIAS.n1645 GND 0.006543f
C2596 CS_BIAS.n1646 GND 0.012603f
C2597 CS_BIAS.n1647 GND 0.006543f
C2598 CS_BIAS.n1648 GND 0.006596f
C2599 CS_BIAS.n1649 GND 0.006543f
C2600 CS_BIAS.n1650 GND 0.012195f
C2601 CS_BIAS.n1651 GND 0.006543f
C2602 CS_BIAS.n1652 GND 0.012195f
C2603 CS_BIAS.n1653 GND 0.006543f
C2604 CS_BIAS.t44 GND 0.226601f
C2605 CS_BIAS.n1654 GND 0.117336f
C2606 CS_BIAS.t42 GND 0.334543f
C2607 CS_BIAS.n1655 GND 0.172165f
C2608 CS_BIAS.n1656 GND 0.079011f
C2609 CS_BIAS.n1657 GND 0.008884f
C2610 CS_BIAS.n1658 GND 0.012195f
C2611 CS_BIAS.n1659 GND 0.012195f
C2612 CS_BIAS.n1660 GND 0.006543f
C2613 CS_BIAS.n1661 GND 0.006543f
C2614 CS_BIAS.n1662 GND 0.006543f
C2615 CS_BIAS.n1663 GND 0.012633f
C2616 CS_BIAS.n1664 GND 0.004276f
C2617 CS_BIAS.n1665 GND 0.009107f
C2618 CS_BIAS.n1666 GND 0.006543f
C2619 CS_BIAS.n1667 GND 0.006543f
C2620 CS_BIAS.n1668 GND 0.006543f
C2621 CS_BIAS.n1669 GND 0.012195f
C2622 CS_BIAS.n1670 GND 0.012195f
C2623 CS_BIAS.t47 GND 0.226601f
C2624 CS_BIAS.n1671 GND 0.091803f
C2625 CS_BIAS.n1672 GND 0.011774f
C2626 CS_BIAS.n1673 GND 0.006543f
C2627 CS_BIAS.n1674 GND 0.006543f
C2628 CS_BIAS.n1675 GND 0.006543f
C2629 CS_BIAS.n1676 GND 0.012195f
C2630 CS_BIAS.n1677 GND 0.012195f
C2631 CS_BIAS.n1678 GND 0.012195f
C2632 CS_BIAS.n1679 GND 0.006543f
C2633 CS_BIAS.n1680 GND 0.006543f
C2634 CS_BIAS.n1681 GND 0.006543f
C2635 CS_BIAS.n1682 GND 0.007464f
C2636 CS_BIAS.n1683 GND 0.005003f
C2637 CS_BIAS.n1684 GND 0.013142f
C2638 CS_BIAS.n1685 GND 0.006543f
C2639 CS_BIAS.n1686 GND 0.006543f
C2640 CS_BIAS.n1687 GND 0.006543f
C2641 CS_BIAS.n1688 GND 0.012195f
C2642 CS_BIAS.n1689 GND 0.012195f
C2643 CS_BIAS.n1690 GND 0.008041f
C2644 CS_BIAS.n1691 GND 0.006543f
C2645 CS_BIAS.n1692 GND 0.006543f
C2646 CS_BIAS.n1693 GND 0.010328f
C2647 CS_BIAS.n1694 GND 0.012195f
C2648 CS_BIAS.n1695 GND 0.012195f
C2649 CS_BIAS.n1696 GND 0.006543f
C2650 CS_BIAS.n1697 GND 0.006543f
C2651 CS_BIAS.n1698 GND 0.006543f
C2652 CS_BIAS.n1699 GND 0.011103f
C2653 CS_BIAS.n1700 GND 0.003811f
C2654 CS_BIAS.n1701 GND 0.011103f
C2655 CS_BIAS.n1702 GND 0.006543f
C2656 CS_BIAS.n1703 GND 0.006543f
C2657 CS_BIAS.n1704 GND 0.006543f
C2658 CS_BIAS.n1705 GND 0.012195f
C2659 CS_BIAS.n1706 GND 0.012195f
C2660 CS_BIAS.t65 GND 0.226601f
C2661 CS_BIAS.n1707 GND 0.091803f
C2662 CS_BIAS.n1708 GND 0.010328f
C2663 CS_BIAS.n1709 GND 0.006543f
C2664 CS_BIAS.n1710 GND 0.006543f
C2665 CS_BIAS.n1711 GND 0.006543f
C2666 CS_BIAS.n1712 GND 0.012195f
C2667 CS_BIAS.n1713 GND 0.012195f
C2668 CS_BIAS.n1714 GND 0.012195f
C2669 CS_BIAS.n1715 GND 0.006543f
C2670 CS_BIAS.n1716 GND 0.006543f
C2671 CS_BIAS.n1717 GND 0.006543f
C2672 CS_BIAS.n1718 GND 0.005003f
C2673 CS_BIAS.n1719 GND 0.007464f
C2674 CS_BIAS.n1720 GND 0.012603f
C2675 CS_BIAS.n1721 GND 0.006543f
C2676 CS_BIAS.n1722 GND 0.006543f
C2677 CS_BIAS.n1723 GND 0.006543f
C2678 CS_BIAS.n1724 GND 0.012195f
C2679 CS_BIAS.n1725 GND 0.012195f
C2680 CS_BIAS.n1726 GND 0.006596f
C2681 CS_BIAS.n1727 GND 0.006543f
C2682 CS_BIAS.n1728 GND 0.006543f
C2683 CS_BIAS.n1729 GND 0.011774f
C2684 CS_BIAS.n1730 GND 0.012195f
C2685 CS_BIAS.n1731 GND 0.012195f
C2686 CS_BIAS.n1732 GND 0.006543f
C2687 CS_BIAS.n1733 GND 0.006543f
C2688 CS_BIAS.n1734 GND 0.006543f
C2689 CS_BIAS.n1735 GND 0.009107f
C2690 CS_BIAS.n1736 GND 0.004276f
C2691 CS_BIAS.n1737 GND 0.012633f
C2692 CS_BIAS.n1738 GND 0.006543f
C2693 CS_BIAS.n1739 GND 0.006543f
C2694 CS_BIAS.n1740 GND 0.006543f
C2695 CS_BIAS.n1741 GND 0.012195f
C2696 CS_BIAS.n1742 GND 0.012195f
C2697 CS_BIAS.n1743 GND 0.008884f
C2698 CS_BIAS.n1744 GND 0.006543f
C2699 CS_BIAS.n1745 GND 0.006543f
C2700 CS_BIAS.n1746 GND 0.009486f
C2701 CS_BIAS.n1747 GND 0.012195f
C2702 CS_BIAS.n1748 GND 0.012195f
C2703 CS_BIAS.n1749 GND 0.006543f
C2704 CS_BIAS.n1750 GND 0.006543f
C2705 CS_BIAS.n1751 GND 0.006543f
C2706 CS_BIAS.n1752 GND 0.012073f
C2707 CS_BIAS.n1753 GND 0.003964f
C2708 CS_BIAS.n1754 GND 0.009979f
C2709 CS_BIAS.n1755 GND 0.006543f
C2710 CS_BIAS.n1756 GND 0.006543f
C2711 CS_BIAS.n1757 GND 0.006543f
C2712 CS_BIAS.n1758 GND 0.012195f
C2713 CS_BIAS.n1759 GND 0.012195f
C2714 CS_BIAS.n1760 GND 0.011172f
C2715 CS_BIAS.n1761 GND 0.013846f
C2716 CS_BIAS.n1762 GND 0.062082f
C2717 CS_BIAS.n1763 GND 0.108829f
C2718 CS_BIAS.n1764 GND 5.69798f
C2719 VDD.t129 GND 0.02549f
C2720 VDD.t141 GND 0.02549f
C2721 VDD.n0 GND 0.145137f
C2722 VDD.t155 GND 0.02549f
C2723 VDD.t138 GND 0.02549f
C2724 VDD.n1 GND 0.140928f
C2725 VDD.n2 GND 0.662777f
C2726 VDD.t147 GND 0.02549f
C2727 VDD.t157 GND 0.02549f
C2728 VDD.n3 GND 0.140928f
C2729 VDD.n4 GND 0.345139f
C2730 VDD.t133 GND 0.02549f
C2731 VDD.t153 GND 0.02549f
C2732 VDD.n5 GND 0.140928f
C2733 VDD.n6 GND 0.293401f
C2734 VDD.t131 GND 0.02549f
C2735 VDD.t145 GND 0.02549f
C2736 VDD.n7 GND 0.145137f
C2737 VDD.t119 GND 0.02549f
C2738 VDD.t149 GND 0.02549f
C2739 VDD.n8 GND 0.140928f
C2740 VDD.n9 GND 0.662778f
C2741 VDD.t151 GND 0.02549f
C2742 VDD.t122 GND 0.02549f
C2743 VDD.n10 GND 0.140928f
C2744 VDD.n11 GND 0.345139f
C2745 VDD.t135 GND 0.02549f
C2746 VDD.t126 GND 0.02549f
C2747 VDD.n12 GND 0.140928f
C2748 VDD.n13 GND 0.293401f
C2749 VDD.n14 GND 0.201231f
C2750 VDD.n15 GND 2.50955f
C2751 VDD.t82 GND 0.147596f
C2752 VDD.t80 GND 0.024054f
C2753 VDD.t104 GND 0.024054f
C2754 VDD.n16 GND 0.106517f
C2755 VDD.n17 GND 0.66799f
C2756 VDD.t102 GND 0.024054f
C2757 VDD.t101 GND 0.024054f
C2758 VDD.n18 GND 0.106517f
C2759 VDD.n19 GND 0.401201f
C2760 VDD.t100 GND 0.142539f
C2761 VDD.n20 GND 0.321523f
C2762 VDD.t113 GND 0.147596f
C2763 VDD.t96 GND 0.024054f
C2764 VDD.t108 GND 0.024054f
C2765 VDD.n21 GND 0.106517f
C2766 VDD.n22 GND 0.66799f
C2767 VDD.t84 GND 0.024054f
C2768 VDD.t71 GND 0.024054f
C2769 VDD.n23 GND 0.106517f
C2770 VDD.n24 GND 0.401201f
C2771 VDD.t114 GND 0.142539f
C2772 VDD.n25 GND 0.298186f
C2773 VDD.n26 GND 0.307678f
C2774 VDD.t112 GND 0.147596f
C2775 VDD.t95 GND 0.024054f
C2776 VDD.t105 GND 0.024054f
C2777 VDD.n27 GND 0.106517f
C2778 VDD.n28 GND 0.66799f
C2779 VDD.t87 GND 0.024054f
C2780 VDD.t72 GND 0.024054f
C2781 VDD.n29 GND 0.106517f
C2782 VDD.n30 GND 0.401201f
C2783 VDD.t115 GND 0.142539f
C2784 VDD.n31 GND 0.298186f
C2785 VDD.n32 GND 0.378384f
C2786 VDD.n33 GND 0.004726f
C2787 VDD.n34 GND 0.006149f
C2788 VDD.n35 GND 0.004949f
C2789 VDD.n36 GND 0.006149f
C2790 VDD.n37 GND 0.004949f
C2791 VDD.n38 GND 0.006149f
C2792 VDD.n39 GND 0.498548f
C2793 VDD.n40 GND 0.006149f
C2794 VDD.n41 GND 0.006149f
C2795 VDD.n42 GND 0.006149f
C2796 VDD.n43 GND 0.498548f
C2797 VDD.n44 GND 0.006149f
C2798 VDD.n45 GND 0.006149f
C2799 VDD.n46 GND 0.006149f
C2800 VDD.n47 GND 0.006149f
C2801 VDD.n48 GND 0.006149f
C2802 VDD.n49 GND 0.004949f
C2803 VDD.n50 GND 0.006149f
C2804 VDD.n51 GND 0.006149f
C2805 VDD.n52 GND 0.006149f
C2806 VDD.n53 GND 0.006149f
C2807 VDD.n54 GND 0.498548f
C2808 VDD.n55 GND 0.006149f
C2809 VDD.n56 GND 0.006149f
C2810 VDD.n57 GND 0.006149f
C2811 VDD.n58 GND 0.006149f
C2812 VDD.n59 GND 0.006149f
C2813 VDD.n60 GND 0.004949f
C2814 VDD.n61 GND 0.006149f
C2815 VDD.n62 GND 0.006149f
C2816 VDD.n63 GND 0.006149f
C2817 VDD.n64 GND 0.006149f
C2818 VDD.n65 GND 0.498548f
C2819 VDD.n66 GND 0.006149f
C2820 VDD.n67 GND 0.006149f
C2821 VDD.n68 GND 0.006149f
C2822 VDD.n69 GND 0.006149f
C2823 VDD.n70 GND 0.006149f
C2824 VDD.n71 GND 0.004949f
C2825 VDD.n72 GND 0.006149f
C2826 VDD.n73 GND 0.006149f
C2827 VDD.n74 GND 0.006149f
C2828 VDD.n75 GND 0.006149f
C2829 VDD.n76 GND 0.498548f
C2830 VDD.n77 GND 0.006149f
C2831 VDD.n78 GND 0.006149f
C2832 VDD.n79 GND 0.006149f
C2833 VDD.n80 GND 0.006149f
C2834 VDD.n81 GND 0.006149f
C2835 VDD.n82 GND 0.004949f
C2836 VDD.n83 GND 0.006149f
C2837 VDD.n84 GND 0.006149f
C2838 VDD.n85 GND 0.006149f
C2839 VDD.n86 GND 0.006149f
C2840 VDD.n87 GND 0.498548f
C2841 VDD.n88 GND 0.006149f
C2842 VDD.n89 GND 0.006149f
C2843 VDD.n90 GND 0.006149f
C2844 VDD.n91 GND 0.006149f
C2845 VDD.n92 GND 0.006149f
C2846 VDD.n93 GND 0.004949f
C2847 VDD.n94 GND 0.006149f
C2848 VDD.n95 GND 0.006149f
C2849 VDD.n96 GND 0.006149f
C2850 VDD.n97 GND 0.006149f
C2851 VDD.n98 GND 0.498548f
C2852 VDD.n99 GND 0.006149f
C2853 VDD.n100 GND 0.006149f
C2854 VDD.n101 GND 0.006149f
C2855 VDD.n102 GND 0.006149f
C2856 VDD.n103 GND 0.006149f
C2857 VDD.n104 GND 0.004949f
C2858 VDD.n105 GND 0.006149f
C2859 VDD.n106 GND 0.006149f
C2860 VDD.n107 GND 0.006149f
C2861 VDD.n108 GND 0.006149f
C2862 VDD.n109 GND 0.498548f
C2863 VDD.n110 GND 0.006149f
C2864 VDD.n111 GND 0.006149f
C2865 VDD.n112 GND 0.006149f
C2866 VDD.n113 GND 0.006149f
C2867 VDD.n114 GND 0.006149f
C2868 VDD.n115 GND 0.004949f
C2869 VDD.n116 GND 0.006149f
C2870 VDD.n117 GND 0.498548f
C2871 VDD.n118 GND 0.006149f
C2872 VDD.n119 GND 0.006149f
C2873 VDD.n120 GND 0.004949f
C2874 VDD.n121 GND 0.006149f
C2875 VDD.n122 GND 0.006149f
C2876 VDD.n123 GND 0.004949f
C2877 VDD.n124 GND 0.006149f
C2878 VDD.n125 GND 0.006149f
C2879 VDD.n126 GND 0.004949f
C2880 VDD.n127 GND 0.006149f
C2881 VDD.n128 GND 0.006149f
C2882 VDD.n129 GND 0.004949f
C2883 VDD.n130 GND 0.006149f
C2884 VDD.n131 GND 0.006149f
C2885 VDD.n132 GND 0.004949f
C2886 VDD.n133 GND 0.006149f
C2887 VDD.n134 GND 0.006149f
C2888 VDD.n135 GND 0.004949f
C2889 VDD.n136 GND 0.006149f
C2890 VDD.n137 GND 0.006149f
C2891 VDD.n138 GND 0.004949f
C2892 VDD.n139 GND 0.006149f
C2893 VDD.n140 GND 0.004949f
C2894 VDD.n141 GND 0.006149f
C2895 VDD.n142 GND 0.004949f
C2896 VDD.n143 GND 0.006149f
C2897 VDD.n144 GND 0.006149f
C2898 VDD.n145 GND 0.498548f
C2899 VDD.n146 GND 0.006149f
C2900 VDD.n147 GND 0.004949f
C2901 VDD.n148 GND 0.006149f
C2902 VDD.n149 GND 0.004949f
C2903 VDD.n150 GND 0.006149f
C2904 VDD.n151 GND 0.498548f
C2905 VDD.n152 GND 0.006149f
C2906 VDD.n153 GND 0.004949f
C2907 VDD.n154 GND 0.006149f
C2908 VDD.n155 GND 0.004949f
C2909 VDD.n156 GND 0.006149f
C2910 VDD.t103 GND 0.249274f
C2911 VDD.n157 GND 0.006149f
C2912 VDD.n158 GND 0.004949f
C2913 VDD.n159 GND 0.006149f
C2914 VDD.n160 GND 0.004949f
C2915 VDD.n161 GND 0.006149f
C2916 VDD.n162 GND 0.498548f
C2917 VDD.n163 GND 0.006149f
C2918 VDD.n164 GND 0.004949f
C2919 VDD.n165 GND 0.006149f
C2920 VDD.n166 GND 0.004949f
C2921 VDD.n167 GND 0.006149f
C2922 VDD.n168 GND 0.498548f
C2923 VDD.n169 GND 0.006149f
C2924 VDD.n170 GND 0.004949f
C2925 VDD.n171 GND 0.006149f
C2926 VDD.n172 GND 0.004949f
C2927 VDD.n173 GND 0.006149f
C2928 VDD.n174 GND 0.498548f
C2929 VDD.n175 GND 0.006149f
C2930 VDD.n176 GND 0.004949f
C2931 VDD.n177 GND 0.006149f
C2932 VDD.n178 GND 0.004949f
C2933 VDD.n179 GND 0.006149f
C2934 VDD.n180 GND 0.498548f
C2935 VDD.n181 GND 0.006149f
C2936 VDD.n182 GND 0.004949f
C2937 VDD.n183 GND 0.006149f
C2938 VDD.n184 GND 0.004949f
C2939 VDD.n185 GND 0.006149f
C2940 VDD.n186 GND 0.498548f
C2941 VDD.n187 GND 0.006149f
C2942 VDD.n188 GND 0.004949f
C2943 VDD.n189 GND 0.006149f
C2944 VDD.n190 GND 0.004949f
C2945 VDD.n191 GND 0.006149f
C2946 VDD.t79 GND 0.249274f
C2947 VDD.n192 GND 0.006149f
C2948 VDD.n193 GND 0.004949f
C2949 VDD.n194 GND 0.006149f
C2950 VDD.n195 GND 0.004949f
C2951 VDD.n196 GND 0.006149f
C2952 VDD.n197 GND 0.498548f
C2953 VDD.n198 GND 0.006149f
C2954 VDD.n199 GND 0.004949f
C2955 VDD.n200 GND 0.006149f
C2956 VDD.n201 GND 0.004949f
C2957 VDD.n202 GND 0.006149f
C2958 VDD.n203 GND 0.498548f
C2959 VDD.n204 GND 0.006149f
C2960 VDD.n205 GND 0.004949f
C2961 VDD.n206 GND 0.006149f
C2962 VDD.n207 GND 0.004949f
C2963 VDD.n208 GND 0.006149f
C2964 VDD.n209 GND 0.498548f
C2965 VDD.n210 GND 0.006149f
C2966 VDD.n211 GND 0.004949f
C2967 VDD.n212 GND 0.006149f
C2968 VDD.n213 GND 0.004949f
C2969 VDD.n214 GND 0.006149f
C2970 VDD.n215 GND 0.498548f
C2971 VDD.n216 GND 0.006149f
C2972 VDD.n217 GND 0.004949f
C2973 VDD.n218 GND 0.006149f
C2974 VDD.n219 GND 0.004949f
C2975 VDD.n220 GND 0.006149f
C2976 VDD.n221 GND 0.498548f
C2977 VDD.n222 GND 0.006149f
C2978 VDD.n223 GND 0.004949f
C2979 VDD.n224 GND 0.006149f
C2980 VDD.n225 GND 0.004949f
C2981 VDD.n226 GND 0.006149f
C2982 VDD.n227 GND 0.498548f
C2983 VDD.n228 GND 0.006149f
C2984 VDD.n229 GND 0.004949f
C2985 VDD.n230 GND 0.006149f
C2986 VDD.n231 GND 0.004949f
C2987 VDD.n232 GND 0.006149f
C2988 VDD.n233 GND 0.498548f
C2989 VDD.n234 GND 0.006149f
C2990 VDD.n235 GND 0.004949f
C2991 VDD.n236 GND 0.006149f
C2992 VDD.n237 GND 0.004949f
C2993 VDD.n238 GND 0.006149f
C2994 VDD.n239 GND 0.498548f
C2995 VDD.n240 GND 0.006149f
C2996 VDD.n241 GND 0.004949f
C2997 VDD.n242 GND 0.006149f
C2998 VDD.n243 GND 0.004949f
C2999 VDD.n244 GND 0.006149f
C3000 VDD.n245 GND 0.498548f
C3001 VDD.n246 GND 0.006149f
C3002 VDD.n247 GND 0.004949f
C3003 VDD.n248 GND 0.006149f
C3004 VDD.n249 GND 0.004949f
C3005 VDD.n250 GND 0.006149f
C3006 VDD.n251 GND 0.498548f
C3007 VDD.n252 GND 0.006149f
C3008 VDD.n253 GND 0.004949f
C3009 VDD.n254 GND 0.006149f
C3010 VDD.n255 GND 0.004949f
C3011 VDD.n256 GND 0.006149f
C3012 VDD.n257 GND 0.498548f
C3013 VDD.n258 GND 0.006149f
C3014 VDD.n259 GND 0.004949f
C3015 VDD.n260 GND 0.006149f
C3016 VDD.n261 GND 0.004949f
C3017 VDD.n262 GND 0.006149f
C3018 VDD.n263 GND 0.498548f
C3019 VDD.n264 GND 0.006149f
C3020 VDD.n265 GND 0.004949f
C3021 VDD.n266 GND 0.006149f
C3022 VDD.n267 GND 0.004949f
C3023 VDD.n268 GND 0.006149f
C3024 VDD.t10 GND 0.249274f
C3025 VDD.n269 GND 0.006149f
C3026 VDD.n270 GND 0.004949f
C3027 VDD.n271 GND 0.006149f
C3028 VDD.n272 GND 0.004949f
C3029 VDD.n273 GND 0.006149f
C3030 VDD.n274 GND 0.498548f
C3031 VDD.n275 GND 0.339013f
C3032 VDD.n276 GND 0.006149f
C3033 VDD.n277 GND 0.004949f
C3034 VDD.n278 GND 0.006149f
C3035 VDD.n279 GND 0.004949f
C3036 VDD.n280 GND 0.006149f
C3037 VDD.n281 GND 0.498548f
C3038 VDD.n282 GND 0.006149f
C3039 VDD.n283 GND 0.004949f
C3040 VDD.n284 GND 0.012337f
C3041 VDD.n285 GND 0.004108f
C3042 VDD.n286 GND 0.013778f
C3043 VDD.n287 GND 0.695475f
C3044 VDD.n288 GND 0.013778f
C3045 VDD.n289 GND 0.004108f
C3046 VDD.n290 GND 0.05129f
C3047 VDD.n291 GND 0.004005f
C3048 VDD.n293 GND 0.006149f
C3049 VDD.n294 GND 0.004949f
C3050 VDD.n295 GND 0.004949f
C3051 VDD.n296 GND 0.006149f
C3052 VDD.n297 GND 0.006149f
C3053 VDD.t0 GND 6.15957f
C3054 VDD.n319 GND 0.006149f
C3055 VDD.n320 GND 0.004182f
C3056 VDD.n321 GND 0.004182f
C3057 VDD.t144 GND 4.95308f
C3058 VDD.n323 GND 2.17866f
C3059 VDD.n324 GND 0.004182f
C3060 VDD.n325 GND 0.004182f
C3061 VDD.n327 GND 0.004182f
C3062 VDD.t59 GND 0.18185f
C3063 VDD.t57 GND 0.551129f
C3064 VDD.n328 GND 0.095638f
C3065 VDD.t60 GND 0.141776f
C3066 VDD.n329 GND 0.095144f
C3067 VDD.n330 GND 0.005159f
C3068 VDD.n332 GND 0.002521f
C3069 VDD.n333 GND 0.004182f
C3070 VDD.n334 GND 0.009844f
C3071 VDD.n336 GND 0.004182f
C3072 VDD.n337 GND 0.339013f
C3073 VDD.n338 GND 0.009324f
C3074 VDD.t130 GND 0.276694f
C3075 VDD.n339 GND 0.009324f
C3076 VDD.n340 GND 0.004182f
C3077 VDD.n341 GND 0.009616f
C3078 VDD.n342 GND 0.004182f
C3079 VDD.n343 GND 0.004182f
C3080 VDD.n344 GND 0.004182f
C3081 VDD.n345 GND 0.004182f
C3082 VDD.n346 GND 0.004182f
C3083 VDD.n348 GND 0.004182f
C3084 VDD.n349 GND 0.004182f
C3085 VDD.n351 GND 0.004182f
C3086 VDD.n352 GND 0.004182f
C3087 VDD.n353 GND 0.004182f
C3088 VDD.n355 GND 0.004182f
C3089 VDD.t62 GND 0.18185f
C3090 VDD.t61 GND 0.551129f
C3091 VDD.n356 GND 0.095638f
C3092 VDD.t63 GND 0.141776f
C3093 VDD.n357 GND 0.095144f
C3094 VDD.n358 GND 0.005159f
C3095 VDD.n360 GND 0.002521f
C3096 VDD.n361 GND 0.004182f
C3097 VDD.n362 GND 0.004182f
C3098 VDD.n363 GND 0.004182f
C3099 VDD.n364 GND 0.339013f
C3100 VDD.n365 GND 0.004182f
C3101 VDD.n366 GND 0.004182f
C3102 VDD.n367 GND 0.004182f
C3103 VDD.n368 GND 0.004182f
C3104 VDD.n369 GND 0.004182f
C3105 VDD.n370 GND 0.339013f
C3106 VDD.n371 GND 0.004182f
C3107 VDD.n372 GND 0.004182f
C3108 VDD.n373 GND 0.004182f
C3109 VDD.n374 GND 0.004182f
C3110 VDD.n375 GND 0.004182f
C3111 VDD.n376 GND 0.004182f
C3112 VDD.n377 GND 0.339013f
C3113 VDD.n378 GND 0.004182f
C3114 VDD.n379 GND 0.004182f
C3115 VDD.n380 GND 0.004182f
C3116 VDD.n381 GND 0.004182f
C3117 VDD.n382 GND 0.004182f
C3118 VDD.t58 GND 0.169506f
C3119 VDD.n383 GND 0.004182f
C3120 VDD.n384 GND 0.004182f
C3121 VDD.n385 GND 0.004182f
C3122 VDD.n386 GND 0.004182f
C3123 VDD.n387 GND 0.004182f
C3124 VDD.n388 GND 0.319071f
C3125 VDD.n389 GND 0.004182f
C3126 VDD.n390 GND 0.004182f
C3127 VDD.n391 GND 0.306607f
C3128 VDD.n392 GND 0.004182f
C3129 VDD.n393 GND 0.004182f
C3130 VDD.n394 GND 0.004182f
C3131 VDD.n395 GND 0.339013f
C3132 VDD.n396 GND 0.004182f
C3133 VDD.n397 GND 0.004182f
C3134 VDD.t148 GND 0.169506f
C3135 VDD.n398 GND 0.004182f
C3136 VDD.n399 GND 0.004182f
C3137 VDD.n400 GND 0.004182f
C3138 VDD.n401 GND 0.339013f
C3139 VDD.n402 GND 0.004182f
C3140 VDD.n403 GND 0.004182f
C3141 VDD.n404 GND 0.004182f
C3142 VDD.n405 GND 0.004182f
C3143 VDD.n406 GND 0.004182f
C3144 VDD.n407 GND 0.339013f
C3145 VDD.n408 GND 0.004182f
C3146 VDD.n409 GND 0.004182f
C3147 VDD.n410 GND 0.004182f
C3148 VDD.n411 GND 0.004182f
C3149 VDD.n412 GND 0.004182f
C3150 VDD.n413 GND 0.339013f
C3151 VDD.n414 GND 0.004182f
C3152 VDD.n415 GND 0.004182f
C3153 VDD.n416 GND 0.004182f
C3154 VDD.n417 GND 0.004182f
C3155 VDD.n418 GND 0.004182f
C3156 VDD.n419 GND 0.339013f
C3157 VDD.n420 GND 0.004182f
C3158 VDD.n421 GND 0.004182f
C3159 VDD.n422 GND 0.004182f
C3160 VDD.n423 GND 0.004182f
C3161 VDD.n424 GND 0.004182f
C3162 VDD.n425 GND 0.339013f
C3163 VDD.n426 GND 0.004182f
C3164 VDD.n427 GND 0.004182f
C3165 VDD.n428 GND 0.004182f
C3166 VDD.n429 GND 0.004182f
C3167 VDD.n430 GND 0.004182f
C3168 VDD.t118 GND 0.169506f
C3169 VDD.n431 GND 0.004182f
C3170 VDD.n432 GND 0.004182f
C3171 VDD.n433 GND 0.004182f
C3172 VDD.n434 GND 0.004182f
C3173 VDD.n435 GND 0.004182f
C3174 VDD.n436 GND 0.339013f
C3175 VDD.n437 GND 0.004182f
C3176 VDD.n438 GND 0.004182f
C3177 VDD.t139 GND 0.169506f
C3178 VDD.n439 GND 0.004182f
C3179 VDD.n440 GND 0.004182f
C3180 VDD.n441 GND 0.004182f
C3181 VDD.n442 GND 0.339013f
C3182 VDD.n443 GND 0.004182f
C3183 VDD.n444 GND 0.004182f
C3184 VDD.n445 GND 0.004182f
C3185 VDD.n446 GND 0.004182f
C3186 VDD.n447 GND 0.004182f
C3187 VDD.n448 GND 0.339013f
C3188 VDD.n449 GND 0.004182f
C3189 VDD.n450 GND 0.004182f
C3190 VDD.n451 GND 0.004182f
C3191 VDD.n452 GND 0.004182f
C3192 VDD.n453 GND 0.004182f
C3193 VDD.n454 GND 0.339013f
C3194 VDD.n455 GND 0.004182f
C3195 VDD.n456 GND 0.004182f
C3196 VDD.n457 GND 0.004182f
C3197 VDD.n458 GND 0.004182f
C3198 VDD.n459 GND 0.004182f
C3199 VDD.n460 GND 0.339013f
C3200 VDD.n461 GND 0.004182f
C3201 VDD.n462 GND 0.004182f
C3202 VDD.n463 GND 0.004182f
C3203 VDD.n464 GND 0.004182f
C3204 VDD.n465 GND 0.004182f
C3205 VDD.n466 GND 0.339013f
C3206 VDD.n467 GND 0.004182f
C3207 VDD.n468 GND 0.004182f
C3208 VDD.n469 GND 0.004182f
C3209 VDD.n470 GND 0.004182f
C3210 VDD.n471 GND 0.004182f
C3211 VDD.t127 GND 0.169506f
C3212 VDD.n472 GND 0.004182f
C3213 VDD.n473 GND 0.004182f
C3214 VDD.n474 GND 0.004182f
C3215 VDD.n475 GND 0.004182f
C3216 VDD.n476 GND 0.004182f
C3217 VDD.n477 GND 0.339013f
C3218 VDD.n478 GND 0.004182f
C3219 VDD.n479 GND 0.004182f
C3220 VDD.n480 GND 0.326549f
C3221 VDD.n481 GND 0.004182f
C3222 VDD.n482 GND 0.004182f
C3223 VDD.n483 GND 0.004182f
C3224 VDD.n484 GND 0.286665f
C3225 VDD.n485 GND 0.004182f
C3226 VDD.n486 GND 0.004182f
C3227 VDD.n487 GND 0.004182f
C3228 VDD.n488 GND 0.004182f
C3229 VDD.n489 GND 0.004182f
C3230 VDD.n490 GND 0.339013f
C3231 VDD.n491 GND 0.004182f
C3232 VDD.n492 GND 0.004182f
C3233 VDD.t121 GND 0.169506f
C3234 VDD.n493 GND 0.004182f
C3235 VDD.n494 GND 0.004182f
C3236 VDD.n495 GND 0.004182f
C3237 VDD.n496 GND 0.339013f
C3238 VDD.n497 GND 0.004182f
C3239 VDD.n498 GND 0.004182f
C3240 VDD.n499 GND 0.004182f
C3241 VDD.n500 GND 0.004182f
C3242 VDD.n501 GND 0.004182f
C3243 VDD.n502 GND 0.339013f
C3244 VDD.n503 GND 0.004182f
C3245 VDD.n504 GND 0.004182f
C3246 VDD.n505 GND 0.004182f
C3247 VDD.n506 GND 0.004182f
C3248 VDD.n507 GND 0.004182f
C3249 VDD.t120 GND 0.169506f
C3250 VDD.n508 GND 0.004182f
C3251 VDD.n509 GND 0.004182f
C3252 VDD.n510 GND 0.004182f
C3253 VDD.n511 GND 0.004182f
C3254 VDD.n512 GND 0.004182f
C3255 VDD.n513 GND 0.339013f
C3256 VDD.n514 GND 0.004182f
C3257 VDD.n515 GND 0.004182f
C3258 VDD.n516 GND 0.18197f
C3259 VDD.n517 GND 0.004182f
C3260 VDD.n518 GND 0.004182f
C3261 VDD.n519 GND 0.004182f
C3262 VDD.n520 GND 0.339013f
C3263 VDD.n521 GND 0.004182f
C3264 VDD.n522 GND 0.004182f
C3265 VDD.n523 GND 0.004182f
C3266 VDD.n524 GND 0.004182f
C3267 VDD.n525 GND 0.004182f
C3268 VDD.t150 GND 0.169506f
C3269 VDD.n526 GND 0.004182f
C3270 VDD.n527 GND 0.004182f
C3271 VDD.n528 GND 0.004182f
C3272 VDD.n529 GND 0.004182f
C3273 VDD.n530 GND 0.004182f
C3274 VDD.n531 GND 0.339013f
C3275 VDD.n532 GND 0.004182f
C3276 VDD.n533 GND 0.004182f
C3277 VDD.n534 GND 0.246781f
C3278 VDD.n535 GND 0.004182f
C3279 VDD.n536 GND 0.004182f
C3280 VDD.n537 GND 0.004182f
C3281 VDD.n538 GND 0.339013f
C3282 VDD.n539 GND 0.004182f
C3283 VDD.n540 GND 0.004182f
C3284 VDD.n541 GND 0.004182f
C3285 VDD.n542 GND 0.004182f
C3286 VDD.n543 GND 0.004182f
C3287 VDD.n544 GND 0.301622f
C3288 VDD.n545 GND 0.004182f
C3289 VDD.n546 GND 0.004182f
C3290 VDD.n547 GND 0.004182f
C3291 VDD.n548 GND 0.004182f
C3292 VDD.n549 GND 0.004182f
C3293 VDD.n550 GND 0.339013f
C3294 VDD.n551 GND 0.004182f
C3295 VDD.n552 GND 0.004182f
C3296 VDD.t136 GND 0.169506f
C3297 VDD.n553 GND 0.004182f
C3298 VDD.n554 GND 0.004182f
C3299 VDD.n555 GND 0.004182f
C3300 VDD.n556 GND 0.339013f
C3301 VDD.n557 GND 0.004182f
C3302 VDD.n558 GND 0.004182f
C3303 VDD.n559 GND 0.004182f
C3304 VDD.n560 GND 0.004182f
C3305 VDD.n561 GND 0.004182f
C3306 VDD.n562 GND 0.23681f
C3307 VDD.n563 GND 0.004182f
C3308 VDD.n564 GND 0.004182f
C3309 VDD.n565 GND 0.004182f
C3310 VDD.n566 GND 0.004182f
C3311 VDD.n567 GND 0.004182f
C3312 VDD.n568 GND 0.339013f
C3313 VDD.n569 GND 0.004182f
C3314 VDD.n570 GND 0.004182f
C3315 VDD.t125 GND 0.169506f
C3316 VDD.n571 GND 0.004182f
C3317 VDD.n572 GND 0.004182f
C3318 VDD.n573 GND 0.004182f
C3319 VDD.n574 GND 0.339013f
C3320 VDD.n575 GND 0.004182f
C3321 VDD.n576 GND 0.004182f
C3322 VDD.n577 GND 0.004182f
C3323 VDD.n578 GND 0.004182f
C3324 VDD.n579 GND 0.004182f
C3325 VDD.n580 GND 0.339013f
C3326 VDD.n581 GND 0.004182f
C3327 VDD.n582 GND 0.004182f
C3328 VDD.n583 GND 0.004182f
C3329 VDD.n584 GND 0.004182f
C3330 VDD.n585 GND 0.004182f
C3331 VDD.n586 GND 0.339013f
C3332 VDD.n587 GND 0.004182f
C3333 VDD.n588 GND 0.004182f
C3334 VDD.n589 GND 0.004182f
C3335 VDD.n590 GND 0.004182f
C3336 VDD.n591 GND 0.004182f
C3337 VDD.n592 GND 0.339013f
C3338 VDD.n593 GND 0.004182f
C3339 VDD.n594 GND 0.004182f
C3340 VDD.n595 GND 0.004182f
C3341 VDD.n596 GND 0.004182f
C3342 VDD.n597 GND 0.004182f
C3343 VDD.t48 GND 0.169506f
C3344 VDD.n598 GND 0.004182f
C3345 VDD.n599 GND 0.004182f
C3346 VDD.n600 GND 0.004182f
C3347 VDD.n601 GND 0.004182f
C3348 VDD.n602 GND 0.004182f
C3349 VDD.t134 GND 0.169506f
C3350 VDD.n603 GND 0.004182f
C3351 VDD.n604 GND 0.004182f
C3352 VDD.n605 GND 0.201912f
C3353 VDD.n606 GND 0.004182f
C3354 VDD.n607 GND 0.004182f
C3355 VDD.n608 GND 0.004182f
C3356 VDD.n609 GND 0.339013f
C3357 VDD.n610 GND 0.004182f
C3358 VDD.n611 GND 0.004182f
C3359 VDD.n612 GND 0.296636f
C3360 VDD.n613 GND 0.004182f
C3361 VDD.n614 GND 0.004182f
C3362 VDD.n615 GND 0.004182f
C3363 VDD.n616 GND 0.339013f
C3364 VDD.n617 GND 0.004182f
C3365 VDD.n618 GND 0.004182f
C3366 VDD.n619 GND 0.004182f
C3367 VDD.n620 GND 0.009324f
C3368 VDD.n621 GND 0.009324f
C3369 VDD.n622 GND 0.446201f
C3370 VDD.n623 GND 0.004182f
C3371 VDD.n624 GND 0.004182f
C3372 VDD.n625 GND 0.009324f
C3373 VDD.n626 GND 0.004182f
C3374 VDD.n627 GND 0.004182f
C3375 VDD.n628 GND 0.446201f
C3376 VDD.n641 GND 0.009616f
C3377 VDD.n654 GND 0.009324f
C3378 VDD.n655 GND 0.004182f
C3379 VDD.n656 GND 0.009324f
C3380 VDD.t19 GND 0.18185f
C3381 VDD.t17 GND 0.551129f
C3382 VDD.n657 GND 0.095638f
C3383 VDD.t20 GND 0.141776f
C3384 VDD.n658 GND 0.095144f
C3385 VDD.n659 GND 0.005159f
C3386 VDD.n660 GND 0.009844f
C3387 VDD.n661 GND 0.004182f
C3388 VDD.n662 GND 0.004182f
C3389 VDD.n663 GND 0.339013f
C3390 VDD.n664 GND 0.004182f
C3391 VDD.n665 GND 0.004182f
C3392 VDD.n666 GND 0.004182f
C3393 VDD.n667 GND 0.004182f
C3394 VDD.n668 GND 0.004182f
C3395 VDD.n669 GND 0.339013f
C3396 VDD.n670 GND 0.004182f
C3397 VDD.n671 GND 0.004182f
C3398 VDD.n672 GND 0.004182f
C3399 VDD.n673 GND 0.004182f
C3400 VDD.n674 GND 0.004182f
C3401 VDD.t32 GND 0.18185f
C3402 VDD.t31 GND 0.551129f
C3403 VDD.n675 GND 0.095638f
C3404 VDD.t33 GND 0.141776f
C3405 VDD.n676 GND 0.095144f
C3406 VDD.n677 GND 0.004182f
C3407 VDD.n678 GND 0.004182f
C3408 VDD.n679 GND 0.296636f
C3409 VDD.n680 GND 0.004182f
C3410 VDD.n681 GND 0.004182f
C3411 VDD.n682 GND 0.004182f
C3412 VDD.n683 GND 0.004182f
C3413 VDD.n684 GND 0.004182f
C3414 VDD.n685 GND 0.201912f
C3415 VDD.n686 GND 0.004182f
C3416 VDD.n687 GND 0.004182f
C3417 VDD.t152 GND 0.169506f
C3418 VDD.n688 GND 0.004182f
C3419 VDD.n689 GND 0.004182f
C3420 VDD.n690 GND 0.004182f
C3421 VDD.n691 GND 0.004182f
C3422 VDD.n692 GND 0.339013f
C3423 VDD.n693 GND 0.004182f
C3424 VDD.n694 GND 0.004182f
C3425 VDD.t18 GND 0.169506f
C3426 VDD.n695 GND 0.004182f
C3427 VDD.n696 GND 0.004182f
C3428 VDD.n697 GND 0.004182f
C3429 VDD.n698 GND 0.339013f
C3430 VDD.n699 GND 0.004182f
C3431 VDD.n700 GND 0.004182f
C3432 VDD.n701 GND 0.004182f
C3433 VDD.n702 GND 0.004182f
C3434 VDD.n703 GND 0.004182f
C3435 VDD.n704 GND 0.339013f
C3436 VDD.n705 GND 0.004182f
C3437 VDD.n706 GND 0.004182f
C3438 VDD.n707 GND 0.004182f
C3439 VDD.n708 GND 0.004182f
C3440 VDD.n709 GND 0.004182f
C3441 VDD.n710 GND 0.339013f
C3442 VDD.n711 GND 0.004182f
C3443 VDD.n712 GND 0.004182f
C3444 VDD.n713 GND 0.004182f
C3445 VDD.n714 GND 0.004182f
C3446 VDD.n715 GND 0.004182f
C3447 VDD.n716 GND 0.339013f
C3448 VDD.n717 GND 0.004182f
C3449 VDD.n718 GND 0.004182f
C3450 VDD.n719 GND 0.004182f
C3451 VDD.n720 GND 0.004182f
C3452 VDD.n721 GND 0.004182f
C3453 VDD.t132 GND 0.169506f
C3454 VDD.n722 GND 0.004182f
C3455 VDD.n723 GND 0.004182f
C3456 VDD.n724 GND 0.004182f
C3457 VDD.n725 GND 0.004182f
C3458 VDD.n726 GND 0.004182f
C3459 VDD.n727 GND 0.339013f
C3460 VDD.n728 GND 0.004182f
C3461 VDD.n729 GND 0.004182f
C3462 VDD.n730 GND 0.23681f
C3463 VDD.n731 GND 0.004182f
C3464 VDD.n732 GND 0.004182f
C3465 VDD.n733 GND 0.004182f
C3466 VDD.n734 GND 0.339013f
C3467 VDD.n735 GND 0.004182f
C3468 VDD.n736 GND 0.004182f
C3469 VDD.n737 GND 0.004182f
C3470 VDD.n738 GND 0.004182f
C3471 VDD.n739 GND 0.004182f
C3472 VDD.t142 GND 0.169506f
C3473 VDD.n740 GND 0.004182f
C3474 VDD.n741 GND 0.004182f
C3475 VDD.n742 GND 0.004182f
C3476 VDD.n743 GND 0.004182f
C3477 VDD.n744 GND 0.004182f
C3478 VDD.n745 GND 0.339013f
C3479 VDD.n746 GND 0.004182f
C3480 VDD.n747 GND 0.004182f
C3481 VDD.n748 GND 0.301622f
C3482 VDD.n749 GND 0.004182f
C3483 VDD.n750 GND 0.004182f
C3484 VDD.n751 GND 0.004182f
C3485 VDD.n752 GND 0.339013f
C3486 VDD.n753 GND 0.004182f
C3487 VDD.n754 GND 0.004182f
C3488 VDD.n755 GND 0.004182f
C3489 VDD.n756 GND 0.004182f
C3490 VDD.n757 GND 0.004182f
C3491 VDD.n758 GND 0.246781f
C3492 VDD.n759 GND 0.004182f
C3493 VDD.n760 GND 0.004182f
C3494 VDD.n761 GND 0.004182f
C3495 VDD.n762 GND 0.004182f
C3496 VDD.n763 GND 0.004182f
C3497 VDD.n764 GND 0.339013f
C3498 VDD.n765 GND 0.004182f
C3499 VDD.n766 GND 0.004182f
C3500 VDD.t156 GND 0.169506f
C3501 VDD.n767 GND 0.004182f
C3502 VDD.n768 GND 0.004182f
C3503 VDD.n769 GND 0.004182f
C3504 VDD.n770 GND 0.339013f
C3505 VDD.n771 GND 0.004182f
C3506 VDD.n772 GND 0.004182f
C3507 VDD.n773 GND 0.004182f
C3508 VDD.n774 GND 0.004182f
C3509 VDD.n775 GND 0.004182f
C3510 VDD.n776 GND 0.18197f
C3511 VDD.n777 GND 0.004182f
C3512 VDD.n778 GND 0.004182f
C3513 VDD.n779 GND 0.004182f
C3514 VDD.n780 GND 0.004182f
C3515 VDD.n781 GND 0.004182f
C3516 VDD.n782 GND 0.339013f
C3517 VDD.n783 GND 0.004182f
C3518 VDD.n784 GND 0.004182f
C3519 VDD.t124 GND 0.169506f
C3520 VDD.n785 GND 0.004182f
C3521 VDD.n786 GND 0.004182f
C3522 VDD.n787 GND 0.004182f
C3523 VDD.n788 GND 0.339013f
C3524 VDD.n789 GND 0.004182f
C3525 VDD.n790 GND 0.004182f
C3526 VDD.n791 GND 0.004182f
C3527 VDD.n792 GND 0.004182f
C3528 VDD.n793 GND 0.004182f
C3529 VDD.n794 GND 0.339013f
C3530 VDD.n795 GND 0.004182f
C3531 VDD.n796 GND 0.004182f
C3532 VDD.n797 GND 0.004182f
C3533 VDD.n798 GND 0.004182f
C3534 VDD.n799 GND 0.004182f
C3535 VDD.t146 GND 0.169506f
C3536 VDD.n800 GND 0.004182f
C3537 VDD.n801 GND 0.004182f
C3538 VDD.n802 GND 0.004182f
C3539 VDD.n803 GND 0.004182f
C3540 VDD.n804 GND 0.004182f
C3541 VDD.n805 GND 0.339013f
C3542 VDD.n806 GND 0.004182f
C3543 VDD.n807 GND 0.004182f
C3544 VDD.n808 GND 0.286665f
C3545 VDD.n809 GND 0.004182f
C3546 VDD.n810 GND 0.004182f
C3547 VDD.n811 GND 0.004182f
C3548 VDD.n812 GND 0.326549f
C3549 VDD.n813 GND 0.004182f
C3550 VDD.n814 GND 0.004182f
C3551 VDD.n815 GND 0.004182f
C3552 VDD.n816 GND 0.004182f
C3553 VDD.n817 GND 0.004182f
C3554 VDD.n818 GND 0.339013f
C3555 VDD.n819 GND 0.004182f
C3556 VDD.n820 GND 0.004182f
C3557 VDD.t123 GND 0.169506f
C3558 VDD.n821 GND 0.004182f
C3559 VDD.n822 GND 0.004182f
C3560 VDD.n823 GND 0.004182f
C3561 VDD.n824 GND 0.339013f
C3562 VDD.n825 GND 0.004182f
C3563 VDD.n826 GND 0.004182f
C3564 VDD.n827 GND 0.004182f
C3565 VDD.n828 GND 0.004182f
C3566 VDD.n829 GND 0.004182f
C3567 VDD.n830 GND 0.339013f
C3568 VDD.n831 GND 0.004182f
C3569 VDD.n832 GND 0.004182f
C3570 VDD.n833 GND 0.004182f
C3571 VDD.n834 GND 0.004182f
C3572 VDD.n835 GND 0.004182f
C3573 VDD.n836 GND 0.339013f
C3574 VDD.n837 GND 0.004182f
C3575 VDD.n838 GND 0.004182f
C3576 VDD.n839 GND 0.004182f
C3577 VDD.n840 GND 0.004182f
C3578 VDD.n841 GND 0.004182f
C3579 VDD.n842 GND 0.339013f
C3580 VDD.n843 GND 0.004182f
C3581 VDD.n844 GND 0.004182f
C3582 VDD.n845 GND 0.004182f
C3583 VDD.n846 GND 0.004182f
C3584 VDD.n847 GND 0.004182f
C3585 VDD.n848 GND 0.339013f
C3586 VDD.n849 GND 0.004182f
C3587 VDD.n850 GND 0.004182f
C3588 VDD.n851 GND 0.004182f
C3589 VDD.n852 GND 0.004182f
C3590 VDD.n853 GND 0.004182f
C3591 VDD.t143 GND 0.169506f
C3592 VDD.n854 GND 0.004182f
C3593 VDD.n855 GND 0.004182f
C3594 VDD.n856 GND 0.004182f
C3595 VDD.n857 GND 0.004182f
C3596 VDD.n858 GND 0.004182f
C3597 VDD.n859 GND 0.339013f
C3598 VDD.n860 GND 0.004182f
C3599 VDD.n861 GND 0.004182f
C3600 VDD.t137 GND 0.169506f
C3601 VDD.n862 GND 0.004182f
C3602 VDD.n863 GND 0.004182f
C3603 VDD.n864 GND 0.004182f
C3604 VDD.n865 GND 0.339013f
C3605 VDD.n866 GND 0.004182f
C3606 VDD.n867 GND 0.004182f
C3607 VDD.n868 GND 0.004182f
C3608 VDD.n869 GND 0.004182f
C3609 VDD.n870 GND 0.004182f
C3610 VDD.n871 GND 0.339013f
C3611 VDD.n872 GND 0.004182f
C3612 VDD.n873 GND 0.004182f
C3613 VDD.n874 GND 0.004182f
C3614 VDD.n875 GND 0.004182f
C3615 VDD.n876 GND 0.004182f
C3616 VDD.n877 GND 0.339013f
C3617 VDD.n878 GND 0.004182f
C3618 VDD.n879 GND 0.004182f
C3619 VDD.n880 GND 0.004182f
C3620 VDD.n881 GND 0.004182f
C3621 VDD.n882 GND 0.004182f
C3622 VDD.n883 GND 0.339013f
C3623 VDD.n884 GND 0.004182f
C3624 VDD.n885 GND 0.004182f
C3625 VDD.n886 GND 0.004182f
C3626 VDD.n887 GND 0.004182f
C3627 VDD.n888 GND 0.004182f
C3628 VDD.n889 GND 0.339013f
C3629 VDD.n890 GND 0.004182f
C3630 VDD.n891 GND 0.004182f
C3631 VDD.n892 GND 0.004182f
C3632 VDD.n893 GND 0.004182f
C3633 VDD.n894 GND 0.004182f
C3634 VDD.t154 GND 0.169506f
C3635 VDD.n895 GND 0.004182f
C3636 VDD.n896 GND 0.004182f
C3637 VDD.n897 GND 0.004182f
C3638 VDD.n898 GND 0.004182f
C3639 VDD.n899 GND 0.004182f
C3640 VDD.n900 GND 0.306607f
C3641 VDD.n901 GND 0.004182f
C3642 VDD.n902 GND 0.004182f
C3643 VDD.n903 GND 0.319071f
C3644 VDD.n904 GND 0.004182f
C3645 VDD.n905 GND 0.004182f
C3646 VDD.n906 GND 0.004182f
C3647 VDD.n907 GND 0.339013f
C3648 VDD.n908 GND 0.004182f
C3649 VDD.n909 GND 0.004182f
C3650 VDD.t41 GND 0.169506f
C3651 VDD.n910 GND 0.004182f
C3652 VDD.n911 GND 0.004182f
C3653 VDD.n912 GND 0.004182f
C3654 VDD.n913 GND 0.339013f
C3655 VDD.n914 GND 0.004182f
C3656 VDD.n915 GND 0.004182f
C3657 VDD.n916 GND 0.004182f
C3658 VDD.n917 GND 0.004182f
C3659 VDD.n918 GND 0.004182f
C3660 VDD.n919 GND 0.339013f
C3661 VDD.n920 GND 0.004182f
C3662 VDD.n921 GND 0.004182f
C3663 VDD.n922 GND 0.004182f
C3664 VDD.n923 GND 0.004182f
C3665 VDD.n924 GND 0.004182f
C3666 VDD.n925 GND 0.339013f
C3667 VDD.n926 GND 0.004182f
C3668 VDD.n927 GND 0.004182f
C3669 VDD.n928 GND 0.004182f
C3670 VDD.n929 GND 0.009616f
C3671 VDD.n930 GND 0.009616f
C3672 VDD.t140 GND 0.276694f
C3673 VDD.n931 GND 0.009324f
C3674 VDD.n932 GND 0.009324f
C3675 VDD.n933 GND 0.009616f
C3676 VDD.n934 GND 0.004182f
C3677 VDD.n935 GND 0.004182f
C3678 VDD.t128 GND 4.95308f
C3679 VDD.n959 GND 0.004182f
C3680 VDD.n960 GND 0.004182f
C3681 VDD.n961 GND 0.004182f
C3682 VDD.n962 GND 0.004182f
C3683 VDD.n963 GND 0.004182f
C3684 VDD.n964 GND 0.004182f
C3685 VDD.n965 GND 0.004182f
C3686 VDD.n966 GND 0.004182f
C3687 VDD.n967 GND 0.004182f
C3688 VDD.n968 GND 0.004182f
C3689 VDD.n969 GND 0.004182f
C3690 VDD.n970 GND 0.004182f
C3691 VDD.n971 GND 0.004182f
C3692 VDD.n972 GND 0.004182f
C3693 VDD.n973 GND 0.004182f
C3694 VDD.n974 GND 0.004182f
C3695 VDD.n975 GND 0.004182f
C3696 VDD.n976 GND 0.004182f
C3697 VDD.n977 GND 0.004182f
C3698 VDD.n978 GND 0.004182f
C3699 VDD.n979 GND 0.004182f
C3700 VDD.n980 GND 0.004182f
C3701 VDD.n981 GND 0.004182f
C3702 VDD.n982 GND 0.004182f
C3703 VDD.n983 GND 0.004182f
C3704 VDD.n984 GND 0.004182f
C3705 VDD.n985 GND 0.004182f
C3706 VDD.n986 GND 0.004182f
C3707 VDD.n987 GND 0.004182f
C3708 VDD.n988 GND 0.004182f
C3709 VDD.n989 GND 0.004182f
C3710 VDD.n990 GND 0.004182f
C3711 VDD.n991 GND 0.004182f
C3712 VDD.n992 GND 0.004182f
C3713 VDD.n993 GND 0.004182f
C3714 VDD.n994 GND 0.004182f
C3715 VDD.n995 GND 0.004182f
C3716 VDD.n996 GND 0.004182f
C3717 VDD.n997 GND 0.004182f
C3718 VDD.n998 GND 0.004182f
C3719 VDD.n999 GND 0.004182f
C3720 VDD.n1000 GND 0.004182f
C3721 VDD.n1001 GND 0.004182f
C3722 VDD.n1002 GND 0.004182f
C3723 VDD.n1003 GND 0.004182f
C3724 VDD.n1004 GND 0.004182f
C3725 VDD.n1005 GND 0.004182f
C3726 VDD.n1006 GND 0.004182f
C3727 VDD.n1007 GND 0.004182f
C3728 VDD.n1008 GND 0.004182f
C3729 VDD.n1009 GND 0.004182f
C3730 VDD.n1010 GND 0.004182f
C3731 VDD.n1011 GND 0.004182f
C3732 VDD.n1012 GND 0.004182f
C3733 VDD.n1013 GND 0.004182f
C3734 VDD.n1014 GND 0.004182f
C3735 VDD.n1015 GND 0.004182f
C3736 VDD.n1016 GND 0.004182f
C3737 VDD.n1017 GND 0.004182f
C3738 VDD.n1018 GND 0.004182f
C3739 VDD.n1019 GND 0.004182f
C3740 VDD.n1020 GND 0.004182f
C3741 VDD.n1021 GND 0.004182f
C3742 VDD.n1022 GND 0.004182f
C3743 VDD.n1023 GND 0.004182f
C3744 VDD.n1024 GND 0.004182f
C3745 VDD.n1025 GND 0.004182f
C3746 VDD.n1026 GND 0.004182f
C3747 VDD.n1027 GND 0.004182f
C3748 VDD.n1028 GND 0.004182f
C3749 VDD.n1029 GND 0.004182f
C3750 VDD.n1030 GND 0.004182f
C3751 VDD.n1031 GND 0.004182f
C3752 VDD.n1032 GND 0.004182f
C3753 VDD.n1033 GND 0.004182f
C3754 VDD.n1034 GND 0.004182f
C3755 VDD.n1035 GND 0.004182f
C3756 VDD.n1036 GND 0.004182f
C3757 VDD.n1037 GND 0.004182f
C3758 VDD.n1038 GND 0.004182f
C3759 VDD.n1039 GND 0.004182f
C3760 VDD.n1040 GND 0.004182f
C3761 VDD.n1041 GND 0.004182f
C3762 VDD.n1042 GND 0.004182f
C3763 VDD.n1043 GND 0.004182f
C3764 VDD.n1044 GND 0.004182f
C3765 VDD.n1045 GND 0.004182f
C3766 VDD.n1046 GND 0.004182f
C3767 VDD.t43 GND 0.18185f
C3768 VDD.t40 GND 0.551129f
C3769 VDD.n1047 GND 0.095638f
C3770 VDD.t42 GND 0.141776f
C3771 VDD.n1048 GND 0.095144f
C3772 VDD.n1049 GND 0.005159f
C3773 VDD.n1050 GND 0.004182f
C3774 VDD.n1051 GND 0.004182f
C3775 VDD.n1052 GND 0.004182f
C3776 VDD.n1053 GND 0.004182f
C3777 VDD.n1054 GND 0.004182f
C3778 VDD.n1055 GND 0.004182f
C3779 VDD.n1056 GND 0.004182f
C3780 VDD.n1057 GND 0.004182f
C3781 VDD.n1058 GND 0.004182f
C3782 VDD.n1059 GND 0.004182f
C3783 VDD.n1060 GND 0.004182f
C3784 VDD.n1061 GND 0.004182f
C3785 VDD.n1062 GND 0.004182f
C3786 VDD.n1063 GND 0.004182f
C3787 VDD.n1064 GND 0.004182f
C3788 VDD.n1065 GND 0.004182f
C3789 VDD.n1066 GND 0.004182f
C3790 VDD.n1067 GND 0.004182f
C3791 VDD.n1068 GND 0.004305f
C3792 VDD.n1070 GND 0.004005f
C3793 VDD.n1071 GND 0.006149f
C3794 VDD.n1072 GND 0.004949f
C3795 VDD.n1073 GND 0.006149f
C3796 VDD.n1074 GND 0.014243f
C3797 VDD.n1075 GND 0.498548f
C3798 VDD.n1076 GND 0.013778f
C3799 VDD.t1 GND 6.15957f
C3800 VDD.n1100 GND 0.006149f
C3801 VDD.n1101 GND 0.006149f
C3802 VDD.n1102 GND 0.006149f
C3803 VDD.n1103 GND 0.006149f
C3804 VDD.n1104 GND 0.006149f
C3805 VDD.n1105 GND 0.006149f
C3806 VDD.n1106 GND 0.006149f
C3807 VDD.n1107 GND 0.006149f
C3808 VDD.n1108 GND 0.006149f
C3809 VDD.n1109 GND 0.006149f
C3810 VDD.n1110 GND 0.003984f
C3811 VDD.t4 GND 0.179673f
C3812 VDD.t2 GND 0.743196f
C3813 VDD.n1111 GND 0.095879f
C3814 VDD.t5 GND 0.131174f
C3815 VDD.n1112 GND 0.098395f
C3816 VDD.n1113 GND 0.006149f
C3817 VDD.n1114 GND 0.006149f
C3818 VDD.n1115 GND 0.006149f
C3819 VDD.n1116 GND 0.006149f
C3820 VDD.n1117 GND 0.006149f
C3821 VDD.n1118 GND 0.006149f
C3822 VDD.n1119 GND 0.006149f
C3823 VDD.n1120 GND 0.006149f
C3824 VDD.n1121 GND 0.006149f
C3825 VDD.n1122 GND 0.006149f
C3826 VDD.n1123 GND 0.006149f
C3827 VDD.n1124 GND 0.006149f
C3828 VDD.n1125 GND 0.006149f
C3829 VDD.n1126 GND 0.006149f
C3830 VDD.n1127 GND 0.006149f
C3831 VDD.n1128 GND 0.006149f
C3832 VDD.t7 GND 0.179673f
C3833 VDD.t6 GND 0.743196f
C3834 VDD.n1129 GND 0.095879f
C3835 VDD.t8 GND 0.131174f
C3836 VDD.n1130 GND 0.098395f
C3837 VDD.n1131 GND 0.006806f
C3838 VDD.n1132 GND 0.006149f
C3839 VDD.n1133 GND 0.006149f
C3840 VDD.n1134 GND 0.006149f
C3841 VDD.n1135 GND 0.006149f
C3842 VDD.n1136 GND 0.006149f
C3843 VDD.n1137 GND 0.006149f
C3844 VDD.n1138 GND 0.006149f
C3845 VDD.n1139 GND 0.006149f
C3846 VDD.n1140 GND 0.006149f
C3847 VDD.n1141 GND 0.006149f
C3848 VDD.n1142 GND 0.006149f
C3849 VDD.n1143 GND 0.006149f
C3850 VDD.n1144 GND 0.006149f
C3851 VDD.n1145 GND 0.004305f
C3852 VDD.n1146 GND 0.004628f
C3853 VDD.n1147 GND 0.004182f
C3854 VDD.n1148 GND 0.004182f
C3855 VDD.n1149 GND 0.004182f
C3856 VDD.n1150 GND 0.004182f
C3857 VDD.n1151 GND 0.004182f
C3858 VDD.n1152 GND 0.004182f
C3859 VDD.n1153 GND 0.004182f
C3860 VDD.n1154 GND 0.004182f
C3861 VDD.n1155 GND 0.004182f
C3862 VDD.n1156 GND 0.004182f
C3863 VDD.n1157 GND 0.004182f
C3864 VDD.n1158 GND 0.004182f
C3865 VDD.n1159 GND 0.004182f
C3866 VDD.n1160 GND 0.004182f
C3867 VDD.n1161 GND 0.004182f
C3868 VDD.n1162 GND 0.004182f
C3869 VDD.n1163 GND 0.004182f
C3870 VDD.n1164 GND 0.004182f
C3871 VDD.n1165 GND 0.004182f
C3872 VDD.n1166 GND 0.004182f
C3873 VDD.n1167 GND 0.004182f
C3874 VDD.n1168 GND 0.004182f
C3875 VDD.n1169 GND 0.004182f
C3876 VDD.t56 GND 0.18185f
C3877 VDD.t54 GND 0.551129f
C3878 VDD.n1170 GND 0.095638f
C3879 VDD.t55 GND 0.141776f
C3880 VDD.n1171 GND 0.095144f
C3881 VDD.n1172 GND 0.004182f
C3882 VDD.n1173 GND 0.004182f
C3883 VDD.n1174 GND 0.004182f
C3884 VDD.n1175 GND 0.002521f
C3885 VDD.n1176 GND 0.005159f
C3886 VDD.n1177 GND 0.003751f
C3887 VDD.n1178 GND 0.004182f
C3888 VDD.n1179 GND 0.004182f
C3889 VDD.n1180 GND 0.004182f
C3890 VDD.n1181 GND 0.004182f
C3891 VDD.n1182 GND 0.004182f
C3892 VDD.n1183 GND 0.004182f
C3893 VDD.n1184 GND 0.004182f
C3894 VDD.n1185 GND 0.004182f
C3895 VDD.n1186 GND 0.004182f
C3896 VDD.n1187 GND 0.004182f
C3897 VDD.n1188 GND 0.004182f
C3898 VDD.n1189 GND 0.004182f
C3899 VDD.n1190 GND 0.004182f
C3900 VDD.n1191 GND 0.004182f
C3901 VDD.n1192 GND 0.004182f
C3902 VDD.n1193 GND 0.053563f
C3903 VDD.n1194 GND 0.014186f
C3904 VDD.t45 GND 0.179673f
C3905 VDD.t44 GND 0.743196f
C3906 VDD.n1195 GND 0.095879f
C3907 VDD.t46 GND 0.131174f
C3908 VDD.n1196 GND 0.098395f
C3909 VDD.n1197 GND 0.006149f
C3910 VDD.n1198 GND 0.006149f
C3911 VDD.n1199 GND 0.00928f
C3912 VDD.n1200 GND 0.002751f
C3913 VDD.n1201 GND 0.006149f
C3914 VDD.n1202 GND 0.004949f
C3915 VDD.n1203 GND 0.006149f
C3916 VDD.n1204 GND 0.498548f
C3917 VDD.n1205 GND 0.006149f
C3918 VDD.n1206 GND 0.004949f
C3919 VDD.n1207 GND 0.006149f
C3920 VDD.n1208 GND 0.004949f
C3921 VDD.n1209 GND 0.006149f
C3922 VDD.n1210 GND 0.498548f
C3923 VDD.n1211 GND 0.006149f
C3924 VDD.n1212 GND 0.004949f
C3925 VDD.n1213 GND 0.004949f
C3926 VDD.n1214 GND 0.006149f
C3927 VDD.n1215 GND 0.004949f
C3928 VDD.n1216 GND 0.006149f
C3929 VDD.t3 GND 0.249274f
C3930 VDD.n1217 GND 0.006149f
C3931 VDD.n1218 GND 0.004949f
C3932 VDD.n1219 GND 0.006149f
C3933 VDD.n1220 GND 0.004949f
C3934 VDD.n1221 GND 0.006149f
C3935 VDD.n1222 GND 0.498548f
C3936 VDD.n1223 GND 0.006149f
C3937 VDD.n1224 GND 0.004949f
C3938 VDD.n1225 GND 0.006149f
C3939 VDD.n1226 GND 0.004949f
C3940 VDD.n1227 GND 0.006149f
C3941 VDD.n1228 GND 0.498548f
C3942 VDD.n1229 GND 0.006149f
C3943 VDD.n1230 GND 0.004949f
C3944 VDD.n1231 GND 0.006149f
C3945 VDD.n1232 GND 0.004949f
C3946 VDD.n1233 GND 0.006149f
C3947 VDD.n1234 GND 0.498548f
C3948 VDD.n1235 GND 0.006149f
C3949 VDD.n1236 GND 0.004949f
C3950 VDD.n1237 GND 0.006149f
C3951 VDD.n1238 GND 0.004949f
C3952 VDD.n1239 GND 0.006149f
C3953 VDD.n1240 GND 0.498548f
C3954 VDD.n1241 GND 0.006149f
C3955 VDD.n1242 GND 0.004949f
C3956 VDD.n1243 GND 0.006149f
C3957 VDD.n1244 GND 0.004949f
C3958 VDD.n1245 GND 0.006149f
C3959 VDD.n1246 GND 0.498548f
C3960 VDD.n1247 GND 0.006149f
C3961 VDD.n1248 GND 0.004949f
C3962 VDD.n1249 GND 0.006149f
C3963 VDD.n1250 GND 0.004949f
C3964 VDD.n1251 GND 0.006149f
C3965 VDD.n1252 GND 0.498548f
C3966 VDD.n1253 GND 0.006149f
C3967 VDD.n1254 GND 0.004949f
C3968 VDD.n1255 GND 0.006149f
C3969 VDD.n1256 GND 0.004949f
C3970 VDD.n1257 GND 0.006149f
C3971 VDD.t77 GND 0.498548f
C3972 VDD.n1258 GND 0.006149f
C3973 VDD.n1259 GND 0.004949f
C3974 VDD.n1260 GND 0.006149f
C3975 VDD.n1261 GND 0.004949f
C3976 VDD.n1262 GND 0.006149f
C3977 VDD.n1263 GND 0.498548f
C3978 VDD.n1264 GND 0.006149f
C3979 VDD.n1265 GND 0.004949f
C3980 VDD.n1266 GND 0.006149f
C3981 VDD.n1267 GND 0.004949f
C3982 VDD.n1268 GND 0.006149f
C3983 VDD.n1269 GND 0.498548f
C3984 VDD.n1270 GND 0.006149f
C3985 VDD.n1271 GND 0.004949f
C3986 VDD.n1272 GND 0.006149f
C3987 VDD.n1273 GND 0.004949f
C3988 VDD.n1274 GND 0.006149f
C3989 VDD.n1275 GND 0.498548f
C3990 VDD.n1276 GND 0.006149f
C3991 VDD.n1277 GND 0.004949f
C3992 VDD.n1278 GND 0.006149f
C3993 VDD.n1279 GND 0.004949f
C3994 VDD.n1280 GND 0.006149f
C3995 VDD.n1281 GND 0.498548f
C3996 VDD.n1282 GND 0.006149f
C3997 VDD.n1283 GND 0.004949f
C3998 VDD.n1284 GND 0.006149f
C3999 VDD.n1285 GND 0.004949f
C4000 VDD.n1286 GND 0.006149f
C4001 VDD.n1287 GND 0.498548f
C4002 VDD.n1288 GND 0.006149f
C4003 VDD.n1289 GND 0.004949f
C4004 VDD.n1290 GND 0.006149f
C4005 VDD.n1291 GND 0.004949f
C4006 VDD.n1292 GND 0.006149f
C4007 VDD.t73 GND 0.249274f
C4008 VDD.n1293 GND 0.006149f
C4009 VDD.n1294 GND 0.004949f
C4010 VDD.n1295 GND 0.006149f
C4011 VDD.n1296 GND 0.004949f
C4012 VDD.n1297 GND 0.006149f
C4013 VDD.n1298 GND 0.498548f
C4014 VDD.n1299 GND 0.299129f
C4015 VDD.n1300 GND 0.006149f
C4016 VDD.n1301 GND 0.004949f
C4017 VDD.n1302 GND 0.006149f
C4018 VDD.n1303 GND 0.004949f
C4019 VDD.n1304 GND 0.006149f
C4020 VDD.n1305 GND 0.498548f
C4021 VDD.n1306 GND 0.006149f
C4022 VDD.n1307 GND 0.004949f
C4023 VDD.n1308 GND 0.006149f
C4024 VDD.n1309 GND 0.004949f
C4025 VDD.n1310 GND 0.006149f
C4026 VDD.n1311 GND 0.498548f
C4027 VDD.n1312 GND 0.006149f
C4028 VDD.n1313 GND 0.004949f
C4029 VDD.n1314 GND 0.006149f
C4030 VDD.n1315 GND 0.004949f
C4031 VDD.n1316 GND 0.006149f
C4032 VDD.n1317 GND 0.498548f
C4033 VDD.n1318 GND 0.006149f
C4034 VDD.n1319 GND 0.004949f
C4035 VDD.n1320 GND 0.006149f
C4036 VDD.n1321 GND 0.004949f
C4037 VDD.n1322 GND 0.006149f
C4038 VDD.n1323 GND 0.498548f
C4039 VDD.n1324 GND 0.006149f
C4040 VDD.n1325 GND 0.004949f
C4041 VDD.n1326 GND 0.006149f
C4042 VDD.n1327 GND 0.004949f
C4043 VDD.n1328 GND 0.006149f
C4044 VDD.t110 GND 0.249274f
C4045 VDD.n1329 GND 0.006149f
C4046 VDD.n1330 GND 0.004949f
C4047 VDD.n1331 GND 0.006149f
C4048 VDD.n1332 GND 0.004949f
C4049 VDD.n1333 GND 0.006149f
C4050 VDD.n1334 GND 0.498548f
C4051 VDD.n1335 GND 0.348984f
C4052 VDD.n1336 GND 0.006149f
C4053 VDD.n1337 GND 0.004949f
C4054 VDD.n1338 GND 0.006149f
C4055 VDD.n1339 GND 0.004949f
C4056 VDD.n1340 GND 0.006149f
C4057 VDD.n1341 GND 0.498548f
C4058 VDD.n1342 GND 0.006149f
C4059 VDD.n1343 GND 0.004949f
C4060 VDD.n1344 GND 0.006149f
C4061 VDD.n1345 GND 0.004949f
C4062 VDD.n1346 GND 0.006149f
C4063 VDD.n1347 GND 0.498548f
C4064 VDD.n1348 GND 0.006149f
C4065 VDD.n1349 GND 0.004949f
C4066 VDD.n1350 GND 0.006149f
C4067 VDD.n1351 GND 0.004949f
C4068 VDD.n1352 GND 0.006149f
C4069 VDD.n1353 GND 0.498548f
C4070 VDD.n1354 GND 0.006149f
C4071 VDD.n1355 GND 0.004949f
C4072 VDD.n1356 GND 0.006149f
C4073 VDD.n1357 GND 0.004949f
C4074 VDD.n1358 GND 0.006149f
C4075 VDD.n1359 GND 0.498548f
C4076 VDD.n1360 GND 0.006149f
C4077 VDD.n1361 GND 0.004949f
C4078 VDD.n1362 GND 0.006149f
C4079 VDD.n1363 GND 0.004949f
C4080 VDD.n1364 GND 0.006149f
C4081 VDD.t97 GND 0.249274f
C4082 VDD.n1365 GND 0.006149f
C4083 VDD.n1366 GND 0.004949f
C4084 VDD.n1367 GND 0.006149f
C4085 VDD.n1368 GND 0.004949f
C4086 VDD.n1369 GND 0.006149f
C4087 VDD.n1370 GND 0.498548f
C4088 VDD.n1371 GND 0.398839f
C4089 VDD.n1372 GND 0.006149f
C4090 VDD.n1373 GND 0.004949f
C4091 VDD.n1374 GND 0.006149f
C4092 VDD.n1375 GND 0.004949f
C4093 VDD.n1376 GND 0.006149f
C4094 VDD.n1377 GND 0.498548f
C4095 VDD.n1378 GND 0.006149f
C4096 VDD.n1379 GND 0.004949f
C4097 VDD.n1380 GND 0.006149f
C4098 VDD.n1381 GND 0.004949f
C4099 VDD.n1382 GND 0.006149f
C4100 VDD.n1383 GND 0.498548f
C4101 VDD.n1384 GND 0.006149f
C4102 VDD.n1385 GND 0.004949f
C4103 VDD.n1386 GND 0.006149f
C4104 VDD.n1387 GND 0.004949f
C4105 VDD.n1388 GND 0.006149f
C4106 VDD.n1389 GND 0.498548f
C4107 VDD.n1390 GND 0.006149f
C4108 VDD.n1391 GND 0.004949f
C4109 VDD.n1392 GND 0.006149f
C4110 VDD.n1393 GND 0.004949f
C4111 VDD.n1394 GND 0.006149f
C4112 VDD.n1395 GND 0.498548f
C4113 VDD.n1396 GND 0.006149f
C4114 VDD.n1397 GND 0.004949f
C4115 VDD.n1398 GND 0.006149f
C4116 VDD.n1399 GND 0.004949f
C4117 VDD.n1400 GND 0.006149f
C4118 VDD.t85 GND 0.249274f
C4119 VDD.n1401 GND 0.006149f
C4120 VDD.n1402 GND 0.004949f
C4121 VDD.n1403 GND 0.006149f
C4122 VDD.n1404 GND 0.004949f
C4123 VDD.n1405 GND 0.006149f
C4124 VDD.n1406 GND 0.498548f
C4125 VDD.n1407 GND 0.448694f
C4126 VDD.n1408 GND 0.006149f
C4127 VDD.n1409 GND 0.004949f
C4128 VDD.n1410 GND 0.006149f
C4129 VDD.n1411 GND 0.004949f
C4130 VDD.n1412 GND 0.006149f
C4131 VDD.n1413 GND 0.498548f
C4132 VDD.n1414 GND 0.006149f
C4133 VDD.n1415 GND 0.004949f
C4134 VDD.n1416 GND 0.006149f
C4135 VDD.n1417 GND 0.004949f
C4136 VDD.n1418 GND 0.006149f
C4137 VDD.n1419 GND 0.498548f
C4138 VDD.n1420 GND 0.006149f
C4139 VDD.n1421 GND 0.004949f
C4140 VDD.n1422 GND 0.006149f
C4141 VDD.n1423 GND 0.004949f
C4142 VDD.n1424 GND 0.006149f
C4143 VDD.n1425 GND 0.498548f
C4144 VDD.n1426 GND 0.006149f
C4145 VDD.n1427 GND 0.004949f
C4146 VDD.n1428 GND 0.006149f
C4147 VDD.n1429 GND 0.004949f
C4148 VDD.n1430 GND 0.006149f
C4149 VDD.n1431 GND 0.498548f
C4150 VDD.n1432 GND 0.006149f
C4151 VDD.n1433 GND 0.004949f
C4152 VDD.n1434 GND 0.006149f
C4153 VDD.n1435 GND 0.004949f
C4154 VDD.n1436 GND 0.006149f
C4155 VDD.n1437 GND 0.498548f
C4156 VDD.n1438 GND 0.006149f
C4157 VDD.n1439 GND 0.004949f
C4158 VDD.n1440 GND 0.006149f
C4159 VDD.n1441 GND 0.004949f
C4160 VDD.n1442 GND 0.006149f
C4161 VDD.n1443 GND 0.498548f
C4162 VDD.n1444 GND 0.006149f
C4163 VDD.n1445 GND 0.004949f
C4164 VDD.n1446 GND 0.006149f
C4165 VDD.n1447 GND 0.004949f
C4166 VDD.n1448 GND 0.006149f
C4167 VDD.n1449 GND 0.498548f
C4168 VDD.n1450 GND 0.006149f
C4169 VDD.n1451 GND 0.004949f
C4170 VDD.n1452 GND 0.006149f
C4171 VDD.n1453 GND 0.004949f
C4172 VDD.n1454 GND 0.006149f
C4173 VDD.n1455 GND 0.498548f
C4174 VDD.n1456 GND 0.006149f
C4175 VDD.n1457 GND 0.004949f
C4176 VDD.n1458 GND 0.006149f
C4177 VDD.n1459 GND 0.004949f
C4178 VDD.n1460 GND 0.006149f
C4179 VDD.n1461 GND 0.498548f
C4180 VDD.n1462 GND 0.006149f
C4181 VDD.n1463 GND 0.004949f
C4182 VDD.n1464 GND 0.006149f
C4183 VDD.n1465 GND 0.004949f
C4184 VDD.n1466 GND 0.006149f
C4185 VDD.n1467 GND 0.498548f
C4186 VDD.n1468 GND 0.006149f
C4187 VDD.n1469 GND 0.004949f
C4188 VDD.n1470 GND 0.006149f
C4189 VDD.n1471 GND 0.004949f
C4190 VDD.n1472 GND 0.006149f
C4191 VDD.n1473 GND 0.498548f
C4192 VDD.n1474 GND 0.006149f
C4193 VDD.n1475 GND 0.004949f
C4194 VDD.n1476 GND 0.006149f
C4195 VDD.n1477 GND 0.004949f
C4196 VDD.n1478 GND 0.006149f
C4197 VDD.t14 GND 0.249274f
C4198 VDD.n1479 GND 0.006149f
C4199 VDD.n1480 GND 0.004949f
C4200 VDD.n1481 GND 0.006149f
C4201 VDD.n1482 GND 0.004949f
C4202 VDD.n1483 GND 0.006149f
C4203 VDD.n1484 GND 0.498548f
C4204 VDD.n1485 GND 0.006149f
C4205 VDD.n1486 GND 0.004949f
C4206 VDD.n1487 GND 0.006149f
C4207 VDD.n1488 GND 0.004949f
C4208 VDD.n1489 GND 0.006149f
C4209 VDD.n1490 GND 0.498548f
C4210 VDD.n1491 GND 0.006149f
C4211 VDD.n1492 GND 0.004949f
C4212 VDD.n1493 GND 0.013778f
C4213 VDD.n1494 GND 0.004108f
C4214 VDD.n1495 GND 0.013778f
C4215 VDD.n1496 GND 0.695475f
C4216 VDD.n1497 GND 0.013778f
C4217 VDD.n1498 GND 0.004108f
C4218 VDD.n1499 GND 0.006149f
C4219 VDD.t16 GND 0.179673f
C4220 VDD.t13 GND 0.743196f
C4221 VDD.n1500 GND 0.095879f
C4222 VDD.t15 GND 0.131174f
C4223 VDD.n1501 GND 0.098395f
C4224 VDD.n1502 GND 0.00928f
C4225 VDD.n1503 GND 0.006149f
C4226 VDD.n1526 GND 0.006149f
C4227 VDD.n1527 GND 0.006149f
C4228 VDD.n1528 GND 0.01414f
C4229 VDD.n1529 GND 0.004949f
C4230 VDD.n1530 GND 0.006149f
C4231 VDD.n1531 GND 0.006149f
C4232 VDD.n1532 GND 0.006149f
C4233 VDD.n1533 GND 0.006149f
C4234 VDD.n1534 GND 0.004949f
C4235 VDD.n1535 GND 0.006149f
C4236 VDD.n1536 GND 0.006149f
C4237 VDD.n1537 GND 0.006149f
C4238 VDD.n1538 GND 0.006149f
C4239 VDD.n1539 GND 0.006149f
C4240 VDD.n1540 GND 0.004949f
C4241 VDD.n1541 GND 0.006149f
C4242 VDD.n1542 GND 0.006149f
C4243 VDD.n1543 GND 0.006149f
C4244 VDD.n1544 GND 0.006149f
C4245 VDD.n1545 GND 0.006149f
C4246 VDD.t30 GND 0.179673f
C4247 VDD.t28 GND 0.743196f
C4248 VDD.n1546 GND 0.095879f
C4249 VDD.t29 GND 0.131174f
C4250 VDD.n1547 GND 0.098395f
C4251 VDD.n1548 GND 0.00928f
C4252 VDD.n1549 GND 0.006149f
C4253 VDD.n1550 GND 0.006149f
C4254 VDD.n1551 GND 0.006149f
C4255 VDD.n1552 GND 0.006149f
C4256 VDD.n1553 GND 0.006149f
C4257 VDD.n1554 GND 0.004949f
C4258 VDD.n1555 GND 0.006149f
C4259 VDD.n1556 GND 0.006149f
C4260 VDD.n1557 GND 0.006149f
C4261 VDD.n1558 GND 0.006149f
C4262 VDD.n1559 GND 0.006149f
C4263 VDD.n1560 GND 0.004949f
C4264 VDD.n1561 GND 0.006149f
C4265 VDD.n1562 GND 0.006149f
C4266 VDD.n1563 GND 0.006149f
C4267 VDD.n1564 GND 0.006149f
C4268 VDD.n1565 GND 0.006149f
C4269 VDD.n1566 GND 0.004949f
C4270 VDD.n1567 GND 0.006149f
C4271 VDD.n1568 GND 0.006149f
C4272 VDD.n1569 GND 0.006149f
C4273 VDD.n1570 GND 0.006149f
C4274 VDD.n1571 GND 0.006149f
C4275 VDD.n1572 GND 0.003217f
C4276 VDD.n1573 GND 0.006149f
C4277 VDD.t27 GND 0.179673f
C4278 VDD.t25 GND 0.743196f
C4279 VDD.n1574 GND 0.095879f
C4280 VDD.t26 GND 0.131174f
C4281 VDD.n1575 GND 0.098395f
C4282 VDD.n1576 GND 0.006806f
C4283 VDD.n1577 GND 0.006149f
C4284 VDD.n1578 GND 0.006149f
C4285 VDD.n1579 GND 0.006149f
C4286 VDD.n1580 GND 0.006149f
C4287 VDD.n1581 GND 0.004949f
C4288 VDD.n1582 GND 0.006149f
C4289 VDD.n1583 GND 0.006149f
C4290 VDD.n1584 GND 0.006149f
C4291 VDD.n1585 GND 0.006149f
C4292 VDD.n1586 GND 0.006149f
C4293 VDD.n1587 GND 0.004949f
C4294 VDD.n1588 GND 0.006149f
C4295 VDD.n1589 GND 0.006149f
C4296 VDD.n1590 GND 0.006149f
C4297 VDD.n1591 GND 0.006149f
C4298 VDD.n1592 GND 0.006149f
C4299 VDD.n1593 GND 0.004949f
C4300 VDD.n1594 GND 0.006149f
C4301 VDD.n1595 GND 0.006149f
C4302 VDD.n1596 GND 0.006149f
C4303 VDD.n1597 GND 0.006149f
C4304 VDD.n1598 GND 0.006149f
C4305 VDD.n1599 GND 0.006149f
C4306 VDD.n1600 GND 0.004628f
C4307 VDD.n1601 GND 0.006149f
C4308 VDD.n1602 GND 0.006149f
C4309 VDD.n1603 GND 0.004949f
C4310 VDD.n1604 GND 0.004949f
C4311 VDD.n1605 GND 0.004949f
C4312 VDD.n1606 GND 0.006149f
C4313 VDD.n1607 GND 0.006149f
C4314 VDD.n1608 GND 0.006149f
C4315 VDD.n1609 GND 0.004949f
C4316 VDD.n1610 GND 0.004949f
C4317 VDD.n1611 GND 0.004949f
C4318 VDD.n1612 GND 0.006149f
C4319 VDD.n1613 GND 0.006149f
C4320 VDD.n1614 GND 0.006149f
C4321 VDD.n1615 GND 0.004949f
C4322 VDD.n1616 GND 0.004949f
C4323 VDD.n1617 GND 0.004949f
C4324 VDD.n1618 GND 0.006149f
C4325 VDD.n1619 GND 0.006149f
C4326 VDD.n1620 GND 0.006149f
C4327 VDD.n1621 GND 0.004949f
C4328 VDD.n1622 GND 0.004949f
C4329 VDD.n1623 GND 0.002574f
C4330 VDD.n1624 GND 0.006149f
C4331 VDD.n1625 GND 0.006149f
C4332 VDD.n1626 GND 0.006149f
C4333 VDD.n1627 GND 0.004949f
C4334 VDD.n1628 GND 0.004949f
C4335 VDD.n1629 GND 0.004949f
C4336 VDD.n1630 GND 0.006149f
C4337 VDD.n1631 GND 0.006149f
C4338 VDD.n1632 GND 0.006149f
C4339 VDD.n1633 GND 0.004949f
C4340 VDD.n1634 GND 0.004949f
C4341 VDD.n1635 GND 0.004949f
C4342 VDD.n1636 GND 0.006149f
C4343 VDD.n1637 GND 0.006149f
C4344 VDD.n1638 GND 0.006149f
C4345 VDD.n1639 GND 0.004949f
C4346 VDD.n1640 GND 0.004949f
C4347 VDD.n1641 GND 0.004949f
C4348 VDD.n1642 GND 0.006149f
C4349 VDD.n1643 GND 0.006149f
C4350 VDD.n1644 GND 0.006149f
C4351 VDD.n1645 GND 0.004949f
C4352 VDD.n1646 GND 0.004949f
C4353 VDD.n1647 GND 0.003984f
C4354 VDD.n1648 GND 0.006149f
C4355 VDD.n1649 GND 0.006149f
C4356 VDD.n1650 GND 0.006149f
C4357 VDD.n1651 GND 0.004281f
C4358 VDD.n1652 GND 0.004949f
C4359 VDD.n1653 GND 0.004949f
C4360 VDD.n1654 GND 0.006149f
C4361 VDD.n1655 GND 0.006149f
C4362 VDD.n1656 GND 0.006149f
C4363 VDD.n1657 GND 0.004949f
C4364 VDD.n1658 GND 0.004949f
C4365 VDD.n1659 GND 0.004949f
C4366 VDD.n1660 GND 0.006149f
C4367 VDD.n1661 GND 0.006149f
C4368 VDD.n1662 GND 0.006149f
C4369 VDD.n1663 GND 0.004949f
C4370 VDD.n1664 GND 0.004949f
C4371 VDD.n1665 GND 0.004949f
C4372 VDD.n1666 GND 0.006149f
C4373 VDD.n1667 GND 0.006149f
C4374 VDD.n1668 GND 0.006149f
C4375 VDD.n1669 GND 0.004949f
C4376 VDD.n1670 GND 0.004108f
C4377 VDD.n1671 GND 0.01414f
C4378 VDD.n1673 GND 1.13918f
C4379 VDD.n1675 GND 0.01414f
C4380 VDD.n1676 GND 0.002796f
C4381 VDD.n1677 GND 0.01414f
C4382 VDD.n1678 GND 0.013778f
C4383 VDD.n1679 GND 0.006149f
C4384 VDD.n1680 GND 0.004949f
C4385 VDD.n1681 GND 0.006149f
C4386 VDD.n1682 GND 0.498548f
C4387 VDD.n1683 GND 0.006149f
C4388 VDD.n1684 GND 0.004949f
C4389 VDD.n1685 GND 0.006149f
C4390 VDD.n1686 GND 0.006149f
C4391 VDD.n1687 GND 0.006149f
C4392 VDD.n1688 GND 0.004949f
C4393 VDD.n1689 GND 0.006149f
C4394 VDD.n1690 GND 0.498548f
C4395 VDD.n1691 GND 0.006149f
C4396 VDD.n1692 GND 0.004949f
C4397 VDD.n1693 GND 0.006149f
C4398 VDD.n1694 GND 0.006149f
C4399 VDD.n1695 GND 0.006149f
C4400 VDD.n1696 GND 0.004949f
C4401 VDD.n1697 GND 0.006149f
C4402 VDD.n1698 GND 0.339013f
C4403 VDD.n1699 GND 0.498548f
C4404 VDD.n1700 GND 0.006149f
C4405 VDD.n1701 GND 0.004949f
C4406 VDD.n1702 GND 0.006149f
C4407 VDD.n1703 GND 0.006149f
C4408 VDD.n1704 GND 0.006149f
C4409 VDD.n1705 GND 0.004949f
C4410 VDD.n1706 GND 0.006149f
C4411 VDD.n1707 GND 0.40881f
C4412 VDD.n1708 GND 0.006149f
C4413 VDD.n1709 GND 0.004949f
C4414 VDD.n1710 GND 0.006149f
C4415 VDD.n1711 GND 0.006149f
C4416 VDD.n1712 GND 0.006149f
C4417 VDD.n1713 GND 0.004949f
C4418 VDD.n1714 GND 0.006149f
C4419 VDD.n1715 GND 0.498548f
C4420 VDD.n1716 GND 0.006149f
C4421 VDD.n1717 GND 0.004949f
C4422 VDD.n1718 GND 0.006149f
C4423 VDD.n1719 GND 0.006149f
C4424 VDD.n1720 GND 0.006149f
C4425 VDD.n1721 GND 0.004949f
C4426 VDD.n1722 GND 0.006149f
C4427 VDD.n1723 GND 0.498548f
C4428 VDD.n1724 GND 0.006149f
C4429 VDD.n1725 GND 0.004949f
C4430 VDD.n1726 GND 0.006149f
C4431 VDD.n1727 GND 0.006149f
C4432 VDD.n1728 GND 0.006149f
C4433 VDD.n1729 GND 0.004949f
C4434 VDD.n1730 GND 0.006149f
C4435 VDD.n1731 GND 0.498548f
C4436 VDD.n1732 GND 0.006149f
C4437 VDD.n1733 GND 0.004949f
C4438 VDD.n1734 GND 0.006149f
C4439 VDD.n1735 GND 0.006149f
C4440 VDD.n1736 GND 0.006149f
C4441 VDD.n1737 GND 0.004949f
C4442 VDD.n1738 GND 0.006149f
C4443 VDD.n1739 GND 0.498548f
C4444 VDD.n1740 GND 0.006149f
C4445 VDD.n1741 GND 0.004949f
C4446 VDD.n1742 GND 0.006149f
C4447 VDD.n1743 GND 0.006149f
C4448 VDD.n1744 GND 0.006149f
C4449 VDD.n1745 GND 0.004949f
C4450 VDD.n1746 GND 0.006149f
C4451 VDD.n1747 GND 0.498548f
C4452 VDD.n1748 GND 0.006149f
C4453 VDD.n1749 GND 0.004949f
C4454 VDD.n1750 GND 0.006149f
C4455 VDD.n1751 GND 0.006149f
C4456 VDD.n1752 GND 0.006149f
C4457 VDD.n1753 GND 0.004949f
C4458 VDD.n1754 GND 0.006149f
C4459 VDD.n1755 GND 0.498548f
C4460 VDD.n1756 GND 0.006149f
C4461 VDD.n1757 GND 0.004949f
C4462 VDD.n1758 GND 0.006149f
C4463 VDD.n1759 GND 0.006149f
C4464 VDD.n1760 GND 0.006149f
C4465 VDD.n1761 GND 0.004949f
C4466 VDD.n1762 GND 0.006149f
C4467 VDD.t91 GND 0.498548f
C4468 VDD.n1763 GND 0.006149f
C4469 VDD.n1764 GND 0.004949f
C4470 VDD.n1765 GND 0.006149f
C4471 VDD.n1766 GND 0.006149f
C4472 VDD.n1767 GND 0.006149f
C4473 VDD.n1768 GND 0.004949f
C4474 VDD.n1769 GND 0.006149f
C4475 VDD.n1770 GND 0.498548f
C4476 VDD.n1771 GND 0.006149f
C4477 VDD.n1772 GND 0.004949f
C4478 VDD.n1773 GND 0.006149f
C4479 VDD.n1774 GND 0.006149f
C4480 VDD.n1775 GND 0.006149f
C4481 VDD.n1776 GND 0.004949f
C4482 VDD.n1777 GND 0.006149f
C4483 VDD.n1778 GND 0.498548f
C4484 VDD.n1779 GND 0.006149f
C4485 VDD.n1780 GND 0.004949f
C4486 VDD.n1781 GND 0.006149f
C4487 VDD.n1782 GND 0.006149f
C4488 VDD.n1783 GND 0.006149f
C4489 VDD.n1784 GND 0.004949f
C4490 VDD.n1785 GND 0.006149f
C4491 VDD.n1786 GND 0.498548f
C4492 VDD.n1787 GND 0.006149f
C4493 VDD.n1788 GND 0.004949f
C4494 VDD.n1789 GND 0.006149f
C4495 VDD.n1790 GND 0.006149f
C4496 VDD.n1791 GND 0.006149f
C4497 VDD.n1792 GND 0.004949f
C4498 VDD.n1793 GND 0.006149f
C4499 VDD.n1794 GND 0.498548f
C4500 VDD.n1795 GND 0.006149f
C4501 VDD.n1796 GND 0.004949f
C4502 VDD.n1797 GND 0.006149f
C4503 VDD.n1798 GND 0.006149f
C4504 VDD.n1799 GND 0.006149f
C4505 VDD.n1800 GND 0.004949f
C4506 VDD.n1801 GND 0.006149f
C4507 VDD.n1802 GND 0.498548f
C4508 VDD.n1803 GND 0.006149f
C4509 VDD.n1804 GND 0.004949f
C4510 VDD.n1805 GND 0.006149f
C4511 VDD.n1806 GND 0.006149f
C4512 VDD.n1807 GND 0.006149f
C4513 VDD.n1808 GND 0.004949f
C4514 VDD.n1809 GND 0.006149f
C4515 VDD.n1810 GND 0.299129f
C4516 VDD.n1811 GND 0.006149f
C4517 VDD.n1812 GND 0.004949f
C4518 VDD.n1813 GND 0.006149f
C4519 VDD.n1814 GND 0.006149f
C4520 VDD.n1815 GND 0.006149f
C4521 VDD.n1816 GND 0.004949f
C4522 VDD.n1817 GND 0.006149f
C4523 VDD.n1818 GND 0.498548f
C4524 VDD.n1819 GND 0.006149f
C4525 VDD.n1820 GND 0.004949f
C4526 VDD.n1821 GND 0.006149f
C4527 VDD.n1822 GND 0.006149f
C4528 VDD.n1823 GND 0.006149f
C4529 VDD.n1824 GND 0.004949f
C4530 VDD.n1825 GND 0.006149f
C4531 VDD.n1826 GND 0.498548f
C4532 VDD.n1827 GND 0.006149f
C4533 VDD.n1828 GND 0.004949f
C4534 VDD.n1829 GND 0.006149f
C4535 VDD.n1830 GND 0.006149f
C4536 VDD.n1831 GND 0.006149f
C4537 VDD.n1832 GND 0.004949f
C4538 VDD.n1833 GND 0.006149f
C4539 VDD.n1834 GND 0.498548f
C4540 VDD.n1835 GND 0.006149f
C4541 VDD.n1836 GND 0.004949f
C4542 VDD.n1837 GND 0.006149f
C4543 VDD.n1838 GND 0.006149f
C4544 VDD.n1839 GND 0.006149f
C4545 VDD.n1840 GND 0.004949f
C4546 VDD.n1841 GND 0.006149f
C4547 VDD.n1842 GND 0.498548f
C4548 VDD.n1843 GND 0.006149f
C4549 VDD.n1844 GND 0.004949f
C4550 VDD.n1845 GND 0.006149f
C4551 VDD.n1846 GND 0.006149f
C4552 VDD.n1847 GND 0.006149f
C4553 VDD.n1848 GND 0.004949f
C4554 VDD.n1849 GND 0.006149f
C4555 VDD.n1850 GND 0.498548f
C4556 VDD.n1851 GND 0.006149f
C4557 VDD.n1852 GND 0.004949f
C4558 VDD.n1853 GND 0.006149f
C4559 VDD.n1854 GND 0.006149f
C4560 VDD.n1855 GND 0.006149f
C4561 VDD.n1856 GND 0.004949f
C4562 VDD.n1857 GND 0.006149f
C4563 VDD.n1858 GND 0.348984f
C4564 VDD.n1859 GND 0.006149f
C4565 VDD.n1860 GND 0.004949f
C4566 VDD.n1861 GND 0.006149f
C4567 VDD.n1862 GND 0.006149f
C4568 VDD.n1863 GND 0.006149f
C4569 VDD.n1864 GND 0.004949f
C4570 VDD.n1865 GND 0.006149f
C4571 VDD.n1866 GND 0.498548f
C4572 VDD.n1867 GND 0.006149f
C4573 VDD.n1868 GND 0.004949f
C4574 VDD.n1869 GND 0.006149f
C4575 VDD.n1870 GND 0.006149f
C4576 VDD.n1871 GND 0.006149f
C4577 VDD.n1872 GND 0.004949f
C4578 VDD.n1873 GND 0.006149f
C4579 VDD.n1874 GND 0.498548f
C4580 VDD.n1875 GND 0.006149f
C4581 VDD.n1876 GND 0.004949f
C4582 VDD.n1877 GND 0.006149f
C4583 VDD.n1878 GND 0.004726f
C4584 VDD.t78 GND 0.147596f
C4585 VDD.t111 GND 0.024054f
C4586 VDD.t74 GND 0.024054f
C4587 VDD.n1879 GND 0.106517f
C4588 VDD.n1880 GND 0.66799f
C4589 VDD.t109 GND 0.024054f
C4590 VDD.t107 GND 0.024054f
C4591 VDD.n1881 GND 0.106517f
C4592 VDD.n1882 GND 0.401201f
C4593 VDD.t92 GND 0.142539f
C4594 VDD.n1883 GND 0.321523f
C4595 VDD.t89 GND 0.147596f
C4596 VDD.t117 GND 0.024054f
C4597 VDD.t75 GND 0.024054f
C4598 VDD.n1884 GND 0.106517f
C4599 VDD.n1885 GND 0.66799f
C4600 VDD.t88 GND 0.024054f
C4601 VDD.t106 GND 0.024054f
C4602 VDD.n1886 GND 0.106517f
C4603 VDD.n1887 GND 0.401201f
C4604 VDD.t94 GND 0.142539f
C4605 VDD.n1888 GND 0.298186f
C4606 VDD.n1889 GND 0.307678f
C4607 VDD.t90 GND 0.147596f
C4608 VDD.t116 GND 0.024054f
C4609 VDD.t76 GND 0.024054f
C4610 VDD.n1890 GND 0.106517f
C4611 VDD.n1891 GND 0.66799f
C4612 VDD.t86 GND 0.024054f
C4613 VDD.t98 GND 0.024054f
C4614 VDD.n1892 GND 0.106517f
C4615 VDD.n1893 GND 0.401201f
C4616 VDD.t93 GND 0.142539f
C4617 VDD.n1894 GND 0.298186f
C4618 VDD.n1895 GND 0.378384f
C4619 VDD.n1896 GND 2.95068f
C4620 VDD.n1897 GND 0.330844f
C4621 VDD.n1898 GND 0.004726f
C4622 VDD.n1899 GND 0.004949f
C4623 VDD.n1900 GND 0.006149f
C4624 VDD.n1901 GND 0.498548f
C4625 VDD.n1902 GND 0.006149f
C4626 VDD.n1903 GND 0.004949f
C4627 VDD.n1904 GND 0.006149f
C4628 VDD.n1905 GND 0.006149f
C4629 VDD.n1906 GND 0.006149f
C4630 VDD.n1907 GND 0.004949f
C4631 VDD.n1908 GND 0.006149f
C4632 VDD.n1909 GND 0.498548f
C4633 VDD.n1910 GND 0.006149f
C4634 VDD.n1911 GND 0.004949f
C4635 VDD.n1912 GND 0.006149f
C4636 VDD.n1913 GND 0.006149f
C4637 VDD.n1914 GND 0.006149f
C4638 VDD.n1915 GND 0.004949f
C4639 VDD.n1916 GND 0.006149f
C4640 VDD.n1917 GND 0.498548f
C4641 VDD.n1918 GND 0.006149f
C4642 VDD.n1919 GND 0.004949f
C4643 VDD.n1920 GND 0.006149f
C4644 VDD.n1921 GND 0.006149f
C4645 VDD.n1922 GND 0.006149f
C4646 VDD.n1923 GND 0.004949f
C4647 VDD.n1924 GND 0.006149f
C4648 VDD.n1925 GND 0.398839f
C4649 VDD.n1926 GND 0.006149f
C4650 VDD.n1927 GND 0.004949f
C4651 VDD.n1928 GND 0.006149f
C4652 VDD.n1929 GND 0.006149f
C4653 VDD.n1930 GND 0.006149f
C4654 VDD.n1931 GND 0.004949f
C4655 VDD.n1932 GND 0.006149f
C4656 VDD.n1933 GND 0.498548f
C4657 VDD.n1934 GND 0.006149f
C4658 VDD.n1935 GND 0.004949f
C4659 VDD.n1936 GND 0.006149f
C4660 VDD.n1937 GND 0.006149f
C4661 VDD.n1938 GND 0.006149f
C4662 VDD.n1939 GND 0.004949f
C4663 VDD.n1940 GND 0.006149f
C4664 VDD.n1941 GND 0.498548f
C4665 VDD.n1942 GND 0.006149f
C4666 VDD.n1943 GND 0.004949f
C4667 VDD.n1944 GND 0.006149f
C4668 VDD.n1945 GND 0.006149f
C4669 VDD.n1946 GND 0.006149f
C4670 VDD.n1947 GND 0.004949f
C4671 VDD.n1948 GND 0.006149f
C4672 VDD.n1949 GND 0.498548f
C4673 VDD.n1950 GND 0.006149f
C4674 VDD.n1951 GND 0.004949f
C4675 VDD.n1952 GND 0.006149f
C4676 VDD.n1953 GND 0.006149f
C4677 VDD.n1954 GND 0.006149f
C4678 VDD.n1955 GND 0.004949f
C4679 VDD.n1956 GND 0.006149f
C4680 VDD.n1957 GND 0.498548f
C4681 VDD.n1958 GND 0.006149f
C4682 VDD.n1959 GND 0.004949f
C4683 VDD.n1960 GND 0.006149f
C4684 VDD.n1961 GND 0.006149f
C4685 VDD.n1962 GND 0.006149f
C4686 VDD.n1963 GND 0.004949f
C4687 VDD.n1964 GND 0.006149f
C4688 VDD.n1965 GND 0.498548f
C4689 VDD.n1966 GND 0.006149f
C4690 VDD.n1967 GND 0.004949f
C4691 VDD.n1968 GND 0.006149f
C4692 VDD.n1969 GND 0.006149f
C4693 VDD.n1970 GND 0.006149f
C4694 VDD.n1971 GND 0.004949f
C4695 VDD.n1972 GND 0.006149f
C4696 VDD.n1973 GND 0.448694f
C4697 VDD.n1974 GND 0.006149f
C4698 VDD.n1975 GND 0.004949f
C4699 VDD.n1976 GND 0.006149f
C4700 VDD.n1977 GND 0.006149f
C4701 VDD.n1978 GND 0.006149f
C4702 VDD.n1979 GND 0.004949f
C4703 VDD.n1980 GND 0.006149f
C4704 VDD.n1981 GND 0.498548f
C4705 VDD.n1982 GND 0.006149f
C4706 VDD.n1983 GND 0.004949f
C4707 VDD.n1984 GND 0.006149f
C4708 VDD.n1985 GND 0.006149f
C4709 VDD.n1986 GND 0.006149f
C4710 VDD.n1987 GND 0.004949f
C4711 VDD.n1988 GND 0.006149f
C4712 VDD.n1989 GND 0.498548f
C4713 VDD.n1990 GND 0.006149f
C4714 VDD.n1991 GND 0.004949f
C4715 VDD.n1992 GND 0.006149f
C4716 VDD.n1993 GND 0.006149f
C4717 VDD.n1994 GND 0.006149f
C4718 VDD.n1995 GND 0.004949f
C4719 VDD.n1996 GND 0.006149f
C4720 VDD.n1997 GND 0.498548f
C4721 VDD.n1998 GND 0.006149f
C4722 VDD.n1999 GND 0.004949f
C4723 VDD.n2000 GND 0.006149f
C4724 VDD.n2001 GND 0.006149f
C4725 VDD.n2002 GND 0.006149f
C4726 VDD.n2003 GND 0.004949f
C4727 VDD.n2004 GND 0.006149f
C4728 VDD.n2005 GND 0.498548f
C4729 VDD.n2006 GND 0.006149f
C4730 VDD.n2007 GND 0.004949f
C4731 VDD.n2008 GND 0.006149f
C4732 VDD.n2009 GND 0.006149f
C4733 VDD.n2010 GND 0.006149f
C4734 VDD.n2011 GND 0.004949f
C4735 VDD.n2012 GND 0.006149f
C4736 VDD.n2013 GND 0.498548f
C4737 VDD.n2014 GND 0.006149f
C4738 VDD.n2015 GND 0.004949f
C4739 VDD.n2016 GND 0.006149f
C4740 VDD.n2017 GND 0.006149f
C4741 VDD.n2018 GND 0.006149f
C4742 VDD.n2019 GND 0.004949f
C4743 VDD.n2020 GND 0.006149f
C4744 VDD.n2021 GND 0.498548f
C4745 VDD.n2022 GND 0.006149f
C4746 VDD.n2023 GND 0.004949f
C4747 VDD.n2024 GND 0.006149f
C4748 VDD.n2025 GND 0.006149f
C4749 VDD.n2026 GND 0.006149f
C4750 VDD.n2027 GND 0.004949f
C4751 VDD.n2028 GND 0.006149f
C4752 VDD.n2029 GND 0.498548f
C4753 VDD.n2030 GND 0.006149f
C4754 VDD.n2031 GND 0.004949f
C4755 VDD.n2032 GND 0.006149f
C4756 VDD.n2033 GND 0.006149f
C4757 VDD.n2034 GND 0.006149f
C4758 VDD.n2035 GND 0.004949f
C4759 VDD.n2036 GND 0.006149f
C4760 VDD.n2037 GND 0.498548f
C4761 VDD.n2038 GND 0.006149f
C4762 VDD.n2039 GND 0.004949f
C4763 VDD.n2040 GND 0.006149f
C4764 VDD.n2041 GND 0.006149f
C4765 VDD.n2042 GND 0.006149f
C4766 VDD.n2043 GND 0.004949f
C4767 VDD.n2044 GND 0.006149f
C4768 VDD.n2045 GND 0.498548f
C4769 VDD.n2046 GND 0.006149f
C4770 VDD.n2047 GND 0.004949f
C4771 VDD.n2048 GND 0.006149f
C4772 VDD.n2049 GND 0.006149f
C4773 VDD.n2050 GND 0.006149f
C4774 VDD.n2051 GND 0.004949f
C4775 VDD.n2052 GND 0.006149f
C4776 VDD.n2053 GND 0.498548f
C4777 VDD.n2054 GND 0.006149f
C4778 VDD.n2055 GND 0.004949f
C4779 VDD.n2056 GND 0.006149f
C4780 VDD.n2057 GND 0.006149f
C4781 VDD.n2058 GND 0.006149f
C4782 VDD.n2059 GND 0.004949f
C4783 VDD.n2060 GND 0.006149f
C4784 VDD.n2061 GND 0.498548f
C4785 VDD.n2062 GND 0.006149f
C4786 VDD.n2063 GND 0.004949f
C4787 VDD.n2064 GND 0.006149f
C4788 VDD.n2065 GND 0.006149f
C4789 VDD.n2066 GND 0.006149f
C4790 VDD.n2067 GND 0.004949f
C4791 VDD.n2068 GND 0.006149f
C4792 VDD.n2069 GND 0.40881f
C4793 VDD.n2070 GND 0.498548f
C4794 VDD.n2071 GND 0.006149f
C4795 VDD.n2072 GND 0.004949f
C4796 VDD.n2073 GND 0.006149f
C4797 VDD.n2074 GND 0.006149f
C4798 VDD.n2075 GND 0.006149f
C4799 VDD.n2076 GND 0.004949f
C4800 VDD.n2077 GND 0.006149f
C4801 VDD.n2078 GND 0.339013f
C4802 VDD.n2079 GND 0.006149f
C4803 VDD.n2080 GND 0.004949f
C4804 VDD.n2081 GND 0.006149f
C4805 VDD.n2082 GND 0.006149f
C4806 VDD.n2083 GND 0.006149f
C4807 VDD.n2084 GND 0.006149f
C4808 VDD.n2085 GND 0.006149f
C4809 VDD.n2086 GND 0.004949f
C4810 VDD.n2087 GND 0.006149f
C4811 VDD.n2088 GND 0.498548f
C4812 VDD.n2089 GND 0.006149f
C4813 VDD.n2090 GND 0.004949f
C4814 VDD.n2091 GND 0.006149f
C4815 VDD.n2092 GND 0.006149f
C4816 VDD.n2093 GND 0.006149f
C4817 VDD.n2094 GND 0.004949f
C4818 VDD.n2095 GND 0.006149f
C4819 VDD.n2096 GND 0.498548f
C4820 VDD.n2097 GND 0.006149f
C4821 VDD.n2098 GND 0.006149f
C4822 VDD.n2099 GND 0.004949f
C4823 VDD.n2100 GND 0.004108f
C4824 VDD.n2101 GND 0.012337f
C4825 VDD.n2102 GND 0.951793f
C4826 VDD.n2104 GND 0.004949f
C4827 VDD.n2105 GND 0.006149f
C4828 VDD.n2106 GND 0.006149f
C4829 VDD.n2107 GND 0.004949f
C4830 VDD.n2108 GND 0.004949f
C4831 VDD.n2109 GND 0.006149f
C4832 VDD.n2110 GND 0.006149f
C4833 VDD.n2111 GND 0.004949f
C4834 VDD.n2112 GND 0.004949f
C4835 VDD.n2113 GND 0.006149f
C4836 VDD.n2114 GND 0.006149f
C4837 VDD.n2115 GND 0.004949f
C4838 VDD.n2116 GND 0.004949f
C4839 VDD.n2117 GND 0.006149f
C4840 VDD.n2118 GND 0.006149f
C4841 VDD.n2119 GND 0.004949f
C4842 VDD.n2120 GND 0.004949f
C4843 VDD.n2121 GND 0.006149f
C4844 VDD.n2122 GND 0.006149f
C4845 VDD.n2123 GND 0.004949f
C4846 VDD.n2124 GND 0.004949f
C4847 VDD.n2125 GND 0.006149f
C4848 VDD.n2126 GND 0.006149f
C4849 VDD.n2127 GND 0.004949f
C4850 VDD.n2128 GND 0.004949f
C4851 VDD.n2129 GND 0.006149f
C4852 VDD.n2130 GND 0.006149f
C4853 VDD.n2131 GND 0.004949f
C4854 VDD.n2132 GND 0.002574f
C4855 VDD.n2133 GND 0.006149f
C4856 VDD.n2134 GND 0.006149f
C4857 VDD.n2135 GND 0.003217f
C4858 VDD.n2136 GND 0.004949f
C4859 VDD.n2137 GND 0.006149f
C4860 VDD.n2138 GND 0.006149f
C4861 VDD.n2139 GND 0.004949f
C4862 VDD.n2140 GND 0.004949f
C4863 VDD.n2141 GND 0.006149f
C4864 VDD.n2142 GND 0.006149f
C4865 VDD.n2143 GND 0.004949f
C4866 VDD.n2144 GND 0.004949f
C4867 VDD.n2145 GND 0.006149f
C4868 VDD.n2146 GND 0.006149f
C4869 VDD.n2147 GND 0.004949f
C4870 VDD.n2148 GND 0.004949f
C4871 VDD.n2149 GND 0.006149f
C4872 VDD.n2150 GND 0.006149f
C4873 VDD.n2151 GND 0.004949f
C4874 VDD.n2152 GND 0.004949f
C4875 VDD.n2153 GND 0.006149f
C4876 VDD.n2154 GND 0.006149f
C4877 VDD.n2155 GND 0.004949f
C4878 VDD.n2156 GND 0.004949f
C4879 VDD.n2157 GND 0.006149f
C4880 VDD.n2158 GND 0.006149f
C4881 VDD.n2159 GND 0.004949f
C4882 VDD.n2160 GND 0.004949f
C4883 VDD.n2161 GND 0.006149f
C4884 VDD.n2162 GND 0.006149f
C4885 VDD.n2163 GND 0.004949f
C4886 VDD.n2164 GND 0.006149f
C4887 VDD.n2165 GND 0.006149f
C4888 VDD.n2166 GND 0.006149f
C4889 VDD.n2167 GND 0.00928f
C4890 VDD.n2168 GND 0.004281f
C4891 VDD.n2169 GND 0.006149f
C4892 VDD.n2170 GND 0.006149f
C4893 VDD.n2171 GND 0.004949f
C4894 VDD.n2172 GND 0.004949f
C4895 VDD.n2173 GND 0.006149f
C4896 VDD.n2174 GND 0.006149f
C4897 VDD.n2175 GND 0.004949f
C4898 VDD.n2176 GND 0.004949f
C4899 VDD.n2177 GND 0.006149f
C4900 VDD.n2178 GND 0.006149f
C4901 VDD.n2179 GND 0.004949f
C4902 VDD.n2180 GND 0.004949f
C4903 VDD.n2181 GND 0.006149f
C4904 VDD.n2182 GND 0.006149f
C4905 VDD.n2183 GND 0.004949f
C4906 VDD.n2184 GND 0.004949f
C4907 VDD.n2185 GND 0.006149f
C4908 VDD.n2186 GND 0.006149f
C4909 VDD.n2187 GND 0.004949f
C4910 VDD.n2188 GND 0.004949f
C4911 VDD.n2189 GND 0.006149f
C4912 VDD.n2190 GND 0.004949f
C4913 VDD.n2191 GND 0.004949f
C4914 VDD.n2192 GND 0.006149f
C4915 VDD.n2194 GND 3.71917f
C4916 VDD.n2195 GND 0.695475f
C4917 VDD.n2196 GND 0.013778f
C4918 VDD.n2197 GND 0.004108f
C4919 VDD.n2198 GND 0.012337f
C4920 VDD.n2199 GND 0.951793f
C4921 VDD.n2200 GND 0.053563f
C4922 VDD.n2201 GND 0.004182f
C4923 VDD.n2202 GND 0.004182f
C4924 VDD.n2203 GND 0.004182f
C4925 VDD.n2204 GND 0.004182f
C4926 VDD.n2205 GND 0.004182f
C4927 VDD.n2206 GND 0.004182f
C4928 VDD.n2207 GND 0.004182f
C4929 VDD.n2208 GND 0.004182f
C4930 VDD.n2209 GND 0.004182f
C4931 VDD.n2210 GND 0.004182f
C4932 VDD.n2211 GND 0.004182f
C4933 VDD.n2212 GND 0.004182f
C4934 VDD.n2213 GND 0.004182f
C4935 VDD.n2214 GND 0.004182f
C4936 VDD.n2215 GND 0.004182f
C4937 VDD.n2216 GND 0.003751f
C4938 VDD.n2217 GND 0.004182f
C4939 VDD.n2218 GND 0.004182f
C4940 VDD.n2219 GND 0.002521f
C4941 VDD.n2220 GND 0.004182f
C4942 VDD.n2221 GND 0.004182f
C4943 VDD.n2222 GND 0.004182f
C4944 VDD.n2223 GND 0.004182f
C4945 VDD.n2224 GND 0.009616f
C4946 VDD.n2225 GND 0.009616f
C4947 VDD.n2226 GND 0.009324f
C4948 VDD.n2227 GND 0.004182f
C4949 VDD.n2228 GND 0.004182f
C4950 VDD.n2229 GND 0.004182f
C4951 VDD.n2230 GND 0.004182f
C4952 VDD.n2231 GND 0.004182f
C4953 VDD.n2232 GND 0.004182f
C4954 VDD.n2233 GND 0.004182f
C4955 VDD.n2234 GND 0.004182f
C4956 VDD.n2235 GND 0.004182f
C4957 VDD.n2236 GND 0.004182f
C4958 VDD.n2237 GND 0.004182f
C4959 VDD.n2238 GND 0.004182f
C4960 VDD.n2239 GND 0.004182f
C4961 VDD.n2240 GND 0.004182f
C4962 VDD.n2241 GND 0.004182f
C4963 VDD.n2242 GND 0.004182f
C4964 VDD.n2243 GND 0.004182f
C4965 VDD.n2244 GND 0.004182f
C4966 VDD.n2245 GND 0.004182f
C4967 VDD.n2246 GND 0.004182f
C4968 VDD.n2247 GND 0.004182f
C4969 VDD.n2248 GND 0.004182f
C4970 VDD.n2249 GND 0.004182f
C4971 VDD.n2250 GND 0.004182f
C4972 VDD.n2251 GND 0.004182f
C4973 VDD.n2252 GND 0.004182f
C4974 VDD.n2253 GND 0.004182f
C4975 VDD.n2254 GND 0.004182f
C4976 VDD.n2255 GND 0.004182f
C4977 VDD.n2256 GND 0.004182f
C4978 VDD.n2257 GND 0.004182f
C4979 VDD.n2258 GND 0.004182f
C4980 VDD.n2259 GND 0.004182f
C4981 VDD.n2260 GND 0.004182f
C4982 VDD.n2261 GND 0.004182f
C4983 VDD.n2262 GND 0.004182f
C4984 VDD.n2263 GND 0.004182f
C4985 VDD.n2264 GND 0.004182f
C4986 VDD.n2265 GND 0.004182f
C4987 VDD.n2266 GND 0.004182f
C4988 VDD.n2267 GND 0.004182f
C4989 VDD.n2268 GND 0.004182f
C4990 VDD.n2269 GND 0.004182f
C4991 VDD.n2270 GND 0.004182f
C4992 VDD.n2271 GND 0.004182f
C4993 VDD.n2272 GND 0.004182f
C4994 VDD.n2273 GND 0.004182f
C4995 VDD.n2274 GND 0.004182f
C4996 VDD.n2275 GND 0.004182f
C4997 VDD.n2276 GND 0.004182f
C4998 VDD.n2277 GND 0.004182f
C4999 VDD.n2278 GND 0.004182f
C5000 VDD.n2279 GND 0.004182f
C5001 VDD.n2280 GND 0.004182f
C5002 VDD.n2281 GND 0.004182f
C5003 VDD.n2282 GND 0.004182f
C5004 VDD.n2283 GND 0.004182f
C5005 VDD.n2284 GND 0.004182f
C5006 VDD.n2285 GND 0.004182f
C5007 VDD.n2286 GND 0.004182f
C5008 VDD.n2287 GND 0.004182f
C5009 VDD.n2288 GND 0.004182f
C5010 VDD.n2289 GND 0.004182f
C5011 VDD.n2290 GND 0.004182f
C5012 VDD.n2291 GND 0.004182f
C5013 VDD.n2292 GND 0.004182f
C5014 VDD.n2293 GND 0.004182f
C5015 VDD.n2294 GND 0.004182f
C5016 VDD.n2295 GND 0.004182f
C5017 VDD.n2296 GND 0.004182f
C5018 VDD.n2297 GND 0.004182f
C5019 VDD.n2298 GND 0.004182f
C5020 VDD.n2299 GND 0.004182f
C5021 VDD.n2300 GND 0.004182f
C5022 VDD.n2301 GND 0.004182f
C5023 VDD.n2302 GND 0.004182f
C5024 VDD.n2303 GND 0.004182f
C5025 VDD.n2304 GND 0.004182f
C5026 VDD.n2305 GND 0.004182f
C5027 VDD.n2306 GND 0.004182f
C5028 VDD.n2307 GND 0.004182f
C5029 VDD.n2308 GND 0.004182f
C5030 VDD.n2309 GND 0.004182f
C5031 VDD.n2310 GND 0.004182f
C5032 VDD.n2311 GND 0.004182f
C5033 VDD.n2312 GND 0.004182f
C5034 VDD.n2313 GND 0.004182f
C5035 VDD.n2314 GND 0.004182f
C5036 VDD.n2315 GND 0.004182f
C5037 VDD.n2316 GND 0.004182f
C5038 VDD.n2317 GND 0.004182f
C5039 VDD.n2318 GND 0.004182f
C5040 VDD.n2319 GND 0.004182f
C5041 VDD.n2320 GND 0.004182f
C5042 VDD.n2321 GND 0.004182f
C5043 VDD.n2322 GND 0.004182f
C5044 VDD.n2323 GND 0.004182f
C5045 VDD.n2324 GND 0.004182f
C5046 VDD.n2325 GND 0.004182f
C5047 VDD.n2326 GND 0.004182f
C5048 VDD.n2327 GND 0.004182f
C5049 VDD.n2328 GND 0.004182f
C5050 VDD.n2329 GND 0.004182f
C5051 VDD.n2330 GND 0.004182f
C5052 VDD.n2331 GND 0.004182f
C5053 VDD.n2332 GND 0.004182f
C5054 VDD.n2333 GND 0.004182f
C5055 VDD.n2334 GND 0.004182f
C5056 VDD.n2335 GND 0.004182f
C5057 VDD.n2336 GND 0.004182f
C5058 VDD.n2337 GND 0.004182f
C5059 VDD.n2338 GND 0.004182f
C5060 VDD.n2339 GND 0.004182f
C5061 VDD.n2340 GND 0.004182f
C5062 VDD.n2341 GND 0.004182f
C5063 VDD.n2342 GND 0.004182f
C5064 VDD.n2343 GND 0.004182f
C5065 VDD.n2344 GND 0.004182f
C5066 VDD.n2345 GND 0.004182f
C5067 VDD.n2346 GND 0.004182f
C5068 VDD.n2347 GND 0.004182f
C5069 VDD.n2348 GND 0.004182f
C5070 VDD.n2349 GND 0.004182f
C5071 VDD.n2350 GND 0.004182f
C5072 VDD.n2351 GND 0.004182f
C5073 VDD.n2352 GND 0.004182f
C5074 VDD.n2353 GND 0.004182f
C5075 VDD.n2354 GND 0.004182f
C5076 VDD.n2355 GND 0.004182f
C5077 VDD.n2356 GND 0.004182f
C5078 VDD.n2357 GND 0.08226f
C5079 VDD.n2358 GND 0.004182f
C5080 VDD.n2359 GND 0.004182f
C5081 VDD.n2360 GND 0.004182f
C5082 VDD.n2361 GND 0.004182f
C5083 VDD.n2362 GND 0.004182f
C5084 VDD.n2363 GND 0.004182f
C5085 VDD.n2364 GND 0.004182f
C5086 VDD.n2365 GND 0.004182f
C5087 VDD.n2366 GND 0.004182f
C5088 VDD.n2367 GND 0.004182f
C5089 VDD.n2368 GND 0.004182f
C5090 VDD.n2369 GND 0.004182f
C5091 VDD.n2370 GND 0.004182f
C5092 VDD.n2371 GND 0.004182f
C5093 VDD.n2372 GND 0.004182f
C5094 VDD.n2373 GND 0.004182f
C5095 VDD.n2374 GND 0.004182f
C5096 VDD.n2375 GND 0.004182f
C5097 VDD.n2376 GND 0.004182f
C5098 VDD.n2377 GND 0.004182f
C5099 VDD.n2378 GND 0.004182f
C5100 VDD.n2379 GND 0.004182f
C5101 VDD.n2380 GND 0.004182f
C5102 VDD.n2381 GND 0.004182f
C5103 VDD.n2382 GND 0.004182f
C5104 VDD.n2383 GND 0.004182f
C5105 VDD.n2384 GND 0.004182f
C5106 VDD.n2385 GND 0.004182f
C5107 VDD.n2386 GND 0.004182f
C5108 VDD.n2387 GND 0.004182f
C5109 VDD.n2388 GND 0.004182f
C5110 VDD.n2389 GND 0.004182f
C5111 VDD.n2390 GND 0.004182f
C5112 VDD.n2391 GND 0.004182f
C5113 VDD.n2392 GND 0.004182f
C5114 VDD.n2393 GND 0.004182f
C5115 VDD.n2394 GND 0.004182f
C5116 VDD.n2395 GND 0.004182f
C5117 VDD.n2396 GND 0.009324f
C5118 VDD.n2397 GND 0.009616f
C5119 VDD.n2398 GND 0.009616f
C5120 VDD.n2399 GND 2.17866f
C5121 VDD.n2401 GND 0.004182f
C5122 VDD.n2402 GND 0.004182f
C5123 VDD.n2403 GND 0.009616f
C5124 VDD.n2404 GND 0.009324f
C5125 VDD.n2405 GND 0.009324f
C5126 VDD.n2406 GND 0.334027f
C5127 VDD.n2407 GND 0.009324f
C5128 VDD.n2408 GND 0.009324f
C5129 VDD.n2409 GND 0.004182f
C5130 VDD.n2410 GND 0.004182f
C5131 VDD.n2411 GND 0.004182f
C5132 VDD.n2412 GND 0.339013f
C5133 VDD.n2413 GND 0.004182f
C5134 VDD.n2414 GND 0.004182f
C5135 VDD.n2415 GND 0.004182f
C5136 VDD.n2416 GND 0.004182f
C5137 VDD.n2417 GND 0.004182f
C5138 VDD.n2418 GND 0.339013f
C5139 VDD.n2419 GND 0.004182f
C5140 VDD.n2420 GND 0.004182f
C5141 VDD.n2421 GND 0.004182f
C5142 VDD.n2422 GND 0.004182f
C5143 VDD.n2423 GND 0.004182f
C5144 VDD.n2424 GND 0.339013f
C5145 VDD.n2425 GND 0.004182f
C5146 VDD.n2426 GND 0.004182f
C5147 VDD.n2427 GND 0.004182f
C5148 VDD.n2428 GND 0.004182f
C5149 VDD.n2429 GND 0.004182f
C5150 VDD.n2430 GND 0.201912f
C5151 VDD.n2431 GND 0.004182f
C5152 VDD.n2432 GND 0.004182f
C5153 VDD.n2433 GND 0.004182f
C5154 VDD.n2434 GND 0.004182f
C5155 VDD.n2435 GND 0.004182f
C5156 VDD.n2436 GND 0.339013f
C5157 VDD.n2437 GND 0.004182f
C5158 VDD.n2438 GND 0.004182f
C5159 VDD.n2439 GND 0.004182f
C5160 VDD.n2440 GND 0.004182f
C5161 VDD.n2441 GND 0.004182f
C5162 VDD.n2442 GND 0.189448f
C5163 VDD.n2443 GND 0.004182f
C5164 VDD.n2444 GND 0.004182f
C5165 VDD.n2445 GND 0.004182f
C5166 VDD.n2446 GND 0.004182f
C5167 VDD.n2447 GND 0.004182f
C5168 VDD.n2448 GND 0.339013f
C5169 VDD.n2449 GND 0.004182f
C5170 VDD.n2450 GND 0.004182f
C5171 VDD.n2451 GND 0.004182f
C5172 VDD.n2452 GND 0.004182f
C5173 VDD.n2453 GND 0.004182f
C5174 VDD.n2454 GND 0.339013f
C5175 VDD.n2455 GND 0.004182f
C5176 VDD.n2456 GND 0.004182f
C5177 VDD.n2457 GND 0.004182f
C5178 VDD.n2458 GND 0.004182f
C5179 VDD.n2459 GND 0.004182f
C5180 VDD.n2460 GND 0.339013f
C5181 VDD.n2461 GND 0.004182f
C5182 VDD.n2462 GND 0.004182f
C5183 VDD.n2463 GND 0.004182f
C5184 VDD.n2464 GND 0.004182f
C5185 VDD.n2465 GND 0.004182f
C5186 VDD.n2466 GND 0.339013f
C5187 VDD.n2467 GND 0.004182f
C5188 VDD.n2468 GND 0.004182f
C5189 VDD.n2469 GND 0.004182f
C5190 VDD.n2470 GND 0.004182f
C5191 VDD.n2471 GND 0.004182f
C5192 VDD.n2472 GND 0.339013f
C5193 VDD.n2473 GND 0.004182f
C5194 VDD.n2474 GND 0.004182f
C5195 VDD.n2475 GND 0.004182f
C5196 VDD.n2476 GND 0.004182f
C5197 VDD.n2477 GND 0.004182f
C5198 VDD.n2478 GND 0.294144f
C5199 VDD.n2479 GND 0.004182f
C5200 VDD.n2480 GND 0.004182f
C5201 VDD.n2481 GND 0.004182f
C5202 VDD.n2482 GND 0.004182f
C5203 VDD.n2483 GND 0.004182f
C5204 VDD.n2484 GND 0.301622f
C5205 VDD.n2485 GND 0.004182f
C5206 VDD.n2486 GND 0.004182f
C5207 VDD.n2487 GND 0.004182f
C5208 VDD.n2488 GND 0.004182f
C5209 VDD.n2489 GND 0.004182f
C5210 VDD.n2490 GND 0.339013f
C5211 VDD.n2491 GND 0.004182f
C5212 VDD.n2492 GND 0.004182f
C5213 VDD.n2493 GND 0.004182f
C5214 VDD.n2494 GND 0.004182f
C5215 VDD.n2495 GND 0.004182f
C5216 VDD.n2496 GND 0.339013f
C5217 VDD.n2497 GND 0.004182f
C5218 VDD.n2498 GND 0.004182f
C5219 VDD.n2499 GND 0.004182f
C5220 VDD.n2500 GND 0.004182f
C5221 VDD.n2501 GND 0.004182f
C5222 VDD.n2502 GND 0.339013f
C5223 VDD.n2503 GND 0.004182f
C5224 VDD.n2504 GND 0.004182f
C5225 VDD.n2505 GND 0.004182f
C5226 VDD.n2506 GND 0.004182f
C5227 VDD.n2507 GND 0.004182f
C5228 VDD.n2508 GND 0.339013f
C5229 VDD.n2509 GND 0.004182f
C5230 VDD.n2510 GND 0.004182f
C5231 VDD.n2511 GND 0.004182f
C5232 VDD.n2512 GND 0.004182f
C5233 VDD.n2513 GND 0.004182f
C5234 VDD.n2514 GND 0.339013f
C5235 VDD.n2515 GND 0.004182f
C5236 VDD.n2516 GND 0.004182f
C5237 VDD.n2517 GND 0.004182f
C5238 VDD.n2518 GND 0.004182f
C5239 VDD.n2519 GND 0.004182f
C5240 VDD.n2520 GND 0.18197f
C5241 VDD.n2521 GND 0.004182f
C5242 VDD.n2522 GND 0.004182f
C5243 VDD.n2523 GND 0.004182f
C5244 VDD.n2524 GND 0.004182f
C5245 VDD.n2525 GND 0.004182f
C5246 VDD.n2526 GND 0.339013f
C5247 VDD.n2527 GND 0.004182f
C5248 VDD.n2528 GND 0.004182f
C5249 VDD.n2529 GND 0.004182f
C5250 VDD.n2530 GND 0.004182f
C5251 VDD.n2531 GND 0.004182f
C5252 VDD.n2532 GND 0.339013f
C5253 VDD.n2533 GND 0.004182f
C5254 VDD.n2534 GND 0.004182f
C5255 VDD.n2535 GND 0.004182f
C5256 VDD.n2536 GND 0.004182f
C5257 VDD.n2537 GND 0.004182f
C5258 VDD.n2538 GND 0.221854f
C5259 VDD.n2539 GND 0.004182f
C5260 VDD.n2540 GND 0.004182f
C5261 VDD.n2541 GND 0.004182f
C5262 VDD.n2542 GND 0.004182f
C5263 VDD.n2543 GND 0.004182f
C5264 VDD.n2544 GND 0.339013f
C5265 VDD.n2545 GND 0.004182f
C5266 VDD.n2546 GND 0.004182f
C5267 VDD.n2547 GND 0.004182f
C5268 VDD.n2548 GND 0.004182f
C5269 VDD.n2549 GND 0.004182f
C5270 VDD.n2550 GND 0.339013f
C5271 VDD.n2551 GND 0.004182f
C5272 VDD.n2552 GND 0.004182f
C5273 VDD.n2553 GND 0.004182f
C5274 VDD.n2554 GND 0.004182f
C5275 VDD.n2555 GND 0.004182f
C5276 VDD.n2556 GND 0.326549f
C5277 VDD.n2557 GND 0.004182f
C5278 VDD.n2558 GND 0.004182f
C5279 VDD.n2559 GND 0.004182f
C5280 VDD.n2560 GND 0.004182f
C5281 VDD.n2561 GND 0.004182f
C5282 VDD.n2562 GND 0.339013f
C5283 VDD.n2563 GND 0.004182f
C5284 VDD.n2564 GND 0.004182f
C5285 VDD.n2565 GND 0.004182f
C5286 VDD.n2566 GND 0.004182f
C5287 VDD.n2567 GND 0.004182f
C5288 VDD.n2568 GND 0.339013f
C5289 VDD.n2569 GND 0.004182f
C5290 VDD.n2570 GND 0.004182f
C5291 VDD.n2571 GND 0.004182f
C5292 VDD.n2572 GND 0.004182f
C5293 VDD.n2573 GND 0.004182f
C5294 VDD.n2574 GND 0.261738f
C5295 VDD.n2575 GND 0.004182f
C5296 VDD.n2576 GND 0.004182f
C5297 VDD.n2577 GND 0.004182f
C5298 VDD.n2578 GND 0.004182f
C5299 VDD.n2579 GND 0.004182f
C5300 VDD.n2580 GND 0.339013f
C5301 VDD.n2581 GND 0.004182f
C5302 VDD.n2582 GND 0.004182f
C5303 VDD.n2583 GND 0.004182f
C5304 VDD.n2584 GND 0.004182f
C5305 VDD.n2585 GND 0.004182f
C5306 VDD.n2586 GND 0.339013f
C5307 VDD.n2587 GND 0.004182f
C5308 VDD.n2588 GND 0.004182f
C5309 VDD.n2589 GND 0.004182f
C5310 VDD.n2590 GND 0.004182f
C5311 VDD.n2591 GND 0.004182f
C5312 VDD.n2592 GND 0.339013f
C5313 VDD.n2593 GND 0.004182f
C5314 VDD.n2594 GND 0.004182f
C5315 VDD.n2595 GND 0.004182f
C5316 VDD.n2596 GND 0.004182f
C5317 VDD.n2597 GND 0.004182f
C5318 VDD.n2598 GND 0.206898f
C5319 VDD.n2599 GND 0.004182f
C5320 VDD.n2600 GND 0.004182f
C5321 VDD.n2601 GND 0.004182f
C5322 VDD.n2602 GND 0.004182f
C5323 VDD.n2603 GND 0.004182f
C5324 VDD.n2604 GND 0.339013f
C5325 VDD.n2605 GND 0.004182f
C5326 VDD.n2606 GND 0.004182f
C5327 VDD.n2607 GND 0.004182f
C5328 VDD.n2608 GND 0.004182f
C5329 VDD.n2609 GND 0.004182f
C5330 VDD.n2610 GND 0.339013f
C5331 VDD.n2611 GND 0.004182f
C5332 VDD.n2612 GND 0.004182f
C5333 VDD.n2613 GND 0.004182f
C5334 VDD.n2614 GND 0.004182f
C5335 VDD.n2615 GND 0.004182f
C5336 VDD.n2616 GND 0.271709f
C5337 VDD.n2617 GND 0.004182f
C5338 VDD.n2618 GND 0.004182f
C5339 VDD.n2619 GND 0.004182f
C5340 VDD.n2620 GND 0.004182f
C5341 VDD.n2621 GND 0.004182f
C5342 VDD.n2622 GND 0.339013f
C5343 VDD.n2623 GND 0.004182f
C5344 VDD.n2624 GND 0.004182f
C5345 VDD.n2625 GND 0.004182f
C5346 VDD.n2626 GND 0.004182f
C5347 VDD.n2627 GND 0.004182f
C5348 VDD.n2628 GND 0.339013f
C5349 VDD.n2629 GND 0.004182f
C5350 VDD.n2630 GND 0.004182f
C5351 VDD.n2631 GND 0.004182f
C5352 VDD.n2632 GND 0.004182f
C5353 VDD.n2633 GND 0.004182f
C5354 VDD.n2634 GND 0.339013f
C5355 VDD.n2635 GND 0.004182f
C5356 VDD.n2636 GND 0.004182f
C5357 VDD.n2637 GND 0.004182f
C5358 VDD.n2638 GND 0.004182f
C5359 VDD.n2639 GND 0.004182f
C5360 VDD.n2640 GND 0.339013f
C5361 VDD.n2641 GND 0.004182f
C5362 VDD.n2642 GND 0.004182f
C5363 VDD.n2643 GND 0.004182f
C5364 VDD.n2644 GND 0.004182f
C5365 VDD.n2645 GND 0.004182f
C5366 VDD.n2646 GND 0.306607f
C5367 VDD.n2647 GND 0.004182f
C5368 VDD.n2648 GND 0.004182f
C5369 VDD.n2649 GND 0.004182f
C5370 VDD.n2650 GND 0.004182f
C5371 VDD.n2651 GND 0.004182f
C5372 VDD.n2652 GND 0.004182f
C5373 VDD.n2653 GND 0.004182f
C5374 VDD.n2654 GND 0.211883f
C5375 VDD.n2655 GND 0.004182f
C5376 VDD.n2656 GND 0.004182f
C5377 VDD.n2657 GND 0.004182f
C5378 VDD.n2658 GND 0.004182f
C5379 VDD.n2659 GND 0.004182f
C5380 VDD.n2660 GND 0.339013f
C5381 VDD.n2661 GND 0.004182f
C5382 VDD.n2662 GND 0.004182f
C5383 VDD.n2663 GND 0.004182f
C5384 VDD.n2664 GND 0.004182f
C5385 VDD.n2665 GND 0.004182f
C5386 VDD.n2666 GND 0.004182f
C5387 VDD.n2667 GND 0.004182f
C5388 VDD.n2668 GND 0.009324f
C5389 VDD.n2669 GND 0.009844f
C5390 VDD.n2670 GND 0.009096f
C5391 VDD.n2671 GND 0.004182f
C5392 VDD.n2672 GND 0.004182f
C5393 VDD.n2673 GND 0.004182f
C5394 VDD.n2674 GND 0.004182f
C5395 VDD.n2675 GND 0.004182f
C5396 VDD.n2676 GND 0.002521f
C5397 VDD.n2677 GND 0.005159f
C5398 VDD.n2678 GND 0.003751f
C5399 VDD.n2679 GND 0.004182f
C5400 VDD.n2680 GND 0.004182f
C5401 VDD.n2681 GND 0.004182f
C5402 VDD.n2682 GND 0.004182f
C5403 VDD.n2683 GND 0.004182f
C5404 VDD.n2684 GND 0.004182f
C5405 VDD.n2685 GND 0.004182f
C5406 VDD.n2686 GND 0.004182f
C5407 VDD.n2687 GND 0.004182f
C5408 VDD.n2688 GND 0.004182f
C5409 VDD.n2689 GND 0.004182f
C5410 VDD.n2690 GND 0.004182f
C5411 VDD.n2691 GND 0.004182f
C5412 VDD.n2692 GND 0.004182f
C5413 VDD.n2693 GND 0.004182f
C5414 VDD.n2694 GND 0.004182f
C5415 VDD.n2695 GND 0.004182f
C5416 VDD.n2696 GND 0.004182f
C5417 VDD.n2697 GND 0.004182f
C5418 VDD.n2698 GND 0.004182f
C5419 VDD.n2699 GND 0.004182f
C5420 VDD.n2700 GND 0.004182f
C5421 VDD.n2701 GND 0.004182f
C5422 VDD.n2702 GND 0.004182f
C5423 VDD.n2703 GND 0.004182f
C5424 VDD.n2704 GND 0.004182f
C5425 VDD.n2705 GND 0.004182f
C5426 VDD.n2706 GND 0.004182f
C5427 VDD.n2707 GND 0.004182f
C5428 VDD.n2708 GND 0.004182f
C5429 VDD.n2709 GND 0.004182f
C5430 VDD.n2710 GND 0.004182f
C5431 VDD.n2711 GND 0.004182f
C5432 VDD.n2712 GND 0.004182f
C5433 VDD.n2713 GND 0.004182f
C5434 VDD.n2714 GND 0.004182f
C5435 VDD.n2715 GND 0.004182f
C5436 VDD.n2716 GND 0.004182f
C5437 VDD.n2717 GND 0.004182f
C5438 VDD.n2718 GND 0.009616f
C5439 VDD.n2719 GND 0.009616f
C5440 VDD.n2720 GND 0.009324f
C5441 VDD.n2721 GND 0.009324f
C5442 VDD.n2722 GND 0.004182f
C5443 VDD.n2723 GND 0.004182f
C5444 VDD.n2724 GND 0.004182f
C5445 VDD.n2725 GND 0.004182f
C5446 VDD.n2726 GND 0.339013f
C5447 VDD.n2727 GND 0.004182f
C5448 VDD.n2728 GND 0.004182f
C5449 VDD.n2729 GND 0.004182f
C5450 VDD.n2730 GND 0.004182f
C5451 VDD.n2731 GND 0.004182f
C5452 VDD.n2732 GND 0.339013f
C5453 VDD.n2733 GND 0.004182f
C5454 VDD.n2734 GND 0.009324f
C5455 VDD.n2735 GND 0.009616f
C5456 VDD.n2736 GND 0.009096f
C5457 VDD.n2737 GND 0.004182f
C5458 VDD.n2738 GND 0.004182f
C5459 VDD.n2739 GND 0.004182f
C5460 VDD.n2740 GND 0.004182f
C5461 VDD.n2741 GND 0.002521f
C5462 VDD.n2742 GND 0.004182f
C5463 VDD.n2743 GND 0.004182f
C5464 VDD.n2744 GND 0.003751f
C5465 VDD.n2745 GND 0.004182f
C5466 VDD.n2746 GND 0.004182f
C5467 VDD.n2747 GND 0.004182f
C5468 VDD.n2748 GND 0.004182f
C5469 VDD.n2749 GND 0.004182f
C5470 VDD.n2750 GND 0.004182f
C5471 VDD.n2751 GND 0.004182f
C5472 VDD.n2752 GND 0.004182f
C5473 VDD.n2753 GND 0.004182f
C5474 VDD.n2754 GND 0.004182f
C5475 VDD.n2755 GND 0.004182f
C5476 VDD.n2756 GND 0.004182f
C5477 VDD.n2757 GND 0.004182f
C5478 VDD.n2758 GND 0.004182f
C5479 VDD.n2759 GND 0.004182f
C5480 VDD.n2760 GND 0.004182f
C5481 VDD.n2761 GND 0.004182f
C5482 VDD.n2762 GND 0.004182f
C5483 VDD.n2763 GND 0.004182f
C5484 VDD.n2764 GND 0.004182f
C5485 VDD.n2765 GND 0.004182f
C5486 VDD.n2766 GND 0.004182f
C5487 VDD.n2767 GND 0.004182f
C5488 VDD.n2768 GND 0.004182f
C5489 VDD.n2769 GND 0.004182f
C5490 VDD.n2770 GND 0.004182f
C5491 VDD.n2771 GND 0.004182f
C5492 VDD.n2772 GND 0.004182f
C5493 VDD.n2773 GND 0.004182f
C5494 VDD.n2774 GND 0.004182f
C5495 VDD.n2775 GND 0.004182f
C5496 VDD.n2776 GND 0.004182f
C5497 VDD.n2777 GND 0.004182f
C5498 VDD.n2778 GND 0.004182f
C5499 VDD.n2779 GND 0.004182f
C5500 VDD.n2780 GND 0.004182f
C5501 VDD.n2781 GND 0.004182f
C5502 VDD.n2782 GND 0.009616f
C5503 VDD.n2783 GND 0.009616f
C5504 VDD.n2784 GND 2.08643f
C5505 VDD.n2807 GND 0.009616f
C5506 VDD.n2808 GND 0.004182f
C5507 VDD.n2809 GND 0.004182f
C5508 VDD.t53 GND 0.18185f
C5509 VDD.t51 GND 0.551129f
C5510 VDD.n2810 GND 0.095638f
C5511 VDD.t52 GND 0.141776f
C5512 VDD.n2811 GND 0.095144f
C5513 VDD.n2812 GND 0.005159f
C5514 VDD.n2813 GND 0.004182f
C5515 VDD.n2814 GND 0.004182f
C5516 VDD.n2815 GND 0.004182f
C5517 VDD.n2816 GND 0.004182f
C5518 VDD.n2817 GND 0.004182f
C5519 VDD.n2818 GND 0.004182f
C5520 VDD.n2819 GND 0.004182f
C5521 VDD.n2820 GND 0.004182f
C5522 VDD.n2821 GND 0.004182f
C5523 VDD.n2822 GND 0.004182f
C5524 VDD.n2823 GND 0.004182f
C5525 VDD.n2824 GND 0.004182f
C5526 VDD.n2825 GND 0.004182f
C5527 VDD.n2826 GND 0.004182f
C5528 VDD.n2827 GND 0.004182f
C5529 VDD.n2828 GND 0.004182f
C5530 VDD.n2829 GND 0.004182f
C5531 VDD.n2830 GND 0.004182f
C5532 VDD.n2831 GND 0.004182f
C5533 VDD.n2832 GND 0.004182f
C5534 VDD.n2833 GND 0.004182f
C5535 VDD.n2834 GND 0.004182f
C5536 VDD.n2835 GND 0.004182f
C5537 VDD.n2836 GND 0.004182f
C5538 VDD.n2837 GND 0.004182f
C5539 VDD.n2838 GND 0.004182f
C5540 VDD.n2839 GND 0.004182f
C5541 VDD.n2840 GND 0.004182f
C5542 VDD.n2841 GND 0.004182f
C5543 VDD.n2842 GND 0.004182f
C5544 VDD.n2843 GND 0.004182f
C5545 VDD.n2844 GND 0.004182f
C5546 VDD.t50 GND 0.18185f
C5547 VDD.t47 GND 0.551129f
C5548 VDD.n2845 GND 0.095638f
C5549 VDD.t49 GND 0.141776f
C5550 VDD.n2846 GND 0.095144f
C5551 VDD.n2847 GND 0.004182f
C5552 VDD.n2848 GND 0.004182f
C5553 VDD.n2849 GND 0.004182f
C5554 VDD.n2850 GND 0.004182f
C5555 VDD.n2851 GND 0.004182f
C5556 VDD.n2852 GND 0.004182f
C5557 VDD.n2853 GND 0.004182f
C5558 VDD.n2854 GND 0.004182f
C5559 VDD.n2855 GND 0.004182f
C5560 VDD.n2856 GND 0.004182f
C5561 VDD.n2857 GND 0.004182f
C5562 VDD.n2858 GND 0.004182f
C5563 VDD.n2859 GND 0.004182f
C5564 VDD.n2860 GND 0.004182f
C5565 VDD.n2861 GND 0.004182f
C5566 VDD.n2862 GND 0.004182f
C5567 VDD.n2863 GND 0.004182f
C5568 VDD.n2864 GND 0.004182f
C5569 VDD.n2865 GND 0.004182f
C5570 VDD.n2866 GND 0.004182f
C5571 VDD.n2867 GND 0.004182f
C5572 VDD.n2868 GND 0.004182f
C5573 VDD.n2869 GND 0.004182f
C5574 VDD.n2870 GND 0.004182f
C5575 VDD.n2871 GND 0.004182f
C5576 VDD.n2872 GND 0.004182f
C5577 VDD.n2873 GND 0.004182f
C5578 VDD.n2874 GND 0.004182f
C5579 VDD.n2875 GND 0.004182f
C5580 VDD.n2876 GND 0.004182f
C5581 VDD.n2877 GND 0.004182f
C5582 VDD.n2878 GND 0.004182f
C5583 VDD.n2879 GND 0.004182f
C5584 VDD.n2880 GND 0.004182f
C5585 VDD.n2881 GND 0.004182f
C5586 VDD.n2882 GND 0.004182f
C5587 VDD.n2883 GND 0.004182f
C5588 VDD.n2884 GND 0.003751f
C5589 VDD.n2885 GND 0.005159f
C5590 VDD.n2886 GND 0.002521f
C5591 VDD.n2887 GND 0.004182f
C5592 VDD.n2888 GND 0.004182f
C5593 VDD.n2889 GND 0.004182f
C5594 VDD.n2890 GND 0.004182f
C5595 VDD.n2891 GND 0.004182f
C5596 VDD.n2892 GND 0.009616f
C5597 VDD.n2893 GND 0.009324f
C5598 VDD.n2894 GND 0.009324f
C5599 VDD.n2895 GND 0.004182f
C5600 VDD.n2896 GND 0.004182f
C5601 VDD.n2897 GND 0.004182f
C5602 VDD.n2898 GND 0.004182f
C5603 VDD.n2899 GND 0.004182f
C5604 VDD.n2900 GND 0.004182f
C5605 VDD.n2901 GND 0.004182f
C5606 VDD.n2902 GND 0.004182f
C5607 VDD.n2903 GND 0.004182f
C5608 VDD.n2904 GND 0.004182f
C5609 VDD.n2905 GND 0.004182f
C5610 VDD.n2906 GND 0.004182f
C5611 VDD.n2907 GND 0.004182f
C5612 VDD.n2908 GND 0.004182f
C5613 VDD.n2909 GND 0.004182f
C5614 VDD.n2910 GND 0.004182f
C5615 VDD.n2911 GND 0.004182f
C5616 VDD.n2912 GND 0.004182f
C5617 VDD.n2913 GND 0.004182f
C5618 VDD.n2914 GND 0.004182f
C5619 VDD.n2915 GND 0.004182f
C5620 VDD.n2916 GND 0.004182f
C5621 VDD.n2917 GND 0.004182f
C5622 VDD.n2918 GND 0.004182f
C5623 VDD.n2919 GND 0.004182f
C5624 VDD.n2920 GND 0.004182f
C5625 VDD.n2921 GND 0.004182f
C5626 VDD.n2922 GND 0.004182f
C5627 VDD.n2923 GND 0.004182f
C5628 VDD.n2924 GND 0.004182f
C5629 VDD.n2925 GND 0.004182f
C5630 VDD.n2926 GND 0.004182f
C5631 VDD.n2927 GND 0.004182f
C5632 VDD.n2928 GND 0.004182f
C5633 VDD.n2929 GND 0.004182f
C5634 VDD.n2930 GND 0.004182f
C5635 VDD.n2931 GND 0.004182f
C5636 VDD.n2932 GND 0.004182f
C5637 VDD.n2933 GND 0.004182f
C5638 VDD.n2934 GND 0.004182f
C5639 VDD.n2935 GND 0.004182f
C5640 VDD.n2936 GND 0.004182f
C5641 VDD.n2937 GND 0.004182f
C5642 VDD.n2938 GND 0.004182f
C5643 VDD.n2939 GND 0.004182f
C5644 VDD.n2940 GND 0.004182f
C5645 VDD.n2941 GND 0.004182f
C5646 VDD.n2942 GND 0.004182f
C5647 VDD.n2943 GND 0.004182f
C5648 VDD.n2944 GND 0.004182f
C5649 VDD.n2945 GND 0.004182f
C5650 VDD.n2946 GND 0.004182f
C5651 VDD.n2947 GND 0.004182f
C5652 VDD.n2948 GND 0.004182f
C5653 VDD.n2949 GND 0.004182f
C5654 VDD.n2950 GND 0.004182f
C5655 VDD.n2951 GND 0.004182f
C5656 VDD.n2952 GND 0.004182f
C5657 VDD.n2953 GND 0.004182f
C5658 VDD.n2954 GND 0.004182f
C5659 VDD.n2955 GND 0.004182f
C5660 VDD.n2956 GND 0.004182f
C5661 VDD.n2957 GND 0.004182f
C5662 VDD.n2958 GND 0.004182f
C5663 VDD.n2959 GND 0.004182f
C5664 VDD.n2960 GND 0.004182f
C5665 VDD.n2961 GND 0.004182f
C5666 VDD.n2962 GND 0.004182f
C5667 VDD.n2963 GND 0.004182f
C5668 VDD.n2964 GND 0.004182f
C5669 VDD.n2965 GND 0.004182f
C5670 VDD.n2966 GND 0.004182f
C5671 VDD.n2967 GND 0.004182f
C5672 VDD.n2968 GND 0.004182f
C5673 VDD.n2969 GND 0.004182f
C5674 VDD.n2970 GND 0.004182f
C5675 VDD.n2971 GND 0.004182f
C5676 VDD.n2972 GND 0.004182f
C5677 VDD.n2973 GND 0.004182f
C5678 VDD.n2974 GND 0.004182f
C5679 VDD.n2975 GND 0.004182f
C5680 VDD.n2976 GND 0.004182f
C5681 VDD.n2977 GND 0.004182f
C5682 VDD.n2978 GND 0.004182f
C5683 VDD.n2979 GND 0.004182f
C5684 VDD.n2980 GND 0.004182f
C5685 VDD.n2981 GND 0.004182f
C5686 VDD.n2982 GND 0.004182f
C5687 VDD.n2983 GND 0.004182f
C5688 VDD.n2984 GND 0.004182f
C5689 VDD.n2985 GND 0.004182f
C5690 VDD.n2986 GND 0.004182f
C5691 VDD.n2987 GND 0.004182f
C5692 VDD.n2988 GND 0.004182f
C5693 VDD.n2989 GND 0.004182f
C5694 VDD.n2990 GND 0.004182f
C5695 VDD.n2991 GND 0.004182f
C5696 VDD.n2992 GND 0.004182f
C5697 VDD.n2993 GND 0.004182f
C5698 VDD.n2994 GND 0.004182f
C5699 VDD.n2995 GND 0.004182f
C5700 VDD.n2996 GND 0.004182f
C5701 VDD.n2997 GND 0.004182f
C5702 VDD.n2998 GND 0.004182f
C5703 VDD.n2999 GND 0.004182f
C5704 VDD.n3000 GND 0.004182f
C5705 VDD.n3001 GND 0.004182f
C5706 VDD.n3002 GND 0.004182f
C5707 VDD.n3003 GND 0.004182f
C5708 VDD.n3004 GND 0.004182f
C5709 VDD.n3005 GND 0.004182f
C5710 VDD.n3006 GND 0.004182f
C5711 VDD.n3007 GND 0.004182f
C5712 VDD.n3008 GND 0.004182f
C5713 VDD.n3009 GND 0.004182f
C5714 VDD.n3010 GND 0.004182f
C5715 VDD.n3011 GND 0.004182f
C5716 VDD.n3012 GND 0.004182f
C5717 VDD.n3013 GND 0.004182f
C5718 VDD.n3014 GND 0.004182f
C5719 VDD.n3015 GND 0.004182f
C5720 VDD.n3016 GND 0.004182f
C5721 VDD.n3017 GND 0.004182f
C5722 VDD.n3018 GND 0.004182f
C5723 VDD.n3019 GND 0.004182f
C5724 VDD.n3020 GND 0.004182f
C5725 VDD.n3021 GND 0.004182f
C5726 VDD.n3022 GND 0.004182f
C5727 VDD.n3023 GND 0.004182f
C5728 VDD.n3024 GND 0.004182f
C5729 VDD.n3025 GND 0.004182f
C5730 VDD.n3026 GND 0.08226f
C5731 VDD.n3027 GND 0.004182f
C5732 VDD.n3028 GND 0.004182f
C5733 VDD.n3029 GND 0.004182f
C5734 VDD.n3030 GND 0.004182f
C5735 VDD.n3031 GND 0.004182f
C5736 VDD.n3032 GND 0.004182f
C5737 VDD.n3033 GND 0.004182f
C5738 VDD.n3034 GND 0.004182f
C5739 VDD.n3035 GND 0.004182f
C5740 VDD.n3036 GND 0.004182f
C5741 VDD.n3037 GND 0.004182f
C5742 VDD.n3038 GND 0.004182f
C5743 VDD.n3039 GND 0.004182f
C5744 VDD.n3040 GND 0.004182f
C5745 VDD.n3041 GND 0.004182f
C5746 VDD.n3042 GND 0.004182f
C5747 VDD.n3043 GND 0.004182f
C5748 VDD.n3044 GND 0.004182f
C5749 VDD.n3045 GND 0.004182f
C5750 VDD.n3046 GND 0.004182f
C5751 VDD.n3047 GND 0.004182f
C5752 VDD.n3048 GND 0.004182f
C5753 VDD.n3049 GND 0.004182f
C5754 VDD.n3050 GND 0.004182f
C5755 VDD.n3051 GND 0.004182f
C5756 VDD.n3052 GND 0.004182f
C5757 VDD.n3053 GND 0.004182f
C5758 VDD.n3054 GND 0.004182f
C5759 VDD.n3055 GND 0.004182f
C5760 VDD.n3056 GND 0.004182f
C5761 VDD.n3057 GND 0.004182f
C5762 VDD.n3058 GND 0.004182f
C5763 VDD.n3059 GND 0.004182f
C5764 VDD.n3060 GND 0.004182f
C5765 VDD.n3061 GND 0.004182f
C5766 VDD.n3062 GND 0.004182f
C5767 VDD.n3063 GND 0.004182f
C5768 VDD.n3064 GND 0.004182f
C5769 VDD.n3065 GND 0.004182f
C5770 VDD.n3066 GND 0.004182f
C5771 VDD.n3067 GND 0.004182f
C5772 VDD.n3068 GND 0.004182f
C5773 VDD.n3069 GND 0.004182f
C5774 VDD.n3070 GND 0.004182f
C5775 VDD.n3071 GND 0.004182f
C5776 VDD.n3072 GND 0.004182f
C5777 VDD.n3073 GND 0.004182f
C5778 VDD.n3074 GND 0.004182f
C5779 VDD.n3075 GND 0.004182f
C5780 VDD.n3076 GND 0.004182f
C5781 VDD.n3077 GND 0.004182f
C5782 VDD.n3078 GND 0.004182f
C5783 VDD.n3079 GND 0.004182f
C5784 VDD.n3080 GND 0.004182f
C5785 VDD.n3081 GND 0.004182f
C5786 VDD.n3082 GND 0.004182f
C5787 VDD.n3083 GND 0.004182f
C5788 VDD.n3084 GND 0.004182f
C5789 VDD.n3085 GND 0.004182f
C5790 VDD.n3086 GND 0.004182f
C5791 VDD.n3087 GND 0.004182f
C5792 VDD.n3088 GND 0.004182f
C5793 VDD.n3089 GND 0.004182f
C5794 VDD.n3090 GND 0.004182f
C5795 VDD.n3091 GND 0.004182f
C5796 VDD.n3092 GND 0.004182f
C5797 VDD.n3093 GND 0.004182f
C5798 VDD.n3094 GND 0.004182f
C5799 VDD.n3095 GND 0.004182f
C5800 VDD.n3096 GND 0.004182f
C5801 VDD.n3097 GND 0.004182f
C5802 VDD.n3098 GND 0.004182f
C5803 VDD.n3099 GND 0.004182f
C5804 VDD.n3100 GND 0.004182f
C5805 VDD.n3101 GND 0.004182f
C5806 VDD.n3102 GND 0.004182f
C5807 VDD.n3103 GND 0.004182f
C5808 VDD.n3104 GND 0.004182f
C5809 VDD.n3105 GND 0.004182f
C5810 VDD.n3106 GND 0.004182f
C5811 VDD.n3107 GND 0.004182f
C5812 VDD.n3108 GND 0.004182f
C5813 VDD.n3109 GND 0.004182f
C5814 VDD.n3110 GND 0.004182f
C5815 VDD.n3111 GND 0.004182f
C5816 VDD.n3112 GND 0.004182f
C5817 VDD.n3113 GND 0.004182f
C5818 VDD.n3114 GND 0.004182f
C5819 VDD.n3115 GND 0.004182f
C5820 VDD.n3116 GND 0.004182f
C5821 VDD.n3117 GND 0.004182f
C5822 VDD.n3118 GND 0.004182f
C5823 VDD.n3119 GND 0.004182f
C5824 VDD.n3120 GND 0.004182f
C5825 VDD.n3121 GND 0.004182f
C5826 VDD.n3122 GND 0.004182f
C5827 VDD.n3123 GND 0.009324f
C5828 VDD.n3124 GND 0.009324f
C5829 VDD.n3125 GND 0.009616f
C5830 VDD.n3126 GND 0.009616f
C5831 VDD.n3127 GND 0.004182f
C5832 VDD.n3128 GND 0.004182f
C5833 VDD.n3129 GND 0.004182f
C5834 VDD.n3130 GND 0.004182f
C5835 VDD.n3131 GND 0.002521f
C5836 VDD.n3132 GND 0.004182f
C5837 VDD.n3133 GND 0.004182f
C5838 VDD.n3134 GND 0.003751f
C5839 VDD.n3135 GND 0.004182f
C5840 VDD.n3136 GND 0.004182f
C5841 VDD.n3137 GND 0.004182f
C5842 VDD.n3138 GND 0.004182f
C5843 VDD.n3139 GND 0.004182f
C5844 VDD.n3140 GND 0.004182f
C5845 VDD.n3141 GND 0.004182f
C5846 VDD.n3142 GND 0.004182f
C5847 VDD.n3143 GND 0.004182f
C5848 VDD.n3144 GND 0.004182f
C5849 VDD.n3145 GND 0.004182f
C5850 VDD.n3146 GND 0.004182f
C5851 VDD.n3147 GND 0.004182f
C5852 VDD.n3148 GND 0.004182f
C5853 VDD.n3149 GND 0.004182f
C5854 VDD.n3150 GND 0.004182f
C5855 VDD.n3151 GND 0.004182f
C5856 VDD.n3152 GND 0.004182f
C5857 VDD.n3153 GND 0.004182f
C5858 VDD.n3154 GND 0.004182f
C5859 VDD.n3155 GND 0.004182f
C5860 VDD.n3156 GND 0.004182f
C5861 VDD.n3157 GND 0.004182f
C5862 VDD.n3158 GND 0.004182f
C5863 VDD.n3159 GND 0.004182f
C5864 VDD.n3160 GND 0.004182f
C5865 VDD.n3161 GND 0.004182f
C5866 VDD.n3162 GND 0.004182f
C5867 VDD.n3163 GND 0.004182f
C5868 VDD.n3164 GND 0.004182f
C5869 VDD.n3165 GND 0.004182f
C5870 VDD.n3166 GND 0.004182f
C5871 VDD.n3167 GND 0.004182f
C5872 VDD.n3168 GND 0.004182f
C5873 VDD.n3169 GND 0.004182f
C5874 VDD.n3170 GND 0.004182f
C5875 VDD.n3171 GND 0.009616f
C5876 VDD.n3172 GND 0.009616f
C5877 VDD.n3174 GND 2.08643f
C5878 VDD.n3176 GND 0.009616f
C5879 VDD.n3177 GND 0.009616f
C5880 VDD.n3178 GND 0.009324f
C5881 VDD.n3179 GND 0.004182f
C5882 VDD.n3180 GND 0.004182f
C5883 VDD.n3181 GND 0.339013f
C5884 VDD.n3182 GND 0.004182f
C5885 VDD.n3183 GND 0.004182f
C5886 VDD.n3184 GND 0.004182f
C5887 VDD.n3185 GND 0.004182f
C5888 VDD.n3186 GND 0.004182f
C5889 VDD.n3187 GND 0.339013f
C5890 VDD.n3188 GND 0.004182f
C5891 VDD.n3189 GND 0.004182f
C5892 VDD.n3190 GND 0.004182f
C5893 VDD.n3191 GND 0.004182f
C5894 VDD.n3192 GND 0.004182f
C5895 VDD.n3193 GND 0.339013f
C5896 VDD.n3194 GND 0.004182f
C5897 VDD.n3195 GND 0.004182f
C5898 VDD.n3196 GND 0.004182f
C5899 VDD.n3197 GND 0.004182f
C5900 VDD.n3198 GND 0.004182f
C5901 VDD.n3199 GND 0.211883f
C5902 VDD.n3200 GND 0.004182f
C5903 VDD.n3201 GND 0.004182f
C5904 VDD.n3202 GND 0.004182f
C5905 VDD.n3203 GND 0.004182f
C5906 VDD.n3204 GND 0.004182f
C5907 VDD.n3205 GND 0.306607f
C5908 VDD.n3206 GND 0.004182f
C5909 VDD.n3207 GND 0.004182f
C5910 VDD.n3208 GND 0.004182f
C5911 VDD.n3209 GND 0.004182f
C5912 VDD.n3210 GND 0.004182f
C5913 VDD.n3211 GND 0.339013f
C5914 VDD.n3212 GND 0.004182f
C5915 VDD.n3213 GND 0.004182f
C5916 VDD.n3214 GND 0.004182f
C5917 VDD.n3215 GND 0.004182f
C5918 VDD.n3216 GND 0.004182f
C5919 VDD.n3217 GND 0.339013f
C5920 VDD.n3218 GND 0.004182f
C5921 VDD.n3219 GND 0.004182f
C5922 VDD.n3220 GND 0.004182f
C5923 VDD.n3221 GND 0.004182f
C5924 VDD.n3222 GND 0.004182f
C5925 VDD.n3223 GND 0.339013f
C5926 VDD.n3224 GND 0.004182f
C5927 VDD.n3225 GND 0.004182f
C5928 VDD.n3226 GND 0.004182f
C5929 VDD.n3227 GND 0.004182f
C5930 VDD.n3228 GND 0.004182f
C5931 VDD.n3229 GND 0.339013f
C5932 VDD.n3230 GND 0.004182f
C5933 VDD.n3231 GND 0.004182f
C5934 VDD.n3232 GND 0.004182f
C5935 VDD.n3233 GND 0.004182f
C5936 VDD.n3234 GND 0.004182f
C5937 VDD.n3235 GND 0.271709f
C5938 VDD.n3236 GND 0.004182f
C5939 VDD.n3237 GND 0.004182f
C5940 VDD.n3238 GND 0.004182f
C5941 VDD.n3239 GND 0.004182f
C5942 VDD.n3240 GND 0.004182f
C5943 VDD.n3241 GND 0.339013f
C5944 VDD.n3242 GND 0.004182f
C5945 VDD.n3243 GND 0.004182f
C5946 VDD.n3244 GND 0.004182f
C5947 VDD.n3245 GND 0.004182f
C5948 VDD.n3246 GND 0.004182f
C5949 VDD.n3247 GND 0.339013f
C5950 VDD.n3248 GND 0.004182f
C5951 VDD.n3249 GND 0.004182f
C5952 VDD.n3250 GND 0.004182f
C5953 VDD.n3251 GND 0.004182f
C5954 VDD.n3252 GND 0.004182f
C5955 VDD.n3253 GND 0.206898f
C5956 VDD.n3254 GND 0.004182f
C5957 VDD.n3255 GND 0.004182f
C5958 VDD.n3256 GND 0.004182f
C5959 VDD.n3257 GND 0.004182f
C5960 VDD.n3258 GND 0.004182f
C5961 VDD.n3259 GND 0.339013f
C5962 VDD.n3260 GND 0.004182f
C5963 VDD.n3261 GND 0.004182f
C5964 VDD.n3262 GND 0.004182f
C5965 VDD.n3263 GND 0.004182f
C5966 VDD.n3264 GND 0.004182f
C5967 VDD.n3265 GND 0.339013f
C5968 VDD.n3266 GND 0.004182f
C5969 VDD.n3267 GND 0.004182f
C5970 VDD.n3268 GND 0.004182f
C5971 VDD.n3269 GND 0.004182f
C5972 VDD.n3270 GND 0.004182f
C5973 VDD.n3271 GND 0.339013f
C5974 VDD.n3272 GND 0.004182f
C5975 VDD.n3273 GND 0.004182f
C5976 VDD.n3274 GND 0.004182f
C5977 VDD.n3275 GND 0.004182f
C5978 VDD.n3276 GND 0.004182f
C5979 VDD.n3277 GND 0.261738f
C5980 VDD.n3278 GND 0.004182f
C5981 VDD.n3279 GND 0.004182f
C5982 VDD.n3280 GND 0.004182f
C5983 VDD.n3281 GND 0.004182f
C5984 VDD.n3282 GND 0.004182f
C5985 VDD.n3283 GND 0.339013f
C5986 VDD.n3284 GND 0.004182f
C5987 VDD.n3285 GND 0.004182f
C5988 VDD.n3286 GND 0.004182f
C5989 VDD.n3287 GND 0.004182f
C5990 VDD.n3288 GND 0.004182f
C5991 VDD.n3289 GND 0.339013f
C5992 VDD.n3290 GND 0.004182f
C5993 VDD.n3291 GND 0.004182f
C5994 VDD.n3292 GND 0.004182f
C5995 VDD.n3293 GND 0.004182f
C5996 VDD.n3294 GND 0.004182f
C5997 VDD.n3295 GND 0.326549f
C5998 VDD.n3296 GND 0.004182f
C5999 VDD.n3297 GND 0.004182f
C6000 VDD.n3298 GND 0.004182f
C6001 VDD.n3299 GND 0.004182f
C6002 VDD.n3300 GND 0.004182f
C6003 VDD.n3301 GND 0.339013f
C6004 VDD.n3302 GND 0.004182f
C6005 VDD.n3303 GND 0.004182f
C6006 VDD.n3304 GND 0.004182f
C6007 VDD.n3305 GND 0.004182f
C6008 VDD.n3306 GND 0.004182f
C6009 VDD.n3307 GND 0.339013f
C6010 VDD.n3308 GND 0.004182f
C6011 VDD.n3309 GND 0.004182f
C6012 VDD.n3310 GND 0.004182f
C6013 VDD.n3311 GND 0.004182f
C6014 VDD.n3312 GND 0.004182f
C6015 VDD.n3313 GND 0.221854f
C6016 VDD.n3314 GND 0.004182f
C6017 VDD.n3315 GND 0.004182f
C6018 VDD.n3316 GND 0.004182f
C6019 VDD.n3317 GND 0.004182f
C6020 VDD.n3318 GND 0.004182f
C6021 VDD.n3319 GND 0.339013f
C6022 VDD.n3320 GND 0.004182f
C6023 VDD.n3321 GND 0.004182f
C6024 VDD.n3322 GND 0.004182f
C6025 VDD.n3323 GND 0.004182f
C6026 VDD.n3324 GND 0.004182f
C6027 VDD.n3325 GND 0.339013f
C6028 VDD.n3326 GND 0.004182f
C6029 VDD.n3327 GND 0.004182f
C6030 VDD.n3328 GND 0.004182f
C6031 VDD.n3329 GND 0.004182f
C6032 VDD.n3330 GND 0.004182f
C6033 VDD.n3331 GND 0.18197f
C6034 VDD.n3332 GND 0.004182f
C6035 VDD.n3333 GND 0.004182f
C6036 VDD.n3334 GND 0.004182f
C6037 VDD.n3335 GND 0.004182f
C6038 VDD.n3336 GND 0.004182f
C6039 VDD.n3337 GND 0.339013f
C6040 VDD.n3338 GND 0.004182f
C6041 VDD.n3339 GND 0.004182f
C6042 VDD.n3340 GND 0.004182f
C6043 VDD.n3341 GND 0.004182f
C6044 VDD.n3342 GND 0.004182f
C6045 VDD.n3343 GND 0.339013f
C6046 VDD.n3344 GND 0.004182f
C6047 VDD.n3345 GND 0.004182f
C6048 VDD.n3346 GND 0.004182f
C6049 VDD.n3347 GND 0.004182f
C6050 VDD.n3348 GND 0.004182f
C6051 VDD.n3349 GND 0.339013f
C6052 VDD.n3350 GND 0.004182f
C6053 VDD.n3351 GND 0.004182f
C6054 VDD.n3352 GND 0.004182f
C6055 VDD.n3353 GND 0.004182f
C6056 VDD.n3354 GND 0.004182f
C6057 VDD.n3355 GND 0.339013f
C6058 VDD.n3356 GND 0.004182f
C6059 VDD.n3357 GND 0.004182f
C6060 VDD.n3358 GND 0.004182f
C6061 VDD.n3359 GND 0.004182f
C6062 VDD.n3360 GND 0.004182f
C6063 VDD.n3361 GND 0.339013f
C6064 VDD.n3362 GND 0.004182f
C6065 VDD.n3363 GND 0.004182f
C6066 VDD.n3364 GND 0.004182f
C6067 VDD.n3365 GND 0.004182f
C6068 VDD.n3366 GND 0.004182f
C6069 VDD.n3367 GND 0.301622f
C6070 VDD.n3368 GND 0.004182f
C6071 VDD.n3369 GND 0.004182f
C6072 VDD.n3370 GND 0.004182f
C6073 VDD.n3371 GND 0.004182f
C6074 VDD.n3372 GND 0.004182f
C6075 VDD.n3373 GND 0.294144f
C6076 VDD.n3374 GND 0.004182f
C6077 VDD.n3375 GND 0.004182f
C6078 VDD.n3376 GND 0.004182f
C6079 VDD.n3377 GND 0.004182f
C6080 VDD.n3378 GND 0.004182f
C6081 VDD.n3379 GND 0.339013f
C6082 VDD.n3380 GND 0.004182f
C6083 VDD.n3381 GND 0.004182f
C6084 VDD.n3382 GND 0.004182f
C6085 VDD.n3383 GND 0.004182f
C6086 VDD.n3384 GND 0.004182f
C6087 VDD.n3385 GND 0.339013f
C6088 VDD.n3386 GND 0.004182f
C6089 VDD.n3387 GND 0.004182f
C6090 VDD.n3388 GND 0.004182f
C6091 VDD.n3389 GND 0.004182f
C6092 VDD.n3390 GND 0.004182f
C6093 VDD.n3391 GND 0.339013f
C6094 VDD.n3392 GND 0.004182f
C6095 VDD.n3393 GND 0.004182f
C6096 VDD.n3394 GND 0.004182f
C6097 VDD.n3395 GND 0.004182f
C6098 VDD.n3396 GND 0.004182f
C6099 VDD.n3397 GND 0.339013f
C6100 VDD.n3398 GND 0.004182f
C6101 VDD.n3399 GND 0.004182f
C6102 VDD.n3400 GND 0.004182f
C6103 VDD.n3401 GND 0.004182f
C6104 VDD.n3402 GND 0.004182f
C6105 VDD.n3403 GND 0.339013f
C6106 VDD.n3404 GND 0.004182f
C6107 VDD.n3405 GND 0.004182f
C6108 VDD.n3406 GND 0.004182f
C6109 VDD.n3407 GND 0.004182f
C6110 VDD.n3408 GND 0.004182f
C6111 VDD.n3409 GND 0.189448f
C6112 VDD.n3410 GND 0.004182f
C6113 VDD.n3411 GND 0.004182f
C6114 VDD.n3412 GND 0.004182f
C6115 VDD.n3413 GND 0.004182f
C6116 VDD.n3414 GND 0.004182f
C6117 VDD.n3415 GND 0.339013f
C6118 VDD.n3416 GND 0.004182f
C6119 VDD.n3417 GND 0.004182f
C6120 VDD.n3418 GND 0.004182f
C6121 VDD.n3419 GND 0.004182f
C6122 VDD.n3420 GND 0.004182f
C6123 VDD.n3421 GND 0.201912f
C6124 VDD.n3422 GND 0.004182f
C6125 VDD.n3423 GND 0.004182f
C6126 VDD.n3424 GND 0.004182f
C6127 VDD.n3425 GND 0.004182f
C6128 VDD.n3426 GND 0.004182f
C6129 VDD.n3427 GND 0.339013f
C6130 VDD.n3428 GND 0.004182f
C6131 VDD.n3429 GND 0.004182f
C6132 VDD.n3430 GND 0.004182f
C6133 VDD.n3431 GND 0.004182f
C6134 VDD.n3432 GND 0.004182f
C6135 VDD.n3433 GND 0.004182f
C6136 VDD.n3435 GND 0.004182f
C6137 VDD.n3436 GND 0.004182f
C6138 VDD.n3438 GND 0.004182f
C6139 VDD.n3439 GND 0.004182f
C6140 VDD.n3440 GND 0.004182f
C6141 VDD.n3442 GND 0.004182f
C6142 VDD.n3443 GND 0.004182f
C6143 VDD.n3444 GND 0.004182f
C6144 VDD.n3445 GND 0.004182f
C6145 VDD.n3446 GND 0.004182f
C6146 VDD.n3447 GND 0.004182f
C6147 VDD.n3449 GND 0.004182f
C6148 VDD.n3450 GND 0.004182f
C6149 VDD.n3451 GND 0.004182f
C6150 VDD.n3452 GND 0.004182f
C6151 VDD.n3453 GND 0.004182f
C6152 VDD.n3454 GND 0.004182f
C6153 VDD.n3456 GND 0.004182f
C6154 VDD.n3457 GND 0.009616f
C6155 VDD.n3458 GND 0.009616f
C6156 VDD.n3459 GND 0.009324f
C6157 VDD.n3460 GND 0.004182f
C6158 VDD.n3461 GND 0.004182f
C6159 VDD.n3462 GND 0.004182f
C6160 VDD.n3463 GND 0.004182f
C6161 VDD.n3464 GND 0.004182f
C6162 VDD.n3465 GND 0.004182f
C6163 VDD.n3466 GND 0.339013f
C6164 VDD.n3467 GND 0.004182f
C6165 VDD.n3468 GND 0.004182f
C6166 VDD.n3469 GND 0.004182f
C6167 VDD.n3470 GND 0.004182f
C6168 VDD.n3471 GND 0.004182f
C6169 VDD.n3472 GND 0.339013f
C6170 VDD.n3473 GND 0.004182f
C6171 VDD.n3474 GND 0.004182f
C6172 VDD.n3475 GND 0.004182f
C6173 VDD.n3476 GND 0.009844f
C6174 VDD.n3478 GND 0.009616f
C6175 VDD.n3479 GND 0.009096f
C6176 VDD.n3480 GND 0.004182f
C6177 VDD.n3481 GND 0.004182f
C6178 VDD.n3482 GND 0.004182f
C6179 VDD.n3484 GND 0.004182f
C6180 VDD.n3485 GND 0.004182f
C6181 VDD.n3486 GND 0.003751f
C6182 VDD.n3487 GND 0.004182f
C6183 VDD.n3488 GND 0.004182f
C6184 VDD.n3489 GND 0.004182f
C6185 VDD.n3491 GND 0.004182f
C6186 VDD.n3492 GND 0.004182f
C6187 VDD.n3493 GND 0.004182f
C6188 VDD.n3494 GND 0.004182f
C6189 VDD.n3495 GND 0.004182f
C6190 VDD.n3496 GND 0.004182f
C6191 VDD.n3498 GND 0.004182f
C6192 VDD.n3499 GND 0.004182f
C6193 VDD.n3501 GND 0.004182f
C6194 VDD.n3502 GND 0.004182f
C6195 VDD.n3503 GND 0.004182f
C6196 VDD.n3504 GND 0.004182f
C6197 VDD.n3505 GND 0.004182f
C6198 VDD.n3506 GND 0.004182f
C6199 VDD.n3508 GND 0.004182f
C6200 VDD.n3509 GND 0.004182f
C6201 VDD.n3510 GND 0.004182f
C6202 VDD.n3511 GND 0.004182f
C6203 VDD.n3512 GND 0.004182f
C6204 VDD.n3513 GND 0.004182f
C6205 VDD.n3515 GND 0.004182f
C6206 VDD.n3516 GND 0.004182f
C6207 VDD.n3518 GND 0.004182f
C6208 VDD.n3519 GND 0.004182f
C6209 VDD.n3520 GND 0.009616f
C6210 VDD.n3521 GND 0.009324f
C6211 VDD.n3522 GND 0.009324f
C6212 VDD.n3523 GND 0.334027f
C6213 VDD.n3524 GND 0.009324f
C6214 VDD.n3525 GND 0.009616f
C6215 VDD.n3526 GND 0.009096f
C6216 VDD.n3527 GND 0.004182f
C6217 VDD.n3528 GND 0.004182f
C6218 VDD.n3529 GND 0.004182f
C6219 VDD.n3531 GND 0.004182f
C6220 VDD.n3532 GND 0.004182f
C6221 VDD.n3533 GND 0.003751f
C6222 VDD.n3534 GND 0.004182f
C6223 VDD.n3535 GND 0.004182f
C6224 VDD.n3536 GND 0.004182f
C6225 VDD.n3538 GND 0.004182f
C6226 VDD.n3539 GND 0.004182f
C6227 VDD.n3540 GND 0.004182f
C6228 VDD.n3541 GND 0.004182f
C6229 VDD.n3542 GND 0.004182f
C6230 VDD.n3543 GND 0.004182f
C6231 VDD.n3545 GND 0.004182f
C6232 VDD.n3546 GND 0.004182f
C6233 VDD.n3547 GND 0.05129f
C6234 VDD.n3548 GND 0.954066f
C6235 VDD.t12 GND 0.179673f
C6236 VDD.t9 GND 0.743196f
C6237 VDD.n3549 GND 0.095879f
C6238 VDD.t11 GND 0.131174f
C6239 VDD.n3550 GND 0.098395f
C6240 VDD.n3551 GND 0.004949f
C6241 VDD.n3552 GND 0.006149f
C6242 VDD.n3553 GND 0.004949f
C6243 VDD.n3554 GND 0.006149f
C6244 VDD.n3555 GND 0.004949f
C6245 VDD.n3556 GND 0.006149f
C6246 VDD.n3557 GND 0.002574f
C6247 VDD.n3558 GND 0.006149f
C6248 VDD.n3559 GND 0.004949f
C6249 VDD.n3560 GND 0.006149f
C6250 VDD.n3561 GND 0.004949f
C6251 VDD.n3562 GND 0.006149f
C6252 VDD.n3563 GND 0.004949f
C6253 VDD.n3564 GND 0.006149f
C6254 VDD.n3565 GND 0.003984f
C6255 VDD.n3566 GND 0.006149f
C6256 VDD.n3567 GND 0.004949f
C6257 VDD.n3568 GND 0.006149f
C6258 VDD.n3569 GND 0.004949f
C6259 VDD.n3570 GND 0.006149f
C6260 VDD.n3571 GND 0.006149f
C6261 VDD.n3572 GND 0.004949f
C6262 VDD.n3573 GND 0.006149f
C6263 VDD.n3574 GND 0.006149f
C6264 VDD.n3575 GND 0.006149f
C6265 VDD.n3576 GND 0.004949f
C6266 VDD.n3577 GND 0.006149f
C6267 VDD.n3578 GND 0.006149f
C6268 VDD.n3579 GND 0.004949f
C6269 VDD.n3580 GND 0.006149f
C6270 VDD.n3581 GND 0.006149f
C6271 VDD.n3582 GND 0.004949f
C6272 VDD.n3583 GND 0.006149f
C6273 VDD.n3584 GND 0.006149f
C6274 VDD.n3585 GND 0.006149f
C6275 VDD.n3586 GND 0.004949f
C6276 VDD.n3587 GND 0.006149f
C6277 VDD.n3588 GND 0.006149f
C6278 VDD.n3589 GND 0.004281f
C6279 VDD.n3590 GND 0.006149f
C6280 VDD.n3591 GND 0.006149f
C6281 VDD.t66 GND 0.179673f
C6282 VDD.t64 GND 0.743196f
C6283 VDD.n3592 GND 0.095879f
C6284 VDD.t65 GND 0.131174f
C6285 VDD.n3593 GND 0.098395f
C6286 VDD.n3594 GND 0.00928f
C6287 VDD.n3595 GND 0.006149f
C6288 VDD.n3596 GND 0.006149f
C6289 VDD.n3597 GND 0.006149f
C6290 VDD.n3598 GND 0.004949f
C6291 VDD.n3599 GND 0.006149f
C6292 VDD.n3600 GND 0.006149f
C6293 VDD.n3601 GND 0.004949f
C6294 VDD.n3602 GND 0.006149f
C6295 VDD.n3603 GND 0.006149f
C6296 VDD.n3604 GND 0.004949f
C6297 VDD.n3605 GND 0.006149f
C6298 VDD.n3606 GND 0.006149f
C6299 VDD.n3607 GND 0.006149f
C6300 VDD.n3608 GND 0.004949f
C6301 VDD.n3609 GND 0.006149f
C6302 VDD.n3610 GND 0.006149f
C6303 VDD.n3611 GND 0.004949f
C6304 VDD.n3612 GND 0.006149f
C6305 VDD.n3613 GND 0.006149f
C6306 VDD.n3614 GND 0.004949f
C6307 VDD.n3615 GND 0.006149f
C6308 VDD.n3616 GND 0.006149f
C6309 VDD.n3617 GND 0.006149f
C6310 VDD.n3618 GND 0.004949f
C6311 VDD.n3619 GND 0.006149f
C6312 VDD.n3620 GND 0.006149f
C6313 VDD.n3621 GND 0.004949f
C6314 VDD.n3622 GND 0.006149f
C6315 VDD.n3623 GND 0.006149f
C6316 VDD.n3624 GND 0.004949f
C6317 VDD.n3625 GND 0.006149f
C6318 VDD.n3626 GND 0.006149f
C6319 VDD.n3627 GND 0.006149f
C6320 VDD.n3628 GND 0.004949f
C6321 VDD.n3629 GND 0.006149f
C6322 VDD.n3630 GND 0.006149f
C6323 VDD.n3631 GND 0.004949f
C6324 VDD.t69 GND 0.179673f
C6325 VDD.t67 GND 0.743196f
C6326 VDD.n3632 GND 0.095879f
C6327 VDD.t68 GND 0.131174f
C6328 VDD.n3633 GND 0.098395f
C6329 VDD.n3634 GND 0.006806f
C6330 VDD.n3635 GND 0.006149f
C6331 VDD.n3636 GND 0.006149f
C6332 VDD.n3637 GND 0.003217f
C6333 VDD.n3638 GND 0.006149f
C6334 VDD.n3639 GND 0.006149f
C6335 VDD.n3640 GND 0.006149f
C6336 VDD.n3641 GND 0.004949f
C6337 VDD.n3642 GND 0.006149f
C6338 VDD.n3643 GND 0.006149f
C6339 VDD.n3644 GND 0.004949f
C6340 VDD.n3645 GND 0.006149f
C6341 VDD.n3646 GND 0.006149f
C6342 VDD.n3647 GND 0.004949f
C6343 VDD.n3648 GND 0.006149f
C6344 VDD.n3649 GND 0.006149f
C6345 VDD.n3650 GND 0.006149f
C6346 VDD.n3651 GND 0.004949f
C6347 VDD.n3652 GND 0.006149f
C6348 VDD.n3653 GND 0.006149f
C6349 VDD.n3654 GND 0.004949f
C6350 VDD.n3655 GND 0.006149f
C6351 VDD.n3656 GND 0.006149f
C6352 VDD.n3657 GND 0.004949f
C6353 VDD.n3658 GND 0.006149f
C6354 VDD.n3659 GND 0.006149f
C6355 VDD.n3660 GND 0.006149f
C6356 VDD.n3661 GND 0.004949f
C6357 VDD.n3662 GND 0.006149f
C6358 VDD.n3663 GND 0.006149f
C6359 VDD.n3664 GND 0.004949f
C6360 VDD.n3665 GND 0.006149f
C6361 VDD.n3666 GND 0.006149f
C6362 VDD.n3667 GND 0.004949f
C6363 VDD.n3668 GND 0.006149f
C6364 VDD.n3669 GND 0.006149f
C6365 VDD.n3670 GND 0.004305f
C6366 VDD.n3671 GND 0.004949f
C6367 VDD.n3672 GND 0.006149f
C6368 VDD.n3673 GND 0.006149f
C6369 VDD.n3674 GND 0.004949f
C6370 VDD.n3676 GND 0.006149f
C6371 VDD.n3677 GND 0.004628f
C6372 VDD.n3678 GND 0.00928f
C6373 VDD.n3679 GND 0.002751f
C6374 VDD.n3680 GND 0.014186f
C6375 VDD.n3682 GND 0.006149f
C6376 VDD.n3683 GND 0.004949f
C6377 VDD.n3684 GND 0.004949f
C6378 VDD.n3685 GND 0.006149f
C6379 VDD.n3686 GND 0.014243f
C6380 VDD.n3688 GND 3.71917f
C6381 VDD.n3690 GND 0.006149f
C6382 VDD.n3691 GND 0.004949f
C6383 VDD.n3692 GND 0.004305f
C6384 VDD.n3693 GND 0.954066f
C6385 VDD.n3694 GND 0.012337f
C6386 VDD.n3695 GND 0.006149f
C6387 VDD.n3696 GND 0.004949f
C6388 VDD.n3697 GND 0.006149f
C6389 VDD.n3698 GND 0.498548f
C6390 VDD.n3699 GND 0.006149f
C6391 VDD.n3700 GND 0.004949f
C6392 VDD.n3701 GND 0.006149f
C6393 VDD.n3702 GND 0.006149f
C6394 VDD.n3703 GND 0.006149f
C6395 VDD.n3704 GND 0.004949f
C6396 VDD.n3705 GND 0.006149f
C6397 VDD.n3706 GND 0.498548f
C6398 VDD.n3707 GND 0.006149f
C6399 VDD.n3708 GND 0.004949f
C6400 VDD.n3709 GND 0.006149f
C6401 VDD.n3710 GND 0.006149f
C6402 VDD.n3711 GND 0.006149f
C6403 VDD.n3712 GND 0.004949f
C6404 VDD.n3713 GND 0.006149f
C6405 VDD.n3714 GND 0.498548f
C6406 VDD.n3715 GND 0.006149f
C6407 VDD.n3716 GND 0.004949f
C6408 VDD.n3717 GND 0.006149f
C6409 VDD.n3718 GND 0.006149f
C6410 VDD.n3719 GND 0.006149f
C6411 VDD.n3720 GND 0.004949f
C6412 VDD.n3721 GND 0.006149f
C6413 VDD.n3722 GND 0.40881f
C6414 VDD.n3723 GND 0.006149f
C6415 VDD.n3724 GND 0.004949f
C6416 VDD.n3725 GND 0.006149f
C6417 VDD.n3726 GND 0.006149f
C6418 VDD.n3727 GND 0.006149f
C6419 VDD.n3728 GND 0.004949f
C6420 VDD.n3729 GND 0.006149f
C6421 VDD.n3730 GND 0.498548f
C6422 VDD.n3731 GND 0.006149f
C6423 VDD.n3732 GND 0.004949f
C6424 VDD.n3733 GND 0.006149f
C6425 VDD.n3734 GND 0.006149f
C6426 VDD.n3735 GND 0.006149f
C6427 VDD.n3736 GND 0.004949f
C6428 VDD.n3737 GND 0.006149f
C6429 VDD.n3738 GND 0.498548f
C6430 VDD.n3739 GND 0.006149f
C6431 VDD.n3740 GND 0.004949f
C6432 VDD.n3741 GND 0.006149f
C6433 VDD.n3742 GND 0.006149f
C6434 VDD.n3743 GND 0.006149f
C6435 VDD.n3744 GND 0.004949f
C6436 VDD.n3745 GND 0.006149f
C6437 VDD.n3746 GND 0.498548f
C6438 VDD.n3747 GND 0.006149f
C6439 VDD.n3748 GND 0.004949f
C6440 VDD.n3749 GND 0.006149f
C6441 VDD.n3750 GND 0.006149f
C6442 VDD.n3751 GND 0.006149f
C6443 VDD.n3752 GND 0.004949f
C6444 VDD.n3753 GND 0.006149f
C6445 VDD.n3754 GND 0.498548f
C6446 VDD.n3755 GND 0.006149f
C6447 VDD.n3756 GND 0.004949f
C6448 VDD.n3757 GND 0.006149f
C6449 VDD.n3758 GND 0.006149f
C6450 VDD.n3759 GND 0.006149f
C6451 VDD.n3760 GND 0.004949f
C6452 VDD.n3761 GND 0.006149f
C6453 VDD.n3762 GND 0.498548f
C6454 VDD.n3763 GND 0.006149f
C6455 VDD.n3764 GND 0.004949f
C6456 VDD.n3765 GND 0.006149f
C6457 VDD.n3766 GND 0.006149f
C6458 VDD.n3767 GND 0.006149f
C6459 VDD.n3768 GND 0.004949f
C6460 VDD.n3769 GND 0.006149f
C6461 VDD.n3770 GND 0.498548f
C6462 VDD.n3771 GND 0.006149f
C6463 VDD.n3772 GND 0.004949f
C6464 VDD.n3773 GND 0.006149f
C6465 VDD.n3774 GND 0.006149f
C6466 VDD.n3775 GND 0.006149f
C6467 VDD.n3776 GND 0.004949f
C6468 VDD.n3777 GND 0.006149f
C6469 VDD.t81 GND 0.498548f
C6470 VDD.n3778 GND 0.006149f
C6471 VDD.n3779 GND 0.004949f
C6472 VDD.n3780 GND 0.006149f
C6473 VDD.n3781 GND 0.006149f
C6474 VDD.n3782 GND 0.006149f
C6475 VDD.n3783 GND 0.004949f
C6476 VDD.n3784 GND 0.006149f
C6477 VDD.n3785 GND 0.498548f
C6478 VDD.n3786 GND 0.006149f
C6479 VDD.n3787 GND 0.004949f
C6480 VDD.n3788 GND 0.006149f
C6481 VDD.n3789 GND 0.006149f
C6482 VDD.n3790 GND 0.006149f
C6483 VDD.n3791 GND 0.004949f
C6484 VDD.n3792 GND 0.006149f
C6485 VDD.n3793 GND 0.498548f
C6486 VDD.n3794 GND 0.006149f
C6487 VDD.n3795 GND 0.004949f
C6488 VDD.n3796 GND 0.006149f
C6489 VDD.n3797 GND 0.006149f
C6490 VDD.n3798 GND 0.006149f
C6491 VDD.n3799 GND 0.004949f
C6492 VDD.n3800 GND 0.006149f
C6493 VDD.n3801 GND 0.498548f
C6494 VDD.n3802 GND 0.006149f
C6495 VDD.n3803 GND 0.004949f
C6496 VDD.n3804 GND 0.006149f
C6497 VDD.n3805 GND 0.006149f
C6498 VDD.n3806 GND 0.006149f
C6499 VDD.n3807 GND 0.004949f
C6500 VDD.n3808 GND 0.006149f
C6501 VDD.n3809 GND 0.498548f
C6502 VDD.n3810 GND 0.006149f
C6503 VDD.n3811 GND 0.004949f
C6504 VDD.n3812 GND 0.006149f
C6505 VDD.n3813 GND 0.006149f
C6506 VDD.n3814 GND 0.006149f
C6507 VDD.n3815 GND 0.004949f
C6508 VDD.n3816 GND 0.006149f
C6509 VDD.n3817 GND 0.448694f
C6510 VDD.n3818 GND 0.498548f
C6511 VDD.n3819 GND 0.006149f
C6512 VDD.n3820 GND 0.004949f
C6513 VDD.n3821 GND 0.006149f
C6514 VDD.n3822 GND 0.006149f
C6515 VDD.n3823 GND 0.006149f
C6516 VDD.n3824 GND 0.004949f
C6517 VDD.n3825 GND 0.006149f
C6518 VDD.n3826 GND 0.299129f
C6519 VDD.n3827 GND 0.006149f
C6520 VDD.n3828 GND 0.004949f
C6521 VDD.n3829 GND 0.006149f
C6522 VDD.n3830 GND 0.006149f
C6523 VDD.n3831 GND 0.006149f
C6524 VDD.n3832 GND 0.004949f
C6525 VDD.n3833 GND 0.006149f
C6526 VDD.n3834 GND 0.498548f
C6527 VDD.n3835 GND 0.006149f
C6528 VDD.n3836 GND 0.004949f
C6529 VDD.n3837 GND 0.006149f
C6530 VDD.n3838 GND 0.006149f
C6531 VDD.n3839 GND 0.006149f
C6532 VDD.n3840 GND 0.004949f
C6533 VDD.n3841 GND 0.006149f
C6534 VDD.n3842 GND 0.498548f
C6535 VDD.n3843 GND 0.006149f
C6536 VDD.n3844 GND 0.004949f
C6537 VDD.n3845 GND 0.006149f
C6538 VDD.n3846 GND 0.006149f
C6539 VDD.n3847 GND 0.006149f
C6540 VDD.n3848 GND 0.004949f
C6541 VDD.n3849 GND 0.006149f
C6542 VDD.n3850 GND 0.498548f
C6543 VDD.n3851 GND 0.006149f
C6544 VDD.n3852 GND 0.004949f
C6545 VDD.n3853 GND 0.006149f
C6546 VDD.n3854 GND 0.006149f
C6547 VDD.n3855 GND 0.006149f
C6548 VDD.n3856 GND 0.004949f
C6549 VDD.n3857 GND 0.006149f
C6550 VDD.n3858 GND 0.498548f
C6551 VDD.n3859 GND 0.006149f
C6552 VDD.n3860 GND 0.004949f
C6553 VDD.n3861 GND 0.006149f
C6554 VDD.n3862 GND 0.006149f
C6555 VDD.n3863 GND 0.006149f
C6556 VDD.n3864 GND 0.006149f
C6557 VDD.n3865 GND 0.004949f
C6558 VDD.n3866 GND 0.004949f
C6559 VDD.n3867 GND 0.006149f
C6560 VDD.n3868 GND 0.398839f
C6561 VDD.n3869 GND 0.498548f
C6562 VDD.n3870 GND 0.006149f
C6563 VDD.n3871 GND 0.004949f
C6564 VDD.n3872 GND 0.006149f
C6565 VDD.n3873 GND 0.006149f
C6566 VDD.n3874 GND 0.006149f
C6567 VDD.n3875 GND 0.004949f
C6568 VDD.n3876 GND 0.006149f
C6569 VDD.n3877 GND 0.348984f
C6570 VDD.n3878 GND 0.006149f
C6571 VDD.n3879 GND 0.006149f
C6572 VDD.n3880 GND 0.004949f
C6573 VDD.n3881 GND 0.006149f
C6574 VDD.n3882 GND 0.006149f
C6575 VDD.n3883 GND 0.006149f
C6576 VDD.n3884 GND 0.004949f
C6577 VDD.n3885 GND 0.006149f
C6578 VDD.n3886 GND 0.498548f
C6579 VDD.n3887 GND 0.498548f
C6580 VDD.n3888 GND 0.006149f
C6581 VDD.n3889 GND 0.004949f
C6582 VDD.n3890 GND 0.006149f
C6583 VDD.n3891 GND 0.006149f
C6584 VDD.n3892 GND 0.006149f
C6585 VDD.n3893 GND 0.004949f
C6586 VDD.n3894 GND 0.006149f
C6587 VDD.n3895 GND 0.006149f
C6588 VDD.n3896 GND 0.498548f
C6589 VDD.n3897 GND 0.006149f
C6590 VDD.n3898 GND 0.004949f
C6591 VDD.n3899 GND 0.006149f
C6592 VDD.n3900 GND 0.006149f
C6593 VDD.n3901 GND 0.006149f
C6594 VDD.n3902 GND 0.004949f
C6595 VDD.n3903 GND 0.004949f
C6596 VDD.n3904 GND 0.004949f
C6597 VDD.n3905 GND 0.006149f
C6598 VDD.n3906 GND 0.006149f
C6599 VDD.n3907 GND 0.006149f
C6600 VDD.n3908 GND 0.004949f
C6601 VDD.n3909 GND 0.004949f
C6602 VDD.n3910 GND 0.004949f
C6603 VDD.n3911 GND 0.006149f
C6604 VDD.n3912 GND 0.006149f
C6605 VDD.n3913 GND 0.006149f
C6606 VDD.n3914 GND 0.004949f
C6607 VDD.n3915 GND 0.004949f
C6608 VDD.n3916 GND 0.004949f
C6609 VDD.n3917 GND 0.006149f
C6610 VDD.n3918 GND 0.006149f
C6611 VDD.n3919 GND 0.006149f
C6612 VDD.n3920 GND 0.004949f
C6613 VDD.n3921 GND 0.004949f
C6614 VDD.n3922 GND 0.004949f
C6615 VDD.n3923 GND 0.006149f
C6616 VDD.n3924 GND 0.006149f
C6617 VDD.n3925 GND 0.006149f
C6618 VDD.n3926 GND 0.004949f
C6619 VDD.n3927 GND 0.004949f
C6620 VDD.n3928 GND 0.004949f
C6621 VDD.n3929 GND 0.006149f
C6622 VDD.n3930 GND 0.006149f
C6623 VDD.n3931 GND 0.006149f
C6624 VDD.n3932 GND 0.004949f
C6625 VDD.n3933 GND 0.004949f
C6626 VDD.n3934 GND 0.004949f
C6627 VDD.n3935 GND 0.006149f
C6628 VDD.n3936 GND 0.006149f
C6629 VDD.n3937 GND 0.006149f
C6630 VDD.n3938 GND 0.004949f
C6631 VDD.n3939 GND 0.004949f
C6632 VDD.n3940 GND 0.004949f
C6633 VDD.n3941 GND 0.006149f
C6634 VDD.n3942 GND 0.006149f
C6635 VDD.n3943 GND 0.006149f
C6636 VDD.n3944 GND 0.006149f
C6637 VDD.n3945 GND 0.006149f
C6638 VDD.n3946 GND 0.004949f
C6639 VDD.n3947 GND 0.006149f
C6640 VDD.n3948 GND 0.498548f
C6641 VDD.n3949 GND 0.006149f
C6642 VDD.n3950 GND 0.006149f
C6643 VDD.n3951 GND 0.006149f
C6644 VDD.n3952 GND 0.006149f
C6645 VDD.n3953 GND 0.006149f
C6646 VDD.n3954 GND 0.004949f
C6647 VDD.n3955 GND 0.006149f
C6648 VDD.n3956 GND 0.006149f
C6649 VDD.n3957 GND 0.006149f
C6650 VDD.n3958 GND 0.006149f
C6651 VDD.n3959 GND 0.498548f
C6652 VDD.n3960 GND 0.006149f
C6653 VDD.n3961 GND 0.006149f
C6654 VDD.n3962 GND 0.006149f
C6655 VDD.n3963 GND 0.006149f
C6656 VDD.n3964 GND 0.006149f
C6657 VDD.n3965 GND 0.004949f
C6658 VDD.n3966 GND 0.006149f
C6659 VDD.n3967 GND 0.006149f
C6660 VDD.n3968 GND 0.006149f
C6661 VDD.n3969 GND 0.006149f
C6662 VDD.n3970 GND 0.498548f
C6663 VDD.n3971 GND 0.006149f
C6664 VDD.n3972 GND 0.006149f
C6665 VDD.n3973 GND 0.006149f
C6666 VDD.n3974 GND 0.006149f
C6667 VDD.n3975 GND 0.006149f
C6668 VDD.n3976 GND 0.004949f
C6669 VDD.n3977 GND 0.006149f
C6670 VDD.n3978 GND 0.006149f
C6671 VDD.n3979 GND 0.006149f
C6672 VDD.n3980 GND 0.006149f
C6673 VDD.t22 GND 0.249274f
C6674 VDD.n3981 GND 0.006149f
C6675 VDD.n3982 GND 0.006149f
C6676 VDD.n3983 GND 0.006149f
C6677 VDD.n3984 GND 0.006149f
C6678 VDD.n3985 GND 0.006149f
C6679 VDD.n3986 GND 0.004949f
C6680 VDD.n3987 GND 0.006149f
C6681 VDD.n3988 GND 0.339013f
C6682 VDD.n3989 GND 0.006149f
C6683 VDD.n3990 GND 0.006149f
C6684 VDD.n3991 GND 0.006149f
C6685 VDD.n3992 GND 0.498548f
C6686 VDD.n3993 GND 0.006149f
C6687 VDD.n3994 GND 0.006149f
C6688 VDD.n3995 GND 0.006149f
C6689 VDD.n3996 GND 0.006149f
C6690 VDD.n3997 GND 0.006149f
C6691 VDD.n3998 GND 0.004108f
C6692 VDD.n3999 GND 0.013778f
C6693 VDD.n4000 GND 0.006149f
C6694 VDD.n4001 GND 0.013778f
C6695 VDD.n4026 GND 0.006149f
C6696 VDD.n4027 GND 0.013778f
C6697 VDD.n4028 GND 0.01414f
C6698 VDD.n4029 GND 0.004949f
C6699 VDD.n4030 GND 0.006149f
C6700 VDD.n4031 GND 0.006149f
C6701 VDD.n4032 GND 0.006149f
C6702 VDD.n4033 GND 0.006149f
C6703 VDD.n4034 GND 0.006149f
C6704 VDD.n4035 GND 0.006149f
C6705 VDD.n4036 GND 0.006149f
C6706 VDD.n4037 GND 0.006149f
C6707 VDD.n4038 GND 0.006149f
C6708 VDD.n4039 GND 0.006149f
C6709 VDD.n4040 GND 0.003984f
C6710 VDD.t35 GND 0.179673f
C6711 VDD.t34 GND 0.743196f
C6712 VDD.n4041 GND 0.095879f
C6713 VDD.t36 GND 0.131174f
C6714 VDD.n4042 GND 0.098395f
C6715 VDD.n4043 GND 0.006149f
C6716 VDD.n4044 GND 0.006149f
C6717 VDD.n4045 GND 0.006149f
C6718 VDD.n4046 GND 0.006149f
C6719 VDD.n4047 GND 0.006149f
C6720 VDD.n4048 GND 0.006149f
C6721 VDD.n4049 GND 0.006149f
C6722 VDD.n4050 GND 0.006149f
C6723 VDD.n4051 GND 0.006149f
C6724 VDD.n4052 GND 0.006149f
C6725 VDD.n4053 GND 0.006149f
C6726 VDD.n4054 GND 0.006149f
C6727 VDD.n4055 GND 0.006149f
C6728 VDD.n4056 GND 0.006149f
C6729 VDD.n4057 GND 0.006149f
C6730 VDD.n4058 GND 0.006149f
C6731 VDD.t38 GND 0.179673f
C6732 VDD.t37 GND 0.743196f
C6733 VDD.n4059 GND 0.095879f
C6734 VDD.t39 GND 0.131174f
C6735 VDD.n4060 GND 0.098395f
C6736 VDD.n4061 GND 0.006806f
C6737 VDD.n4062 GND 0.006149f
C6738 VDD.n4063 GND 0.006149f
C6739 VDD.n4064 GND 0.006149f
C6740 VDD.n4065 GND 0.006149f
C6741 VDD.n4066 GND 0.006149f
C6742 VDD.n4067 GND 0.006149f
C6743 VDD.n4068 GND 0.006149f
C6744 VDD.n4069 GND 0.006149f
C6745 VDD.n4070 GND 0.006149f
C6746 VDD.n4071 GND 0.006149f
C6747 VDD.n4072 GND 0.006149f
C6748 VDD.n4073 GND 0.006149f
C6749 VDD.n4074 GND 0.006149f
C6750 VDD.n4075 GND 0.006149f
C6751 VDD.n4076 GND 0.006149f
C6752 VDD.n4077 GND 0.006149f
C6753 VDD.n4078 GND 0.01414f
C6754 VDD.n4079 GND 0.002796f
C6755 VDD.t23 GND 0.179673f
C6756 VDD.t21 GND 0.743196f
C6757 VDD.n4080 GND 0.095879f
C6758 VDD.t24 GND 0.131174f
C6759 VDD.n4081 GND 0.098395f
C6760 VDD.n4082 GND 0.006149f
C6761 VDD.n4083 GND 0.004949f
C6762 VDD.n4084 GND 0.006149f
C6763 VDD.n4085 GND 0.004949f
C6764 VDD.n4086 GND 0.006149f
C6765 VDD.n4087 GND 0.004949f
C6766 VDD.n4088 GND 0.006149f
C6767 VDD.n4089 GND 0.004949f
C6768 VDD.n4090 GND 0.006149f
C6769 VDD.n4091 GND 0.006149f
C6770 VDD.n4092 GND 0.004949f
C6771 VDD.n4093 GND 0.004949f
C6772 VDD.n4094 GND 0.006149f
C6773 VDD.n4095 GND 0.006149f
C6774 VDD.n4096 GND 0.006149f
C6775 VDD.n4097 GND 0.006149f
C6776 VDD.n4098 GND 0.004949f
C6777 VDD.n4099 GND 0.004949f
C6778 VDD.n4100 GND 0.004949f
C6779 VDD.n4101 GND 0.006149f
C6780 VDD.n4102 GND 0.006149f
C6781 VDD.n4103 GND 0.006149f
C6782 VDD.n4104 GND 0.006149f
C6783 VDD.n4105 GND 0.004949f
C6784 VDD.n4106 GND 0.004949f
C6785 VDD.n4107 GND 0.004949f
C6786 VDD.n4108 GND 0.006149f
C6787 VDD.n4109 GND 0.006149f
C6788 VDD.n4110 GND 0.006149f
C6789 VDD.n4111 GND 0.006149f
C6790 VDD.n4112 GND 0.004949f
C6791 VDD.n4113 GND 0.004949f
C6792 VDD.n4114 GND 0.004949f
C6793 VDD.n4115 GND 0.006149f
C6794 VDD.n4116 GND 0.006149f
C6795 VDD.n4117 GND 0.006149f
C6796 VDD.n4118 GND 0.006149f
C6797 VDD.n4119 GND 0.004949f
C6798 VDD.n4120 GND 0.004949f
C6799 VDD.n4121 GND 0.004108f
C6800 VDD.n4122 GND 0.013778f
C6801 VDD.n4123 GND 0.01414f
C6802 VDD.n4124 GND 0.006149f
C6803 VDD.n4125 GND 0.00928f
C6804 VDD.n4126 GND 0.006149f
C6805 VDD.n4127 GND 0.006149f
C6806 VDD.n4128 GND 0.004628f
C6807 VDD.n4129 GND 0.004949f
C6808 VDD.n4130 GND 0.006149f
C6809 VDD.n4131 GND 0.006149f
C6810 VDD.n4132 GND 0.004949f
C6811 VDD.n4133 GND 0.004949f
C6812 VDD.n4134 GND 0.006149f
C6813 VDD.n4135 GND 0.006149f
C6814 VDD.n4136 GND 0.004949f
C6815 VDD.n4137 GND 0.004949f
C6816 VDD.n4138 GND 0.006149f
C6817 VDD.n4139 GND 0.006149f
C6818 VDD.n4140 GND 0.004949f
C6819 VDD.n4141 GND 0.004949f
C6820 VDD.n4142 GND 0.006149f
C6821 VDD.n4143 GND 0.006149f
C6822 VDD.n4144 GND 0.004949f
C6823 VDD.n4145 GND 0.004949f
C6824 VDD.n4146 GND 0.006149f
C6825 VDD.n4147 GND 0.006149f
C6826 VDD.n4148 GND 0.004949f
C6827 VDD.n4149 GND 0.004949f
C6828 VDD.n4150 GND 0.006149f
C6829 VDD.n4151 GND 0.006149f
C6830 VDD.n4152 GND 0.004949f
C6831 VDD.n4153 GND 0.004949f
C6832 VDD.n4154 GND 0.006149f
C6833 VDD.n4155 GND 0.006149f
C6834 VDD.n4156 GND 0.004949f
C6835 VDD.n4157 GND 0.002574f
C6836 VDD.n4158 GND 0.006149f
C6837 VDD.n4159 GND 0.006149f
C6838 VDD.n4160 GND 0.003217f
C6839 VDD.n4161 GND 0.004949f
C6840 VDD.n4162 GND 0.006149f
C6841 VDD.n4163 GND 0.006149f
C6842 VDD.n4164 GND 0.004949f
C6843 VDD.n4165 GND 0.004949f
C6844 VDD.n4166 GND 0.006149f
C6845 VDD.n4167 GND 0.006149f
C6846 VDD.n4168 GND 0.004949f
C6847 VDD.n4169 GND 0.004949f
C6848 VDD.n4170 GND 0.006149f
C6849 VDD.n4171 GND 0.006149f
C6850 VDD.n4172 GND 0.004949f
C6851 VDD.n4173 GND 0.004949f
C6852 VDD.n4174 GND 0.006149f
C6853 VDD.n4175 GND 0.006149f
C6854 VDD.n4176 GND 0.004949f
C6855 VDD.n4177 GND 0.004949f
C6856 VDD.n4178 GND 0.006149f
C6857 VDD.n4179 GND 0.006149f
C6858 VDD.n4180 GND 0.004949f
C6859 VDD.n4181 GND 0.004949f
C6860 VDD.n4182 GND 0.006149f
C6861 VDD.n4183 GND 0.006149f
C6862 VDD.n4184 GND 0.004949f
C6863 VDD.n4185 GND 0.004949f
C6864 VDD.n4186 GND 0.006149f
C6865 VDD.n4187 GND 0.006149f
C6866 VDD.n4188 GND 0.004949f
C6867 VDD.n4189 GND 0.006149f
C6868 VDD.n4190 GND 0.006149f
C6869 VDD.n4191 GND 0.006149f
C6870 VDD.n4192 GND 0.00928f
C6871 VDD.n4193 GND 0.004281f
C6872 VDD.n4194 GND 0.006149f
C6873 VDD.n4195 GND 0.006149f
C6874 VDD.n4196 GND 0.004949f
C6875 VDD.n4197 GND 0.004949f
C6876 VDD.n4198 GND 0.006149f
C6877 VDD.n4199 GND 0.006149f
C6878 VDD.n4200 GND 0.004949f
C6879 VDD.n4201 GND 0.004949f
C6880 VDD.n4202 GND 0.006149f
C6881 VDD.n4203 GND 0.006149f
C6882 VDD.n4204 GND 0.004949f
C6883 VDD.n4205 GND 0.004949f
C6884 VDD.n4206 GND 0.006149f
C6885 VDD.n4207 GND 0.006149f
C6886 VDD.n4208 GND 0.004949f
C6887 VDD.n4209 GND 0.004949f
C6888 VDD.n4210 GND 0.006149f
C6889 VDD.n4211 GND 0.006149f
C6890 VDD.n4212 GND 0.004949f
C6891 VDD.n4213 GND 0.006149f
C6892 VDD.n4214 GND 0.006149f
C6893 VDD.n4215 GND 0.004949f
C6894 VDD.n4216 GND 0.006149f
C6895 VDD.n4217 GND 0.006149f
C6896 VDD.n4218 GND 0.006149f
C6897 VDD.n4219 GND 0.004949f
C6898 VDD.n4220 GND 0.004108f
C6899 VDD.n4221 GND 0.01414f
C6900 VDD.n4222 GND 1.13918f
C6901 VDD.n4223 GND 0.695475f
C6902 VDD.n4224 GND 0.498548f
C6903 VDD.n4225 GND 0.006149f
C6904 VDD.n4226 GND 0.004949f
C6905 VDD.n4227 GND 0.004949f
C6906 VDD.n4228 GND 0.004949f
C6907 VDD.n4229 GND 0.006149f
C6908 VDD.n4230 GND 0.498548f
C6909 VDD.n4231 GND 0.498548f
C6910 VDD.n4232 GND 0.498548f
C6911 VDD.n4233 GND 0.006149f
C6912 VDD.n4234 GND 0.004949f
C6913 VDD.n4235 GND 0.004949f
C6914 VDD.n4236 GND 0.004949f
C6915 VDD.n4237 GND 0.006149f
C6916 VDD.n4238 GND 0.40881f
C6917 VDD.n4239 GND 0.498548f
C6918 VDD.n4240 GND 0.498548f
C6919 VDD.n4241 GND 0.006149f
C6920 VDD.n4242 GND 0.004949f
C6921 VDD.n4243 GND 0.004949f
C6922 VDD.n4244 GND 0.004949f
C6923 VDD.n4245 GND 0.006149f
C6924 VDD.n4246 GND 0.498548f
C6925 VDD.n4247 GND 0.498548f
C6926 VDD.n4248 GND 0.498548f
C6927 VDD.n4249 GND 0.006149f
C6928 VDD.n4250 GND 0.004949f
C6929 VDD.n4251 GND 0.004949f
C6930 VDD.n4252 GND 0.004949f
C6931 VDD.n4253 GND 0.006149f
C6932 VDD.n4254 GND 0.498548f
C6933 VDD.n4255 GND 0.498548f
C6934 VDD.n4256 GND 0.498548f
C6935 VDD.n4257 GND 0.006149f
C6936 VDD.n4258 GND 0.004949f
C6937 VDD.n4259 GND 0.004949f
C6938 VDD.n4260 GND 0.004949f
C6939 VDD.n4261 GND 0.006149f
C6940 VDD.n4262 GND 0.498548f
C6941 VDD.n4263 GND 0.006149f
C6942 VDD.n4264 GND 0.004949f
C6943 VDD.n4265 GND 0.004949f
C6944 VDD.n4266 GND 0.004949f
C6945 VDD.n4267 GND 0.006149f
C6946 VDD.t99 GND 0.498548f
C6947 VDD.n4268 GND 0.006149f
C6948 VDD.n4269 GND 0.004949f
C6949 VDD.n4270 GND 0.004949f
C6950 VDD.n4271 GND 0.004949f
C6951 VDD.n4272 GND 0.006149f
C6952 VDD.n4273 GND 0.498548f
C6953 VDD.n4274 GND 0.498548f
C6954 VDD.n4275 GND 0.498548f
C6955 VDD.n4276 GND 0.006149f
C6956 VDD.n4277 GND 0.004949f
C6957 VDD.n4278 GND 0.004949f
C6958 VDD.n4279 GND 0.004949f
C6959 VDD.n4280 GND 0.006149f
C6960 VDD.n4281 GND 0.498548f
C6961 VDD.n4282 GND 0.498548f
C6962 VDD.n4283 GND 0.498548f
C6963 VDD.n4284 GND 0.006149f
C6964 VDD.n4285 GND 0.004949f
C6965 VDD.n4286 GND 0.004949f
C6966 VDD.n4287 GND 0.004949f
C6967 VDD.n4288 GND 0.006149f
C6968 VDD.n4289 GND 0.498548f
C6969 VDD.n4290 GND 0.448694f
C6970 VDD.t70 GND 0.249274f
C6971 VDD.n4291 GND 0.299129f
C6972 VDD.n4292 GND 0.006149f
C6973 VDD.n4293 GND 0.004949f
C6974 VDD.n4294 GND 0.004949f
C6975 VDD.n4295 GND 0.004949f
C6976 VDD.n4296 GND 0.006149f
C6977 VDD.n4297 GND 0.498548f
C6978 VDD.n4298 GND 0.498548f
C6979 VDD.n4299 GND 0.498548f
C6980 VDD.n4300 GND 0.006149f
C6981 VDD.n4301 GND 0.004949f
C6982 VDD.n4302 GND 0.004949f
C6983 VDD.n4303 GND 0.004949f
C6984 VDD.n4304 GND 0.006149f
C6985 VDD.n4305 GND 0.498548f
C6986 VDD.n4306 GND 0.498548f
C6987 VDD.n4307 GND 0.498548f
C6988 VDD.n4308 GND 0.006149f
C6989 VDD.n4309 GND 0.004949f
C6990 VDD.n4310 GND 0.004949f
C6991 VDD.n4311 GND 0.004949f
C6992 VDD.n4312 GND 0.006149f
C6993 VDD.n4313 GND 0.498548f
C6994 VDD.n4314 GND 0.398839f
C6995 VDD.t83 GND 0.249274f
C6996 VDD.n4315 GND 0.348984f
C6997 VDD.n4316 GND 0.006149f
C6998 VDD.n4317 GND 0.004949f
C6999 VDD.n4318 GND 0.004949f
C7000 VDD.n4319 GND 0.004949f
C7001 VDD.n4320 GND 0.006149f
C7002 VDD.n4321 GND 0.498548f
C7003 VDD.n4322 GND 0.498548f
C7004 VDD.n4323 GND 0.498548f
C7005 VDD.n4324 GND 0.006149f
C7006 VDD.n4325 GND 0.004949f
C7007 VDD.n4326 GND 0.004949f
C7008 VDD.n4327 GND 0.004726f
C7009 VDD.n4328 GND 0.330844f
C7010 VDD.n4329 GND 2.94455f
C7011 a_n18640_8567.n0 GND 0.537469f
C7012 a_n18640_8567.n1 GND 0.616917f
C7013 a_n18640_8567.n2 GND 0.537469f
C7014 a_n18640_8567.n3 GND 0.616917f
C7015 a_n18640_8567.n4 GND 0.60089f
C7016 a_n18640_8567.n5 GND 0.616917f
C7017 a_n18640_8567.n6 GND 0.226382f
C7018 a_n18640_8567.n7 GND 0.226382f
C7019 a_n18640_8567.n8 GND 0.253594f
C7020 a_n18640_8567.n9 GND 0.226382f
C7021 a_n18640_8567.n10 GND 0.218418f
C7022 a_n18640_8567.n11 GND 0.226382f
C7023 a_n18640_8567.n12 GND 0.175419f
C7024 a_n18640_8567.n13 GND 0.226382f
C7025 a_n18640_8567.n14 GND 0.23713f
C7026 a_n18640_8567.n15 GND 0.406708f
C7027 a_n18640_8567.n16 GND 0.218661f
C7028 a_n18640_8567.n17 GND 0.226382f
C7029 a_n18640_8567.n18 GND 0.226382f
C7030 a_n18640_8567.n19 GND 0.253594f
C7031 a_n18640_8567.n20 GND 0.226382f
C7032 a_n18640_8567.n21 GND 0.218418f
C7033 a_n18640_8567.n22 GND 0.226382f
C7034 a_n18640_8567.n23 GND 0.175419f
C7035 a_n18640_8567.n24 GND 0.226382f
C7036 a_n18640_8567.n25 GND 0.23713f
C7037 a_n18640_8567.n26 GND 0.406708f
C7038 a_n18640_8567.n27 GND 0.218661f
C7039 a_n18640_8567.n28 GND 0.226382f
C7040 a_n18640_8567.n29 GND 0.226382f
C7041 a_n18640_8567.n30 GND 0.253594f
C7042 a_n18640_8567.n31 GND 0.226382f
C7043 a_n18640_8567.n32 GND 0.218418f
C7044 a_n18640_8567.n33 GND 0.226382f
C7045 a_n18640_8567.n34 GND 0.175419f
C7046 a_n18640_8567.n35 GND 0.226382f
C7047 a_n18640_8567.n36 GND 0.23713f
C7048 a_n18640_8567.n37 GND 0.406708f
C7049 a_n18640_8567.n38 GND 0.218661f
C7050 a_n18640_8567.n39 GND 0.491601f
C7051 a_n18640_8567.n40 GND 0.218418f
C7052 a_n18640_8567.n41 GND 0.226382f
C7053 a_n18640_8567.n42 GND 0.175419f
C7054 a_n18640_8567.n43 GND 0.226382f
C7055 a_n18640_8567.n44 GND 0.23713f
C7056 a_n18640_8567.n45 GND 0.226382f
C7057 a_n18640_8567.n46 GND 0.218661f
C7058 a_n18640_8567.n47 GND 0.226382f
C7059 a_n18640_8567.n48 GND 0.491601f
C7060 a_n18640_8567.n49 GND 0.218418f
C7061 a_n18640_8567.n50 GND 0.226382f
C7062 a_n18640_8567.n51 GND 0.175419f
C7063 a_n18640_8567.n52 GND 0.226382f
C7064 a_n18640_8567.n53 GND 0.23713f
C7065 a_n18640_8567.n54 GND 0.226382f
C7066 a_n18640_8567.n55 GND 0.218661f
C7067 a_n18640_8567.n56 GND 0.226382f
C7068 a_n18640_8567.n57 GND 0.491601f
C7069 a_n18640_8567.n58 GND 0.218418f
C7070 a_n18640_8567.n59 GND 0.226382f
C7071 a_n18640_8567.n60 GND 0.175419f
C7072 a_n18640_8567.n61 GND 0.226382f
C7073 a_n18640_8567.n62 GND 0.23713f
C7074 a_n18640_8567.n63 GND 0.226382f
C7075 a_n18640_8567.n64 GND 0.218661f
C7076 a_n18640_8567.n65 GND 0.226382f
C7077 a_n18640_8567.n66 GND 0.395981f
C7078 a_n18640_8567.n67 GND 0.644823f
C7079 a_n18640_8567.n68 GND 0.395981f
C7080 a_n18640_8567.n69 GND 0.644823f
C7081 a_n18640_8567.n70 GND 0.459401f
C7082 a_n18640_8567.n71 GND 0.644823f
C7083 a_n18640_8567.n72 GND 0.170044f
C7084 a_n18640_8567.n73 GND 0.178108f
C7085 a_n18640_8567.n74 GND 0.165381f
C7086 a_n18640_8567.n75 GND 0.170044f
C7087 a_n18640_8567.n76 GND 0.178108f
C7088 a_n18640_8567.n77 GND 0.165381f
C7089 a_n18640_8567.n78 GND 0.170044f
C7090 a_n18640_8567.n79 GND 0.178108f
C7091 a_n18640_8567.n80 GND 0.165381f
C7092 a_n18640_8567.n81 GND 0.178108f
C7093 a_n18640_8567.n82 GND 0.165381f
C7094 a_n18640_8567.n83 GND 0.178108f
C7095 a_n18640_8567.n84 GND 0.165381f
C7096 a_n18640_8567.n85 GND 0.178108f
C7097 a_n18640_8567.n86 GND 0.165381f
C7098 a_n18640_8567.n87 GND 0.123489f
C7099 a_n18640_8567.n88 GND 0.123489f
C7100 a_n18640_8567.n89 GND 0.123489f
C7101 a_n18640_8567.t17 GND 0.089851f
C7102 a_n18640_8567.t14 GND 0.089851f
C7103 a_n18640_8567.t13 GND 0.089851f
C7104 a_n18640_8567.n90 GND 0.511603f
C7105 a_n18640_8567.t12 GND 0.089851f
C7106 a_n18640_8567.t18 GND 0.089851f
C7107 a_n18640_8567.n91 GND 0.496767f
C7108 a_n18640_8567.n92 GND 4.47007f
C7109 a_n18640_8567.t9 GND 0.09491f
C7110 a_n18640_8567.t11 GND 0.09491f
C7111 a_n18640_8567.n93 GND 0.706068f
C7112 a_n18640_8567.t4 GND 0.09491f
C7113 a_n18640_8567.t0 GND 0.09491f
C7114 a_n18640_8567.n94 GND 0.673066f
C7115 a_n18640_8567.t8 GND 0.09491f
C7116 a_n18640_8567.t1 GND 0.09491f
C7117 a_n18640_8567.n95 GND 0.706067f
C7118 a_n18640_8567.t6 GND 0.09491f
C7119 a_n18640_8567.t7 GND 0.09491f
C7120 a_n18640_8567.n96 GND 0.673065f
C7121 a_n18640_8567.t10 GND 0.09491f
C7122 a_n18640_8567.t2 GND 0.09491f
C7123 a_n18640_8567.n97 GND 0.706067f
C7124 a_n18640_8567.n98 GND 7.79829f
C7125 a_n18640_8567.t3 GND 0.09491f
C7126 a_n18640_8567.t5 GND 0.09491f
C7127 a_n18640_8567.n99 GND 0.673066f
C7128 a_n18640_8567.n100 GND 4.8645f
C7129 a_n18640_8567.n101 GND 2.72007f
C7130 a_n18640_8567.t42 GND 2.41267f
C7131 a_n18640_8567.t32 GND 1.88106f
C7132 a_n18640_8567.n102 GND 0.802165f
C7133 a_n18640_8567.t46 GND 1.88106f
C7134 a_n18640_8567.n103 GND 0.905314f
C7135 a_n18640_8567.t40 GND 2.45823f
C7136 a_n18640_8567.n104 GND 1.01156f
C7137 a_n18640_8567.t21 GND 1.88106f
C7138 a_n18640_8567.n105 GND 0.898629f
C7139 a_n18640_8567.t51 GND 1.88106f
C7140 a_n18640_8567.n106 GND 0.800712f
C7141 a_n18640_8567.t43 GND 2.41267f
C7142 a_n18640_8567.t30 GND 1.88106f
C7143 a_n18640_8567.n107 GND 0.802165f
C7144 a_n18640_8567.t44 GND 1.88106f
C7145 a_n18640_8567.n108 GND 0.905314f
C7146 a_n18640_8567.t39 GND 2.45823f
C7147 a_n18640_8567.n109 GND 1.01156f
C7148 a_n18640_8567.t20 GND 1.88106f
C7149 a_n18640_8567.n110 GND 0.898629f
C7150 a_n18640_8567.t52 GND 1.88106f
C7151 a_n18640_8567.n111 GND 0.800712f
C7152 a_n18640_8567.n112 GND 0.421957f
C7153 a_n18640_8567.t50 GND 2.41267f
C7154 a_n18640_8567.t27 GND 1.88106f
C7155 a_n18640_8567.n113 GND 0.802165f
C7156 a_n18640_8567.t28 GND 1.88106f
C7157 a_n18640_8567.n114 GND 0.905314f
C7158 a_n18640_8567.t41 GND 2.45823f
C7159 a_n18640_8567.n115 GND 1.01156f
C7160 a_n18640_8567.t26 GND 1.88106f
C7161 a_n18640_8567.n116 GND 0.898629f
C7162 a_n18640_8567.t53 GND 1.88106f
C7163 a_n18640_8567.n117 GND 0.800712f
C7164 a_n18640_8567.n118 GND 2.30302f
C7165 a_n18640_8567.t25 GND 2.23087f
C7166 a_n18640_8567.t38 GND 1.88106f
C7167 a_n18640_8567.n119 GND 0.788108f
C7168 a_n18640_8567.t31 GND 1.88106f
C7169 a_n18640_8567.n120 GND 0.802165f
C7170 a_n18640_8567.t45 GND 1.88106f
C7171 a_n18640_8567.n121 GND 0.898629f
C7172 a_n18640_8567.t22 GND 2.45823f
C7173 a_n18640_8567.t54 GND 1.88106f
C7174 a_n18640_8567.n122 GND 0.864778f
C7175 a_n18640_8567.n123 GND 1.01157f
C7176 a_n18640_8567.t24 GND 2.23087f
C7177 a_n18640_8567.t37 GND 1.88106f
C7178 a_n18640_8567.n124 GND 0.788108f
C7179 a_n18640_8567.t29 GND 1.88106f
C7180 a_n18640_8567.n125 GND 0.802165f
C7181 a_n18640_8567.t47 GND 1.88106f
C7182 a_n18640_8567.n126 GND 0.898629f
C7183 a_n18640_8567.t23 GND 2.45823f
C7184 a_n18640_8567.t55 GND 1.88106f
C7185 a_n18640_8567.n127 GND 0.864778f
C7186 a_n18640_8567.n128 GND 1.01157f
C7187 a_n18640_8567.n129 GND 0.421957f
C7188 a_n18640_8567.t48 GND 2.23087f
C7189 a_n18640_8567.t49 GND 1.88106f
C7190 a_n18640_8567.n130 GND 0.788108f
C7191 a_n18640_8567.t33 GND 1.88106f
C7192 a_n18640_8567.n131 GND 0.802165f
C7193 a_n18640_8567.t34 GND 1.88106f
C7194 a_n18640_8567.n132 GND 0.898629f
C7195 a_n18640_8567.t36 GND 2.45823f
C7196 a_n18640_8567.t35 GND 1.88106f
C7197 a_n18640_8567.n133 GND 0.864778f
C7198 a_n18640_8567.n134 GND 1.01157f
C7199 a_n18640_8567.n135 GND 1.05436f
C7200 a_n18640_8567.n136 GND 16.2107f
C7201 a_n18640_8567.n137 GND 2.42898f
C7202 a_n18640_8567.n138 GND 8.8814f
C7203 a_n18640_8567.t15 GND 0.089851f
C7204 a_n18640_8567.t16 GND 0.089851f
C7205 a_n18640_8567.n139 GND 0.511601f
C7206 a_n18640_8567.n140 GND 5.61685f
C7207 a_n18640_8567.n141 GND 0.496767f
C7208 a_n18640_8567.t19 GND 0.089851f
C7209 a_n5326_8245.n0 GND 4.969f
C7210 a_n5326_8245.n1 GND 5.41733f
C7211 a_n5326_8245.n2 GND 3.67239f
C7212 a_n5326_8245.n3 GND 4.72852f
C7213 a_n5326_8245.t0 GND 0.171142p
C7214 a_n5326_8245.t10 GND 0.483862f
C7215 a_n5326_8245.t15 GND 0.077269f
C7216 a_n5326_8245.t6 GND 0.077269f
C7217 a_n5326_8245.n4 GND 0.35788f
C7218 a_n5326_8245.t13 GND 0.473922f
C7219 a_n5326_8245.t5 GND 0.483865f
C7220 a_n5326_8245.t7 GND 0.077269f
C7221 a_n5326_8245.t16 GND 0.077269f
C7222 a_n5326_8245.n5 GND 0.35788f
C7223 a_n5326_8245.t9 GND 0.473922f
C7224 a_n5326_8245.t8 GND 0.473922f
C7225 a_n5326_8245.t2 GND 0.077269f
C7226 a_n5326_8245.t11 GND 0.077269f
C7227 a_n5326_8245.n6 GND 0.35788f
C7228 a_n5326_8245.t3 GND 0.483865f
C7229 a_n5326_8245.t12 GND 0.077269f
C7230 a_n5326_8245.t14 GND 0.077269f
C7231 a_n5326_8245.n7 GND 0.35788f
C7232 a_n5326_8245.t4 GND 0.473922f
C7233 a_n5326_8245.t1 GND 0.473922f
C7234 a_n7837_10186.n0 GND 4.46585f
C7235 a_n7837_10186.n1 GND 0.648796f
C7236 a_n7837_10186.n2 GND 3.54323f
C7237 a_n7837_10186.n3 GND 1.05432f
C7238 a_n7837_10186.n4 GND 3.55849f
C7239 a_n7837_10186.n5 GND 1.05432f
C7240 a_n7837_10186.n6 GND 3.42272f
C7241 a_n7837_10186.n7 GND 1.05432f
C7242 a_n7837_10186.n8 GND 10.9807f
C7243 a_n7837_10186.n9 GND 1.05626f
C7244 a_n7837_10186.n10 GND 1.05685f
C7245 a_n7837_10186.n11 GND 1.91784f
C7246 a_n7837_10186.n12 GND 1.05897f
C7247 a_n7837_10186.n13 GND 1.05635f
C7248 a_n7837_10186.n14 GND 0.646788f
C7249 a_n7837_10186.n15 GND 9.99096f
C7250 a_n7837_10186.n16 GND 1.72118f
C7251 a_n7837_10186.n17 GND 4.93917f
C7252 a_n7837_10186.n18 GND 4.80522f
C7253 a_n7837_10186.t21 GND 2.03429f
C7254 a_n7837_10186.t19 GND 1.61672f
C7255 a_n7837_10186.t2 GND 0.108277f
C7256 a_n7837_10186.t1 GND 0.108277f
C7257 a_n7837_10186.n19 GND 0.805502f
C7258 a_n7837_10186.t10 GND 0.108277f
C7259 a_n7837_10186.t3 GND 0.108277f
C7260 a_n7837_10186.n20 GND 0.767852f
C7261 a_n7837_10186.t27 GND 0.108277f
C7262 a_n7837_10186.t0 GND 0.108277f
C7263 a_n7837_10186.n21 GND 0.805502f
C7264 a_n7837_10186.n22 GND 8.876571f
C7265 a_n7837_10186.t5 GND 0.108277f
C7266 a_n7837_10186.t8 GND 0.108277f
C7267 a_n7837_10186.n23 GND 0.767854f
C7268 a_n7837_10186.t6 GND 0.108277f
C7269 a_n7837_10186.t7 GND 0.108277f
C7270 a_n7837_10186.n24 GND 0.767854f
C7271 a_n7837_10186.t9 GND 0.108277f
C7272 a_n7837_10186.t4 GND 0.108277f
C7273 a_n7837_10186.n25 GND 0.805503f
C7274 a_n7837_10186.t13 GND 2.01747f
C7275 a_n7837_10186.t11 GND 2.03429f
C7276 a_n7837_10186.t40 GND 2.03429f
C7277 a_n7837_10186.t47 GND 2.01981f
C7278 a_n7837_10186.t48 GND 2.04622f
C7279 a_n7837_10186.t35 GND 2.03428f
C7280 a_n7837_10186.t18 GND 0.64189f
C7281 a_n7837_10186.t16 GND 0.102505f
C7282 a_n7837_10186.t24 GND 0.102505f
C7283 a_n7837_10186.n26 GND 0.474759f
C7284 a_n7837_10186.t26 GND 0.628695f
C7285 a_n7837_10186.t25 GND 2.03428f
C7286 a_n7837_10186.t23 GND 2.04622f
C7287 a_n7837_10186.t15 GND 2.01981f
C7288 a_n7837_10186.t17 GND 2.03429f
C7289 a_n7837_10186.t38 GND 2.03428f
C7290 a_n7837_10186.t39 GND 2.04622f
C7291 a_n7837_10186.t28 GND 2.01981f
C7292 a_n7837_10186.t37 GND 2.03429f
C7293 a_n7837_10186.t36 GND 2.03428f
C7294 a_n7837_10186.t45 GND 2.01976f
C7295 a_n7837_10186.t33 GND 2.04424f
C7296 a_n7837_10186.t51 GND 2.03429f
C7297 a_n7837_10186.t50 GND 2.03428f
C7298 a_n7837_10186.t32 GND 2.04401f
C7299 a_n7837_10186.t49 GND 2.01948f
C7300 a_n7837_10186.t43 GND 2.03429f
C7301 a_n7837_10186.t31 GND 2.03428f
C7302 a_n7837_10186.t44 GND 2.02079f
C7303 a_n7837_10186.t29 GND 2.04059f
C7304 a_n7837_10186.t34 GND 2.03429f
C7305 a_n7837_10186.t42 GND 2.03428f
C7306 a_n7837_10186.t30 GND 2.04498f
C7307 a_n7837_10186.t41 GND 2.01911f
C7308 a_n7837_10186.t46 GND 2.03429f
C7309 a_n7837_10186.n27 GND 0.837367f
C7310 a_n7837_10186.t22 GND 0.628699f
C7311 a_n7837_10186.t20 GND 0.102505f
C7312 a_n7837_10186.t14 GND 0.102505f
C7313 a_n7837_10186.n28 GND 0.474759f
C7314 a_n7837_10186.t12 GND 0.64189f
.ends

