* NGSPICE file created from diff_pair_sample_1527.ext - technology: sky130A

.subckt diff_pair_sample_1527 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t19 B.t0 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X1 VDD1.t9 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X2 VDD1.t8 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=2.36445 ps=14.66 w=14.33 l=3.94
X3 VTAIL.t18 VN.t1 VDD2.t8 B.t9 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X4 VTAIL.t17 VN.t2 VDD2.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X5 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=0 ps=0 w=14.33 l=3.94
X6 VDD2.t6 VN.t3 VTAIL.t16 B.t3 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X7 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=0 ps=0 w=14.33 l=3.94
X8 VDD1.t7 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=2.36445 ps=14.66 w=14.33 l=3.94
X9 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=0 ps=0 w=14.33 l=3.94
X10 VDD1.t6 VP.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X11 VDD2.t5 VN.t4 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=2.36445 ps=14.66 w=14.33 l=3.94
X12 VDD2.t4 VN.t5 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=5.5887 ps=29.44 w=14.33 l=3.94
X13 VTAIL.t9 VP.t4 VDD1.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X14 VTAIL.t15 VN.t6 VDD2.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X15 VTAIL.t10 VN.t7 VDD2.t2 B.t7 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X16 VTAIL.t7 VP.t5 VDD1.t4 B.t7 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X17 VTAIL.t8 VP.t6 VDD1.t3 B.t8 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
X18 VDD1.t2 VP.t7 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=5.5887 ps=29.44 w=14.33 l=3.94
X19 VDD2.t1 VN.t8 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=2.36445 ps=14.66 w=14.33 l=3.94
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.5887 pd=29.44 as=0 ps=0 w=14.33 l=3.94
X21 VDD2.t0 VN.t9 VTAIL.t12 B.t6 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=5.5887 ps=29.44 w=14.33 l=3.94
X22 VDD1.t1 VP.t8 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=5.5887 ps=29.44 w=14.33 l=3.94
X23 VTAIL.t4 VP.t9 VDD1.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=2.36445 pd=14.66 as=2.36445 ps=14.66 w=14.33 l=3.94
R0 VN.n112 VN.n111 161.3
R1 VN.n110 VN.n58 161.3
R2 VN.n109 VN.n108 161.3
R3 VN.n107 VN.n59 161.3
R4 VN.n106 VN.n105 161.3
R5 VN.n104 VN.n60 161.3
R6 VN.n103 VN.n102 161.3
R7 VN.n101 VN.n61 161.3
R8 VN.n100 VN.n99 161.3
R9 VN.n97 VN.n62 161.3
R10 VN.n96 VN.n95 161.3
R11 VN.n94 VN.n63 161.3
R12 VN.n93 VN.n92 161.3
R13 VN.n91 VN.n64 161.3
R14 VN.n90 VN.n89 161.3
R15 VN.n88 VN.n65 161.3
R16 VN.n87 VN.n86 161.3
R17 VN.n85 VN.n66 161.3
R18 VN.n84 VN.n83 161.3
R19 VN.n82 VN.n67 161.3
R20 VN.n81 VN.n80 161.3
R21 VN.n79 VN.n68 161.3
R22 VN.n78 VN.n77 161.3
R23 VN.n76 VN.n69 161.3
R24 VN.n75 VN.n74 161.3
R25 VN.n73 VN.n70 161.3
R26 VN.n55 VN.n54 161.3
R27 VN.n53 VN.n1 161.3
R28 VN.n52 VN.n51 161.3
R29 VN.n50 VN.n2 161.3
R30 VN.n49 VN.n48 161.3
R31 VN.n47 VN.n3 161.3
R32 VN.n46 VN.n45 161.3
R33 VN.n44 VN.n4 161.3
R34 VN.n43 VN.n42 161.3
R35 VN.n40 VN.n5 161.3
R36 VN.n39 VN.n38 161.3
R37 VN.n37 VN.n6 161.3
R38 VN.n36 VN.n35 161.3
R39 VN.n34 VN.n7 161.3
R40 VN.n33 VN.n32 161.3
R41 VN.n31 VN.n8 161.3
R42 VN.n30 VN.n29 161.3
R43 VN.n28 VN.n9 161.3
R44 VN.n27 VN.n26 161.3
R45 VN.n25 VN.n10 161.3
R46 VN.n24 VN.n23 161.3
R47 VN.n22 VN.n11 161.3
R48 VN.n21 VN.n20 161.3
R49 VN.n19 VN.n12 161.3
R50 VN.n18 VN.n17 161.3
R51 VN.n16 VN.n13 161.3
R52 VN.n71 VN.t5 120.222
R53 VN.n14 VN.t4 120.222
R54 VN.n56 VN.n0 88.1101
R55 VN.n113 VN.n57 88.1101
R56 VN.n28 VN.t3 87.6535
R57 VN.n15 VN.t2 87.6535
R58 VN.n41 VN.t7 87.6535
R59 VN.n0 VN.t9 87.6535
R60 VN.n85 VN.t0 87.6535
R61 VN.n72 VN.t6 87.6535
R62 VN.n98 VN.t1 87.6535
R63 VN.n57 VN.t8 87.6535
R64 VN VN.n113 62.4033
R65 VN.n15 VN.n14 61.9406
R66 VN.n72 VN.n71 61.9406
R67 VN.n22 VN.n21 53.6055
R68 VN.n35 VN.n34 53.6055
R69 VN.n79 VN.n78 53.6055
R70 VN.n92 VN.n91 53.6055
R71 VN.n48 VN.n47 49.7204
R72 VN.n105 VN.n104 49.7204
R73 VN.n48 VN.n2 31.2664
R74 VN.n105 VN.n59 31.2664
R75 VN.n23 VN.n22 27.3813
R76 VN.n34 VN.n33 27.3813
R77 VN.n80 VN.n79 27.3813
R78 VN.n91 VN.n90 27.3813
R79 VN.n17 VN.n16 24.4675
R80 VN.n17 VN.n12 24.4675
R81 VN.n21 VN.n12 24.4675
R82 VN.n23 VN.n10 24.4675
R83 VN.n27 VN.n10 24.4675
R84 VN.n28 VN.n27 24.4675
R85 VN.n29 VN.n28 24.4675
R86 VN.n29 VN.n8 24.4675
R87 VN.n33 VN.n8 24.4675
R88 VN.n35 VN.n6 24.4675
R89 VN.n39 VN.n6 24.4675
R90 VN.n40 VN.n39 24.4675
R91 VN.n42 VN.n4 24.4675
R92 VN.n46 VN.n4 24.4675
R93 VN.n47 VN.n46 24.4675
R94 VN.n52 VN.n2 24.4675
R95 VN.n53 VN.n52 24.4675
R96 VN.n54 VN.n53 24.4675
R97 VN.n78 VN.n69 24.4675
R98 VN.n74 VN.n69 24.4675
R99 VN.n74 VN.n73 24.4675
R100 VN.n90 VN.n65 24.4675
R101 VN.n86 VN.n65 24.4675
R102 VN.n86 VN.n85 24.4675
R103 VN.n85 VN.n84 24.4675
R104 VN.n84 VN.n67 24.4675
R105 VN.n80 VN.n67 24.4675
R106 VN.n104 VN.n103 24.4675
R107 VN.n103 VN.n61 24.4675
R108 VN.n99 VN.n61 24.4675
R109 VN.n97 VN.n96 24.4675
R110 VN.n96 VN.n63 24.4675
R111 VN.n92 VN.n63 24.4675
R112 VN.n111 VN.n110 24.4675
R113 VN.n110 VN.n109 24.4675
R114 VN.n109 VN.n59 24.4675
R115 VN.n16 VN.n15 13.2127
R116 VN.n41 VN.n40 13.2127
R117 VN.n73 VN.n72 13.2127
R118 VN.n98 VN.n97 13.2127
R119 VN.n42 VN.n41 11.2553
R120 VN.n99 VN.n98 11.2553
R121 VN.n71 VN.n70 2.48786
R122 VN.n14 VN.n13 2.48786
R123 VN.n54 VN.n0 1.95786
R124 VN.n111 VN.n57 1.95786
R125 VN.n113 VN.n112 0.354971
R126 VN.n56 VN.n55 0.354971
R127 VN VN.n56 0.26696
R128 VN.n112 VN.n58 0.189894
R129 VN.n108 VN.n58 0.189894
R130 VN.n108 VN.n107 0.189894
R131 VN.n107 VN.n106 0.189894
R132 VN.n106 VN.n60 0.189894
R133 VN.n102 VN.n60 0.189894
R134 VN.n102 VN.n101 0.189894
R135 VN.n101 VN.n100 0.189894
R136 VN.n100 VN.n62 0.189894
R137 VN.n95 VN.n62 0.189894
R138 VN.n95 VN.n94 0.189894
R139 VN.n94 VN.n93 0.189894
R140 VN.n93 VN.n64 0.189894
R141 VN.n89 VN.n64 0.189894
R142 VN.n89 VN.n88 0.189894
R143 VN.n88 VN.n87 0.189894
R144 VN.n87 VN.n66 0.189894
R145 VN.n83 VN.n66 0.189894
R146 VN.n83 VN.n82 0.189894
R147 VN.n82 VN.n81 0.189894
R148 VN.n81 VN.n68 0.189894
R149 VN.n77 VN.n68 0.189894
R150 VN.n77 VN.n76 0.189894
R151 VN.n76 VN.n75 0.189894
R152 VN.n75 VN.n70 0.189894
R153 VN.n18 VN.n13 0.189894
R154 VN.n19 VN.n18 0.189894
R155 VN.n20 VN.n19 0.189894
R156 VN.n20 VN.n11 0.189894
R157 VN.n24 VN.n11 0.189894
R158 VN.n25 VN.n24 0.189894
R159 VN.n26 VN.n25 0.189894
R160 VN.n26 VN.n9 0.189894
R161 VN.n30 VN.n9 0.189894
R162 VN.n31 VN.n30 0.189894
R163 VN.n32 VN.n31 0.189894
R164 VN.n32 VN.n7 0.189894
R165 VN.n36 VN.n7 0.189894
R166 VN.n37 VN.n36 0.189894
R167 VN.n38 VN.n37 0.189894
R168 VN.n38 VN.n5 0.189894
R169 VN.n43 VN.n5 0.189894
R170 VN.n44 VN.n43 0.189894
R171 VN.n45 VN.n44 0.189894
R172 VN.n45 VN.n3 0.189894
R173 VN.n49 VN.n3 0.189894
R174 VN.n50 VN.n49 0.189894
R175 VN.n51 VN.n50 0.189894
R176 VN.n51 VN.n1 0.189894
R177 VN.n55 VN.n1 0.189894
R178 VTAIL.n11 VTAIL.t11 46.6385
R179 VTAIL.n17 VTAIL.t12 46.6384
R180 VTAIL.n2 VTAIL.t5 46.6384
R181 VTAIL.n16 VTAIL.t6 46.6384
R182 VTAIL.n15 VTAIL.n14 45.2568
R183 VTAIL.n13 VTAIL.n12 45.2568
R184 VTAIL.n10 VTAIL.n9 45.2568
R185 VTAIL.n8 VTAIL.n7 45.2568
R186 VTAIL.n19 VTAIL.n18 45.2566
R187 VTAIL.n1 VTAIL.n0 45.2566
R188 VTAIL.n4 VTAIL.n3 45.2566
R189 VTAIL.n6 VTAIL.n5 45.2566
R190 VTAIL.n8 VTAIL.n6 32.0824
R191 VTAIL.n17 VTAIL.n16 28.4014
R192 VTAIL.n10 VTAIL.n8 3.68153
R193 VTAIL.n11 VTAIL.n10 3.68153
R194 VTAIL.n15 VTAIL.n13 3.68153
R195 VTAIL.n16 VTAIL.n15 3.68153
R196 VTAIL.n6 VTAIL.n4 3.68153
R197 VTAIL.n4 VTAIL.n2 3.68153
R198 VTAIL.n19 VTAIL.n17 3.68153
R199 VTAIL VTAIL.n1 2.81947
R200 VTAIL.n13 VTAIL.n11 2.31084
R201 VTAIL.n2 VTAIL.n1 2.31084
R202 VTAIL.n18 VTAIL.t16 1.38222
R203 VTAIL.n18 VTAIL.t10 1.38222
R204 VTAIL.n0 VTAIL.t13 1.38222
R205 VTAIL.n0 VTAIL.t17 1.38222
R206 VTAIL.n3 VTAIL.t0 1.38222
R207 VTAIL.n3 VTAIL.t8 1.38222
R208 VTAIL.n5 VTAIL.t2 1.38222
R209 VTAIL.n5 VTAIL.t9 1.38222
R210 VTAIL.n14 VTAIL.t3 1.38222
R211 VTAIL.n14 VTAIL.t7 1.38222
R212 VTAIL.n12 VTAIL.t1 1.38222
R213 VTAIL.n12 VTAIL.t4 1.38222
R214 VTAIL.n9 VTAIL.t19 1.38222
R215 VTAIL.n9 VTAIL.t15 1.38222
R216 VTAIL.n7 VTAIL.t14 1.38222
R217 VTAIL.n7 VTAIL.t18 1.38222
R218 VTAIL VTAIL.n19 0.862569
R219 VDD2.n1 VDD2.t5 66.9982
R220 VDD2.n3 VDD2.n2 64.6408
R221 VDD2 VDD2.n7 64.638
R222 VDD2.n4 VDD2.t1 63.3172
R223 VDD2.n6 VDD2.n5 61.9356
R224 VDD2.n1 VDD2.n0 61.9353
R225 VDD2.n4 VDD2.n3 53.5537
R226 VDD2.n6 VDD2.n4 3.68153
R227 VDD2.n7 VDD2.t3 1.38222
R228 VDD2.n7 VDD2.t4 1.38222
R229 VDD2.n5 VDD2.t8 1.38222
R230 VDD2.n5 VDD2.t9 1.38222
R231 VDD2.n2 VDD2.t2 1.38222
R232 VDD2.n2 VDD2.t0 1.38222
R233 VDD2.n0 VDD2.t7 1.38222
R234 VDD2.n0 VDD2.t6 1.38222
R235 VDD2 VDD2.n6 0.978948
R236 VDD2.n3 VDD2.n1 0.865413
R237 B.n1207 B.n1206 585
R238 B.n416 B.n204 585
R239 B.n415 B.n414 585
R240 B.n413 B.n412 585
R241 B.n411 B.n410 585
R242 B.n409 B.n408 585
R243 B.n407 B.n406 585
R244 B.n405 B.n404 585
R245 B.n403 B.n402 585
R246 B.n401 B.n400 585
R247 B.n399 B.n398 585
R248 B.n397 B.n396 585
R249 B.n395 B.n394 585
R250 B.n393 B.n392 585
R251 B.n391 B.n390 585
R252 B.n389 B.n388 585
R253 B.n387 B.n386 585
R254 B.n385 B.n384 585
R255 B.n383 B.n382 585
R256 B.n381 B.n380 585
R257 B.n379 B.n378 585
R258 B.n377 B.n376 585
R259 B.n375 B.n374 585
R260 B.n373 B.n372 585
R261 B.n371 B.n370 585
R262 B.n369 B.n368 585
R263 B.n367 B.n366 585
R264 B.n365 B.n364 585
R265 B.n363 B.n362 585
R266 B.n361 B.n360 585
R267 B.n359 B.n358 585
R268 B.n357 B.n356 585
R269 B.n355 B.n354 585
R270 B.n353 B.n352 585
R271 B.n351 B.n350 585
R272 B.n349 B.n348 585
R273 B.n347 B.n346 585
R274 B.n345 B.n344 585
R275 B.n343 B.n342 585
R276 B.n341 B.n340 585
R277 B.n339 B.n338 585
R278 B.n337 B.n336 585
R279 B.n335 B.n334 585
R280 B.n333 B.n332 585
R281 B.n331 B.n330 585
R282 B.n329 B.n328 585
R283 B.n327 B.n326 585
R284 B.n325 B.n324 585
R285 B.n323 B.n322 585
R286 B.n321 B.n320 585
R287 B.n319 B.n318 585
R288 B.n317 B.n316 585
R289 B.n315 B.n314 585
R290 B.n313 B.n312 585
R291 B.n311 B.n310 585
R292 B.n309 B.n308 585
R293 B.n307 B.n306 585
R294 B.n305 B.n304 585
R295 B.n303 B.n302 585
R296 B.n301 B.n300 585
R297 B.n299 B.n298 585
R298 B.n297 B.n296 585
R299 B.n295 B.n294 585
R300 B.n293 B.n292 585
R301 B.n291 B.n290 585
R302 B.n289 B.n288 585
R303 B.n287 B.n286 585
R304 B.n285 B.n284 585
R305 B.n283 B.n282 585
R306 B.n281 B.n280 585
R307 B.n279 B.n278 585
R308 B.n277 B.n276 585
R309 B.n275 B.n274 585
R310 B.n273 B.n272 585
R311 B.n271 B.n270 585
R312 B.n269 B.n268 585
R313 B.n267 B.n266 585
R314 B.n265 B.n264 585
R315 B.n263 B.n262 585
R316 B.n261 B.n260 585
R317 B.n259 B.n258 585
R318 B.n257 B.n256 585
R319 B.n255 B.n254 585
R320 B.n253 B.n252 585
R321 B.n251 B.n250 585
R322 B.n249 B.n248 585
R323 B.n247 B.n246 585
R324 B.n245 B.n244 585
R325 B.n243 B.n242 585
R326 B.n241 B.n240 585
R327 B.n239 B.n238 585
R328 B.n237 B.n236 585
R329 B.n235 B.n234 585
R330 B.n233 B.n232 585
R331 B.n231 B.n230 585
R332 B.n229 B.n228 585
R333 B.n227 B.n226 585
R334 B.n225 B.n224 585
R335 B.n223 B.n222 585
R336 B.n221 B.n220 585
R337 B.n219 B.n218 585
R338 B.n217 B.n216 585
R339 B.n215 B.n214 585
R340 B.n213 B.n212 585
R341 B.n152 B.n151 585
R342 B.n1212 B.n1211 585
R343 B.n1205 B.n205 585
R344 B.n205 B.n149 585
R345 B.n1204 B.n148 585
R346 B.n1216 B.n148 585
R347 B.n1203 B.n147 585
R348 B.n1217 B.n147 585
R349 B.n1202 B.n146 585
R350 B.n1218 B.n146 585
R351 B.n1201 B.n1200 585
R352 B.n1200 B.n142 585
R353 B.n1199 B.n141 585
R354 B.n1224 B.n141 585
R355 B.n1198 B.n140 585
R356 B.n1225 B.n140 585
R357 B.n1197 B.n139 585
R358 B.n1226 B.n139 585
R359 B.n1196 B.n1195 585
R360 B.n1195 B.n135 585
R361 B.n1194 B.n134 585
R362 B.n1232 B.n134 585
R363 B.n1193 B.n133 585
R364 B.n1233 B.n133 585
R365 B.n1192 B.n132 585
R366 B.n1234 B.n132 585
R367 B.n1191 B.n1190 585
R368 B.n1190 B.n128 585
R369 B.n1189 B.n127 585
R370 B.n1240 B.n127 585
R371 B.n1188 B.n126 585
R372 B.n1241 B.n126 585
R373 B.n1187 B.n125 585
R374 B.n1242 B.n125 585
R375 B.n1186 B.n1185 585
R376 B.n1185 B.n121 585
R377 B.n1184 B.n120 585
R378 B.n1248 B.n120 585
R379 B.n1183 B.n119 585
R380 B.n1249 B.n119 585
R381 B.n1182 B.n118 585
R382 B.n1250 B.n118 585
R383 B.n1181 B.n1180 585
R384 B.n1180 B.n114 585
R385 B.n1179 B.n113 585
R386 B.n1256 B.n113 585
R387 B.n1178 B.n112 585
R388 B.n1257 B.n112 585
R389 B.n1177 B.n111 585
R390 B.n1258 B.n111 585
R391 B.n1176 B.n1175 585
R392 B.n1175 B.n107 585
R393 B.n1174 B.n106 585
R394 B.n1264 B.n106 585
R395 B.n1173 B.n105 585
R396 B.n1265 B.n105 585
R397 B.n1172 B.n104 585
R398 B.n1266 B.n104 585
R399 B.n1171 B.n1170 585
R400 B.n1170 B.n100 585
R401 B.n1169 B.n99 585
R402 B.n1272 B.n99 585
R403 B.n1168 B.n98 585
R404 B.n1273 B.n98 585
R405 B.n1167 B.n97 585
R406 B.n1274 B.n97 585
R407 B.n1166 B.n1165 585
R408 B.n1165 B.n93 585
R409 B.n1164 B.n92 585
R410 B.n1280 B.n92 585
R411 B.n1163 B.n91 585
R412 B.n1281 B.n91 585
R413 B.n1162 B.n90 585
R414 B.n1282 B.n90 585
R415 B.n1161 B.n1160 585
R416 B.n1160 B.n86 585
R417 B.n1159 B.n85 585
R418 B.n1288 B.n85 585
R419 B.n1158 B.n84 585
R420 B.n1289 B.n84 585
R421 B.n1157 B.n83 585
R422 B.n1290 B.n83 585
R423 B.n1156 B.n1155 585
R424 B.n1155 B.n79 585
R425 B.n1154 B.n78 585
R426 B.n1296 B.n78 585
R427 B.n1153 B.n77 585
R428 B.n1297 B.n77 585
R429 B.n1152 B.n76 585
R430 B.n1298 B.n76 585
R431 B.n1151 B.n1150 585
R432 B.n1150 B.n72 585
R433 B.n1149 B.n71 585
R434 B.n1304 B.n71 585
R435 B.n1148 B.n70 585
R436 B.n1305 B.n70 585
R437 B.n1147 B.n69 585
R438 B.n1306 B.n69 585
R439 B.n1146 B.n1145 585
R440 B.n1145 B.n65 585
R441 B.n1144 B.n64 585
R442 B.n1312 B.n64 585
R443 B.n1143 B.n63 585
R444 B.n1313 B.n63 585
R445 B.n1142 B.n62 585
R446 B.n1314 B.n62 585
R447 B.n1141 B.n1140 585
R448 B.n1140 B.n58 585
R449 B.n1139 B.n57 585
R450 B.n1320 B.n57 585
R451 B.n1138 B.n56 585
R452 B.n1321 B.n56 585
R453 B.n1137 B.n55 585
R454 B.n1322 B.n55 585
R455 B.n1136 B.n1135 585
R456 B.n1135 B.n51 585
R457 B.n1134 B.n50 585
R458 B.n1328 B.n50 585
R459 B.n1133 B.n49 585
R460 B.n1329 B.n49 585
R461 B.n1132 B.n48 585
R462 B.n1330 B.n48 585
R463 B.n1131 B.n1130 585
R464 B.n1130 B.n44 585
R465 B.n1129 B.n43 585
R466 B.n1336 B.n43 585
R467 B.n1128 B.n42 585
R468 B.n1337 B.n42 585
R469 B.n1127 B.n41 585
R470 B.n1338 B.n41 585
R471 B.n1126 B.n1125 585
R472 B.n1125 B.n37 585
R473 B.n1124 B.n36 585
R474 B.n1344 B.n36 585
R475 B.n1123 B.n35 585
R476 B.n1345 B.n35 585
R477 B.n1122 B.n34 585
R478 B.n1346 B.n34 585
R479 B.n1121 B.n1120 585
R480 B.n1120 B.n30 585
R481 B.n1119 B.n29 585
R482 B.n1352 B.n29 585
R483 B.n1118 B.n28 585
R484 B.n1353 B.n28 585
R485 B.n1117 B.n27 585
R486 B.n1354 B.n27 585
R487 B.n1116 B.n1115 585
R488 B.n1115 B.n23 585
R489 B.n1114 B.n22 585
R490 B.n1360 B.n22 585
R491 B.n1113 B.n21 585
R492 B.n1361 B.n21 585
R493 B.n1112 B.n20 585
R494 B.n1362 B.n20 585
R495 B.n1111 B.n1110 585
R496 B.n1110 B.n16 585
R497 B.n1109 B.n15 585
R498 B.n1368 B.n15 585
R499 B.n1108 B.n14 585
R500 B.n1369 B.n14 585
R501 B.n1107 B.n13 585
R502 B.n1370 B.n13 585
R503 B.n1106 B.n1105 585
R504 B.n1105 B.n12 585
R505 B.n1104 B.n1103 585
R506 B.n1104 B.n8 585
R507 B.n1102 B.n7 585
R508 B.n1377 B.n7 585
R509 B.n1101 B.n6 585
R510 B.n1378 B.n6 585
R511 B.n1100 B.n5 585
R512 B.n1379 B.n5 585
R513 B.n1099 B.n1098 585
R514 B.n1098 B.n4 585
R515 B.n1097 B.n417 585
R516 B.n1097 B.n1096 585
R517 B.n1087 B.n418 585
R518 B.n419 B.n418 585
R519 B.n1089 B.n1088 585
R520 B.n1090 B.n1089 585
R521 B.n1086 B.n424 585
R522 B.n424 B.n423 585
R523 B.n1085 B.n1084 585
R524 B.n1084 B.n1083 585
R525 B.n426 B.n425 585
R526 B.n427 B.n426 585
R527 B.n1076 B.n1075 585
R528 B.n1077 B.n1076 585
R529 B.n1074 B.n432 585
R530 B.n432 B.n431 585
R531 B.n1073 B.n1072 585
R532 B.n1072 B.n1071 585
R533 B.n434 B.n433 585
R534 B.n435 B.n434 585
R535 B.n1064 B.n1063 585
R536 B.n1065 B.n1064 585
R537 B.n1062 B.n440 585
R538 B.n440 B.n439 585
R539 B.n1061 B.n1060 585
R540 B.n1060 B.n1059 585
R541 B.n442 B.n441 585
R542 B.n443 B.n442 585
R543 B.n1052 B.n1051 585
R544 B.n1053 B.n1052 585
R545 B.n1050 B.n448 585
R546 B.n448 B.n447 585
R547 B.n1049 B.n1048 585
R548 B.n1048 B.n1047 585
R549 B.n450 B.n449 585
R550 B.n451 B.n450 585
R551 B.n1040 B.n1039 585
R552 B.n1041 B.n1040 585
R553 B.n1038 B.n456 585
R554 B.n456 B.n455 585
R555 B.n1037 B.n1036 585
R556 B.n1036 B.n1035 585
R557 B.n458 B.n457 585
R558 B.n459 B.n458 585
R559 B.n1028 B.n1027 585
R560 B.n1029 B.n1028 585
R561 B.n1026 B.n464 585
R562 B.n464 B.n463 585
R563 B.n1025 B.n1024 585
R564 B.n1024 B.n1023 585
R565 B.n466 B.n465 585
R566 B.n467 B.n466 585
R567 B.n1016 B.n1015 585
R568 B.n1017 B.n1016 585
R569 B.n1014 B.n472 585
R570 B.n472 B.n471 585
R571 B.n1013 B.n1012 585
R572 B.n1012 B.n1011 585
R573 B.n474 B.n473 585
R574 B.n475 B.n474 585
R575 B.n1004 B.n1003 585
R576 B.n1005 B.n1004 585
R577 B.n1002 B.n479 585
R578 B.n483 B.n479 585
R579 B.n1001 B.n1000 585
R580 B.n1000 B.n999 585
R581 B.n481 B.n480 585
R582 B.n482 B.n481 585
R583 B.n992 B.n991 585
R584 B.n993 B.n992 585
R585 B.n990 B.n488 585
R586 B.n488 B.n487 585
R587 B.n989 B.n988 585
R588 B.n988 B.n987 585
R589 B.n490 B.n489 585
R590 B.n491 B.n490 585
R591 B.n980 B.n979 585
R592 B.n981 B.n980 585
R593 B.n978 B.n496 585
R594 B.n496 B.n495 585
R595 B.n977 B.n976 585
R596 B.n976 B.n975 585
R597 B.n498 B.n497 585
R598 B.n499 B.n498 585
R599 B.n968 B.n967 585
R600 B.n969 B.n968 585
R601 B.n966 B.n504 585
R602 B.n504 B.n503 585
R603 B.n965 B.n964 585
R604 B.n964 B.n963 585
R605 B.n506 B.n505 585
R606 B.n507 B.n506 585
R607 B.n956 B.n955 585
R608 B.n957 B.n956 585
R609 B.n954 B.n512 585
R610 B.n512 B.n511 585
R611 B.n953 B.n952 585
R612 B.n952 B.n951 585
R613 B.n514 B.n513 585
R614 B.n515 B.n514 585
R615 B.n944 B.n943 585
R616 B.n945 B.n944 585
R617 B.n942 B.n520 585
R618 B.n520 B.n519 585
R619 B.n941 B.n940 585
R620 B.n940 B.n939 585
R621 B.n522 B.n521 585
R622 B.n523 B.n522 585
R623 B.n932 B.n931 585
R624 B.n933 B.n932 585
R625 B.n930 B.n528 585
R626 B.n528 B.n527 585
R627 B.n929 B.n928 585
R628 B.n928 B.n927 585
R629 B.n530 B.n529 585
R630 B.n531 B.n530 585
R631 B.n920 B.n919 585
R632 B.n921 B.n920 585
R633 B.n918 B.n536 585
R634 B.n536 B.n535 585
R635 B.n917 B.n916 585
R636 B.n916 B.n915 585
R637 B.n538 B.n537 585
R638 B.n539 B.n538 585
R639 B.n908 B.n907 585
R640 B.n909 B.n908 585
R641 B.n906 B.n544 585
R642 B.n544 B.n543 585
R643 B.n905 B.n904 585
R644 B.n904 B.n903 585
R645 B.n546 B.n545 585
R646 B.n547 B.n546 585
R647 B.n896 B.n895 585
R648 B.n897 B.n896 585
R649 B.n894 B.n552 585
R650 B.n552 B.n551 585
R651 B.n893 B.n892 585
R652 B.n892 B.n891 585
R653 B.n554 B.n553 585
R654 B.n555 B.n554 585
R655 B.n884 B.n883 585
R656 B.n885 B.n884 585
R657 B.n882 B.n560 585
R658 B.n560 B.n559 585
R659 B.n881 B.n880 585
R660 B.n880 B.n879 585
R661 B.n562 B.n561 585
R662 B.n563 B.n562 585
R663 B.n872 B.n871 585
R664 B.n873 B.n872 585
R665 B.n870 B.n568 585
R666 B.n568 B.n567 585
R667 B.n869 B.n868 585
R668 B.n868 B.n867 585
R669 B.n570 B.n569 585
R670 B.n571 B.n570 585
R671 B.n860 B.n859 585
R672 B.n861 B.n860 585
R673 B.n858 B.n576 585
R674 B.n576 B.n575 585
R675 B.n857 B.n856 585
R676 B.n856 B.n855 585
R677 B.n578 B.n577 585
R678 B.n579 B.n578 585
R679 B.n851 B.n850 585
R680 B.n582 B.n581 585
R681 B.n847 B.n846 585
R682 B.n848 B.n847 585
R683 B.n845 B.n635 585
R684 B.n844 B.n843 585
R685 B.n842 B.n841 585
R686 B.n840 B.n839 585
R687 B.n838 B.n837 585
R688 B.n836 B.n835 585
R689 B.n834 B.n833 585
R690 B.n832 B.n831 585
R691 B.n830 B.n829 585
R692 B.n828 B.n827 585
R693 B.n826 B.n825 585
R694 B.n824 B.n823 585
R695 B.n822 B.n821 585
R696 B.n820 B.n819 585
R697 B.n818 B.n817 585
R698 B.n816 B.n815 585
R699 B.n814 B.n813 585
R700 B.n812 B.n811 585
R701 B.n810 B.n809 585
R702 B.n808 B.n807 585
R703 B.n806 B.n805 585
R704 B.n804 B.n803 585
R705 B.n802 B.n801 585
R706 B.n800 B.n799 585
R707 B.n798 B.n797 585
R708 B.n796 B.n795 585
R709 B.n794 B.n793 585
R710 B.n792 B.n791 585
R711 B.n790 B.n789 585
R712 B.n788 B.n787 585
R713 B.n786 B.n785 585
R714 B.n784 B.n783 585
R715 B.n782 B.n781 585
R716 B.n780 B.n779 585
R717 B.n778 B.n777 585
R718 B.n776 B.n775 585
R719 B.n774 B.n773 585
R720 B.n772 B.n771 585
R721 B.n770 B.n769 585
R722 B.n768 B.n767 585
R723 B.n766 B.n765 585
R724 B.n764 B.n763 585
R725 B.n762 B.n761 585
R726 B.n760 B.n759 585
R727 B.n758 B.n757 585
R728 B.n755 B.n754 585
R729 B.n753 B.n752 585
R730 B.n751 B.n750 585
R731 B.n749 B.n748 585
R732 B.n747 B.n746 585
R733 B.n745 B.n744 585
R734 B.n743 B.n742 585
R735 B.n741 B.n740 585
R736 B.n739 B.n738 585
R737 B.n737 B.n736 585
R738 B.n734 B.n733 585
R739 B.n732 B.n731 585
R740 B.n730 B.n729 585
R741 B.n728 B.n727 585
R742 B.n726 B.n725 585
R743 B.n724 B.n723 585
R744 B.n722 B.n721 585
R745 B.n720 B.n719 585
R746 B.n718 B.n717 585
R747 B.n716 B.n715 585
R748 B.n714 B.n713 585
R749 B.n712 B.n711 585
R750 B.n710 B.n709 585
R751 B.n708 B.n707 585
R752 B.n706 B.n705 585
R753 B.n704 B.n703 585
R754 B.n702 B.n701 585
R755 B.n700 B.n699 585
R756 B.n698 B.n697 585
R757 B.n696 B.n695 585
R758 B.n694 B.n693 585
R759 B.n692 B.n691 585
R760 B.n690 B.n689 585
R761 B.n688 B.n687 585
R762 B.n686 B.n685 585
R763 B.n684 B.n683 585
R764 B.n682 B.n681 585
R765 B.n680 B.n679 585
R766 B.n678 B.n677 585
R767 B.n676 B.n675 585
R768 B.n674 B.n673 585
R769 B.n672 B.n671 585
R770 B.n670 B.n669 585
R771 B.n668 B.n667 585
R772 B.n666 B.n665 585
R773 B.n664 B.n663 585
R774 B.n662 B.n661 585
R775 B.n660 B.n659 585
R776 B.n658 B.n657 585
R777 B.n656 B.n655 585
R778 B.n654 B.n653 585
R779 B.n652 B.n651 585
R780 B.n650 B.n649 585
R781 B.n648 B.n647 585
R782 B.n646 B.n645 585
R783 B.n644 B.n643 585
R784 B.n642 B.n641 585
R785 B.n640 B.n634 585
R786 B.n848 B.n634 585
R787 B.n852 B.n580 585
R788 B.n580 B.n579 585
R789 B.n854 B.n853 585
R790 B.n855 B.n854 585
R791 B.n574 B.n573 585
R792 B.n575 B.n574 585
R793 B.n863 B.n862 585
R794 B.n862 B.n861 585
R795 B.n864 B.n572 585
R796 B.n572 B.n571 585
R797 B.n866 B.n865 585
R798 B.n867 B.n866 585
R799 B.n566 B.n565 585
R800 B.n567 B.n566 585
R801 B.n875 B.n874 585
R802 B.n874 B.n873 585
R803 B.n876 B.n564 585
R804 B.n564 B.n563 585
R805 B.n878 B.n877 585
R806 B.n879 B.n878 585
R807 B.n558 B.n557 585
R808 B.n559 B.n558 585
R809 B.n887 B.n886 585
R810 B.n886 B.n885 585
R811 B.n888 B.n556 585
R812 B.n556 B.n555 585
R813 B.n890 B.n889 585
R814 B.n891 B.n890 585
R815 B.n550 B.n549 585
R816 B.n551 B.n550 585
R817 B.n899 B.n898 585
R818 B.n898 B.n897 585
R819 B.n900 B.n548 585
R820 B.n548 B.n547 585
R821 B.n902 B.n901 585
R822 B.n903 B.n902 585
R823 B.n542 B.n541 585
R824 B.n543 B.n542 585
R825 B.n911 B.n910 585
R826 B.n910 B.n909 585
R827 B.n912 B.n540 585
R828 B.n540 B.n539 585
R829 B.n914 B.n913 585
R830 B.n915 B.n914 585
R831 B.n534 B.n533 585
R832 B.n535 B.n534 585
R833 B.n923 B.n922 585
R834 B.n922 B.n921 585
R835 B.n924 B.n532 585
R836 B.n532 B.n531 585
R837 B.n926 B.n925 585
R838 B.n927 B.n926 585
R839 B.n526 B.n525 585
R840 B.n527 B.n526 585
R841 B.n935 B.n934 585
R842 B.n934 B.n933 585
R843 B.n936 B.n524 585
R844 B.n524 B.n523 585
R845 B.n938 B.n937 585
R846 B.n939 B.n938 585
R847 B.n518 B.n517 585
R848 B.n519 B.n518 585
R849 B.n947 B.n946 585
R850 B.n946 B.n945 585
R851 B.n948 B.n516 585
R852 B.n516 B.n515 585
R853 B.n950 B.n949 585
R854 B.n951 B.n950 585
R855 B.n510 B.n509 585
R856 B.n511 B.n510 585
R857 B.n959 B.n958 585
R858 B.n958 B.n957 585
R859 B.n960 B.n508 585
R860 B.n508 B.n507 585
R861 B.n962 B.n961 585
R862 B.n963 B.n962 585
R863 B.n502 B.n501 585
R864 B.n503 B.n502 585
R865 B.n971 B.n970 585
R866 B.n970 B.n969 585
R867 B.n972 B.n500 585
R868 B.n500 B.n499 585
R869 B.n974 B.n973 585
R870 B.n975 B.n974 585
R871 B.n494 B.n493 585
R872 B.n495 B.n494 585
R873 B.n983 B.n982 585
R874 B.n982 B.n981 585
R875 B.n984 B.n492 585
R876 B.n492 B.n491 585
R877 B.n986 B.n985 585
R878 B.n987 B.n986 585
R879 B.n486 B.n485 585
R880 B.n487 B.n486 585
R881 B.n995 B.n994 585
R882 B.n994 B.n993 585
R883 B.n996 B.n484 585
R884 B.n484 B.n482 585
R885 B.n998 B.n997 585
R886 B.n999 B.n998 585
R887 B.n478 B.n477 585
R888 B.n483 B.n478 585
R889 B.n1007 B.n1006 585
R890 B.n1006 B.n1005 585
R891 B.n1008 B.n476 585
R892 B.n476 B.n475 585
R893 B.n1010 B.n1009 585
R894 B.n1011 B.n1010 585
R895 B.n470 B.n469 585
R896 B.n471 B.n470 585
R897 B.n1019 B.n1018 585
R898 B.n1018 B.n1017 585
R899 B.n1020 B.n468 585
R900 B.n468 B.n467 585
R901 B.n1022 B.n1021 585
R902 B.n1023 B.n1022 585
R903 B.n462 B.n461 585
R904 B.n463 B.n462 585
R905 B.n1031 B.n1030 585
R906 B.n1030 B.n1029 585
R907 B.n1032 B.n460 585
R908 B.n460 B.n459 585
R909 B.n1034 B.n1033 585
R910 B.n1035 B.n1034 585
R911 B.n454 B.n453 585
R912 B.n455 B.n454 585
R913 B.n1043 B.n1042 585
R914 B.n1042 B.n1041 585
R915 B.n1044 B.n452 585
R916 B.n452 B.n451 585
R917 B.n1046 B.n1045 585
R918 B.n1047 B.n1046 585
R919 B.n446 B.n445 585
R920 B.n447 B.n446 585
R921 B.n1055 B.n1054 585
R922 B.n1054 B.n1053 585
R923 B.n1056 B.n444 585
R924 B.n444 B.n443 585
R925 B.n1058 B.n1057 585
R926 B.n1059 B.n1058 585
R927 B.n438 B.n437 585
R928 B.n439 B.n438 585
R929 B.n1067 B.n1066 585
R930 B.n1066 B.n1065 585
R931 B.n1068 B.n436 585
R932 B.n436 B.n435 585
R933 B.n1070 B.n1069 585
R934 B.n1071 B.n1070 585
R935 B.n430 B.n429 585
R936 B.n431 B.n430 585
R937 B.n1079 B.n1078 585
R938 B.n1078 B.n1077 585
R939 B.n1080 B.n428 585
R940 B.n428 B.n427 585
R941 B.n1082 B.n1081 585
R942 B.n1083 B.n1082 585
R943 B.n422 B.n421 585
R944 B.n423 B.n422 585
R945 B.n1092 B.n1091 585
R946 B.n1091 B.n1090 585
R947 B.n1093 B.n420 585
R948 B.n420 B.n419 585
R949 B.n1095 B.n1094 585
R950 B.n1096 B.n1095 585
R951 B.n3 B.n0 585
R952 B.n4 B.n3 585
R953 B.n1376 B.n1 585
R954 B.n1377 B.n1376 585
R955 B.n1375 B.n1374 585
R956 B.n1375 B.n8 585
R957 B.n1373 B.n9 585
R958 B.n12 B.n9 585
R959 B.n1372 B.n1371 585
R960 B.n1371 B.n1370 585
R961 B.n11 B.n10 585
R962 B.n1369 B.n11 585
R963 B.n1367 B.n1366 585
R964 B.n1368 B.n1367 585
R965 B.n1365 B.n17 585
R966 B.n17 B.n16 585
R967 B.n1364 B.n1363 585
R968 B.n1363 B.n1362 585
R969 B.n19 B.n18 585
R970 B.n1361 B.n19 585
R971 B.n1359 B.n1358 585
R972 B.n1360 B.n1359 585
R973 B.n1357 B.n24 585
R974 B.n24 B.n23 585
R975 B.n1356 B.n1355 585
R976 B.n1355 B.n1354 585
R977 B.n26 B.n25 585
R978 B.n1353 B.n26 585
R979 B.n1351 B.n1350 585
R980 B.n1352 B.n1351 585
R981 B.n1349 B.n31 585
R982 B.n31 B.n30 585
R983 B.n1348 B.n1347 585
R984 B.n1347 B.n1346 585
R985 B.n33 B.n32 585
R986 B.n1345 B.n33 585
R987 B.n1343 B.n1342 585
R988 B.n1344 B.n1343 585
R989 B.n1341 B.n38 585
R990 B.n38 B.n37 585
R991 B.n1340 B.n1339 585
R992 B.n1339 B.n1338 585
R993 B.n40 B.n39 585
R994 B.n1337 B.n40 585
R995 B.n1335 B.n1334 585
R996 B.n1336 B.n1335 585
R997 B.n1333 B.n45 585
R998 B.n45 B.n44 585
R999 B.n1332 B.n1331 585
R1000 B.n1331 B.n1330 585
R1001 B.n47 B.n46 585
R1002 B.n1329 B.n47 585
R1003 B.n1327 B.n1326 585
R1004 B.n1328 B.n1327 585
R1005 B.n1325 B.n52 585
R1006 B.n52 B.n51 585
R1007 B.n1324 B.n1323 585
R1008 B.n1323 B.n1322 585
R1009 B.n54 B.n53 585
R1010 B.n1321 B.n54 585
R1011 B.n1319 B.n1318 585
R1012 B.n1320 B.n1319 585
R1013 B.n1317 B.n59 585
R1014 B.n59 B.n58 585
R1015 B.n1316 B.n1315 585
R1016 B.n1315 B.n1314 585
R1017 B.n61 B.n60 585
R1018 B.n1313 B.n61 585
R1019 B.n1311 B.n1310 585
R1020 B.n1312 B.n1311 585
R1021 B.n1309 B.n66 585
R1022 B.n66 B.n65 585
R1023 B.n1308 B.n1307 585
R1024 B.n1307 B.n1306 585
R1025 B.n68 B.n67 585
R1026 B.n1305 B.n68 585
R1027 B.n1303 B.n1302 585
R1028 B.n1304 B.n1303 585
R1029 B.n1301 B.n73 585
R1030 B.n73 B.n72 585
R1031 B.n1300 B.n1299 585
R1032 B.n1299 B.n1298 585
R1033 B.n75 B.n74 585
R1034 B.n1297 B.n75 585
R1035 B.n1295 B.n1294 585
R1036 B.n1296 B.n1295 585
R1037 B.n1293 B.n80 585
R1038 B.n80 B.n79 585
R1039 B.n1292 B.n1291 585
R1040 B.n1291 B.n1290 585
R1041 B.n82 B.n81 585
R1042 B.n1289 B.n82 585
R1043 B.n1287 B.n1286 585
R1044 B.n1288 B.n1287 585
R1045 B.n1285 B.n87 585
R1046 B.n87 B.n86 585
R1047 B.n1284 B.n1283 585
R1048 B.n1283 B.n1282 585
R1049 B.n89 B.n88 585
R1050 B.n1281 B.n89 585
R1051 B.n1279 B.n1278 585
R1052 B.n1280 B.n1279 585
R1053 B.n1277 B.n94 585
R1054 B.n94 B.n93 585
R1055 B.n1276 B.n1275 585
R1056 B.n1275 B.n1274 585
R1057 B.n96 B.n95 585
R1058 B.n1273 B.n96 585
R1059 B.n1271 B.n1270 585
R1060 B.n1272 B.n1271 585
R1061 B.n1269 B.n101 585
R1062 B.n101 B.n100 585
R1063 B.n1268 B.n1267 585
R1064 B.n1267 B.n1266 585
R1065 B.n103 B.n102 585
R1066 B.n1265 B.n103 585
R1067 B.n1263 B.n1262 585
R1068 B.n1264 B.n1263 585
R1069 B.n1261 B.n108 585
R1070 B.n108 B.n107 585
R1071 B.n1260 B.n1259 585
R1072 B.n1259 B.n1258 585
R1073 B.n110 B.n109 585
R1074 B.n1257 B.n110 585
R1075 B.n1255 B.n1254 585
R1076 B.n1256 B.n1255 585
R1077 B.n1253 B.n115 585
R1078 B.n115 B.n114 585
R1079 B.n1252 B.n1251 585
R1080 B.n1251 B.n1250 585
R1081 B.n117 B.n116 585
R1082 B.n1249 B.n117 585
R1083 B.n1247 B.n1246 585
R1084 B.n1248 B.n1247 585
R1085 B.n1245 B.n122 585
R1086 B.n122 B.n121 585
R1087 B.n1244 B.n1243 585
R1088 B.n1243 B.n1242 585
R1089 B.n124 B.n123 585
R1090 B.n1241 B.n124 585
R1091 B.n1239 B.n1238 585
R1092 B.n1240 B.n1239 585
R1093 B.n1237 B.n129 585
R1094 B.n129 B.n128 585
R1095 B.n1236 B.n1235 585
R1096 B.n1235 B.n1234 585
R1097 B.n131 B.n130 585
R1098 B.n1233 B.n131 585
R1099 B.n1231 B.n1230 585
R1100 B.n1232 B.n1231 585
R1101 B.n1229 B.n136 585
R1102 B.n136 B.n135 585
R1103 B.n1228 B.n1227 585
R1104 B.n1227 B.n1226 585
R1105 B.n138 B.n137 585
R1106 B.n1225 B.n138 585
R1107 B.n1223 B.n1222 585
R1108 B.n1224 B.n1223 585
R1109 B.n1221 B.n143 585
R1110 B.n143 B.n142 585
R1111 B.n1220 B.n1219 585
R1112 B.n1219 B.n1218 585
R1113 B.n145 B.n144 585
R1114 B.n1217 B.n145 585
R1115 B.n1215 B.n1214 585
R1116 B.n1216 B.n1215 585
R1117 B.n1213 B.n150 585
R1118 B.n150 B.n149 585
R1119 B.n1380 B.n1379 585
R1120 B.n1378 B.n2 585
R1121 B.n1211 B.n150 535.745
R1122 B.n1207 B.n205 535.745
R1123 B.n634 B.n578 535.745
R1124 B.n850 B.n580 535.745
R1125 B.n209 B.t14 297.101
R1126 B.n206 B.t10 297.101
R1127 B.n638 B.t21 297.101
R1128 B.n636 B.t17 297.101
R1129 B.n1209 B.n1208 256.663
R1130 B.n1209 B.n203 256.663
R1131 B.n1209 B.n202 256.663
R1132 B.n1209 B.n201 256.663
R1133 B.n1209 B.n200 256.663
R1134 B.n1209 B.n199 256.663
R1135 B.n1209 B.n198 256.663
R1136 B.n1209 B.n197 256.663
R1137 B.n1209 B.n196 256.663
R1138 B.n1209 B.n195 256.663
R1139 B.n1209 B.n194 256.663
R1140 B.n1209 B.n193 256.663
R1141 B.n1209 B.n192 256.663
R1142 B.n1209 B.n191 256.663
R1143 B.n1209 B.n190 256.663
R1144 B.n1209 B.n189 256.663
R1145 B.n1209 B.n188 256.663
R1146 B.n1209 B.n187 256.663
R1147 B.n1209 B.n186 256.663
R1148 B.n1209 B.n185 256.663
R1149 B.n1209 B.n184 256.663
R1150 B.n1209 B.n183 256.663
R1151 B.n1209 B.n182 256.663
R1152 B.n1209 B.n181 256.663
R1153 B.n1209 B.n180 256.663
R1154 B.n1209 B.n179 256.663
R1155 B.n1209 B.n178 256.663
R1156 B.n1209 B.n177 256.663
R1157 B.n1209 B.n176 256.663
R1158 B.n1209 B.n175 256.663
R1159 B.n1209 B.n174 256.663
R1160 B.n1209 B.n173 256.663
R1161 B.n1209 B.n172 256.663
R1162 B.n1209 B.n171 256.663
R1163 B.n1209 B.n170 256.663
R1164 B.n1209 B.n169 256.663
R1165 B.n1209 B.n168 256.663
R1166 B.n1209 B.n167 256.663
R1167 B.n1209 B.n166 256.663
R1168 B.n1209 B.n165 256.663
R1169 B.n1209 B.n164 256.663
R1170 B.n1209 B.n163 256.663
R1171 B.n1209 B.n162 256.663
R1172 B.n1209 B.n161 256.663
R1173 B.n1209 B.n160 256.663
R1174 B.n1209 B.n159 256.663
R1175 B.n1209 B.n158 256.663
R1176 B.n1209 B.n157 256.663
R1177 B.n1209 B.n156 256.663
R1178 B.n1209 B.n155 256.663
R1179 B.n1209 B.n154 256.663
R1180 B.n1209 B.n153 256.663
R1181 B.n1210 B.n1209 256.663
R1182 B.n849 B.n848 256.663
R1183 B.n848 B.n583 256.663
R1184 B.n848 B.n584 256.663
R1185 B.n848 B.n585 256.663
R1186 B.n848 B.n586 256.663
R1187 B.n848 B.n587 256.663
R1188 B.n848 B.n588 256.663
R1189 B.n848 B.n589 256.663
R1190 B.n848 B.n590 256.663
R1191 B.n848 B.n591 256.663
R1192 B.n848 B.n592 256.663
R1193 B.n848 B.n593 256.663
R1194 B.n848 B.n594 256.663
R1195 B.n848 B.n595 256.663
R1196 B.n848 B.n596 256.663
R1197 B.n848 B.n597 256.663
R1198 B.n848 B.n598 256.663
R1199 B.n848 B.n599 256.663
R1200 B.n848 B.n600 256.663
R1201 B.n848 B.n601 256.663
R1202 B.n848 B.n602 256.663
R1203 B.n848 B.n603 256.663
R1204 B.n848 B.n604 256.663
R1205 B.n848 B.n605 256.663
R1206 B.n848 B.n606 256.663
R1207 B.n848 B.n607 256.663
R1208 B.n848 B.n608 256.663
R1209 B.n848 B.n609 256.663
R1210 B.n848 B.n610 256.663
R1211 B.n848 B.n611 256.663
R1212 B.n848 B.n612 256.663
R1213 B.n848 B.n613 256.663
R1214 B.n848 B.n614 256.663
R1215 B.n848 B.n615 256.663
R1216 B.n848 B.n616 256.663
R1217 B.n848 B.n617 256.663
R1218 B.n848 B.n618 256.663
R1219 B.n848 B.n619 256.663
R1220 B.n848 B.n620 256.663
R1221 B.n848 B.n621 256.663
R1222 B.n848 B.n622 256.663
R1223 B.n848 B.n623 256.663
R1224 B.n848 B.n624 256.663
R1225 B.n848 B.n625 256.663
R1226 B.n848 B.n626 256.663
R1227 B.n848 B.n627 256.663
R1228 B.n848 B.n628 256.663
R1229 B.n848 B.n629 256.663
R1230 B.n848 B.n630 256.663
R1231 B.n848 B.n631 256.663
R1232 B.n848 B.n632 256.663
R1233 B.n848 B.n633 256.663
R1234 B.n1382 B.n1381 256.663
R1235 B.n212 B.n152 163.367
R1236 B.n216 B.n215 163.367
R1237 B.n220 B.n219 163.367
R1238 B.n224 B.n223 163.367
R1239 B.n228 B.n227 163.367
R1240 B.n232 B.n231 163.367
R1241 B.n236 B.n235 163.367
R1242 B.n240 B.n239 163.367
R1243 B.n244 B.n243 163.367
R1244 B.n248 B.n247 163.367
R1245 B.n252 B.n251 163.367
R1246 B.n256 B.n255 163.367
R1247 B.n260 B.n259 163.367
R1248 B.n264 B.n263 163.367
R1249 B.n268 B.n267 163.367
R1250 B.n272 B.n271 163.367
R1251 B.n276 B.n275 163.367
R1252 B.n280 B.n279 163.367
R1253 B.n284 B.n283 163.367
R1254 B.n288 B.n287 163.367
R1255 B.n292 B.n291 163.367
R1256 B.n296 B.n295 163.367
R1257 B.n300 B.n299 163.367
R1258 B.n304 B.n303 163.367
R1259 B.n308 B.n307 163.367
R1260 B.n312 B.n311 163.367
R1261 B.n316 B.n315 163.367
R1262 B.n320 B.n319 163.367
R1263 B.n324 B.n323 163.367
R1264 B.n328 B.n327 163.367
R1265 B.n332 B.n331 163.367
R1266 B.n336 B.n335 163.367
R1267 B.n340 B.n339 163.367
R1268 B.n344 B.n343 163.367
R1269 B.n348 B.n347 163.367
R1270 B.n352 B.n351 163.367
R1271 B.n356 B.n355 163.367
R1272 B.n360 B.n359 163.367
R1273 B.n364 B.n363 163.367
R1274 B.n368 B.n367 163.367
R1275 B.n372 B.n371 163.367
R1276 B.n376 B.n375 163.367
R1277 B.n380 B.n379 163.367
R1278 B.n384 B.n383 163.367
R1279 B.n388 B.n387 163.367
R1280 B.n392 B.n391 163.367
R1281 B.n396 B.n395 163.367
R1282 B.n400 B.n399 163.367
R1283 B.n404 B.n403 163.367
R1284 B.n408 B.n407 163.367
R1285 B.n412 B.n411 163.367
R1286 B.n414 B.n204 163.367
R1287 B.n856 B.n578 163.367
R1288 B.n856 B.n576 163.367
R1289 B.n860 B.n576 163.367
R1290 B.n860 B.n570 163.367
R1291 B.n868 B.n570 163.367
R1292 B.n868 B.n568 163.367
R1293 B.n872 B.n568 163.367
R1294 B.n872 B.n562 163.367
R1295 B.n880 B.n562 163.367
R1296 B.n880 B.n560 163.367
R1297 B.n884 B.n560 163.367
R1298 B.n884 B.n554 163.367
R1299 B.n892 B.n554 163.367
R1300 B.n892 B.n552 163.367
R1301 B.n896 B.n552 163.367
R1302 B.n896 B.n546 163.367
R1303 B.n904 B.n546 163.367
R1304 B.n904 B.n544 163.367
R1305 B.n908 B.n544 163.367
R1306 B.n908 B.n538 163.367
R1307 B.n916 B.n538 163.367
R1308 B.n916 B.n536 163.367
R1309 B.n920 B.n536 163.367
R1310 B.n920 B.n530 163.367
R1311 B.n928 B.n530 163.367
R1312 B.n928 B.n528 163.367
R1313 B.n932 B.n528 163.367
R1314 B.n932 B.n522 163.367
R1315 B.n940 B.n522 163.367
R1316 B.n940 B.n520 163.367
R1317 B.n944 B.n520 163.367
R1318 B.n944 B.n514 163.367
R1319 B.n952 B.n514 163.367
R1320 B.n952 B.n512 163.367
R1321 B.n956 B.n512 163.367
R1322 B.n956 B.n506 163.367
R1323 B.n964 B.n506 163.367
R1324 B.n964 B.n504 163.367
R1325 B.n968 B.n504 163.367
R1326 B.n968 B.n498 163.367
R1327 B.n976 B.n498 163.367
R1328 B.n976 B.n496 163.367
R1329 B.n980 B.n496 163.367
R1330 B.n980 B.n490 163.367
R1331 B.n988 B.n490 163.367
R1332 B.n988 B.n488 163.367
R1333 B.n992 B.n488 163.367
R1334 B.n992 B.n481 163.367
R1335 B.n1000 B.n481 163.367
R1336 B.n1000 B.n479 163.367
R1337 B.n1004 B.n479 163.367
R1338 B.n1004 B.n474 163.367
R1339 B.n1012 B.n474 163.367
R1340 B.n1012 B.n472 163.367
R1341 B.n1016 B.n472 163.367
R1342 B.n1016 B.n466 163.367
R1343 B.n1024 B.n466 163.367
R1344 B.n1024 B.n464 163.367
R1345 B.n1028 B.n464 163.367
R1346 B.n1028 B.n458 163.367
R1347 B.n1036 B.n458 163.367
R1348 B.n1036 B.n456 163.367
R1349 B.n1040 B.n456 163.367
R1350 B.n1040 B.n450 163.367
R1351 B.n1048 B.n450 163.367
R1352 B.n1048 B.n448 163.367
R1353 B.n1052 B.n448 163.367
R1354 B.n1052 B.n442 163.367
R1355 B.n1060 B.n442 163.367
R1356 B.n1060 B.n440 163.367
R1357 B.n1064 B.n440 163.367
R1358 B.n1064 B.n434 163.367
R1359 B.n1072 B.n434 163.367
R1360 B.n1072 B.n432 163.367
R1361 B.n1076 B.n432 163.367
R1362 B.n1076 B.n426 163.367
R1363 B.n1084 B.n426 163.367
R1364 B.n1084 B.n424 163.367
R1365 B.n1089 B.n424 163.367
R1366 B.n1089 B.n418 163.367
R1367 B.n1097 B.n418 163.367
R1368 B.n1098 B.n1097 163.367
R1369 B.n1098 B.n5 163.367
R1370 B.n6 B.n5 163.367
R1371 B.n7 B.n6 163.367
R1372 B.n1104 B.n7 163.367
R1373 B.n1105 B.n1104 163.367
R1374 B.n1105 B.n13 163.367
R1375 B.n14 B.n13 163.367
R1376 B.n15 B.n14 163.367
R1377 B.n1110 B.n15 163.367
R1378 B.n1110 B.n20 163.367
R1379 B.n21 B.n20 163.367
R1380 B.n22 B.n21 163.367
R1381 B.n1115 B.n22 163.367
R1382 B.n1115 B.n27 163.367
R1383 B.n28 B.n27 163.367
R1384 B.n29 B.n28 163.367
R1385 B.n1120 B.n29 163.367
R1386 B.n1120 B.n34 163.367
R1387 B.n35 B.n34 163.367
R1388 B.n36 B.n35 163.367
R1389 B.n1125 B.n36 163.367
R1390 B.n1125 B.n41 163.367
R1391 B.n42 B.n41 163.367
R1392 B.n43 B.n42 163.367
R1393 B.n1130 B.n43 163.367
R1394 B.n1130 B.n48 163.367
R1395 B.n49 B.n48 163.367
R1396 B.n50 B.n49 163.367
R1397 B.n1135 B.n50 163.367
R1398 B.n1135 B.n55 163.367
R1399 B.n56 B.n55 163.367
R1400 B.n57 B.n56 163.367
R1401 B.n1140 B.n57 163.367
R1402 B.n1140 B.n62 163.367
R1403 B.n63 B.n62 163.367
R1404 B.n64 B.n63 163.367
R1405 B.n1145 B.n64 163.367
R1406 B.n1145 B.n69 163.367
R1407 B.n70 B.n69 163.367
R1408 B.n71 B.n70 163.367
R1409 B.n1150 B.n71 163.367
R1410 B.n1150 B.n76 163.367
R1411 B.n77 B.n76 163.367
R1412 B.n78 B.n77 163.367
R1413 B.n1155 B.n78 163.367
R1414 B.n1155 B.n83 163.367
R1415 B.n84 B.n83 163.367
R1416 B.n85 B.n84 163.367
R1417 B.n1160 B.n85 163.367
R1418 B.n1160 B.n90 163.367
R1419 B.n91 B.n90 163.367
R1420 B.n92 B.n91 163.367
R1421 B.n1165 B.n92 163.367
R1422 B.n1165 B.n97 163.367
R1423 B.n98 B.n97 163.367
R1424 B.n99 B.n98 163.367
R1425 B.n1170 B.n99 163.367
R1426 B.n1170 B.n104 163.367
R1427 B.n105 B.n104 163.367
R1428 B.n106 B.n105 163.367
R1429 B.n1175 B.n106 163.367
R1430 B.n1175 B.n111 163.367
R1431 B.n112 B.n111 163.367
R1432 B.n113 B.n112 163.367
R1433 B.n1180 B.n113 163.367
R1434 B.n1180 B.n118 163.367
R1435 B.n119 B.n118 163.367
R1436 B.n120 B.n119 163.367
R1437 B.n1185 B.n120 163.367
R1438 B.n1185 B.n125 163.367
R1439 B.n126 B.n125 163.367
R1440 B.n127 B.n126 163.367
R1441 B.n1190 B.n127 163.367
R1442 B.n1190 B.n132 163.367
R1443 B.n133 B.n132 163.367
R1444 B.n134 B.n133 163.367
R1445 B.n1195 B.n134 163.367
R1446 B.n1195 B.n139 163.367
R1447 B.n140 B.n139 163.367
R1448 B.n141 B.n140 163.367
R1449 B.n1200 B.n141 163.367
R1450 B.n1200 B.n146 163.367
R1451 B.n147 B.n146 163.367
R1452 B.n148 B.n147 163.367
R1453 B.n205 B.n148 163.367
R1454 B.n847 B.n582 163.367
R1455 B.n847 B.n635 163.367
R1456 B.n843 B.n842 163.367
R1457 B.n839 B.n838 163.367
R1458 B.n835 B.n834 163.367
R1459 B.n831 B.n830 163.367
R1460 B.n827 B.n826 163.367
R1461 B.n823 B.n822 163.367
R1462 B.n819 B.n818 163.367
R1463 B.n815 B.n814 163.367
R1464 B.n811 B.n810 163.367
R1465 B.n807 B.n806 163.367
R1466 B.n803 B.n802 163.367
R1467 B.n799 B.n798 163.367
R1468 B.n795 B.n794 163.367
R1469 B.n791 B.n790 163.367
R1470 B.n787 B.n786 163.367
R1471 B.n783 B.n782 163.367
R1472 B.n779 B.n778 163.367
R1473 B.n775 B.n774 163.367
R1474 B.n771 B.n770 163.367
R1475 B.n767 B.n766 163.367
R1476 B.n763 B.n762 163.367
R1477 B.n759 B.n758 163.367
R1478 B.n754 B.n753 163.367
R1479 B.n750 B.n749 163.367
R1480 B.n746 B.n745 163.367
R1481 B.n742 B.n741 163.367
R1482 B.n738 B.n737 163.367
R1483 B.n733 B.n732 163.367
R1484 B.n729 B.n728 163.367
R1485 B.n725 B.n724 163.367
R1486 B.n721 B.n720 163.367
R1487 B.n717 B.n716 163.367
R1488 B.n713 B.n712 163.367
R1489 B.n709 B.n708 163.367
R1490 B.n705 B.n704 163.367
R1491 B.n701 B.n700 163.367
R1492 B.n697 B.n696 163.367
R1493 B.n693 B.n692 163.367
R1494 B.n689 B.n688 163.367
R1495 B.n685 B.n684 163.367
R1496 B.n681 B.n680 163.367
R1497 B.n677 B.n676 163.367
R1498 B.n673 B.n672 163.367
R1499 B.n669 B.n668 163.367
R1500 B.n665 B.n664 163.367
R1501 B.n661 B.n660 163.367
R1502 B.n657 B.n656 163.367
R1503 B.n653 B.n652 163.367
R1504 B.n649 B.n648 163.367
R1505 B.n645 B.n644 163.367
R1506 B.n641 B.n634 163.367
R1507 B.n854 B.n580 163.367
R1508 B.n854 B.n574 163.367
R1509 B.n862 B.n574 163.367
R1510 B.n862 B.n572 163.367
R1511 B.n866 B.n572 163.367
R1512 B.n866 B.n566 163.367
R1513 B.n874 B.n566 163.367
R1514 B.n874 B.n564 163.367
R1515 B.n878 B.n564 163.367
R1516 B.n878 B.n558 163.367
R1517 B.n886 B.n558 163.367
R1518 B.n886 B.n556 163.367
R1519 B.n890 B.n556 163.367
R1520 B.n890 B.n550 163.367
R1521 B.n898 B.n550 163.367
R1522 B.n898 B.n548 163.367
R1523 B.n902 B.n548 163.367
R1524 B.n902 B.n542 163.367
R1525 B.n910 B.n542 163.367
R1526 B.n910 B.n540 163.367
R1527 B.n914 B.n540 163.367
R1528 B.n914 B.n534 163.367
R1529 B.n922 B.n534 163.367
R1530 B.n922 B.n532 163.367
R1531 B.n926 B.n532 163.367
R1532 B.n926 B.n526 163.367
R1533 B.n934 B.n526 163.367
R1534 B.n934 B.n524 163.367
R1535 B.n938 B.n524 163.367
R1536 B.n938 B.n518 163.367
R1537 B.n946 B.n518 163.367
R1538 B.n946 B.n516 163.367
R1539 B.n950 B.n516 163.367
R1540 B.n950 B.n510 163.367
R1541 B.n958 B.n510 163.367
R1542 B.n958 B.n508 163.367
R1543 B.n962 B.n508 163.367
R1544 B.n962 B.n502 163.367
R1545 B.n970 B.n502 163.367
R1546 B.n970 B.n500 163.367
R1547 B.n974 B.n500 163.367
R1548 B.n974 B.n494 163.367
R1549 B.n982 B.n494 163.367
R1550 B.n982 B.n492 163.367
R1551 B.n986 B.n492 163.367
R1552 B.n986 B.n486 163.367
R1553 B.n994 B.n486 163.367
R1554 B.n994 B.n484 163.367
R1555 B.n998 B.n484 163.367
R1556 B.n998 B.n478 163.367
R1557 B.n1006 B.n478 163.367
R1558 B.n1006 B.n476 163.367
R1559 B.n1010 B.n476 163.367
R1560 B.n1010 B.n470 163.367
R1561 B.n1018 B.n470 163.367
R1562 B.n1018 B.n468 163.367
R1563 B.n1022 B.n468 163.367
R1564 B.n1022 B.n462 163.367
R1565 B.n1030 B.n462 163.367
R1566 B.n1030 B.n460 163.367
R1567 B.n1034 B.n460 163.367
R1568 B.n1034 B.n454 163.367
R1569 B.n1042 B.n454 163.367
R1570 B.n1042 B.n452 163.367
R1571 B.n1046 B.n452 163.367
R1572 B.n1046 B.n446 163.367
R1573 B.n1054 B.n446 163.367
R1574 B.n1054 B.n444 163.367
R1575 B.n1058 B.n444 163.367
R1576 B.n1058 B.n438 163.367
R1577 B.n1066 B.n438 163.367
R1578 B.n1066 B.n436 163.367
R1579 B.n1070 B.n436 163.367
R1580 B.n1070 B.n430 163.367
R1581 B.n1078 B.n430 163.367
R1582 B.n1078 B.n428 163.367
R1583 B.n1082 B.n428 163.367
R1584 B.n1082 B.n422 163.367
R1585 B.n1091 B.n422 163.367
R1586 B.n1091 B.n420 163.367
R1587 B.n1095 B.n420 163.367
R1588 B.n1095 B.n3 163.367
R1589 B.n1380 B.n3 163.367
R1590 B.n1376 B.n2 163.367
R1591 B.n1376 B.n1375 163.367
R1592 B.n1375 B.n9 163.367
R1593 B.n1371 B.n9 163.367
R1594 B.n1371 B.n11 163.367
R1595 B.n1367 B.n11 163.367
R1596 B.n1367 B.n17 163.367
R1597 B.n1363 B.n17 163.367
R1598 B.n1363 B.n19 163.367
R1599 B.n1359 B.n19 163.367
R1600 B.n1359 B.n24 163.367
R1601 B.n1355 B.n24 163.367
R1602 B.n1355 B.n26 163.367
R1603 B.n1351 B.n26 163.367
R1604 B.n1351 B.n31 163.367
R1605 B.n1347 B.n31 163.367
R1606 B.n1347 B.n33 163.367
R1607 B.n1343 B.n33 163.367
R1608 B.n1343 B.n38 163.367
R1609 B.n1339 B.n38 163.367
R1610 B.n1339 B.n40 163.367
R1611 B.n1335 B.n40 163.367
R1612 B.n1335 B.n45 163.367
R1613 B.n1331 B.n45 163.367
R1614 B.n1331 B.n47 163.367
R1615 B.n1327 B.n47 163.367
R1616 B.n1327 B.n52 163.367
R1617 B.n1323 B.n52 163.367
R1618 B.n1323 B.n54 163.367
R1619 B.n1319 B.n54 163.367
R1620 B.n1319 B.n59 163.367
R1621 B.n1315 B.n59 163.367
R1622 B.n1315 B.n61 163.367
R1623 B.n1311 B.n61 163.367
R1624 B.n1311 B.n66 163.367
R1625 B.n1307 B.n66 163.367
R1626 B.n1307 B.n68 163.367
R1627 B.n1303 B.n68 163.367
R1628 B.n1303 B.n73 163.367
R1629 B.n1299 B.n73 163.367
R1630 B.n1299 B.n75 163.367
R1631 B.n1295 B.n75 163.367
R1632 B.n1295 B.n80 163.367
R1633 B.n1291 B.n80 163.367
R1634 B.n1291 B.n82 163.367
R1635 B.n1287 B.n82 163.367
R1636 B.n1287 B.n87 163.367
R1637 B.n1283 B.n87 163.367
R1638 B.n1283 B.n89 163.367
R1639 B.n1279 B.n89 163.367
R1640 B.n1279 B.n94 163.367
R1641 B.n1275 B.n94 163.367
R1642 B.n1275 B.n96 163.367
R1643 B.n1271 B.n96 163.367
R1644 B.n1271 B.n101 163.367
R1645 B.n1267 B.n101 163.367
R1646 B.n1267 B.n103 163.367
R1647 B.n1263 B.n103 163.367
R1648 B.n1263 B.n108 163.367
R1649 B.n1259 B.n108 163.367
R1650 B.n1259 B.n110 163.367
R1651 B.n1255 B.n110 163.367
R1652 B.n1255 B.n115 163.367
R1653 B.n1251 B.n115 163.367
R1654 B.n1251 B.n117 163.367
R1655 B.n1247 B.n117 163.367
R1656 B.n1247 B.n122 163.367
R1657 B.n1243 B.n122 163.367
R1658 B.n1243 B.n124 163.367
R1659 B.n1239 B.n124 163.367
R1660 B.n1239 B.n129 163.367
R1661 B.n1235 B.n129 163.367
R1662 B.n1235 B.n131 163.367
R1663 B.n1231 B.n131 163.367
R1664 B.n1231 B.n136 163.367
R1665 B.n1227 B.n136 163.367
R1666 B.n1227 B.n138 163.367
R1667 B.n1223 B.n138 163.367
R1668 B.n1223 B.n143 163.367
R1669 B.n1219 B.n143 163.367
R1670 B.n1219 B.n145 163.367
R1671 B.n1215 B.n145 163.367
R1672 B.n1215 B.n150 163.367
R1673 B.n206 B.t12 151.308
R1674 B.n638 B.t23 151.308
R1675 B.n209 B.t15 151.288
R1676 B.n636 B.t20 151.288
R1677 B.n210 B.n209 82.8126
R1678 B.n207 B.n206 82.8126
R1679 B.n639 B.n638 82.8126
R1680 B.n637 B.n636 82.8126
R1681 B.n1211 B.n1210 71.676
R1682 B.n212 B.n153 71.676
R1683 B.n216 B.n154 71.676
R1684 B.n220 B.n155 71.676
R1685 B.n224 B.n156 71.676
R1686 B.n228 B.n157 71.676
R1687 B.n232 B.n158 71.676
R1688 B.n236 B.n159 71.676
R1689 B.n240 B.n160 71.676
R1690 B.n244 B.n161 71.676
R1691 B.n248 B.n162 71.676
R1692 B.n252 B.n163 71.676
R1693 B.n256 B.n164 71.676
R1694 B.n260 B.n165 71.676
R1695 B.n264 B.n166 71.676
R1696 B.n268 B.n167 71.676
R1697 B.n272 B.n168 71.676
R1698 B.n276 B.n169 71.676
R1699 B.n280 B.n170 71.676
R1700 B.n284 B.n171 71.676
R1701 B.n288 B.n172 71.676
R1702 B.n292 B.n173 71.676
R1703 B.n296 B.n174 71.676
R1704 B.n300 B.n175 71.676
R1705 B.n304 B.n176 71.676
R1706 B.n308 B.n177 71.676
R1707 B.n312 B.n178 71.676
R1708 B.n316 B.n179 71.676
R1709 B.n320 B.n180 71.676
R1710 B.n324 B.n181 71.676
R1711 B.n328 B.n182 71.676
R1712 B.n332 B.n183 71.676
R1713 B.n336 B.n184 71.676
R1714 B.n340 B.n185 71.676
R1715 B.n344 B.n186 71.676
R1716 B.n348 B.n187 71.676
R1717 B.n352 B.n188 71.676
R1718 B.n356 B.n189 71.676
R1719 B.n360 B.n190 71.676
R1720 B.n364 B.n191 71.676
R1721 B.n368 B.n192 71.676
R1722 B.n372 B.n193 71.676
R1723 B.n376 B.n194 71.676
R1724 B.n380 B.n195 71.676
R1725 B.n384 B.n196 71.676
R1726 B.n388 B.n197 71.676
R1727 B.n392 B.n198 71.676
R1728 B.n396 B.n199 71.676
R1729 B.n400 B.n200 71.676
R1730 B.n404 B.n201 71.676
R1731 B.n408 B.n202 71.676
R1732 B.n412 B.n203 71.676
R1733 B.n1208 B.n204 71.676
R1734 B.n1208 B.n1207 71.676
R1735 B.n414 B.n203 71.676
R1736 B.n411 B.n202 71.676
R1737 B.n407 B.n201 71.676
R1738 B.n403 B.n200 71.676
R1739 B.n399 B.n199 71.676
R1740 B.n395 B.n198 71.676
R1741 B.n391 B.n197 71.676
R1742 B.n387 B.n196 71.676
R1743 B.n383 B.n195 71.676
R1744 B.n379 B.n194 71.676
R1745 B.n375 B.n193 71.676
R1746 B.n371 B.n192 71.676
R1747 B.n367 B.n191 71.676
R1748 B.n363 B.n190 71.676
R1749 B.n359 B.n189 71.676
R1750 B.n355 B.n188 71.676
R1751 B.n351 B.n187 71.676
R1752 B.n347 B.n186 71.676
R1753 B.n343 B.n185 71.676
R1754 B.n339 B.n184 71.676
R1755 B.n335 B.n183 71.676
R1756 B.n331 B.n182 71.676
R1757 B.n327 B.n181 71.676
R1758 B.n323 B.n180 71.676
R1759 B.n319 B.n179 71.676
R1760 B.n315 B.n178 71.676
R1761 B.n311 B.n177 71.676
R1762 B.n307 B.n176 71.676
R1763 B.n303 B.n175 71.676
R1764 B.n299 B.n174 71.676
R1765 B.n295 B.n173 71.676
R1766 B.n291 B.n172 71.676
R1767 B.n287 B.n171 71.676
R1768 B.n283 B.n170 71.676
R1769 B.n279 B.n169 71.676
R1770 B.n275 B.n168 71.676
R1771 B.n271 B.n167 71.676
R1772 B.n267 B.n166 71.676
R1773 B.n263 B.n165 71.676
R1774 B.n259 B.n164 71.676
R1775 B.n255 B.n163 71.676
R1776 B.n251 B.n162 71.676
R1777 B.n247 B.n161 71.676
R1778 B.n243 B.n160 71.676
R1779 B.n239 B.n159 71.676
R1780 B.n235 B.n158 71.676
R1781 B.n231 B.n157 71.676
R1782 B.n227 B.n156 71.676
R1783 B.n223 B.n155 71.676
R1784 B.n219 B.n154 71.676
R1785 B.n215 B.n153 71.676
R1786 B.n1210 B.n152 71.676
R1787 B.n850 B.n849 71.676
R1788 B.n635 B.n583 71.676
R1789 B.n842 B.n584 71.676
R1790 B.n838 B.n585 71.676
R1791 B.n834 B.n586 71.676
R1792 B.n830 B.n587 71.676
R1793 B.n826 B.n588 71.676
R1794 B.n822 B.n589 71.676
R1795 B.n818 B.n590 71.676
R1796 B.n814 B.n591 71.676
R1797 B.n810 B.n592 71.676
R1798 B.n806 B.n593 71.676
R1799 B.n802 B.n594 71.676
R1800 B.n798 B.n595 71.676
R1801 B.n794 B.n596 71.676
R1802 B.n790 B.n597 71.676
R1803 B.n786 B.n598 71.676
R1804 B.n782 B.n599 71.676
R1805 B.n778 B.n600 71.676
R1806 B.n774 B.n601 71.676
R1807 B.n770 B.n602 71.676
R1808 B.n766 B.n603 71.676
R1809 B.n762 B.n604 71.676
R1810 B.n758 B.n605 71.676
R1811 B.n753 B.n606 71.676
R1812 B.n749 B.n607 71.676
R1813 B.n745 B.n608 71.676
R1814 B.n741 B.n609 71.676
R1815 B.n737 B.n610 71.676
R1816 B.n732 B.n611 71.676
R1817 B.n728 B.n612 71.676
R1818 B.n724 B.n613 71.676
R1819 B.n720 B.n614 71.676
R1820 B.n716 B.n615 71.676
R1821 B.n712 B.n616 71.676
R1822 B.n708 B.n617 71.676
R1823 B.n704 B.n618 71.676
R1824 B.n700 B.n619 71.676
R1825 B.n696 B.n620 71.676
R1826 B.n692 B.n621 71.676
R1827 B.n688 B.n622 71.676
R1828 B.n684 B.n623 71.676
R1829 B.n680 B.n624 71.676
R1830 B.n676 B.n625 71.676
R1831 B.n672 B.n626 71.676
R1832 B.n668 B.n627 71.676
R1833 B.n664 B.n628 71.676
R1834 B.n660 B.n629 71.676
R1835 B.n656 B.n630 71.676
R1836 B.n652 B.n631 71.676
R1837 B.n648 B.n632 71.676
R1838 B.n644 B.n633 71.676
R1839 B.n849 B.n582 71.676
R1840 B.n843 B.n583 71.676
R1841 B.n839 B.n584 71.676
R1842 B.n835 B.n585 71.676
R1843 B.n831 B.n586 71.676
R1844 B.n827 B.n587 71.676
R1845 B.n823 B.n588 71.676
R1846 B.n819 B.n589 71.676
R1847 B.n815 B.n590 71.676
R1848 B.n811 B.n591 71.676
R1849 B.n807 B.n592 71.676
R1850 B.n803 B.n593 71.676
R1851 B.n799 B.n594 71.676
R1852 B.n795 B.n595 71.676
R1853 B.n791 B.n596 71.676
R1854 B.n787 B.n597 71.676
R1855 B.n783 B.n598 71.676
R1856 B.n779 B.n599 71.676
R1857 B.n775 B.n600 71.676
R1858 B.n771 B.n601 71.676
R1859 B.n767 B.n602 71.676
R1860 B.n763 B.n603 71.676
R1861 B.n759 B.n604 71.676
R1862 B.n754 B.n605 71.676
R1863 B.n750 B.n606 71.676
R1864 B.n746 B.n607 71.676
R1865 B.n742 B.n608 71.676
R1866 B.n738 B.n609 71.676
R1867 B.n733 B.n610 71.676
R1868 B.n729 B.n611 71.676
R1869 B.n725 B.n612 71.676
R1870 B.n721 B.n613 71.676
R1871 B.n717 B.n614 71.676
R1872 B.n713 B.n615 71.676
R1873 B.n709 B.n616 71.676
R1874 B.n705 B.n617 71.676
R1875 B.n701 B.n618 71.676
R1876 B.n697 B.n619 71.676
R1877 B.n693 B.n620 71.676
R1878 B.n689 B.n621 71.676
R1879 B.n685 B.n622 71.676
R1880 B.n681 B.n623 71.676
R1881 B.n677 B.n624 71.676
R1882 B.n673 B.n625 71.676
R1883 B.n669 B.n626 71.676
R1884 B.n665 B.n627 71.676
R1885 B.n661 B.n628 71.676
R1886 B.n657 B.n629 71.676
R1887 B.n653 B.n630 71.676
R1888 B.n649 B.n631 71.676
R1889 B.n645 B.n632 71.676
R1890 B.n641 B.n633 71.676
R1891 B.n1381 B.n1380 71.676
R1892 B.n1381 B.n2 71.676
R1893 B.n207 B.t13 68.4948
R1894 B.n639 B.t22 68.4948
R1895 B.n210 B.t16 68.4761
R1896 B.n637 B.t19 68.4761
R1897 B.n848 B.n579 67.8913
R1898 B.n1209 B.n149 67.8913
R1899 B.n211 B.n210 59.5399
R1900 B.n208 B.n207 59.5399
R1901 B.n735 B.n639 59.5399
R1902 B.n756 B.n637 59.5399
R1903 B.n855 B.n579 38.154
R1904 B.n855 B.n575 38.154
R1905 B.n861 B.n575 38.154
R1906 B.n861 B.n571 38.154
R1907 B.n867 B.n571 38.154
R1908 B.n867 B.n567 38.154
R1909 B.n873 B.n567 38.154
R1910 B.n873 B.n563 38.154
R1911 B.n879 B.n563 38.154
R1912 B.n885 B.n559 38.154
R1913 B.n885 B.n555 38.154
R1914 B.n891 B.n555 38.154
R1915 B.n891 B.n551 38.154
R1916 B.n897 B.n551 38.154
R1917 B.n897 B.n547 38.154
R1918 B.n903 B.n547 38.154
R1919 B.n903 B.n543 38.154
R1920 B.n909 B.n543 38.154
R1921 B.n909 B.n539 38.154
R1922 B.n915 B.n539 38.154
R1923 B.n915 B.n535 38.154
R1924 B.n921 B.n535 38.154
R1925 B.n921 B.n531 38.154
R1926 B.n927 B.n531 38.154
R1927 B.n933 B.n527 38.154
R1928 B.n933 B.n523 38.154
R1929 B.n939 B.n523 38.154
R1930 B.n939 B.n519 38.154
R1931 B.n945 B.n519 38.154
R1932 B.n945 B.n515 38.154
R1933 B.n951 B.n515 38.154
R1934 B.n951 B.n511 38.154
R1935 B.n957 B.n511 38.154
R1936 B.n957 B.n507 38.154
R1937 B.n963 B.n507 38.154
R1938 B.n969 B.n503 38.154
R1939 B.n969 B.n499 38.154
R1940 B.n975 B.n499 38.154
R1941 B.n975 B.n495 38.154
R1942 B.n981 B.n495 38.154
R1943 B.n981 B.n491 38.154
R1944 B.n987 B.n491 38.154
R1945 B.n987 B.n487 38.154
R1946 B.n993 B.n487 38.154
R1947 B.n993 B.n482 38.154
R1948 B.n999 B.n482 38.154
R1949 B.n999 B.n483 38.154
R1950 B.n1005 B.n475 38.154
R1951 B.n1011 B.n475 38.154
R1952 B.n1011 B.n471 38.154
R1953 B.n1017 B.n471 38.154
R1954 B.n1017 B.n467 38.154
R1955 B.n1023 B.n467 38.154
R1956 B.n1023 B.n463 38.154
R1957 B.n1029 B.n463 38.154
R1958 B.n1029 B.n459 38.154
R1959 B.n1035 B.n459 38.154
R1960 B.n1035 B.n455 38.154
R1961 B.n1041 B.n455 38.154
R1962 B.n1047 B.n451 38.154
R1963 B.n1047 B.n447 38.154
R1964 B.n1053 B.n447 38.154
R1965 B.n1053 B.n443 38.154
R1966 B.n1059 B.n443 38.154
R1967 B.n1059 B.n439 38.154
R1968 B.n1065 B.n439 38.154
R1969 B.n1065 B.n435 38.154
R1970 B.n1071 B.n435 38.154
R1971 B.n1071 B.n431 38.154
R1972 B.n1077 B.n431 38.154
R1973 B.n1083 B.n427 38.154
R1974 B.n1083 B.n423 38.154
R1975 B.n1090 B.n423 38.154
R1976 B.n1090 B.n419 38.154
R1977 B.n1096 B.n419 38.154
R1978 B.n1096 B.n4 38.154
R1979 B.n1379 B.n4 38.154
R1980 B.n1379 B.n1378 38.154
R1981 B.n1378 B.n1377 38.154
R1982 B.n1377 B.n8 38.154
R1983 B.n12 B.n8 38.154
R1984 B.n1370 B.n12 38.154
R1985 B.n1370 B.n1369 38.154
R1986 B.n1369 B.n1368 38.154
R1987 B.n1368 B.n16 38.154
R1988 B.n1362 B.n1361 38.154
R1989 B.n1361 B.n1360 38.154
R1990 B.n1360 B.n23 38.154
R1991 B.n1354 B.n23 38.154
R1992 B.n1354 B.n1353 38.154
R1993 B.n1353 B.n1352 38.154
R1994 B.n1352 B.n30 38.154
R1995 B.n1346 B.n30 38.154
R1996 B.n1346 B.n1345 38.154
R1997 B.n1345 B.n1344 38.154
R1998 B.n1344 B.n37 38.154
R1999 B.n1338 B.n1337 38.154
R2000 B.n1337 B.n1336 38.154
R2001 B.n1336 B.n44 38.154
R2002 B.n1330 B.n44 38.154
R2003 B.n1330 B.n1329 38.154
R2004 B.n1329 B.n1328 38.154
R2005 B.n1328 B.n51 38.154
R2006 B.n1322 B.n51 38.154
R2007 B.n1322 B.n1321 38.154
R2008 B.n1321 B.n1320 38.154
R2009 B.n1320 B.n58 38.154
R2010 B.n1314 B.n58 38.154
R2011 B.n1313 B.n1312 38.154
R2012 B.n1312 B.n65 38.154
R2013 B.n1306 B.n65 38.154
R2014 B.n1306 B.n1305 38.154
R2015 B.n1305 B.n1304 38.154
R2016 B.n1304 B.n72 38.154
R2017 B.n1298 B.n72 38.154
R2018 B.n1298 B.n1297 38.154
R2019 B.n1297 B.n1296 38.154
R2020 B.n1296 B.n79 38.154
R2021 B.n1290 B.n79 38.154
R2022 B.n1290 B.n1289 38.154
R2023 B.n1288 B.n86 38.154
R2024 B.n1282 B.n86 38.154
R2025 B.n1282 B.n1281 38.154
R2026 B.n1281 B.n1280 38.154
R2027 B.n1280 B.n93 38.154
R2028 B.n1274 B.n93 38.154
R2029 B.n1274 B.n1273 38.154
R2030 B.n1273 B.n1272 38.154
R2031 B.n1272 B.n100 38.154
R2032 B.n1266 B.n100 38.154
R2033 B.n1266 B.n1265 38.154
R2034 B.n1264 B.n107 38.154
R2035 B.n1258 B.n107 38.154
R2036 B.n1258 B.n1257 38.154
R2037 B.n1257 B.n1256 38.154
R2038 B.n1256 B.n114 38.154
R2039 B.n1250 B.n114 38.154
R2040 B.n1250 B.n1249 38.154
R2041 B.n1249 B.n1248 38.154
R2042 B.n1248 B.n121 38.154
R2043 B.n1242 B.n121 38.154
R2044 B.n1242 B.n1241 38.154
R2045 B.n1241 B.n1240 38.154
R2046 B.n1240 B.n128 38.154
R2047 B.n1234 B.n128 38.154
R2048 B.n1234 B.n1233 38.154
R2049 B.n1232 B.n135 38.154
R2050 B.n1226 B.n135 38.154
R2051 B.n1226 B.n1225 38.154
R2052 B.n1225 B.n1224 38.154
R2053 B.n1224 B.n142 38.154
R2054 B.n1218 B.n142 38.154
R2055 B.n1218 B.n1217 38.154
R2056 B.n1217 B.n1216 38.154
R2057 B.n1216 B.n149 38.154
R2058 B.n963 B.t9 35.9097
R2059 B.t8 B.n451 35.9097
R2060 B.t4 B.n37 35.9097
R2061 B.t7 B.n1288 35.9097
R2062 B.n852 B.n851 34.8103
R2063 B.n640 B.n577 34.8103
R2064 B.n1206 B.n1205 34.8103
R2065 B.n1213 B.n1212 34.8103
R2066 B.n879 B.t18 23.5659
R2067 B.t2 B.n527 23.5659
R2068 B.n1077 B.t5 23.5659
R2069 B.n1362 B.t1 23.5659
R2070 B.n1265 B.t6 23.5659
R2071 B.t11 B.n1232 23.5659
R2072 B.n483 B.t0 19.0773
R2073 B.n1005 B.t0 19.0773
R2074 B.n1314 B.t3 19.0773
R2075 B.t3 B.n1313 19.0773
R2076 B B.n1382 18.0485
R2077 B.t18 B.n559 14.5886
R2078 B.n927 B.t2 14.5886
R2079 B.t5 B.n427 14.5886
R2080 B.t1 B.n16 14.5886
R2081 B.t6 B.n1264 14.5886
R2082 B.n1233 B.t11 14.5886
R2083 B.n853 B.n852 10.6151
R2084 B.n853 B.n573 10.6151
R2085 B.n863 B.n573 10.6151
R2086 B.n864 B.n863 10.6151
R2087 B.n865 B.n864 10.6151
R2088 B.n865 B.n565 10.6151
R2089 B.n875 B.n565 10.6151
R2090 B.n876 B.n875 10.6151
R2091 B.n877 B.n876 10.6151
R2092 B.n877 B.n557 10.6151
R2093 B.n887 B.n557 10.6151
R2094 B.n888 B.n887 10.6151
R2095 B.n889 B.n888 10.6151
R2096 B.n889 B.n549 10.6151
R2097 B.n899 B.n549 10.6151
R2098 B.n900 B.n899 10.6151
R2099 B.n901 B.n900 10.6151
R2100 B.n901 B.n541 10.6151
R2101 B.n911 B.n541 10.6151
R2102 B.n912 B.n911 10.6151
R2103 B.n913 B.n912 10.6151
R2104 B.n913 B.n533 10.6151
R2105 B.n923 B.n533 10.6151
R2106 B.n924 B.n923 10.6151
R2107 B.n925 B.n924 10.6151
R2108 B.n925 B.n525 10.6151
R2109 B.n935 B.n525 10.6151
R2110 B.n936 B.n935 10.6151
R2111 B.n937 B.n936 10.6151
R2112 B.n937 B.n517 10.6151
R2113 B.n947 B.n517 10.6151
R2114 B.n948 B.n947 10.6151
R2115 B.n949 B.n948 10.6151
R2116 B.n949 B.n509 10.6151
R2117 B.n959 B.n509 10.6151
R2118 B.n960 B.n959 10.6151
R2119 B.n961 B.n960 10.6151
R2120 B.n961 B.n501 10.6151
R2121 B.n971 B.n501 10.6151
R2122 B.n972 B.n971 10.6151
R2123 B.n973 B.n972 10.6151
R2124 B.n973 B.n493 10.6151
R2125 B.n983 B.n493 10.6151
R2126 B.n984 B.n983 10.6151
R2127 B.n985 B.n984 10.6151
R2128 B.n985 B.n485 10.6151
R2129 B.n995 B.n485 10.6151
R2130 B.n996 B.n995 10.6151
R2131 B.n997 B.n996 10.6151
R2132 B.n997 B.n477 10.6151
R2133 B.n1007 B.n477 10.6151
R2134 B.n1008 B.n1007 10.6151
R2135 B.n1009 B.n1008 10.6151
R2136 B.n1009 B.n469 10.6151
R2137 B.n1019 B.n469 10.6151
R2138 B.n1020 B.n1019 10.6151
R2139 B.n1021 B.n1020 10.6151
R2140 B.n1021 B.n461 10.6151
R2141 B.n1031 B.n461 10.6151
R2142 B.n1032 B.n1031 10.6151
R2143 B.n1033 B.n1032 10.6151
R2144 B.n1033 B.n453 10.6151
R2145 B.n1043 B.n453 10.6151
R2146 B.n1044 B.n1043 10.6151
R2147 B.n1045 B.n1044 10.6151
R2148 B.n1045 B.n445 10.6151
R2149 B.n1055 B.n445 10.6151
R2150 B.n1056 B.n1055 10.6151
R2151 B.n1057 B.n1056 10.6151
R2152 B.n1057 B.n437 10.6151
R2153 B.n1067 B.n437 10.6151
R2154 B.n1068 B.n1067 10.6151
R2155 B.n1069 B.n1068 10.6151
R2156 B.n1069 B.n429 10.6151
R2157 B.n1079 B.n429 10.6151
R2158 B.n1080 B.n1079 10.6151
R2159 B.n1081 B.n1080 10.6151
R2160 B.n1081 B.n421 10.6151
R2161 B.n1092 B.n421 10.6151
R2162 B.n1093 B.n1092 10.6151
R2163 B.n1094 B.n1093 10.6151
R2164 B.n1094 B.n0 10.6151
R2165 B.n851 B.n581 10.6151
R2166 B.n846 B.n581 10.6151
R2167 B.n846 B.n845 10.6151
R2168 B.n845 B.n844 10.6151
R2169 B.n844 B.n841 10.6151
R2170 B.n841 B.n840 10.6151
R2171 B.n840 B.n837 10.6151
R2172 B.n837 B.n836 10.6151
R2173 B.n836 B.n833 10.6151
R2174 B.n833 B.n832 10.6151
R2175 B.n832 B.n829 10.6151
R2176 B.n829 B.n828 10.6151
R2177 B.n828 B.n825 10.6151
R2178 B.n825 B.n824 10.6151
R2179 B.n824 B.n821 10.6151
R2180 B.n821 B.n820 10.6151
R2181 B.n820 B.n817 10.6151
R2182 B.n817 B.n816 10.6151
R2183 B.n816 B.n813 10.6151
R2184 B.n813 B.n812 10.6151
R2185 B.n812 B.n809 10.6151
R2186 B.n809 B.n808 10.6151
R2187 B.n808 B.n805 10.6151
R2188 B.n805 B.n804 10.6151
R2189 B.n804 B.n801 10.6151
R2190 B.n801 B.n800 10.6151
R2191 B.n800 B.n797 10.6151
R2192 B.n797 B.n796 10.6151
R2193 B.n796 B.n793 10.6151
R2194 B.n793 B.n792 10.6151
R2195 B.n792 B.n789 10.6151
R2196 B.n789 B.n788 10.6151
R2197 B.n788 B.n785 10.6151
R2198 B.n785 B.n784 10.6151
R2199 B.n784 B.n781 10.6151
R2200 B.n781 B.n780 10.6151
R2201 B.n780 B.n777 10.6151
R2202 B.n777 B.n776 10.6151
R2203 B.n776 B.n773 10.6151
R2204 B.n773 B.n772 10.6151
R2205 B.n772 B.n769 10.6151
R2206 B.n769 B.n768 10.6151
R2207 B.n768 B.n765 10.6151
R2208 B.n765 B.n764 10.6151
R2209 B.n764 B.n761 10.6151
R2210 B.n761 B.n760 10.6151
R2211 B.n760 B.n757 10.6151
R2212 B.n755 B.n752 10.6151
R2213 B.n752 B.n751 10.6151
R2214 B.n751 B.n748 10.6151
R2215 B.n748 B.n747 10.6151
R2216 B.n747 B.n744 10.6151
R2217 B.n744 B.n743 10.6151
R2218 B.n743 B.n740 10.6151
R2219 B.n740 B.n739 10.6151
R2220 B.n739 B.n736 10.6151
R2221 B.n734 B.n731 10.6151
R2222 B.n731 B.n730 10.6151
R2223 B.n730 B.n727 10.6151
R2224 B.n727 B.n726 10.6151
R2225 B.n726 B.n723 10.6151
R2226 B.n723 B.n722 10.6151
R2227 B.n722 B.n719 10.6151
R2228 B.n719 B.n718 10.6151
R2229 B.n718 B.n715 10.6151
R2230 B.n715 B.n714 10.6151
R2231 B.n714 B.n711 10.6151
R2232 B.n711 B.n710 10.6151
R2233 B.n710 B.n707 10.6151
R2234 B.n707 B.n706 10.6151
R2235 B.n706 B.n703 10.6151
R2236 B.n703 B.n702 10.6151
R2237 B.n702 B.n699 10.6151
R2238 B.n699 B.n698 10.6151
R2239 B.n698 B.n695 10.6151
R2240 B.n695 B.n694 10.6151
R2241 B.n694 B.n691 10.6151
R2242 B.n691 B.n690 10.6151
R2243 B.n690 B.n687 10.6151
R2244 B.n687 B.n686 10.6151
R2245 B.n686 B.n683 10.6151
R2246 B.n683 B.n682 10.6151
R2247 B.n682 B.n679 10.6151
R2248 B.n679 B.n678 10.6151
R2249 B.n678 B.n675 10.6151
R2250 B.n675 B.n674 10.6151
R2251 B.n674 B.n671 10.6151
R2252 B.n671 B.n670 10.6151
R2253 B.n670 B.n667 10.6151
R2254 B.n667 B.n666 10.6151
R2255 B.n666 B.n663 10.6151
R2256 B.n663 B.n662 10.6151
R2257 B.n662 B.n659 10.6151
R2258 B.n659 B.n658 10.6151
R2259 B.n658 B.n655 10.6151
R2260 B.n655 B.n654 10.6151
R2261 B.n654 B.n651 10.6151
R2262 B.n651 B.n650 10.6151
R2263 B.n650 B.n647 10.6151
R2264 B.n647 B.n646 10.6151
R2265 B.n646 B.n643 10.6151
R2266 B.n643 B.n642 10.6151
R2267 B.n642 B.n640 10.6151
R2268 B.n857 B.n577 10.6151
R2269 B.n858 B.n857 10.6151
R2270 B.n859 B.n858 10.6151
R2271 B.n859 B.n569 10.6151
R2272 B.n869 B.n569 10.6151
R2273 B.n870 B.n869 10.6151
R2274 B.n871 B.n870 10.6151
R2275 B.n871 B.n561 10.6151
R2276 B.n881 B.n561 10.6151
R2277 B.n882 B.n881 10.6151
R2278 B.n883 B.n882 10.6151
R2279 B.n883 B.n553 10.6151
R2280 B.n893 B.n553 10.6151
R2281 B.n894 B.n893 10.6151
R2282 B.n895 B.n894 10.6151
R2283 B.n895 B.n545 10.6151
R2284 B.n905 B.n545 10.6151
R2285 B.n906 B.n905 10.6151
R2286 B.n907 B.n906 10.6151
R2287 B.n907 B.n537 10.6151
R2288 B.n917 B.n537 10.6151
R2289 B.n918 B.n917 10.6151
R2290 B.n919 B.n918 10.6151
R2291 B.n919 B.n529 10.6151
R2292 B.n929 B.n529 10.6151
R2293 B.n930 B.n929 10.6151
R2294 B.n931 B.n930 10.6151
R2295 B.n931 B.n521 10.6151
R2296 B.n941 B.n521 10.6151
R2297 B.n942 B.n941 10.6151
R2298 B.n943 B.n942 10.6151
R2299 B.n943 B.n513 10.6151
R2300 B.n953 B.n513 10.6151
R2301 B.n954 B.n953 10.6151
R2302 B.n955 B.n954 10.6151
R2303 B.n955 B.n505 10.6151
R2304 B.n965 B.n505 10.6151
R2305 B.n966 B.n965 10.6151
R2306 B.n967 B.n966 10.6151
R2307 B.n967 B.n497 10.6151
R2308 B.n977 B.n497 10.6151
R2309 B.n978 B.n977 10.6151
R2310 B.n979 B.n978 10.6151
R2311 B.n979 B.n489 10.6151
R2312 B.n989 B.n489 10.6151
R2313 B.n990 B.n989 10.6151
R2314 B.n991 B.n990 10.6151
R2315 B.n991 B.n480 10.6151
R2316 B.n1001 B.n480 10.6151
R2317 B.n1002 B.n1001 10.6151
R2318 B.n1003 B.n1002 10.6151
R2319 B.n1003 B.n473 10.6151
R2320 B.n1013 B.n473 10.6151
R2321 B.n1014 B.n1013 10.6151
R2322 B.n1015 B.n1014 10.6151
R2323 B.n1015 B.n465 10.6151
R2324 B.n1025 B.n465 10.6151
R2325 B.n1026 B.n1025 10.6151
R2326 B.n1027 B.n1026 10.6151
R2327 B.n1027 B.n457 10.6151
R2328 B.n1037 B.n457 10.6151
R2329 B.n1038 B.n1037 10.6151
R2330 B.n1039 B.n1038 10.6151
R2331 B.n1039 B.n449 10.6151
R2332 B.n1049 B.n449 10.6151
R2333 B.n1050 B.n1049 10.6151
R2334 B.n1051 B.n1050 10.6151
R2335 B.n1051 B.n441 10.6151
R2336 B.n1061 B.n441 10.6151
R2337 B.n1062 B.n1061 10.6151
R2338 B.n1063 B.n1062 10.6151
R2339 B.n1063 B.n433 10.6151
R2340 B.n1073 B.n433 10.6151
R2341 B.n1074 B.n1073 10.6151
R2342 B.n1075 B.n1074 10.6151
R2343 B.n1075 B.n425 10.6151
R2344 B.n1085 B.n425 10.6151
R2345 B.n1086 B.n1085 10.6151
R2346 B.n1088 B.n1086 10.6151
R2347 B.n1088 B.n1087 10.6151
R2348 B.n1087 B.n417 10.6151
R2349 B.n1099 B.n417 10.6151
R2350 B.n1100 B.n1099 10.6151
R2351 B.n1101 B.n1100 10.6151
R2352 B.n1102 B.n1101 10.6151
R2353 B.n1103 B.n1102 10.6151
R2354 B.n1106 B.n1103 10.6151
R2355 B.n1107 B.n1106 10.6151
R2356 B.n1108 B.n1107 10.6151
R2357 B.n1109 B.n1108 10.6151
R2358 B.n1111 B.n1109 10.6151
R2359 B.n1112 B.n1111 10.6151
R2360 B.n1113 B.n1112 10.6151
R2361 B.n1114 B.n1113 10.6151
R2362 B.n1116 B.n1114 10.6151
R2363 B.n1117 B.n1116 10.6151
R2364 B.n1118 B.n1117 10.6151
R2365 B.n1119 B.n1118 10.6151
R2366 B.n1121 B.n1119 10.6151
R2367 B.n1122 B.n1121 10.6151
R2368 B.n1123 B.n1122 10.6151
R2369 B.n1124 B.n1123 10.6151
R2370 B.n1126 B.n1124 10.6151
R2371 B.n1127 B.n1126 10.6151
R2372 B.n1128 B.n1127 10.6151
R2373 B.n1129 B.n1128 10.6151
R2374 B.n1131 B.n1129 10.6151
R2375 B.n1132 B.n1131 10.6151
R2376 B.n1133 B.n1132 10.6151
R2377 B.n1134 B.n1133 10.6151
R2378 B.n1136 B.n1134 10.6151
R2379 B.n1137 B.n1136 10.6151
R2380 B.n1138 B.n1137 10.6151
R2381 B.n1139 B.n1138 10.6151
R2382 B.n1141 B.n1139 10.6151
R2383 B.n1142 B.n1141 10.6151
R2384 B.n1143 B.n1142 10.6151
R2385 B.n1144 B.n1143 10.6151
R2386 B.n1146 B.n1144 10.6151
R2387 B.n1147 B.n1146 10.6151
R2388 B.n1148 B.n1147 10.6151
R2389 B.n1149 B.n1148 10.6151
R2390 B.n1151 B.n1149 10.6151
R2391 B.n1152 B.n1151 10.6151
R2392 B.n1153 B.n1152 10.6151
R2393 B.n1154 B.n1153 10.6151
R2394 B.n1156 B.n1154 10.6151
R2395 B.n1157 B.n1156 10.6151
R2396 B.n1158 B.n1157 10.6151
R2397 B.n1159 B.n1158 10.6151
R2398 B.n1161 B.n1159 10.6151
R2399 B.n1162 B.n1161 10.6151
R2400 B.n1163 B.n1162 10.6151
R2401 B.n1164 B.n1163 10.6151
R2402 B.n1166 B.n1164 10.6151
R2403 B.n1167 B.n1166 10.6151
R2404 B.n1168 B.n1167 10.6151
R2405 B.n1169 B.n1168 10.6151
R2406 B.n1171 B.n1169 10.6151
R2407 B.n1172 B.n1171 10.6151
R2408 B.n1173 B.n1172 10.6151
R2409 B.n1174 B.n1173 10.6151
R2410 B.n1176 B.n1174 10.6151
R2411 B.n1177 B.n1176 10.6151
R2412 B.n1178 B.n1177 10.6151
R2413 B.n1179 B.n1178 10.6151
R2414 B.n1181 B.n1179 10.6151
R2415 B.n1182 B.n1181 10.6151
R2416 B.n1183 B.n1182 10.6151
R2417 B.n1184 B.n1183 10.6151
R2418 B.n1186 B.n1184 10.6151
R2419 B.n1187 B.n1186 10.6151
R2420 B.n1188 B.n1187 10.6151
R2421 B.n1189 B.n1188 10.6151
R2422 B.n1191 B.n1189 10.6151
R2423 B.n1192 B.n1191 10.6151
R2424 B.n1193 B.n1192 10.6151
R2425 B.n1194 B.n1193 10.6151
R2426 B.n1196 B.n1194 10.6151
R2427 B.n1197 B.n1196 10.6151
R2428 B.n1198 B.n1197 10.6151
R2429 B.n1199 B.n1198 10.6151
R2430 B.n1201 B.n1199 10.6151
R2431 B.n1202 B.n1201 10.6151
R2432 B.n1203 B.n1202 10.6151
R2433 B.n1204 B.n1203 10.6151
R2434 B.n1205 B.n1204 10.6151
R2435 B.n1374 B.n1 10.6151
R2436 B.n1374 B.n1373 10.6151
R2437 B.n1373 B.n1372 10.6151
R2438 B.n1372 B.n10 10.6151
R2439 B.n1366 B.n10 10.6151
R2440 B.n1366 B.n1365 10.6151
R2441 B.n1365 B.n1364 10.6151
R2442 B.n1364 B.n18 10.6151
R2443 B.n1358 B.n18 10.6151
R2444 B.n1358 B.n1357 10.6151
R2445 B.n1357 B.n1356 10.6151
R2446 B.n1356 B.n25 10.6151
R2447 B.n1350 B.n25 10.6151
R2448 B.n1350 B.n1349 10.6151
R2449 B.n1349 B.n1348 10.6151
R2450 B.n1348 B.n32 10.6151
R2451 B.n1342 B.n32 10.6151
R2452 B.n1342 B.n1341 10.6151
R2453 B.n1341 B.n1340 10.6151
R2454 B.n1340 B.n39 10.6151
R2455 B.n1334 B.n39 10.6151
R2456 B.n1334 B.n1333 10.6151
R2457 B.n1333 B.n1332 10.6151
R2458 B.n1332 B.n46 10.6151
R2459 B.n1326 B.n46 10.6151
R2460 B.n1326 B.n1325 10.6151
R2461 B.n1325 B.n1324 10.6151
R2462 B.n1324 B.n53 10.6151
R2463 B.n1318 B.n53 10.6151
R2464 B.n1318 B.n1317 10.6151
R2465 B.n1317 B.n1316 10.6151
R2466 B.n1316 B.n60 10.6151
R2467 B.n1310 B.n60 10.6151
R2468 B.n1310 B.n1309 10.6151
R2469 B.n1309 B.n1308 10.6151
R2470 B.n1308 B.n67 10.6151
R2471 B.n1302 B.n67 10.6151
R2472 B.n1302 B.n1301 10.6151
R2473 B.n1301 B.n1300 10.6151
R2474 B.n1300 B.n74 10.6151
R2475 B.n1294 B.n74 10.6151
R2476 B.n1294 B.n1293 10.6151
R2477 B.n1293 B.n1292 10.6151
R2478 B.n1292 B.n81 10.6151
R2479 B.n1286 B.n81 10.6151
R2480 B.n1286 B.n1285 10.6151
R2481 B.n1285 B.n1284 10.6151
R2482 B.n1284 B.n88 10.6151
R2483 B.n1278 B.n88 10.6151
R2484 B.n1278 B.n1277 10.6151
R2485 B.n1277 B.n1276 10.6151
R2486 B.n1276 B.n95 10.6151
R2487 B.n1270 B.n95 10.6151
R2488 B.n1270 B.n1269 10.6151
R2489 B.n1269 B.n1268 10.6151
R2490 B.n1268 B.n102 10.6151
R2491 B.n1262 B.n102 10.6151
R2492 B.n1262 B.n1261 10.6151
R2493 B.n1261 B.n1260 10.6151
R2494 B.n1260 B.n109 10.6151
R2495 B.n1254 B.n109 10.6151
R2496 B.n1254 B.n1253 10.6151
R2497 B.n1253 B.n1252 10.6151
R2498 B.n1252 B.n116 10.6151
R2499 B.n1246 B.n116 10.6151
R2500 B.n1246 B.n1245 10.6151
R2501 B.n1245 B.n1244 10.6151
R2502 B.n1244 B.n123 10.6151
R2503 B.n1238 B.n123 10.6151
R2504 B.n1238 B.n1237 10.6151
R2505 B.n1237 B.n1236 10.6151
R2506 B.n1236 B.n130 10.6151
R2507 B.n1230 B.n130 10.6151
R2508 B.n1230 B.n1229 10.6151
R2509 B.n1229 B.n1228 10.6151
R2510 B.n1228 B.n137 10.6151
R2511 B.n1222 B.n137 10.6151
R2512 B.n1222 B.n1221 10.6151
R2513 B.n1221 B.n1220 10.6151
R2514 B.n1220 B.n144 10.6151
R2515 B.n1214 B.n144 10.6151
R2516 B.n1214 B.n1213 10.6151
R2517 B.n1212 B.n151 10.6151
R2518 B.n213 B.n151 10.6151
R2519 B.n214 B.n213 10.6151
R2520 B.n217 B.n214 10.6151
R2521 B.n218 B.n217 10.6151
R2522 B.n221 B.n218 10.6151
R2523 B.n222 B.n221 10.6151
R2524 B.n225 B.n222 10.6151
R2525 B.n226 B.n225 10.6151
R2526 B.n229 B.n226 10.6151
R2527 B.n230 B.n229 10.6151
R2528 B.n233 B.n230 10.6151
R2529 B.n234 B.n233 10.6151
R2530 B.n237 B.n234 10.6151
R2531 B.n238 B.n237 10.6151
R2532 B.n241 B.n238 10.6151
R2533 B.n242 B.n241 10.6151
R2534 B.n245 B.n242 10.6151
R2535 B.n246 B.n245 10.6151
R2536 B.n249 B.n246 10.6151
R2537 B.n250 B.n249 10.6151
R2538 B.n253 B.n250 10.6151
R2539 B.n254 B.n253 10.6151
R2540 B.n257 B.n254 10.6151
R2541 B.n258 B.n257 10.6151
R2542 B.n261 B.n258 10.6151
R2543 B.n262 B.n261 10.6151
R2544 B.n265 B.n262 10.6151
R2545 B.n266 B.n265 10.6151
R2546 B.n269 B.n266 10.6151
R2547 B.n270 B.n269 10.6151
R2548 B.n273 B.n270 10.6151
R2549 B.n274 B.n273 10.6151
R2550 B.n277 B.n274 10.6151
R2551 B.n278 B.n277 10.6151
R2552 B.n281 B.n278 10.6151
R2553 B.n282 B.n281 10.6151
R2554 B.n285 B.n282 10.6151
R2555 B.n286 B.n285 10.6151
R2556 B.n289 B.n286 10.6151
R2557 B.n290 B.n289 10.6151
R2558 B.n293 B.n290 10.6151
R2559 B.n294 B.n293 10.6151
R2560 B.n297 B.n294 10.6151
R2561 B.n298 B.n297 10.6151
R2562 B.n301 B.n298 10.6151
R2563 B.n302 B.n301 10.6151
R2564 B.n306 B.n305 10.6151
R2565 B.n309 B.n306 10.6151
R2566 B.n310 B.n309 10.6151
R2567 B.n313 B.n310 10.6151
R2568 B.n314 B.n313 10.6151
R2569 B.n317 B.n314 10.6151
R2570 B.n318 B.n317 10.6151
R2571 B.n321 B.n318 10.6151
R2572 B.n322 B.n321 10.6151
R2573 B.n326 B.n325 10.6151
R2574 B.n329 B.n326 10.6151
R2575 B.n330 B.n329 10.6151
R2576 B.n333 B.n330 10.6151
R2577 B.n334 B.n333 10.6151
R2578 B.n337 B.n334 10.6151
R2579 B.n338 B.n337 10.6151
R2580 B.n341 B.n338 10.6151
R2581 B.n342 B.n341 10.6151
R2582 B.n345 B.n342 10.6151
R2583 B.n346 B.n345 10.6151
R2584 B.n349 B.n346 10.6151
R2585 B.n350 B.n349 10.6151
R2586 B.n353 B.n350 10.6151
R2587 B.n354 B.n353 10.6151
R2588 B.n357 B.n354 10.6151
R2589 B.n358 B.n357 10.6151
R2590 B.n361 B.n358 10.6151
R2591 B.n362 B.n361 10.6151
R2592 B.n365 B.n362 10.6151
R2593 B.n366 B.n365 10.6151
R2594 B.n369 B.n366 10.6151
R2595 B.n370 B.n369 10.6151
R2596 B.n373 B.n370 10.6151
R2597 B.n374 B.n373 10.6151
R2598 B.n377 B.n374 10.6151
R2599 B.n378 B.n377 10.6151
R2600 B.n381 B.n378 10.6151
R2601 B.n382 B.n381 10.6151
R2602 B.n385 B.n382 10.6151
R2603 B.n386 B.n385 10.6151
R2604 B.n389 B.n386 10.6151
R2605 B.n390 B.n389 10.6151
R2606 B.n393 B.n390 10.6151
R2607 B.n394 B.n393 10.6151
R2608 B.n397 B.n394 10.6151
R2609 B.n398 B.n397 10.6151
R2610 B.n401 B.n398 10.6151
R2611 B.n402 B.n401 10.6151
R2612 B.n405 B.n402 10.6151
R2613 B.n406 B.n405 10.6151
R2614 B.n409 B.n406 10.6151
R2615 B.n410 B.n409 10.6151
R2616 B.n413 B.n410 10.6151
R2617 B.n415 B.n413 10.6151
R2618 B.n416 B.n415 10.6151
R2619 B.n1206 B.n416 10.6151
R2620 B.n757 B.n756 9.36635
R2621 B.n735 B.n734 9.36635
R2622 B.n302 B.n211 9.36635
R2623 B.n325 B.n208 9.36635
R2624 B.n1382 B.n0 8.11757
R2625 B.n1382 B.n1 8.11757
R2626 B.t9 B.n503 2.24483
R2627 B.n1041 B.t8 2.24483
R2628 B.n1338 B.t4 2.24483
R2629 B.n1289 B.t7 2.24483
R2630 B.n756 B.n755 1.24928
R2631 B.n736 B.n735 1.24928
R2632 B.n305 B.n211 1.24928
R2633 B.n322 B.n208 1.24928
R2634 VP.n35 VP.n32 161.3
R2635 VP.n37 VP.n36 161.3
R2636 VP.n38 VP.n31 161.3
R2637 VP.n40 VP.n39 161.3
R2638 VP.n41 VP.n30 161.3
R2639 VP.n43 VP.n42 161.3
R2640 VP.n44 VP.n29 161.3
R2641 VP.n46 VP.n45 161.3
R2642 VP.n47 VP.n28 161.3
R2643 VP.n49 VP.n48 161.3
R2644 VP.n50 VP.n27 161.3
R2645 VP.n52 VP.n51 161.3
R2646 VP.n53 VP.n26 161.3
R2647 VP.n55 VP.n54 161.3
R2648 VP.n56 VP.n25 161.3
R2649 VP.n58 VP.n57 161.3
R2650 VP.n59 VP.n24 161.3
R2651 VP.n62 VP.n61 161.3
R2652 VP.n63 VP.n23 161.3
R2653 VP.n65 VP.n64 161.3
R2654 VP.n66 VP.n22 161.3
R2655 VP.n68 VP.n67 161.3
R2656 VP.n69 VP.n21 161.3
R2657 VP.n71 VP.n70 161.3
R2658 VP.n72 VP.n20 161.3
R2659 VP.n74 VP.n73 161.3
R2660 VP.n131 VP.n130 161.3
R2661 VP.n129 VP.n1 161.3
R2662 VP.n128 VP.n127 161.3
R2663 VP.n126 VP.n2 161.3
R2664 VP.n125 VP.n124 161.3
R2665 VP.n123 VP.n3 161.3
R2666 VP.n122 VP.n121 161.3
R2667 VP.n120 VP.n4 161.3
R2668 VP.n119 VP.n118 161.3
R2669 VP.n116 VP.n5 161.3
R2670 VP.n115 VP.n114 161.3
R2671 VP.n113 VP.n6 161.3
R2672 VP.n112 VP.n111 161.3
R2673 VP.n110 VP.n7 161.3
R2674 VP.n109 VP.n108 161.3
R2675 VP.n107 VP.n8 161.3
R2676 VP.n106 VP.n105 161.3
R2677 VP.n104 VP.n9 161.3
R2678 VP.n103 VP.n102 161.3
R2679 VP.n101 VP.n10 161.3
R2680 VP.n100 VP.n99 161.3
R2681 VP.n98 VP.n11 161.3
R2682 VP.n97 VP.n96 161.3
R2683 VP.n95 VP.n12 161.3
R2684 VP.n94 VP.n93 161.3
R2685 VP.n92 VP.n13 161.3
R2686 VP.n90 VP.n89 161.3
R2687 VP.n88 VP.n14 161.3
R2688 VP.n87 VP.n86 161.3
R2689 VP.n85 VP.n15 161.3
R2690 VP.n84 VP.n83 161.3
R2691 VP.n82 VP.n16 161.3
R2692 VP.n81 VP.n80 161.3
R2693 VP.n79 VP.n17 161.3
R2694 VP.n78 VP.n77 161.3
R2695 VP.n33 VP.t1 120.221
R2696 VP.n76 VP.n18 88.1101
R2697 VP.n132 VP.n0 88.1101
R2698 VP.n75 VP.n19 88.1101
R2699 VP.n104 VP.t3 87.6535
R2700 VP.n18 VP.t2 87.6535
R2701 VP.n91 VP.t4 87.6535
R2702 VP.n117 VP.t6 87.6535
R2703 VP.n0 VP.t8 87.6535
R2704 VP.n47 VP.t0 87.6535
R2705 VP.n19 VP.t7 87.6535
R2706 VP.n60 VP.t5 87.6535
R2707 VP.n34 VP.t9 87.6535
R2708 VP.n76 VP.n75 62.238
R2709 VP.n34 VP.n33 61.9406
R2710 VP.n98 VP.n97 53.6055
R2711 VP.n111 VP.n110 53.6055
R2712 VP.n54 VP.n53 53.6055
R2713 VP.n41 VP.n40 53.6055
R2714 VP.n85 VP.n84 49.7204
R2715 VP.n124 VP.n123 49.7204
R2716 VP.n67 VP.n66 49.7204
R2717 VP.n84 VP.n16 31.2664
R2718 VP.n124 VP.n2 31.2664
R2719 VP.n67 VP.n21 31.2664
R2720 VP.n99 VP.n98 27.3813
R2721 VP.n110 VP.n109 27.3813
R2722 VP.n53 VP.n52 27.3813
R2723 VP.n42 VP.n41 27.3813
R2724 VP.n79 VP.n78 24.4675
R2725 VP.n80 VP.n79 24.4675
R2726 VP.n80 VP.n16 24.4675
R2727 VP.n86 VP.n85 24.4675
R2728 VP.n86 VP.n14 24.4675
R2729 VP.n90 VP.n14 24.4675
R2730 VP.n93 VP.n92 24.4675
R2731 VP.n93 VP.n12 24.4675
R2732 VP.n97 VP.n12 24.4675
R2733 VP.n99 VP.n10 24.4675
R2734 VP.n103 VP.n10 24.4675
R2735 VP.n104 VP.n103 24.4675
R2736 VP.n105 VP.n104 24.4675
R2737 VP.n105 VP.n8 24.4675
R2738 VP.n109 VP.n8 24.4675
R2739 VP.n111 VP.n6 24.4675
R2740 VP.n115 VP.n6 24.4675
R2741 VP.n116 VP.n115 24.4675
R2742 VP.n118 VP.n4 24.4675
R2743 VP.n122 VP.n4 24.4675
R2744 VP.n123 VP.n122 24.4675
R2745 VP.n128 VP.n2 24.4675
R2746 VP.n129 VP.n128 24.4675
R2747 VP.n130 VP.n129 24.4675
R2748 VP.n71 VP.n21 24.4675
R2749 VP.n72 VP.n71 24.4675
R2750 VP.n73 VP.n72 24.4675
R2751 VP.n54 VP.n25 24.4675
R2752 VP.n58 VP.n25 24.4675
R2753 VP.n59 VP.n58 24.4675
R2754 VP.n61 VP.n23 24.4675
R2755 VP.n65 VP.n23 24.4675
R2756 VP.n66 VP.n65 24.4675
R2757 VP.n42 VP.n29 24.4675
R2758 VP.n46 VP.n29 24.4675
R2759 VP.n47 VP.n46 24.4675
R2760 VP.n48 VP.n47 24.4675
R2761 VP.n48 VP.n27 24.4675
R2762 VP.n52 VP.n27 24.4675
R2763 VP.n36 VP.n35 24.4675
R2764 VP.n36 VP.n31 24.4675
R2765 VP.n40 VP.n31 24.4675
R2766 VP.n92 VP.n91 13.2127
R2767 VP.n117 VP.n116 13.2127
R2768 VP.n60 VP.n59 13.2127
R2769 VP.n35 VP.n34 13.2127
R2770 VP.n91 VP.n90 11.2553
R2771 VP.n118 VP.n117 11.2553
R2772 VP.n61 VP.n60 11.2553
R2773 VP.n33 VP.n32 2.48785
R2774 VP.n78 VP.n18 1.95786
R2775 VP.n130 VP.n0 1.95786
R2776 VP.n73 VP.n19 1.95786
R2777 VP.n75 VP.n74 0.354971
R2778 VP.n77 VP.n76 0.354971
R2779 VP.n132 VP.n131 0.354971
R2780 VP VP.n132 0.26696
R2781 VP.n37 VP.n32 0.189894
R2782 VP.n38 VP.n37 0.189894
R2783 VP.n39 VP.n38 0.189894
R2784 VP.n39 VP.n30 0.189894
R2785 VP.n43 VP.n30 0.189894
R2786 VP.n44 VP.n43 0.189894
R2787 VP.n45 VP.n44 0.189894
R2788 VP.n45 VP.n28 0.189894
R2789 VP.n49 VP.n28 0.189894
R2790 VP.n50 VP.n49 0.189894
R2791 VP.n51 VP.n50 0.189894
R2792 VP.n51 VP.n26 0.189894
R2793 VP.n55 VP.n26 0.189894
R2794 VP.n56 VP.n55 0.189894
R2795 VP.n57 VP.n56 0.189894
R2796 VP.n57 VP.n24 0.189894
R2797 VP.n62 VP.n24 0.189894
R2798 VP.n63 VP.n62 0.189894
R2799 VP.n64 VP.n63 0.189894
R2800 VP.n64 VP.n22 0.189894
R2801 VP.n68 VP.n22 0.189894
R2802 VP.n69 VP.n68 0.189894
R2803 VP.n70 VP.n69 0.189894
R2804 VP.n70 VP.n20 0.189894
R2805 VP.n74 VP.n20 0.189894
R2806 VP.n77 VP.n17 0.189894
R2807 VP.n81 VP.n17 0.189894
R2808 VP.n82 VP.n81 0.189894
R2809 VP.n83 VP.n82 0.189894
R2810 VP.n83 VP.n15 0.189894
R2811 VP.n87 VP.n15 0.189894
R2812 VP.n88 VP.n87 0.189894
R2813 VP.n89 VP.n88 0.189894
R2814 VP.n89 VP.n13 0.189894
R2815 VP.n94 VP.n13 0.189894
R2816 VP.n95 VP.n94 0.189894
R2817 VP.n96 VP.n95 0.189894
R2818 VP.n96 VP.n11 0.189894
R2819 VP.n100 VP.n11 0.189894
R2820 VP.n101 VP.n100 0.189894
R2821 VP.n102 VP.n101 0.189894
R2822 VP.n102 VP.n9 0.189894
R2823 VP.n106 VP.n9 0.189894
R2824 VP.n107 VP.n106 0.189894
R2825 VP.n108 VP.n107 0.189894
R2826 VP.n108 VP.n7 0.189894
R2827 VP.n112 VP.n7 0.189894
R2828 VP.n113 VP.n112 0.189894
R2829 VP.n114 VP.n113 0.189894
R2830 VP.n114 VP.n5 0.189894
R2831 VP.n119 VP.n5 0.189894
R2832 VP.n120 VP.n119 0.189894
R2833 VP.n121 VP.n120 0.189894
R2834 VP.n121 VP.n3 0.189894
R2835 VP.n125 VP.n3 0.189894
R2836 VP.n126 VP.n125 0.189894
R2837 VP.n127 VP.n126 0.189894
R2838 VP.n127 VP.n1 0.189894
R2839 VP.n131 VP.n1 0.189894
R2840 VDD1.n1 VDD1.t8 66.9983
R2841 VDD1.n3 VDD1.t7 66.9982
R2842 VDD1.n5 VDD1.n4 64.6408
R2843 VDD1.n1 VDD1.n0 61.9356
R2844 VDD1.n7 VDD1.n6 61.9354
R2845 VDD1.n3 VDD1.n2 61.9353
R2846 VDD1.n7 VDD1.n5 55.9772
R2847 VDD1 VDD1.n7 2.70309
R2848 VDD1.n6 VDD1.t4 1.38222
R2849 VDD1.n6 VDD1.t2 1.38222
R2850 VDD1.n0 VDD1.t0 1.38222
R2851 VDD1.n0 VDD1.t9 1.38222
R2852 VDD1.n4 VDD1.t3 1.38222
R2853 VDD1.n4 VDD1.t1 1.38222
R2854 VDD1.n2 VDD1.t5 1.38222
R2855 VDD1.n2 VDD1.t6 1.38222
R2856 VDD1 VDD1.n1 0.978948
R2857 VDD1.n5 VDD1.n3 0.865413
C0 VP VN 10.8049f
C1 VTAIL VP 14.6614f
C2 VP VDD2 0.753897f
C3 VDD1 VP 14.136499f
C4 VTAIL VN 14.6464f
C5 VN VDD2 13.5425f
C6 VDD1 VN 0.156412f
C7 VTAIL VDD2 12.0667f
C8 VTAIL VDD1 12.006f
C9 VDD1 VDD2 3.04761f
C10 VDD2 B 9.170935f
C11 VDD1 B 9.160812f
C12 VTAIL B 10.15655f
C13 VN B 24.70798f
C14 VP B 23.289326f
C15 VDD1.t8 B 3.2538f
C16 VDD1.t0 B 0.279831f
C17 VDD1.t9 B 0.279831f
C18 VDD1.n0 B 2.52499f
C19 VDD1.n1 B 1.10947f
C20 VDD1.t7 B 3.25378f
C21 VDD1.t5 B 0.279831f
C22 VDD1.t6 B 0.279831f
C23 VDD1.n2 B 2.52499f
C24 VDD1.n3 B 1.10111f
C25 VDD1.t3 B 0.279831f
C26 VDD1.t1 B 0.279831f
C27 VDD1.n4 B 2.55509f
C28 VDD1.n5 B 3.86356f
C29 VDD1.t4 B 0.279831f
C30 VDD1.t2 B 0.279831f
C31 VDD1.n6 B 2.52498f
C32 VDD1.n7 B 3.85648f
C33 VP.t8 B 2.49633f
C34 VP.n0 B 0.928728f
C35 VP.n1 B 0.016152f
C36 VP.n2 B 0.032431f
C37 VP.n3 B 0.016152f
C38 VP.n4 B 0.030104f
C39 VP.n5 B 0.016152f
C40 VP.t6 B 2.49633f
C41 VP.n6 B 0.030104f
C42 VP.n7 B 0.016152f
C43 VP.n8 B 0.030104f
C44 VP.n9 B 0.016152f
C45 VP.t3 B 2.49633f
C46 VP.n10 B 0.030104f
C47 VP.n11 B 0.016152f
C48 VP.n12 B 0.030104f
C49 VP.n13 B 0.016152f
C50 VP.t4 B 2.49633f
C51 VP.n14 B 0.030104f
C52 VP.n15 B 0.016152f
C53 VP.n16 B 0.032431f
C54 VP.n17 B 0.016152f
C55 VP.t2 B 2.49633f
C56 VP.n18 B 0.928728f
C57 VP.t7 B 2.49633f
C58 VP.n19 B 0.928728f
C59 VP.n20 B 0.016152f
C60 VP.n21 B 0.032431f
C61 VP.n22 B 0.016152f
C62 VP.n23 B 0.030104f
C63 VP.n24 B 0.016152f
C64 VP.t5 B 2.49633f
C65 VP.n25 B 0.030104f
C66 VP.n26 B 0.016152f
C67 VP.n27 B 0.030104f
C68 VP.n28 B 0.016152f
C69 VP.t0 B 2.49633f
C70 VP.n29 B 0.030104f
C71 VP.n30 B 0.016152f
C72 VP.n31 B 0.030104f
C73 VP.n32 B 0.210842f
C74 VP.t9 B 2.49633f
C75 VP.t1 B 2.76664f
C76 VP.n33 B 0.88221f
C77 VP.n34 B 0.926154f
C78 VP.n35 B 0.023268f
C79 VP.n36 B 0.030104f
C80 VP.n37 B 0.016152f
C81 VP.n38 B 0.016152f
C82 VP.n39 B 0.016152f
C83 VP.n40 B 0.028489f
C84 VP.n41 B 0.017282f
C85 VP.n42 B 0.031496f
C86 VP.n43 B 0.016152f
C87 VP.n44 B 0.016152f
C88 VP.n45 B 0.016152f
C89 VP.n46 B 0.030104f
C90 VP.n47 B 0.882032f
C91 VP.n48 B 0.030104f
C92 VP.n49 B 0.016152f
C93 VP.n50 B 0.016152f
C94 VP.n51 B 0.016152f
C95 VP.n52 B 0.031496f
C96 VP.n53 B 0.017282f
C97 VP.n54 B 0.028489f
C98 VP.n55 B 0.016152f
C99 VP.n56 B 0.016152f
C100 VP.n57 B 0.016152f
C101 VP.n58 B 0.030104f
C102 VP.n59 B 0.023268f
C103 VP.n60 B 0.866791f
C104 VP.n61 B 0.022079f
C105 VP.n62 B 0.016152f
C106 VP.n63 B 0.016152f
C107 VP.n64 B 0.016152f
C108 VP.n65 B 0.030104f
C109 VP.n66 B 0.029802f
C110 VP.n67 B 0.015033f
C111 VP.n68 B 0.016152f
C112 VP.n69 B 0.016152f
C113 VP.n70 B 0.016152f
C114 VP.n71 B 0.030104f
C115 VP.n72 B 0.030104f
C116 VP.n73 B 0.016431f
C117 VP.n74 B 0.02607f
C118 VP.n75 B 1.25476f
C119 VP.n76 B 1.26409f
C120 VP.n77 B 0.02607f
C121 VP.n78 B 0.016431f
C122 VP.n79 B 0.030104f
C123 VP.n80 B 0.030104f
C124 VP.n81 B 0.016152f
C125 VP.n82 B 0.016152f
C126 VP.n83 B 0.016152f
C127 VP.n84 B 0.015033f
C128 VP.n85 B 0.029802f
C129 VP.n86 B 0.030104f
C130 VP.n87 B 0.016152f
C131 VP.n88 B 0.016152f
C132 VP.n89 B 0.016152f
C133 VP.n90 B 0.022079f
C134 VP.n91 B 0.866791f
C135 VP.n92 B 0.023268f
C136 VP.n93 B 0.030104f
C137 VP.n94 B 0.016152f
C138 VP.n95 B 0.016152f
C139 VP.n96 B 0.016152f
C140 VP.n97 B 0.028489f
C141 VP.n98 B 0.017282f
C142 VP.n99 B 0.031496f
C143 VP.n100 B 0.016152f
C144 VP.n101 B 0.016152f
C145 VP.n102 B 0.016152f
C146 VP.n103 B 0.030104f
C147 VP.n104 B 0.882032f
C148 VP.n105 B 0.030104f
C149 VP.n106 B 0.016152f
C150 VP.n107 B 0.016152f
C151 VP.n108 B 0.016152f
C152 VP.n109 B 0.031496f
C153 VP.n110 B 0.017282f
C154 VP.n111 B 0.028489f
C155 VP.n112 B 0.016152f
C156 VP.n113 B 0.016152f
C157 VP.n114 B 0.016152f
C158 VP.n115 B 0.030104f
C159 VP.n116 B 0.023268f
C160 VP.n117 B 0.866791f
C161 VP.n118 B 0.022079f
C162 VP.n119 B 0.016152f
C163 VP.n120 B 0.016152f
C164 VP.n121 B 0.016152f
C165 VP.n122 B 0.030104f
C166 VP.n123 B 0.029802f
C167 VP.n124 B 0.015033f
C168 VP.n125 B 0.016152f
C169 VP.n126 B 0.016152f
C170 VP.n127 B 0.016152f
C171 VP.n128 B 0.030104f
C172 VP.n129 B 0.030104f
C173 VP.n130 B 0.016431f
C174 VP.n131 B 0.02607f
C175 VP.n132 B 0.051339f
C176 VDD2.t5 B 3.20794f
C177 VDD2.t7 B 0.275888f
C178 VDD2.t6 B 0.275888f
C179 VDD2.n0 B 2.48941f
C180 VDD2.n1 B 1.0856f
C181 VDD2.t2 B 0.275888f
C182 VDD2.t0 B 0.275888f
C183 VDD2.n2 B 2.51909f
C184 VDD2.n3 B 3.64932f
C185 VDD2.t1 B 3.17712f
C186 VDD2.n4 B 3.7245f
C187 VDD2.t8 B 0.275888f
C188 VDD2.t9 B 0.275888f
C189 VDD2.n5 B 2.48941f
C190 VDD2.n6 B 0.563478f
C191 VDD2.t3 B 0.275888f
C192 VDD2.t4 B 0.275888f
C193 VDD2.n7 B 2.51903f
C194 VTAIL.t13 B 0.285746f
C195 VTAIL.t17 B 0.285746f
C196 VTAIL.n0 B 2.50468f
C197 VTAIL.n1 B 0.661211f
C198 VTAIL.t5 B 3.19515f
C199 VTAIL.n2 B 0.820141f
C200 VTAIL.t0 B 0.285746f
C201 VTAIL.t8 B 0.285746f
C202 VTAIL.n3 B 2.50468f
C203 VTAIL.n4 B 0.842753f
C204 VTAIL.t2 B 0.285746f
C205 VTAIL.t9 B 0.285746f
C206 VTAIL.n5 B 2.50468f
C207 VTAIL.n6 B 2.48927f
C208 VTAIL.t14 B 0.285746f
C209 VTAIL.t18 B 0.285746f
C210 VTAIL.n7 B 2.50468f
C211 VTAIL.n8 B 2.48926f
C212 VTAIL.t19 B 0.285746f
C213 VTAIL.t15 B 0.285746f
C214 VTAIL.n9 B 2.50468f
C215 VTAIL.n10 B 0.84275f
C216 VTAIL.t11 B 3.19517f
C217 VTAIL.n11 B 0.820119f
C218 VTAIL.t1 B 0.285746f
C219 VTAIL.t4 B 0.285746f
C220 VTAIL.n12 B 2.50468f
C221 VTAIL.n13 B 0.731301f
C222 VTAIL.t3 B 0.285746f
C223 VTAIL.t7 B 0.285746f
C224 VTAIL.n14 B 2.50468f
C225 VTAIL.n15 B 0.84275f
C226 VTAIL.t6 B 3.19515f
C227 VTAIL.n16 B 2.2788f
C228 VTAIL.t12 B 3.19515f
C229 VTAIL.n17 B 2.2788f
C230 VTAIL.t16 B 0.285746f
C231 VTAIL.t10 B 0.285746f
C232 VTAIL.n18 B 2.50468f
C233 VTAIL.n19 B 0.613547f
C234 VN.t9 B 2.4508f
C235 VN.n0 B 0.911789f
C236 VN.n1 B 0.015858f
C237 VN.n2 B 0.03184f
C238 VN.n3 B 0.015858f
C239 VN.n4 B 0.029555f
C240 VN.n5 B 0.015858f
C241 VN.t7 B 2.4508f
C242 VN.n6 B 0.029555f
C243 VN.n7 B 0.015858f
C244 VN.n8 B 0.029555f
C245 VN.n9 B 0.015858f
C246 VN.t3 B 2.4508f
C247 VN.n10 B 0.029555f
C248 VN.n11 B 0.015858f
C249 VN.n12 B 0.029555f
C250 VN.n13 B 0.206996f
C251 VN.t2 B 2.4508f
C252 VN.t4 B 2.71618f
C253 VN.n14 B 0.866118f
C254 VN.n15 B 0.909261f
C255 VN.n16 B 0.022843f
C256 VN.n17 B 0.029555f
C257 VN.n18 B 0.015858f
C258 VN.n19 B 0.015858f
C259 VN.n20 B 0.015858f
C260 VN.n21 B 0.027969f
C261 VN.n22 B 0.016967f
C262 VN.n23 B 0.030922f
C263 VN.n24 B 0.015858f
C264 VN.n25 B 0.015858f
C265 VN.n26 B 0.015858f
C266 VN.n27 B 0.029555f
C267 VN.n28 B 0.865945f
C268 VN.n29 B 0.029555f
C269 VN.n30 B 0.015858f
C270 VN.n31 B 0.015858f
C271 VN.n32 B 0.015858f
C272 VN.n33 B 0.030922f
C273 VN.n34 B 0.016967f
C274 VN.n35 B 0.027969f
C275 VN.n36 B 0.015858f
C276 VN.n37 B 0.015858f
C277 VN.n38 B 0.015858f
C278 VN.n39 B 0.029555f
C279 VN.n40 B 0.022843f
C280 VN.n41 B 0.850981f
C281 VN.n42 B 0.021676f
C282 VN.n43 B 0.015858f
C283 VN.n44 B 0.015858f
C284 VN.n45 B 0.015858f
C285 VN.n46 B 0.029555f
C286 VN.n47 B 0.029259f
C287 VN.n48 B 0.014759f
C288 VN.n49 B 0.015858f
C289 VN.n50 B 0.015858f
C290 VN.n51 B 0.015858f
C291 VN.n52 B 0.029555f
C292 VN.n53 B 0.029555f
C293 VN.n54 B 0.016131f
C294 VN.n55 B 0.025594f
C295 VN.n56 B 0.050402f
C296 VN.t8 B 2.4508f
C297 VN.n57 B 0.911789f
C298 VN.n58 B 0.015858f
C299 VN.n59 B 0.03184f
C300 VN.n60 B 0.015858f
C301 VN.n61 B 0.029555f
C302 VN.n62 B 0.015858f
C303 VN.t1 B 2.4508f
C304 VN.n63 B 0.029555f
C305 VN.n64 B 0.015858f
C306 VN.n65 B 0.029555f
C307 VN.n66 B 0.015858f
C308 VN.t0 B 2.4508f
C309 VN.n67 B 0.029555f
C310 VN.n68 B 0.015858f
C311 VN.n69 B 0.029555f
C312 VN.n70 B 0.206996f
C313 VN.t6 B 2.4508f
C314 VN.t5 B 2.71618f
C315 VN.n71 B 0.866118f
C316 VN.n72 B 0.909261f
C317 VN.n73 B 0.022843f
C318 VN.n74 B 0.029555f
C319 VN.n75 B 0.015858f
C320 VN.n76 B 0.015858f
C321 VN.n77 B 0.015858f
C322 VN.n78 B 0.027969f
C323 VN.n79 B 0.016967f
C324 VN.n80 B 0.030922f
C325 VN.n81 B 0.015858f
C326 VN.n82 B 0.015858f
C327 VN.n83 B 0.015858f
C328 VN.n84 B 0.029555f
C329 VN.n85 B 0.865945f
C330 VN.n86 B 0.029555f
C331 VN.n87 B 0.015858f
C332 VN.n88 B 0.015858f
C333 VN.n89 B 0.015858f
C334 VN.n90 B 0.030922f
C335 VN.n91 B 0.016967f
C336 VN.n92 B 0.027969f
C337 VN.n93 B 0.015858f
C338 VN.n94 B 0.015858f
C339 VN.n95 B 0.015858f
C340 VN.n96 B 0.029555f
C341 VN.n97 B 0.022843f
C342 VN.n98 B 0.850981f
C343 VN.n99 B 0.021676f
C344 VN.n100 B 0.015858f
C345 VN.n101 B 0.015858f
C346 VN.n102 B 0.015858f
C347 VN.n103 B 0.029555f
C348 VN.n104 B 0.029259f
C349 VN.n105 B 0.014759f
C350 VN.n106 B 0.015858f
C351 VN.n107 B 0.015858f
C352 VN.n108 B 0.015858f
C353 VN.n109 B 0.029555f
C354 VN.n110 B 0.029555f
C355 VN.n111 B 0.016131f
C356 VN.n112 B 0.025594f
C357 VN.n113 B 1.23792f
.ends

