* NGSPICE file created from diff_pair_sample_0622.ext - technology: sky130A

.subckt diff_pair_sample_0622 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.17
X1 VDD1.t1 VP.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0.8424 ps=5.1 w=2.16 l=2.17
X2 VDD1.t0 VP.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0.8424 ps=5.1 w=2.16 l=2.17
X3 VDD2.t1 VN.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0.8424 ps=5.1 w=2.16 l=2.17
X4 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.17
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.17
X6 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0.8424 ps=5.1 w=2.16 l=2.17
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.8424 pd=5.1 as=0 ps=0 w=2.16 l=2.17
R0 B.n370 B.n369 585
R1 B.n371 B.n370 585
R2 B.n133 B.n63 585
R3 B.n132 B.n131 585
R4 B.n130 B.n129 585
R5 B.n128 B.n127 585
R6 B.n126 B.n125 585
R7 B.n124 B.n123 585
R8 B.n122 B.n121 585
R9 B.n120 B.n119 585
R10 B.n118 B.n117 585
R11 B.n116 B.n115 585
R12 B.n114 B.n113 585
R13 B.n112 B.n111 585
R14 B.n110 B.n109 585
R15 B.n108 B.n107 585
R16 B.n106 B.n105 585
R17 B.n104 B.n103 585
R18 B.n102 B.n101 585
R19 B.n100 B.n99 585
R20 B.n98 B.n97 585
R21 B.n96 B.n95 585
R22 B.n94 B.n93 585
R23 B.n91 B.n90 585
R24 B.n89 B.n88 585
R25 B.n87 B.n86 585
R26 B.n85 B.n84 585
R27 B.n83 B.n82 585
R28 B.n81 B.n80 585
R29 B.n79 B.n78 585
R30 B.n77 B.n76 585
R31 B.n75 B.n74 585
R32 B.n73 B.n72 585
R33 B.n71 B.n70 585
R34 B.n46 B.n45 585
R35 B.n374 B.n373 585
R36 B.n368 B.n64 585
R37 B.n64 B.n43 585
R38 B.n367 B.n42 585
R39 B.n378 B.n42 585
R40 B.n366 B.n41 585
R41 B.n379 B.n41 585
R42 B.n365 B.n40 585
R43 B.n380 B.n40 585
R44 B.n364 B.n363 585
R45 B.n363 B.n36 585
R46 B.n362 B.n35 585
R47 B.n386 B.n35 585
R48 B.n361 B.n34 585
R49 B.n387 B.n34 585
R50 B.n360 B.n33 585
R51 B.n388 B.n33 585
R52 B.n359 B.n358 585
R53 B.n358 B.n29 585
R54 B.n357 B.n28 585
R55 B.n394 B.n28 585
R56 B.n356 B.n27 585
R57 B.n395 B.n27 585
R58 B.n355 B.n26 585
R59 B.n396 B.n26 585
R60 B.n354 B.n353 585
R61 B.n353 B.n22 585
R62 B.n352 B.n21 585
R63 B.n402 B.n21 585
R64 B.n351 B.n20 585
R65 B.n403 B.n20 585
R66 B.n350 B.n19 585
R67 B.n404 B.n19 585
R68 B.n349 B.n348 585
R69 B.n348 B.n15 585
R70 B.n347 B.n14 585
R71 B.n410 B.n14 585
R72 B.n346 B.n13 585
R73 B.n411 B.n13 585
R74 B.n345 B.n12 585
R75 B.n412 B.n12 585
R76 B.n344 B.n343 585
R77 B.n343 B.n8 585
R78 B.n342 B.n7 585
R79 B.n418 B.n7 585
R80 B.n341 B.n6 585
R81 B.n419 B.n6 585
R82 B.n340 B.n5 585
R83 B.n420 B.n5 585
R84 B.n339 B.n338 585
R85 B.n338 B.n4 585
R86 B.n337 B.n134 585
R87 B.n337 B.n336 585
R88 B.n327 B.n135 585
R89 B.n136 B.n135 585
R90 B.n329 B.n328 585
R91 B.n330 B.n329 585
R92 B.n326 B.n141 585
R93 B.n141 B.n140 585
R94 B.n325 B.n324 585
R95 B.n324 B.n323 585
R96 B.n143 B.n142 585
R97 B.n144 B.n143 585
R98 B.n316 B.n315 585
R99 B.n317 B.n316 585
R100 B.n314 B.n149 585
R101 B.n149 B.n148 585
R102 B.n313 B.n312 585
R103 B.n312 B.n311 585
R104 B.n151 B.n150 585
R105 B.n152 B.n151 585
R106 B.n304 B.n303 585
R107 B.n305 B.n304 585
R108 B.n302 B.n157 585
R109 B.n157 B.n156 585
R110 B.n301 B.n300 585
R111 B.n300 B.n299 585
R112 B.n159 B.n158 585
R113 B.n160 B.n159 585
R114 B.n292 B.n291 585
R115 B.n293 B.n292 585
R116 B.n290 B.n165 585
R117 B.n165 B.n164 585
R118 B.n289 B.n288 585
R119 B.n288 B.n287 585
R120 B.n167 B.n166 585
R121 B.n168 B.n167 585
R122 B.n280 B.n279 585
R123 B.n281 B.n280 585
R124 B.n278 B.n173 585
R125 B.n173 B.n172 585
R126 B.n277 B.n276 585
R127 B.n276 B.n275 585
R128 B.n175 B.n174 585
R129 B.n176 B.n175 585
R130 B.n271 B.n270 585
R131 B.n179 B.n178 585
R132 B.n267 B.n266 585
R133 B.n268 B.n267 585
R134 B.n265 B.n196 585
R135 B.n264 B.n263 585
R136 B.n262 B.n261 585
R137 B.n260 B.n259 585
R138 B.n258 B.n257 585
R139 B.n256 B.n255 585
R140 B.n254 B.n253 585
R141 B.n252 B.n251 585
R142 B.n250 B.n249 585
R143 B.n248 B.n247 585
R144 B.n246 B.n245 585
R145 B.n244 B.n243 585
R146 B.n242 B.n241 585
R147 B.n240 B.n239 585
R148 B.n238 B.n237 585
R149 B.n236 B.n235 585
R150 B.n234 B.n233 585
R151 B.n232 B.n231 585
R152 B.n230 B.n229 585
R153 B.n227 B.n226 585
R154 B.n225 B.n224 585
R155 B.n223 B.n222 585
R156 B.n221 B.n220 585
R157 B.n219 B.n218 585
R158 B.n217 B.n216 585
R159 B.n215 B.n214 585
R160 B.n213 B.n212 585
R161 B.n211 B.n210 585
R162 B.n209 B.n208 585
R163 B.n207 B.n206 585
R164 B.n205 B.n204 585
R165 B.n203 B.n202 585
R166 B.n272 B.n177 585
R167 B.n177 B.n176 585
R168 B.n274 B.n273 585
R169 B.n275 B.n274 585
R170 B.n171 B.n170 585
R171 B.n172 B.n171 585
R172 B.n283 B.n282 585
R173 B.n282 B.n281 585
R174 B.n284 B.n169 585
R175 B.n169 B.n168 585
R176 B.n286 B.n285 585
R177 B.n287 B.n286 585
R178 B.n163 B.n162 585
R179 B.n164 B.n163 585
R180 B.n295 B.n294 585
R181 B.n294 B.n293 585
R182 B.n296 B.n161 585
R183 B.n161 B.n160 585
R184 B.n298 B.n297 585
R185 B.n299 B.n298 585
R186 B.n155 B.n154 585
R187 B.n156 B.n155 585
R188 B.n307 B.n306 585
R189 B.n306 B.n305 585
R190 B.n308 B.n153 585
R191 B.n153 B.n152 585
R192 B.n310 B.n309 585
R193 B.n311 B.n310 585
R194 B.n147 B.n146 585
R195 B.n148 B.n147 585
R196 B.n319 B.n318 585
R197 B.n318 B.n317 585
R198 B.n320 B.n145 585
R199 B.n145 B.n144 585
R200 B.n322 B.n321 585
R201 B.n323 B.n322 585
R202 B.n139 B.n138 585
R203 B.n140 B.n139 585
R204 B.n332 B.n331 585
R205 B.n331 B.n330 585
R206 B.n333 B.n137 585
R207 B.n137 B.n136 585
R208 B.n335 B.n334 585
R209 B.n336 B.n335 585
R210 B.n2 B.n0 585
R211 B.n4 B.n2 585
R212 B.n3 B.n1 585
R213 B.n419 B.n3 585
R214 B.n417 B.n416 585
R215 B.n418 B.n417 585
R216 B.n415 B.n9 585
R217 B.n9 B.n8 585
R218 B.n414 B.n413 585
R219 B.n413 B.n412 585
R220 B.n11 B.n10 585
R221 B.n411 B.n11 585
R222 B.n409 B.n408 585
R223 B.n410 B.n409 585
R224 B.n407 B.n16 585
R225 B.n16 B.n15 585
R226 B.n406 B.n405 585
R227 B.n405 B.n404 585
R228 B.n18 B.n17 585
R229 B.n403 B.n18 585
R230 B.n401 B.n400 585
R231 B.n402 B.n401 585
R232 B.n399 B.n23 585
R233 B.n23 B.n22 585
R234 B.n398 B.n397 585
R235 B.n397 B.n396 585
R236 B.n25 B.n24 585
R237 B.n395 B.n25 585
R238 B.n393 B.n392 585
R239 B.n394 B.n393 585
R240 B.n391 B.n30 585
R241 B.n30 B.n29 585
R242 B.n390 B.n389 585
R243 B.n389 B.n388 585
R244 B.n32 B.n31 585
R245 B.n387 B.n32 585
R246 B.n385 B.n384 585
R247 B.n386 B.n385 585
R248 B.n383 B.n37 585
R249 B.n37 B.n36 585
R250 B.n382 B.n381 585
R251 B.n381 B.n380 585
R252 B.n39 B.n38 585
R253 B.n379 B.n39 585
R254 B.n377 B.n376 585
R255 B.n378 B.n377 585
R256 B.n375 B.n44 585
R257 B.n44 B.n43 585
R258 B.n422 B.n421 585
R259 B.n421 B.n420 585
R260 B.n270 B.n177 463.671
R261 B.n373 B.n44 463.671
R262 B.n202 B.n175 463.671
R263 B.n370 B.n64 463.671
R264 B.n371 B.n62 256.663
R265 B.n371 B.n61 256.663
R266 B.n371 B.n60 256.663
R267 B.n371 B.n59 256.663
R268 B.n371 B.n58 256.663
R269 B.n371 B.n57 256.663
R270 B.n371 B.n56 256.663
R271 B.n371 B.n55 256.663
R272 B.n371 B.n54 256.663
R273 B.n371 B.n53 256.663
R274 B.n371 B.n52 256.663
R275 B.n371 B.n51 256.663
R276 B.n371 B.n50 256.663
R277 B.n371 B.n49 256.663
R278 B.n371 B.n48 256.663
R279 B.n371 B.n47 256.663
R280 B.n372 B.n371 256.663
R281 B.n269 B.n268 256.663
R282 B.n268 B.n180 256.663
R283 B.n268 B.n181 256.663
R284 B.n268 B.n182 256.663
R285 B.n268 B.n183 256.663
R286 B.n268 B.n184 256.663
R287 B.n268 B.n185 256.663
R288 B.n268 B.n186 256.663
R289 B.n268 B.n187 256.663
R290 B.n268 B.n188 256.663
R291 B.n268 B.n189 256.663
R292 B.n268 B.n190 256.663
R293 B.n268 B.n191 256.663
R294 B.n268 B.n192 256.663
R295 B.n268 B.n193 256.663
R296 B.n268 B.n194 256.663
R297 B.n268 B.n195 256.663
R298 B.n200 B.t10 231.28
R299 B.n197 B.t6 231.28
R300 B.n68 B.t13 231.28
R301 B.n65 B.t2 231.28
R302 B.n268 B.n176 164.224
R303 B.n371 B.n43 164.224
R304 B.n274 B.n177 163.367
R305 B.n274 B.n171 163.367
R306 B.n282 B.n171 163.367
R307 B.n282 B.n169 163.367
R308 B.n286 B.n169 163.367
R309 B.n286 B.n163 163.367
R310 B.n294 B.n163 163.367
R311 B.n294 B.n161 163.367
R312 B.n298 B.n161 163.367
R313 B.n298 B.n155 163.367
R314 B.n306 B.n155 163.367
R315 B.n306 B.n153 163.367
R316 B.n310 B.n153 163.367
R317 B.n310 B.n147 163.367
R318 B.n318 B.n147 163.367
R319 B.n318 B.n145 163.367
R320 B.n322 B.n145 163.367
R321 B.n322 B.n139 163.367
R322 B.n331 B.n139 163.367
R323 B.n331 B.n137 163.367
R324 B.n335 B.n137 163.367
R325 B.n335 B.n2 163.367
R326 B.n421 B.n2 163.367
R327 B.n421 B.n3 163.367
R328 B.n417 B.n3 163.367
R329 B.n417 B.n9 163.367
R330 B.n413 B.n9 163.367
R331 B.n413 B.n11 163.367
R332 B.n409 B.n11 163.367
R333 B.n409 B.n16 163.367
R334 B.n405 B.n16 163.367
R335 B.n405 B.n18 163.367
R336 B.n401 B.n18 163.367
R337 B.n401 B.n23 163.367
R338 B.n397 B.n23 163.367
R339 B.n397 B.n25 163.367
R340 B.n393 B.n25 163.367
R341 B.n393 B.n30 163.367
R342 B.n389 B.n30 163.367
R343 B.n389 B.n32 163.367
R344 B.n385 B.n32 163.367
R345 B.n385 B.n37 163.367
R346 B.n381 B.n37 163.367
R347 B.n381 B.n39 163.367
R348 B.n377 B.n39 163.367
R349 B.n377 B.n44 163.367
R350 B.n267 B.n179 163.367
R351 B.n267 B.n196 163.367
R352 B.n263 B.n262 163.367
R353 B.n259 B.n258 163.367
R354 B.n255 B.n254 163.367
R355 B.n251 B.n250 163.367
R356 B.n247 B.n246 163.367
R357 B.n243 B.n242 163.367
R358 B.n239 B.n238 163.367
R359 B.n235 B.n234 163.367
R360 B.n231 B.n230 163.367
R361 B.n226 B.n225 163.367
R362 B.n222 B.n221 163.367
R363 B.n218 B.n217 163.367
R364 B.n214 B.n213 163.367
R365 B.n210 B.n209 163.367
R366 B.n206 B.n205 163.367
R367 B.n276 B.n175 163.367
R368 B.n276 B.n173 163.367
R369 B.n280 B.n173 163.367
R370 B.n280 B.n167 163.367
R371 B.n288 B.n167 163.367
R372 B.n288 B.n165 163.367
R373 B.n292 B.n165 163.367
R374 B.n292 B.n159 163.367
R375 B.n300 B.n159 163.367
R376 B.n300 B.n157 163.367
R377 B.n304 B.n157 163.367
R378 B.n304 B.n151 163.367
R379 B.n312 B.n151 163.367
R380 B.n312 B.n149 163.367
R381 B.n316 B.n149 163.367
R382 B.n316 B.n143 163.367
R383 B.n324 B.n143 163.367
R384 B.n324 B.n141 163.367
R385 B.n329 B.n141 163.367
R386 B.n329 B.n135 163.367
R387 B.n337 B.n135 163.367
R388 B.n338 B.n337 163.367
R389 B.n338 B.n5 163.367
R390 B.n6 B.n5 163.367
R391 B.n7 B.n6 163.367
R392 B.n343 B.n7 163.367
R393 B.n343 B.n12 163.367
R394 B.n13 B.n12 163.367
R395 B.n14 B.n13 163.367
R396 B.n348 B.n14 163.367
R397 B.n348 B.n19 163.367
R398 B.n20 B.n19 163.367
R399 B.n21 B.n20 163.367
R400 B.n353 B.n21 163.367
R401 B.n353 B.n26 163.367
R402 B.n27 B.n26 163.367
R403 B.n28 B.n27 163.367
R404 B.n358 B.n28 163.367
R405 B.n358 B.n33 163.367
R406 B.n34 B.n33 163.367
R407 B.n35 B.n34 163.367
R408 B.n363 B.n35 163.367
R409 B.n363 B.n40 163.367
R410 B.n41 B.n40 163.367
R411 B.n42 B.n41 163.367
R412 B.n64 B.n42 163.367
R413 B.n70 B.n46 163.367
R414 B.n74 B.n73 163.367
R415 B.n78 B.n77 163.367
R416 B.n82 B.n81 163.367
R417 B.n86 B.n85 163.367
R418 B.n90 B.n89 163.367
R419 B.n95 B.n94 163.367
R420 B.n99 B.n98 163.367
R421 B.n103 B.n102 163.367
R422 B.n107 B.n106 163.367
R423 B.n111 B.n110 163.367
R424 B.n115 B.n114 163.367
R425 B.n119 B.n118 163.367
R426 B.n123 B.n122 163.367
R427 B.n127 B.n126 163.367
R428 B.n131 B.n130 163.367
R429 B.n370 B.n63 163.367
R430 B.n200 B.t12 133.583
R431 B.n65 B.t4 133.583
R432 B.n197 B.t9 133.583
R433 B.n68 B.t14 133.583
R434 B.n275 B.n176 100.606
R435 B.n275 B.n172 100.606
R436 B.n281 B.n172 100.606
R437 B.n281 B.n168 100.606
R438 B.n287 B.n168 100.606
R439 B.n287 B.n164 100.606
R440 B.n293 B.n164 100.606
R441 B.n299 B.n160 100.606
R442 B.n299 B.n156 100.606
R443 B.n305 B.n156 100.606
R444 B.n305 B.n152 100.606
R445 B.n311 B.n152 100.606
R446 B.n311 B.n148 100.606
R447 B.n317 B.n148 100.606
R448 B.n317 B.n144 100.606
R449 B.n323 B.n144 100.606
R450 B.n330 B.n140 100.606
R451 B.n330 B.n136 100.606
R452 B.n336 B.n136 100.606
R453 B.n336 B.n4 100.606
R454 B.n420 B.n4 100.606
R455 B.n420 B.n419 100.606
R456 B.n419 B.n418 100.606
R457 B.n418 B.n8 100.606
R458 B.n412 B.n8 100.606
R459 B.n412 B.n411 100.606
R460 B.n410 B.n15 100.606
R461 B.n404 B.n15 100.606
R462 B.n404 B.n403 100.606
R463 B.n403 B.n402 100.606
R464 B.n402 B.n22 100.606
R465 B.n396 B.n22 100.606
R466 B.n396 B.n395 100.606
R467 B.n395 B.n394 100.606
R468 B.n394 B.n29 100.606
R469 B.n388 B.n387 100.606
R470 B.n387 B.n386 100.606
R471 B.n386 B.n36 100.606
R472 B.n380 B.n36 100.606
R473 B.n380 B.n379 100.606
R474 B.n379 B.n378 100.606
R475 B.n378 B.n43 100.606
R476 B.n201 B.t11 85.0987
R477 B.n66 B.t5 85.0987
R478 B.n198 B.t8 85.0984
R479 B.n69 B.t15 85.0984
R480 B.t7 B.n160 84.3314
R481 B.t3 B.n29 84.3314
R482 B.n323 B.t1 72.4954
R483 B.t0 B.n410 72.4954
R484 B.n270 B.n269 71.676
R485 B.n196 B.n180 71.676
R486 B.n262 B.n181 71.676
R487 B.n258 B.n182 71.676
R488 B.n254 B.n183 71.676
R489 B.n250 B.n184 71.676
R490 B.n246 B.n185 71.676
R491 B.n242 B.n186 71.676
R492 B.n238 B.n187 71.676
R493 B.n234 B.n188 71.676
R494 B.n230 B.n189 71.676
R495 B.n225 B.n190 71.676
R496 B.n221 B.n191 71.676
R497 B.n217 B.n192 71.676
R498 B.n213 B.n193 71.676
R499 B.n209 B.n194 71.676
R500 B.n205 B.n195 71.676
R501 B.n373 B.n372 71.676
R502 B.n70 B.n47 71.676
R503 B.n74 B.n48 71.676
R504 B.n78 B.n49 71.676
R505 B.n82 B.n50 71.676
R506 B.n86 B.n51 71.676
R507 B.n90 B.n52 71.676
R508 B.n95 B.n53 71.676
R509 B.n99 B.n54 71.676
R510 B.n103 B.n55 71.676
R511 B.n107 B.n56 71.676
R512 B.n111 B.n57 71.676
R513 B.n115 B.n58 71.676
R514 B.n119 B.n59 71.676
R515 B.n123 B.n60 71.676
R516 B.n127 B.n61 71.676
R517 B.n131 B.n62 71.676
R518 B.n63 B.n62 71.676
R519 B.n130 B.n61 71.676
R520 B.n126 B.n60 71.676
R521 B.n122 B.n59 71.676
R522 B.n118 B.n58 71.676
R523 B.n114 B.n57 71.676
R524 B.n110 B.n56 71.676
R525 B.n106 B.n55 71.676
R526 B.n102 B.n54 71.676
R527 B.n98 B.n53 71.676
R528 B.n94 B.n52 71.676
R529 B.n89 B.n51 71.676
R530 B.n85 B.n50 71.676
R531 B.n81 B.n49 71.676
R532 B.n77 B.n48 71.676
R533 B.n73 B.n47 71.676
R534 B.n372 B.n46 71.676
R535 B.n269 B.n179 71.676
R536 B.n263 B.n180 71.676
R537 B.n259 B.n181 71.676
R538 B.n255 B.n182 71.676
R539 B.n251 B.n183 71.676
R540 B.n247 B.n184 71.676
R541 B.n243 B.n185 71.676
R542 B.n239 B.n186 71.676
R543 B.n235 B.n187 71.676
R544 B.n231 B.n188 71.676
R545 B.n226 B.n189 71.676
R546 B.n222 B.n190 71.676
R547 B.n218 B.n191 71.676
R548 B.n214 B.n192 71.676
R549 B.n210 B.n193 71.676
R550 B.n206 B.n194 71.676
R551 B.n202 B.n195 71.676
R552 B.n228 B.n201 59.5399
R553 B.n199 B.n198 59.5399
R554 B.n92 B.n69 59.5399
R555 B.n67 B.n66 59.5399
R556 B.n201 B.n200 48.4853
R557 B.n198 B.n197 48.4853
R558 B.n69 B.n68 48.4853
R559 B.n66 B.n65 48.4853
R560 B.n375 B.n374 30.1273
R561 B.n203 B.n174 30.1273
R562 B.n272 B.n271 30.1273
R563 B.n369 B.n368 30.1273
R564 B.t1 B.n140 28.1108
R565 B.n411 B.t0 28.1108
R566 B B.n422 18.0485
R567 B.n293 B.t7 16.2749
R568 B.n388 B.t3 16.2749
R569 B.n374 B.n45 10.6151
R570 B.n71 B.n45 10.6151
R571 B.n72 B.n71 10.6151
R572 B.n75 B.n72 10.6151
R573 B.n76 B.n75 10.6151
R574 B.n79 B.n76 10.6151
R575 B.n80 B.n79 10.6151
R576 B.n83 B.n80 10.6151
R577 B.n84 B.n83 10.6151
R578 B.n87 B.n84 10.6151
R579 B.n88 B.n87 10.6151
R580 B.n91 B.n88 10.6151
R581 B.n96 B.n93 10.6151
R582 B.n97 B.n96 10.6151
R583 B.n100 B.n97 10.6151
R584 B.n101 B.n100 10.6151
R585 B.n104 B.n101 10.6151
R586 B.n105 B.n104 10.6151
R587 B.n108 B.n105 10.6151
R588 B.n109 B.n108 10.6151
R589 B.n113 B.n112 10.6151
R590 B.n116 B.n113 10.6151
R591 B.n117 B.n116 10.6151
R592 B.n120 B.n117 10.6151
R593 B.n121 B.n120 10.6151
R594 B.n124 B.n121 10.6151
R595 B.n125 B.n124 10.6151
R596 B.n128 B.n125 10.6151
R597 B.n129 B.n128 10.6151
R598 B.n132 B.n129 10.6151
R599 B.n133 B.n132 10.6151
R600 B.n369 B.n133 10.6151
R601 B.n277 B.n174 10.6151
R602 B.n278 B.n277 10.6151
R603 B.n279 B.n278 10.6151
R604 B.n279 B.n166 10.6151
R605 B.n289 B.n166 10.6151
R606 B.n290 B.n289 10.6151
R607 B.n291 B.n290 10.6151
R608 B.n291 B.n158 10.6151
R609 B.n301 B.n158 10.6151
R610 B.n302 B.n301 10.6151
R611 B.n303 B.n302 10.6151
R612 B.n303 B.n150 10.6151
R613 B.n313 B.n150 10.6151
R614 B.n314 B.n313 10.6151
R615 B.n315 B.n314 10.6151
R616 B.n315 B.n142 10.6151
R617 B.n325 B.n142 10.6151
R618 B.n326 B.n325 10.6151
R619 B.n328 B.n326 10.6151
R620 B.n328 B.n327 10.6151
R621 B.n327 B.n134 10.6151
R622 B.n339 B.n134 10.6151
R623 B.n340 B.n339 10.6151
R624 B.n341 B.n340 10.6151
R625 B.n342 B.n341 10.6151
R626 B.n344 B.n342 10.6151
R627 B.n345 B.n344 10.6151
R628 B.n346 B.n345 10.6151
R629 B.n347 B.n346 10.6151
R630 B.n349 B.n347 10.6151
R631 B.n350 B.n349 10.6151
R632 B.n351 B.n350 10.6151
R633 B.n352 B.n351 10.6151
R634 B.n354 B.n352 10.6151
R635 B.n355 B.n354 10.6151
R636 B.n356 B.n355 10.6151
R637 B.n357 B.n356 10.6151
R638 B.n359 B.n357 10.6151
R639 B.n360 B.n359 10.6151
R640 B.n361 B.n360 10.6151
R641 B.n362 B.n361 10.6151
R642 B.n364 B.n362 10.6151
R643 B.n365 B.n364 10.6151
R644 B.n366 B.n365 10.6151
R645 B.n367 B.n366 10.6151
R646 B.n368 B.n367 10.6151
R647 B.n271 B.n178 10.6151
R648 B.n266 B.n178 10.6151
R649 B.n266 B.n265 10.6151
R650 B.n265 B.n264 10.6151
R651 B.n264 B.n261 10.6151
R652 B.n261 B.n260 10.6151
R653 B.n260 B.n257 10.6151
R654 B.n257 B.n256 10.6151
R655 B.n256 B.n253 10.6151
R656 B.n253 B.n252 10.6151
R657 B.n252 B.n249 10.6151
R658 B.n249 B.n248 10.6151
R659 B.n245 B.n244 10.6151
R660 B.n244 B.n241 10.6151
R661 B.n241 B.n240 10.6151
R662 B.n240 B.n237 10.6151
R663 B.n237 B.n236 10.6151
R664 B.n236 B.n233 10.6151
R665 B.n233 B.n232 10.6151
R666 B.n232 B.n229 10.6151
R667 B.n227 B.n224 10.6151
R668 B.n224 B.n223 10.6151
R669 B.n223 B.n220 10.6151
R670 B.n220 B.n219 10.6151
R671 B.n219 B.n216 10.6151
R672 B.n216 B.n215 10.6151
R673 B.n215 B.n212 10.6151
R674 B.n212 B.n211 10.6151
R675 B.n211 B.n208 10.6151
R676 B.n208 B.n207 10.6151
R677 B.n207 B.n204 10.6151
R678 B.n204 B.n203 10.6151
R679 B.n273 B.n272 10.6151
R680 B.n273 B.n170 10.6151
R681 B.n283 B.n170 10.6151
R682 B.n284 B.n283 10.6151
R683 B.n285 B.n284 10.6151
R684 B.n285 B.n162 10.6151
R685 B.n295 B.n162 10.6151
R686 B.n296 B.n295 10.6151
R687 B.n297 B.n296 10.6151
R688 B.n297 B.n154 10.6151
R689 B.n307 B.n154 10.6151
R690 B.n308 B.n307 10.6151
R691 B.n309 B.n308 10.6151
R692 B.n309 B.n146 10.6151
R693 B.n319 B.n146 10.6151
R694 B.n320 B.n319 10.6151
R695 B.n321 B.n320 10.6151
R696 B.n321 B.n138 10.6151
R697 B.n332 B.n138 10.6151
R698 B.n333 B.n332 10.6151
R699 B.n334 B.n333 10.6151
R700 B.n334 B.n0 10.6151
R701 B.n416 B.n1 10.6151
R702 B.n416 B.n415 10.6151
R703 B.n415 B.n414 10.6151
R704 B.n414 B.n10 10.6151
R705 B.n408 B.n10 10.6151
R706 B.n408 B.n407 10.6151
R707 B.n407 B.n406 10.6151
R708 B.n406 B.n17 10.6151
R709 B.n400 B.n17 10.6151
R710 B.n400 B.n399 10.6151
R711 B.n399 B.n398 10.6151
R712 B.n398 B.n24 10.6151
R713 B.n392 B.n24 10.6151
R714 B.n392 B.n391 10.6151
R715 B.n391 B.n390 10.6151
R716 B.n390 B.n31 10.6151
R717 B.n384 B.n31 10.6151
R718 B.n384 B.n383 10.6151
R719 B.n383 B.n382 10.6151
R720 B.n382 B.n38 10.6151
R721 B.n376 B.n38 10.6151
R722 B.n376 B.n375 10.6151
R723 B.n93 B.n92 6.5566
R724 B.n109 B.n67 6.5566
R725 B.n245 B.n199 6.5566
R726 B.n229 B.n228 6.5566
R727 B.n92 B.n91 4.05904
R728 B.n112 B.n67 4.05904
R729 B.n248 B.n199 4.05904
R730 B.n228 B.n227 4.05904
R731 B.n422 B.n0 2.81026
R732 B.n422 B.n1 2.81026
R733 VP.n0 VP.t0 109.266
R734 VP.n0 VP.t1 73.2045
R735 VP VP.n0 0.336784
R736 VTAIL.n3 VTAIL.t0 85.5676
R737 VTAIL.n0 VTAIL.t2 85.5676
R738 VTAIL.n2 VTAIL.t3 85.5676
R739 VTAIL.n1 VTAIL.t1 85.5675
R740 VTAIL.n1 VTAIL.n0 18.5393
R741 VTAIL.n3 VTAIL.n2 16.3841
R742 VTAIL.n2 VTAIL.n1 1.54791
R743 VTAIL VTAIL.n0 1.06731
R744 VTAIL VTAIL.n3 0.481103
R745 VDD1 VDD1.t0 133.142
R746 VDD1 VDD1.t1 102.844
R747 VN VN.t0 109.362
R748 VN VN.t1 73.5407
R749 VDD2.n0 VDD2.t0 132.078
R750 VDD2.n0 VDD2.t1 102.246
R751 VDD2 VDD2.n0 0.597483
C0 VDD2 VTAIL 2.3825f
C1 VN VDD1 0.154339f
C2 VN VP 3.43934f
C3 VDD1 VP 0.858044f
C4 VDD2 VN 0.692708f
C5 VDD2 VDD1 0.621979f
C6 VTAIL VN 0.90846f
C7 VDD2 VP 0.321247f
C8 VTAIL VDD1 2.33259f
C9 VTAIL VP 0.922607f
C10 VDD2 B 2.477676f
C11 VDD1 B 4.22168f
C12 VTAIL B 2.926331f
C13 VN B 7.044059f
C14 VP B 5.016919f
C15 VDD2.t0 B 0.425423f
C16 VDD2.t1 B 0.257409f
C17 VDD2.n0 B 1.62379f
C18 VN.t1 B 0.539718f
C19 VN.t0 B 0.914978f
C20 VDD1.t1 B 0.241326f
C21 VDD1.t0 B 0.412518f
C22 VTAIL.t2 B 0.274527f
C23 VTAIL.n0 B 0.940079f
C24 VTAIL.t1 B 0.274529f
C25 VTAIL.n1 B 0.971962f
C26 VTAIL.t3 B 0.274527f
C27 VTAIL.n2 B 0.828982f
C28 VTAIL.t0 B 0.274527f
C29 VTAIL.n3 B 0.758207f
C30 VP.t0 B 0.921557f
C31 VP.t1 B 0.545315f
C32 VP.n0 B 1.87432f
.ends

