* NGSPICE file created from diff_pair_sample_0014.ext - technology: sky130A

.subckt diff_pair_sample_0014 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=1.5951 ps=8.96 w=4.09 l=2.45
X1 VDD1.t8 VP.t1 VTAIL.t16 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0.67485 ps=4.42 w=4.09 l=2.45
X2 VDD1.t7 VP.t2 VTAIL.t12 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0.67485 ps=4.42 w=4.09 l=2.45
X3 VDD2.t9 VN.t0 VTAIL.t8 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0.67485 ps=4.42 w=4.09 l=2.45
X4 B.t11 B.t9 B.t10 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0 ps=0 w=4.09 l=2.45
X5 VDD2.t8 VN.t1 VTAIL.t1 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X6 VTAIL.t11 VP.t3 VDD1.t6 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X7 VDD2.t7 VN.t2 VTAIL.t0 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=1.5951 ps=8.96 w=4.09 l=2.45
X8 VDD2.t6 VN.t3 VTAIL.t7 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X9 VDD1.t5 VP.t4 VTAIL.t10 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=1.5951 ps=8.96 w=4.09 l=2.45
X10 VDD2.t5 VN.t4 VTAIL.t4 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=1.5951 ps=8.96 w=4.09 l=2.45
X11 B.t8 B.t6 B.t7 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0 ps=0 w=4.09 l=2.45
X12 VTAIL.t17 VP.t5 VDD1.t4 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X13 VTAIL.t3 VN.t5 VDD2.t4 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X14 VTAIL.t14 VP.t6 VDD1.t3 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X15 B.t5 B.t3 B.t4 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0 ps=0 w=4.09 l=2.45
X16 VTAIL.t9 VN.t6 VDD2.t3 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X17 VTAIL.t5 VN.t7 VDD2.t2 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X18 VDD1.t2 VP.t7 VTAIL.t13 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X19 VTAIL.t19 VP.t8 VDD1.t1 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X20 VTAIL.t6 VN.t8 VDD2.t1 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
X21 VDD2.t0 VN.t9 VTAIL.t2 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0.67485 ps=4.42 w=4.09 l=2.45
X22 B.t2 B.t0 B.t1 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=1.5951 pd=8.96 as=0 ps=0 w=4.09 l=2.45
X23 VDD1.t0 VP.t9 VTAIL.t18 w_n4306_n1786# sky130_fd_pr__pfet_01v8 ad=0.67485 pd=4.42 as=0.67485 ps=4.42 w=4.09 l=2.45
R0 VP.n23 VP.n20 161.3
R1 VP.n25 VP.n24 161.3
R2 VP.n26 VP.n19 161.3
R3 VP.n28 VP.n27 161.3
R4 VP.n29 VP.n18 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n17 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n36 VP.n16 161.3
R9 VP.n38 VP.n37 161.3
R10 VP.n39 VP.n15 161.3
R11 VP.n41 VP.n40 161.3
R12 VP.n43 VP.n14 161.3
R13 VP.n45 VP.n44 161.3
R14 VP.n46 VP.n13 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n49 VP.n12 161.3
R17 VP.n88 VP.n0 161.3
R18 VP.n87 VP.n86 161.3
R19 VP.n85 VP.n1 161.3
R20 VP.n84 VP.n83 161.3
R21 VP.n82 VP.n2 161.3
R22 VP.n80 VP.n79 161.3
R23 VP.n78 VP.n3 161.3
R24 VP.n77 VP.n76 161.3
R25 VP.n75 VP.n4 161.3
R26 VP.n74 VP.n73 161.3
R27 VP.n72 VP.n5 161.3
R28 VP.n71 VP.n70 161.3
R29 VP.n68 VP.n6 161.3
R30 VP.n67 VP.n66 161.3
R31 VP.n65 VP.n7 161.3
R32 VP.n64 VP.n63 161.3
R33 VP.n62 VP.n8 161.3
R34 VP.n60 VP.n59 161.3
R35 VP.n58 VP.n9 161.3
R36 VP.n57 VP.n56 161.3
R37 VP.n55 VP.n10 161.3
R38 VP.n54 VP.n53 161.3
R39 VP.n52 VP.n11 95.5869
R40 VP.n90 VP.n89 95.5869
R41 VP.n51 VP.n50 95.5869
R42 VP.n21 VP.t2 72.6457
R43 VP.n22 VP.n21 70.9722
R44 VP.n67 VP.n7 54.0911
R45 VP.n76 VP.n75 54.0911
R46 VP.n37 VP.n36 54.0911
R47 VP.n28 VP.n19 54.0911
R48 VP.n56 VP.n9 48.2635
R49 VP.n83 VP.n1 48.2635
R50 VP.n44 VP.n13 48.2635
R51 VP.n52 VP.n51 46.3708
R52 VP.n11 VP.t1 40.2327
R53 VP.n61 VP.t6 40.2327
R54 VP.n69 VP.t9 40.2327
R55 VP.n81 VP.t5 40.2327
R56 VP.n89 VP.t0 40.2327
R57 VP.n50 VP.t4 40.2327
R58 VP.n42 VP.t8 40.2327
R59 VP.n30 VP.t7 40.2327
R60 VP.n22 VP.t3 40.2327
R61 VP.n56 VP.n55 32.7233
R62 VP.n87 VP.n1 32.7233
R63 VP.n48 VP.n13 32.7233
R64 VP.n68 VP.n67 26.8957
R65 VP.n75 VP.n74 26.8957
R66 VP.n36 VP.n35 26.8957
R67 VP.n29 VP.n28 26.8957
R68 VP.n55 VP.n54 24.4675
R69 VP.n60 VP.n9 24.4675
R70 VP.n63 VP.n62 24.4675
R71 VP.n63 VP.n7 24.4675
R72 VP.n70 VP.n68 24.4675
R73 VP.n74 VP.n5 24.4675
R74 VP.n76 VP.n3 24.4675
R75 VP.n80 VP.n3 24.4675
R76 VP.n83 VP.n82 24.4675
R77 VP.n88 VP.n87 24.4675
R78 VP.n49 VP.n48 24.4675
R79 VP.n37 VP.n15 24.4675
R80 VP.n41 VP.n15 24.4675
R81 VP.n44 VP.n43 24.4675
R82 VP.n31 VP.n29 24.4675
R83 VP.n35 VP.n17 24.4675
R84 VP.n24 VP.n23 24.4675
R85 VP.n24 VP.n19 24.4675
R86 VP.n61 VP.n60 22.9995
R87 VP.n82 VP.n81 22.9995
R88 VP.n43 VP.n42 22.9995
R89 VP.n54 VP.n11 15.17
R90 VP.n89 VP.n88 15.17
R91 VP.n50 VP.n49 15.17
R92 VP.n70 VP.n69 12.234
R93 VP.n69 VP.n5 12.234
R94 VP.n31 VP.n30 12.234
R95 VP.n30 VP.n17 12.234
R96 VP.n21 VP.n20 9.50148
R97 VP.n62 VP.n61 1.46852
R98 VP.n81 VP.n80 1.46852
R99 VP.n42 VP.n41 1.46852
R100 VP.n23 VP.n22 1.46852
R101 VP.n51 VP.n12 0.278367
R102 VP.n53 VP.n52 0.278367
R103 VP.n90 VP.n0 0.278367
R104 VP.n25 VP.n20 0.189894
R105 VP.n26 VP.n25 0.189894
R106 VP.n27 VP.n26 0.189894
R107 VP.n27 VP.n18 0.189894
R108 VP.n32 VP.n18 0.189894
R109 VP.n33 VP.n32 0.189894
R110 VP.n34 VP.n33 0.189894
R111 VP.n34 VP.n16 0.189894
R112 VP.n38 VP.n16 0.189894
R113 VP.n39 VP.n38 0.189894
R114 VP.n40 VP.n39 0.189894
R115 VP.n40 VP.n14 0.189894
R116 VP.n45 VP.n14 0.189894
R117 VP.n46 VP.n45 0.189894
R118 VP.n47 VP.n46 0.189894
R119 VP.n47 VP.n12 0.189894
R120 VP.n53 VP.n10 0.189894
R121 VP.n57 VP.n10 0.189894
R122 VP.n58 VP.n57 0.189894
R123 VP.n59 VP.n58 0.189894
R124 VP.n59 VP.n8 0.189894
R125 VP.n64 VP.n8 0.189894
R126 VP.n65 VP.n64 0.189894
R127 VP.n66 VP.n65 0.189894
R128 VP.n66 VP.n6 0.189894
R129 VP.n71 VP.n6 0.189894
R130 VP.n72 VP.n71 0.189894
R131 VP.n73 VP.n72 0.189894
R132 VP.n73 VP.n4 0.189894
R133 VP.n77 VP.n4 0.189894
R134 VP.n78 VP.n77 0.189894
R135 VP.n79 VP.n78 0.189894
R136 VP.n79 VP.n2 0.189894
R137 VP.n84 VP.n2 0.189894
R138 VP.n85 VP.n84 0.189894
R139 VP.n86 VP.n85 0.189894
R140 VP.n86 VP.n0 0.189894
R141 VP VP.n90 0.153454
R142 VTAIL.n11 VTAIL.t4 97.5219
R143 VTAIL.n17 VTAIL.t0 97.5217
R144 VTAIL.n2 VTAIL.t15 97.5217
R145 VTAIL.n16 VTAIL.t10 97.5217
R146 VTAIL.n15 VTAIL.n14 89.5745
R147 VTAIL.n13 VTAIL.n12 89.5745
R148 VTAIL.n10 VTAIL.n9 89.5745
R149 VTAIL.n8 VTAIL.n7 89.5745
R150 VTAIL.n19 VTAIL.n18 89.5743
R151 VTAIL.n1 VTAIL.n0 89.5743
R152 VTAIL.n4 VTAIL.n3 89.5743
R153 VTAIL.n6 VTAIL.n5 89.5743
R154 VTAIL.n8 VTAIL.n6 20.6858
R155 VTAIL.n17 VTAIL.n16 18.2893
R156 VTAIL.n18 VTAIL.t1 7.94793
R157 VTAIL.n18 VTAIL.t9 7.94793
R158 VTAIL.n0 VTAIL.t8 7.94793
R159 VTAIL.n0 VTAIL.t3 7.94793
R160 VTAIL.n3 VTAIL.t18 7.94793
R161 VTAIL.n3 VTAIL.t17 7.94793
R162 VTAIL.n5 VTAIL.t16 7.94793
R163 VTAIL.n5 VTAIL.t14 7.94793
R164 VTAIL.n14 VTAIL.t13 7.94793
R165 VTAIL.n14 VTAIL.t19 7.94793
R166 VTAIL.n12 VTAIL.t12 7.94793
R167 VTAIL.n12 VTAIL.t11 7.94793
R168 VTAIL.n9 VTAIL.t7 7.94793
R169 VTAIL.n9 VTAIL.t5 7.94793
R170 VTAIL.n7 VTAIL.t2 7.94793
R171 VTAIL.n7 VTAIL.t6 7.94793
R172 VTAIL.n10 VTAIL.n8 2.39705
R173 VTAIL.n11 VTAIL.n10 2.39705
R174 VTAIL.n15 VTAIL.n13 2.39705
R175 VTAIL.n16 VTAIL.n15 2.39705
R176 VTAIL.n6 VTAIL.n4 2.39705
R177 VTAIL.n4 VTAIL.n2 2.39705
R178 VTAIL.n19 VTAIL.n17 2.39705
R179 VTAIL VTAIL.n1 1.8561
R180 VTAIL.n13 VTAIL.n11 1.6686
R181 VTAIL.n2 VTAIL.n1 1.6686
R182 VTAIL VTAIL.n19 0.541448
R183 VDD1.n1 VDD1.t7 116.597
R184 VDD1.n3 VDD1.t8 116.597
R185 VDD1.n5 VDD1.n4 107.996
R186 VDD1.n1 VDD1.n0 106.254
R187 VDD1.n7 VDD1.n6 106.254
R188 VDD1.n3 VDD1.n2 106.254
R189 VDD1.n7 VDD1.n5 40.4061
R190 VDD1.n6 VDD1.t1 7.94793
R191 VDD1.n6 VDD1.t5 7.94793
R192 VDD1.n0 VDD1.t6 7.94793
R193 VDD1.n0 VDD1.t2 7.94793
R194 VDD1.n4 VDD1.t4 7.94793
R195 VDD1.n4 VDD1.t9 7.94793
R196 VDD1.n2 VDD1.t3 7.94793
R197 VDD1.n2 VDD1.t0 7.94793
R198 VDD1 VDD1.n7 1.73972
R199 VDD1 VDD1.n1 0.657828
R200 VDD1.n5 VDD1.n3 0.544292
R201 VN.n77 VN.n40 161.3
R202 VN.n76 VN.n75 161.3
R203 VN.n74 VN.n41 161.3
R204 VN.n73 VN.n72 161.3
R205 VN.n71 VN.n42 161.3
R206 VN.n69 VN.n68 161.3
R207 VN.n67 VN.n43 161.3
R208 VN.n66 VN.n65 161.3
R209 VN.n64 VN.n44 161.3
R210 VN.n63 VN.n62 161.3
R211 VN.n61 VN.n45 161.3
R212 VN.n60 VN.n59 161.3
R213 VN.n58 VN.n46 161.3
R214 VN.n57 VN.n56 161.3
R215 VN.n55 VN.n48 161.3
R216 VN.n54 VN.n53 161.3
R217 VN.n52 VN.n49 161.3
R218 VN.n37 VN.n0 161.3
R219 VN.n36 VN.n35 161.3
R220 VN.n34 VN.n1 161.3
R221 VN.n33 VN.n32 161.3
R222 VN.n31 VN.n2 161.3
R223 VN.n29 VN.n28 161.3
R224 VN.n27 VN.n3 161.3
R225 VN.n26 VN.n25 161.3
R226 VN.n24 VN.n4 161.3
R227 VN.n23 VN.n22 161.3
R228 VN.n21 VN.n5 161.3
R229 VN.n20 VN.n19 161.3
R230 VN.n17 VN.n6 161.3
R231 VN.n16 VN.n15 161.3
R232 VN.n14 VN.n7 161.3
R233 VN.n13 VN.n12 161.3
R234 VN.n11 VN.n8 161.3
R235 VN.n39 VN.n38 95.5869
R236 VN.n79 VN.n78 95.5869
R237 VN.n9 VN.t0 72.6457
R238 VN.n50 VN.t4 72.6457
R239 VN.n10 VN.n9 70.9722
R240 VN.n51 VN.n50 70.9722
R241 VN.n16 VN.n7 54.0911
R242 VN.n25 VN.n24 54.0911
R243 VN.n57 VN.n48 54.0911
R244 VN.n65 VN.n64 54.0911
R245 VN.n32 VN.n1 48.2635
R246 VN.n72 VN.n41 48.2635
R247 VN VN.n79 46.6497
R248 VN.n10 VN.t5 40.2327
R249 VN.n18 VN.t1 40.2327
R250 VN.n30 VN.t6 40.2327
R251 VN.n38 VN.t2 40.2327
R252 VN.n51 VN.t7 40.2327
R253 VN.n47 VN.t3 40.2327
R254 VN.n70 VN.t8 40.2327
R255 VN.n78 VN.t9 40.2327
R256 VN.n36 VN.n1 32.7233
R257 VN.n76 VN.n41 32.7233
R258 VN.n17 VN.n16 26.8957
R259 VN.n24 VN.n23 26.8957
R260 VN.n58 VN.n57 26.8957
R261 VN.n64 VN.n63 26.8957
R262 VN.n12 VN.n11 24.4675
R263 VN.n12 VN.n7 24.4675
R264 VN.n19 VN.n17 24.4675
R265 VN.n23 VN.n5 24.4675
R266 VN.n25 VN.n3 24.4675
R267 VN.n29 VN.n3 24.4675
R268 VN.n32 VN.n31 24.4675
R269 VN.n37 VN.n36 24.4675
R270 VN.n53 VN.n48 24.4675
R271 VN.n53 VN.n52 24.4675
R272 VN.n63 VN.n45 24.4675
R273 VN.n59 VN.n58 24.4675
R274 VN.n72 VN.n71 24.4675
R275 VN.n69 VN.n43 24.4675
R276 VN.n65 VN.n43 24.4675
R277 VN.n77 VN.n76 24.4675
R278 VN.n31 VN.n30 22.9995
R279 VN.n71 VN.n70 22.9995
R280 VN.n38 VN.n37 15.17
R281 VN.n78 VN.n77 15.17
R282 VN.n19 VN.n18 12.234
R283 VN.n18 VN.n5 12.234
R284 VN.n47 VN.n45 12.234
R285 VN.n59 VN.n47 12.234
R286 VN.n50 VN.n49 9.50148
R287 VN.n9 VN.n8 9.50148
R288 VN.n11 VN.n10 1.46852
R289 VN.n30 VN.n29 1.46852
R290 VN.n52 VN.n51 1.46852
R291 VN.n70 VN.n69 1.46852
R292 VN.n79 VN.n40 0.278367
R293 VN.n39 VN.n0 0.278367
R294 VN.n75 VN.n40 0.189894
R295 VN.n75 VN.n74 0.189894
R296 VN.n74 VN.n73 0.189894
R297 VN.n73 VN.n42 0.189894
R298 VN.n68 VN.n42 0.189894
R299 VN.n68 VN.n67 0.189894
R300 VN.n67 VN.n66 0.189894
R301 VN.n66 VN.n44 0.189894
R302 VN.n62 VN.n44 0.189894
R303 VN.n62 VN.n61 0.189894
R304 VN.n61 VN.n60 0.189894
R305 VN.n60 VN.n46 0.189894
R306 VN.n56 VN.n46 0.189894
R307 VN.n56 VN.n55 0.189894
R308 VN.n55 VN.n54 0.189894
R309 VN.n54 VN.n49 0.189894
R310 VN.n13 VN.n8 0.189894
R311 VN.n14 VN.n13 0.189894
R312 VN.n15 VN.n14 0.189894
R313 VN.n15 VN.n6 0.189894
R314 VN.n20 VN.n6 0.189894
R315 VN.n21 VN.n20 0.189894
R316 VN.n22 VN.n21 0.189894
R317 VN.n22 VN.n4 0.189894
R318 VN.n26 VN.n4 0.189894
R319 VN.n27 VN.n26 0.189894
R320 VN.n28 VN.n27 0.189894
R321 VN.n28 VN.n2 0.189894
R322 VN.n33 VN.n2 0.189894
R323 VN.n34 VN.n33 0.189894
R324 VN.n35 VN.n34 0.189894
R325 VN.n35 VN.n0 0.189894
R326 VN VN.n39 0.153454
R327 VDD2.n1 VDD2.t9 116.597
R328 VDD2.n4 VDD2.t0 114.201
R329 VDD2.n3 VDD2.n2 107.996
R330 VDD2 VDD2.n7 107.993
R331 VDD2.n6 VDD2.n5 106.254
R332 VDD2.n1 VDD2.n0 106.254
R333 VDD2.n4 VDD2.n3 38.6248
R334 VDD2.n7 VDD2.t2 7.94793
R335 VDD2.n7 VDD2.t5 7.94793
R336 VDD2.n5 VDD2.t1 7.94793
R337 VDD2.n5 VDD2.t6 7.94793
R338 VDD2.n2 VDD2.t3 7.94793
R339 VDD2.n2 VDD2.t7 7.94793
R340 VDD2.n0 VDD2.t4 7.94793
R341 VDD2.n0 VDD2.t8 7.94793
R342 VDD2.n6 VDD2.n4 2.39705
R343 VDD2 VDD2.n6 0.657828
R344 VDD2.n3 VDD2.n1 0.544292
R345 B.n499 B.n58 585
R346 B.n501 B.n500 585
R347 B.n502 B.n57 585
R348 B.n504 B.n503 585
R349 B.n505 B.n56 585
R350 B.n507 B.n506 585
R351 B.n508 B.n55 585
R352 B.n510 B.n509 585
R353 B.n511 B.n54 585
R354 B.n513 B.n512 585
R355 B.n514 B.n53 585
R356 B.n516 B.n515 585
R357 B.n517 B.n52 585
R358 B.n519 B.n518 585
R359 B.n520 B.n51 585
R360 B.n522 B.n521 585
R361 B.n523 B.n47 585
R362 B.n525 B.n524 585
R363 B.n526 B.n46 585
R364 B.n528 B.n527 585
R365 B.n529 B.n45 585
R366 B.n531 B.n530 585
R367 B.n532 B.n44 585
R368 B.n534 B.n533 585
R369 B.n535 B.n43 585
R370 B.n537 B.n536 585
R371 B.n538 B.n42 585
R372 B.n540 B.n539 585
R373 B.n542 B.n39 585
R374 B.n544 B.n543 585
R375 B.n545 B.n38 585
R376 B.n547 B.n546 585
R377 B.n548 B.n37 585
R378 B.n550 B.n549 585
R379 B.n551 B.n36 585
R380 B.n553 B.n552 585
R381 B.n554 B.n35 585
R382 B.n556 B.n555 585
R383 B.n557 B.n34 585
R384 B.n559 B.n558 585
R385 B.n560 B.n33 585
R386 B.n562 B.n561 585
R387 B.n563 B.n32 585
R388 B.n565 B.n564 585
R389 B.n566 B.n31 585
R390 B.n568 B.n567 585
R391 B.n498 B.n497 585
R392 B.n496 B.n59 585
R393 B.n495 B.n494 585
R394 B.n493 B.n60 585
R395 B.n492 B.n491 585
R396 B.n490 B.n61 585
R397 B.n489 B.n488 585
R398 B.n487 B.n62 585
R399 B.n486 B.n485 585
R400 B.n484 B.n63 585
R401 B.n483 B.n482 585
R402 B.n481 B.n64 585
R403 B.n480 B.n479 585
R404 B.n478 B.n65 585
R405 B.n477 B.n476 585
R406 B.n475 B.n66 585
R407 B.n474 B.n473 585
R408 B.n472 B.n67 585
R409 B.n471 B.n470 585
R410 B.n469 B.n68 585
R411 B.n468 B.n467 585
R412 B.n466 B.n69 585
R413 B.n465 B.n464 585
R414 B.n463 B.n70 585
R415 B.n462 B.n461 585
R416 B.n460 B.n71 585
R417 B.n459 B.n458 585
R418 B.n457 B.n72 585
R419 B.n456 B.n455 585
R420 B.n454 B.n73 585
R421 B.n453 B.n452 585
R422 B.n451 B.n74 585
R423 B.n450 B.n449 585
R424 B.n448 B.n75 585
R425 B.n447 B.n446 585
R426 B.n445 B.n76 585
R427 B.n444 B.n443 585
R428 B.n442 B.n77 585
R429 B.n441 B.n440 585
R430 B.n439 B.n78 585
R431 B.n438 B.n437 585
R432 B.n436 B.n79 585
R433 B.n435 B.n434 585
R434 B.n433 B.n80 585
R435 B.n432 B.n431 585
R436 B.n430 B.n81 585
R437 B.n429 B.n428 585
R438 B.n427 B.n82 585
R439 B.n426 B.n425 585
R440 B.n424 B.n83 585
R441 B.n423 B.n422 585
R442 B.n421 B.n84 585
R443 B.n420 B.n419 585
R444 B.n418 B.n85 585
R445 B.n417 B.n416 585
R446 B.n415 B.n86 585
R447 B.n414 B.n413 585
R448 B.n412 B.n87 585
R449 B.n411 B.n410 585
R450 B.n409 B.n88 585
R451 B.n408 B.n407 585
R452 B.n406 B.n89 585
R453 B.n405 B.n404 585
R454 B.n403 B.n90 585
R455 B.n402 B.n401 585
R456 B.n400 B.n91 585
R457 B.n399 B.n398 585
R458 B.n397 B.n92 585
R459 B.n396 B.n395 585
R460 B.n394 B.n93 585
R461 B.n393 B.n392 585
R462 B.n391 B.n94 585
R463 B.n390 B.n389 585
R464 B.n388 B.n95 585
R465 B.n387 B.n386 585
R466 B.n385 B.n96 585
R467 B.n384 B.n383 585
R468 B.n382 B.n97 585
R469 B.n381 B.n380 585
R470 B.n379 B.n98 585
R471 B.n378 B.n377 585
R472 B.n376 B.n99 585
R473 B.n375 B.n374 585
R474 B.n373 B.n100 585
R475 B.n372 B.n371 585
R476 B.n370 B.n101 585
R477 B.n369 B.n368 585
R478 B.n367 B.n102 585
R479 B.n366 B.n365 585
R480 B.n364 B.n103 585
R481 B.n363 B.n362 585
R482 B.n361 B.n104 585
R483 B.n360 B.n359 585
R484 B.n358 B.n105 585
R485 B.n357 B.n356 585
R486 B.n355 B.n106 585
R487 B.n354 B.n353 585
R488 B.n352 B.n107 585
R489 B.n351 B.n350 585
R490 B.n349 B.n108 585
R491 B.n348 B.n347 585
R492 B.n346 B.n109 585
R493 B.n345 B.n344 585
R494 B.n343 B.n110 585
R495 B.n342 B.n341 585
R496 B.n340 B.n111 585
R497 B.n339 B.n338 585
R498 B.n337 B.n112 585
R499 B.n336 B.n335 585
R500 B.n334 B.n113 585
R501 B.n333 B.n332 585
R502 B.n331 B.n114 585
R503 B.n330 B.n329 585
R504 B.n328 B.n115 585
R505 B.n327 B.n326 585
R506 B.n256 B.n143 585
R507 B.n258 B.n257 585
R508 B.n259 B.n142 585
R509 B.n261 B.n260 585
R510 B.n262 B.n141 585
R511 B.n264 B.n263 585
R512 B.n265 B.n140 585
R513 B.n267 B.n266 585
R514 B.n268 B.n139 585
R515 B.n270 B.n269 585
R516 B.n271 B.n138 585
R517 B.n273 B.n272 585
R518 B.n274 B.n137 585
R519 B.n276 B.n275 585
R520 B.n277 B.n136 585
R521 B.n279 B.n278 585
R522 B.n280 B.n135 585
R523 B.n282 B.n281 585
R524 B.n284 B.n132 585
R525 B.n286 B.n285 585
R526 B.n287 B.n131 585
R527 B.n289 B.n288 585
R528 B.n290 B.n130 585
R529 B.n292 B.n291 585
R530 B.n293 B.n129 585
R531 B.n295 B.n294 585
R532 B.n296 B.n128 585
R533 B.n298 B.n297 585
R534 B.n300 B.n299 585
R535 B.n301 B.n124 585
R536 B.n303 B.n302 585
R537 B.n304 B.n123 585
R538 B.n306 B.n305 585
R539 B.n307 B.n122 585
R540 B.n309 B.n308 585
R541 B.n310 B.n121 585
R542 B.n312 B.n311 585
R543 B.n313 B.n120 585
R544 B.n315 B.n314 585
R545 B.n316 B.n119 585
R546 B.n318 B.n317 585
R547 B.n319 B.n118 585
R548 B.n321 B.n320 585
R549 B.n322 B.n117 585
R550 B.n324 B.n323 585
R551 B.n325 B.n116 585
R552 B.n255 B.n254 585
R553 B.n253 B.n144 585
R554 B.n252 B.n251 585
R555 B.n250 B.n145 585
R556 B.n249 B.n248 585
R557 B.n247 B.n146 585
R558 B.n246 B.n245 585
R559 B.n244 B.n147 585
R560 B.n243 B.n242 585
R561 B.n241 B.n148 585
R562 B.n240 B.n239 585
R563 B.n238 B.n149 585
R564 B.n237 B.n236 585
R565 B.n235 B.n150 585
R566 B.n234 B.n233 585
R567 B.n232 B.n151 585
R568 B.n231 B.n230 585
R569 B.n229 B.n152 585
R570 B.n228 B.n227 585
R571 B.n226 B.n153 585
R572 B.n225 B.n224 585
R573 B.n223 B.n154 585
R574 B.n222 B.n221 585
R575 B.n220 B.n155 585
R576 B.n219 B.n218 585
R577 B.n217 B.n156 585
R578 B.n216 B.n215 585
R579 B.n214 B.n157 585
R580 B.n213 B.n212 585
R581 B.n211 B.n158 585
R582 B.n210 B.n209 585
R583 B.n208 B.n159 585
R584 B.n207 B.n206 585
R585 B.n205 B.n160 585
R586 B.n204 B.n203 585
R587 B.n202 B.n161 585
R588 B.n201 B.n200 585
R589 B.n199 B.n162 585
R590 B.n198 B.n197 585
R591 B.n196 B.n163 585
R592 B.n195 B.n194 585
R593 B.n193 B.n164 585
R594 B.n192 B.n191 585
R595 B.n190 B.n165 585
R596 B.n189 B.n188 585
R597 B.n187 B.n166 585
R598 B.n186 B.n185 585
R599 B.n184 B.n167 585
R600 B.n183 B.n182 585
R601 B.n181 B.n168 585
R602 B.n180 B.n179 585
R603 B.n178 B.n169 585
R604 B.n177 B.n176 585
R605 B.n175 B.n170 585
R606 B.n174 B.n173 585
R607 B.n172 B.n171 585
R608 B.n2 B.n0 585
R609 B.n653 B.n1 585
R610 B.n652 B.n651 585
R611 B.n650 B.n3 585
R612 B.n649 B.n648 585
R613 B.n647 B.n4 585
R614 B.n646 B.n645 585
R615 B.n644 B.n5 585
R616 B.n643 B.n642 585
R617 B.n641 B.n6 585
R618 B.n640 B.n639 585
R619 B.n638 B.n7 585
R620 B.n637 B.n636 585
R621 B.n635 B.n8 585
R622 B.n634 B.n633 585
R623 B.n632 B.n9 585
R624 B.n631 B.n630 585
R625 B.n629 B.n10 585
R626 B.n628 B.n627 585
R627 B.n626 B.n11 585
R628 B.n625 B.n624 585
R629 B.n623 B.n12 585
R630 B.n622 B.n621 585
R631 B.n620 B.n13 585
R632 B.n619 B.n618 585
R633 B.n617 B.n14 585
R634 B.n616 B.n615 585
R635 B.n614 B.n15 585
R636 B.n613 B.n612 585
R637 B.n611 B.n16 585
R638 B.n610 B.n609 585
R639 B.n608 B.n17 585
R640 B.n607 B.n606 585
R641 B.n605 B.n18 585
R642 B.n604 B.n603 585
R643 B.n602 B.n19 585
R644 B.n601 B.n600 585
R645 B.n599 B.n20 585
R646 B.n598 B.n597 585
R647 B.n596 B.n21 585
R648 B.n595 B.n594 585
R649 B.n593 B.n22 585
R650 B.n592 B.n591 585
R651 B.n590 B.n23 585
R652 B.n589 B.n588 585
R653 B.n587 B.n24 585
R654 B.n586 B.n585 585
R655 B.n584 B.n25 585
R656 B.n583 B.n582 585
R657 B.n581 B.n26 585
R658 B.n580 B.n579 585
R659 B.n578 B.n27 585
R660 B.n577 B.n576 585
R661 B.n575 B.n28 585
R662 B.n574 B.n573 585
R663 B.n572 B.n29 585
R664 B.n571 B.n570 585
R665 B.n569 B.n30 585
R666 B.n655 B.n654 585
R667 B.n256 B.n255 550.159
R668 B.n569 B.n568 550.159
R669 B.n327 B.n116 550.159
R670 B.n497 B.n58 550.159
R671 B.n125 B.t6 248.042
R672 B.n133 B.t3 248.042
R673 B.n40 B.t9 248.042
R674 B.n48 B.t0 248.042
R675 B.n125 B.t8 173.18
R676 B.n48 B.t1 173.18
R677 B.n133 B.t5 173.177
R678 B.n40 B.t10 173.177
R679 B.n255 B.n144 163.367
R680 B.n251 B.n144 163.367
R681 B.n251 B.n250 163.367
R682 B.n250 B.n249 163.367
R683 B.n249 B.n146 163.367
R684 B.n245 B.n146 163.367
R685 B.n245 B.n244 163.367
R686 B.n244 B.n243 163.367
R687 B.n243 B.n148 163.367
R688 B.n239 B.n148 163.367
R689 B.n239 B.n238 163.367
R690 B.n238 B.n237 163.367
R691 B.n237 B.n150 163.367
R692 B.n233 B.n150 163.367
R693 B.n233 B.n232 163.367
R694 B.n232 B.n231 163.367
R695 B.n231 B.n152 163.367
R696 B.n227 B.n152 163.367
R697 B.n227 B.n226 163.367
R698 B.n226 B.n225 163.367
R699 B.n225 B.n154 163.367
R700 B.n221 B.n154 163.367
R701 B.n221 B.n220 163.367
R702 B.n220 B.n219 163.367
R703 B.n219 B.n156 163.367
R704 B.n215 B.n156 163.367
R705 B.n215 B.n214 163.367
R706 B.n214 B.n213 163.367
R707 B.n213 B.n158 163.367
R708 B.n209 B.n158 163.367
R709 B.n209 B.n208 163.367
R710 B.n208 B.n207 163.367
R711 B.n207 B.n160 163.367
R712 B.n203 B.n160 163.367
R713 B.n203 B.n202 163.367
R714 B.n202 B.n201 163.367
R715 B.n201 B.n162 163.367
R716 B.n197 B.n162 163.367
R717 B.n197 B.n196 163.367
R718 B.n196 B.n195 163.367
R719 B.n195 B.n164 163.367
R720 B.n191 B.n164 163.367
R721 B.n191 B.n190 163.367
R722 B.n190 B.n189 163.367
R723 B.n189 B.n166 163.367
R724 B.n185 B.n166 163.367
R725 B.n185 B.n184 163.367
R726 B.n184 B.n183 163.367
R727 B.n183 B.n168 163.367
R728 B.n179 B.n168 163.367
R729 B.n179 B.n178 163.367
R730 B.n178 B.n177 163.367
R731 B.n177 B.n170 163.367
R732 B.n173 B.n170 163.367
R733 B.n173 B.n172 163.367
R734 B.n172 B.n2 163.367
R735 B.n654 B.n2 163.367
R736 B.n654 B.n653 163.367
R737 B.n653 B.n652 163.367
R738 B.n652 B.n3 163.367
R739 B.n648 B.n3 163.367
R740 B.n648 B.n647 163.367
R741 B.n647 B.n646 163.367
R742 B.n646 B.n5 163.367
R743 B.n642 B.n5 163.367
R744 B.n642 B.n641 163.367
R745 B.n641 B.n640 163.367
R746 B.n640 B.n7 163.367
R747 B.n636 B.n7 163.367
R748 B.n636 B.n635 163.367
R749 B.n635 B.n634 163.367
R750 B.n634 B.n9 163.367
R751 B.n630 B.n9 163.367
R752 B.n630 B.n629 163.367
R753 B.n629 B.n628 163.367
R754 B.n628 B.n11 163.367
R755 B.n624 B.n11 163.367
R756 B.n624 B.n623 163.367
R757 B.n623 B.n622 163.367
R758 B.n622 B.n13 163.367
R759 B.n618 B.n13 163.367
R760 B.n618 B.n617 163.367
R761 B.n617 B.n616 163.367
R762 B.n616 B.n15 163.367
R763 B.n612 B.n15 163.367
R764 B.n612 B.n611 163.367
R765 B.n611 B.n610 163.367
R766 B.n610 B.n17 163.367
R767 B.n606 B.n17 163.367
R768 B.n606 B.n605 163.367
R769 B.n605 B.n604 163.367
R770 B.n604 B.n19 163.367
R771 B.n600 B.n19 163.367
R772 B.n600 B.n599 163.367
R773 B.n599 B.n598 163.367
R774 B.n598 B.n21 163.367
R775 B.n594 B.n21 163.367
R776 B.n594 B.n593 163.367
R777 B.n593 B.n592 163.367
R778 B.n592 B.n23 163.367
R779 B.n588 B.n23 163.367
R780 B.n588 B.n587 163.367
R781 B.n587 B.n586 163.367
R782 B.n586 B.n25 163.367
R783 B.n582 B.n25 163.367
R784 B.n582 B.n581 163.367
R785 B.n581 B.n580 163.367
R786 B.n580 B.n27 163.367
R787 B.n576 B.n27 163.367
R788 B.n576 B.n575 163.367
R789 B.n575 B.n574 163.367
R790 B.n574 B.n29 163.367
R791 B.n570 B.n29 163.367
R792 B.n570 B.n569 163.367
R793 B.n257 B.n256 163.367
R794 B.n257 B.n142 163.367
R795 B.n261 B.n142 163.367
R796 B.n262 B.n261 163.367
R797 B.n263 B.n262 163.367
R798 B.n263 B.n140 163.367
R799 B.n267 B.n140 163.367
R800 B.n268 B.n267 163.367
R801 B.n269 B.n268 163.367
R802 B.n269 B.n138 163.367
R803 B.n273 B.n138 163.367
R804 B.n274 B.n273 163.367
R805 B.n275 B.n274 163.367
R806 B.n275 B.n136 163.367
R807 B.n279 B.n136 163.367
R808 B.n280 B.n279 163.367
R809 B.n281 B.n280 163.367
R810 B.n281 B.n132 163.367
R811 B.n286 B.n132 163.367
R812 B.n287 B.n286 163.367
R813 B.n288 B.n287 163.367
R814 B.n288 B.n130 163.367
R815 B.n292 B.n130 163.367
R816 B.n293 B.n292 163.367
R817 B.n294 B.n293 163.367
R818 B.n294 B.n128 163.367
R819 B.n298 B.n128 163.367
R820 B.n299 B.n298 163.367
R821 B.n299 B.n124 163.367
R822 B.n303 B.n124 163.367
R823 B.n304 B.n303 163.367
R824 B.n305 B.n304 163.367
R825 B.n305 B.n122 163.367
R826 B.n309 B.n122 163.367
R827 B.n310 B.n309 163.367
R828 B.n311 B.n310 163.367
R829 B.n311 B.n120 163.367
R830 B.n315 B.n120 163.367
R831 B.n316 B.n315 163.367
R832 B.n317 B.n316 163.367
R833 B.n317 B.n118 163.367
R834 B.n321 B.n118 163.367
R835 B.n322 B.n321 163.367
R836 B.n323 B.n322 163.367
R837 B.n323 B.n116 163.367
R838 B.n328 B.n327 163.367
R839 B.n329 B.n328 163.367
R840 B.n329 B.n114 163.367
R841 B.n333 B.n114 163.367
R842 B.n334 B.n333 163.367
R843 B.n335 B.n334 163.367
R844 B.n335 B.n112 163.367
R845 B.n339 B.n112 163.367
R846 B.n340 B.n339 163.367
R847 B.n341 B.n340 163.367
R848 B.n341 B.n110 163.367
R849 B.n345 B.n110 163.367
R850 B.n346 B.n345 163.367
R851 B.n347 B.n346 163.367
R852 B.n347 B.n108 163.367
R853 B.n351 B.n108 163.367
R854 B.n352 B.n351 163.367
R855 B.n353 B.n352 163.367
R856 B.n353 B.n106 163.367
R857 B.n357 B.n106 163.367
R858 B.n358 B.n357 163.367
R859 B.n359 B.n358 163.367
R860 B.n359 B.n104 163.367
R861 B.n363 B.n104 163.367
R862 B.n364 B.n363 163.367
R863 B.n365 B.n364 163.367
R864 B.n365 B.n102 163.367
R865 B.n369 B.n102 163.367
R866 B.n370 B.n369 163.367
R867 B.n371 B.n370 163.367
R868 B.n371 B.n100 163.367
R869 B.n375 B.n100 163.367
R870 B.n376 B.n375 163.367
R871 B.n377 B.n376 163.367
R872 B.n377 B.n98 163.367
R873 B.n381 B.n98 163.367
R874 B.n382 B.n381 163.367
R875 B.n383 B.n382 163.367
R876 B.n383 B.n96 163.367
R877 B.n387 B.n96 163.367
R878 B.n388 B.n387 163.367
R879 B.n389 B.n388 163.367
R880 B.n389 B.n94 163.367
R881 B.n393 B.n94 163.367
R882 B.n394 B.n393 163.367
R883 B.n395 B.n394 163.367
R884 B.n395 B.n92 163.367
R885 B.n399 B.n92 163.367
R886 B.n400 B.n399 163.367
R887 B.n401 B.n400 163.367
R888 B.n401 B.n90 163.367
R889 B.n405 B.n90 163.367
R890 B.n406 B.n405 163.367
R891 B.n407 B.n406 163.367
R892 B.n407 B.n88 163.367
R893 B.n411 B.n88 163.367
R894 B.n412 B.n411 163.367
R895 B.n413 B.n412 163.367
R896 B.n413 B.n86 163.367
R897 B.n417 B.n86 163.367
R898 B.n418 B.n417 163.367
R899 B.n419 B.n418 163.367
R900 B.n419 B.n84 163.367
R901 B.n423 B.n84 163.367
R902 B.n424 B.n423 163.367
R903 B.n425 B.n424 163.367
R904 B.n425 B.n82 163.367
R905 B.n429 B.n82 163.367
R906 B.n430 B.n429 163.367
R907 B.n431 B.n430 163.367
R908 B.n431 B.n80 163.367
R909 B.n435 B.n80 163.367
R910 B.n436 B.n435 163.367
R911 B.n437 B.n436 163.367
R912 B.n437 B.n78 163.367
R913 B.n441 B.n78 163.367
R914 B.n442 B.n441 163.367
R915 B.n443 B.n442 163.367
R916 B.n443 B.n76 163.367
R917 B.n447 B.n76 163.367
R918 B.n448 B.n447 163.367
R919 B.n449 B.n448 163.367
R920 B.n449 B.n74 163.367
R921 B.n453 B.n74 163.367
R922 B.n454 B.n453 163.367
R923 B.n455 B.n454 163.367
R924 B.n455 B.n72 163.367
R925 B.n459 B.n72 163.367
R926 B.n460 B.n459 163.367
R927 B.n461 B.n460 163.367
R928 B.n461 B.n70 163.367
R929 B.n465 B.n70 163.367
R930 B.n466 B.n465 163.367
R931 B.n467 B.n466 163.367
R932 B.n467 B.n68 163.367
R933 B.n471 B.n68 163.367
R934 B.n472 B.n471 163.367
R935 B.n473 B.n472 163.367
R936 B.n473 B.n66 163.367
R937 B.n477 B.n66 163.367
R938 B.n478 B.n477 163.367
R939 B.n479 B.n478 163.367
R940 B.n479 B.n64 163.367
R941 B.n483 B.n64 163.367
R942 B.n484 B.n483 163.367
R943 B.n485 B.n484 163.367
R944 B.n485 B.n62 163.367
R945 B.n489 B.n62 163.367
R946 B.n490 B.n489 163.367
R947 B.n491 B.n490 163.367
R948 B.n491 B.n60 163.367
R949 B.n495 B.n60 163.367
R950 B.n496 B.n495 163.367
R951 B.n497 B.n496 163.367
R952 B.n568 B.n31 163.367
R953 B.n564 B.n31 163.367
R954 B.n564 B.n563 163.367
R955 B.n563 B.n562 163.367
R956 B.n562 B.n33 163.367
R957 B.n558 B.n33 163.367
R958 B.n558 B.n557 163.367
R959 B.n557 B.n556 163.367
R960 B.n556 B.n35 163.367
R961 B.n552 B.n35 163.367
R962 B.n552 B.n551 163.367
R963 B.n551 B.n550 163.367
R964 B.n550 B.n37 163.367
R965 B.n546 B.n37 163.367
R966 B.n546 B.n545 163.367
R967 B.n545 B.n544 163.367
R968 B.n544 B.n39 163.367
R969 B.n539 B.n39 163.367
R970 B.n539 B.n538 163.367
R971 B.n538 B.n537 163.367
R972 B.n537 B.n43 163.367
R973 B.n533 B.n43 163.367
R974 B.n533 B.n532 163.367
R975 B.n532 B.n531 163.367
R976 B.n531 B.n45 163.367
R977 B.n527 B.n45 163.367
R978 B.n527 B.n526 163.367
R979 B.n526 B.n525 163.367
R980 B.n525 B.n47 163.367
R981 B.n521 B.n47 163.367
R982 B.n521 B.n520 163.367
R983 B.n520 B.n519 163.367
R984 B.n519 B.n52 163.367
R985 B.n515 B.n52 163.367
R986 B.n515 B.n514 163.367
R987 B.n514 B.n513 163.367
R988 B.n513 B.n54 163.367
R989 B.n509 B.n54 163.367
R990 B.n509 B.n508 163.367
R991 B.n508 B.n507 163.367
R992 B.n507 B.n56 163.367
R993 B.n503 B.n56 163.367
R994 B.n503 B.n502 163.367
R995 B.n502 B.n501 163.367
R996 B.n501 B.n58 163.367
R997 B.n126 B.t7 119.266
R998 B.n49 B.t2 119.266
R999 B.n134 B.t4 119.261
R1000 B.n41 B.t11 119.261
R1001 B.n127 B.n126 59.5399
R1002 B.n283 B.n134 59.5399
R1003 B.n541 B.n41 59.5399
R1004 B.n50 B.n49 59.5399
R1005 B.n126 B.n125 53.9157
R1006 B.n134 B.n133 53.9157
R1007 B.n41 B.n40 53.9157
R1008 B.n49 B.n48 53.9157
R1009 B.n567 B.n30 35.7468
R1010 B.n499 B.n498 35.7468
R1011 B.n326 B.n325 35.7468
R1012 B.n254 B.n143 35.7468
R1013 B B.n655 18.0485
R1014 B.n567 B.n566 10.6151
R1015 B.n566 B.n565 10.6151
R1016 B.n565 B.n32 10.6151
R1017 B.n561 B.n32 10.6151
R1018 B.n561 B.n560 10.6151
R1019 B.n560 B.n559 10.6151
R1020 B.n559 B.n34 10.6151
R1021 B.n555 B.n34 10.6151
R1022 B.n555 B.n554 10.6151
R1023 B.n554 B.n553 10.6151
R1024 B.n553 B.n36 10.6151
R1025 B.n549 B.n36 10.6151
R1026 B.n549 B.n548 10.6151
R1027 B.n548 B.n547 10.6151
R1028 B.n547 B.n38 10.6151
R1029 B.n543 B.n38 10.6151
R1030 B.n543 B.n542 10.6151
R1031 B.n540 B.n42 10.6151
R1032 B.n536 B.n42 10.6151
R1033 B.n536 B.n535 10.6151
R1034 B.n535 B.n534 10.6151
R1035 B.n534 B.n44 10.6151
R1036 B.n530 B.n44 10.6151
R1037 B.n530 B.n529 10.6151
R1038 B.n529 B.n528 10.6151
R1039 B.n528 B.n46 10.6151
R1040 B.n524 B.n523 10.6151
R1041 B.n523 B.n522 10.6151
R1042 B.n522 B.n51 10.6151
R1043 B.n518 B.n51 10.6151
R1044 B.n518 B.n517 10.6151
R1045 B.n517 B.n516 10.6151
R1046 B.n516 B.n53 10.6151
R1047 B.n512 B.n53 10.6151
R1048 B.n512 B.n511 10.6151
R1049 B.n511 B.n510 10.6151
R1050 B.n510 B.n55 10.6151
R1051 B.n506 B.n55 10.6151
R1052 B.n506 B.n505 10.6151
R1053 B.n505 B.n504 10.6151
R1054 B.n504 B.n57 10.6151
R1055 B.n500 B.n57 10.6151
R1056 B.n500 B.n499 10.6151
R1057 B.n326 B.n115 10.6151
R1058 B.n330 B.n115 10.6151
R1059 B.n331 B.n330 10.6151
R1060 B.n332 B.n331 10.6151
R1061 B.n332 B.n113 10.6151
R1062 B.n336 B.n113 10.6151
R1063 B.n337 B.n336 10.6151
R1064 B.n338 B.n337 10.6151
R1065 B.n338 B.n111 10.6151
R1066 B.n342 B.n111 10.6151
R1067 B.n343 B.n342 10.6151
R1068 B.n344 B.n343 10.6151
R1069 B.n344 B.n109 10.6151
R1070 B.n348 B.n109 10.6151
R1071 B.n349 B.n348 10.6151
R1072 B.n350 B.n349 10.6151
R1073 B.n350 B.n107 10.6151
R1074 B.n354 B.n107 10.6151
R1075 B.n355 B.n354 10.6151
R1076 B.n356 B.n355 10.6151
R1077 B.n356 B.n105 10.6151
R1078 B.n360 B.n105 10.6151
R1079 B.n361 B.n360 10.6151
R1080 B.n362 B.n361 10.6151
R1081 B.n362 B.n103 10.6151
R1082 B.n366 B.n103 10.6151
R1083 B.n367 B.n366 10.6151
R1084 B.n368 B.n367 10.6151
R1085 B.n368 B.n101 10.6151
R1086 B.n372 B.n101 10.6151
R1087 B.n373 B.n372 10.6151
R1088 B.n374 B.n373 10.6151
R1089 B.n374 B.n99 10.6151
R1090 B.n378 B.n99 10.6151
R1091 B.n379 B.n378 10.6151
R1092 B.n380 B.n379 10.6151
R1093 B.n380 B.n97 10.6151
R1094 B.n384 B.n97 10.6151
R1095 B.n385 B.n384 10.6151
R1096 B.n386 B.n385 10.6151
R1097 B.n386 B.n95 10.6151
R1098 B.n390 B.n95 10.6151
R1099 B.n391 B.n390 10.6151
R1100 B.n392 B.n391 10.6151
R1101 B.n392 B.n93 10.6151
R1102 B.n396 B.n93 10.6151
R1103 B.n397 B.n396 10.6151
R1104 B.n398 B.n397 10.6151
R1105 B.n398 B.n91 10.6151
R1106 B.n402 B.n91 10.6151
R1107 B.n403 B.n402 10.6151
R1108 B.n404 B.n403 10.6151
R1109 B.n404 B.n89 10.6151
R1110 B.n408 B.n89 10.6151
R1111 B.n409 B.n408 10.6151
R1112 B.n410 B.n409 10.6151
R1113 B.n410 B.n87 10.6151
R1114 B.n414 B.n87 10.6151
R1115 B.n415 B.n414 10.6151
R1116 B.n416 B.n415 10.6151
R1117 B.n416 B.n85 10.6151
R1118 B.n420 B.n85 10.6151
R1119 B.n421 B.n420 10.6151
R1120 B.n422 B.n421 10.6151
R1121 B.n422 B.n83 10.6151
R1122 B.n426 B.n83 10.6151
R1123 B.n427 B.n426 10.6151
R1124 B.n428 B.n427 10.6151
R1125 B.n428 B.n81 10.6151
R1126 B.n432 B.n81 10.6151
R1127 B.n433 B.n432 10.6151
R1128 B.n434 B.n433 10.6151
R1129 B.n434 B.n79 10.6151
R1130 B.n438 B.n79 10.6151
R1131 B.n439 B.n438 10.6151
R1132 B.n440 B.n439 10.6151
R1133 B.n440 B.n77 10.6151
R1134 B.n444 B.n77 10.6151
R1135 B.n445 B.n444 10.6151
R1136 B.n446 B.n445 10.6151
R1137 B.n446 B.n75 10.6151
R1138 B.n450 B.n75 10.6151
R1139 B.n451 B.n450 10.6151
R1140 B.n452 B.n451 10.6151
R1141 B.n452 B.n73 10.6151
R1142 B.n456 B.n73 10.6151
R1143 B.n457 B.n456 10.6151
R1144 B.n458 B.n457 10.6151
R1145 B.n458 B.n71 10.6151
R1146 B.n462 B.n71 10.6151
R1147 B.n463 B.n462 10.6151
R1148 B.n464 B.n463 10.6151
R1149 B.n464 B.n69 10.6151
R1150 B.n468 B.n69 10.6151
R1151 B.n469 B.n468 10.6151
R1152 B.n470 B.n469 10.6151
R1153 B.n470 B.n67 10.6151
R1154 B.n474 B.n67 10.6151
R1155 B.n475 B.n474 10.6151
R1156 B.n476 B.n475 10.6151
R1157 B.n476 B.n65 10.6151
R1158 B.n480 B.n65 10.6151
R1159 B.n481 B.n480 10.6151
R1160 B.n482 B.n481 10.6151
R1161 B.n482 B.n63 10.6151
R1162 B.n486 B.n63 10.6151
R1163 B.n487 B.n486 10.6151
R1164 B.n488 B.n487 10.6151
R1165 B.n488 B.n61 10.6151
R1166 B.n492 B.n61 10.6151
R1167 B.n493 B.n492 10.6151
R1168 B.n494 B.n493 10.6151
R1169 B.n494 B.n59 10.6151
R1170 B.n498 B.n59 10.6151
R1171 B.n258 B.n143 10.6151
R1172 B.n259 B.n258 10.6151
R1173 B.n260 B.n259 10.6151
R1174 B.n260 B.n141 10.6151
R1175 B.n264 B.n141 10.6151
R1176 B.n265 B.n264 10.6151
R1177 B.n266 B.n265 10.6151
R1178 B.n266 B.n139 10.6151
R1179 B.n270 B.n139 10.6151
R1180 B.n271 B.n270 10.6151
R1181 B.n272 B.n271 10.6151
R1182 B.n272 B.n137 10.6151
R1183 B.n276 B.n137 10.6151
R1184 B.n277 B.n276 10.6151
R1185 B.n278 B.n277 10.6151
R1186 B.n278 B.n135 10.6151
R1187 B.n282 B.n135 10.6151
R1188 B.n285 B.n284 10.6151
R1189 B.n285 B.n131 10.6151
R1190 B.n289 B.n131 10.6151
R1191 B.n290 B.n289 10.6151
R1192 B.n291 B.n290 10.6151
R1193 B.n291 B.n129 10.6151
R1194 B.n295 B.n129 10.6151
R1195 B.n296 B.n295 10.6151
R1196 B.n297 B.n296 10.6151
R1197 B.n301 B.n300 10.6151
R1198 B.n302 B.n301 10.6151
R1199 B.n302 B.n123 10.6151
R1200 B.n306 B.n123 10.6151
R1201 B.n307 B.n306 10.6151
R1202 B.n308 B.n307 10.6151
R1203 B.n308 B.n121 10.6151
R1204 B.n312 B.n121 10.6151
R1205 B.n313 B.n312 10.6151
R1206 B.n314 B.n313 10.6151
R1207 B.n314 B.n119 10.6151
R1208 B.n318 B.n119 10.6151
R1209 B.n319 B.n318 10.6151
R1210 B.n320 B.n319 10.6151
R1211 B.n320 B.n117 10.6151
R1212 B.n324 B.n117 10.6151
R1213 B.n325 B.n324 10.6151
R1214 B.n254 B.n253 10.6151
R1215 B.n253 B.n252 10.6151
R1216 B.n252 B.n145 10.6151
R1217 B.n248 B.n145 10.6151
R1218 B.n248 B.n247 10.6151
R1219 B.n247 B.n246 10.6151
R1220 B.n246 B.n147 10.6151
R1221 B.n242 B.n147 10.6151
R1222 B.n242 B.n241 10.6151
R1223 B.n241 B.n240 10.6151
R1224 B.n240 B.n149 10.6151
R1225 B.n236 B.n149 10.6151
R1226 B.n236 B.n235 10.6151
R1227 B.n235 B.n234 10.6151
R1228 B.n234 B.n151 10.6151
R1229 B.n230 B.n151 10.6151
R1230 B.n230 B.n229 10.6151
R1231 B.n229 B.n228 10.6151
R1232 B.n228 B.n153 10.6151
R1233 B.n224 B.n153 10.6151
R1234 B.n224 B.n223 10.6151
R1235 B.n223 B.n222 10.6151
R1236 B.n222 B.n155 10.6151
R1237 B.n218 B.n155 10.6151
R1238 B.n218 B.n217 10.6151
R1239 B.n217 B.n216 10.6151
R1240 B.n216 B.n157 10.6151
R1241 B.n212 B.n157 10.6151
R1242 B.n212 B.n211 10.6151
R1243 B.n211 B.n210 10.6151
R1244 B.n210 B.n159 10.6151
R1245 B.n206 B.n159 10.6151
R1246 B.n206 B.n205 10.6151
R1247 B.n205 B.n204 10.6151
R1248 B.n204 B.n161 10.6151
R1249 B.n200 B.n161 10.6151
R1250 B.n200 B.n199 10.6151
R1251 B.n199 B.n198 10.6151
R1252 B.n198 B.n163 10.6151
R1253 B.n194 B.n163 10.6151
R1254 B.n194 B.n193 10.6151
R1255 B.n193 B.n192 10.6151
R1256 B.n192 B.n165 10.6151
R1257 B.n188 B.n165 10.6151
R1258 B.n188 B.n187 10.6151
R1259 B.n187 B.n186 10.6151
R1260 B.n186 B.n167 10.6151
R1261 B.n182 B.n167 10.6151
R1262 B.n182 B.n181 10.6151
R1263 B.n181 B.n180 10.6151
R1264 B.n180 B.n169 10.6151
R1265 B.n176 B.n169 10.6151
R1266 B.n176 B.n175 10.6151
R1267 B.n175 B.n174 10.6151
R1268 B.n174 B.n171 10.6151
R1269 B.n171 B.n0 10.6151
R1270 B.n651 B.n1 10.6151
R1271 B.n651 B.n650 10.6151
R1272 B.n650 B.n649 10.6151
R1273 B.n649 B.n4 10.6151
R1274 B.n645 B.n4 10.6151
R1275 B.n645 B.n644 10.6151
R1276 B.n644 B.n643 10.6151
R1277 B.n643 B.n6 10.6151
R1278 B.n639 B.n6 10.6151
R1279 B.n639 B.n638 10.6151
R1280 B.n638 B.n637 10.6151
R1281 B.n637 B.n8 10.6151
R1282 B.n633 B.n8 10.6151
R1283 B.n633 B.n632 10.6151
R1284 B.n632 B.n631 10.6151
R1285 B.n631 B.n10 10.6151
R1286 B.n627 B.n10 10.6151
R1287 B.n627 B.n626 10.6151
R1288 B.n626 B.n625 10.6151
R1289 B.n625 B.n12 10.6151
R1290 B.n621 B.n12 10.6151
R1291 B.n621 B.n620 10.6151
R1292 B.n620 B.n619 10.6151
R1293 B.n619 B.n14 10.6151
R1294 B.n615 B.n14 10.6151
R1295 B.n615 B.n614 10.6151
R1296 B.n614 B.n613 10.6151
R1297 B.n613 B.n16 10.6151
R1298 B.n609 B.n16 10.6151
R1299 B.n609 B.n608 10.6151
R1300 B.n608 B.n607 10.6151
R1301 B.n607 B.n18 10.6151
R1302 B.n603 B.n18 10.6151
R1303 B.n603 B.n602 10.6151
R1304 B.n602 B.n601 10.6151
R1305 B.n601 B.n20 10.6151
R1306 B.n597 B.n20 10.6151
R1307 B.n597 B.n596 10.6151
R1308 B.n596 B.n595 10.6151
R1309 B.n595 B.n22 10.6151
R1310 B.n591 B.n22 10.6151
R1311 B.n591 B.n590 10.6151
R1312 B.n590 B.n589 10.6151
R1313 B.n589 B.n24 10.6151
R1314 B.n585 B.n24 10.6151
R1315 B.n585 B.n584 10.6151
R1316 B.n584 B.n583 10.6151
R1317 B.n583 B.n26 10.6151
R1318 B.n579 B.n26 10.6151
R1319 B.n579 B.n578 10.6151
R1320 B.n578 B.n577 10.6151
R1321 B.n577 B.n28 10.6151
R1322 B.n573 B.n28 10.6151
R1323 B.n573 B.n572 10.6151
R1324 B.n572 B.n571 10.6151
R1325 B.n571 B.n30 10.6151
R1326 B.n542 B.n541 9.36635
R1327 B.n524 B.n50 9.36635
R1328 B.n283 B.n282 9.36635
R1329 B.n300 B.n127 9.36635
R1330 B.n655 B.n0 2.81026
R1331 B.n655 B.n1 2.81026
R1332 B.n541 B.n540 1.24928
R1333 B.n50 B.n46 1.24928
R1334 B.n284 B.n283 1.24928
R1335 B.n297 B.n127 1.24928
C0 B VN 1.18606f
C1 VDD2 VN 3.93236f
C2 VDD1 VN 0.157224f
C3 w_n4306_n1786# VN 9.024651f
C4 VDD2 B 1.91031f
C5 B VDD1 1.7981f
C6 VDD2 VDD1 2.07543f
C7 VTAIL VN 5.084681f
C8 B w_n4306_n1786# 8.09682f
C9 VDD2 w_n4306_n1786# 2.31396f
C10 w_n4306_n1786# VDD1 2.17851f
C11 VP VN 6.71579f
C12 VTAIL B 1.88093f
C13 VTAIL VDD2 6.66542f
C14 VTAIL VDD1 6.6137f
C15 VP B 2.12698f
C16 VDD2 VP 0.568614f
C17 VP VDD1 4.34057f
C18 VTAIL w_n4306_n1786# 2.06274f
C19 VP w_n4306_n1786# 9.58404f
C20 VTAIL VP 5.09885f
C21 VDD2 VSUBS 1.842804f
C22 VDD1 VSUBS 1.677882f
C23 VTAIL VSUBS 0.594388f
C24 VN VSUBS 7.17451f
C25 VP VSUBS 3.469129f
C26 B VSUBS 4.246393f
C27 w_n4306_n1786# VSUBS 96.7817f
C28 B.n0 VSUBS 0.005483f
C29 B.n1 VSUBS 0.005483f
C30 B.n2 VSUBS 0.008671f
C31 B.n3 VSUBS 0.008671f
C32 B.n4 VSUBS 0.008671f
C33 B.n5 VSUBS 0.008671f
C34 B.n6 VSUBS 0.008671f
C35 B.n7 VSUBS 0.008671f
C36 B.n8 VSUBS 0.008671f
C37 B.n9 VSUBS 0.008671f
C38 B.n10 VSUBS 0.008671f
C39 B.n11 VSUBS 0.008671f
C40 B.n12 VSUBS 0.008671f
C41 B.n13 VSUBS 0.008671f
C42 B.n14 VSUBS 0.008671f
C43 B.n15 VSUBS 0.008671f
C44 B.n16 VSUBS 0.008671f
C45 B.n17 VSUBS 0.008671f
C46 B.n18 VSUBS 0.008671f
C47 B.n19 VSUBS 0.008671f
C48 B.n20 VSUBS 0.008671f
C49 B.n21 VSUBS 0.008671f
C50 B.n22 VSUBS 0.008671f
C51 B.n23 VSUBS 0.008671f
C52 B.n24 VSUBS 0.008671f
C53 B.n25 VSUBS 0.008671f
C54 B.n26 VSUBS 0.008671f
C55 B.n27 VSUBS 0.008671f
C56 B.n28 VSUBS 0.008671f
C57 B.n29 VSUBS 0.008671f
C58 B.n30 VSUBS 0.021081f
C59 B.n31 VSUBS 0.008671f
C60 B.n32 VSUBS 0.008671f
C61 B.n33 VSUBS 0.008671f
C62 B.n34 VSUBS 0.008671f
C63 B.n35 VSUBS 0.008671f
C64 B.n36 VSUBS 0.008671f
C65 B.n37 VSUBS 0.008671f
C66 B.n38 VSUBS 0.008671f
C67 B.n39 VSUBS 0.008671f
C68 B.t11 VSUBS 0.134223f
C69 B.t10 VSUBS 0.156555f
C70 B.t9 VSUBS 0.595391f
C71 B.n40 VSUBS 0.11259f
C72 B.n41 VSUBS 0.084096f
C73 B.n42 VSUBS 0.008671f
C74 B.n43 VSUBS 0.008671f
C75 B.n44 VSUBS 0.008671f
C76 B.n45 VSUBS 0.008671f
C77 B.n46 VSUBS 0.004845f
C78 B.n47 VSUBS 0.008671f
C79 B.t2 VSUBS 0.134223f
C80 B.t1 VSUBS 0.156554f
C81 B.t0 VSUBS 0.595391f
C82 B.n48 VSUBS 0.112591f
C83 B.n49 VSUBS 0.084096f
C84 B.n50 VSUBS 0.020089f
C85 B.n51 VSUBS 0.008671f
C86 B.n52 VSUBS 0.008671f
C87 B.n53 VSUBS 0.008671f
C88 B.n54 VSUBS 0.008671f
C89 B.n55 VSUBS 0.008671f
C90 B.n56 VSUBS 0.008671f
C91 B.n57 VSUBS 0.008671f
C92 B.n58 VSUBS 0.022017f
C93 B.n59 VSUBS 0.008671f
C94 B.n60 VSUBS 0.008671f
C95 B.n61 VSUBS 0.008671f
C96 B.n62 VSUBS 0.008671f
C97 B.n63 VSUBS 0.008671f
C98 B.n64 VSUBS 0.008671f
C99 B.n65 VSUBS 0.008671f
C100 B.n66 VSUBS 0.008671f
C101 B.n67 VSUBS 0.008671f
C102 B.n68 VSUBS 0.008671f
C103 B.n69 VSUBS 0.008671f
C104 B.n70 VSUBS 0.008671f
C105 B.n71 VSUBS 0.008671f
C106 B.n72 VSUBS 0.008671f
C107 B.n73 VSUBS 0.008671f
C108 B.n74 VSUBS 0.008671f
C109 B.n75 VSUBS 0.008671f
C110 B.n76 VSUBS 0.008671f
C111 B.n77 VSUBS 0.008671f
C112 B.n78 VSUBS 0.008671f
C113 B.n79 VSUBS 0.008671f
C114 B.n80 VSUBS 0.008671f
C115 B.n81 VSUBS 0.008671f
C116 B.n82 VSUBS 0.008671f
C117 B.n83 VSUBS 0.008671f
C118 B.n84 VSUBS 0.008671f
C119 B.n85 VSUBS 0.008671f
C120 B.n86 VSUBS 0.008671f
C121 B.n87 VSUBS 0.008671f
C122 B.n88 VSUBS 0.008671f
C123 B.n89 VSUBS 0.008671f
C124 B.n90 VSUBS 0.008671f
C125 B.n91 VSUBS 0.008671f
C126 B.n92 VSUBS 0.008671f
C127 B.n93 VSUBS 0.008671f
C128 B.n94 VSUBS 0.008671f
C129 B.n95 VSUBS 0.008671f
C130 B.n96 VSUBS 0.008671f
C131 B.n97 VSUBS 0.008671f
C132 B.n98 VSUBS 0.008671f
C133 B.n99 VSUBS 0.008671f
C134 B.n100 VSUBS 0.008671f
C135 B.n101 VSUBS 0.008671f
C136 B.n102 VSUBS 0.008671f
C137 B.n103 VSUBS 0.008671f
C138 B.n104 VSUBS 0.008671f
C139 B.n105 VSUBS 0.008671f
C140 B.n106 VSUBS 0.008671f
C141 B.n107 VSUBS 0.008671f
C142 B.n108 VSUBS 0.008671f
C143 B.n109 VSUBS 0.008671f
C144 B.n110 VSUBS 0.008671f
C145 B.n111 VSUBS 0.008671f
C146 B.n112 VSUBS 0.008671f
C147 B.n113 VSUBS 0.008671f
C148 B.n114 VSUBS 0.008671f
C149 B.n115 VSUBS 0.008671f
C150 B.n116 VSUBS 0.022017f
C151 B.n117 VSUBS 0.008671f
C152 B.n118 VSUBS 0.008671f
C153 B.n119 VSUBS 0.008671f
C154 B.n120 VSUBS 0.008671f
C155 B.n121 VSUBS 0.008671f
C156 B.n122 VSUBS 0.008671f
C157 B.n123 VSUBS 0.008671f
C158 B.n124 VSUBS 0.008671f
C159 B.t7 VSUBS 0.134223f
C160 B.t8 VSUBS 0.156554f
C161 B.t6 VSUBS 0.595391f
C162 B.n125 VSUBS 0.112591f
C163 B.n126 VSUBS 0.084096f
C164 B.n127 VSUBS 0.020089f
C165 B.n128 VSUBS 0.008671f
C166 B.n129 VSUBS 0.008671f
C167 B.n130 VSUBS 0.008671f
C168 B.n131 VSUBS 0.008671f
C169 B.n132 VSUBS 0.008671f
C170 B.t4 VSUBS 0.134223f
C171 B.t5 VSUBS 0.156555f
C172 B.t3 VSUBS 0.595391f
C173 B.n133 VSUBS 0.11259f
C174 B.n134 VSUBS 0.084096f
C175 B.n135 VSUBS 0.008671f
C176 B.n136 VSUBS 0.008671f
C177 B.n137 VSUBS 0.008671f
C178 B.n138 VSUBS 0.008671f
C179 B.n139 VSUBS 0.008671f
C180 B.n140 VSUBS 0.008671f
C181 B.n141 VSUBS 0.008671f
C182 B.n142 VSUBS 0.008671f
C183 B.n143 VSUBS 0.022017f
C184 B.n144 VSUBS 0.008671f
C185 B.n145 VSUBS 0.008671f
C186 B.n146 VSUBS 0.008671f
C187 B.n147 VSUBS 0.008671f
C188 B.n148 VSUBS 0.008671f
C189 B.n149 VSUBS 0.008671f
C190 B.n150 VSUBS 0.008671f
C191 B.n151 VSUBS 0.008671f
C192 B.n152 VSUBS 0.008671f
C193 B.n153 VSUBS 0.008671f
C194 B.n154 VSUBS 0.008671f
C195 B.n155 VSUBS 0.008671f
C196 B.n156 VSUBS 0.008671f
C197 B.n157 VSUBS 0.008671f
C198 B.n158 VSUBS 0.008671f
C199 B.n159 VSUBS 0.008671f
C200 B.n160 VSUBS 0.008671f
C201 B.n161 VSUBS 0.008671f
C202 B.n162 VSUBS 0.008671f
C203 B.n163 VSUBS 0.008671f
C204 B.n164 VSUBS 0.008671f
C205 B.n165 VSUBS 0.008671f
C206 B.n166 VSUBS 0.008671f
C207 B.n167 VSUBS 0.008671f
C208 B.n168 VSUBS 0.008671f
C209 B.n169 VSUBS 0.008671f
C210 B.n170 VSUBS 0.008671f
C211 B.n171 VSUBS 0.008671f
C212 B.n172 VSUBS 0.008671f
C213 B.n173 VSUBS 0.008671f
C214 B.n174 VSUBS 0.008671f
C215 B.n175 VSUBS 0.008671f
C216 B.n176 VSUBS 0.008671f
C217 B.n177 VSUBS 0.008671f
C218 B.n178 VSUBS 0.008671f
C219 B.n179 VSUBS 0.008671f
C220 B.n180 VSUBS 0.008671f
C221 B.n181 VSUBS 0.008671f
C222 B.n182 VSUBS 0.008671f
C223 B.n183 VSUBS 0.008671f
C224 B.n184 VSUBS 0.008671f
C225 B.n185 VSUBS 0.008671f
C226 B.n186 VSUBS 0.008671f
C227 B.n187 VSUBS 0.008671f
C228 B.n188 VSUBS 0.008671f
C229 B.n189 VSUBS 0.008671f
C230 B.n190 VSUBS 0.008671f
C231 B.n191 VSUBS 0.008671f
C232 B.n192 VSUBS 0.008671f
C233 B.n193 VSUBS 0.008671f
C234 B.n194 VSUBS 0.008671f
C235 B.n195 VSUBS 0.008671f
C236 B.n196 VSUBS 0.008671f
C237 B.n197 VSUBS 0.008671f
C238 B.n198 VSUBS 0.008671f
C239 B.n199 VSUBS 0.008671f
C240 B.n200 VSUBS 0.008671f
C241 B.n201 VSUBS 0.008671f
C242 B.n202 VSUBS 0.008671f
C243 B.n203 VSUBS 0.008671f
C244 B.n204 VSUBS 0.008671f
C245 B.n205 VSUBS 0.008671f
C246 B.n206 VSUBS 0.008671f
C247 B.n207 VSUBS 0.008671f
C248 B.n208 VSUBS 0.008671f
C249 B.n209 VSUBS 0.008671f
C250 B.n210 VSUBS 0.008671f
C251 B.n211 VSUBS 0.008671f
C252 B.n212 VSUBS 0.008671f
C253 B.n213 VSUBS 0.008671f
C254 B.n214 VSUBS 0.008671f
C255 B.n215 VSUBS 0.008671f
C256 B.n216 VSUBS 0.008671f
C257 B.n217 VSUBS 0.008671f
C258 B.n218 VSUBS 0.008671f
C259 B.n219 VSUBS 0.008671f
C260 B.n220 VSUBS 0.008671f
C261 B.n221 VSUBS 0.008671f
C262 B.n222 VSUBS 0.008671f
C263 B.n223 VSUBS 0.008671f
C264 B.n224 VSUBS 0.008671f
C265 B.n225 VSUBS 0.008671f
C266 B.n226 VSUBS 0.008671f
C267 B.n227 VSUBS 0.008671f
C268 B.n228 VSUBS 0.008671f
C269 B.n229 VSUBS 0.008671f
C270 B.n230 VSUBS 0.008671f
C271 B.n231 VSUBS 0.008671f
C272 B.n232 VSUBS 0.008671f
C273 B.n233 VSUBS 0.008671f
C274 B.n234 VSUBS 0.008671f
C275 B.n235 VSUBS 0.008671f
C276 B.n236 VSUBS 0.008671f
C277 B.n237 VSUBS 0.008671f
C278 B.n238 VSUBS 0.008671f
C279 B.n239 VSUBS 0.008671f
C280 B.n240 VSUBS 0.008671f
C281 B.n241 VSUBS 0.008671f
C282 B.n242 VSUBS 0.008671f
C283 B.n243 VSUBS 0.008671f
C284 B.n244 VSUBS 0.008671f
C285 B.n245 VSUBS 0.008671f
C286 B.n246 VSUBS 0.008671f
C287 B.n247 VSUBS 0.008671f
C288 B.n248 VSUBS 0.008671f
C289 B.n249 VSUBS 0.008671f
C290 B.n250 VSUBS 0.008671f
C291 B.n251 VSUBS 0.008671f
C292 B.n252 VSUBS 0.008671f
C293 B.n253 VSUBS 0.008671f
C294 B.n254 VSUBS 0.021081f
C295 B.n255 VSUBS 0.021081f
C296 B.n256 VSUBS 0.022017f
C297 B.n257 VSUBS 0.008671f
C298 B.n258 VSUBS 0.008671f
C299 B.n259 VSUBS 0.008671f
C300 B.n260 VSUBS 0.008671f
C301 B.n261 VSUBS 0.008671f
C302 B.n262 VSUBS 0.008671f
C303 B.n263 VSUBS 0.008671f
C304 B.n264 VSUBS 0.008671f
C305 B.n265 VSUBS 0.008671f
C306 B.n266 VSUBS 0.008671f
C307 B.n267 VSUBS 0.008671f
C308 B.n268 VSUBS 0.008671f
C309 B.n269 VSUBS 0.008671f
C310 B.n270 VSUBS 0.008671f
C311 B.n271 VSUBS 0.008671f
C312 B.n272 VSUBS 0.008671f
C313 B.n273 VSUBS 0.008671f
C314 B.n274 VSUBS 0.008671f
C315 B.n275 VSUBS 0.008671f
C316 B.n276 VSUBS 0.008671f
C317 B.n277 VSUBS 0.008671f
C318 B.n278 VSUBS 0.008671f
C319 B.n279 VSUBS 0.008671f
C320 B.n280 VSUBS 0.008671f
C321 B.n281 VSUBS 0.008671f
C322 B.n282 VSUBS 0.008161f
C323 B.n283 VSUBS 0.020089f
C324 B.n284 VSUBS 0.004845f
C325 B.n285 VSUBS 0.008671f
C326 B.n286 VSUBS 0.008671f
C327 B.n287 VSUBS 0.008671f
C328 B.n288 VSUBS 0.008671f
C329 B.n289 VSUBS 0.008671f
C330 B.n290 VSUBS 0.008671f
C331 B.n291 VSUBS 0.008671f
C332 B.n292 VSUBS 0.008671f
C333 B.n293 VSUBS 0.008671f
C334 B.n294 VSUBS 0.008671f
C335 B.n295 VSUBS 0.008671f
C336 B.n296 VSUBS 0.008671f
C337 B.n297 VSUBS 0.004845f
C338 B.n298 VSUBS 0.008671f
C339 B.n299 VSUBS 0.008671f
C340 B.n300 VSUBS 0.008161f
C341 B.n301 VSUBS 0.008671f
C342 B.n302 VSUBS 0.008671f
C343 B.n303 VSUBS 0.008671f
C344 B.n304 VSUBS 0.008671f
C345 B.n305 VSUBS 0.008671f
C346 B.n306 VSUBS 0.008671f
C347 B.n307 VSUBS 0.008671f
C348 B.n308 VSUBS 0.008671f
C349 B.n309 VSUBS 0.008671f
C350 B.n310 VSUBS 0.008671f
C351 B.n311 VSUBS 0.008671f
C352 B.n312 VSUBS 0.008671f
C353 B.n313 VSUBS 0.008671f
C354 B.n314 VSUBS 0.008671f
C355 B.n315 VSUBS 0.008671f
C356 B.n316 VSUBS 0.008671f
C357 B.n317 VSUBS 0.008671f
C358 B.n318 VSUBS 0.008671f
C359 B.n319 VSUBS 0.008671f
C360 B.n320 VSUBS 0.008671f
C361 B.n321 VSUBS 0.008671f
C362 B.n322 VSUBS 0.008671f
C363 B.n323 VSUBS 0.008671f
C364 B.n324 VSUBS 0.008671f
C365 B.n325 VSUBS 0.022017f
C366 B.n326 VSUBS 0.021081f
C367 B.n327 VSUBS 0.021081f
C368 B.n328 VSUBS 0.008671f
C369 B.n329 VSUBS 0.008671f
C370 B.n330 VSUBS 0.008671f
C371 B.n331 VSUBS 0.008671f
C372 B.n332 VSUBS 0.008671f
C373 B.n333 VSUBS 0.008671f
C374 B.n334 VSUBS 0.008671f
C375 B.n335 VSUBS 0.008671f
C376 B.n336 VSUBS 0.008671f
C377 B.n337 VSUBS 0.008671f
C378 B.n338 VSUBS 0.008671f
C379 B.n339 VSUBS 0.008671f
C380 B.n340 VSUBS 0.008671f
C381 B.n341 VSUBS 0.008671f
C382 B.n342 VSUBS 0.008671f
C383 B.n343 VSUBS 0.008671f
C384 B.n344 VSUBS 0.008671f
C385 B.n345 VSUBS 0.008671f
C386 B.n346 VSUBS 0.008671f
C387 B.n347 VSUBS 0.008671f
C388 B.n348 VSUBS 0.008671f
C389 B.n349 VSUBS 0.008671f
C390 B.n350 VSUBS 0.008671f
C391 B.n351 VSUBS 0.008671f
C392 B.n352 VSUBS 0.008671f
C393 B.n353 VSUBS 0.008671f
C394 B.n354 VSUBS 0.008671f
C395 B.n355 VSUBS 0.008671f
C396 B.n356 VSUBS 0.008671f
C397 B.n357 VSUBS 0.008671f
C398 B.n358 VSUBS 0.008671f
C399 B.n359 VSUBS 0.008671f
C400 B.n360 VSUBS 0.008671f
C401 B.n361 VSUBS 0.008671f
C402 B.n362 VSUBS 0.008671f
C403 B.n363 VSUBS 0.008671f
C404 B.n364 VSUBS 0.008671f
C405 B.n365 VSUBS 0.008671f
C406 B.n366 VSUBS 0.008671f
C407 B.n367 VSUBS 0.008671f
C408 B.n368 VSUBS 0.008671f
C409 B.n369 VSUBS 0.008671f
C410 B.n370 VSUBS 0.008671f
C411 B.n371 VSUBS 0.008671f
C412 B.n372 VSUBS 0.008671f
C413 B.n373 VSUBS 0.008671f
C414 B.n374 VSUBS 0.008671f
C415 B.n375 VSUBS 0.008671f
C416 B.n376 VSUBS 0.008671f
C417 B.n377 VSUBS 0.008671f
C418 B.n378 VSUBS 0.008671f
C419 B.n379 VSUBS 0.008671f
C420 B.n380 VSUBS 0.008671f
C421 B.n381 VSUBS 0.008671f
C422 B.n382 VSUBS 0.008671f
C423 B.n383 VSUBS 0.008671f
C424 B.n384 VSUBS 0.008671f
C425 B.n385 VSUBS 0.008671f
C426 B.n386 VSUBS 0.008671f
C427 B.n387 VSUBS 0.008671f
C428 B.n388 VSUBS 0.008671f
C429 B.n389 VSUBS 0.008671f
C430 B.n390 VSUBS 0.008671f
C431 B.n391 VSUBS 0.008671f
C432 B.n392 VSUBS 0.008671f
C433 B.n393 VSUBS 0.008671f
C434 B.n394 VSUBS 0.008671f
C435 B.n395 VSUBS 0.008671f
C436 B.n396 VSUBS 0.008671f
C437 B.n397 VSUBS 0.008671f
C438 B.n398 VSUBS 0.008671f
C439 B.n399 VSUBS 0.008671f
C440 B.n400 VSUBS 0.008671f
C441 B.n401 VSUBS 0.008671f
C442 B.n402 VSUBS 0.008671f
C443 B.n403 VSUBS 0.008671f
C444 B.n404 VSUBS 0.008671f
C445 B.n405 VSUBS 0.008671f
C446 B.n406 VSUBS 0.008671f
C447 B.n407 VSUBS 0.008671f
C448 B.n408 VSUBS 0.008671f
C449 B.n409 VSUBS 0.008671f
C450 B.n410 VSUBS 0.008671f
C451 B.n411 VSUBS 0.008671f
C452 B.n412 VSUBS 0.008671f
C453 B.n413 VSUBS 0.008671f
C454 B.n414 VSUBS 0.008671f
C455 B.n415 VSUBS 0.008671f
C456 B.n416 VSUBS 0.008671f
C457 B.n417 VSUBS 0.008671f
C458 B.n418 VSUBS 0.008671f
C459 B.n419 VSUBS 0.008671f
C460 B.n420 VSUBS 0.008671f
C461 B.n421 VSUBS 0.008671f
C462 B.n422 VSUBS 0.008671f
C463 B.n423 VSUBS 0.008671f
C464 B.n424 VSUBS 0.008671f
C465 B.n425 VSUBS 0.008671f
C466 B.n426 VSUBS 0.008671f
C467 B.n427 VSUBS 0.008671f
C468 B.n428 VSUBS 0.008671f
C469 B.n429 VSUBS 0.008671f
C470 B.n430 VSUBS 0.008671f
C471 B.n431 VSUBS 0.008671f
C472 B.n432 VSUBS 0.008671f
C473 B.n433 VSUBS 0.008671f
C474 B.n434 VSUBS 0.008671f
C475 B.n435 VSUBS 0.008671f
C476 B.n436 VSUBS 0.008671f
C477 B.n437 VSUBS 0.008671f
C478 B.n438 VSUBS 0.008671f
C479 B.n439 VSUBS 0.008671f
C480 B.n440 VSUBS 0.008671f
C481 B.n441 VSUBS 0.008671f
C482 B.n442 VSUBS 0.008671f
C483 B.n443 VSUBS 0.008671f
C484 B.n444 VSUBS 0.008671f
C485 B.n445 VSUBS 0.008671f
C486 B.n446 VSUBS 0.008671f
C487 B.n447 VSUBS 0.008671f
C488 B.n448 VSUBS 0.008671f
C489 B.n449 VSUBS 0.008671f
C490 B.n450 VSUBS 0.008671f
C491 B.n451 VSUBS 0.008671f
C492 B.n452 VSUBS 0.008671f
C493 B.n453 VSUBS 0.008671f
C494 B.n454 VSUBS 0.008671f
C495 B.n455 VSUBS 0.008671f
C496 B.n456 VSUBS 0.008671f
C497 B.n457 VSUBS 0.008671f
C498 B.n458 VSUBS 0.008671f
C499 B.n459 VSUBS 0.008671f
C500 B.n460 VSUBS 0.008671f
C501 B.n461 VSUBS 0.008671f
C502 B.n462 VSUBS 0.008671f
C503 B.n463 VSUBS 0.008671f
C504 B.n464 VSUBS 0.008671f
C505 B.n465 VSUBS 0.008671f
C506 B.n466 VSUBS 0.008671f
C507 B.n467 VSUBS 0.008671f
C508 B.n468 VSUBS 0.008671f
C509 B.n469 VSUBS 0.008671f
C510 B.n470 VSUBS 0.008671f
C511 B.n471 VSUBS 0.008671f
C512 B.n472 VSUBS 0.008671f
C513 B.n473 VSUBS 0.008671f
C514 B.n474 VSUBS 0.008671f
C515 B.n475 VSUBS 0.008671f
C516 B.n476 VSUBS 0.008671f
C517 B.n477 VSUBS 0.008671f
C518 B.n478 VSUBS 0.008671f
C519 B.n479 VSUBS 0.008671f
C520 B.n480 VSUBS 0.008671f
C521 B.n481 VSUBS 0.008671f
C522 B.n482 VSUBS 0.008671f
C523 B.n483 VSUBS 0.008671f
C524 B.n484 VSUBS 0.008671f
C525 B.n485 VSUBS 0.008671f
C526 B.n486 VSUBS 0.008671f
C527 B.n487 VSUBS 0.008671f
C528 B.n488 VSUBS 0.008671f
C529 B.n489 VSUBS 0.008671f
C530 B.n490 VSUBS 0.008671f
C531 B.n491 VSUBS 0.008671f
C532 B.n492 VSUBS 0.008671f
C533 B.n493 VSUBS 0.008671f
C534 B.n494 VSUBS 0.008671f
C535 B.n495 VSUBS 0.008671f
C536 B.n496 VSUBS 0.008671f
C537 B.n497 VSUBS 0.021081f
C538 B.n498 VSUBS 0.022017f
C539 B.n499 VSUBS 0.021081f
C540 B.n500 VSUBS 0.008671f
C541 B.n501 VSUBS 0.008671f
C542 B.n502 VSUBS 0.008671f
C543 B.n503 VSUBS 0.008671f
C544 B.n504 VSUBS 0.008671f
C545 B.n505 VSUBS 0.008671f
C546 B.n506 VSUBS 0.008671f
C547 B.n507 VSUBS 0.008671f
C548 B.n508 VSUBS 0.008671f
C549 B.n509 VSUBS 0.008671f
C550 B.n510 VSUBS 0.008671f
C551 B.n511 VSUBS 0.008671f
C552 B.n512 VSUBS 0.008671f
C553 B.n513 VSUBS 0.008671f
C554 B.n514 VSUBS 0.008671f
C555 B.n515 VSUBS 0.008671f
C556 B.n516 VSUBS 0.008671f
C557 B.n517 VSUBS 0.008671f
C558 B.n518 VSUBS 0.008671f
C559 B.n519 VSUBS 0.008671f
C560 B.n520 VSUBS 0.008671f
C561 B.n521 VSUBS 0.008671f
C562 B.n522 VSUBS 0.008671f
C563 B.n523 VSUBS 0.008671f
C564 B.n524 VSUBS 0.008161f
C565 B.n525 VSUBS 0.008671f
C566 B.n526 VSUBS 0.008671f
C567 B.n527 VSUBS 0.008671f
C568 B.n528 VSUBS 0.008671f
C569 B.n529 VSUBS 0.008671f
C570 B.n530 VSUBS 0.008671f
C571 B.n531 VSUBS 0.008671f
C572 B.n532 VSUBS 0.008671f
C573 B.n533 VSUBS 0.008671f
C574 B.n534 VSUBS 0.008671f
C575 B.n535 VSUBS 0.008671f
C576 B.n536 VSUBS 0.008671f
C577 B.n537 VSUBS 0.008671f
C578 B.n538 VSUBS 0.008671f
C579 B.n539 VSUBS 0.008671f
C580 B.n540 VSUBS 0.004845f
C581 B.n541 VSUBS 0.020089f
C582 B.n542 VSUBS 0.008161f
C583 B.n543 VSUBS 0.008671f
C584 B.n544 VSUBS 0.008671f
C585 B.n545 VSUBS 0.008671f
C586 B.n546 VSUBS 0.008671f
C587 B.n547 VSUBS 0.008671f
C588 B.n548 VSUBS 0.008671f
C589 B.n549 VSUBS 0.008671f
C590 B.n550 VSUBS 0.008671f
C591 B.n551 VSUBS 0.008671f
C592 B.n552 VSUBS 0.008671f
C593 B.n553 VSUBS 0.008671f
C594 B.n554 VSUBS 0.008671f
C595 B.n555 VSUBS 0.008671f
C596 B.n556 VSUBS 0.008671f
C597 B.n557 VSUBS 0.008671f
C598 B.n558 VSUBS 0.008671f
C599 B.n559 VSUBS 0.008671f
C600 B.n560 VSUBS 0.008671f
C601 B.n561 VSUBS 0.008671f
C602 B.n562 VSUBS 0.008671f
C603 B.n563 VSUBS 0.008671f
C604 B.n564 VSUBS 0.008671f
C605 B.n565 VSUBS 0.008671f
C606 B.n566 VSUBS 0.008671f
C607 B.n567 VSUBS 0.022017f
C608 B.n568 VSUBS 0.022017f
C609 B.n569 VSUBS 0.021081f
C610 B.n570 VSUBS 0.008671f
C611 B.n571 VSUBS 0.008671f
C612 B.n572 VSUBS 0.008671f
C613 B.n573 VSUBS 0.008671f
C614 B.n574 VSUBS 0.008671f
C615 B.n575 VSUBS 0.008671f
C616 B.n576 VSUBS 0.008671f
C617 B.n577 VSUBS 0.008671f
C618 B.n578 VSUBS 0.008671f
C619 B.n579 VSUBS 0.008671f
C620 B.n580 VSUBS 0.008671f
C621 B.n581 VSUBS 0.008671f
C622 B.n582 VSUBS 0.008671f
C623 B.n583 VSUBS 0.008671f
C624 B.n584 VSUBS 0.008671f
C625 B.n585 VSUBS 0.008671f
C626 B.n586 VSUBS 0.008671f
C627 B.n587 VSUBS 0.008671f
C628 B.n588 VSUBS 0.008671f
C629 B.n589 VSUBS 0.008671f
C630 B.n590 VSUBS 0.008671f
C631 B.n591 VSUBS 0.008671f
C632 B.n592 VSUBS 0.008671f
C633 B.n593 VSUBS 0.008671f
C634 B.n594 VSUBS 0.008671f
C635 B.n595 VSUBS 0.008671f
C636 B.n596 VSUBS 0.008671f
C637 B.n597 VSUBS 0.008671f
C638 B.n598 VSUBS 0.008671f
C639 B.n599 VSUBS 0.008671f
C640 B.n600 VSUBS 0.008671f
C641 B.n601 VSUBS 0.008671f
C642 B.n602 VSUBS 0.008671f
C643 B.n603 VSUBS 0.008671f
C644 B.n604 VSUBS 0.008671f
C645 B.n605 VSUBS 0.008671f
C646 B.n606 VSUBS 0.008671f
C647 B.n607 VSUBS 0.008671f
C648 B.n608 VSUBS 0.008671f
C649 B.n609 VSUBS 0.008671f
C650 B.n610 VSUBS 0.008671f
C651 B.n611 VSUBS 0.008671f
C652 B.n612 VSUBS 0.008671f
C653 B.n613 VSUBS 0.008671f
C654 B.n614 VSUBS 0.008671f
C655 B.n615 VSUBS 0.008671f
C656 B.n616 VSUBS 0.008671f
C657 B.n617 VSUBS 0.008671f
C658 B.n618 VSUBS 0.008671f
C659 B.n619 VSUBS 0.008671f
C660 B.n620 VSUBS 0.008671f
C661 B.n621 VSUBS 0.008671f
C662 B.n622 VSUBS 0.008671f
C663 B.n623 VSUBS 0.008671f
C664 B.n624 VSUBS 0.008671f
C665 B.n625 VSUBS 0.008671f
C666 B.n626 VSUBS 0.008671f
C667 B.n627 VSUBS 0.008671f
C668 B.n628 VSUBS 0.008671f
C669 B.n629 VSUBS 0.008671f
C670 B.n630 VSUBS 0.008671f
C671 B.n631 VSUBS 0.008671f
C672 B.n632 VSUBS 0.008671f
C673 B.n633 VSUBS 0.008671f
C674 B.n634 VSUBS 0.008671f
C675 B.n635 VSUBS 0.008671f
C676 B.n636 VSUBS 0.008671f
C677 B.n637 VSUBS 0.008671f
C678 B.n638 VSUBS 0.008671f
C679 B.n639 VSUBS 0.008671f
C680 B.n640 VSUBS 0.008671f
C681 B.n641 VSUBS 0.008671f
C682 B.n642 VSUBS 0.008671f
C683 B.n643 VSUBS 0.008671f
C684 B.n644 VSUBS 0.008671f
C685 B.n645 VSUBS 0.008671f
C686 B.n646 VSUBS 0.008671f
C687 B.n647 VSUBS 0.008671f
C688 B.n648 VSUBS 0.008671f
C689 B.n649 VSUBS 0.008671f
C690 B.n650 VSUBS 0.008671f
C691 B.n651 VSUBS 0.008671f
C692 B.n652 VSUBS 0.008671f
C693 B.n653 VSUBS 0.008671f
C694 B.n654 VSUBS 0.008671f
C695 B.n655 VSUBS 0.019634f
C696 VDD2.t9 VSUBS 0.857492f
C697 VDD2.t4 VSUBS 0.104157f
C698 VDD2.t8 VSUBS 0.104157f
C699 VDD2.n0 VSUBS 0.6126f
C700 VDD2.n1 VSUBS 1.52865f
C701 VDD2.t3 VSUBS 0.104157f
C702 VDD2.t7 VSUBS 0.104157f
C703 VDD2.n2 VSUBS 0.627177f
C704 VDD2.n3 VSUBS 3.22768f
C705 VDD2.t0 VSUBS 0.841514f
C706 VDD2.n4 VSUBS 3.31708f
C707 VDD2.t1 VSUBS 0.104157f
C708 VDD2.t6 VSUBS 0.104157f
C709 VDD2.n5 VSUBS 0.612602f
C710 VDD2.n6 VSUBS 0.777583f
C711 VDD2.t2 VSUBS 0.104157f
C712 VDD2.t5 VSUBS 0.104157f
C713 VDD2.n7 VSUBS 0.627141f
C714 VN.n0 VSUBS 0.054705f
C715 VN.t2 VSUBS 1.07026f
C716 VN.n1 VSUBS 0.037085f
C717 VN.n2 VSUBS 0.041494f
C718 VN.t6 VSUBS 1.07026f
C719 VN.n3 VSUBS 0.077334f
C720 VN.n4 VSUBS 0.041494f
C721 VN.n5 VSUBS 0.058244f
C722 VN.n6 VSUBS 0.041494f
C723 VN.n7 VSUBS 0.07273f
C724 VN.n8 VSUBS 0.363508f
C725 VN.t5 VSUBS 1.07026f
C726 VN.t0 VSUBS 1.36841f
C727 VN.n9 VSUBS 0.521782f
C728 VN.n10 VSUBS 0.527138f
C729 VN.n11 VSUBS 0.041444f
C730 VN.n12 VSUBS 0.077334f
C731 VN.n13 VSUBS 0.041494f
C732 VN.n14 VSUBS 0.041494f
C733 VN.n15 VSUBS 0.041494f
C734 VN.n16 VSUBS 0.045316f
C735 VN.n17 VSUBS 0.080434f
C736 VN.t1 VSUBS 1.07026f
C737 VN.n18 VSUBS 0.426589f
C738 VN.n19 VSUBS 0.058244f
C739 VN.n20 VSUBS 0.041494f
C740 VN.n21 VSUBS 0.041494f
C741 VN.n22 VSUBS 0.041494f
C742 VN.n23 VSUBS 0.080434f
C743 VN.n24 VSUBS 0.045316f
C744 VN.n25 VSUBS 0.07273f
C745 VN.n26 VSUBS 0.041494f
C746 VN.n27 VSUBS 0.041494f
C747 VN.n28 VSUBS 0.041494f
C748 VN.n29 VSUBS 0.041444f
C749 VN.n30 VSUBS 0.426589f
C750 VN.n31 VSUBS 0.075043f
C751 VN.n32 VSUBS 0.077707f
C752 VN.n33 VSUBS 0.041494f
C753 VN.n34 VSUBS 0.041494f
C754 VN.n35 VSUBS 0.041494f
C755 VN.n36 VSUBS 0.083688f
C756 VN.n37 VSUBS 0.062825f
C757 VN.n38 VSUBS 0.569765f
C758 VN.n39 VSUBS 0.059781f
C759 VN.n40 VSUBS 0.054705f
C760 VN.t9 VSUBS 1.07026f
C761 VN.n41 VSUBS 0.037085f
C762 VN.n42 VSUBS 0.041494f
C763 VN.t8 VSUBS 1.07026f
C764 VN.n43 VSUBS 0.077334f
C765 VN.n44 VSUBS 0.041494f
C766 VN.n45 VSUBS 0.058244f
C767 VN.n46 VSUBS 0.041494f
C768 VN.t3 VSUBS 1.07026f
C769 VN.n47 VSUBS 0.426589f
C770 VN.n48 VSUBS 0.07273f
C771 VN.n49 VSUBS 0.363508f
C772 VN.t7 VSUBS 1.07026f
C773 VN.t4 VSUBS 1.36841f
C774 VN.n50 VSUBS 0.521782f
C775 VN.n51 VSUBS 0.527138f
C776 VN.n52 VSUBS 0.041444f
C777 VN.n53 VSUBS 0.077334f
C778 VN.n54 VSUBS 0.041494f
C779 VN.n55 VSUBS 0.041494f
C780 VN.n56 VSUBS 0.041494f
C781 VN.n57 VSUBS 0.045316f
C782 VN.n58 VSUBS 0.080434f
C783 VN.n59 VSUBS 0.058244f
C784 VN.n60 VSUBS 0.041494f
C785 VN.n61 VSUBS 0.041494f
C786 VN.n62 VSUBS 0.041494f
C787 VN.n63 VSUBS 0.080434f
C788 VN.n64 VSUBS 0.045316f
C789 VN.n65 VSUBS 0.07273f
C790 VN.n66 VSUBS 0.041494f
C791 VN.n67 VSUBS 0.041494f
C792 VN.n68 VSUBS 0.041494f
C793 VN.n69 VSUBS 0.041444f
C794 VN.n70 VSUBS 0.426589f
C795 VN.n71 VSUBS 0.075043f
C796 VN.n72 VSUBS 0.077707f
C797 VN.n73 VSUBS 0.041494f
C798 VN.n74 VSUBS 0.041494f
C799 VN.n75 VSUBS 0.041494f
C800 VN.n76 VSUBS 0.083688f
C801 VN.n77 VSUBS 0.062825f
C802 VN.n78 VSUBS 0.569765f
C803 VN.n79 VSUBS 2.07804f
C804 VDD1.t7 VSUBS 0.862087f
C805 VDD1.t6 VSUBS 0.104715f
C806 VDD1.t2 VSUBS 0.104715f
C807 VDD1.n0 VSUBS 0.615883f
C808 VDD1.n1 VSUBS 1.5473f
C809 VDD1.t8 VSUBS 0.862084f
C810 VDD1.t3 VSUBS 0.104715f
C811 VDD1.t0 VSUBS 0.104715f
C812 VDD1.n2 VSUBS 0.615881f
C813 VDD1.n3 VSUBS 1.53684f
C814 VDD1.t4 VSUBS 0.104715f
C815 VDD1.t9 VSUBS 0.104715f
C816 VDD1.n4 VSUBS 0.630535f
C817 VDD1.n5 VSUBS 3.39322f
C818 VDD1.t1 VSUBS 0.104715f
C819 VDD1.t5 VSUBS 0.104715f
C820 VDD1.n6 VSUBS 0.61588f
C821 VDD1.n7 VSUBS 3.43238f
C822 VTAIL.t8 VSUBS 0.108668f
C823 VTAIL.t3 VSUBS 0.108668f
C824 VTAIL.n0 VSUBS 0.550871f
C825 VTAIL.n1 VSUBS 0.904726f
C826 VTAIL.t15 VSUBS 0.787048f
C827 VTAIL.n2 VSUBS 1.02352f
C828 VTAIL.t18 VSUBS 0.108668f
C829 VTAIL.t17 VSUBS 0.108668f
C830 VTAIL.n3 VSUBS 0.550871f
C831 VTAIL.n4 VSUBS 1.04225f
C832 VTAIL.t16 VSUBS 0.108668f
C833 VTAIL.t14 VSUBS 0.108668f
C834 VTAIL.n5 VSUBS 0.550871f
C835 VTAIL.n6 VSUBS 2.14059f
C836 VTAIL.t2 VSUBS 0.108668f
C837 VTAIL.t6 VSUBS 0.108668f
C838 VTAIL.n7 VSUBS 0.550874f
C839 VTAIL.n8 VSUBS 2.14058f
C840 VTAIL.t7 VSUBS 0.108668f
C841 VTAIL.t5 VSUBS 0.108668f
C842 VTAIL.n9 VSUBS 0.550874f
C843 VTAIL.n10 VSUBS 1.04225f
C844 VTAIL.t4 VSUBS 0.787052f
C845 VTAIL.n11 VSUBS 1.02352f
C846 VTAIL.t12 VSUBS 0.108668f
C847 VTAIL.t11 VSUBS 0.108668f
C848 VTAIL.n12 VSUBS 0.550874f
C849 VTAIL.n13 VSUBS 0.963328f
C850 VTAIL.t13 VSUBS 0.108668f
C851 VTAIL.t19 VSUBS 0.108668f
C852 VTAIL.n14 VSUBS 0.550874f
C853 VTAIL.n15 VSUBS 1.04225f
C854 VTAIL.t10 VSUBS 0.787048f
C855 VTAIL.n16 VSUBS 1.94114f
C856 VTAIL.t0 VSUBS 0.787048f
C857 VTAIL.n17 VSUBS 1.94114f
C858 VTAIL.t1 VSUBS 0.108668f
C859 VTAIL.t9 VSUBS 0.108668f
C860 VTAIL.n18 VSUBS 0.550871f
C861 VTAIL.n19 VSUBS 0.841218f
C862 VP.n0 VSUBS 0.061717f
C863 VP.t0 VSUBS 1.20744f
C864 VP.n1 VSUBS 0.041838f
C865 VP.n2 VSUBS 0.046812f
C866 VP.t5 VSUBS 1.20744f
C867 VP.n3 VSUBS 0.087245f
C868 VP.n4 VSUBS 0.046812f
C869 VP.n5 VSUBS 0.065709f
C870 VP.n6 VSUBS 0.046812f
C871 VP.n7 VSUBS 0.082052f
C872 VP.n8 VSUBS 0.046812f
C873 VP.t6 VSUBS 1.20744f
C874 VP.n9 VSUBS 0.087666f
C875 VP.n10 VSUBS 0.046812f
C876 VP.t1 VSUBS 1.20744f
C877 VP.n11 VSUBS 0.642792f
C878 VP.n12 VSUBS 0.061717f
C879 VP.t4 VSUBS 1.20744f
C880 VP.n13 VSUBS 0.041838f
C881 VP.n14 VSUBS 0.046812f
C882 VP.t8 VSUBS 1.20744f
C883 VP.n15 VSUBS 0.087245f
C884 VP.n16 VSUBS 0.046812f
C885 VP.n17 VSUBS 0.065709f
C886 VP.n18 VSUBS 0.046812f
C887 VP.n19 VSUBS 0.082052f
C888 VP.n20 VSUBS 0.410099f
C889 VP.t3 VSUBS 1.20744f
C890 VP.t2 VSUBS 1.5438f
C891 VP.n21 VSUBS 0.588659f
C892 VP.n22 VSUBS 0.594702f
C893 VP.n23 VSUBS 0.046756f
C894 VP.n24 VSUBS 0.087245f
C895 VP.n25 VSUBS 0.046812f
C896 VP.n26 VSUBS 0.046812f
C897 VP.n27 VSUBS 0.046812f
C898 VP.n28 VSUBS 0.051124f
C899 VP.n29 VSUBS 0.090743f
C900 VP.t7 VSUBS 1.20744f
C901 VP.n30 VSUBS 0.481265f
C902 VP.n31 VSUBS 0.065709f
C903 VP.n32 VSUBS 0.046812f
C904 VP.n33 VSUBS 0.046812f
C905 VP.n34 VSUBS 0.046812f
C906 VP.n35 VSUBS 0.090743f
C907 VP.n36 VSUBS 0.051124f
C908 VP.n37 VSUBS 0.082052f
C909 VP.n38 VSUBS 0.046812f
C910 VP.n39 VSUBS 0.046812f
C911 VP.n40 VSUBS 0.046812f
C912 VP.n41 VSUBS 0.046756f
C913 VP.n42 VSUBS 0.481265f
C914 VP.n43 VSUBS 0.084661f
C915 VP.n44 VSUBS 0.087666f
C916 VP.n45 VSUBS 0.046812f
C917 VP.n46 VSUBS 0.046812f
C918 VP.n47 VSUBS 0.046812f
C919 VP.n48 VSUBS 0.094415f
C920 VP.n49 VSUBS 0.070877f
C921 VP.n50 VSUBS 0.642792f
C922 VP.n51 VSUBS 2.31892f
C923 VP.n52 VSUBS 2.35521f
C924 VP.n53 VSUBS 0.061717f
C925 VP.n54 VSUBS 0.070877f
C926 VP.n55 VSUBS 0.094415f
C927 VP.n56 VSUBS 0.041838f
C928 VP.n57 VSUBS 0.046812f
C929 VP.n58 VSUBS 0.046812f
C930 VP.n59 VSUBS 0.046812f
C931 VP.n60 VSUBS 0.084661f
C932 VP.n61 VSUBS 0.481265f
C933 VP.n62 VSUBS 0.046756f
C934 VP.n63 VSUBS 0.087245f
C935 VP.n64 VSUBS 0.046812f
C936 VP.n65 VSUBS 0.046812f
C937 VP.n66 VSUBS 0.046812f
C938 VP.n67 VSUBS 0.051124f
C939 VP.n68 VSUBS 0.090743f
C940 VP.t9 VSUBS 1.20744f
C941 VP.n69 VSUBS 0.481265f
C942 VP.n70 VSUBS 0.065709f
C943 VP.n71 VSUBS 0.046812f
C944 VP.n72 VSUBS 0.046812f
C945 VP.n73 VSUBS 0.046812f
C946 VP.n74 VSUBS 0.090743f
C947 VP.n75 VSUBS 0.051124f
C948 VP.n76 VSUBS 0.082052f
C949 VP.n77 VSUBS 0.046812f
C950 VP.n78 VSUBS 0.046812f
C951 VP.n79 VSUBS 0.046812f
C952 VP.n80 VSUBS 0.046756f
C953 VP.n81 VSUBS 0.481265f
C954 VP.n82 VSUBS 0.084661f
C955 VP.n83 VSUBS 0.087666f
C956 VP.n84 VSUBS 0.046812f
C957 VP.n85 VSUBS 0.046812f
C958 VP.n86 VSUBS 0.046812f
C959 VP.n87 VSUBS 0.094415f
C960 VP.n88 VSUBS 0.070877f
C961 VP.n89 VSUBS 0.642792f
C962 VP.n90 VSUBS 0.067443f
.ends

