* NGSPICE file created from diff_pair_sample_0779.ext - technology: sky130A

.subckt diff_pair_sample_0779 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=0.48
X1 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=0.48
X2 VDD1.t2 VP.t1 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=0.48
X3 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=0.48
X4 VTAIL.t7 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=0.48
X5 VTAIL.t0 VN.t0 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=0.48
X6 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=0.48
X7 VTAIL.t6 VP.t3 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=0.48
X8 VDD2.t2 VN.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=0.48
X9 VDD2.t1 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.51975 pd=3.48 as=1.2285 ps=7.08 w=3.15 l=0.48
X10 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0 ps=0 w=3.15 l=0.48
X11 VTAIL.t3 VN.t3 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2285 pd=7.08 as=0.51975 ps=3.48 w=3.15 l=0.48
R0 VP.n0 VP.t3 261.481
R1 VP.n0 VP.t0 261.455
R2 VP.n2 VP.t2 240.499
R3 VP.n3 VP.t1 240.499
R4 VP.n4 VP.n3 161.3
R5 VP.n2 VP.n1 161.3
R6 VP.n1 VP.n0 103.275
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n122 VTAIL.n112 289.615
R11 VTAIL.n10 VTAIL.n0 289.615
R12 VTAIL.n26 VTAIL.n16 289.615
R13 VTAIL.n42 VTAIL.n32 289.615
R14 VTAIL.n106 VTAIL.n96 289.615
R15 VTAIL.n90 VTAIL.n80 289.615
R16 VTAIL.n74 VTAIL.n64 289.615
R17 VTAIL.n58 VTAIL.n48 289.615
R18 VTAIL.n116 VTAIL.n115 185
R19 VTAIL.n121 VTAIL.n120 185
R20 VTAIL.n123 VTAIL.n122 185
R21 VTAIL.n4 VTAIL.n3 185
R22 VTAIL.n9 VTAIL.n8 185
R23 VTAIL.n11 VTAIL.n10 185
R24 VTAIL.n20 VTAIL.n19 185
R25 VTAIL.n25 VTAIL.n24 185
R26 VTAIL.n27 VTAIL.n26 185
R27 VTAIL.n36 VTAIL.n35 185
R28 VTAIL.n41 VTAIL.n40 185
R29 VTAIL.n43 VTAIL.n42 185
R30 VTAIL.n107 VTAIL.n106 185
R31 VTAIL.n105 VTAIL.n104 185
R32 VTAIL.n100 VTAIL.n99 185
R33 VTAIL.n91 VTAIL.n90 185
R34 VTAIL.n89 VTAIL.n88 185
R35 VTAIL.n84 VTAIL.n83 185
R36 VTAIL.n75 VTAIL.n74 185
R37 VTAIL.n73 VTAIL.n72 185
R38 VTAIL.n68 VTAIL.n67 185
R39 VTAIL.n59 VTAIL.n58 185
R40 VTAIL.n57 VTAIL.n56 185
R41 VTAIL.n52 VTAIL.n51 185
R42 VTAIL.n117 VTAIL.t1 148.606
R43 VTAIL.n5 VTAIL.t3 148.606
R44 VTAIL.n21 VTAIL.t4 148.606
R45 VTAIL.n37 VTAIL.t7 148.606
R46 VTAIL.n101 VTAIL.t5 148.606
R47 VTAIL.n85 VTAIL.t6 148.606
R48 VTAIL.n69 VTAIL.t2 148.606
R49 VTAIL.n53 VTAIL.t0 148.606
R50 VTAIL.n121 VTAIL.n115 104.615
R51 VTAIL.n122 VTAIL.n121 104.615
R52 VTAIL.n9 VTAIL.n3 104.615
R53 VTAIL.n10 VTAIL.n9 104.615
R54 VTAIL.n25 VTAIL.n19 104.615
R55 VTAIL.n26 VTAIL.n25 104.615
R56 VTAIL.n41 VTAIL.n35 104.615
R57 VTAIL.n42 VTAIL.n41 104.615
R58 VTAIL.n106 VTAIL.n105 104.615
R59 VTAIL.n105 VTAIL.n99 104.615
R60 VTAIL.n90 VTAIL.n89 104.615
R61 VTAIL.n89 VTAIL.n83 104.615
R62 VTAIL.n74 VTAIL.n73 104.615
R63 VTAIL.n73 VTAIL.n67 104.615
R64 VTAIL.n58 VTAIL.n57 104.615
R65 VTAIL.n57 VTAIL.n51 104.615
R66 VTAIL.t1 VTAIL.n115 52.3082
R67 VTAIL.t3 VTAIL.n3 52.3082
R68 VTAIL.t4 VTAIL.n19 52.3082
R69 VTAIL.t7 VTAIL.n35 52.3082
R70 VTAIL.t5 VTAIL.n99 52.3082
R71 VTAIL.t6 VTAIL.n83 52.3082
R72 VTAIL.t2 VTAIL.n67 52.3082
R73 VTAIL.t0 VTAIL.n51 52.3082
R74 VTAIL.n127 VTAIL.n126 32.7672
R75 VTAIL.n15 VTAIL.n14 32.7672
R76 VTAIL.n31 VTAIL.n30 32.7672
R77 VTAIL.n47 VTAIL.n46 32.7672
R78 VTAIL.n111 VTAIL.n110 32.7672
R79 VTAIL.n95 VTAIL.n94 32.7672
R80 VTAIL.n79 VTAIL.n78 32.7672
R81 VTAIL.n63 VTAIL.n62 32.7672
R82 VTAIL.n127 VTAIL.n111 15.7807
R83 VTAIL.n63 VTAIL.n47 15.7807
R84 VTAIL.n117 VTAIL.n116 15.5966
R85 VTAIL.n5 VTAIL.n4 15.5966
R86 VTAIL.n21 VTAIL.n20 15.5966
R87 VTAIL.n37 VTAIL.n36 15.5966
R88 VTAIL.n101 VTAIL.n100 15.5966
R89 VTAIL.n85 VTAIL.n84 15.5966
R90 VTAIL.n69 VTAIL.n68 15.5966
R91 VTAIL.n53 VTAIL.n52 15.5966
R92 VTAIL.n120 VTAIL.n119 12.8005
R93 VTAIL.n8 VTAIL.n7 12.8005
R94 VTAIL.n24 VTAIL.n23 12.8005
R95 VTAIL.n40 VTAIL.n39 12.8005
R96 VTAIL.n104 VTAIL.n103 12.8005
R97 VTAIL.n88 VTAIL.n87 12.8005
R98 VTAIL.n72 VTAIL.n71 12.8005
R99 VTAIL.n56 VTAIL.n55 12.8005
R100 VTAIL.n123 VTAIL.n114 12.0247
R101 VTAIL.n11 VTAIL.n2 12.0247
R102 VTAIL.n27 VTAIL.n18 12.0247
R103 VTAIL.n43 VTAIL.n34 12.0247
R104 VTAIL.n107 VTAIL.n98 12.0247
R105 VTAIL.n91 VTAIL.n82 12.0247
R106 VTAIL.n75 VTAIL.n66 12.0247
R107 VTAIL.n59 VTAIL.n50 12.0247
R108 VTAIL.n124 VTAIL.n112 11.249
R109 VTAIL.n12 VTAIL.n0 11.249
R110 VTAIL.n28 VTAIL.n16 11.249
R111 VTAIL.n44 VTAIL.n32 11.249
R112 VTAIL.n108 VTAIL.n96 11.249
R113 VTAIL.n92 VTAIL.n80 11.249
R114 VTAIL.n76 VTAIL.n64 11.249
R115 VTAIL.n60 VTAIL.n48 11.249
R116 VTAIL.n126 VTAIL.n125 9.45567
R117 VTAIL.n14 VTAIL.n13 9.45567
R118 VTAIL.n30 VTAIL.n29 9.45567
R119 VTAIL.n46 VTAIL.n45 9.45567
R120 VTAIL.n110 VTAIL.n109 9.45567
R121 VTAIL.n94 VTAIL.n93 9.45567
R122 VTAIL.n78 VTAIL.n77 9.45567
R123 VTAIL.n62 VTAIL.n61 9.45567
R124 VTAIL.n125 VTAIL.n124 9.3005
R125 VTAIL.n114 VTAIL.n113 9.3005
R126 VTAIL.n119 VTAIL.n118 9.3005
R127 VTAIL.n13 VTAIL.n12 9.3005
R128 VTAIL.n2 VTAIL.n1 9.3005
R129 VTAIL.n7 VTAIL.n6 9.3005
R130 VTAIL.n29 VTAIL.n28 9.3005
R131 VTAIL.n18 VTAIL.n17 9.3005
R132 VTAIL.n23 VTAIL.n22 9.3005
R133 VTAIL.n45 VTAIL.n44 9.3005
R134 VTAIL.n34 VTAIL.n33 9.3005
R135 VTAIL.n39 VTAIL.n38 9.3005
R136 VTAIL.n109 VTAIL.n108 9.3005
R137 VTAIL.n98 VTAIL.n97 9.3005
R138 VTAIL.n103 VTAIL.n102 9.3005
R139 VTAIL.n93 VTAIL.n92 9.3005
R140 VTAIL.n82 VTAIL.n81 9.3005
R141 VTAIL.n87 VTAIL.n86 9.3005
R142 VTAIL.n77 VTAIL.n76 9.3005
R143 VTAIL.n66 VTAIL.n65 9.3005
R144 VTAIL.n71 VTAIL.n70 9.3005
R145 VTAIL.n61 VTAIL.n60 9.3005
R146 VTAIL.n50 VTAIL.n49 9.3005
R147 VTAIL.n55 VTAIL.n54 9.3005
R148 VTAIL.n118 VTAIL.n117 4.46457
R149 VTAIL.n6 VTAIL.n5 4.46457
R150 VTAIL.n22 VTAIL.n21 4.46457
R151 VTAIL.n38 VTAIL.n37 4.46457
R152 VTAIL.n102 VTAIL.n101 4.46457
R153 VTAIL.n86 VTAIL.n85 4.46457
R154 VTAIL.n70 VTAIL.n69 4.46457
R155 VTAIL.n54 VTAIL.n53 4.46457
R156 VTAIL.n126 VTAIL.n112 2.71565
R157 VTAIL.n14 VTAIL.n0 2.71565
R158 VTAIL.n30 VTAIL.n16 2.71565
R159 VTAIL.n46 VTAIL.n32 2.71565
R160 VTAIL.n110 VTAIL.n96 2.71565
R161 VTAIL.n94 VTAIL.n80 2.71565
R162 VTAIL.n78 VTAIL.n64 2.71565
R163 VTAIL.n62 VTAIL.n48 2.71565
R164 VTAIL.n124 VTAIL.n123 1.93989
R165 VTAIL.n12 VTAIL.n11 1.93989
R166 VTAIL.n28 VTAIL.n27 1.93989
R167 VTAIL.n44 VTAIL.n43 1.93989
R168 VTAIL.n108 VTAIL.n107 1.93989
R169 VTAIL.n92 VTAIL.n91 1.93989
R170 VTAIL.n76 VTAIL.n75 1.93989
R171 VTAIL.n60 VTAIL.n59 1.93989
R172 VTAIL.n120 VTAIL.n114 1.16414
R173 VTAIL.n8 VTAIL.n2 1.16414
R174 VTAIL.n24 VTAIL.n18 1.16414
R175 VTAIL.n40 VTAIL.n34 1.16414
R176 VTAIL.n104 VTAIL.n98 1.16414
R177 VTAIL.n88 VTAIL.n82 1.16414
R178 VTAIL.n72 VTAIL.n66 1.16414
R179 VTAIL.n56 VTAIL.n50 1.16414
R180 VTAIL.n79 VTAIL.n63 0.698776
R181 VTAIL.n111 VTAIL.n95 0.698776
R182 VTAIL.n47 VTAIL.n31 0.698776
R183 VTAIL.n95 VTAIL.n79 0.470328
R184 VTAIL.n31 VTAIL.n15 0.470328
R185 VTAIL VTAIL.n15 0.407828
R186 VTAIL.n119 VTAIL.n116 0.388379
R187 VTAIL.n7 VTAIL.n4 0.388379
R188 VTAIL.n23 VTAIL.n20 0.388379
R189 VTAIL.n39 VTAIL.n36 0.388379
R190 VTAIL.n103 VTAIL.n100 0.388379
R191 VTAIL.n87 VTAIL.n84 0.388379
R192 VTAIL.n71 VTAIL.n68 0.388379
R193 VTAIL.n55 VTAIL.n52 0.388379
R194 VTAIL VTAIL.n127 0.291448
R195 VTAIL.n118 VTAIL.n113 0.155672
R196 VTAIL.n125 VTAIL.n113 0.155672
R197 VTAIL.n6 VTAIL.n1 0.155672
R198 VTAIL.n13 VTAIL.n1 0.155672
R199 VTAIL.n22 VTAIL.n17 0.155672
R200 VTAIL.n29 VTAIL.n17 0.155672
R201 VTAIL.n38 VTAIL.n33 0.155672
R202 VTAIL.n45 VTAIL.n33 0.155672
R203 VTAIL.n109 VTAIL.n97 0.155672
R204 VTAIL.n102 VTAIL.n97 0.155672
R205 VTAIL.n93 VTAIL.n81 0.155672
R206 VTAIL.n86 VTAIL.n81 0.155672
R207 VTAIL.n77 VTAIL.n65 0.155672
R208 VTAIL.n70 VTAIL.n65 0.155672
R209 VTAIL.n61 VTAIL.n49 0.155672
R210 VTAIL.n54 VTAIL.n49 0.155672
R211 VDD1 VDD1.n1 107.38
R212 VDD1 VDD1.n0 78.3891
R213 VDD1.n0 VDD1.t0 6.28621
R214 VDD1.n0 VDD1.t3 6.28621
R215 VDD1.n1 VDD1.t1 6.28621
R216 VDD1.n1 VDD1.t2 6.28621
R217 B.n336 B.n335 585
R218 B.n337 B.n336 585
R219 B.n134 B.n52 585
R220 B.n133 B.n132 585
R221 B.n131 B.n130 585
R222 B.n129 B.n128 585
R223 B.n127 B.n126 585
R224 B.n125 B.n124 585
R225 B.n123 B.n122 585
R226 B.n121 B.n120 585
R227 B.n119 B.n118 585
R228 B.n117 B.n116 585
R229 B.n115 B.n114 585
R230 B.n113 B.n112 585
R231 B.n111 B.n110 585
R232 B.n109 B.n108 585
R233 B.n107 B.n106 585
R234 B.n104 B.n103 585
R235 B.n102 B.n101 585
R236 B.n100 B.n99 585
R237 B.n98 B.n97 585
R238 B.n96 B.n95 585
R239 B.n94 B.n93 585
R240 B.n92 B.n91 585
R241 B.n90 B.n89 585
R242 B.n88 B.n87 585
R243 B.n86 B.n85 585
R244 B.n84 B.n83 585
R245 B.n82 B.n81 585
R246 B.n80 B.n79 585
R247 B.n78 B.n77 585
R248 B.n76 B.n75 585
R249 B.n74 B.n73 585
R250 B.n72 B.n71 585
R251 B.n70 B.n69 585
R252 B.n68 B.n67 585
R253 B.n66 B.n65 585
R254 B.n64 B.n63 585
R255 B.n62 B.n61 585
R256 B.n60 B.n59 585
R257 B.n32 B.n31 585
R258 B.n340 B.n339 585
R259 B.n334 B.n53 585
R260 B.n53 B.n29 585
R261 B.n333 B.n28 585
R262 B.n344 B.n28 585
R263 B.n332 B.n27 585
R264 B.n345 B.n27 585
R265 B.n331 B.n26 585
R266 B.n346 B.n26 585
R267 B.n330 B.n329 585
R268 B.n329 B.n25 585
R269 B.n328 B.n21 585
R270 B.n352 B.n21 585
R271 B.n327 B.n20 585
R272 B.n353 B.n20 585
R273 B.n326 B.n19 585
R274 B.n354 B.n19 585
R275 B.n325 B.n324 585
R276 B.n324 B.n15 585
R277 B.n323 B.n14 585
R278 B.n360 B.n14 585
R279 B.n322 B.n13 585
R280 B.n361 B.n13 585
R281 B.n321 B.n12 585
R282 B.n362 B.n12 585
R283 B.n320 B.n319 585
R284 B.n319 B.n11 585
R285 B.n318 B.n7 585
R286 B.n368 B.n7 585
R287 B.n317 B.n6 585
R288 B.n369 B.n6 585
R289 B.n316 B.n5 585
R290 B.n370 B.n5 585
R291 B.n315 B.n314 585
R292 B.n314 B.n4 585
R293 B.n313 B.n135 585
R294 B.n313 B.n312 585
R295 B.n302 B.n136 585
R296 B.n305 B.n136 585
R297 B.n304 B.n303 585
R298 B.n306 B.n304 585
R299 B.n301 B.n141 585
R300 B.n141 B.n140 585
R301 B.n300 B.n299 585
R302 B.n299 B.n298 585
R303 B.n143 B.n142 585
R304 B.n144 B.n143 585
R305 B.n291 B.n290 585
R306 B.n292 B.n291 585
R307 B.n289 B.n149 585
R308 B.n149 B.n148 585
R309 B.n288 B.n287 585
R310 B.n287 B.n286 585
R311 B.n151 B.n150 585
R312 B.n279 B.n151 585
R313 B.n278 B.n277 585
R314 B.n280 B.n278 585
R315 B.n276 B.n156 585
R316 B.n156 B.n155 585
R317 B.n275 B.n274 585
R318 B.n274 B.n273 585
R319 B.n158 B.n157 585
R320 B.n159 B.n158 585
R321 B.n269 B.n268 585
R322 B.n162 B.n161 585
R323 B.n265 B.n264 585
R324 B.n266 B.n265 585
R325 B.n263 B.n182 585
R326 B.n262 B.n261 585
R327 B.n260 B.n259 585
R328 B.n258 B.n257 585
R329 B.n256 B.n255 585
R330 B.n254 B.n253 585
R331 B.n252 B.n251 585
R332 B.n250 B.n249 585
R333 B.n248 B.n247 585
R334 B.n246 B.n245 585
R335 B.n244 B.n243 585
R336 B.n242 B.n241 585
R337 B.n240 B.n239 585
R338 B.n237 B.n236 585
R339 B.n235 B.n234 585
R340 B.n233 B.n232 585
R341 B.n231 B.n230 585
R342 B.n229 B.n228 585
R343 B.n227 B.n226 585
R344 B.n225 B.n224 585
R345 B.n223 B.n222 585
R346 B.n221 B.n220 585
R347 B.n219 B.n218 585
R348 B.n217 B.n216 585
R349 B.n215 B.n214 585
R350 B.n213 B.n212 585
R351 B.n211 B.n210 585
R352 B.n209 B.n208 585
R353 B.n207 B.n206 585
R354 B.n205 B.n204 585
R355 B.n203 B.n202 585
R356 B.n201 B.n200 585
R357 B.n199 B.n198 585
R358 B.n197 B.n196 585
R359 B.n195 B.n194 585
R360 B.n193 B.n192 585
R361 B.n191 B.n190 585
R362 B.n189 B.n188 585
R363 B.n270 B.n160 585
R364 B.n160 B.n159 585
R365 B.n272 B.n271 585
R366 B.n273 B.n272 585
R367 B.n154 B.n153 585
R368 B.n155 B.n154 585
R369 B.n282 B.n281 585
R370 B.n281 B.n280 585
R371 B.n283 B.n152 585
R372 B.n279 B.n152 585
R373 B.n285 B.n284 585
R374 B.n286 B.n285 585
R375 B.n147 B.n146 585
R376 B.n148 B.n147 585
R377 B.n294 B.n293 585
R378 B.n293 B.n292 585
R379 B.n295 B.n145 585
R380 B.n145 B.n144 585
R381 B.n297 B.n296 585
R382 B.n298 B.n297 585
R383 B.n139 B.n138 585
R384 B.n140 B.n139 585
R385 B.n308 B.n307 585
R386 B.n307 B.n306 585
R387 B.n309 B.n137 585
R388 B.n305 B.n137 585
R389 B.n311 B.n310 585
R390 B.n312 B.n311 585
R391 B.n2 B.n0 585
R392 B.n4 B.n2 585
R393 B.n3 B.n1 585
R394 B.n369 B.n3 585
R395 B.n367 B.n366 585
R396 B.n368 B.n367 585
R397 B.n365 B.n8 585
R398 B.n11 B.n8 585
R399 B.n364 B.n363 585
R400 B.n363 B.n362 585
R401 B.n10 B.n9 585
R402 B.n361 B.n10 585
R403 B.n359 B.n358 585
R404 B.n360 B.n359 585
R405 B.n357 B.n16 585
R406 B.n16 B.n15 585
R407 B.n356 B.n355 585
R408 B.n355 B.n354 585
R409 B.n18 B.n17 585
R410 B.n353 B.n18 585
R411 B.n351 B.n350 585
R412 B.n352 B.n351 585
R413 B.n349 B.n22 585
R414 B.n25 B.n22 585
R415 B.n348 B.n347 585
R416 B.n347 B.n346 585
R417 B.n24 B.n23 585
R418 B.n345 B.n24 585
R419 B.n343 B.n342 585
R420 B.n344 B.n343 585
R421 B.n341 B.n30 585
R422 B.n30 B.n29 585
R423 B.n372 B.n371 585
R424 B.n371 B.n370 585
R425 B.n268 B.n160 521.33
R426 B.n339 B.n30 521.33
R427 B.n188 B.n158 521.33
R428 B.n336 B.n53 521.33
R429 B.n185 B.t15 365.067
R430 B.n183 B.t8 365.067
R431 B.n56 B.t12 365.067
R432 B.n54 B.t4 365.067
R433 B.n337 B.n51 256.663
R434 B.n337 B.n50 256.663
R435 B.n337 B.n49 256.663
R436 B.n337 B.n48 256.663
R437 B.n337 B.n47 256.663
R438 B.n337 B.n46 256.663
R439 B.n337 B.n45 256.663
R440 B.n337 B.n44 256.663
R441 B.n337 B.n43 256.663
R442 B.n337 B.n42 256.663
R443 B.n337 B.n41 256.663
R444 B.n337 B.n40 256.663
R445 B.n337 B.n39 256.663
R446 B.n337 B.n38 256.663
R447 B.n337 B.n37 256.663
R448 B.n337 B.n36 256.663
R449 B.n337 B.n35 256.663
R450 B.n337 B.n34 256.663
R451 B.n337 B.n33 256.663
R452 B.n338 B.n337 256.663
R453 B.n267 B.n266 256.663
R454 B.n266 B.n163 256.663
R455 B.n266 B.n164 256.663
R456 B.n266 B.n165 256.663
R457 B.n266 B.n166 256.663
R458 B.n266 B.n167 256.663
R459 B.n266 B.n168 256.663
R460 B.n266 B.n169 256.663
R461 B.n266 B.n170 256.663
R462 B.n266 B.n171 256.663
R463 B.n266 B.n172 256.663
R464 B.n266 B.n173 256.663
R465 B.n266 B.n174 256.663
R466 B.n266 B.n175 256.663
R467 B.n266 B.n176 256.663
R468 B.n266 B.n177 256.663
R469 B.n266 B.n178 256.663
R470 B.n266 B.n179 256.663
R471 B.n266 B.n180 256.663
R472 B.n266 B.n181 256.663
R473 B.n266 B.n159 184.095
R474 B.n337 B.n29 184.095
R475 B.n272 B.n160 163.367
R476 B.n272 B.n154 163.367
R477 B.n281 B.n154 163.367
R478 B.n281 B.n152 163.367
R479 B.n285 B.n152 163.367
R480 B.n285 B.n147 163.367
R481 B.n293 B.n147 163.367
R482 B.n293 B.n145 163.367
R483 B.n297 B.n145 163.367
R484 B.n297 B.n139 163.367
R485 B.n307 B.n139 163.367
R486 B.n307 B.n137 163.367
R487 B.n311 B.n137 163.367
R488 B.n311 B.n2 163.367
R489 B.n371 B.n2 163.367
R490 B.n371 B.n3 163.367
R491 B.n367 B.n3 163.367
R492 B.n367 B.n8 163.367
R493 B.n363 B.n8 163.367
R494 B.n363 B.n10 163.367
R495 B.n359 B.n10 163.367
R496 B.n359 B.n16 163.367
R497 B.n355 B.n16 163.367
R498 B.n355 B.n18 163.367
R499 B.n351 B.n18 163.367
R500 B.n351 B.n22 163.367
R501 B.n347 B.n22 163.367
R502 B.n347 B.n24 163.367
R503 B.n343 B.n24 163.367
R504 B.n343 B.n30 163.367
R505 B.n265 B.n162 163.367
R506 B.n265 B.n182 163.367
R507 B.n261 B.n260 163.367
R508 B.n257 B.n256 163.367
R509 B.n253 B.n252 163.367
R510 B.n249 B.n248 163.367
R511 B.n245 B.n244 163.367
R512 B.n241 B.n240 163.367
R513 B.n236 B.n235 163.367
R514 B.n232 B.n231 163.367
R515 B.n228 B.n227 163.367
R516 B.n224 B.n223 163.367
R517 B.n220 B.n219 163.367
R518 B.n216 B.n215 163.367
R519 B.n212 B.n211 163.367
R520 B.n208 B.n207 163.367
R521 B.n204 B.n203 163.367
R522 B.n200 B.n199 163.367
R523 B.n196 B.n195 163.367
R524 B.n192 B.n191 163.367
R525 B.n274 B.n158 163.367
R526 B.n274 B.n156 163.367
R527 B.n278 B.n156 163.367
R528 B.n278 B.n151 163.367
R529 B.n287 B.n151 163.367
R530 B.n287 B.n149 163.367
R531 B.n291 B.n149 163.367
R532 B.n291 B.n143 163.367
R533 B.n299 B.n143 163.367
R534 B.n299 B.n141 163.367
R535 B.n304 B.n141 163.367
R536 B.n304 B.n136 163.367
R537 B.n313 B.n136 163.367
R538 B.n314 B.n313 163.367
R539 B.n314 B.n5 163.367
R540 B.n6 B.n5 163.367
R541 B.n7 B.n6 163.367
R542 B.n319 B.n7 163.367
R543 B.n319 B.n12 163.367
R544 B.n13 B.n12 163.367
R545 B.n14 B.n13 163.367
R546 B.n324 B.n14 163.367
R547 B.n324 B.n19 163.367
R548 B.n20 B.n19 163.367
R549 B.n21 B.n20 163.367
R550 B.n329 B.n21 163.367
R551 B.n329 B.n26 163.367
R552 B.n27 B.n26 163.367
R553 B.n28 B.n27 163.367
R554 B.n53 B.n28 163.367
R555 B.n59 B.n32 163.367
R556 B.n63 B.n62 163.367
R557 B.n67 B.n66 163.367
R558 B.n71 B.n70 163.367
R559 B.n75 B.n74 163.367
R560 B.n79 B.n78 163.367
R561 B.n83 B.n82 163.367
R562 B.n87 B.n86 163.367
R563 B.n91 B.n90 163.367
R564 B.n95 B.n94 163.367
R565 B.n99 B.n98 163.367
R566 B.n103 B.n102 163.367
R567 B.n108 B.n107 163.367
R568 B.n112 B.n111 163.367
R569 B.n116 B.n115 163.367
R570 B.n120 B.n119 163.367
R571 B.n124 B.n123 163.367
R572 B.n128 B.n127 163.367
R573 B.n132 B.n131 163.367
R574 B.n336 B.n52 163.367
R575 B.n185 B.t17 146.918
R576 B.n54 B.t6 146.918
R577 B.n183 B.t11 146.918
R578 B.n56 B.t13 146.918
R579 B.n186 B.t16 131.209
R580 B.n55 B.t7 131.209
R581 B.n184 B.t10 131.209
R582 B.n57 B.t14 131.209
R583 B.n273 B.n159 88.7839
R584 B.n273 B.n155 88.7839
R585 B.n280 B.n155 88.7839
R586 B.n280 B.n279 88.7839
R587 B.n286 B.n148 88.7839
R588 B.n292 B.n148 88.7839
R589 B.n292 B.n144 88.7839
R590 B.n298 B.n144 88.7839
R591 B.n306 B.n140 88.7839
R592 B.n306 B.n305 88.7839
R593 B.n312 B.n4 88.7839
R594 B.n370 B.n4 88.7839
R595 B.n370 B.n369 88.7839
R596 B.n369 B.n368 88.7839
R597 B.n362 B.n11 88.7839
R598 B.n362 B.n361 88.7839
R599 B.n360 B.n15 88.7839
R600 B.n354 B.n15 88.7839
R601 B.n354 B.n353 88.7839
R602 B.n353 B.n352 88.7839
R603 B.n346 B.n25 88.7839
R604 B.n346 B.n345 88.7839
R605 B.n345 B.n344 88.7839
R606 B.n344 B.n29 88.7839
R607 B.n298 B.t0 73.1162
R608 B.t1 B.n360 73.1162
R609 B.n268 B.n267 71.676
R610 B.n182 B.n163 71.676
R611 B.n260 B.n164 71.676
R612 B.n256 B.n165 71.676
R613 B.n252 B.n166 71.676
R614 B.n248 B.n167 71.676
R615 B.n244 B.n168 71.676
R616 B.n240 B.n169 71.676
R617 B.n235 B.n170 71.676
R618 B.n231 B.n171 71.676
R619 B.n227 B.n172 71.676
R620 B.n223 B.n173 71.676
R621 B.n219 B.n174 71.676
R622 B.n215 B.n175 71.676
R623 B.n211 B.n176 71.676
R624 B.n207 B.n177 71.676
R625 B.n203 B.n178 71.676
R626 B.n199 B.n179 71.676
R627 B.n195 B.n180 71.676
R628 B.n191 B.n181 71.676
R629 B.n339 B.n338 71.676
R630 B.n59 B.n33 71.676
R631 B.n63 B.n34 71.676
R632 B.n67 B.n35 71.676
R633 B.n71 B.n36 71.676
R634 B.n75 B.n37 71.676
R635 B.n79 B.n38 71.676
R636 B.n83 B.n39 71.676
R637 B.n87 B.n40 71.676
R638 B.n91 B.n41 71.676
R639 B.n95 B.n42 71.676
R640 B.n99 B.n43 71.676
R641 B.n103 B.n44 71.676
R642 B.n108 B.n45 71.676
R643 B.n112 B.n46 71.676
R644 B.n116 B.n47 71.676
R645 B.n120 B.n48 71.676
R646 B.n124 B.n49 71.676
R647 B.n128 B.n50 71.676
R648 B.n132 B.n51 71.676
R649 B.n52 B.n51 71.676
R650 B.n131 B.n50 71.676
R651 B.n127 B.n49 71.676
R652 B.n123 B.n48 71.676
R653 B.n119 B.n47 71.676
R654 B.n115 B.n46 71.676
R655 B.n111 B.n45 71.676
R656 B.n107 B.n44 71.676
R657 B.n102 B.n43 71.676
R658 B.n98 B.n42 71.676
R659 B.n94 B.n41 71.676
R660 B.n90 B.n40 71.676
R661 B.n86 B.n39 71.676
R662 B.n82 B.n38 71.676
R663 B.n78 B.n37 71.676
R664 B.n74 B.n36 71.676
R665 B.n70 B.n35 71.676
R666 B.n66 B.n34 71.676
R667 B.n62 B.n33 71.676
R668 B.n338 B.n32 71.676
R669 B.n267 B.n162 71.676
R670 B.n261 B.n163 71.676
R671 B.n257 B.n164 71.676
R672 B.n253 B.n165 71.676
R673 B.n249 B.n166 71.676
R674 B.n245 B.n167 71.676
R675 B.n241 B.n168 71.676
R676 B.n236 B.n169 71.676
R677 B.n232 B.n170 71.676
R678 B.n228 B.n171 71.676
R679 B.n224 B.n172 71.676
R680 B.n220 B.n173 71.676
R681 B.n216 B.n174 71.676
R682 B.n212 B.n175 71.676
R683 B.n208 B.n176 71.676
R684 B.n204 B.n177 71.676
R685 B.n200 B.n178 71.676
R686 B.n196 B.n179 71.676
R687 B.n192 B.n180 71.676
R688 B.n188 B.n181 71.676
R689 B.n312 B.t2 70.505
R690 B.n368 B.t3 70.505
R691 B.n286 B.t9 67.8937
R692 B.n352 B.t5 67.8937
R693 B.n187 B.n186 59.5399
R694 B.n238 B.n184 59.5399
R695 B.n58 B.n57 59.5399
R696 B.n105 B.n55 59.5399
R697 B.n341 B.n340 33.8737
R698 B.n335 B.n334 33.8737
R699 B.n189 B.n157 33.8737
R700 B.n270 B.n269 33.8737
R701 B.n279 B.t9 20.8907
R702 B.n25 B.t5 20.8907
R703 B.n305 B.t2 18.2794
R704 B.n11 B.t3 18.2794
R705 B B.n372 18.0485
R706 B.n186 B.n185 15.7096
R707 B.n184 B.n183 15.7096
R708 B.n57 B.n56 15.7096
R709 B.n55 B.n54 15.7096
R710 B.t0 B.n140 15.6682
R711 B.n361 B.t1 15.6682
R712 B.n340 B.n31 10.6151
R713 B.n60 B.n31 10.6151
R714 B.n61 B.n60 10.6151
R715 B.n64 B.n61 10.6151
R716 B.n65 B.n64 10.6151
R717 B.n68 B.n65 10.6151
R718 B.n69 B.n68 10.6151
R719 B.n72 B.n69 10.6151
R720 B.n73 B.n72 10.6151
R721 B.n76 B.n73 10.6151
R722 B.n77 B.n76 10.6151
R723 B.n80 B.n77 10.6151
R724 B.n81 B.n80 10.6151
R725 B.n84 B.n81 10.6151
R726 B.n85 B.n84 10.6151
R727 B.n89 B.n88 10.6151
R728 B.n92 B.n89 10.6151
R729 B.n93 B.n92 10.6151
R730 B.n96 B.n93 10.6151
R731 B.n97 B.n96 10.6151
R732 B.n100 B.n97 10.6151
R733 B.n101 B.n100 10.6151
R734 B.n104 B.n101 10.6151
R735 B.n109 B.n106 10.6151
R736 B.n110 B.n109 10.6151
R737 B.n113 B.n110 10.6151
R738 B.n114 B.n113 10.6151
R739 B.n117 B.n114 10.6151
R740 B.n118 B.n117 10.6151
R741 B.n121 B.n118 10.6151
R742 B.n122 B.n121 10.6151
R743 B.n125 B.n122 10.6151
R744 B.n126 B.n125 10.6151
R745 B.n129 B.n126 10.6151
R746 B.n130 B.n129 10.6151
R747 B.n133 B.n130 10.6151
R748 B.n134 B.n133 10.6151
R749 B.n335 B.n134 10.6151
R750 B.n275 B.n157 10.6151
R751 B.n276 B.n275 10.6151
R752 B.n277 B.n276 10.6151
R753 B.n277 B.n150 10.6151
R754 B.n288 B.n150 10.6151
R755 B.n289 B.n288 10.6151
R756 B.n290 B.n289 10.6151
R757 B.n290 B.n142 10.6151
R758 B.n300 B.n142 10.6151
R759 B.n301 B.n300 10.6151
R760 B.n303 B.n301 10.6151
R761 B.n303 B.n302 10.6151
R762 B.n302 B.n135 10.6151
R763 B.n315 B.n135 10.6151
R764 B.n316 B.n315 10.6151
R765 B.n317 B.n316 10.6151
R766 B.n318 B.n317 10.6151
R767 B.n320 B.n318 10.6151
R768 B.n321 B.n320 10.6151
R769 B.n322 B.n321 10.6151
R770 B.n323 B.n322 10.6151
R771 B.n325 B.n323 10.6151
R772 B.n326 B.n325 10.6151
R773 B.n327 B.n326 10.6151
R774 B.n328 B.n327 10.6151
R775 B.n330 B.n328 10.6151
R776 B.n331 B.n330 10.6151
R777 B.n332 B.n331 10.6151
R778 B.n333 B.n332 10.6151
R779 B.n334 B.n333 10.6151
R780 B.n269 B.n161 10.6151
R781 B.n264 B.n161 10.6151
R782 B.n264 B.n263 10.6151
R783 B.n263 B.n262 10.6151
R784 B.n262 B.n259 10.6151
R785 B.n259 B.n258 10.6151
R786 B.n258 B.n255 10.6151
R787 B.n255 B.n254 10.6151
R788 B.n254 B.n251 10.6151
R789 B.n251 B.n250 10.6151
R790 B.n250 B.n247 10.6151
R791 B.n247 B.n246 10.6151
R792 B.n246 B.n243 10.6151
R793 B.n243 B.n242 10.6151
R794 B.n242 B.n239 10.6151
R795 B.n237 B.n234 10.6151
R796 B.n234 B.n233 10.6151
R797 B.n233 B.n230 10.6151
R798 B.n230 B.n229 10.6151
R799 B.n229 B.n226 10.6151
R800 B.n226 B.n225 10.6151
R801 B.n225 B.n222 10.6151
R802 B.n222 B.n221 10.6151
R803 B.n218 B.n217 10.6151
R804 B.n217 B.n214 10.6151
R805 B.n214 B.n213 10.6151
R806 B.n213 B.n210 10.6151
R807 B.n210 B.n209 10.6151
R808 B.n209 B.n206 10.6151
R809 B.n206 B.n205 10.6151
R810 B.n205 B.n202 10.6151
R811 B.n202 B.n201 10.6151
R812 B.n201 B.n198 10.6151
R813 B.n198 B.n197 10.6151
R814 B.n197 B.n194 10.6151
R815 B.n194 B.n193 10.6151
R816 B.n193 B.n190 10.6151
R817 B.n190 B.n189 10.6151
R818 B.n271 B.n270 10.6151
R819 B.n271 B.n153 10.6151
R820 B.n282 B.n153 10.6151
R821 B.n283 B.n282 10.6151
R822 B.n284 B.n283 10.6151
R823 B.n284 B.n146 10.6151
R824 B.n294 B.n146 10.6151
R825 B.n295 B.n294 10.6151
R826 B.n296 B.n295 10.6151
R827 B.n296 B.n138 10.6151
R828 B.n308 B.n138 10.6151
R829 B.n309 B.n308 10.6151
R830 B.n310 B.n309 10.6151
R831 B.n310 B.n0 10.6151
R832 B.n366 B.n1 10.6151
R833 B.n366 B.n365 10.6151
R834 B.n365 B.n364 10.6151
R835 B.n364 B.n9 10.6151
R836 B.n358 B.n9 10.6151
R837 B.n358 B.n357 10.6151
R838 B.n357 B.n356 10.6151
R839 B.n356 B.n17 10.6151
R840 B.n350 B.n17 10.6151
R841 B.n350 B.n349 10.6151
R842 B.n349 B.n348 10.6151
R843 B.n348 B.n23 10.6151
R844 B.n342 B.n23 10.6151
R845 B.n342 B.n341 10.6151
R846 B.n88 B.n58 6.5566
R847 B.n105 B.n104 6.5566
R848 B.n238 B.n237 6.5566
R849 B.n221 B.n187 6.5566
R850 B.n85 B.n58 4.05904
R851 B.n106 B.n105 4.05904
R852 B.n239 B.n238 4.05904
R853 B.n218 B.n187 4.05904
R854 B.n372 B.n0 2.81026
R855 B.n372 B.n1 2.81026
R856 VN.n0 VN.t3 261.481
R857 VN.n1 VN.t1 261.481
R858 VN.n0 VN.t2 261.455
R859 VN.n1 VN.t0 261.455
R860 VN VN.n1 103.656
R861 VN VN.n0 70.265
R862 VDD2.n2 VDD2.n0 106.856
R863 VDD2.n2 VDD2.n1 78.3309
R864 VDD2.n1 VDD2.t3 6.28621
R865 VDD2.n1 VDD2.t2 6.28621
R866 VDD2.n0 VDD2.t0 6.28621
R867 VDD2.n0 VDD2.t1 6.28621
R868 VDD2 VDD2.n2 0.0586897
C0 VN VDD2 0.8954f
C1 VN VP 3.03177f
C2 VDD2 VP 0.264745f
C3 VN VDD1 0.151982f
C4 VDD2 VDD1 0.519117f
C5 VP VDD1 1.00751f
C6 VN VTAIL 0.877706f
C7 VDD2 VTAIL 3.09248f
C8 VP VTAIL 0.891812f
C9 VTAIL VDD1 3.05248f
C10 VDD2 B 1.861199f
C11 VDD1 B 3.81694f
C12 VTAIL B 3.519144f
C13 VN B 5.50536f
C14 VP B 3.717188f
C15 VDD2.t0 B 0.054796f
C16 VDD2.t1 B 0.054796f
C17 VDD2.n0 B 0.621534f
C18 VDD2.t3 B 0.054796f
C19 VDD2.t2 B 0.054796f
C20 VDD2.n1 B 0.411724f
C21 VDD2.n2 B 1.79329f
C22 VN.t3 B 0.163679f
C23 VN.t2 B 0.163667f
C24 VN.n0 B 0.169791f
C25 VN.t1 B 0.163679f
C26 VN.t0 B 0.163667f
C27 VN.n1 B 0.486853f
C28 VDD1.t0 B 0.053396f
C29 VDD1.t3 B 0.053396f
C30 VDD1.n0 B 0.401367f
C31 VDD1.t1 B 0.053396f
C32 VDD1.t2 B 0.053396f
C33 VDD1.n1 B 0.62041f
C34 VTAIL.n0 B 0.02175f
C35 VTAIL.n1 B 0.016504f
C36 VTAIL.n2 B 0.008869f
C37 VTAIL.n3 B 0.015721f
C38 VTAIL.n4 B 0.012223f
C39 VTAIL.t3 B 0.035146f
C40 VTAIL.n5 B 0.060436f
C41 VTAIL.n6 B 0.174541f
C42 VTAIL.n7 B 0.008869f
C43 VTAIL.n8 B 0.00939f
C44 VTAIL.n9 B 0.020962f
C45 VTAIL.n10 B 0.042819f
C46 VTAIL.n11 B 0.00939f
C47 VTAIL.n12 B 0.008869f
C48 VTAIL.n13 B 0.038825f
C49 VTAIL.n14 B 0.023717f
C50 VTAIL.n15 B 0.061124f
C51 VTAIL.n16 B 0.02175f
C52 VTAIL.n17 B 0.016504f
C53 VTAIL.n18 B 0.008869f
C54 VTAIL.n19 B 0.015721f
C55 VTAIL.n20 B 0.012223f
C56 VTAIL.t4 B 0.035146f
C57 VTAIL.n21 B 0.060436f
C58 VTAIL.n22 B 0.174541f
C59 VTAIL.n23 B 0.008869f
C60 VTAIL.n24 B 0.00939f
C61 VTAIL.n25 B 0.020962f
C62 VTAIL.n26 B 0.042819f
C63 VTAIL.n27 B 0.00939f
C64 VTAIL.n28 B 0.008869f
C65 VTAIL.n29 B 0.038825f
C66 VTAIL.n30 B 0.023717f
C67 VTAIL.n31 B 0.076597f
C68 VTAIL.n32 B 0.02175f
C69 VTAIL.n33 B 0.016504f
C70 VTAIL.n34 B 0.008869f
C71 VTAIL.n35 B 0.015721f
C72 VTAIL.n36 B 0.012223f
C73 VTAIL.t7 B 0.035146f
C74 VTAIL.n37 B 0.060436f
C75 VTAIL.n38 B 0.174541f
C76 VTAIL.n39 B 0.008869f
C77 VTAIL.n40 B 0.00939f
C78 VTAIL.n41 B 0.020962f
C79 VTAIL.n42 B 0.042819f
C80 VTAIL.n43 B 0.00939f
C81 VTAIL.n44 B 0.008869f
C82 VTAIL.n45 B 0.038825f
C83 VTAIL.n46 B 0.023717f
C84 VTAIL.n47 B 0.457342f
C85 VTAIL.n48 B 0.02175f
C86 VTAIL.n49 B 0.016504f
C87 VTAIL.n50 B 0.008869f
C88 VTAIL.n51 B 0.015721f
C89 VTAIL.n52 B 0.012223f
C90 VTAIL.t0 B 0.035146f
C91 VTAIL.n53 B 0.060436f
C92 VTAIL.n54 B 0.174541f
C93 VTAIL.n55 B 0.008869f
C94 VTAIL.n56 B 0.00939f
C95 VTAIL.n57 B 0.020962f
C96 VTAIL.n58 B 0.042819f
C97 VTAIL.n59 B 0.00939f
C98 VTAIL.n60 B 0.008869f
C99 VTAIL.n61 B 0.038825f
C100 VTAIL.n62 B 0.023717f
C101 VTAIL.n63 B 0.457343f
C102 VTAIL.n64 B 0.02175f
C103 VTAIL.n65 B 0.016504f
C104 VTAIL.n66 B 0.008869f
C105 VTAIL.n67 B 0.015721f
C106 VTAIL.n68 B 0.012223f
C107 VTAIL.t2 B 0.035146f
C108 VTAIL.n69 B 0.060436f
C109 VTAIL.n70 B 0.174541f
C110 VTAIL.n71 B 0.008869f
C111 VTAIL.n72 B 0.00939f
C112 VTAIL.n73 B 0.020962f
C113 VTAIL.n74 B 0.042819f
C114 VTAIL.n75 B 0.00939f
C115 VTAIL.n76 B 0.008869f
C116 VTAIL.n77 B 0.038825f
C117 VTAIL.n78 B 0.023717f
C118 VTAIL.n79 B 0.076597f
C119 VTAIL.n80 B 0.02175f
C120 VTAIL.n81 B 0.016504f
C121 VTAIL.n82 B 0.008869f
C122 VTAIL.n83 B 0.015721f
C123 VTAIL.n84 B 0.012223f
C124 VTAIL.t6 B 0.035146f
C125 VTAIL.n85 B 0.060436f
C126 VTAIL.n86 B 0.174541f
C127 VTAIL.n87 B 0.008869f
C128 VTAIL.n88 B 0.00939f
C129 VTAIL.n89 B 0.020962f
C130 VTAIL.n90 B 0.042819f
C131 VTAIL.n91 B 0.00939f
C132 VTAIL.n92 B 0.008869f
C133 VTAIL.n93 B 0.038825f
C134 VTAIL.n94 B 0.023717f
C135 VTAIL.n95 B 0.076597f
C136 VTAIL.n96 B 0.02175f
C137 VTAIL.n97 B 0.016504f
C138 VTAIL.n98 B 0.008869f
C139 VTAIL.n99 B 0.015721f
C140 VTAIL.n100 B 0.012223f
C141 VTAIL.t5 B 0.035146f
C142 VTAIL.n101 B 0.060436f
C143 VTAIL.n102 B 0.174541f
C144 VTAIL.n103 B 0.008869f
C145 VTAIL.n104 B 0.00939f
C146 VTAIL.n105 B 0.020962f
C147 VTAIL.n106 B 0.042819f
C148 VTAIL.n107 B 0.00939f
C149 VTAIL.n108 B 0.008869f
C150 VTAIL.n109 B 0.038825f
C151 VTAIL.n110 B 0.023717f
C152 VTAIL.n111 B 0.457342f
C153 VTAIL.n112 B 0.02175f
C154 VTAIL.n113 B 0.016504f
C155 VTAIL.n114 B 0.008869f
C156 VTAIL.n115 B 0.015721f
C157 VTAIL.n116 B 0.012223f
C158 VTAIL.t1 B 0.035146f
C159 VTAIL.n117 B 0.060436f
C160 VTAIL.n118 B 0.174541f
C161 VTAIL.n119 B 0.008869f
C162 VTAIL.n120 B 0.00939f
C163 VTAIL.n121 B 0.020962f
C164 VTAIL.n122 B 0.042819f
C165 VTAIL.n123 B 0.00939f
C166 VTAIL.n124 B 0.008869f
C167 VTAIL.n125 B 0.038825f
C168 VTAIL.n126 B 0.023717f
C169 VTAIL.n127 B 0.435681f
C170 VP.t0 B 0.16636f
C171 VP.t3 B 0.166372f
C172 VP.n0 B 0.484864f
C173 VP.n1 B 1.6358f
C174 VP.t2 B 0.158844f
C175 VP.n2 B 0.093765f
C176 VP.t1 B 0.158844f
C177 VP.n3 B 0.093765f
C178 VP.n4 B 0.027208f
.ends

