* NGSPICE file created from diff_pair_sample_0821.ext - technology: sky130A

.subckt diff_pair_sample_0821 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.7527 ps=4.64 w=1.93 l=0.65
X1 VTAIL.t9 VP.t1 VDD1.t8 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X2 B.t11 B.t9 B.t10 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0 ps=0 w=1.93 l=0.65
X3 VTAIL.t18 VN.t0 VDD2.t9 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X4 B.t8 B.t6 B.t7 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0 ps=0 w=1.93 l=0.65
X5 B.t5 B.t3 B.t4 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0 ps=0 w=1.93 l=0.65
X6 VDD1.t7 VP.t2 VTAIL.t14 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0.31845 ps=2.26 w=1.93 l=0.65
X7 VDD2.t8 VN.t1 VTAIL.t19 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0.31845 ps=2.26 w=1.93 l=0.65
X8 VDD1.t6 VP.t3 VTAIL.t16 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0.31845 ps=2.26 w=1.93 l=0.65
X9 VTAIL.t15 VP.t4 VDD1.t5 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X10 VDD2.t7 VN.t2 VTAIL.t4 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.7527 ps=4.64 w=1.93 l=0.65
X11 VDD2.t6 VN.t3 VTAIL.t3 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.7527 ps=4.64 w=1.93 l=0.65
X12 VDD1.t4 VP.t5 VTAIL.t13 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X13 VDD2.t5 VN.t4 VTAIL.t6 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X14 VTAIL.t1 VN.t5 VDD2.t4 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X15 B.t2 B.t0 B.t1 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0 ps=0 w=1.93 l=0.65
X16 VDD1.t3 VP.t6 VTAIL.t10 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X17 VDD1.t2 VP.t7 VTAIL.t7 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.7527 ps=4.64 w=1.93 l=0.65
X18 VDD2.t3 VN.t6 VTAIL.t2 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.7527 pd=4.64 as=0.31845 ps=2.26 w=1.93 l=0.65
X19 VTAIL.t5 VN.t7 VDD2.t2 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X20 VDD2.t1 VN.t8 VTAIL.t0 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X21 VTAIL.t11 VP.t8 VDD1.t1 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X22 VTAIL.t8 VP.t9 VDD1.t0 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
X23 VTAIL.t17 VN.t9 VDD2.t0 w_n2146_n1354# sky130_fd_pr__pfet_01v8 ad=0.31845 pd=2.26 as=0.31845 ps=2.26 w=1.93 l=0.65
R0 VP.n17 VP.n16 161.3
R1 VP.n9 VP.n8 161.3
R2 VP.n11 VP.n10 161.3
R3 VP.n4 VP.t2 159.186
R4 VP.n10 VP.t3 132.365
R5 VP.n1 VP.t1 132.365
R6 VP.n14 VP.t5 132.365
R7 VP.n15 VP.t8 132.365
R8 VP.n16 VP.t7 132.365
R9 VP.n8 VP.t0 132.365
R10 VP.n7 VP.t4 132.365
R11 VP.n6 VP.t6 132.365
R12 VP.n5 VP.t9 132.365
R13 VP.n6 VP.n3 80.6037
R14 VP.n7 VP.n2 80.6037
R15 VP.n15 VP.n0 80.6037
R16 VP.n14 VP.n13 80.6037
R17 VP.n12 VP.n1 80.6037
R18 VP.n10 VP.n1 48.2005
R19 VP.n14 VP.n1 48.2005
R20 VP.n15 VP.n14 48.2005
R21 VP.n16 VP.n15 48.2005
R22 VP.n8 VP.n7 48.2005
R23 VP.n7 VP.n6 48.2005
R24 VP.n6 VP.n5 48.2005
R25 VP.n4 VP.n3 45.2318
R26 VP.n11 VP.n9 34.9853
R27 VP.n5 VP.n4 13.3799
R28 VP.n3 VP.n2 0.380177
R29 VP.n13 VP.n12 0.380177
R30 VP.n13 VP.n0 0.380177
R31 VP.n9 VP.n2 0.285035
R32 VP.n12 VP.n11 0.285035
R33 VP.n17 VP.n0 0.285035
R34 VP VP.n17 0.0516364
R35 VTAIL.n40 VTAIL.n38 756.745
R36 VTAIL.n4 VTAIL.n2 756.745
R37 VTAIL.n32 VTAIL.n30 756.745
R38 VTAIL.n20 VTAIL.n18 756.745
R39 VTAIL.n41 VTAIL.n40 585
R40 VTAIL.n5 VTAIL.n4 585
R41 VTAIL.n33 VTAIL.n32 585
R42 VTAIL.n21 VTAIL.n20 585
R43 VTAIL.t4 VTAIL.n39 417.779
R44 VTAIL.t7 VTAIL.n3 417.779
R45 VTAIL.t12 VTAIL.n31 417.779
R46 VTAIL.t3 VTAIL.n19 417.779
R47 VTAIL.n29 VTAIL.n28 182.794
R48 VTAIL.n27 VTAIL.n26 182.794
R49 VTAIL.n17 VTAIL.n16 182.794
R50 VTAIL.n15 VTAIL.n14 182.794
R51 VTAIL.n47 VTAIL.n46 182.794
R52 VTAIL.n1 VTAIL.n0 182.794
R53 VTAIL.n11 VTAIL.n10 182.794
R54 VTAIL.n13 VTAIL.n12 182.794
R55 VTAIL.n40 VTAIL.t4 85.8723
R56 VTAIL.n4 VTAIL.t7 85.8723
R57 VTAIL.n32 VTAIL.t12 85.8723
R58 VTAIL.n20 VTAIL.t3 85.8723
R59 VTAIL.n45 VTAIL.n44 30.052
R60 VTAIL.n9 VTAIL.n8 30.052
R61 VTAIL.n37 VTAIL.n36 30.052
R62 VTAIL.n25 VTAIL.n24 30.052
R63 VTAIL.n46 VTAIL.t6 16.8425
R64 VTAIL.n46 VTAIL.t5 16.8425
R65 VTAIL.n0 VTAIL.t2 16.8425
R66 VTAIL.n0 VTAIL.t17 16.8425
R67 VTAIL.n10 VTAIL.t13 16.8425
R68 VTAIL.n10 VTAIL.t11 16.8425
R69 VTAIL.n12 VTAIL.t16 16.8425
R70 VTAIL.n12 VTAIL.t9 16.8425
R71 VTAIL.n28 VTAIL.t10 16.8425
R72 VTAIL.n28 VTAIL.t15 16.8425
R73 VTAIL.n26 VTAIL.t14 16.8425
R74 VTAIL.n26 VTAIL.t8 16.8425
R75 VTAIL.n16 VTAIL.t0 16.8425
R76 VTAIL.n16 VTAIL.t18 16.8425
R77 VTAIL.n14 VTAIL.t19 16.8425
R78 VTAIL.n14 VTAIL.t1 16.8425
R79 VTAIL.n15 VTAIL.n13 15.7203
R80 VTAIL.n45 VTAIL.n37 14.8755
R81 VTAIL.n41 VTAIL.n39 9.84608
R82 VTAIL.n5 VTAIL.n3 9.84608
R83 VTAIL.n33 VTAIL.n31 9.84608
R84 VTAIL.n21 VTAIL.n19 9.84608
R85 VTAIL.n44 VTAIL.n43 9.45567
R86 VTAIL.n8 VTAIL.n7 9.45567
R87 VTAIL.n36 VTAIL.n35 9.45567
R88 VTAIL.n24 VTAIL.n23 9.45567
R89 VTAIL.n43 VTAIL.n42 9.3005
R90 VTAIL.n7 VTAIL.n6 9.3005
R91 VTAIL.n35 VTAIL.n34 9.3005
R92 VTAIL.n23 VTAIL.n22 9.3005
R93 VTAIL.n44 VTAIL.n38 8.14595
R94 VTAIL.n8 VTAIL.n2 8.14595
R95 VTAIL.n36 VTAIL.n30 8.14595
R96 VTAIL.n24 VTAIL.n18 8.14595
R97 VTAIL.n42 VTAIL.n41 7.3702
R98 VTAIL.n6 VTAIL.n5 7.3702
R99 VTAIL.n34 VTAIL.n33 7.3702
R100 VTAIL.n22 VTAIL.n21 7.3702
R101 VTAIL.n42 VTAIL.n38 5.81868
R102 VTAIL.n6 VTAIL.n2 5.81868
R103 VTAIL.n34 VTAIL.n30 5.81868
R104 VTAIL.n22 VTAIL.n18 5.81868
R105 VTAIL.n23 VTAIL.n19 3.32369
R106 VTAIL.n43 VTAIL.n39 3.32369
R107 VTAIL.n7 VTAIL.n3 3.32369
R108 VTAIL.n35 VTAIL.n31 3.32369
R109 VTAIL.n27 VTAIL.n25 0.892741
R110 VTAIL.n9 VTAIL.n1 0.892741
R111 VTAIL.n17 VTAIL.n15 0.845328
R112 VTAIL.n25 VTAIL.n17 0.845328
R113 VTAIL.n29 VTAIL.n27 0.845328
R114 VTAIL.n37 VTAIL.n29 0.845328
R115 VTAIL.n13 VTAIL.n11 0.845328
R116 VTAIL.n11 VTAIL.n9 0.845328
R117 VTAIL.n47 VTAIL.n45 0.845328
R118 VTAIL VTAIL.n1 0.69231
R119 VTAIL VTAIL.n47 0.153517
R120 VDD1.n2 VDD1.n0 756.745
R121 VDD1.n11 VDD1.n9 756.745
R122 VDD1.n3 VDD1.n2 585
R123 VDD1.n12 VDD1.n11 585
R124 VDD1.t6 VDD1.n10 417.779
R125 VDD1.t7 VDD1.n1 417.779
R126 VDD1.n19 VDD1.n18 200.052
R127 VDD1.n21 VDD1.n20 199.474
R128 VDD1.n8 VDD1.n7 199.474
R129 VDD1.n17 VDD1.n16 199.474
R130 VDD1.n2 VDD1.t7 85.8723
R131 VDD1.n11 VDD1.t6 85.8723
R132 VDD1.n8 VDD1.n6 47.5756
R133 VDD1.n17 VDD1.n15 47.5756
R134 VDD1.n21 VDD1.n19 30.3974
R135 VDD1.n20 VDD1.t5 16.8425
R136 VDD1.n20 VDD1.t9 16.8425
R137 VDD1.n7 VDD1.t0 16.8425
R138 VDD1.n7 VDD1.t3 16.8425
R139 VDD1.n18 VDD1.t1 16.8425
R140 VDD1.n18 VDD1.t2 16.8425
R141 VDD1.n16 VDD1.t8 16.8425
R142 VDD1.n16 VDD1.t4 16.8425
R143 VDD1.n3 VDD1.n1 9.84608
R144 VDD1.n12 VDD1.n10 9.84608
R145 VDD1.n6 VDD1.n5 9.45567
R146 VDD1.n15 VDD1.n14 9.45567
R147 VDD1.n5 VDD1.n4 9.3005
R148 VDD1.n14 VDD1.n13 9.3005
R149 VDD1.n6 VDD1.n0 8.14595
R150 VDD1.n15 VDD1.n9 8.14595
R151 VDD1.n4 VDD1.n3 7.3702
R152 VDD1.n13 VDD1.n12 7.3702
R153 VDD1.n4 VDD1.n0 5.81868
R154 VDD1.n13 VDD1.n9 5.81868
R155 VDD1.n5 VDD1.n1 3.32369
R156 VDD1.n14 VDD1.n10 3.32369
R157 VDD1 VDD1.n21 0.575931
R158 VDD1 VDD1.n8 0.269897
R159 VDD1.n19 VDD1.n17 0.156361
R160 B.n184 B.n183 585
R161 B.n182 B.n63 585
R162 B.n181 B.n180 585
R163 B.n179 B.n64 585
R164 B.n178 B.n177 585
R165 B.n176 B.n65 585
R166 B.n175 B.n174 585
R167 B.n173 B.n66 585
R168 B.n172 B.n171 585
R169 B.n170 B.n67 585
R170 B.n169 B.n168 585
R171 B.n167 B.n68 585
R172 B.n165 B.n164 585
R173 B.n163 B.n71 585
R174 B.n162 B.n161 585
R175 B.n160 B.n72 585
R176 B.n159 B.n158 585
R177 B.n157 B.n73 585
R178 B.n156 B.n155 585
R179 B.n154 B.n74 585
R180 B.n153 B.n152 585
R181 B.n151 B.n75 585
R182 B.n150 B.n149 585
R183 B.n145 B.n76 585
R184 B.n144 B.n143 585
R185 B.n142 B.n77 585
R186 B.n141 B.n140 585
R187 B.n139 B.n78 585
R188 B.n138 B.n137 585
R189 B.n136 B.n79 585
R190 B.n135 B.n134 585
R191 B.n133 B.n80 585
R192 B.n132 B.n131 585
R193 B.n130 B.n81 585
R194 B.n185 B.n62 585
R195 B.n187 B.n186 585
R196 B.n188 B.n61 585
R197 B.n190 B.n189 585
R198 B.n191 B.n60 585
R199 B.n193 B.n192 585
R200 B.n194 B.n59 585
R201 B.n196 B.n195 585
R202 B.n197 B.n58 585
R203 B.n199 B.n198 585
R204 B.n200 B.n57 585
R205 B.n202 B.n201 585
R206 B.n203 B.n56 585
R207 B.n205 B.n204 585
R208 B.n206 B.n55 585
R209 B.n208 B.n207 585
R210 B.n209 B.n54 585
R211 B.n211 B.n210 585
R212 B.n212 B.n53 585
R213 B.n214 B.n213 585
R214 B.n215 B.n52 585
R215 B.n217 B.n216 585
R216 B.n218 B.n51 585
R217 B.n220 B.n219 585
R218 B.n221 B.n50 585
R219 B.n223 B.n222 585
R220 B.n224 B.n49 585
R221 B.n226 B.n225 585
R222 B.n227 B.n48 585
R223 B.n229 B.n228 585
R224 B.n230 B.n47 585
R225 B.n232 B.n231 585
R226 B.n233 B.n46 585
R227 B.n235 B.n234 585
R228 B.n236 B.n45 585
R229 B.n238 B.n237 585
R230 B.n239 B.n44 585
R231 B.n241 B.n240 585
R232 B.n242 B.n43 585
R233 B.n244 B.n243 585
R234 B.n245 B.n42 585
R235 B.n247 B.n246 585
R236 B.n248 B.n41 585
R237 B.n250 B.n249 585
R238 B.n251 B.n40 585
R239 B.n253 B.n252 585
R240 B.n254 B.n39 585
R241 B.n256 B.n255 585
R242 B.n257 B.n38 585
R243 B.n259 B.n258 585
R244 B.n260 B.n37 585
R245 B.n262 B.n261 585
R246 B.n314 B.n313 585
R247 B.n312 B.n15 585
R248 B.n311 B.n310 585
R249 B.n309 B.n16 585
R250 B.n308 B.n307 585
R251 B.n306 B.n17 585
R252 B.n305 B.n304 585
R253 B.n303 B.n18 585
R254 B.n302 B.n301 585
R255 B.n300 B.n19 585
R256 B.n299 B.n298 585
R257 B.n297 B.n20 585
R258 B.n296 B.n295 585
R259 B.n294 B.n21 585
R260 B.n293 B.n292 585
R261 B.n291 B.n25 585
R262 B.n290 B.n289 585
R263 B.n288 B.n26 585
R264 B.n287 B.n286 585
R265 B.n285 B.n27 585
R266 B.n284 B.n283 585
R267 B.n282 B.n28 585
R268 B.n280 B.n279 585
R269 B.n278 B.n31 585
R270 B.n277 B.n276 585
R271 B.n275 B.n32 585
R272 B.n274 B.n273 585
R273 B.n272 B.n33 585
R274 B.n271 B.n270 585
R275 B.n269 B.n34 585
R276 B.n268 B.n267 585
R277 B.n266 B.n35 585
R278 B.n265 B.n264 585
R279 B.n263 B.n36 585
R280 B.n315 B.n14 585
R281 B.n317 B.n316 585
R282 B.n318 B.n13 585
R283 B.n320 B.n319 585
R284 B.n321 B.n12 585
R285 B.n323 B.n322 585
R286 B.n324 B.n11 585
R287 B.n326 B.n325 585
R288 B.n327 B.n10 585
R289 B.n329 B.n328 585
R290 B.n330 B.n9 585
R291 B.n332 B.n331 585
R292 B.n333 B.n8 585
R293 B.n335 B.n334 585
R294 B.n336 B.n7 585
R295 B.n338 B.n337 585
R296 B.n339 B.n6 585
R297 B.n341 B.n340 585
R298 B.n342 B.n5 585
R299 B.n344 B.n343 585
R300 B.n345 B.n4 585
R301 B.n347 B.n346 585
R302 B.n348 B.n3 585
R303 B.n350 B.n349 585
R304 B.n351 B.n0 585
R305 B.n2 B.n1 585
R306 B.n94 B.n93 585
R307 B.n96 B.n95 585
R308 B.n97 B.n92 585
R309 B.n99 B.n98 585
R310 B.n100 B.n91 585
R311 B.n102 B.n101 585
R312 B.n103 B.n90 585
R313 B.n105 B.n104 585
R314 B.n106 B.n89 585
R315 B.n108 B.n107 585
R316 B.n109 B.n88 585
R317 B.n111 B.n110 585
R318 B.n112 B.n87 585
R319 B.n114 B.n113 585
R320 B.n115 B.n86 585
R321 B.n117 B.n116 585
R322 B.n118 B.n85 585
R323 B.n120 B.n119 585
R324 B.n121 B.n84 585
R325 B.n123 B.n122 585
R326 B.n124 B.n83 585
R327 B.n126 B.n125 585
R328 B.n127 B.n82 585
R329 B.n129 B.n128 585
R330 B.n130 B.n129 449.257
R331 B.n183 B.n62 449.257
R332 B.n261 B.n36 449.257
R333 B.n315 B.n314 449.257
R334 B.n146 B.t3 275.185
R335 B.n69 B.t9 275.185
R336 B.n29 B.t6 275.185
R337 B.n22 B.t0 275.185
R338 B.n69 B.t10 265.986
R339 B.n29 B.t8 265.986
R340 B.n146 B.t4 265.986
R341 B.n22 B.t2 265.986
R342 B.n353 B.n352 256.663
R343 B.n70 B.t11 246.981
R344 B.n30 B.t7 246.981
R345 B.n147 B.t5 246.98
R346 B.n23 B.t1 246.98
R347 B.n352 B.n351 235.042
R348 B.n352 B.n2 235.042
R349 B.n131 B.n130 163.367
R350 B.n131 B.n80 163.367
R351 B.n135 B.n80 163.367
R352 B.n136 B.n135 163.367
R353 B.n137 B.n136 163.367
R354 B.n137 B.n78 163.367
R355 B.n141 B.n78 163.367
R356 B.n142 B.n141 163.367
R357 B.n143 B.n142 163.367
R358 B.n143 B.n76 163.367
R359 B.n150 B.n76 163.367
R360 B.n151 B.n150 163.367
R361 B.n152 B.n151 163.367
R362 B.n152 B.n74 163.367
R363 B.n156 B.n74 163.367
R364 B.n157 B.n156 163.367
R365 B.n158 B.n157 163.367
R366 B.n158 B.n72 163.367
R367 B.n162 B.n72 163.367
R368 B.n163 B.n162 163.367
R369 B.n164 B.n163 163.367
R370 B.n164 B.n68 163.367
R371 B.n169 B.n68 163.367
R372 B.n170 B.n169 163.367
R373 B.n171 B.n170 163.367
R374 B.n171 B.n66 163.367
R375 B.n175 B.n66 163.367
R376 B.n176 B.n175 163.367
R377 B.n177 B.n176 163.367
R378 B.n177 B.n64 163.367
R379 B.n181 B.n64 163.367
R380 B.n182 B.n181 163.367
R381 B.n183 B.n182 163.367
R382 B.n261 B.n260 163.367
R383 B.n260 B.n259 163.367
R384 B.n259 B.n38 163.367
R385 B.n255 B.n38 163.367
R386 B.n255 B.n254 163.367
R387 B.n254 B.n253 163.367
R388 B.n253 B.n40 163.367
R389 B.n249 B.n40 163.367
R390 B.n249 B.n248 163.367
R391 B.n248 B.n247 163.367
R392 B.n247 B.n42 163.367
R393 B.n243 B.n42 163.367
R394 B.n243 B.n242 163.367
R395 B.n242 B.n241 163.367
R396 B.n241 B.n44 163.367
R397 B.n237 B.n44 163.367
R398 B.n237 B.n236 163.367
R399 B.n236 B.n235 163.367
R400 B.n235 B.n46 163.367
R401 B.n231 B.n46 163.367
R402 B.n231 B.n230 163.367
R403 B.n230 B.n229 163.367
R404 B.n229 B.n48 163.367
R405 B.n225 B.n48 163.367
R406 B.n225 B.n224 163.367
R407 B.n224 B.n223 163.367
R408 B.n223 B.n50 163.367
R409 B.n219 B.n50 163.367
R410 B.n219 B.n218 163.367
R411 B.n218 B.n217 163.367
R412 B.n217 B.n52 163.367
R413 B.n213 B.n52 163.367
R414 B.n213 B.n212 163.367
R415 B.n212 B.n211 163.367
R416 B.n211 B.n54 163.367
R417 B.n207 B.n54 163.367
R418 B.n207 B.n206 163.367
R419 B.n206 B.n205 163.367
R420 B.n205 B.n56 163.367
R421 B.n201 B.n56 163.367
R422 B.n201 B.n200 163.367
R423 B.n200 B.n199 163.367
R424 B.n199 B.n58 163.367
R425 B.n195 B.n58 163.367
R426 B.n195 B.n194 163.367
R427 B.n194 B.n193 163.367
R428 B.n193 B.n60 163.367
R429 B.n189 B.n60 163.367
R430 B.n189 B.n188 163.367
R431 B.n188 B.n187 163.367
R432 B.n187 B.n62 163.367
R433 B.n314 B.n15 163.367
R434 B.n310 B.n15 163.367
R435 B.n310 B.n309 163.367
R436 B.n309 B.n308 163.367
R437 B.n308 B.n17 163.367
R438 B.n304 B.n17 163.367
R439 B.n304 B.n303 163.367
R440 B.n303 B.n302 163.367
R441 B.n302 B.n19 163.367
R442 B.n298 B.n19 163.367
R443 B.n298 B.n297 163.367
R444 B.n297 B.n296 163.367
R445 B.n296 B.n21 163.367
R446 B.n292 B.n21 163.367
R447 B.n292 B.n291 163.367
R448 B.n291 B.n290 163.367
R449 B.n290 B.n26 163.367
R450 B.n286 B.n26 163.367
R451 B.n286 B.n285 163.367
R452 B.n285 B.n284 163.367
R453 B.n284 B.n28 163.367
R454 B.n279 B.n28 163.367
R455 B.n279 B.n278 163.367
R456 B.n278 B.n277 163.367
R457 B.n277 B.n32 163.367
R458 B.n273 B.n32 163.367
R459 B.n273 B.n272 163.367
R460 B.n272 B.n271 163.367
R461 B.n271 B.n34 163.367
R462 B.n267 B.n34 163.367
R463 B.n267 B.n266 163.367
R464 B.n266 B.n265 163.367
R465 B.n265 B.n36 163.367
R466 B.n316 B.n315 163.367
R467 B.n316 B.n13 163.367
R468 B.n320 B.n13 163.367
R469 B.n321 B.n320 163.367
R470 B.n322 B.n321 163.367
R471 B.n322 B.n11 163.367
R472 B.n326 B.n11 163.367
R473 B.n327 B.n326 163.367
R474 B.n328 B.n327 163.367
R475 B.n328 B.n9 163.367
R476 B.n332 B.n9 163.367
R477 B.n333 B.n332 163.367
R478 B.n334 B.n333 163.367
R479 B.n334 B.n7 163.367
R480 B.n338 B.n7 163.367
R481 B.n339 B.n338 163.367
R482 B.n340 B.n339 163.367
R483 B.n340 B.n5 163.367
R484 B.n344 B.n5 163.367
R485 B.n345 B.n344 163.367
R486 B.n346 B.n345 163.367
R487 B.n346 B.n3 163.367
R488 B.n350 B.n3 163.367
R489 B.n351 B.n350 163.367
R490 B.n94 B.n2 163.367
R491 B.n95 B.n94 163.367
R492 B.n95 B.n92 163.367
R493 B.n99 B.n92 163.367
R494 B.n100 B.n99 163.367
R495 B.n101 B.n100 163.367
R496 B.n101 B.n90 163.367
R497 B.n105 B.n90 163.367
R498 B.n106 B.n105 163.367
R499 B.n107 B.n106 163.367
R500 B.n107 B.n88 163.367
R501 B.n111 B.n88 163.367
R502 B.n112 B.n111 163.367
R503 B.n113 B.n112 163.367
R504 B.n113 B.n86 163.367
R505 B.n117 B.n86 163.367
R506 B.n118 B.n117 163.367
R507 B.n119 B.n118 163.367
R508 B.n119 B.n84 163.367
R509 B.n123 B.n84 163.367
R510 B.n124 B.n123 163.367
R511 B.n125 B.n124 163.367
R512 B.n125 B.n82 163.367
R513 B.n129 B.n82 163.367
R514 B.n148 B.n147 59.5399
R515 B.n166 B.n70 59.5399
R516 B.n281 B.n30 59.5399
R517 B.n24 B.n23 59.5399
R518 B.n185 B.n184 29.1907
R519 B.n313 B.n14 29.1907
R520 B.n263 B.n262 29.1907
R521 B.n128 B.n81 29.1907
R522 B.n147 B.n146 19.0066
R523 B.n70 B.n69 19.0066
R524 B.n30 B.n29 19.0066
R525 B.n23 B.n22 19.0066
R526 B B.n353 18.0485
R527 B.n317 B.n14 10.6151
R528 B.n318 B.n317 10.6151
R529 B.n319 B.n318 10.6151
R530 B.n319 B.n12 10.6151
R531 B.n323 B.n12 10.6151
R532 B.n324 B.n323 10.6151
R533 B.n325 B.n324 10.6151
R534 B.n325 B.n10 10.6151
R535 B.n329 B.n10 10.6151
R536 B.n330 B.n329 10.6151
R537 B.n331 B.n330 10.6151
R538 B.n331 B.n8 10.6151
R539 B.n335 B.n8 10.6151
R540 B.n336 B.n335 10.6151
R541 B.n337 B.n336 10.6151
R542 B.n337 B.n6 10.6151
R543 B.n341 B.n6 10.6151
R544 B.n342 B.n341 10.6151
R545 B.n343 B.n342 10.6151
R546 B.n343 B.n4 10.6151
R547 B.n347 B.n4 10.6151
R548 B.n348 B.n347 10.6151
R549 B.n349 B.n348 10.6151
R550 B.n349 B.n0 10.6151
R551 B.n313 B.n312 10.6151
R552 B.n312 B.n311 10.6151
R553 B.n311 B.n16 10.6151
R554 B.n307 B.n16 10.6151
R555 B.n307 B.n306 10.6151
R556 B.n306 B.n305 10.6151
R557 B.n305 B.n18 10.6151
R558 B.n301 B.n18 10.6151
R559 B.n301 B.n300 10.6151
R560 B.n300 B.n299 10.6151
R561 B.n299 B.n20 10.6151
R562 B.n295 B.n294 10.6151
R563 B.n294 B.n293 10.6151
R564 B.n293 B.n25 10.6151
R565 B.n289 B.n25 10.6151
R566 B.n289 B.n288 10.6151
R567 B.n288 B.n287 10.6151
R568 B.n287 B.n27 10.6151
R569 B.n283 B.n27 10.6151
R570 B.n283 B.n282 10.6151
R571 B.n280 B.n31 10.6151
R572 B.n276 B.n31 10.6151
R573 B.n276 B.n275 10.6151
R574 B.n275 B.n274 10.6151
R575 B.n274 B.n33 10.6151
R576 B.n270 B.n33 10.6151
R577 B.n270 B.n269 10.6151
R578 B.n269 B.n268 10.6151
R579 B.n268 B.n35 10.6151
R580 B.n264 B.n35 10.6151
R581 B.n264 B.n263 10.6151
R582 B.n262 B.n37 10.6151
R583 B.n258 B.n37 10.6151
R584 B.n258 B.n257 10.6151
R585 B.n257 B.n256 10.6151
R586 B.n256 B.n39 10.6151
R587 B.n252 B.n39 10.6151
R588 B.n252 B.n251 10.6151
R589 B.n251 B.n250 10.6151
R590 B.n250 B.n41 10.6151
R591 B.n246 B.n41 10.6151
R592 B.n246 B.n245 10.6151
R593 B.n245 B.n244 10.6151
R594 B.n244 B.n43 10.6151
R595 B.n240 B.n43 10.6151
R596 B.n240 B.n239 10.6151
R597 B.n239 B.n238 10.6151
R598 B.n238 B.n45 10.6151
R599 B.n234 B.n45 10.6151
R600 B.n234 B.n233 10.6151
R601 B.n233 B.n232 10.6151
R602 B.n232 B.n47 10.6151
R603 B.n228 B.n47 10.6151
R604 B.n228 B.n227 10.6151
R605 B.n227 B.n226 10.6151
R606 B.n226 B.n49 10.6151
R607 B.n222 B.n49 10.6151
R608 B.n222 B.n221 10.6151
R609 B.n221 B.n220 10.6151
R610 B.n220 B.n51 10.6151
R611 B.n216 B.n51 10.6151
R612 B.n216 B.n215 10.6151
R613 B.n215 B.n214 10.6151
R614 B.n214 B.n53 10.6151
R615 B.n210 B.n53 10.6151
R616 B.n210 B.n209 10.6151
R617 B.n209 B.n208 10.6151
R618 B.n208 B.n55 10.6151
R619 B.n204 B.n55 10.6151
R620 B.n204 B.n203 10.6151
R621 B.n203 B.n202 10.6151
R622 B.n202 B.n57 10.6151
R623 B.n198 B.n57 10.6151
R624 B.n198 B.n197 10.6151
R625 B.n197 B.n196 10.6151
R626 B.n196 B.n59 10.6151
R627 B.n192 B.n59 10.6151
R628 B.n192 B.n191 10.6151
R629 B.n191 B.n190 10.6151
R630 B.n190 B.n61 10.6151
R631 B.n186 B.n61 10.6151
R632 B.n186 B.n185 10.6151
R633 B.n93 B.n1 10.6151
R634 B.n96 B.n93 10.6151
R635 B.n97 B.n96 10.6151
R636 B.n98 B.n97 10.6151
R637 B.n98 B.n91 10.6151
R638 B.n102 B.n91 10.6151
R639 B.n103 B.n102 10.6151
R640 B.n104 B.n103 10.6151
R641 B.n104 B.n89 10.6151
R642 B.n108 B.n89 10.6151
R643 B.n109 B.n108 10.6151
R644 B.n110 B.n109 10.6151
R645 B.n110 B.n87 10.6151
R646 B.n114 B.n87 10.6151
R647 B.n115 B.n114 10.6151
R648 B.n116 B.n115 10.6151
R649 B.n116 B.n85 10.6151
R650 B.n120 B.n85 10.6151
R651 B.n121 B.n120 10.6151
R652 B.n122 B.n121 10.6151
R653 B.n122 B.n83 10.6151
R654 B.n126 B.n83 10.6151
R655 B.n127 B.n126 10.6151
R656 B.n128 B.n127 10.6151
R657 B.n132 B.n81 10.6151
R658 B.n133 B.n132 10.6151
R659 B.n134 B.n133 10.6151
R660 B.n134 B.n79 10.6151
R661 B.n138 B.n79 10.6151
R662 B.n139 B.n138 10.6151
R663 B.n140 B.n139 10.6151
R664 B.n140 B.n77 10.6151
R665 B.n144 B.n77 10.6151
R666 B.n145 B.n144 10.6151
R667 B.n149 B.n145 10.6151
R668 B.n153 B.n75 10.6151
R669 B.n154 B.n153 10.6151
R670 B.n155 B.n154 10.6151
R671 B.n155 B.n73 10.6151
R672 B.n159 B.n73 10.6151
R673 B.n160 B.n159 10.6151
R674 B.n161 B.n160 10.6151
R675 B.n161 B.n71 10.6151
R676 B.n165 B.n71 10.6151
R677 B.n168 B.n167 10.6151
R678 B.n168 B.n67 10.6151
R679 B.n172 B.n67 10.6151
R680 B.n173 B.n172 10.6151
R681 B.n174 B.n173 10.6151
R682 B.n174 B.n65 10.6151
R683 B.n178 B.n65 10.6151
R684 B.n179 B.n178 10.6151
R685 B.n180 B.n179 10.6151
R686 B.n180 B.n63 10.6151
R687 B.n184 B.n63 10.6151
R688 B.n24 B.n20 9.36635
R689 B.n281 B.n280 9.36635
R690 B.n149 B.n148 9.36635
R691 B.n167 B.n166 9.36635
R692 B.n353 B.n0 8.11757
R693 B.n353 B.n1 8.11757
R694 B.n295 B.n24 1.24928
R695 B.n282 B.n281 1.24928
R696 B.n148 B.n75 1.24928
R697 B.n166 B.n165 1.24928
R698 VN.n7 VN.n6 161.3
R699 VN.n15 VN.n14 161.3
R700 VN.n2 VN.t6 159.186
R701 VN.n10 VN.t3 159.186
R702 VN.n1 VN.t9 132.365
R703 VN.n4 VN.t4 132.365
R704 VN.n5 VN.t7 132.365
R705 VN.n6 VN.t2 132.365
R706 VN.n9 VN.t0 132.365
R707 VN.n12 VN.t8 132.365
R708 VN.n13 VN.t5 132.365
R709 VN.n14 VN.t1 132.365
R710 VN.n13 VN.n8 80.6037
R711 VN.n12 VN.n11 80.6037
R712 VN.n5 VN.n0 80.6037
R713 VN.n4 VN.n3 80.6037
R714 VN.n4 VN.n1 48.2005
R715 VN.n5 VN.n4 48.2005
R716 VN.n6 VN.n5 48.2005
R717 VN.n12 VN.n9 48.2005
R718 VN.n13 VN.n12 48.2005
R719 VN.n14 VN.n13 48.2005
R720 VN.n11 VN.n10 45.2318
R721 VN.n3 VN.n2 45.2318
R722 VN VN.n15 35.366
R723 VN.n10 VN.n9 13.3799
R724 VN.n2 VN.n1 13.3799
R725 VN.n11 VN.n8 0.380177
R726 VN.n3 VN.n0 0.380177
R727 VN.n15 VN.n8 0.285035
R728 VN.n7 VN.n0 0.285035
R729 VN VN.n7 0.0516364
R730 VDD2.n13 VDD2.n11 756.745
R731 VDD2.n2 VDD2.n0 756.745
R732 VDD2.n14 VDD2.n13 585
R733 VDD2.n3 VDD2.n2 585
R734 VDD2.t3 VDD2.n1 417.779
R735 VDD2.t8 VDD2.n12 417.779
R736 VDD2.n10 VDD2.n9 200.052
R737 VDD2 VDD2.n21 200.048
R738 VDD2.n20 VDD2.n19 199.474
R739 VDD2.n8 VDD2.n7 199.474
R740 VDD2.n13 VDD2.t8 85.8723
R741 VDD2.n2 VDD2.t3 85.8723
R742 VDD2.n8 VDD2.n6 47.5756
R743 VDD2.n18 VDD2.n17 46.7308
R744 VDD2.n18 VDD2.n10 29.392
R745 VDD2.n21 VDD2.t9 16.8425
R746 VDD2.n21 VDD2.t6 16.8425
R747 VDD2.n19 VDD2.t4 16.8425
R748 VDD2.n19 VDD2.t1 16.8425
R749 VDD2.n9 VDD2.t2 16.8425
R750 VDD2.n9 VDD2.t7 16.8425
R751 VDD2.n7 VDD2.t0 16.8425
R752 VDD2.n7 VDD2.t5 16.8425
R753 VDD2.n14 VDD2.n12 9.84608
R754 VDD2.n3 VDD2.n1 9.84608
R755 VDD2.n17 VDD2.n16 9.45567
R756 VDD2.n6 VDD2.n5 9.45567
R757 VDD2.n16 VDD2.n15 9.3005
R758 VDD2.n5 VDD2.n4 9.3005
R759 VDD2.n17 VDD2.n11 8.14595
R760 VDD2.n6 VDD2.n0 8.14595
R761 VDD2.n15 VDD2.n14 7.3702
R762 VDD2.n4 VDD2.n3 7.3702
R763 VDD2.n15 VDD2.n11 5.81868
R764 VDD2.n4 VDD2.n0 5.81868
R765 VDD2.n16 VDD2.n12 3.32369
R766 VDD2.n5 VDD2.n1 3.32369
R767 VDD2.n20 VDD2.n18 0.845328
R768 VDD2 VDD2.n20 0.269897
R769 VDD2.n10 VDD2.n8 0.156361
C0 VDD2 B 0.9923f
C1 VDD2 VDD1 0.939278f
C2 VP w_n2146_n1354# 4.03651f
C3 VTAIL VP 1.73367f
C4 VDD1 B 0.949778f
C5 VDD2 w_n2146_n1354# 1.31161f
C6 VDD2 VTAIL 4.46583f
C7 VDD1 w_n2146_n1354# 1.27032f
C8 w_n2146_n1354# B 4.43636f
C9 VTAIL VDD1 4.42641f
C10 VTAIL B 0.881091f
C11 VP VN 3.6631f
C12 VTAIL w_n2146_n1354# 1.40149f
C13 VDD2 VN 1.38961f
C14 VDD1 VN 0.155574f
C15 VN B 0.662354f
C16 VN w_n2146_n1354# 3.76795f
C17 VTAIL VN 1.71948f
C18 VDD2 VP 0.341144f
C19 VP VDD1 1.57307f
C20 VP B 1.11053f
C21 VDD2 VSUBS 0.767928f
C22 VDD1 VSUBS 0.794693f
C23 VTAIL VSUBS 0.301962f
C24 VN VSUBS 3.69054f
C25 VP VSUBS 1.266203f
C26 B VSUBS 1.992952f
C27 w_n2146_n1354# VSUBS 37.1086f
C28 VDD2.n0 VSUBS 0.020993f
C29 VDD2.n1 VSUBS 0.054221f
C30 VDD2.t3 VSUBS 0.054343f
C31 VDD2.n2 VSUBS 0.052681f
C32 VDD2.n3 VSUBS 0.015825f
C33 VDD2.n4 VSUBS 0.010266f
C34 VDD2.n5 VSUBS 0.126877f
C35 VDD2.n6 VSUBS 0.044216f
C36 VDD2.t0 VSUBS 0.029137f
C37 VDD2.t5 VSUBS 0.029137f
C38 VDD2.n7 VSUBS 0.12019f
C39 VDD2.n8 VSUBS 0.355718f
C40 VDD2.t2 VSUBS 0.029137f
C41 VDD2.t7 VSUBS 0.029137f
C42 VDD2.n9 VSUBS 0.121062f
C43 VDD2.n10 VSUBS 1.03543f
C44 VDD2.n11 VSUBS 0.020993f
C45 VDD2.n12 VSUBS 0.054221f
C46 VDD2.t8 VSUBS 0.054343f
C47 VDD2.n13 VSUBS 0.052681f
C48 VDD2.n14 VSUBS 0.015825f
C49 VDD2.n15 VSUBS 0.010266f
C50 VDD2.n16 VSUBS 0.126877f
C51 VDD2.n17 VSUBS 0.042669f
C52 VDD2.n18 VSUBS 1.00976f
C53 VDD2.t4 VSUBS 0.029137f
C54 VDD2.t1 VSUBS 0.029137f
C55 VDD2.n19 VSUBS 0.12019f
C56 VDD2.n20 VSUBS 0.274261f
C57 VDD2.t9 VSUBS 0.029137f
C58 VDD2.t6 VSUBS 0.029137f
C59 VDD2.n21 VSUBS 0.121056f
C60 VN.n0 VSUBS 0.086128f
C61 VN.t9 VSUBS 0.201889f
C62 VN.n1 VSUBS 0.156281f
C63 VN.t6 VSUBS 0.22627f
C64 VN.n2 VSUBS 0.121774f
C65 VN.n3 VSUBS 0.275112f
C66 VN.t4 VSUBS 0.201889f
C67 VN.n4 VSUBS 0.156281f
C68 VN.t7 VSUBS 0.201889f
C69 VN.n5 VSUBS 0.156281f
C70 VN.t2 VSUBS 0.201889f
C71 VN.n6 VSUBS 0.144547f
C72 VN.n7 VSUBS 0.057363f
C73 VN.n8 VSUBS 0.086128f
C74 VN.t0 VSUBS 0.201889f
C75 VN.n9 VSUBS 0.156281f
C76 VN.t8 VSUBS 0.201889f
C77 VN.t3 VSUBS 0.22627f
C78 VN.n10 VSUBS 0.121774f
C79 VN.n11 VSUBS 0.275112f
C80 VN.n12 VSUBS 0.156281f
C81 VN.t5 VSUBS 0.201889f
C82 VN.n13 VSUBS 0.156281f
C83 VN.t1 VSUBS 0.201889f
C84 VN.n14 VSUBS 0.144547f
C85 VN.n15 VSUBS 1.59123f
C86 B.n0 VSUBS 0.007559f
C87 B.n1 VSUBS 0.007559f
C88 B.n2 VSUBS 0.01118f
C89 B.n3 VSUBS 0.008567f
C90 B.n4 VSUBS 0.008567f
C91 B.n5 VSUBS 0.008567f
C92 B.n6 VSUBS 0.008567f
C93 B.n7 VSUBS 0.008567f
C94 B.n8 VSUBS 0.008567f
C95 B.n9 VSUBS 0.008567f
C96 B.n10 VSUBS 0.008567f
C97 B.n11 VSUBS 0.008567f
C98 B.n12 VSUBS 0.008567f
C99 B.n13 VSUBS 0.008567f
C100 B.n14 VSUBS 0.017997f
C101 B.n15 VSUBS 0.008567f
C102 B.n16 VSUBS 0.008567f
C103 B.n17 VSUBS 0.008567f
C104 B.n18 VSUBS 0.008567f
C105 B.n19 VSUBS 0.008567f
C106 B.n20 VSUBS 0.008063f
C107 B.n21 VSUBS 0.008567f
C108 B.t1 VSUBS 0.040164f
C109 B.t2 VSUBS 0.044353f
C110 B.t0 VSUBS 0.072995f
C111 B.n22 VSUBS 0.075164f
C112 B.n23 VSUBS 0.07084f
C113 B.n24 VSUBS 0.019849f
C114 B.n25 VSUBS 0.008567f
C115 B.n26 VSUBS 0.008567f
C116 B.n27 VSUBS 0.008567f
C117 B.n28 VSUBS 0.008567f
C118 B.t7 VSUBS 0.040164f
C119 B.t8 VSUBS 0.044353f
C120 B.t6 VSUBS 0.072995f
C121 B.n29 VSUBS 0.075164f
C122 B.n30 VSUBS 0.07084f
C123 B.n31 VSUBS 0.008567f
C124 B.n32 VSUBS 0.008567f
C125 B.n33 VSUBS 0.008567f
C126 B.n34 VSUBS 0.008567f
C127 B.n35 VSUBS 0.008567f
C128 B.n36 VSUBS 0.019295f
C129 B.n37 VSUBS 0.008567f
C130 B.n38 VSUBS 0.008567f
C131 B.n39 VSUBS 0.008567f
C132 B.n40 VSUBS 0.008567f
C133 B.n41 VSUBS 0.008567f
C134 B.n42 VSUBS 0.008567f
C135 B.n43 VSUBS 0.008567f
C136 B.n44 VSUBS 0.008567f
C137 B.n45 VSUBS 0.008567f
C138 B.n46 VSUBS 0.008567f
C139 B.n47 VSUBS 0.008567f
C140 B.n48 VSUBS 0.008567f
C141 B.n49 VSUBS 0.008567f
C142 B.n50 VSUBS 0.008567f
C143 B.n51 VSUBS 0.008567f
C144 B.n52 VSUBS 0.008567f
C145 B.n53 VSUBS 0.008567f
C146 B.n54 VSUBS 0.008567f
C147 B.n55 VSUBS 0.008567f
C148 B.n56 VSUBS 0.008567f
C149 B.n57 VSUBS 0.008567f
C150 B.n58 VSUBS 0.008567f
C151 B.n59 VSUBS 0.008567f
C152 B.n60 VSUBS 0.008567f
C153 B.n61 VSUBS 0.008567f
C154 B.n62 VSUBS 0.017997f
C155 B.n63 VSUBS 0.008567f
C156 B.n64 VSUBS 0.008567f
C157 B.n65 VSUBS 0.008567f
C158 B.n66 VSUBS 0.008567f
C159 B.n67 VSUBS 0.008567f
C160 B.n68 VSUBS 0.008567f
C161 B.t11 VSUBS 0.040164f
C162 B.t10 VSUBS 0.044353f
C163 B.t9 VSUBS 0.072995f
C164 B.n69 VSUBS 0.075164f
C165 B.n70 VSUBS 0.07084f
C166 B.n71 VSUBS 0.008567f
C167 B.n72 VSUBS 0.008567f
C168 B.n73 VSUBS 0.008567f
C169 B.n74 VSUBS 0.008567f
C170 B.n75 VSUBS 0.004787f
C171 B.n76 VSUBS 0.008567f
C172 B.n77 VSUBS 0.008567f
C173 B.n78 VSUBS 0.008567f
C174 B.n79 VSUBS 0.008567f
C175 B.n80 VSUBS 0.008567f
C176 B.n81 VSUBS 0.019295f
C177 B.n82 VSUBS 0.008567f
C178 B.n83 VSUBS 0.008567f
C179 B.n84 VSUBS 0.008567f
C180 B.n85 VSUBS 0.008567f
C181 B.n86 VSUBS 0.008567f
C182 B.n87 VSUBS 0.008567f
C183 B.n88 VSUBS 0.008567f
C184 B.n89 VSUBS 0.008567f
C185 B.n90 VSUBS 0.008567f
C186 B.n91 VSUBS 0.008567f
C187 B.n92 VSUBS 0.008567f
C188 B.n93 VSUBS 0.008567f
C189 B.n94 VSUBS 0.008567f
C190 B.n95 VSUBS 0.008567f
C191 B.n96 VSUBS 0.008567f
C192 B.n97 VSUBS 0.008567f
C193 B.n98 VSUBS 0.008567f
C194 B.n99 VSUBS 0.008567f
C195 B.n100 VSUBS 0.008567f
C196 B.n101 VSUBS 0.008567f
C197 B.n102 VSUBS 0.008567f
C198 B.n103 VSUBS 0.008567f
C199 B.n104 VSUBS 0.008567f
C200 B.n105 VSUBS 0.008567f
C201 B.n106 VSUBS 0.008567f
C202 B.n107 VSUBS 0.008567f
C203 B.n108 VSUBS 0.008567f
C204 B.n109 VSUBS 0.008567f
C205 B.n110 VSUBS 0.008567f
C206 B.n111 VSUBS 0.008567f
C207 B.n112 VSUBS 0.008567f
C208 B.n113 VSUBS 0.008567f
C209 B.n114 VSUBS 0.008567f
C210 B.n115 VSUBS 0.008567f
C211 B.n116 VSUBS 0.008567f
C212 B.n117 VSUBS 0.008567f
C213 B.n118 VSUBS 0.008567f
C214 B.n119 VSUBS 0.008567f
C215 B.n120 VSUBS 0.008567f
C216 B.n121 VSUBS 0.008567f
C217 B.n122 VSUBS 0.008567f
C218 B.n123 VSUBS 0.008567f
C219 B.n124 VSUBS 0.008567f
C220 B.n125 VSUBS 0.008567f
C221 B.n126 VSUBS 0.008567f
C222 B.n127 VSUBS 0.008567f
C223 B.n128 VSUBS 0.017997f
C224 B.n129 VSUBS 0.017997f
C225 B.n130 VSUBS 0.019295f
C226 B.n131 VSUBS 0.008567f
C227 B.n132 VSUBS 0.008567f
C228 B.n133 VSUBS 0.008567f
C229 B.n134 VSUBS 0.008567f
C230 B.n135 VSUBS 0.008567f
C231 B.n136 VSUBS 0.008567f
C232 B.n137 VSUBS 0.008567f
C233 B.n138 VSUBS 0.008567f
C234 B.n139 VSUBS 0.008567f
C235 B.n140 VSUBS 0.008567f
C236 B.n141 VSUBS 0.008567f
C237 B.n142 VSUBS 0.008567f
C238 B.n143 VSUBS 0.008567f
C239 B.n144 VSUBS 0.008567f
C240 B.n145 VSUBS 0.008567f
C241 B.t5 VSUBS 0.040164f
C242 B.t4 VSUBS 0.044353f
C243 B.t3 VSUBS 0.072995f
C244 B.n146 VSUBS 0.075164f
C245 B.n147 VSUBS 0.07084f
C246 B.n148 VSUBS 0.019849f
C247 B.n149 VSUBS 0.008063f
C248 B.n150 VSUBS 0.008567f
C249 B.n151 VSUBS 0.008567f
C250 B.n152 VSUBS 0.008567f
C251 B.n153 VSUBS 0.008567f
C252 B.n154 VSUBS 0.008567f
C253 B.n155 VSUBS 0.008567f
C254 B.n156 VSUBS 0.008567f
C255 B.n157 VSUBS 0.008567f
C256 B.n158 VSUBS 0.008567f
C257 B.n159 VSUBS 0.008567f
C258 B.n160 VSUBS 0.008567f
C259 B.n161 VSUBS 0.008567f
C260 B.n162 VSUBS 0.008567f
C261 B.n163 VSUBS 0.008567f
C262 B.n164 VSUBS 0.008567f
C263 B.n165 VSUBS 0.004787f
C264 B.n166 VSUBS 0.019849f
C265 B.n167 VSUBS 0.008063f
C266 B.n168 VSUBS 0.008567f
C267 B.n169 VSUBS 0.008567f
C268 B.n170 VSUBS 0.008567f
C269 B.n171 VSUBS 0.008567f
C270 B.n172 VSUBS 0.008567f
C271 B.n173 VSUBS 0.008567f
C272 B.n174 VSUBS 0.008567f
C273 B.n175 VSUBS 0.008567f
C274 B.n176 VSUBS 0.008567f
C275 B.n177 VSUBS 0.008567f
C276 B.n178 VSUBS 0.008567f
C277 B.n179 VSUBS 0.008567f
C278 B.n180 VSUBS 0.008567f
C279 B.n181 VSUBS 0.008567f
C280 B.n182 VSUBS 0.008567f
C281 B.n183 VSUBS 0.019295f
C282 B.n184 VSUBS 0.018162f
C283 B.n185 VSUBS 0.019129f
C284 B.n186 VSUBS 0.008567f
C285 B.n187 VSUBS 0.008567f
C286 B.n188 VSUBS 0.008567f
C287 B.n189 VSUBS 0.008567f
C288 B.n190 VSUBS 0.008567f
C289 B.n191 VSUBS 0.008567f
C290 B.n192 VSUBS 0.008567f
C291 B.n193 VSUBS 0.008567f
C292 B.n194 VSUBS 0.008567f
C293 B.n195 VSUBS 0.008567f
C294 B.n196 VSUBS 0.008567f
C295 B.n197 VSUBS 0.008567f
C296 B.n198 VSUBS 0.008567f
C297 B.n199 VSUBS 0.008567f
C298 B.n200 VSUBS 0.008567f
C299 B.n201 VSUBS 0.008567f
C300 B.n202 VSUBS 0.008567f
C301 B.n203 VSUBS 0.008567f
C302 B.n204 VSUBS 0.008567f
C303 B.n205 VSUBS 0.008567f
C304 B.n206 VSUBS 0.008567f
C305 B.n207 VSUBS 0.008567f
C306 B.n208 VSUBS 0.008567f
C307 B.n209 VSUBS 0.008567f
C308 B.n210 VSUBS 0.008567f
C309 B.n211 VSUBS 0.008567f
C310 B.n212 VSUBS 0.008567f
C311 B.n213 VSUBS 0.008567f
C312 B.n214 VSUBS 0.008567f
C313 B.n215 VSUBS 0.008567f
C314 B.n216 VSUBS 0.008567f
C315 B.n217 VSUBS 0.008567f
C316 B.n218 VSUBS 0.008567f
C317 B.n219 VSUBS 0.008567f
C318 B.n220 VSUBS 0.008567f
C319 B.n221 VSUBS 0.008567f
C320 B.n222 VSUBS 0.008567f
C321 B.n223 VSUBS 0.008567f
C322 B.n224 VSUBS 0.008567f
C323 B.n225 VSUBS 0.008567f
C324 B.n226 VSUBS 0.008567f
C325 B.n227 VSUBS 0.008567f
C326 B.n228 VSUBS 0.008567f
C327 B.n229 VSUBS 0.008567f
C328 B.n230 VSUBS 0.008567f
C329 B.n231 VSUBS 0.008567f
C330 B.n232 VSUBS 0.008567f
C331 B.n233 VSUBS 0.008567f
C332 B.n234 VSUBS 0.008567f
C333 B.n235 VSUBS 0.008567f
C334 B.n236 VSUBS 0.008567f
C335 B.n237 VSUBS 0.008567f
C336 B.n238 VSUBS 0.008567f
C337 B.n239 VSUBS 0.008567f
C338 B.n240 VSUBS 0.008567f
C339 B.n241 VSUBS 0.008567f
C340 B.n242 VSUBS 0.008567f
C341 B.n243 VSUBS 0.008567f
C342 B.n244 VSUBS 0.008567f
C343 B.n245 VSUBS 0.008567f
C344 B.n246 VSUBS 0.008567f
C345 B.n247 VSUBS 0.008567f
C346 B.n248 VSUBS 0.008567f
C347 B.n249 VSUBS 0.008567f
C348 B.n250 VSUBS 0.008567f
C349 B.n251 VSUBS 0.008567f
C350 B.n252 VSUBS 0.008567f
C351 B.n253 VSUBS 0.008567f
C352 B.n254 VSUBS 0.008567f
C353 B.n255 VSUBS 0.008567f
C354 B.n256 VSUBS 0.008567f
C355 B.n257 VSUBS 0.008567f
C356 B.n258 VSUBS 0.008567f
C357 B.n259 VSUBS 0.008567f
C358 B.n260 VSUBS 0.008567f
C359 B.n261 VSUBS 0.017997f
C360 B.n262 VSUBS 0.017997f
C361 B.n263 VSUBS 0.019295f
C362 B.n264 VSUBS 0.008567f
C363 B.n265 VSUBS 0.008567f
C364 B.n266 VSUBS 0.008567f
C365 B.n267 VSUBS 0.008567f
C366 B.n268 VSUBS 0.008567f
C367 B.n269 VSUBS 0.008567f
C368 B.n270 VSUBS 0.008567f
C369 B.n271 VSUBS 0.008567f
C370 B.n272 VSUBS 0.008567f
C371 B.n273 VSUBS 0.008567f
C372 B.n274 VSUBS 0.008567f
C373 B.n275 VSUBS 0.008567f
C374 B.n276 VSUBS 0.008567f
C375 B.n277 VSUBS 0.008567f
C376 B.n278 VSUBS 0.008567f
C377 B.n279 VSUBS 0.008567f
C378 B.n280 VSUBS 0.008063f
C379 B.n281 VSUBS 0.019849f
C380 B.n282 VSUBS 0.004787f
C381 B.n283 VSUBS 0.008567f
C382 B.n284 VSUBS 0.008567f
C383 B.n285 VSUBS 0.008567f
C384 B.n286 VSUBS 0.008567f
C385 B.n287 VSUBS 0.008567f
C386 B.n288 VSUBS 0.008567f
C387 B.n289 VSUBS 0.008567f
C388 B.n290 VSUBS 0.008567f
C389 B.n291 VSUBS 0.008567f
C390 B.n292 VSUBS 0.008567f
C391 B.n293 VSUBS 0.008567f
C392 B.n294 VSUBS 0.008567f
C393 B.n295 VSUBS 0.004787f
C394 B.n296 VSUBS 0.008567f
C395 B.n297 VSUBS 0.008567f
C396 B.n298 VSUBS 0.008567f
C397 B.n299 VSUBS 0.008567f
C398 B.n300 VSUBS 0.008567f
C399 B.n301 VSUBS 0.008567f
C400 B.n302 VSUBS 0.008567f
C401 B.n303 VSUBS 0.008567f
C402 B.n304 VSUBS 0.008567f
C403 B.n305 VSUBS 0.008567f
C404 B.n306 VSUBS 0.008567f
C405 B.n307 VSUBS 0.008567f
C406 B.n308 VSUBS 0.008567f
C407 B.n309 VSUBS 0.008567f
C408 B.n310 VSUBS 0.008567f
C409 B.n311 VSUBS 0.008567f
C410 B.n312 VSUBS 0.008567f
C411 B.n313 VSUBS 0.019295f
C412 B.n314 VSUBS 0.019295f
C413 B.n315 VSUBS 0.017997f
C414 B.n316 VSUBS 0.008567f
C415 B.n317 VSUBS 0.008567f
C416 B.n318 VSUBS 0.008567f
C417 B.n319 VSUBS 0.008567f
C418 B.n320 VSUBS 0.008567f
C419 B.n321 VSUBS 0.008567f
C420 B.n322 VSUBS 0.008567f
C421 B.n323 VSUBS 0.008567f
C422 B.n324 VSUBS 0.008567f
C423 B.n325 VSUBS 0.008567f
C424 B.n326 VSUBS 0.008567f
C425 B.n327 VSUBS 0.008567f
C426 B.n328 VSUBS 0.008567f
C427 B.n329 VSUBS 0.008567f
C428 B.n330 VSUBS 0.008567f
C429 B.n331 VSUBS 0.008567f
C430 B.n332 VSUBS 0.008567f
C431 B.n333 VSUBS 0.008567f
C432 B.n334 VSUBS 0.008567f
C433 B.n335 VSUBS 0.008567f
C434 B.n336 VSUBS 0.008567f
C435 B.n337 VSUBS 0.008567f
C436 B.n338 VSUBS 0.008567f
C437 B.n339 VSUBS 0.008567f
C438 B.n340 VSUBS 0.008567f
C439 B.n341 VSUBS 0.008567f
C440 B.n342 VSUBS 0.008567f
C441 B.n343 VSUBS 0.008567f
C442 B.n344 VSUBS 0.008567f
C443 B.n345 VSUBS 0.008567f
C444 B.n346 VSUBS 0.008567f
C445 B.n347 VSUBS 0.008567f
C446 B.n348 VSUBS 0.008567f
C447 B.n349 VSUBS 0.008567f
C448 B.n350 VSUBS 0.008567f
C449 B.n351 VSUBS 0.01118f
C450 B.n352 VSUBS 0.011909f
C451 B.n353 VSUBS 0.023682f
C452 VDD1.n0 VSUBS 0.02021f
C453 VDD1.n1 VSUBS 0.052198f
C454 VDD1.t7 VSUBS 0.052315f
C455 VDD1.n2 VSUBS 0.050715f
C456 VDD1.n3 VSUBS 0.015235f
C457 VDD1.n4 VSUBS 0.009883f
C458 VDD1.n5 VSUBS 0.122142f
C459 VDD1.n6 VSUBS 0.042566f
C460 VDD1.t0 VSUBS 0.02805f
C461 VDD1.t3 VSUBS 0.02805f
C462 VDD1.n7 VSUBS 0.115705f
C463 VDD1.n8 VSUBS 0.346436f
C464 VDD1.n9 VSUBS 0.02021f
C465 VDD1.n10 VSUBS 0.052198f
C466 VDD1.t6 VSUBS 0.052315f
C467 VDD1.n11 VSUBS 0.050715f
C468 VDD1.n12 VSUBS 0.015235f
C469 VDD1.n13 VSUBS 0.009883f
C470 VDD1.n14 VSUBS 0.122142f
C471 VDD1.n15 VSUBS 0.042566f
C472 VDD1.t8 VSUBS 0.02805f
C473 VDD1.t4 VSUBS 0.02805f
C474 VDD1.n16 VSUBS 0.115705f
C475 VDD1.n17 VSUBS 0.342444f
C476 VDD1.t1 VSUBS 0.02805f
C477 VDD1.t2 VSUBS 0.02805f
C478 VDD1.n18 VSUBS 0.116544f
C479 VDD1.n19 VSUBS 1.04908f
C480 VDD1.t5 VSUBS 0.02805f
C481 VDD1.t9 VSUBS 0.02805f
C482 VDD1.n20 VSUBS 0.115705f
C483 VDD1.n21 VSUBS 1.19338f
C484 VTAIL.t2 VSUBS 0.036045f
C485 VTAIL.t17 VSUBS 0.036045f
C486 VTAIL.n0 VSUBS 0.12588f
C487 VTAIL.n1 VSUBS 0.365742f
C488 VTAIL.n2 VSUBS 0.02597f
C489 VTAIL.n3 VSUBS 0.067075f
C490 VTAIL.t7 VSUBS 0.067226f
C491 VTAIL.n4 VSUBS 0.06517f
C492 VTAIL.n5 VSUBS 0.019577f
C493 VTAIL.n6 VSUBS 0.0127f
C494 VTAIL.n7 VSUBS 0.156957f
C495 VTAIL.n8 VSUBS 0.036435f
C496 VTAIL.n9 VSUBS 0.150469f
C497 VTAIL.t13 VSUBS 0.036045f
C498 VTAIL.t11 VSUBS 0.036045f
C499 VTAIL.n10 VSUBS 0.12588f
C500 VTAIL.n11 VSUBS 0.373784f
C501 VTAIL.t16 VSUBS 0.036045f
C502 VTAIL.t9 VSUBS 0.036045f
C503 VTAIL.n12 VSUBS 0.12588f
C504 VTAIL.n13 VSUBS 0.885865f
C505 VTAIL.t19 VSUBS 0.036045f
C506 VTAIL.t1 VSUBS 0.036045f
C507 VTAIL.n14 VSUBS 0.12588f
C508 VTAIL.n15 VSUBS 0.885864f
C509 VTAIL.t0 VSUBS 0.036045f
C510 VTAIL.t18 VSUBS 0.036045f
C511 VTAIL.n16 VSUBS 0.12588f
C512 VTAIL.n17 VSUBS 0.373784f
C513 VTAIL.n18 VSUBS 0.02597f
C514 VTAIL.n19 VSUBS 0.067075f
C515 VTAIL.t3 VSUBS 0.067226f
C516 VTAIL.n20 VSUBS 0.06517f
C517 VTAIL.n21 VSUBS 0.019577f
C518 VTAIL.n22 VSUBS 0.0127f
C519 VTAIL.n23 VSUBS 0.156957f
C520 VTAIL.n24 VSUBS 0.036435f
C521 VTAIL.n25 VSUBS 0.150469f
C522 VTAIL.t14 VSUBS 0.036045f
C523 VTAIL.t8 VSUBS 0.036045f
C524 VTAIL.n26 VSUBS 0.12588f
C525 VTAIL.n27 VSUBS 0.377394f
C526 VTAIL.t10 VSUBS 0.036045f
C527 VTAIL.t15 VSUBS 0.036045f
C528 VTAIL.n28 VSUBS 0.12588f
C529 VTAIL.n29 VSUBS 0.373784f
C530 VTAIL.n30 VSUBS 0.02597f
C531 VTAIL.n31 VSUBS 0.067075f
C532 VTAIL.t12 VSUBS 0.067226f
C533 VTAIL.n32 VSUBS 0.06517f
C534 VTAIL.n33 VSUBS 0.019577f
C535 VTAIL.n34 VSUBS 0.0127f
C536 VTAIL.n35 VSUBS 0.156957f
C537 VTAIL.n36 VSUBS 0.036435f
C538 VTAIL.n37 VSUBS 0.594602f
C539 VTAIL.n38 VSUBS 0.02597f
C540 VTAIL.n39 VSUBS 0.067075f
C541 VTAIL.t4 VSUBS 0.067226f
C542 VTAIL.n40 VSUBS 0.06517f
C543 VTAIL.n41 VSUBS 0.019577f
C544 VTAIL.n42 VSUBS 0.0127f
C545 VTAIL.n43 VSUBS 0.156957f
C546 VTAIL.n44 VSUBS 0.036435f
C547 VTAIL.n45 VSUBS 0.594602f
C548 VTAIL.t6 VSUBS 0.036045f
C549 VTAIL.t5 VSUBS 0.036045f
C550 VTAIL.n46 VSUBS 0.12588f
C551 VTAIL.n47 VSUBS 0.3211f
C552 VP.n0 VSUBS 0.08929f
C553 VP.t1 VSUBS 0.209301f
C554 VP.n1 VSUBS 0.162019f
C555 VP.n2 VSUBS 0.08929f
C556 VP.t0 VSUBS 0.209301f
C557 VP.t4 VSUBS 0.209301f
C558 VP.t6 VSUBS 0.209301f
C559 VP.n3 VSUBS 0.285212f
C560 VP.t9 VSUBS 0.209301f
C561 VP.t2 VSUBS 0.234577f
C562 VP.n4 VSUBS 0.126245f
C563 VP.n5 VSUBS 0.162019f
C564 VP.n6 VSUBS 0.162019f
C565 VP.n7 VSUBS 0.162019f
C566 VP.n8 VSUBS 0.149854f
C567 VP.n9 VSUBS 1.61402f
C568 VP.t3 VSUBS 0.209301f
C569 VP.n10 VSUBS 0.149854f
C570 VP.n11 VSUBS 1.6691f
C571 VP.n12 VSUBS 0.08929f
C572 VP.n13 VSUBS 0.107216f
C573 VP.t5 VSUBS 0.209301f
C574 VP.n14 VSUBS 0.162019f
C575 VP.t8 VSUBS 0.209301f
C576 VP.n15 VSUBS 0.162019f
C577 VP.t7 VSUBS 0.209301f
C578 VP.n16 VSUBS 0.149854f
C579 VP.n17 VSUBS 0.059469f
.ends

