* NGSPICE file created from diff_pair_sample_0675.ext - technology: sky130A

.subckt diff_pair_sample_0675 VTAIL VN VP B VDD2 VDD1
X0 B.t15 B.t13 B.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=0 ps=0 w=9.17 l=1.31
X1 VDD1.t1 VP.t0 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=3.5763 ps=19.12 w=9.17 l=1.31
X2 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=0 ps=0 w=9.17 l=1.31
X3 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=0 ps=0 w=9.17 l=1.31
X4 VDD2.t1 VN.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=3.5763 ps=19.12 w=9.17 l=1.31
X5 VDD2.t0 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=3.5763 ps=19.12 w=9.17 l=1.31
X6 VDD1.t0 VP.t1 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=3.5763 ps=19.12 w=9.17 l=1.31
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=3.5763 pd=19.12 as=0 ps=0 w=9.17 l=1.31
R0 B.n532 B.n531 585
R1 B.n227 B.n72 585
R2 B.n226 B.n225 585
R3 B.n224 B.n223 585
R4 B.n222 B.n221 585
R5 B.n220 B.n219 585
R6 B.n218 B.n217 585
R7 B.n216 B.n215 585
R8 B.n214 B.n213 585
R9 B.n212 B.n211 585
R10 B.n210 B.n209 585
R11 B.n208 B.n207 585
R12 B.n206 B.n205 585
R13 B.n204 B.n203 585
R14 B.n202 B.n201 585
R15 B.n200 B.n199 585
R16 B.n198 B.n197 585
R17 B.n196 B.n195 585
R18 B.n194 B.n193 585
R19 B.n192 B.n191 585
R20 B.n190 B.n189 585
R21 B.n188 B.n187 585
R22 B.n186 B.n185 585
R23 B.n184 B.n183 585
R24 B.n182 B.n181 585
R25 B.n180 B.n179 585
R26 B.n178 B.n177 585
R27 B.n176 B.n175 585
R28 B.n174 B.n173 585
R29 B.n172 B.n171 585
R30 B.n170 B.n169 585
R31 B.n168 B.n167 585
R32 B.n166 B.n165 585
R33 B.n163 B.n162 585
R34 B.n161 B.n160 585
R35 B.n159 B.n158 585
R36 B.n157 B.n156 585
R37 B.n155 B.n154 585
R38 B.n153 B.n152 585
R39 B.n151 B.n150 585
R40 B.n149 B.n148 585
R41 B.n147 B.n146 585
R42 B.n145 B.n144 585
R43 B.n142 B.n141 585
R44 B.n140 B.n139 585
R45 B.n138 B.n137 585
R46 B.n136 B.n135 585
R47 B.n134 B.n133 585
R48 B.n132 B.n131 585
R49 B.n130 B.n129 585
R50 B.n128 B.n127 585
R51 B.n126 B.n125 585
R52 B.n124 B.n123 585
R53 B.n122 B.n121 585
R54 B.n120 B.n119 585
R55 B.n118 B.n117 585
R56 B.n116 B.n115 585
R57 B.n114 B.n113 585
R58 B.n112 B.n111 585
R59 B.n110 B.n109 585
R60 B.n108 B.n107 585
R61 B.n106 B.n105 585
R62 B.n104 B.n103 585
R63 B.n102 B.n101 585
R64 B.n100 B.n99 585
R65 B.n98 B.n97 585
R66 B.n96 B.n95 585
R67 B.n94 B.n93 585
R68 B.n92 B.n91 585
R69 B.n90 B.n89 585
R70 B.n88 B.n87 585
R71 B.n86 B.n85 585
R72 B.n84 B.n83 585
R73 B.n82 B.n81 585
R74 B.n80 B.n79 585
R75 B.n78 B.n77 585
R76 B.n530 B.n34 585
R77 B.n535 B.n34 585
R78 B.n529 B.n33 585
R79 B.n536 B.n33 585
R80 B.n528 B.n527 585
R81 B.n527 B.n29 585
R82 B.n526 B.n28 585
R83 B.n542 B.n28 585
R84 B.n525 B.n27 585
R85 B.n543 B.n27 585
R86 B.n524 B.n26 585
R87 B.n544 B.n26 585
R88 B.n523 B.n522 585
R89 B.n522 B.n22 585
R90 B.n521 B.n21 585
R91 B.n550 B.n21 585
R92 B.n520 B.n20 585
R93 B.n551 B.n20 585
R94 B.n519 B.n19 585
R95 B.n552 B.n19 585
R96 B.n518 B.n517 585
R97 B.n517 B.n15 585
R98 B.n516 B.n14 585
R99 B.n558 B.n14 585
R100 B.n515 B.n13 585
R101 B.n559 B.n13 585
R102 B.n514 B.n12 585
R103 B.n560 B.n12 585
R104 B.n513 B.n512 585
R105 B.n512 B.n511 585
R106 B.n510 B.n509 585
R107 B.n510 B.n8 585
R108 B.n508 B.n7 585
R109 B.n567 B.n7 585
R110 B.n507 B.n6 585
R111 B.n568 B.n6 585
R112 B.n506 B.n5 585
R113 B.n569 B.n5 585
R114 B.n505 B.n504 585
R115 B.n504 B.n4 585
R116 B.n503 B.n228 585
R117 B.n503 B.n502 585
R118 B.n493 B.n229 585
R119 B.n230 B.n229 585
R120 B.n495 B.n494 585
R121 B.n496 B.n495 585
R122 B.n492 B.n235 585
R123 B.n235 B.n234 585
R124 B.n491 B.n490 585
R125 B.n490 B.n489 585
R126 B.n237 B.n236 585
R127 B.n238 B.n237 585
R128 B.n482 B.n481 585
R129 B.n483 B.n482 585
R130 B.n480 B.n243 585
R131 B.n243 B.n242 585
R132 B.n479 B.n478 585
R133 B.n478 B.n477 585
R134 B.n245 B.n244 585
R135 B.n246 B.n245 585
R136 B.n470 B.n469 585
R137 B.n471 B.n470 585
R138 B.n468 B.n251 585
R139 B.n251 B.n250 585
R140 B.n467 B.n466 585
R141 B.n466 B.n465 585
R142 B.n253 B.n252 585
R143 B.n254 B.n253 585
R144 B.n458 B.n457 585
R145 B.n459 B.n458 585
R146 B.n456 B.n259 585
R147 B.n259 B.n258 585
R148 B.n451 B.n450 585
R149 B.n449 B.n299 585
R150 B.n448 B.n298 585
R151 B.n453 B.n298 585
R152 B.n447 B.n446 585
R153 B.n445 B.n444 585
R154 B.n443 B.n442 585
R155 B.n441 B.n440 585
R156 B.n439 B.n438 585
R157 B.n437 B.n436 585
R158 B.n435 B.n434 585
R159 B.n433 B.n432 585
R160 B.n431 B.n430 585
R161 B.n429 B.n428 585
R162 B.n427 B.n426 585
R163 B.n425 B.n424 585
R164 B.n423 B.n422 585
R165 B.n421 B.n420 585
R166 B.n419 B.n418 585
R167 B.n417 B.n416 585
R168 B.n415 B.n414 585
R169 B.n413 B.n412 585
R170 B.n411 B.n410 585
R171 B.n409 B.n408 585
R172 B.n407 B.n406 585
R173 B.n405 B.n404 585
R174 B.n403 B.n402 585
R175 B.n401 B.n400 585
R176 B.n399 B.n398 585
R177 B.n397 B.n396 585
R178 B.n395 B.n394 585
R179 B.n393 B.n392 585
R180 B.n391 B.n390 585
R181 B.n389 B.n388 585
R182 B.n387 B.n386 585
R183 B.n385 B.n384 585
R184 B.n383 B.n382 585
R185 B.n381 B.n380 585
R186 B.n379 B.n378 585
R187 B.n377 B.n376 585
R188 B.n375 B.n374 585
R189 B.n373 B.n372 585
R190 B.n371 B.n370 585
R191 B.n369 B.n368 585
R192 B.n367 B.n366 585
R193 B.n365 B.n364 585
R194 B.n363 B.n362 585
R195 B.n361 B.n360 585
R196 B.n359 B.n358 585
R197 B.n357 B.n356 585
R198 B.n355 B.n354 585
R199 B.n353 B.n352 585
R200 B.n351 B.n350 585
R201 B.n349 B.n348 585
R202 B.n347 B.n346 585
R203 B.n345 B.n344 585
R204 B.n343 B.n342 585
R205 B.n341 B.n340 585
R206 B.n339 B.n338 585
R207 B.n337 B.n336 585
R208 B.n335 B.n334 585
R209 B.n333 B.n332 585
R210 B.n331 B.n330 585
R211 B.n329 B.n328 585
R212 B.n327 B.n326 585
R213 B.n325 B.n324 585
R214 B.n323 B.n322 585
R215 B.n321 B.n320 585
R216 B.n319 B.n318 585
R217 B.n317 B.n316 585
R218 B.n315 B.n314 585
R219 B.n313 B.n312 585
R220 B.n311 B.n310 585
R221 B.n309 B.n308 585
R222 B.n307 B.n306 585
R223 B.n261 B.n260 585
R224 B.n455 B.n454 585
R225 B.n454 B.n453 585
R226 B.n257 B.n256 585
R227 B.n258 B.n257 585
R228 B.n461 B.n460 585
R229 B.n460 B.n459 585
R230 B.n462 B.n255 585
R231 B.n255 B.n254 585
R232 B.n464 B.n463 585
R233 B.n465 B.n464 585
R234 B.n249 B.n248 585
R235 B.n250 B.n249 585
R236 B.n473 B.n472 585
R237 B.n472 B.n471 585
R238 B.n474 B.n247 585
R239 B.n247 B.n246 585
R240 B.n476 B.n475 585
R241 B.n477 B.n476 585
R242 B.n241 B.n240 585
R243 B.n242 B.n241 585
R244 B.n485 B.n484 585
R245 B.n484 B.n483 585
R246 B.n486 B.n239 585
R247 B.n239 B.n238 585
R248 B.n488 B.n487 585
R249 B.n489 B.n488 585
R250 B.n233 B.n232 585
R251 B.n234 B.n233 585
R252 B.n498 B.n497 585
R253 B.n497 B.n496 585
R254 B.n499 B.n231 585
R255 B.n231 B.n230 585
R256 B.n501 B.n500 585
R257 B.n502 B.n501 585
R258 B.n3 B.n0 585
R259 B.n4 B.n3 585
R260 B.n566 B.n1 585
R261 B.n567 B.n566 585
R262 B.n565 B.n564 585
R263 B.n565 B.n8 585
R264 B.n563 B.n9 585
R265 B.n511 B.n9 585
R266 B.n562 B.n561 585
R267 B.n561 B.n560 585
R268 B.n11 B.n10 585
R269 B.n559 B.n11 585
R270 B.n557 B.n556 585
R271 B.n558 B.n557 585
R272 B.n555 B.n16 585
R273 B.n16 B.n15 585
R274 B.n554 B.n553 585
R275 B.n553 B.n552 585
R276 B.n18 B.n17 585
R277 B.n551 B.n18 585
R278 B.n549 B.n548 585
R279 B.n550 B.n549 585
R280 B.n547 B.n23 585
R281 B.n23 B.n22 585
R282 B.n546 B.n545 585
R283 B.n545 B.n544 585
R284 B.n25 B.n24 585
R285 B.n543 B.n25 585
R286 B.n541 B.n540 585
R287 B.n542 B.n541 585
R288 B.n539 B.n30 585
R289 B.n30 B.n29 585
R290 B.n538 B.n537 585
R291 B.n537 B.n536 585
R292 B.n32 B.n31 585
R293 B.n535 B.n32 585
R294 B.n570 B.n569 585
R295 B.n568 B.n2 585
R296 B.n77 B.n32 554.963
R297 B.n532 B.n34 554.963
R298 B.n454 B.n259 554.963
R299 B.n451 B.n257 554.963
R300 B.n75 B.t6 373.356
R301 B.n73 B.t10 373.356
R302 B.n303 B.t2 373.356
R303 B.n300 B.t13 373.356
R304 B.n534 B.n533 256.663
R305 B.n534 B.n71 256.663
R306 B.n534 B.n70 256.663
R307 B.n534 B.n69 256.663
R308 B.n534 B.n68 256.663
R309 B.n534 B.n67 256.663
R310 B.n534 B.n66 256.663
R311 B.n534 B.n65 256.663
R312 B.n534 B.n64 256.663
R313 B.n534 B.n63 256.663
R314 B.n534 B.n62 256.663
R315 B.n534 B.n61 256.663
R316 B.n534 B.n60 256.663
R317 B.n534 B.n59 256.663
R318 B.n534 B.n58 256.663
R319 B.n534 B.n57 256.663
R320 B.n534 B.n56 256.663
R321 B.n534 B.n55 256.663
R322 B.n534 B.n54 256.663
R323 B.n534 B.n53 256.663
R324 B.n534 B.n52 256.663
R325 B.n534 B.n51 256.663
R326 B.n534 B.n50 256.663
R327 B.n534 B.n49 256.663
R328 B.n534 B.n48 256.663
R329 B.n534 B.n47 256.663
R330 B.n534 B.n46 256.663
R331 B.n534 B.n45 256.663
R332 B.n534 B.n44 256.663
R333 B.n534 B.n43 256.663
R334 B.n534 B.n42 256.663
R335 B.n534 B.n41 256.663
R336 B.n534 B.n40 256.663
R337 B.n534 B.n39 256.663
R338 B.n534 B.n38 256.663
R339 B.n534 B.n37 256.663
R340 B.n534 B.n36 256.663
R341 B.n534 B.n35 256.663
R342 B.n453 B.n452 256.663
R343 B.n453 B.n262 256.663
R344 B.n453 B.n263 256.663
R345 B.n453 B.n264 256.663
R346 B.n453 B.n265 256.663
R347 B.n453 B.n266 256.663
R348 B.n453 B.n267 256.663
R349 B.n453 B.n268 256.663
R350 B.n453 B.n269 256.663
R351 B.n453 B.n270 256.663
R352 B.n453 B.n271 256.663
R353 B.n453 B.n272 256.663
R354 B.n453 B.n273 256.663
R355 B.n453 B.n274 256.663
R356 B.n453 B.n275 256.663
R357 B.n453 B.n276 256.663
R358 B.n453 B.n277 256.663
R359 B.n453 B.n278 256.663
R360 B.n453 B.n279 256.663
R361 B.n453 B.n280 256.663
R362 B.n453 B.n281 256.663
R363 B.n453 B.n282 256.663
R364 B.n453 B.n283 256.663
R365 B.n453 B.n284 256.663
R366 B.n453 B.n285 256.663
R367 B.n453 B.n286 256.663
R368 B.n453 B.n287 256.663
R369 B.n453 B.n288 256.663
R370 B.n453 B.n289 256.663
R371 B.n453 B.n290 256.663
R372 B.n453 B.n291 256.663
R373 B.n453 B.n292 256.663
R374 B.n453 B.n293 256.663
R375 B.n453 B.n294 256.663
R376 B.n453 B.n295 256.663
R377 B.n453 B.n296 256.663
R378 B.n453 B.n297 256.663
R379 B.n572 B.n571 256.663
R380 B.n81 B.n80 163.367
R381 B.n85 B.n84 163.367
R382 B.n89 B.n88 163.367
R383 B.n93 B.n92 163.367
R384 B.n97 B.n96 163.367
R385 B.n101 B.n100 163.367
R386 B.n105 B.n104 163.367
R387 B.n109 B.n108 163.367
R388 B.n113 B.n112 163.367
R389 B.n117 B.n116 163.367
R390 B.n121 B.n120 163.367
R391 B.n125 B.n124 163.367
R392 B.n129 B.n128 163.367
R393 B.n133 B.n132 163.367
R394 B.n137 B.n136 163.367
R395 B.n141 B.n140 163.367
R396 B.n146 B.n145 163.367
R397 B.n150 B.n149 163.367
R398 B.n154 B.n153 163.367
R399 B.n158 B.n157 163.367
R400 B.n162 B.n161 163.367
R401 B.n167 B.n166 163.367
R402 B.n171 B.n170 163.367
R403 B.n175 B.n174 163.367
R404 B.n179 B.n178 163.367
R405 B.n183 B.n182 163.367
R406 B.n187 B.n186 163.367
R407 B.n191 B.n190 163.367
R408 B.n195 B.n194 163.367
R409 B.n199 B.n198 163.367
R410 B.n203 B.n202 163.367
R411 B.n207 B.n206 163.367
R412 B.n211 B.n210 163.367
R413 B.n215 B.n214 163.367
R414 B.n219 B.n218 163.367
R415 B.n223 B.n222 163.367
R416 B.n225 B.n72 163.367
R417 B.n458 B.n259 163.367
R418 B.n458 B.n253 163.367
R419 B.n466 B.n253 163.367
R420 B.n466 B.n251 163.367
R421 B.n470 B.n251 163.367
R422 B.n470 B.n245 163.367
R423 B.n478 B.n245 163.367
R424 B.n478 B.n243 163.367
R425 B.n482 B.n243 163.367
R426 B.n482 B.n237 163.367
R427 B.n490 B.n237 163.367
R428 B.n490 B.n235 163.367
R429 B.n495 B.n235 163.367
R430 B.n495 B.n229 163.367
R431 B.n503 B.n229 163.367
R432 B.n504 B.n503 163.367
R433 B.n504 B.n5 163.367
R434 B.n6 B.n5 163.367
R435 B.n7 B.n6 163.367
R436 B.n510 B.n7 163.367
R437 B.n512 B.n510 163.367
R438 B.n512 B.n12 163.367
R439 B.n13 B.n12 163.367
R440 B.n14 B.n13 163.367
R441 B.n517 B.n14 163.367
R442 B.n517 B.n19 163.367
R443 B.n20 B.n19 163.367
R444 B.n21 B.n20 163.367
R445 B.n522 B.n21 163.367
R446 B.n522 B.n26 163.367
R447 B.n27 B.n26 163.367
R448 B.n28 B.n27 163.367
R449 B.n527 B.n28 163.367
R450 B.n527 B.n33 163.367
R451 B.n34 B.n33 163.367
R452 B.n299 B.n298 163.367
R453 B.n446 B.n298 163.367
R454 B.n444 B.n443 163.367
R455 B.n440 B.n439 163.367
R456 B.n436 B.n435 163.367
R457 B.n432 B.n431 163.367
R458 B.n428 B.n427 163.367
R459 B.n424 B.n423 163.367
R460 B.n420 B.n419 163.367
R461 B.n416 B.n415 163.367
R462 B.n412 B.n411 163.367
R463 B.n408 B.n407 163.367
R464 B.n404 B.n403 163.367
R465 B.n400 B.n399 163.367
R466 B.n396 B.n395 163.367
R467 B.n392 B.n391 163.367
R468 B.n388 B.n387 163.367
R469 B.n384 B.n383 163.367
R470 B.n380 B.n379 163.367
R471 B.n376 B.n375 163.367
R472 B.n372 B.n371 163.367
R473 B.n368 B.n367 163.367
R474 B.n364 B.n363 163.367
R475 B.n360 B.n359 163.367
R476 B.n356 B.n355 163.367
R477 B.n352 B.n351 163.367
R478 B.n348 B.n347 163.367
R479 B.n344 B.n343 163.367
R480 B.n340 B.n339 163.367
R481 B.n336 B.n335 163.367
R482 B.n332 B.n331 163.367
R483 B.n328 B.n327 163.367
R484 B.n324 B.n323 163.367
R485 B.n320 B.n319 163.367
R486 B.n316 B.n315 163.367
R487 B.n312 B.n311 163.367
R488 B.n308 B.n307 163.367
R489 B.n454 B.n261 163.367
R490 B.n460 B.n257 163.367
R491 B.n460 B.n255 163.367
R492 B.n464 B.n255 163.367
R493 B.n464 B.n249 163.367
R494 B.n472 B.n249 163.367
R495 B.n472 B.n247 163.367
R496 B.n476 B.n247 163.367
R497 B.n476 B.n241 163.367
R498 B.n484 B.n241 163.367
R499 B.n484 B.n239 163.367
R500 B.n488 B.n239 163.367
R501 B.n488 B.n233 163.367
R502 B.n497 B.n233 163.367
R503 B.n497 B.n231 163.367
R504 B.n501 B.n231 163.367
R505 B.n501 B.n3 163.367
R506 B.n570 B.n3 163.367
R507 B.n566 B.n2 163.367
R508 B.n566 B.n565 163.367
R509 B.n565 B.n9 163.367
R510 B.n561 B.n9 163.367
R511 B.n561 B.n11 163.367
R512 B.n557 B.n11 163.367
R513 B.n557 B.n16 163.367
R514 B.n553 B.n16 163.367
R515 B.n553 B.n18 163.367
R516 B.n549 B.n18 163.367
R517 B.n549 B.n23 163.367
R518 B.n545 B.n23 163.367
R519 B.n545 B.n25 163.367
R520 B.n541 B.n25 163.367
R521 B.n541 B.n30 163.367
R522 B.n537 B.n30 163.367
R523 B.n537 B.n32 163.367
R524 B.n453 B.n258 107.374
R525 B.n535 B.n534 107.374
R526 B.n73 B.t11 106.501
R527 B.n303 B.t5 106.501
R528 B.n75 B.t8 106.49
R529 B.n300 B.t15 106.49
R530 B.n74 B.t12 74.6948
R531 B.n304 B.t4 74.6948
R532 B.n76 B.t9 74.684
R533 B.n301 B.t14 74.684
R534 B.n77 B.n35 71.676
R535 B.n81 B.n36 71.676
R536 B.n85 B.n37 71.676
R537 B.n89 B.n38 71.676
R538 B.n93 B.n39 71.676
R539 B.n97 B.n40 71.676
R540 B.n101 B.n41 71.676
R541 B.n105 B.n42 71.676
R542 B.n109 B.n43 71.676
R543 B.n113 B.n44 71.676
R544 B.n117 B.n45 71.676
R545 B.n121 B.n46 71.676
R546 B.n125 B.n47 71.676
R547 B.n129 B.n48 71.676
R548 B.n133 B.n49 71.676
R549 B.n137 B.n50 71.676
R550 B.n141 B.n51 71.676
R551 B.n146 B.n52 71.676
R552 B.n150 B.n53 71.676
R553 B.n154 B.n54 71.676
R554 B.n158 B.n55 71.676
R555 B.n162 B.n56 71.676
R556 B.n167 B.n57 71.676
R557 B.n171 B.n58 71.676
R558 B.n175 B.n59 71.676
R559 B.n179 B.n60 71.676
R560 B.n183 B.n61 71.676
R561 B.n187 B.n62 71.676
R562 B.n191 B.n63 71.676
R563 B.n195 B.n64 71.676
R564 B.n199 B.n65 71.676
R565 B.n203 B.n66 71.676
R566 B.n207 B.n67 71.676
R567 B.n211 B.n68 71.676
R568 B.n215 B.n69 71.676
R569 B.n219 B.n70 71.676
R570 B.n223 B.n71 71.676
R571 B.n533 B.n72 71.676
R572 B.n533 B.n532 71.676
R573 B.n225 B.n71 71.676
R574 B.n222 B.n70 71.676
R575 B.n218 B.n69 71.676
R576 B.n214 B.n68 71.676
R577 B.n210 B.n67 71.676
R578 B.n206 B.n66 71.676
R579 B.n202 B.n65 71.676
R580 B.n198 B.n64 71.676
R581 B.n194 B.n63 71.676
R582 B.n190 B.n62 71.676
R583 B.n186 B.n61 71.676
R584 B.n182 B.n60 71.676
R585 B.n178 B.n59 71.676
R586 B.n174 B.n58 71.676
R587 B.n170 B.n57 71.676
R588 B.n166 B.n56 71.676
R589 B.n161 B.n55 71.676
R590 B.n157 B.n54 71.676
R591 B.n153 B.n53 71.676
R592 B.n149 B.n52 71.676
R593 B.n145 B.n51 71.676
R594 B.n140 B.n50 71.676
R595 B.n136 B.n49 71.676
R596 B.n132 B.n48 71.676
R597 B.n128 B.n47 71.676
R598 B.n124 B.n46 71.676
R599 B.n120 B.n45 71.676
R600 B.n116 B.n44 71.676
R601 B.n112 B.n43 71.676
R602 B.n108 B.n42 71.676
R603 B.n104 B.n41 71.676
R604 B.n100 B.n40 71.676
R605 B.n96 B.n39 71.676
R606 B.n92 B.n38 71.676
R607 B.n88 B.n37 71.676
R608 B.n84 B.n36 71.676
R609 B.n80 B.n35 71.676
R610 B.n452 B.n451 71.676
R611 B.n446 B.n262 71.676
R612 B.n443 B.n263 71.676
R613 B.n439 B.n264 71.676
R614 B.n435 B.n265 71.676
R615 B.n431 B.n266 71.676
R616 B.n427 B.n267 71.676
R617 B.n423 B.n268 71.676
R618 B.n419 B.n269 71.676
R619 B.n415 B.n270 71.676
R620 B.n411 B.n271 71.676
R621 B.n407 B.n272 71.676
R622 B.n403 B.n273 71.676
R623 B.n399 B.n274 71.676
R624 B.n395 B.n275 71.676
R625 B.n391 B.n276 71.676
R626 B.n387 B.n277 71.676
R627 B.n383 B.n278 71.676
R628 B.n379 B.n279 71.676
R629 B.n375 B.n280 71.676
R630 B.n371 B.n281 71.676
R631 B.n367 B.n282 71.676
R632 B.n363 B.n283 71.676
R633 B.n359 B.n284 71.676
R634 B.n355 B.n285 71.676
R635 B.n351 B.n286 71.676
R636 B.n347 B.n287 71.676
R637 B.n343 B.n288 71.676
R638 B.n339 B.n289 71.676
R639 B.n335 B.n290 71.676
R640 B.n331 B.n291 71.676
R641 B.n327 B.n292 71.676
R642 B.n323 B.n293 71.676
R643 B.n319 B.n294 71.676
R644 B.n315 B.n295 71.676
R645 B.n311 B.n296 71.676
R646 B.n307 B.n297 71.676
R647 B.n452 B.n299 71.676
R648 B.n444 B.n262 71.676
R649 B.n440 B.n263 71.676
R650 B.n436 B.n264 71.676
R651 B.n432 B.n265 71.676
R652 B.n428 B.n266 71.676
R653 B.n424 B.n267 71.676
R654 B.n420 B.n268 71.676
R655 B.n416 B.n269 71.676
R656 B.n412 B.n270 71.676
R657 B.n408 B.n271 71.676
R658 B.n404 B.n272 71.676
R659 B.n400 B.n273 71.676
R660 B.n396 B.n274 71.676
R661 B.n392 B.n275 71.676
R662 B.n388 B.n276 71.676
R663 B.n384 B.n277 71.676
R664 B.n380 B.n278 71.676
R665 B.n376 B.n279 71.676
R666 B.n372 B.n280 71.676
R667 B.n368 B.n281 71.676
R668 B.n364 B.n282 71.676
R669 B.n360 B.n283 71.676
R670 B.n356 B.n284 71.676
R671 B.n352 B.n285 71.676
R672 B.n348 B.n286 71.676
R673 B.n344 B.n287 71.676
R674 B.n340 B.n288 71.676
R675 B.n336 B.n289 71.676
R676 B.n332 B.n290 71.676
R677 B.n328 B.n291 71.676
R678 B.n324 B.n292 71.676
R679 B.n320 B.n293 71.676
R680 B.n316 B.n294 71.676
R681 B.n312 B.n295 71.676
R682 B.n308 B.n296 71.676
R683 B.n297 B.n261 71.676
R684 B.n571 B.n570 71.676
R685 B.n571 B.n2 71.676
R686 B.n143 B.n76 59.5399
R687 B.n164 B.n74 59.5399
R688 B.n305 B.n304 59.5399
R689 B.n302 B.n301 59.5399
R690 B.n459 B.n258 51.7831
R691 B.n459 B.n254 51.7831
R692 B.n465 B.n254 51.7831
R693 B.n465 B.n250 51.7831
R694 B.n471 B.n250 51.7831
R695 B.n477 B.n246 51.7831
R696 B.n477 B.n242 51.7831
R697 B.n483 B.n242 51.7831
R698 B.n483 B.n238 51.7831
R699 B.n489 B.n238 51.7831
R700 B.n489 B.n234 51.7831
R701 B.n496 B.n234 51.7831
R702 B.n502 B.n230 51.7831
R703 B.n502 B.n4 51.7831
R704 B.n569 B.n4 51.7831
R705 B.n569 B.n568 51.7831
R706 B.n568 B.n567 51.7831
R707 B.n567 B.n8 51.7831
R708 B.n511 B.n8 51.7831
R709 B.n560 B.n559 51.7831
R710 B.n559 B.n558 51.7831
R711 B.n558 B.n15 51.7831
R712 B.n552 B.n15 51.7831
R713 B.n552 B.n551 51.7831
R714 B.n551 B.n550 51.7831
R715 B.n550 B.n22 51.7831
R716 B.n544 B.n543 51.7831
R717 B.n543 B.n542 51.7831
R718 B.n542 B.n29 51.7831
R719 B.n536 B.n29 51.7831
R720 B.n536 B.n535 51.7831
R721 B.n531 B.n530 36.059
R722 B.n450 B.n256 36.059
R723 B.n456 B.n455 36.059
R724 B.n78 B.n31 36.059
R725 B.n76 B.n75 31.8066
R726 B.n74 B.n73 31.8066
R727 B.n304 B.n303 31.8066
R728 B.n301 B.n300 31.8066
R729 B.t3 B.n246 28.1763
R730 B.t7 B.n22 28.1763
R731 B.t1 B.n230 26.6533
R732 B.n511 B.t0 26.6533
R733 B.n496 B.t1 25.1303
R734 B.n560 B.t0 25.1303
R735 B.n471 B.t3 23.6073
R736 B.n544 B.t7 23.6073
R737 B B.n572 18.0485
R738 B.n461 B.n256 10.6151
R739 B.n462 B.n461 10.6151
R740 B.n463 B.n462 10.6151
R741 B.n463 B.n248 10.6151
R742 B.n473 B.n248 10.6151
R743 B.n474 B.n473 10.6151
R744 B.n475 B.n474 10.6151
R745 B.n475 B.n240 10.6151
R746 B.n485 B.n240 10.6151
R747 B.n486 B.n485 10.6151
R748 B.n487 B.n486 10.6151
R749 B.n487 B.n232 10.6151
R750 B.n498 B.n232 10.6151
R751 B.n499 B.n498 10.6151
R752 B.n500 B.n499 10.6151
R753 B.n500 B.n0 10.6151
R754 B.n450 B.n449 10.6151
R755 B.n449 B.n448 10.6151
R756 B.n448 B.n447 10.6151
R757 B.n447 B.n445 10.6151
R758 B.n445 B.n442 10.6151
R759 B.n442 B.n441 10.6151
R760 B.n441 B.n438 10.6151
R761 B.n438 B.n437 10.6151
R762 B.n437 B.n434 10.6151
R763 B.n434 B.n433 10.6151
R764 B.n433 B.n430 10.6151
R765 B.n430 B.n429 10.6151
R766 B.n429 B.n426 10.6151
R767 B.n426 B.n425 10.6151
R768 B.n425 B.n422 10.6151
R769 B.n422 B.n421 10.6151
R770 B.n421 B.n418 10.6151
R771 B.n418 B.n417 10.6151
R772 B.n417 B.n414 10.6151
R773 B.n414 B.n413 10.6151
R774 B.n413 B.n410 10.6151
R775 B.n410 B.n409 10.6151
R776 B.n409 B.n406 10.6151
R777 B.n406 B.n405 10.6151
R778 B.n405 B.n402 10.6151
R779 B.n402 B.n401 10.6151
R780 B.n401 B.n398 10.6151
R781 B.n398 B.n397 10.6151
R782 B.n397 B.n394 10.6151
R783 B.n394 B.n393 10.6151
R784 B.n393 B.n390 10.6151
R785 B.n390 B.n389 10.6151
R786 B.n386 B.n385 10.6151
R787 B.n385 B.n382 10.6151
R788 B.n382 B.n381 10.6151
R789 B.n381 B.n378 10.6151
R790 B.n378 B.n377 10.6151
R791 B.n377 B.n374 10.6151
R792 B.n374 B.n373 10.6151
R793 B.n373 B.n370 10.6151
R794 B.n370 B.n369 10.6151
R795 B.n366 B.n365 10.6151
R796 B.n365 B.n362 10.6151
R797 B.n362 B.n361 10.6151
R798 B.n361 B.n358 10.6151
R799 B.n358 B.n357 10.6151
R800 B.n357 B.n354 10.6151
R801 B.n354 B.n353 10.6151
R802 B.n353 B.n350 10.6151
R803 B.n350 B.n349 10.6151
R804 B.n349 B.n346 10.6151
R805 B.n346 B.n345 10.6151
R806 B.n345 B.n342 10.6151
R807 B.n342 B.n341 10.6151
R808 B.n341 B.n338 10.6151
R809 B.n338 B.n337 10.6151
R810 B.n337 B.n334 10.6151
R811 B.n334 B.n333 10.6151
R812 B.n333 B.n330 10.6151
R813 B.n330 B.n329 10.6151
R814 B.n329 B.n326 10.6151
R815 B.n326 B.n325 10.6151
R816 B.n325 B.n322 10.6151
R817 B.n322 B.n321 10.6151
R818 B.n321 B.n318 10.6151
R819 B.n318 B.n317 10.6151
R820 B.n317 B.n314 10.6151
R821 B.n314 B.n313 10.6151
R822 B.n313 B.n310 10.6151
R823 B.n310 B.n309 10.6151
R824 B.n309 B.n306 10.6151
R825 B.n306 B.n260 10.6151
R826 B.n455 B.n260 10.6151
R827 B.n457 B.n456 10.6151
R828 B.n457 B.n252 10.6151
R829 B.n467 B.n252 10.6151
R830 B.n468 B.n467 10.6151
R831 B.n469 B.n468 10.6151
R832 B.n469 B.n244 10.6151
R833 B.n479 B.n244 10.6151
R834 B.n480 B.n479 10.6151
R835 B.n481 B.n480 10.6151
R836 B.n481 B.n236 10.6151
R837 B.n491 B.n236 10.6151
R838 B.n492 B.n491 10.6151
R839 B.n494 B.n492 10.6151
R840 B.n494 B.n493 10.6151
R841 B.n493 B.n228 10.6151
R842 B.n505 B.n228 10.6151
R843 B.n506 B.n505 10.6151
R844 B.n507 B.n506 10.6151
R845 B.n508 B.n507 10.6151
R846 B.n509 B.n508 10.6151
R847 B.n513 B.n509 10.6151
R848 B.n514 B.n513 10.6151
R849 B.n515 B.n514 10.6151
R850 B.n516 B.n515 10.6151
R851 B.n518 B.n516 10.6151
R852 B.n519 B.n518 10.6151
R853 B.n520 B.n519 10.6151
R854 B.n521 B.n520 10.6151
R855 B.n523 B.n521 10.6151
R856 B.n524 B.n523 10.6151
R857 B.n525 B.n524 10.6151
R858 B.n526 B.n525 10.6151
R859 B.n528 B.n526 10.6151
R860 B.n529 B.n528 10.6151
R861 B.n530 B.n529 10.6151
R862 B.n564 B.n1 10.6151
R863 B.n564 B.n563 10.6151
R864 B.n563 B.n562 10.6151
R865 B.n562 B.n10 10.6151
R866 B.n556 B.n10 10.6151
R867 B.n556 B.n555 10.6151
R868 B.n555 B.n554 10.6151
R869 B.n554 B.n17 10.6151
R870 B.n548 B.n17 10.6151
R871 B.n548 B.n547 10.6151
R872 B.n547 B.n546 10.6151
R873 B.n546 B.n24 10.6151
R874 B.n540 B.n24 10.6151
R875 B.n540 B.n539 10.6151
R876 B.n539 B.n538 10.6151
R877 B.n538 B.n31 10.6151
R878 B.n79 B.n78 10.6151
R879 B.n82 B.n79 10.6151
R880 B.n83 B.n82 10.6151
R881 B.n86 B.n83 10.6151
R882 B.n87 B.n86 10.6151
R883 B.n90 B.n87 10.6151
R884 B.n91 B.n90 10.6151
R885 B.n94 B.n91 10.6151
R886 B.n95 B.n94 10.6151
R887 B.n98 B.n95 10.6151
R888 B.n99 B.n98 10.6151
R889 B.n102 B.n99 10.6151
R890 B.n103 B.n102 10.6151
R891 B.n106 B.n103 10.6151
R892 B.n107 B.n106 10.6151
R893 B.n110 B.n107 10.6151
R894 B.n111 B.n110 10.6151
R895 B.n114 B.n111 10.6151
R896 B.n115 B.n114 10.6151
R897 B.n118 B.n115 10.6151
R898 B.n119 B.n118 10.6151
R899 B.n122 B.n119 10.6151
R900 B.n123 B.n122 10.6151
R901 B.n126 B.n123 10.6151
R902 B.n127 B.n126 10.6151
R903 B.n130 B.n127 10.6151
R904 B.n131 B.n130 10.6151
R905 B.n134 B.n131 10.6151
R906 B.n135 B.n134 10.6151
R907 B.n138 B.n135 10.6151
R908 B.n139 B.n138 10.6151
R909 B.n142 B.n139 10.6151
R910 B.n147 B.n144 10.6151
R911 B.n148 B.n147 10.6151
R912 B.n151 B.n148 10.6151
R913 B.n152 B.n151 10.6151
R914 B.n155 B.n152 10.6151
R915 B.n156 B.n155 10.6151
R916 B.n159 B.n156 10.6151
R917 B.n160 B.n159 10.6151
R918 B.n163 B.n160 10.6151
R919 B.n168 B.n165 10.6151
R920 B.n169 B.n168 10.6151
R921 B.n172 B.n169 10.6151
R922 B.n173 B.n172 10.6151
R923 B.n176 B.n173 10.6151
R924 B.n177 B.n176 10.6151
R925 B.n180 B.n177 10.6151
R926 B.n181 B.n180 10.6151
R927 B.n184 B.n181 10.6151
R928 B.n185 B.n184 10.6151
R929 B.n188 B.n185 10.6151
R930 B.n189 B.n188 10.6151
R931 B.n192 B.n189 10.6151
R932 B.n193 B.n192 10.6151
R933 B.n196 B.n193 10.6151
R934 B.n197 B.n196 10.6151
R935 B.n200 B.n197 10.6151
R936 B.n201 B.n200 10.6151
R937 B.n204 B.n201 10.6151
R938 B.n205 B.n204 10.6151
R939 B.n208 B.n205 10.6151
R940 B.n209 B.n208 10.6151
R941 B.n212 B.n209 10.6151
R942 B.n213 B.n212 10.6151
R943 B.n216 B.n213 10.6151
R944 B.n217 B.n216 10.6151
R945 B.n220 B.n217 10.6151
R946 B.n221 B.n220 10.6151
R947 B.n224 B.n221 10.6151
R948 B.n226 B.n224 10.6151
R949 B.n227 B.n226 10.6151
R950 B.n531 B.n227 10.6151
R951 B.n389 B.n302 9.36635
R952 B.n366 B.n305 9.36635
R953 B.n143 B.n142 9.36635
R954 B.n165 B.n164 9.36635
R955 B.n572 B.n0 8.11757
R956 B.n572 B.n1 8.11757
R957 B.n386 B.n302 1.24928
R958 B.n369 B.n305 1.24928
R959 B.n144 B.n143 1.24928
R960 B.n164 B.n163 1.24928
R961 VP.n0 VP.t1 318.567
R962 VP.n0 VP.t0 279.474
R963 VP VP.n0 0.146778
R964 VTAIL.n2 VTAIL.t3 47.8176
R965 VTAIL.n1 VTAIL.t1 47.8176
R966 VTAIL.n3 VTAIL.t0 47.8174
R967 VTAIL.n0 VTAIL.t2 47.8174
R968 VTAIL.n1 VTAIL.n0 23.0996
R969 VTAIL.n3 VTAIL.n2 21.6858
R970 VTAIL.n2 VTAIL.n1 1.17722
R971 VTAIL VTAIL.n0 0.881965
R972 VTAIL VTAIL.n3 0.295759
R973 VDD1 VDD1.t1 99.7667
R974 VDD1 VDD1.t0 64.908
R975 VN VN.t1 318.853
R976 VN VN.t0 279.62
R977 VDD2.n0 VDD2.t1 98.8884
R978 VDD2.n0 VDD2.t0 64.4964
R979 VDD2 VDD2.n0 0.412138
C0 VTAIL VDD2 4.29581f
C1 VDD1 VDD2 0.524612f
C2 VDD1 VTAIL 4.25482f
C3 VDD2 VP 0.278715f
C4 VDD2 VN 1.90156f
C5 VTAIL VP 1.61279f
C6 VTAIL VN 1.59842f
C7 VDD1 VP 2.02999f
C8 VDD1 VN 0.147531f
C9 VN VP 4.32674f
C10 VDD2 B 3.443923f
C11 VDD1 B 6.10405f
C12 VTAIL B 5.559774f
C13 VN B 6.91503f
C14 VP B 4.591925f
C15 VDD2.t1 B 1.42507f
C16 VDD2.t0 B 1.13829f
C17 VDD2.n0 B 1.68514f
C18 VN.t0 B 0.950875f
C19 VN.t1 B 1.09702f
C20 VDD1.t0 B 1.64932f
C21 VDD1.t1 B 2.0895f
C22 VTAIL.t2 B 1.17842f
C23 VTAIL.n0 B 0.992011f
C24 VTAIL.t1 B 1.17843f
C25 VTAIL.n1 B 1.00666f
C26 VTAIL.t3 B 1.17843f
C27 VTAIL.n2 B 0.936489f
C28 VTAIL.t0 B 1.17842f
C29 VTAIL.n3 B 0.892746f
C30 VP.t1 B 1.61642f
C31 VP.t0 B 1.40426f
C32 VP.n0 B 3.24576f
.ends

