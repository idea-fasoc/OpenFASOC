* NGSPICE file created from diff_pair_sample_0814.ext - technology: sky130A

.subckt diff_pair_sample_0814 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t11 VN.t0 VDD2.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=3.24555 ps=20 w=19.67 l=3.13
X1 VDD1.t5 VP.t0 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.13
X2 VTAIL.t10 VN.t1 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=3.24555 ps=20 w=19.67 l=3.13
X3 VDD2.t3 VN.t2 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.13
X4 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.13
X5 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.13
X6 VDD2.t4 VN.t3 VTAIL.t8 B.t4 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.13
X7 VDD1.t4 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.13
X8 VTAIL.t1 VP.t2 VDD1.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=3.24555 ps=20 w=19.67 l=3.13
X9 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.13
X10 VDD2.t0 VN.t4 VTAIL.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=3.24555 ps=20 w=19.67 l=3.13
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.6713 pd=40.12 as=0 ps=0 w=19.67 l=3.13
X12 VDD1.t2 VP.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.13
X13 VTAIL.t0 VP.t4 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=3.24555 ps=20 w=19.67 l=3.13
X14 VDD2.t2 VN.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.13
X15 VDD1.t0 VP.t5 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=3.24555 pd=20 as=7.6713 ps=40.12 w=19.67 l=3.13
R0 VN.n20 VN.t3 184.864
R1 VN.n4 VN.t2 184.864
R2 VN.n30 VN.n29 161.3
R3 VN.n28 VN.n17 161.3
R4 VN.n27 VN.n26 161.3
R5 VN.n25 VN.n18 161.3
R6 VN.n24 VN.n23 161.3
R7 VN.n22 VN.n19 161.3
R8 VN.n14 VN.n13 161.3
R9 VN.n12 VN.n1 161.3
R10 VN.n11 VN.n10 161.3
R11 VN.n9 VN.n2 161.3
R12 VN.n8 VN.n7 161.3
R13 VN.n6 VN.n3 161.3
R14 VN.n5 VN.t1 151.453
R15 VN.n0 VN.t5 151.453
R16 VN.n21 VN.t0 151.453
R17 VN.n16 VN.t4 151.453
R18 VN.n15 VN.n0 67.5578
R19 VN.n31 VN.n16 67.5578
R20 VN VN.n31 56.9223
R21 VN.n11 VN.n2 56.5193
R22 VN.n27 VN.n18 56.5193
R23 VN.n21 VN.n20 49.5199
R24 VN.n5 VN.n4 49.5199
R25 VN.n6 VN.n5 24.4675
R26 VN.n7 VN.n6 24.4675
R27 VN.n7 VN.n2 24.4675
R28 VN.n12 VN.n11 24.4675
R29 VN.n13 VN.n12 24.4675
R30 VN.n23 VN.n18 24.4675
R31 VN.n23 VN.n22 24.4675
R32 VN.n22 VN.n21 24.4675
R33 VN.n29 VN.n28 24.4675
R34 VN.n28 VN.n27 24.4675
R35 VN.n13 VN.n0 22.5101
R36 VN.n29 VN.n16 22.5101
R37 VN.n20 VN.n19 3.79387
R38 VN.n4 VN.n3 3.79387
R39 VN.n31 VN.n30 0.354971
R40 VN.n15 VN.n14 0.354971
R41 VN VN.n15 0.26696
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VDD2.n215 VDD2.n111 289.615
R53 VDD2.n104 VDD2.n0 289.615
R54 VDD2.n216 VDD2.n215 185
R55 VDD2.n214 VDD2.n213 185
R56 VDD2.n115 VDD2.n114 185
R57 VDD2.n208 VDD2.n207 185
R58 VDD2.n206 VDD2.n205 185
R59 VDD2.n119 VDD2.n118 185
R60 VDD2.n200 VDD2.n199 185
R61 VDD2.n198 VDD2.n197 185
R62 VDD2.n123 VDD2.n122 185
R63 VDD2.n127 VDD2.n125 185
R64 VDD2.n192 VDD2.n191 185
R65 VDD2.n190 VDD2.n189 185
R66 VDD2.n129 VDD2.n128 185
R67 VDD2.n184 VDD2.n183 185
R68 VDD2.n182 VDD2.n181 185
R69 VDD2.n133 VDD2.n132 185
R70 VDD2.n176 VDD2.n175 185
R71 VDD2.n174 VDD2.n173 185
R72 VDD2.n137 VDD2.n136 185
R73 VDD2.n168 VDD2.n167 185
R74 VDD2.n166 VDD2.n165 185
R75 VDD2.n141 VDD2.n140 185
R76 VDD2.n160 VDD2.n159 185
R77 VDD2.n158 VDD2.n157 185
R78 VDD2.n145 VDD2.n144 185
R79 VDD2.n152 VDD2.n151 185
R80 VDD2.n150 VDD2.n149 185
R81 VDD2.n37 VDD2.n36 185
R82 VDD2.n39 VDD2.n38 185
R83 VDD2.n32 VDD2.n31 185
R84 VDD2.n45 VDD2.n44 185
R85 VDD2.n47 VDD2.n46 185
R86 VDD2.n28 VDD2.n27 185
R87 VDD2.n53 VDD2.n52 185
R88 VDD2.n55 VDD2.n54 185
R89 VDD2.n24 VDD2.n23 185
R90 VDD2.n61 VDD2.n60 185
R91 VDD2.n63 VDD2.n62 185
R92 VDD2.n20 VDD2.n19 185
R93 VDD2.n69 VDD2.n68 185
R94 VDD2.n71 VDD2.n70 185
R95 VDD2.n16 VDD2.n15 185
R96 VDD2.n78 VDD2.n77 185
R97 VDD2.n79 VDD2.n14 185
R98 VDD2.n81 VDD2.n80 185
R99 VDD2.n12 VDD2.n11 185
R100 VDD2.n87 VDD2.n86 185
R101 VDD2.n89 VDD2.n88 185
R102 VDD2.n8 VDD2.n7 185
R103 VDD2.n95 VDD2.n94 185
R104 VDD2.n97 VDD2.n96 185
R105 VDD2.n4 VDD2.n3 185
R106 VDD2.n103 VDD2.n102 185
R107 VDD2.n105 VDD2.n104 185
R108 VDD2.n148 VDD2.t0 147.659
R109 VDD2.n35 VDD2.t3 147.659
R110 VDD2.n215 VDD2.n214 104.615
R111 VDD2.n214 VDD2.n114 104.615
R112 VDD2.n207 VDD2.n114 104.615
R113 VDD2.n207 VDD2.n206 104.615
R114 VDD2.n206 VDD2.n118 104.615
R115 VDD2.n199 VDD2.n118 104.615
R116 VDD2.n199 VDD2.n198 104.615
R117 VDD2.n198 VDD2.n122 104.615
R118 VDD2.n127 VDD2.n122 104.615
R119 VDD2.n191 VDD2.n127 104.615
R120 VDD2.n191 VDD2.n190 104.615
R121 VDD2.n190 VDD2.n128 104.615
R122 VDD2.n183 VDD2.n128 104.615
R123 VDD2.n183 VDD2.n182 104.615
R124 VDD2.n182 VDD2.n132 104.615
R125 VDD2.n175 VDD2.n132 104.615
R126 VDD2.n175 VDD2.n174 104.615
R127 VDD2.n174 VDD2.n136 104.615
R128 VDD2.n167 VDD2.n136 104.615
R129 VDD2.n167 VDD2.n166 104.615
R130 VDD2.n166 VDD2.n140 104.615
R131 VDD2.n159 VDD2.n140 104.615
R132 VDD2.n159 VDD2.n158 104.615
R133 VDD2.n158 VDD2.n144 104.615
R134 VDD2.n151 VDD2.n144 104.615
R135 VDD2.n151 VDD2.n150 104.615
R136 VDD2.n38 VDD2.n37 104.615
R137 VDD2.n38 VDD2.n31 104.615
R138 VDD2.n45 VDD2.n31 104.615
R139 VDD2.n46 VDD2.n45 104.615
R140 VDD2.n46 VDD2.n27 104.615
R141 VDD2.n53 VDD2.n27 104.615
R142 VDD2.n54 VDD2.n53 104.615
R143 VDD2.n54 VDD2.n23 104.615
R144 VDD2.n61 VDD2.n23 104.615
R145 VDD2.n62 VDD2.n61 104.615
R146 VDD2.n62 VDD2.n19 104.615
R147 VDD2.n69 VDD2.n19 104.615
R148 VDD2.n70 VDD2.n69 104.615
R149 VDD2.n70 VDD2.n15 104.615
R150 VDD2.n78 VDD2.n15 104.615
R151 VDD2.n79 VDD2.n78 104.615
R152 VDD2.n80 VDD2.n79 104.615
R153 VDD2.n80 VDD2.n11 104.615
R154 VDD2.n87 VDD2.n11 104.615
R155 VDD2.n88 VDD2.n87 104.615
R156 VDD2.n88 VDD2.n7 104.615
R157 VDD2.n95 VDD2.n7 104.615
R158 VDD2.n96 VDD2.n95 104.615
R159 VDD2.n96 VDD2.n3 104.615
R160 VDD2.n103 VDD2.n3 104.615
R161 VDD2.n104 VDD2.n103 104.615
R162 VDD2.n110 VDD2.n109 61.0984
R163 VDD2 VDD2.n221 61.0955
R164 VDD2.n150 VDD2.t0 52.3082
R165 VDD2.n37 VDD2.t3 52.3082
R166 VDD2.n110 VDD2.n108 50.8519
R167 VDD2.n220 VDD2.n110 50.3662
R168 VDD2.n220 VDD2.n219 48.6702
R169 VDD2.n149 VDD2.n148 15.6677
R170 VDD2.n36 VDD2.n35 15.6677
R171 VDD2.n125 VDD2.n123 13.1884
R172 VDD2.n81 VDD2.n12 13.1884
R173 VDD2.n197 VDD2.n196 12.8005
R174 VDD2.n193 VDD2.n192 12.8005
R175 VDD2.n152 VDD2.n147 12.8005
R176 VDD2.n39 VDD2.n34 12.8005
R177 VDD2.n82 VDD2.n14 12.8005
R178 VDD2.n86 VDD2.n85 12.8005
R179 VDD2.n200 VDD2.n121 12.0247
R180 VDD2.n189 VDD2.n126 12.0247
R181 VDD2.n153 VDD2.n145 12.0247
R182 VDD2.n40 VDD2.n32 12.0247
R183 VDD2.n77 VDD2.n76 12.0247
R184 VDD2.n89 VDD2.n10 12.0247
R185 VDD2.n201 VDD2.n119 11.249
R186 VDD2.n188 VDD2.n129 11.249
R187 VDD2.n157 VDD2.n156 11.249
R188 VDD2.n44 VDD2.n43 11.249
R189 VDD2.n75 VDD2.n16 11.249
R190 VDD2.n90 VDD2.n8 11.249
R191 VDD2.n205 VDD2.n204 10.4732
R192 VDD2.n185 VDD2.n184 10.4732
R193 VDD2.n160 VDD2.n143 10.4732
R194 VDD2.n47 VDD2.n30 10.4732
R195 VDD2.n72 VDD2.n71 10.4732
R196 VDD2.n94 VDD2.n93 10.4732
R197 VDD2.n208 VDD2.n117 9.69747
R198 VDD2.n181 VDD2.n131 9.69747
R199 VDD2.n161 VDD2.n141 9.69747
R200 VDD2.n48 VDD2.n28 9.69747
R201 VDD2.n68 VDD2.n18 9.69747
R202 VDD2.n97 VDD2.n6 9.69747
R203 VDD2.n219 VDD2.n218 9.45567
R204 VDD2.n108 VDD2.n107 9.45567
R205 VDD2.n135 VDD2.n134 9.3005
R206 VDD2.n178 VDD2.n177 9.3005
R207 VDD2.n180 VDD2.n179 9.3005
R208 VDD2.n131 VDD2.n130 9.3005
R209 VDD2.n186 VDD2.n185 9.3005
R210 VDD2.n188 VDD2.n187 9.3005
R211 VDD2.n126 VDD2.n124 9.3005
R212 VDD2.n194 VDD2.n193 9.3005
R213 VDD2.n218 VDD2.n217 9.3005
R214 VDD2.n113 VDD2.n112 9.3005
R215 VDD2.n212 VDD2.n211 9.3005
R216 VDD2.n210 VDD2.n209 9.3005
R217 VDD2.n117 VDD2.n116 9.3005
R218 VDD2.n204 VDD2.n203 9.3005
R219 VDD2.n202 VDD2.n201 9.3005
R220 VDD2.n121 VDD2.n120 9.3005
R221 VDD2.n196 VDD2.n195 9.3005
R222 VDD2.n172 VDD2.n171 9.3005
R223 VDD2.n170 VDD2.n169 9.3005
R224 VDD2.n139 VDD2.n138 9.3005
R225 VDD2.n164 VDD2.n163 9.3005
R226 VDD2.n162 VDD2.n161 9.3005
R227 VDD2.n143 VDD2.n142 9.3005
R228 VDD2.n156 VDD2.n155 9.3005
R229 VDD2.n154 VDD2.n153 9.3005
R230 VDD2.n147 VDD2.n146 9.3005
R231 VDD2.n107 VDD2.n106 9.3005
R232 VDD2.n101 VDD2.n100 9.3005
R233 VDD2.n99 VDD2.n98 9.3005
R234 VDD2.n6 VDD2.n5 9.3005
R235 VDD2.n93 VDD2.n92 9.3005
R236 VDD2.n91 VDD2.n90 9.3005
R237 VDD2.n10 VDD2.n9 9.3005
R238 VDD2.n85 VDD2.n84 9.3005
R239 VDD2.n57 VDD2.n56 9.3005
R240 VDD2.n26 VDD2.n25 9.3005
R241 VDD2.n51 VDD2.n50 9.3005
R242 VDD2.n49 VDD2.n48 9.3005
R243 VDD2.n30 VDD2.n29 9.3005
R244 VDD2.n43 VDD2.n42 9.3005
R245 VDD2.n41 VDD2.n40 9.3005
R246 VDD2.n34 VDD2.n33 9.3005
R247 VDD2.n59 VDD2.n58 9.3005
R248 VDD2.n22 VDD2.n21 9.3005
R249 VDD2.n65 VDD2.n64 9.3005
R250 VDD2.n67 VDD2.n66 9.3005
R251 VDD2.n18 VDD2.n17 9.3005
R252 VDD2.n73 VDD2.n72 9.3005
R253 VDD2.n75 VDD2.n74 9.3005
R254 VDD2.n76 VDD2.n13 9.3005
R255 VDD2.n83 VDD2.n82 9.3005
R256 VDD2.n2 VDD2.n1 9.3005
R257 VDD2.n209 VDD2.n115 8.92171
R258 VDD2.n180 VDD2.n133 8.92171
R259 VDD2.n165 VDD2.n164 8.92171
R260 VDD2.n52 VDD2.n51 8.92171
R261 VDD2.n67 VDD2.n20 8.92171
R262 VDD2.n98 VDD2.n4 8.92171
R263 VDD2.n213 VDD2.n212 8.14595
R264 VDD2.n177 VDD2.n176 8.14595
R265 VDD2.n168 VDD2.n139 8.14595
R266 VDD2.n55 VDD2.n26 8.14595
R267 VDD2.n64 VDD2.n63 8.14595
R268 VDD2.n102 VDD2.n101 8.14595
R269 VDD2.n219 VDD2.n111 7.3702
R270 VDD2.n216 VDD2.n113 7.3702
R271 VDD2.n173 VDD2.n135 7.3702
R272 VDD2.n169 VDD2.n137 7.3702
R273 VDD2.n56 VDD2.n24 7.3702
R274 VDD2.n60 VDD2.n22 7.3702
R275 VDD2.n105 VDD2.n2 7.3702
R276 VDD2.n108 VDD2.n0 7.3702
R277 VDD2.n217 VDD2.n111 6.59444
R278 VDD2.n217 VDD2.n216 6.59444
R279 VDD2.n173 VDD2.n172 6.59444
R280 VDD2.n172 VDD2.n137 6.59444
R281 VDD2.n59 VDD2.n24 6.59444
R282 VDD2.n60 VDD2.n59 6.59444
R283 VDD2.n106 VDD2.n105 6.59444
R284 VDD2.n106 VDD2.n0 6.59444
R285 VDD2.n213 VDD2.n113 5.81868
R286 VDD2.n176 VDD2.n135 5.81868
R287 VDD2.n169 VDD2.n168 5.81868
R288 VDD2.n56 VDD2.n55 5.81868
R289 VDD2.n63 VDD2.n22 5.81868
R290 VDD2.n102 VDD2.n2 5.81868
R291 VDD2.n212 VDD2.n115 5.04292
R292 VDD2.n177 VDD2.n133 5.04292
R293 VDD2.n165 VDD2.n139 5.04292
R294 VDD2.n52 VDD2.n26 5.04292
R295 VDD2.n64 VDD2.n20 5.04292
R296 VDD2.n101 VDD2.n4 5.04292
R297 VDD2.n148 VDD2.n146 4.38563
R298 VDD2.n35 VDD2.n33 4.38563
R299 VDD2.n209 VDD2.n208 4.26717
R300 VDD2.n181 VDD2.n180 4.26717
R301 VDD2.n164 VDD2.n141 4.26717
R302 VDD2.n51 VDD2.n28 4.26717
R303 VDD2.n68 VDD2.n67 4.26717
R304 VDD2.n98 VDD2.n97 4.26717
R305 VDD2.n205 VDD2.n117 3.49141
R306 VDD2.n184 VDD2.n131 3.49141
R307 VDD2.n161 VDD2.n160 3.49141
R308 VDD2.n48 VDD2.n47 3.49141
R309 VDD2.n71 VDD2.n18 3.49141
R310 VDD2.n94 VDD2.n6 3.49141
R311 VDD2.n204 VDD2.n119 2.71565
R312 VDD2.n185 VDD2.n129 2.71565
R313 VDD2.n157 VDD2.n143 2.71565
R314 VDD2.n44 VDD2.n30 2.71565
R315 VDD2.n72 VDD2.n16 2.71565
R316 VDD2.n93 VDD2.n8 2.71565
R317 VDD2 VDD2.n220 2.29576
R318 VDD2.n201 VDD2.n200 1.93989
R319 VDD2.n189 VDD2.n188 1.93989
R320 VDD2.n156 VDD2.n145 1.93989
R321 VDD2.n43 VDD2.n32 1.93989
R322 VDD2.n77 VDD2.n75 1.93989
R323 VDD2.n90 VDD2.n89 1.93989
R324 VDD2.n197 VDD2.n121 1.16414
R325 VDD2.n192 VDD2.n126 1.16414
R326 VDD2.n153 VDD2.n152 1.16414
R327 VDD2.n40 VDD2.n39 1.16414
R328 VDD2.n76 VDD2.n14 1.16414
R329 VDD2.n86 VDD2.n10 1.16414
R330 VDD2.n221 VDD2.t5 1.00711
R331 VDD2.n221 VDD2.t4 1.00711
R332 VDD2.n109 VDD2.t1 1.00711
R333 VDD2.n109 VDD2.t2 1.00711
R334 VDD2.n196 VDD2.n123 0.388379
R335 VDD2.n193 VDD2.n125 0.388379
R336 VDD2.n149 VDD2.n147 0.388379
R337 VDD2.n36 VDD2.n34 0.388379
R338 VDD2.n82 VDD2.n81 0.388379
R339 VDD2.n85 VDD2.n12 0.388379
R340 VDD2.n218 VDD2.n112 0.155672
R341 VDD2.n211 VDD2.n112 0.155672
R342 VDD2.n211 VDD2.n210 0.155672
R343 VDD2.n210 VDD2.n116 0.155672
R344 VDD2.n203 VDD2.n116 0.155672
R345 VDD2.n203 VDD2.n202 0.155672
R346 VDD2.n202 VDD2.n120 0.155672
R347 VDD2.n195 VDD2.n120 0.155672
R348 VDD2.n195 VDD2.n194 0.155672
R349 VDD2.n194 VDD2.n124 0.155672
R350 VDD2.n187 VDD2.n124 0.155672
R351 VDD2.n187 VDD2.n186 0.155672
R352 VDD2.n186 VDD2.n130 0.155672
R353 VDD2.n179 VDD2.n130 0.155672
R354 VDD2.n179 VDD2.n178 0.155672
R355 VDD2.n178 VDD2.n134 0.155672
R356 VDD2.n171 VDD2.n134 0.155672
R357 VDD2.n171 VDD2.n170 0.155672
R358 VDD2.n170 VDD2.n138 0.155672
R359 VDD2.n163 VDD2.n138 0.155672
R360 VDD2.n163 VDD2.n162 0.155672
R361 VDD2.n162 VDD2.n142 0.155672
R362 VDD2.n155 VDD2.n142 0.155672
R363 VDD2.n155 VDD2.n154 0.155672
R364 VDD2.n154 VDD2.n146 0.155672
R365 VDD2.n41 VDD2.n33 0.155672
R366 VDD2.n42 VDD2.n41 0.155672
R367 VDD2.n42 VDD2.n29 0.155672
R368 VDD2.n49 VDD2.n29 0.155672
R369 VDD2.n50 VDD2.n49 0.155672
R370 VDD2.n50 VDD2.n25 0.155672
R371 VDD2.n57 VDD2.n25 0.155672
R372 VDD2.n58 VDD2.n57 0.155672
R373 VDD2.n58 VDD2.n21 0.155672
R374 VDD2.n65 VDD2.n21 0.155672
R375 VDD2.n66 VDD2.n65 0.155672
R376 VDD2.n66 VDD2.n17 0.155672
R377 VDD2.n73 VDD2.n17 0.155672
R378 VDD2.n74 VDD2.n73 0.155672
R379 VDD2.n74 VDD2.n13 0.155672
R380 VDD2.n83 VDD2.n13 0.155672
R381 VDD2.n84 VDD2.n83 0.155672
R382 VDD2.n84 VDD2.n9 0.155672
R383 VDD2.n91 VDD2.n9 0.155672
R384 VDD2.n92 VDD2.n91 0.155672
R385 VDD2.n92 VDD2.n5 0.155672
R386 VDD2.n99 VDD2.n5 0.155672
R387 VDD2.n100 VDD2.n99 0.155672
R388 VDD2.n100 VDD2.n1 0.155672
R389 VDD2.n107 VDD2.n1 0.155672
R390 VTAIL.n442 VTAIL.n338 289.615
R391 VTAIL.n106 VTAIL.n2 289.615
R392 VTAIL.n332 VTAIL.n228 289.615
R393 VTAIL.n220 VTAIL.n116 289.615
R394 VTAIL.n375 VTAIL.n374 185
R395 VTAIL.n377 VTAIL.n376 185
R396 VTAIL.n370 VTAIL.n369 185
R397 VTAIL.n383 VTAIL.n382 185
R398 VTAIL.n385 VTAIL.n384 185
R399 VTAIL.n366 VTAIL.n365 185
R400 VTAIL.n391 VTAIL.n390 185
R401 VTAIL.n393 VTAIL.n392 185
R402 VTAIL.n362 VTAIL.n361 185
R403 VTAIL.n399 VTAIL.n398 185
R404 VTAIL.n401 VTAIL.n400 185
R405 VTAIL.n358 VTAIL.n357 185
R406 VTAIL.n407 VTAIL.n406 185
R407 VTAIL.n409 VTAIL.n408 185
R408 VTAIL.n354 VTAIL.n353 185
R409 VTAIL.n416 VTAIL.n415 185
R410 VTAIL.n417 VTAIL.n352 185
R411 VTAIL.n419 VTAIL.n418 185
R412 VTAIL.n350 VTAIL.n349 185
R413 VTAIL.n425 VTAIL.n424 185
R414 VTAIL.n427 VTAIL.n426 185
R415 VTAIL.n346 VTAIL.n345 185
R416 VTAIL.n433 VTAIL.n432 185
R417 VTAIL.n435 VTAIL.n434 185
R418 VTAIL.n342 VTAIL.n341 185
R419 VTAIL.n441 VTAIL.n440 185
R420 VTAIL.n443 VTAIL.n442 185
R421 VTAIL.n39 VTAIL.n38 185
R422 VTAIL.n41 VTAIL.n40 185
R423 VTAIL.n34 VTAIL.n33 185
R424 VTAIL.n47 VTAIL.n46 185
R425 VTAIL.n49 VTAIL.n48 185
R426 VTAIL.n30 VTAIL.n29 185
R427 VTAIL.n55 VTAIL.n54 185
R428 VTAIL.n57 VTAIL.n56 185
R429 VTAIL.n26 VTAIL.n25 185
R430 VTAIL.n63 VTAIL.n62 185
R431 VTAIL.n65 VTAIL.n64 185
R432 VTAIL.n22 VTAIL.n21 185
R433 VTAIL.n71 VTAIL.n70 185
R434 VTAIL.n73 VTAIL.n72 185
R435 VTAIL.n18 VTAIL.n17 185
R436 VTAIL.n80 VTAIL.n79 185
R437 VTAIL.n81 VTAIL.n16 185
R438 VTAIL.n83 VTAIL.n82 185
R439 VTAIL.n14 VTAIL.n13 185
R440 VTAIL.n89 VTAIL.n88 185
R441 VTAIL.n91 VTAIL.n90 185
R442 VTAIL.n10 VTAIL.n9 185
R443 VTAIL.n97 VTAIL.n96 185
R444 VTAIL.n99 VTAIL.n98 185
R445 VTAIL.n6 VTAIL.n5 185
R446 VTAIL.n105 VTAIL.n104 185
R447 VTAIL.n107 VTAIL.n106 185
R448 VTAIL.n333 VTAIL.n332 185
R449 VTAIL.n331 VTAIL.n330 185
R450 VTAIL.n232 VTAIL.n231 185
R451 VTAIL.n325 VTAIL.n324 185
R452 VTAIL.n323 VTAIL.n322 185
R453 VTAIL.n236 VTAIL.n235 185
R454 VTAIL.n317 VTAIL.n316 185
R455 VTAIL.n315 VTAIL.n314 185
R456 VTAIL.n240 VTAIL.n239 185
R457 VTAIL.n244 VTAIL.n242 185
R458 VTAIL.n309 VTAIL.n308 185
R459 VTAIL.n307 VTAIL.n306 185
R460 VTAIL.n246 VTAIL.n245 185
R461 VTAIL.n301 VTAIL.n300 185
R462 VTAIL.n299 VTAIL.n298 185
R463 VTAIL.n250 VTAIL.n249 185
R464 VTAIL.n293 VTAIL.n292 185
R465 VTAIL.n291 VTAIL.n290 185
R466 VTAIL.n254 VTAIL.n253 185
R467 VTAIL.n285 VTAIL.n284 185
R468 VTAIL.n283 VTAIL.n282 185
R469 VTAIL.n258 VTAIL.n257 185
R470 VTAIL.n277 VTAIL.n276 185
R471 VTAIL.n275 VTAIL.n274 185
R472 VTAIL.n262 VTAIL.n261 185
R473 VTAIL.n269 VTAIL.n268 185
R474 VTAIL.n267 VTAIL.n266 185
R475 VTAIL.n221 VTAIL.n220 185
R476 VTAIL.n219 VTAIL.n218 185
R477 VTAIL.n120 VTAIL.n119 185
R478 VTAIL.n213 VTAIL.n212 185
R479 VTAIL.n211 VTAIL.n210 185
R480 VTAIL.n124 VTAIL.n123 185
R481 VTAIL.n205 VTAIL.n204 185
R482 VTAIL.n203 VTAIL.n202 185
R483 VTAIL.n128 VTAIL.n127 185
R484 VTAIL.n132 VTAIL.n130 185
R485 VTAIL.n197 VTAIL.n196 185
R486 VTAIL.n195 VTAIL.n194 185
R487 VTAIL.n134 VTAIL.n133 185
R488 VTAIL.n189 VTAIL.n188 185
R489 VTAIL.n187 VTAIL.n186 185
R490 VTAIL.n138 VTAIL.n137 185
R491 VTAIL.n181 VTAIL.n180 185
R492 VTAIL.n179 VTAIL.n178 185
R493 VTAIL.n142 VTAIL.n141 185
R494 VTAIL.n173 VTAIL.n172 185
R495 VTAIL.n171 VTAIL.n170 185
R496 VTAIL.n146 VTAIL.n145 185
R497 VTAIL.n165 VTAIL.n164 185
R498 VTAIL.n163 VTAIL.n162 185
R499 VTAIL.n150 VTAIL.n149 185
R500 VTAIL.n157 VTAIL.n156 185
R501 VTAIL.n155 VTAIL.n154 185
R502 VTAIL.n373 VTAIL.t6 147.659
R503 VTAIL.n37 VTAIL.t4 147.659
R504 VTAIL.n265 VTAIL.t5 147.659
R505 VTAIL.n153 VTAIL.t8 147.659
R506 VTAIL.n376 VTAIL.n375 104.615
R507 VTAIL.n376 VTAIL.n369 104.615
R508 VTAIL.n383 VTAIL.n369 104.615
R509 VTAIL.n384 VTAIL.n383 104.615
R510 VTAIL.n384 VTAIL.n365 104.615
R511 VTAIL.n391 VTAIL.n365 104.615
R512 VTAIL.n392 VTAIL.n391 104.615
R513 VTAIL.n392 VTAIL.n361 104.615
R514 VTAIL.n399 VTAIL.n361 104.615
R515 VTAIL.n400 VTAIL.n399 104.615
R516 VTAIL.n400 VTAIL.n357 104.615
R517 VTAIL.n407 VTAIL.n357 104.615
R518 VTAIL.n408 VTAIL.n407 104.615
R519 VTAIL.n408 VTAIL.n353 104.615
R520 VTAIL.n416 VTAIL.n353 104.615
R521 VTAIL.n417 VTAIL.n416 104.615
R522 VTAIL.n418 VTAIL.n417 104.615
R523 VTAIL.n418 VTAIL.n349 104.615
R524 VTAIL.n425 VTAIL.n349 104.615
R525 VTAIL.n426 VTAIL.n425 104.615
R526 VTAIL.n426 VTAIL.n345 104.615
R527 VTAIL.n433 VTAIL.n345 104.615
R528 VTAIL.n434 VTAIL.n433 104.615
R529 VTAIL.n434 VTAIL.n341 104.615
R530 VTAIL.n441 VTAIL.n341 104.615
R531 VTAIL.n442 VTAIL.n441 104.615
R532 VTAIL.n40 VTAIL.n39 104.615
R533 VTAIL.n40 VTAIL.n33 104.615
R534 VTAIL.n47 VTAIL.n33 104.615
R535 VTAIL.n48 VTAIL.n47 104.615
R536 VTAIL.n48 VTAIL.n29 104.615
R537 VTAIL.n55 VTAIL.n29 104.615
R538 VTAIL.n56 VTAIL.n55 104.615
R539 VTAIL.n56 VTAIL.n25 104.615
R540 VTAIL.n63 VTAIL.n25 104.615
R541 VTAIL.n64 VTAIL.n63 104.615
R542 VTAIL.n64 VTAIL.n21 104.615
R543 VTAIL.n71 VTAIL.n21 104.615
R544 VTAIL.n72 VTAIL.n71 104.615
R545 VTAIL.n72 VTAIL.n17 104.615
R546 VTAIL.n80 VTAIL.n17 104.615
R547 VTAIL.n81 VTAIL.n80 104.615
R548 VTAIL.n82 VTAIL.n81 104.615
R549 VTAIL.n82 VTAIL.n13 104.615
R550 VTAIL.n89 VTAIL.n13 104.615
R551 VTAIL.n90 VTAIL.n89 104.615
R552 VTAIL.n90 VTAIL.n9 104.615
R553 VTAIL.n97 VTAIL.n9 104.615
R554 VTAIL.n98 VTAIL.n97 104.615
R555 VTAIL.n98 VTAIL.n5 104.615
R556 VTAIL.n105 VTAIL.n5 104.615
R557 VTAIL.n106 VTAIL.n105 104.615
R558 VTAIL.n332 VTAIL.n331 104.615
R559 VTAIL.n331 VTAIL.n231 104.615
R560 VTAIL.n324 VTAIL.n231 104.615
R561 VTAIL.n324 VTAIL.n323 104.615
R562 VTAIL.n323 VTAIL.n235 104.615
R563 VTAIL.n316 VTAIL.n235 104.615
R564 VTAIL.n316 VTAIL.n315 104.615
R565 VTAIL.n315 VTAIL.n239 104.615
R566 VTAIL.n244 VTAIL.n239 104.615
R567 VTAIL.n308 VTAIL.n244 104.615
R568 VTAIL.n308 VTAIL.n307 104.615
R569 VTAIL.n307 VTAIL.n245 104.615
R570 VTAIL.n300 VTAIL.n245 104.615
R571 VTAIL.n300 VTAIL.n299 104.615
R572 VTAIL.n299 VTAIL.n249 104.615
R573 VTAIL.n292 VTAIL.n249 104.615
R574 VTAIL.n292 VTAIL.n291 104.615
R575 VTAIL.n291 VTAIL.n253 104.615
R576 VTAIL.n284 VTAIL.n253 104.615
R577 VTAIL.n284 VTAIL.n283 104.615
R578 VTAIL.n283 VTAIL.n257 104.615
R579 VTAIL.n276 VTAIL.n257 104.615
R580 VTAIL.n276 VTAIL.n275 104.615
R581 VTAIL.n275 VTAIL.n261 104.615
R582 VTAIL.n268 VTAIL.n261 104.615
R583 VTAIL.n268 VTAIL.n267 104.615
R584 VTAIL.n220 VTAIL.n219 104.615
R585 VTAIL.n219 VTAIL.n119 104.615
R586 VTAIL.n212 VTAIL.n119 104.615
R587 VTAIL.n212 VTAIL.n211 104.615
R588 VTAIL.n211 VTAIL.n123 104.615
R589 VTAIL.n204 VTAIL.n123 104.615
R590 VTAIL.n204 VTAIL.n203 104.615
R591 VTAIL.n203 VTAIL.n127 104.615
R592 VTAIL.n132 VTAIL.n127 104.615
R593 VTAIL.n196 VTAIL.n132 104.615
R594 VTAIL.n196 VTAIL.n195 104.615
R595 VTAIL.n195 VTAIL.n133 104.615
R596 VTAIL.n188 VTAIL.n133 104.615
R597 VTAIL.n188 VTAIL.n187 104.615
R598 VTAIL.n187 VTAIL.n137 104.615
R599 VTAIL.n180 VTAIL.n137 104.615
R600 VTAIL.n180 VTAIL.n179 104.615
R601 VTAIL.n179 VTAIL.n141 104.615
R602 VTAIL.n172 VTAIL.n141 104.615
R603 VTAIL.n172 VTAIL.n171 104.615
R604 VTAIL.n171 VTAIL.n145 104.615
R605 VTAIL.n164 VTAIL.n145 104.615
R606 VTAIL.n164 VTAIL.n163 104.615
R607 VTAIL.n163 VTAIL.n149 104.615
R608 VTAIL.n156 VTAIL.n149 104.615
R609 VTAIL.n156 VTAIL.n155 104.615
R610 VTAIL.n375 VTAIL.t6 52.3082
R611 VTAIL.n39 VTAIL.t4 52.3082
R612 VTAIL.n267 VTAIL.t5 52.3082
R613 VTAIL.n155 VTAIL.t8 52.3082
R614 VTAIL.n227 VTAIL.n226 43.7294
R615 VTAIL.n115 VTAIL.n114 43.7294
R616 VTAIL.n1 VTAIL.n0 43.7292
R617 VTAIL.n113 VTAIL.n112 43.7292
R618 VTAIL.n115 VTAIL.n113 35.2893
R619 VTAIL.n447 VTAIL.n337 32.3065
R620 VTAIL.n447 VTAIL.n446 31.9914
R621 VTAIL.n111 VTAIL.n110 31.9914
R622 VTAIL.n337 VTAIL.n336 31.9914
R623 VTAIL.n225 VTAIL.n224 31.9914
R624 VTAIL.n374 VTAIL.n373 15.6677
R625 VTAIL.n38 VTAIL.n37 15.6677
R626 VTAIL.n266 VTAIL.n265 15.6677
R627 VTAIL.n154 VTAIL.n153 15.6677
R628 VTAIL.n419 VTAIL.n350 13.1884
R629 VTAIL.n83 VTAIL.n14 13.1884
R630 VTAIL.n242 VTAIL.n240 13.1884
R631 VTAIL.n130 VTAIL.n128 13.1884
R632 VTAIL.n377 VTAIL.n372 12.8005
R633 VTAIL.n420 VTAIL.n352 12.8005
R634 VTAIL.n424 VTAIL.n423 12.8005
R635 VTAIL.n41 VTAIL.n36 12.8005
R636 VTAIL.n84 VTAIL.n16 12.8005
R637 VTAIL.n88 VTAIL.n87 12.8005
R638 VTAIL.n314 VTAIL.n313 12.8005
R639 VTAIL.n310 VTAIL.n309 12.8005
R640 VTAIL.n269 VTAIL.n264 12.8005
R641 VTAIL.n202 VTAIL.n201 12.8005
R642 VTAIL.n198 VTAIL.n197 12.8005
R643 VTAIL.n157 VTAIL.n152 12.8005
R644 VTAIL.n378 VTAIL.n370 12.0247
R645 VTAIL.n415 VTAIL.n414 12.0247
R646 VTAIL.n427 VTAIL.n348 12.0247
R647 VTAIL.n42 VTAIL.n34 12.0247
R648 VTAIL.n79 VTAIL.n78 12.0247
R649 VTAIL.n91 VTAIL.n12 12.0247
R650 VTAIL.n317 VTAIL.n238 12.0247
R651 VTAIL.n306 VTAIL.n243 12.0247
R652 VTAIL.n270 VTAIL.n262 12.0247
R653 VTAIL.n205 VTAIL.n126 12.0247
R654 VTAIL.n194 VTAIL.n131 12.0247
R655 VTAIL.n158 VTAIL.n150 12.0247
R656 VTAIL.n382 VTAIL.n381 11.249
R657 VTAIL.n413 VTAIL.n354 11.249
R658 VTAIL.n428 VTAIL.n346 11.249
R659 VTAIL.n46 VTAIL.n45 11.249
R660 VTAIL.n77 VTAIL.n18 11.249
R661 VTAIL.n92 VTAIL.n10 11.249
R662 VTAIL.n318 VTAIL.n236 11.249
R663 VTAIL.n305 VTAIL.n246 11.249
R664 VTAIL.n274 VTAIL.n273 11.249
R665 VTAIL.n206 VTAIL.n124 11.249
R666 VTAIL.n193 VTAIL.n134 11.249
R667 VTAIL.n162 VTAIL.n161 11.249
R668 VTAIL.n385 VTAIL.n368 10.4732
R669 VTAIL.n410 VTAIL.n409 10.4732
R670 VTAIL.n432 VTAIL.n431 10.4732
R671 VTAIL.n49 VTAIL.n32 10.4732
R672 VTAIL.n74 VTAIL.n73 10.4732
R673 VTAIL.n96 VTAIL.n95 10.4732
R674 VTAIL.n322 VTAIL.n321 10.4732
R675 VTAIL.n302 VTAIL.n301 10.4732
R676 VTAIL.n277 VTAIL.n260 10.4732
R677 VTAIL.n210 VTAIL.n209 10.4732
R678 VTAIL.n190 VTAIL.n189 10.4732
R679 VTAIL.n165 VTAIL.n148 10.4732
R680 VTAIL.n386 VTAIL.n366 9.69747
R681 VTAIL.n406 VTAIL.n356 9.69747
R682 VTAIL.n435 VTAIL.n344 9.69747
R683 VTAIL.n50 VTAIL.n30 9.69747
R684 VTAIL.n70 VTAIL.n20 9.69747
R685 VTAIL.n99 VTAIL.n8 9.69747
R686 VTAIL.n325 VTAIL.n234 9.69747
R687 VTAIL.n298 VTAIL.n248 9.69747
R688 VTAIL.n278 VTAIL.n258 9.69747
R689 VTAIL.n213 VTAIL.n122 9.69747
R690 VTAIL.n186 VTAIL.n136 9.69747
R691 VTAIL.n166 VTAIL.n146 9.69747
R692 VTAIL.n446 VTAIL.n445 9.45567
R693 VTAIL.n110 VTAIL.n109 9.45567
R694 VTAIL.n336 VTAIL.n335 9.45567
R695 VTAIL.n224 VTAIL.n223 9.45567
R696 VTAIL.n445 VTAIL.n444 9.3005
R697 VTAIL.n439 VTAIL.n438 9.3005
R698 VTAIL.n437 VTAIL.n436 9.3005
R699 VTAIL.n344 VTAIL.n343 9.3005
R700 VTAIL.n431 VTAIL.n430 9.3005
R701 VTAIL.n429 VTAIL.n428 9.3005
R702 VTAIL.n348 VTAIL.n347 9.3005
R703 VTAIL.n423 VTAIL.n422 9.3005
R704 VTAIL.n395 VTAIL.n394 9.3005
R705 VTAIL.n364 VTAIL.n363 9.3005
R706 VTAIL.n389 VTAIL.n388 9.3005
R707 VTAIL.n387 VTAIL.n386 9.3005
R708 VTAIL.n368 VTAIL.n367 9.3005
R709 VTAIL.n381 VTAIL.n380 9.3005
R710 VTAIL.n379 VTAIL.n378 9.3005
R711 VTAIL.n372 VTAIL.n371 9.3005
R712 VTAIL.n397 VTAIL.n396 9.3005
R713 VTAIL.n360 VTAIL.n359 9.3005
R714 VTAIL.n403 VTAIL.n402 9.3005
R715 VTAIL.n405 VTAIL.n404 9.3005
R716 VTAIL.n356 VTAIL.n355 9.3005
R717 VTAIL.n411 VTAIL.n410 9.3005
R718 VTAIL.n413 VTAIL.n412 9.3005
R719 VTAIL.n414 VTAIL.n351 9.3005
R720 VTAIL.n421 VTAIL.n420 9.3005
R721 VTAIL.n340 VTAIL.n339 9.3005
R722 VTAIL.n109 VTAIL.n108 9.3005
R723 VTAIL.n103 VTAIL.n102 9.3005
R724 VTAIL.n101 VTAIL.n100 9.3005
R725 VTAIL.n8 VTAIL.n7 9.3005
R726 VTAIL.n95 VTAIL.n94 9.3005
R727 VTAIL.n93 VTAIL.n92 9.3005
R728 VTAIL.n12 VTAIL.n11 9.3005
R729 VTAIL.n87 VTAIL.n86 9.3005
R730 VTAIL.n59 VTAIL.n58 9.3005
R731 VTAIL.n28 VTAIL.n27 9.3005
R732 VTAIL.n53 VTAIL.n52 9.3005
R733 VTAIL.n51 VTAIL.n50 9.3005
R734 VTAIL.n32 VTAIL.n31 9.3005
R735 VTAIL.n45 VTAIL.n44 9.3005
R736 VTAIL.n43 VTAIL.n42 9.3005
R737 VTAIL.n36 VTAIL.n35 9.3005
R738 VTAIL.n61 VTAIL.n60 9.3005
R739 VTAIL.n24 VTAIL.n23 9.3005
R740 VTAIL.n67 VTAIL.n66 9.3005
R741 VTAIL.n69 VTAIL.n68 9.3005
R742 VTAIL.n20 VTAIL.n19 9.3005
R743 VTAIL.n75 VTAIL.n74 9.3005
R744 VTAIL.n77 VTAIL.n76 9.3005
R745 VTAIL.n78 VTAIL.n15 9.3005
R746 VTAIL.n85 VTAIL.n84 9.3005
R747 VTAIL.n4 VTAIL.n3 9.3005
R748 VTAIL.n252 VTAIL.n251 9.3005
R749 VTAIL.n295 VTAIL.n294 9.3005
R750 VTAIL.n297 VTAIL.n296 9.3005
R751 VTAIL.n248 VTAIL.n247 9.3005
R752 VTAIL.n303 VTAIL.n302 9.3005
R753 VTAIL.n305 VTAIL.n304 9.3005
R754 VTAIL.n243 VTAIL.n241 9.3005
R755 VTAIL.n311 VTAIL.n310 9.3005
R756 VTAIL.n335 VTAIL.n334 9.3005
R757 VTAIL.n230 VTAIL.n229 9.3005
R758 VTAIL.n329 VTAIL.n328 9.3005
R759 VTAIL.n327 VTAIL.n326 9.3005
R760 VTAIL.n234 VTAIL.n233 9.3005
R761 VTAIL.n321 VTAIL.n320 9.3005
R762 VTAIL.n319 VTAIL.n318 9.3005
R763 VTAIL.n238 VTAIL.n237 9.3005
R764 VTAIL.n313 VTAIL.n312 9.3005
R765 VTAIL.n289 VTAIL.n288 9.3005
R766 VTAIL.n287 VTAIL.n286 9.3005
R767 VTAIL.n256 VTAIL.n255 9.3005
R768 VTAIL.n281 VTAIL.n280 9.3005
R769 VTAIL.n279 VTAIL.n278 9.3005
R770 VTAIL.n260 VTAIL.n259 9.3005
R771 VTAIL.n273 VTAIL.n272 9.3005
R772 VTAIL.n271 VTAIL.n270 9.3005
R773 VTAIL.n264 VTAIL.n263 9.3005
R774 VTAIL.n140 VTAIL.n139 9.3005
R775 VTAIL.n183 VTAIL.n182 9.3005
R776 VTAIL.n185 VTAIL.n184 9.3005
R777 VTAIL.n136 VTAIL.n135 9.3005
R778 VTAIL.n191 VTAIL.n190 9.3005
R779 VTAIL.n193 VTAIL.n192 9.3005
R780 VTAIL.n131 VTAIL.n129 9.3005
R781 VTAIL.n199 VTAIL.n198 9.3005
R782 VTAIL.n223 VTAIL.n222 9.3005
R783 VTAIL.n118 VTAIL.n117 9.3005
R784 VTAIL.n217 VTAIL.n216 9.3005
R785 VTAIL.n215 VTAIL.n214 9.3005
R786 VTAIL.n122 VTAIL.n121 9.3005
R787 VTAIL.n209 VTAIL.n208 9.3005
R788 VTAIL.n207 VTAIL.n206 9.3005
R789 VTAIL.n126 VTAIL.n125 9.3005
R790 VTAIL.n201 VTAIL.n200 9.3005
R791 VTAIL.n177 VTAIL.n176 9.3005
R792 VTAIL.n175 VTAIL.n174 9.3005
R793 VTAIL.n144 VTAIL.n143 9.3005
R794 VTAIL.n169 VTAIL.n168 9.3005
R795 VTAIL.n167 VTAIL.n166 9.3005
R796 VTAIL.n148 VTAIL.n147 9.3005
R797 VTAIL.n161 VTAIL.n160 9.3005
R798 VTAIL.n159 VTAIL.n158 9.3005
R799 VTAIL.n152 VTAIL.n151 9.3005
R800 VTAIL.n390 VTAIL.n389 8.92171
R801 VTAIL.n405 VTAIL.n358 8.92171
R802 VTAIL.n436 VTAIL.n342 8.92171
R803 VTAIL.n54 VTAIL.n53 8.92171
R804 VTAIL.n69 VTAIL.n22 8.92171
R805 VTAIL.n100 VTAIL.n6 8.92171
R806 VTAIL.n326 VTAIL.n232 8.92171
R807 VTAIL.n297 VTAIL.n250 8.92171
R808 VTAIL.n282 VTAIL.n281 8.92171
R809 VTAIL.n214 VTAIL.n120 8.92171
R810 VTAIL.n185 VTAIL.n138 8.92171
R811 VTAIL.n170 VTAIL.n169 8.92171
R812 VTAIL.n393 VTAIL.n364 8.14595
R813 VTAIL.n402 VTAIL.n401 8.14595
R814 VTAIL.n440 VTAIL.n439 8.14595
R815 VTAIL.n57 VTAIL.n28 8.14595
R816 VTAIL.n66 VTAIL.n65 8.14595
R817 VTAIL.n104 VTAIL.n103 8.14595
R818 VTAIL.n330 VTAIL.n329 8.14595
R819 VTAIL.n294 VTAIL.n293 8.14595
R820 VTAIL.n285 VTAIL.n256 8.14595
R821 VTAIL.n218 VTAIL.n217 8.14595
R822 VTAIL.n182 VTAIL.n181 8.14595
R823 VTAIL.n173 VTAIL.n144 8.14595
R824 VTAIL.n394 VTAIL.n362 7.3702
R825 VTAIL.n398 VTAIL.n360 7.3702
R826 VTAIL.n443 VTAIL.n340 7.3702
R827 VTAIL.n446 VTAIL.n338 7.3702
R828 VTAIL.n58 VTAIL.n26 7.3702
R829 VTAIL.n62 VTAIL.n24 7.3702
R830 VTAIL.n107 VTAIL.n4 7.3702
R831 VTAIL.n110 VTAIL.n2 7.3702
R832 VTAIL.n336 VTAIL.n228 7.3702
R833 VTAIL.n333 VTAIL.n230 7.3702
R834 VTAIL.n290 VTAIL.n252 7.3702
R835 VTAIL.n286 VTAIL.n254 7.3702
R836 VTAIL.n224 VTAIL.n116 7.3702
R837 VTAIL.n221 VTAIL.n118 7.3702
R838 VTAIL.n178 VTAIL.n140 7.3702
R839 VTAIL.n174 VTAIL.n142 7.3702
R840 VTAIL.n397 VTAIL.n362 6.59444
R841 VTAIL.n398 VTAIL.n397 6.59444
R842 VTAIL.n444 VTAIL.n443 6.59444
R843 VTAIL.n444 VTAIL.n338 6.59444
R844 VTAIL.n61 VTAIL.n26 6.59444
R845 VTAIL.n62 VTAIL.n61 6.59444
R846 VTAIL.n108 VTAIL.n107 6.59444
R847 VTAIL.n108 VTAIL.n2 6.59444
R848 VTAIL.n334 VTAIL.n228 6.59444
R849 VTAIL.n334 VTAIL.n333 6.59444
R850 VTAIL.n290 VTAIL.n289 6.59444
R851 VTAIL.n289 VTAIL.n254 6.59444
R852 VTAIL.n222 VTAIL.n116 6.59444
R853 VTAIL.n222 VTAIL.n221 6.59444
R854 VTAIL.n178 VTAIL.n177 6.59444
R855 VTAIL.n177 VTAIL.n142 6.59444
R856 VTAIL.n394 VTAIL.n393 5.81868
R857 VTAIL.n401 VTAIL.n360 5.81868
R858 VTAIL.n440 VTAIL.n340 5.81868
R859 VTAIL.n58 VTAIL.n57 5.81868
R860 VTAIL.n65 VTAIL.n24 5.81868
R861 VTAIL.n104 VTAIL.n4 5.81868
R862 VTAIL.n330 VTAIL.n230 5.81868
R863 VTAIL.n293 VTAIL.n252 5.81868
R864 VTAIL.n286 VTAIL.n285 5.81868
R865 VTAIL.n218 VTAIL.n118 5.81868
R866 VTAIL.n181 VTAIL.n140 5.81868
R867 VTAIL.n174 VTAIL.n173 5.81868
R868 VTAIL.n390 VTAIL.n364 5.04292
R869 VTAIL.n402 VTAIL.n358 5.04292
R870 VTAIL.n439 VTAIL.n342 5.04292
R871 VTAIL.n54 VTAIL.n28 5.04292
R872 VTAIL.n66 VTAIL.n22 5.04292
R873 VTAIL.n103 VTAIL.n6 5.04292
R874 VTAIL.n329 VTAIL.n232 5.04292
R875 VTAIL.n294 VTAIL.n250 5.04292
R876 VTAIL.n282 VTAIL.n256 5.04292
R877 VTAIL.n217 VTAIL.n120 5.04292
R878 VTAIL.n182 VTAIL.n138 5.04292
R879 VTAIL.n170 VTAIL.n144 5.04292
R880 VTAIL.n373 VTAIL.n371 4.38563
R881 VTAIL.n37 VTAIL.n35 4.38563
R882 VTAIL.n265 VTAIL.n263 4.38563
R883 VTAIL.n153 VTAIL.n151 4.38563
R884 VTAIL.n389 VTAIL.n366 4.26717
R885 VTAIL.n406 VTAIL.n405 4.26717
R886 VTAIL.n436 VTAIL.n435 4.26717
R887 VTAIL.n53 VTAIL.n30 4.26717
R888 VTAIL.n70 VTAIL.n69 4.26717
R889 VTAIL.n100 VTAIL.n99 4.26717
R890 VTAIL.n326 VTAIL.n325 4.26717
R891 VTAIL.n298 VTAIL.n297 4.26717
R892 VTAIL.n281 VTAIL.n258 4.26717
R893 VTAIL.n214 VTAIL.n213 4.26717
R894 VTAIL.n186 VTAIL.n185 4.26717
R895 VTAIL.n169 VTAIL.n146 4.26717
R896 VTAIL.n386 VTAIL.n385 3.49141
R897 VTAIL.n409 VTAIL.n356 3.49141
R898 VTAIL.n432 VTAIL.n344 3.49141
R899 VTAIL.n50 VTAIL.n49 3.49141
R900 VTAIL.n73 VTAIL.n20 3.49141
R901 VTAIL.n96 VTAIL.n8 3.49141
R902 VTAIL.n322 VTAIL.n234 3.49141
R903 VTAIL.n301 VTAIL.n248 3.49141
R904 VTAIL.n278 VTAIL.n277 3.49141
R905 VTAIL.n210 VTAIL.n122 3.49141
R906 VTAIL.n189 VTAIL.n136 3.49141
R907 VTAIL.n166 VTAIL.n165 3.49141
R908 VTAIL.n225 VTAIL.n115 2.98326
R909 VTAIL.n337 VTAIL.n227 2.98326
R910 VTAIL.n113 VTAIL.n111 2.98326
R911 VTAIL.n382 VTAIL.n368 2.71565
R912 VTAIL.n410 VTAIL.n354 2.71565
R913 VTAIL.n431 VTAIL.n346 2.71565
R914 VTAIL.n46 VTAIL.n32 2.71565
R915 VTAIL.n74 VTAIL.n18 2.71565
R916 VTAIL.n95 VTAIL.n10 2.71565
R917 VTAIL.n321 VTAIL.n236 2.71565
R918 VTAIL.n302 VTAIL.n246 2.71565
R919 VTAIL.n274 VTAIL.n260 2.71565
R920 VTAIL.n209 VTAIL.n124 2.71565
R921 VTAIL.n190 VTAIL.n134 2.71565
R922 VTAIL.n162 VTAIL.n148 2.71565
R923 VTAIL VTAIL.n447 2.17938
R924 VTAIL.n227 VTAIL.n225 1.96171
R925 VTAIL.n111 VTAIL.n1 1.96171
R926 VTAIL.n381 VTAIL.n370 1.93989
R927 VTAIL.n415 VTAIL.n413 1.93989
R928 VTAIL.n428 VTAIL.n427 1.93989
R929 VTAIL.n45 VTAIL.n34 1.93989
R930 VTAIL.n79 VTAIL.n77 1.93989
R931 VTAIL.n92 VTAIL.n91 1.93989
R932 VTAIL.n318 VTAIL.n317 1.93989
R933 VTAIL.n306 VTAIL.n305 1.93989
R934 VTAIL.n273 VTAIL.n262 1.93989
R935 VTAIL.n206 VTAIL.n205 1.93989
R936 VTAIL.n194 VTAIL.n193 1.93989
R937 VTAIL.n161 VTAIL.n150 1.93989
R938 VTAIL.n378 VTAIL.n377 1.16414
R939 VTAIL.n414 VTAIL.n352 1.16414
R940 VTAIL.n424 VTAIL.n348 1.16414
R941 VTAIL.n42 VTAIL.n41 1.16414
R942 VTAIL.n78 VTAIL.n16 1.16414
R943 VTAIL.n88 VTAIL.n12 1.16414
R944 VTAIL.n314 VTAIL.n238 1.16414
R945 VTAIL.n309 VTAIL.n243 1.16414
R946 VTAIL.n270 VTAIL.n269 1.16414
R947 VTAIL.n202 VTAIL.n126 1.16414
R948 VTAIL.n197 VTAIL.n131 1.16414
R949 VTAIL.n158 VTAIL.n157 1.16414
R950 VTAIL.n0 VTAIL.t9 1.00711
R951 VTAIL.n0 VTAIL.t10 1.00711
R952 VTAIL.n112 VTAIL.t2 1.00711
R953 VTAIL.n112 VTAIL.t0 1.00711
R954 VTAIL.n226 VTAIL.t3 1.00711
R955 VTAIL.n226 VTAIL.t1 1.00711
R956 VTAIL.n114 VTAIL.t7 1.00711
R957 VTAIL.n114 VTAIL.t11 1.00711
R958 VTAIL VTAIL.n1 0.804379
R959 VTAIL.n374 VTAIL.n372 0.388379
R960 VTAIL.n420 VTAIL.n419 0.388379
R961 VTAIL.n423 VTAIL.n350 0.388379
R962 VTAIL.n38 VTAIL.n36 0.388379
R963 VTAIL.n84 VTAIL.n83 0.388379
R964 VTAIL.n87 VTAIL.n14 0.388379
R965 VTAIL.n313 VTAIL.n240 0.388379
R966 VTAIL.n310 VTAIL.n242 0.388379
R967 VTAIL.n266 VTAIL.n264 0.388379
R968 VTAIL.n201 VTAIL.n128 0.388379
R969 VTAIL.n198 VTAIL.n130 0.388379
R970 VTAIL.n154 VTAIL.n152 0.388379
R971 VTAIL.n379 VTAIL.n371 0.155672
R972 VTAIL.n380 VTAIL.n379 0.155672
R973 VTAIL.n380 VTAIL.n367 0.155672
R974 VTAIL.n387 VTAIL.n367 0.155672
R975 VTAIL.n388 VTAIL.n387 0.155672
R976 VTAIL.n388 VTAIL.n363 0.155672
R977 VTAIL.n395 VTAIL.n363 0.155672
R978 VTAIL.n396 VTAIL.n395 0.155672
R979 VTAIL.n396 VTAIL.n359 0.155672
R980 VTAIL.n403 VTAIL.n359 0.155672
R981 VTAIL.n404 VTAIL.n403 0.155672
R982 VTAIL.n404 VTAIL.n355 0.155672
R983 VTAIL.n411 VTAIL.n355 0.155672
R984 VTAIL.n412 VTAIL.n411 0.155672
R985 VTAIL.n412 VTAIL.n351 0.155672
R986 VTAIL.n421 VTAIL.n351 0.155672
R987 VTAIL.n422 VTAIL.n421 0.155672
R988 VTAIL.n422 VTAIL.n347 0.155672
R989 VTAIL.n429 VTAIL.n347 0.155672
R990 VTAIL.n430 VTAIL.n429 0.155672
R991 VTAIL.n430 VTAIL.n343 0.155672
R992 VTAIL.n437 VTAIL.n343 0.155672
R993 VTAIL.n438 VTAIL.n437 0.155672
R994 VTAIL.n438 VTAIL.n339 0.155672
R995 VTAIL.n445 VTAIL.n339 0.155672
R996 VTAIL.n43 VTAIL.n35 0.155672
R997 VTAIL.n44 VTAIL.n43 0.155672
R998 VTAIL.n44 VTAIL.n31 0.155672
R999 VTAIL.n51 VTAIL.n31 0.155672
R1000 VTAIL.n52 VTAIL.n51 0.155672
R1001 VTAIL.n52 VTAIL.n27 0.155672
R1002 VTAIL.n59 VTAIL.n27 0.155672
R1003 VTAIL.n60 VTAIL.n59 0.155672
R1004 VTAIL.n60 VTAIL.n23 0.155672
R1005 VTAIL.n67 VTAIL.n23 0.155672
R1006 VTAIL.n68 VTAIL.n67 0.155672
R1007 VTAIL.n68 VTAIL.n19 0.155672
R1008 VTAIL.n75 VTAIL.n19 0.155672
R1009 VTAIL.n76 VTAIL.n75 0.155672
R1010 VTAIL.n76 VTAIL.n15 0.155672
R1011 VTAIL.n85 VTAIL.n15 0.155672
R1012 VTAIL.n86 VTAIL.n85 0.155672
R1013 VTAIL.n86 VTAIL.n11 0.155672
R1014 VTAIL.n93 VTAIL.n11 0.155672
R1015 VTAIL.n94 VTAIL.n93 0.155672
R1016 VTAIL.n94 VTAIL.n7 0.155672
R1017 VTAIL.n101 VTAIL.n7 0.155672
R1018 VTAIL.n102 VTAIL.n101 0.155672
R1019 VTAIL.n102 VTAIL.n3 0.155672
R1020 VTAIL.n109 VTAIL.n3 0.155672
R1021 VTAIL.n335 VTAIL.n229 0.155672
R1022 VTAIL.n328 VTAIL.n229 0.155672
R1023 VTAIL.n328 VTAIL.n327 0.155672
R1024 VTAIL.n327 VTAIL.n233 0.155672
R1025 VTAIL.n320 VTAIL.n233 0.155672
R1026 VTAIL.n320 VTAIL.n319 0.155672
R1027 VTAIL.n319 VTAIL.n237 0.155672
R1028 VTAIL.n312 VTAIL.n237 0.155672
R1029 VTAIL.n312 VTAIL.n311 0.155672
R1030 VTAIL.n311 VTAIL.n241 0.155672
R1031 VTAIL.n304 VTAIL.n241 0.155672
R1032 VTAIL.n304 VTAIL.n303 0.155672
R1033 VTAIL.n303 VTAIL.n247 0.155672
R1034 VTAIL.n296 VTAIL.n247 0.155672
R1035 VTAIL.n296 VTAIL.n295 0.155672
R1036 VTAIL.n295 VTAIL.n251 0.155672
R1037 VTAIL.n288 VTAIL.n251 0.155672
R1038 VTAIL.n288 VTAIL.n287 0.155672
R1039 VTAIL.n287 VTAIL.n255 0.155672
R1040 VTAIL.n280 VTAIL.n255 0.155672
R1041 VTAIL.n280 VTAIL.n279 0.155672
R1042 VTAIL.n279 VTAIL.n259 0.155672
R1043 VTAIL.n272 VTAIL.n259 0.155672
R1044 VTAIL.n272 VTAIL.n271 0.155672
R1045 VTAIL.n271 VTAIL.n263 0.155672
R1046 VTAIL.n223 VTAIL.n117 0.155672
R1047 VTAIL.n216 VTAIL.n117 0.155672
R1048 VTAIL.n216 VTAIL.n215 0.155672
R1049 VTAIL.n215 VTAIL.n121 0.155672
R1050 VTAIL.n208 VTAIL.n121 0.155672
R1051 VTAIL.n208 VTAIL.n207 0.155672
R1052 VTAIL.n207 VTAIL.n125 0.155672
R1053 VTAIL.n200 VTAIL.n125 0.155672
R1054 VTAIL.n200 VTAIL.n199 0.155672
R1055 VTAIL.n199 VTAIL.n129 0.155672
R1056 VTAIL.n192 VTAIL.n129 0.155672
R1057 VTAIL.n192 VTAIL.n191 0.155672
R1058 VTAIL.n191 VTAIL.n135 0.155672
R1059 VTAIL.n184 VTAIL.n135 0.155672
R1060 VTAIL.n184 VTAIL.n183 0.155672
R1061 VTAIL.n183 VTAIL.n139 0.155672
R1062 VTAIL.n176 VTAIL.n139 0.155672
R1063 VTAIL.n176 VTAIL.n175 0.155672
R1064 VTAIL.n175 VTAIL.n143 0.155672
R1065 VTAIL.n168 VTAIL.n143 0.155672
R1066 VTAIL.n168 VTAIL.n167 0.155672
R1067 VTAIL.n167 VTAIL.n147 0.155672
R1068 VTAIL.n160 VTAIL.n147 0.155672
R1069 VTAIL.n160 VTAIL.n159 0.155672
R1070 VTAIL.n159 VTAIL.n151 0.155672
R1071 B.n1095 B.n1094 585
R1072 B.n438 B.n159 585
R1073 B.n437 B.n436 585
R1074 B.n435 B.n434 585
R1075 B.n433 B.n432 585
R1076 B.n431 B.n430 585
R1077 B.n429 B.n428 585
R1078 B.n427 B.n426 585
R1079 B.n425 B.n424 585
R1080 B.n423 B.n422 585
R1081 B.n421 B.n420 585
R1082 B.n419 B.n418 585
R1083 B.n417 B.n416 585
R1084 B.n415 B.n414 585
R1085 B.n413 B.n412 585
R1086 B.n411 B.n410 585
R1087 B.n409 B.n408 585
R1088 B.n407 B.n406 585
R1089 B.n405 B.n404 585
R1090 B.n403 B.n402 585
R1091 B.n401 B.n400 585
R1092 B.n399 B.n398 585
R1093 B.n397 B.n396 585
R1094 B.n395 B.n394 585
R1095 B.n393 B.n392 585
R1096 B.n391 B.n390 585
R1097 B.n389 B.n388 585
R1098 B.n387 B.n386 585
R1099 B.n385 B.n384 585
R1100 B.n383 B.n382 585
R1101 B.n381 B.n380 585
R1102 B.n379 B.n378 585
R1103 B.n377 B.n376 585
R1104 B.n375 B.n374 585
R1105 B.n373 B.n372 585
R1106 B.n371 B.n370 585
R1107 B.n369 B.n368 585
R1108 B.n367 B.n366 585
R1109 B.n365 B.n364 585
R1110 B.n363 B.n362 585
R1111 B.n361 B.n360 585
R1112 B.n359 B.n358 585
R1113 B.n357 B.n356 585
R1114 B.n355 B.n354 585
R1115 B.n353 B.n352 585
R1116 B.n351 B.n350 585
R1117 B.n349 B.n348 585
R1118 B.n347 B.n346 585
R1119 B.n345 B.n344 585
R1120 B.n343 B.n342 585
R1121 B.n341 B.n340 585
R1122 B.n339 B.n338 585
R1123 B.n337 B.n336 585
R1124 B.n335 B.n334 585
R1125 B.n333 B.n332 585
R1126 B.n331 B.n330 585
R1127 B.n329 B.n328 585
R1128 B.n327 B.n326 585
R1129 B.n325 B.n324 585
R1130 B.n323 B.n322 585
R1131 B.n321 B.n320 585
R1132 B.n319 B.n318 585
R1133 B.n317 B.n316 585
R1134 B.n315 B.n314 585
R1135 B.n313 B.n312 585
R1136 B.n311 B.n310 585
R1137 B.n309 B.n308 585
R1138 B.n307 B.n306 585
R1139 B.n305 B.n304 585
R1140 B.n303 B.n302 585
R1141 B.n301 B.n300 585
R1142 B.n299 B.n298 585
R1143 B.n297 B.n296 585
R1144 B.n295 B.n294 585
R1145 B.n293 B.n292 585
R1146 B.n291 B.n290 585
R1147 B.n289 B.n288 585
R1148 B.n287 B.n286 585
R1149 B.n285 B.n284 585
R1150 B.n283 B.n282 585
R1151 B.n281 B.n280 585
R1152 B.n279 B.n278 585
R1153 B.n277 B.n276 585
R1154 B.n275 B.n274 585
R1155 B.n273 B.n272 585
R1156 B.n271 B.n270 585
R1157 B.n269 B.n268 585
R1158 B.n267 B.n266 585
R1159 B.n265 B.n264 585
R1160 B.n263 B.n262 585
R1161 B.n261 B.n260 585
R1162 B.n259 B.n258 585
R1163 B.n257 B.n256 585
R1164 B.n255 B.n254 585
R1165 B.n253 B.n252 585
R1166 B.n251 B.n250 585
R1167 B.n249 B.n248 585
R1168 B.n247 B.n246 585
R1169 B.n245 B.n244 585
R1170 B.n243 B.n242 585
R1171 B.n241 B.n240 585
R1172 B.n239 B.n238 585
R1173 B.n237 B.n236 585
R1174 B.n235 B.n234 585
R1175 B.n233 B.n232 585
R1176 B.n231 B.n230 585
R1177 B.n229 B.n228 585
R1178 B.n227 B.n226 585
R1179 B.n225 B.n224 585
R1180 B.n223 B.n222 585
R1181 B.n221 B.n220 585
R1182 B.n219 B.n218 585
R1183 B.n217 B.n216 585
R1184 B.n215 B.n214 585
R1185 B.n213 B.n212 585
R1186 B.n211 B.n210 585
R1187 B.n209 B.n208 585
R1188 B.n207 B.n206 585
R1189 B.n205 B.n204 585
R1190 B.n203 B.n202 585
R1191 B.n201 B.n200 585
R1192 B.n199 B.n198 585
R1193 B.n197 B.n196 585
R1194 B.n195 B.n194 585
R1195 B.n193 B.n192 585
R1196 B.n191 B.n190 585
R1197 B.n189 B.n188 585
R1198 B.n187 B.n186 585
R1199 B.n185 B.n184 585
R1200 B.n183 B.n182 585
R1201 B.n181 B.n180 585
R1202 B.n179 B.n178 585
R1203 B.n177 B.n176 585
R1204 B.n175 B.n174 585
R1205 B.n173 B.n172 585
R1206 B.n171 B.n170 585
R1207 B.n169 B.n168 585
R1208 B.n167 B.n166 585
R1209 B.n1093 B.n90 585
R1210 B.n1098 B.n90 585
R1211 B.n1092 B.n89 585
R1212 B.n1099 B.n89 585
R1213 B.n1091 B.n1090 585
R1214 B.n1090 B.n85 585
R1215 B.n1089 B.n84 585
R1216 B.n1105 B.n84 585
R1217 B.n1088 B.n83 585
R1218 B.n1106 B.n83 585
R1219 B.n1087 B.n82 585
R1220 B.n1107 B.n82 585
R1221 B.n1086 B.n1085 585
R1222 B.n1085 B.n78 585
R1223 B.n1084 B.n77 585
R1224 B.n1113 B.n77 585
R1225 B.n1083 B.n76 585
R1226 B.n1114 B.n76 585
R1227 B.n1082 B.n75 585
R1228 B.n1115 B.n75 585
R1229 B.n1081 B.n1080 585
R1230 B.n1080 B.n71 585
R1231 B.n1079 B.n70 585
R1232 B.n1121 B.n70 585
R1233 B.n1078 B.n69 585
R1234 B.n1122 B.n69 585
R1235 B.n1077 B.n68 585
R1236 B.n1123 B.n68 585
R1237 B.n1076 B.n1075 585
R1238 B.n1075 B.n64 585
R1239 B.n1074 B.n63 585
R1240 B.n1129 B.n63 585
R1241 B.n1073 B.n62 585
R1242 B.n1130 B.n62 585
R1243 B.n1072 B.n61 585
R1244 B.n1131 B.n61 585
R1245 B.n1071 B.n1070 585
R1246 B.n1070 B.n57 585
R1247 B.n1069 B.n56 585
R1248 B.n1137 B.n56 585
R1249 B.n1068 B.n55 585
R1250 B.n1138 B.n55 585
R1251 B.n1067 B.n54 585
R1252 B.n1139 B.n54 585
R1253 B.n1066 B.n1065 585
R1254 B.n1065 B.n50 585
R1255 B.n1064 B.n49 585
R1256 B.n1145 B.n49 585
R1257 B.n1063 B.n48 585
R1258 B.n1146 B.n48 585
R1259 B.n1062 B.n47 585
R1260 B.n1147 B.n47 585
R1261 B.n1061 B.n1060 585
R1262 B.n1060 B.n43 585
R1263 B.n1059 B.n42 585
R1264 B.n1153 B.n42 585
R1265 B.n1058 B.n41 585
R1266 B.n1154 B.n41 585
R1267 B.n1057 B.n40 585
R1268 B.n1155 B.n40 585
R1269 B.n1056 B.n1055 585
R1270 B.n1055 B.n36 585
R1271 B.n1054 B.n35 585
R1272 B.n1161 B.n35 585
R1273 B.n1053 B.n34 585
R1274 B.n1162 B.n34 585
R1275 B.n1052 B.n33 585
R1276 B.n1163 B.n33 585
R1277 B.n1051 B.n1050 585
R1278 B.n1050 B.n29 585
R1279 B.n1049 B.n28 585
R1280 B.n1169 B.n28 585
R1281 B.n1048 B.n27 585
R1282 B.n1170 B.n27 585
R1283 B.n1047 B.n26 585
R1284 B.n1171 B.n26 585
R1285 B.n1046 B.n1045 585
R1286 B.n1045 B.n22 585
R1287 B.n1044 B.n21 585
R1288 B.n1177 B.n21 585
R1289 B.n1043 B.n20 585
R1290 B.n1178 B.n20 585
R1291 B.n1042 B.n19 585
R1292 B.n1179 B.n19 585
R1293 B.n1041 B.n1040 585
R1294 B.n1040 B.n18 585
R1295 B.n1039 B.n14 585
R1296 B.n1185 B.n14 585
R1297 B.n1038 B.n13 585
R1298 B.n1186 B.n13 585
R1299 B.n1037 B.n12 585
R1300 B.n1187 B.n12 585
R1301 B.n1036 B.n1035 585
R1302 B.n1035 B.n8 585
R1303 B.n1034 B.n7 585
R1304 B.n1193 B.n7 585
R1305 B.n1033 B.n6 585
R1306 B.n1194 B.n6 585
R1307 B.n1032 B.n5 585
R1308 B.n1195 B.n5 585
R1309 B.n1031 B.n1030 585
R1310 B.n1030 B.n4 585
R1311 B.n1029 B.n439 585
R1312 B.n1029 B.n1028 585
R1313 B.n1019 B.n440 585
R1314 B.n441 B.n440 585
R1315 B.n1021 B.n1020 585
R1316 B.n1022 B.n1021 585
R1317 B.n1018 B.n446 585
R1318 B.n446 B.n445 585
R1319 B.n1017 B.n1016 585
R1320 B.n1016 B.n1015 585
R1321 B.n448 B.n447 585
R1322 B.n1008 B.n448 585
R1323 B.n1007 B.n1006 585
R1324 B.n1009 B.n1007 585
R1325 B.n1005 B.n453 585
R1326 B.n453 B.n452 585
R1327 B.n1004 B.n1003 585
R1328 B.n1003 B.n1002 585
R1329 B.n455 B.n454 585
R1330 B.n456 B.n455 585
R1331 B.n995 B.n994 585
R1332 B.n996 B.n995 585
R1333 B.n993 B.n461 585
R1334 B.n461 B.n460 585
R1335 B.n992 B.n991 585
R1336 B.n991 B.n990 585
R1337 B.n463 B.n462 585
R1338 B.n464 B.n463 585
R1339 B.n983 B.n982 585
R1340 B.n984 B.n983 585
R1341 B.n981 B.n468 585
R1342 B.n472 B.n468 585
R1343 B.n980 B.n979 585
R1344 B.n979 B.n978 585
R1345 B.n470 B.n469 585
R1346 B.n471 B.n470 585
R1347 B.n971 B.n970 585
R1348 B.n972 B.n971 585
R1349 B.n969 B.n477 585
R1350 B.n477 B.n476 585
R1351 B.n968 B.n967 585
R1352 B.n967 B.n966 585
R1353 B.n479 B.n478 585
R1354 B.n480 B.n479 585
R1355 B.n959 B.n958 585
R1356 B.n960 B.n959 585
R1357 B.n957 B.n485 585
R1358 B.n485 B.n484 585
R1359 B.n956 B.n955 585
R1360 B.n955 B.n954 585
R1361 B.n487 B.n486 585
R1362 B.n488 B.n487 585
R1363 B.n947 B.n946 585
R1364 B.n948 B.n947 585
R1365 B.n945 B.n493 585
R1366 B.n493 B.n492 585
R1367 B.n944 B.n943 585
R1368 B.n943 B.n942 585
R1369 B.n495 B.n494 585
R1370 B.n496 B.n495 585
R1371 B.n935 B.n934 585
R1372 B.n936 B.n935 585
R1373 B.n933 B.n501 585
R1374 B.n501 B.n500 585
R1375 B.n932 B.n931 585
R1376 B.n931 B.n930 585
R1377 B.n503 B.n502 585
R1378 B.n504 B.n503 585
R1379 B.n923 B.n922 585
R1380 B.n924 B.n923 585
R1381 B.n921 B.n509 585
R1382 B.n509 B.n508 585
R1383 B.n920 B.n919 585
R1384 B.n919 B.n918 585
R1385 B.n511 B.n510 585
R1386 B.n512 B.n511 585
R1387 B.n911 B.n910 585
R1388 B.n912 B.n911 585
R1389 B.n909 B.n516 585
R1390 B.n520 B.n516 585
R1391 B.n908 B.n907 585
R1392 B.n907 B.n906 585
R1393 B.n518 B.n517 585
R1394 B.n519 B.n518 585
R1395 B.n899 B.n898 585
R1396 B.n900 B.n899 585
R1397 B.n897 B.n525 585
R1398 B.n525 B.n524 585
R1399 B.n896 B.n895 585
R1400 B.n895 B.n894 585
R1401 B.n527 B.n526 585
R1402 B.n528 B.n527 585
R1403 B.n887 B.n886 585
R1404 B.n888 B.n887 585
R1405 B.n885 B.n533 585
R1406 B.n533 B.n532 585
R1407 B.n880 B.n879 585
R1408 B.n878 B.n604 585
R1409 B.n877 B.n603 585
R1410 B.n882 B.n603 585
R1411 B.n876 B.n875 585
R1412 B.n874 B.n873 585
R1413 B.n872 B.n871 585
R1414 B.n870 B.n869 585
R1415 B.n868 B.n867 585
R1416 B.n866 B.n865 585
R1417 B.n864 B.n863 585
R1418 B.n862 B.n861 585
R1419 B.n860 B.n859 585
R1420 B.n858 B.n857 585
R1421 B.n856 B.n855 585
R1422 B.n854 B.n853 585
R1423 B.n852 B.n851 585
R1424 B.n850 B.n849 585
R1425 B.n848 B.n847 585
R1426 B.n846 B.n845 585
R1427 B.n844 B.n843 585
R1428 B.n842 B.n841 585
R1429 B.n840 B.n839 585
R1430 B.n838 B.n837 585
R1431 B.n836 B.n835 585
R1432 B.n834 B.n833 585
R1433 B.n832 B.n831 585
R1434 B.n830 B.n829 585
R1435 B.n828 B.n827 585
R1436 B.n826 B.n825 585
R1437 B.n824 B.n823 585
R1438 B.n822 B.n821 585
R1439 B.n820 B.n819 585
R1440 B.n818 B.n817 585
R1441 B.n816 B.n815 585
R1442 B.n814 B.n813 585
R1443 B.n812 B.n811 585
R1444 B.n810 B.n809 585
R1445 B.n808 B.n807 585
R1446 B.n806 B.n805 585
R1447 B.n804 B.n803 585
R1448 B.n802 B.n801 585
R1449 B.n800 B.n799 585
R1450 B.n798 B.n797 585
R1451 B.n796 B.n795 585
R1452 B.n794 B.n793 585
R1453 B.n792 B.n791 585
R1454 B.n790 B.n789 585
R1455 B.n788 B.n787 585
R1456 B.n786 B.n785 585
R1457 B.n784 B.n783 585
R1458 B.n782 B.n781 585
R1459 B.n780 B.n779 585
R1460 B.n778 B.n777 585
R1461 B.n776 B.n775 585
R1462 B.n774 B.n773 585
R1463 B.n772 B.n771 585
R1464 B.n770 B.n769 585
R1465 B.n768 B.n767 585
R1466 B.n766 B.n765 585
R1467 B.n764 B.n763 585
R1468 B.n762 B.n761 585
R1469 B.n760 B.n759 585
R1470 B.n758 B.n757 585
R1471 B.n756 B.n755 585
R1472 B.n753 B.n752 585
R1473 B.n751 B.n750 585
R1474 B.n749 B.n748 585
R1475 B.n747 B.n746 585
R1476 B.n745 B.n744 585
R1477 B.n743 B.n742 585
R1478 B.n741 B.n740 585
R1479 B.n739 B.n738 585
R1480 B.n737 B.n736 585
R1481 B.n735 B.n734 585
R1482 B.n732 B.n731 585
R1483 B.n730 B.n729 585
R1484 B.n728 B.n727 585
R1485 B.n726 B.n725 585
R1486 B.n724 B.n723 585
R1487 B.n722 B.n721 585
R1488 B.n720 B.n719 585
R1489 B.n718 B.n717 585
R1490 B.n716 B.n715 585
R1491 B.n714 B.n713 585
R1492 B.n712 B.n711 585
R1493 B.n710 B.n709 585
R1494 B.n708 B.n707 585
R1495 B.n706 B.n705 585
R1496 B.n704 B.n703 585
R1497 B.n702 B.n701 585
R1498 B.n700 B.n699 585
R1499 B.n698 B.n697 585
R1500 B.n696 B.n695 585
R1501 B.n694 B.n693 585
R1502 B.n692 B.n691 585
R1503 B.n690 B.n689 585
R1504 B.n688 B.n687 585
R1505 B.n686 B.n685 585
R1506 B.n684 B.n683 585
R1507 B.n682 B.n681 585
R1508 B.n680 B.n679 585
R1509 B.n678 B.n677 585
R1510 B.n676 B.n675 585
R1511 B.n674 B.n673 585
R1512 B.n672 B.n671 585
R1513 B.n670 B.n669 585
R1514 B.n668 B.n667 585
R1515 B.n666 B.n665 585
R1516 B.n664 B.n663 585
R1517 B.n662 B.n661 585
R1518 B.n660 B.n659 585
R1519 B.n658 B.n657 585
R1520 B.n656 B.n655 585
R1521 B.n654 B.n653 585
R1522 B.n652 B.n651 585
R1523 B.n650 B.n649 585
R1524 B.n648 B.n647 585
R1525 B.n646 B.n645 585
R1526 B.n644 B.n643 585
R1527 B.n642 B.n641 585
R1528 B.n640 B.n639 585
R1529 B.n638 B.n637 585
R1530 B.n636 B.n635 585
R1531 B.n634 B.n633 585
R1532 B.n632 B.n631 585
R1533 B.n630 B.n629 585
R1534 B.n628 B.n627 585
R1535 B.n626 B.n625 585
R1536 B.n624 B.n623 585
R1537 B.n622 B.n621 585
R1538 B.n620 B.n619 585
R1539 B.n618 B.n617 585
R1540 B.n616 B.n615 585
R1541 B.n614 B.n613 585
R1542 B.n612 B.n611 585
R1543 B.n610 B.n609 585
R1544 B.n535 B.n534 585
R1545 B.n884 B.n883 585
R1546 B.n883 B.n882 585
R1547 B.n531 B.n530 585
R1548 B.n532 B.n531 585
R1549 B.n890 B.n889 585
R1550 B.n889 B.n888 585
R1551 B.n891 B.n529 585
R1552 B.n529 B.n528 585
R1553 B.n893 B.n892 585
R1554 B.n894 B.n893 585
R1555 B.n523 B.n522 585
R1556 B.n524 B.n523 585
R1557 B.n902 B.n901 585
R1558 B.n901 B.n900 585
R1559 B.n903 B.n521 585
R1560 B.n521 B.n519 585
R1561 B.n905 B.n904 585
R1562 B.n906 B.n905 585
R1563 B.n515 B.n514 585
R1564 B.n520 B.n515 585
R1565 B.n914 B.n913 585
R1566 B.n913 B.n912 585
R1567 B.n915 B.n513 585
R1568 B.n513 B.n512 585
R1569 B.n917 B.n916 585
R1570 B.n918 B.n917 585
R1571 B.n507 B.n506 585
R1572 B.n508 B.n507 585
R1573 B.n926 B.n925 585
R1574 B.n925 B.n924 585
R1575 B.n927 B.n505 585
R1576 B.n505 B.n504 585
R1577 B.n929 B.n928 585
R1578 B.n930 B.n929 585
R1579 B.n499 B.n498 585
R1580 B.n500 B.n499 585
R1581 B.n938 B.n937 585
R1582 B.n937 B.n936 585
R1583 B.n939 B.n497 585
R1584 B.n497 B.n496 585
R1585 B.n941 B.n940 585
R1586 B.n942 B.n941 585
R1587 B.n491 B.n490 585
R1588 B.n492 B.n491 585
R1589 B.n950 B.n949 585
R1590 B.n949 B.n948 585
R1591 B.n951 B.n489 585
R1592 B.n489 B.n488 585
R1593 B.n953 B.n952 585
R1594 B.n954 B.n953 585
R1595 B.n483 B.n482 585
R1596 B.n484 B.n483 585
R1597 B.n962 B.n961 585
R1598 B.n961 B.n960 585
R1599 B.n963 B.n481 585
R1600 B.n481 B.n480 585
R1601 B.n965 B.n964 585
R1602 B.n966 B.n965 585
R1603 B.n475 B.n474 585
R1604 B.n476 B.n475 585
R1605 B.n974 B.n973 585
R1606 B.n973 B.n972 585
R1607 B.n975 B.n473 585
R1608 B.n473 B.n471 585
R1609 B.n977 B.n976 585
R1610 B.n978 B.n977 585
R1611 B.n467 B.n466 585
R1612 B.n472 B.n467 585
R1613 B.n986 B.n985 585
R1614 B.n985 B.n984 585
R1615 B.n987 B.n465 585
R1616 B.n465 B.n464 585
R1617 B.n989 B.n988 585
R1618 B.n990 B.n989 585
R1619 B.n459 B.n458 585
R1620 B.n460 B.n459 585
R1621 B.n998 B.n997 585
R1622 B.n997 B.n996 585
R1623 B.n999 B.n457 585
R1624 B.n457 B.n456 585
R1625 B.n1001 B.n1000 585
R1626 B.n1002 B.n1001 585
R1627 B.n451 B.n450 585
R1628 B.n452 B.n451 585
R1629 B.n1011 B.n1010 585
R1630 B.n1010 B.n1009 585
R1631 B.n1012 B.n449 585
R1632 B.n1008 B.n449 585
R1633 B.n1014 B.n1013 585
R1634 B.n1015 B.n1014 585
R1635 B.n444 B.n443 585
R1636 B.n445 B.n444 585
R1637 B.n1024 B.n1023 585
R1638 B.n1023 B.n1022 585
R1639 B.n1025 B.n442 585
R1640 B.n442 B.n441 585
R1641 B.n1027 B.n1026 585
R1642 B.n1028 B.n1027 585
R1643 B.n2 B.n0 585
R1644 B.n4 B.n2 585
R1645 B.n3 B.n1 585
R1646 B.n1194 B.n3 585
R1647 B.n1192 B.n1191 585
R1648 B.n1193 B.n1192 585
R1649 B.n1190 B.n9 585
R1650 B.n9 B.n8 585
R1651 B.n1189 B.n1188 585
R1652 B.n1188 B.n1187 585
R1653 B.n11 B.n10 585
R1654 B.n1186 B.n11 585
R1655 B.n1184 B.n1183 585
R1656 B.n1185 B.n1184 585
R1657 B.n1182 B.n15 585
R1658 B.n18 B.n15 585
R1659 B.n1181 B.n1180 585
R1660 B.n1180 B.n1179 585
R1661 B.n17 B.n16 585
R1662 B.n1178 B.n17 585
R1663 B.n1176 B.n1175 585
R1664 B.n1177 B.n1176 585
R1665 B.n1174 B.n23 585
R1666 B.n23 B.n22 585
R1667 B.n1173 B.n1172 585
R1668 B.n1172 B.n1171 585
R1669 B.n25 B.n24 585
R1670 B.n1170 B.n25 585
R1671 B.n1168 B.n1167 585
R1672 B.n1169 B.n1168 585
R1673 B.n1166 B.n30 585
R1674 B.n30 B.n29 585
R1675 B.n1165 B.n1164 585
R1676 B.n1164 B.n1163 585
R1677 B.n32 B.n31 585
R1678 B.n1162 B.n32 585
R1679 B.n1160 B.n1159 585
R1680 B.n1161 B.n1160 585
R1681 B.n1158 B.n37 585
R1682 B.n37 B.n36 585
R1683 B.n1157 B.n1156 585
R1684 B.n1156 B.n1155 585
R1685 B.n39 B.n38 585
R1686 B.n1154 B.n39 585
R1687 B.n1152 B.n1151 585
R1688 B.n1153 B.n1152 585
R1689 B.n1150 B.n44 585
R1690 B.n44 B.n43 585
R1691 B.n1149 B.n1148 585
R1692 B.n1148 B.n1147 585
R1693 B.n46 B.n45 585
R1694 B.n1146 B.n46 585
R1695 B.n1144 B.n1143 585
R1696 B.n1145 B.n1144 585
R1697 B.n1142 B.n51 585
R1698 B.n51 B.n50 585
R1699 B.n1141 B.n1140 585
R1700 B.n1140 B.n1139 585
R1701 B.n53 B.n52 585
R1702 B.n1138 B.n53 585
R1703 B.n1136 B.n1135 585
R1704 B.n1137 B.n1136 585
R1705 B.n1134 B.n58 585
R1706 B.n58 B.n57 585
R1707 B.n1133 B.n1132 585
R1708 B.n1132 B.n1131 585
R1709 B.n60 B.n59 585
R1710 B.n1130 B.n60 585
R1711 B.n1128 B.n1127 585
R1712 B.n1129 B.n1128 585
R1713 B.n1126 B.n65 585
R1714 B.n65 B.n64 585
R1715 B.n1125 B.n1124 585
R1716 B.n1124 B.n1123 585
R1717 B.n67 B.n66 585
R1718 B.n1122 B.n67 585
R1719 B.n1120 B.n1119 585
R1720 B.n1121 B.n1120 585
R1721 B.n1118 B.n72 585
R1722 B.n72 B.n71 585
R1723 B.n1117 B.n1116 585
R1724 B.n1116 B.n1115 585
R1725 B.n74 B.n73 585
R1726 B.n1114 B.n74 585
R1727 B.n1112 B.n1111 585
R1728 B.n1113 B.n1112 585
R1729 B.n1110 B.n79 585
R1730 B.n79 B.n78 585
R1731 B.n1109 B.n1108 585
R1732 B.n1108 B.n1107 585
R1733 B.n81 B.n80 585
R1734 B.n1106 B.n81 585
R1735 B.n1104 B.n1103 585
R1736 B.n1105 B.n1104 585
R1737 B.n1102 B.n86 585
R1738 B.n86 B.n85 585
R1739 B.n1101 B.n1100 585
R1740 B.n1100 B.n1099 585
R1741 B.n88 B.n87 585
R1742 B.n1098 B.n88 585
R1743 B.n1197 B.n1196 585
R1744 B.n1196 B.n1195 585
R1745 B.n607 B.t19 481.632
R1746 B.n160 B.t8 481.632
R1747 B.n605 B.t16 481.632
R1748 B.n163 B.t11 481.632
R1749 B.n880 B.n531 463.671
R1750 B.n166 B.n88 463.671
R1751 B.n883 B.n533 463.671
R1752 B.n1095 B.n90 463.671
R1753 B.n608 B.t18 414.529
R1754 B.n161 B.t9 414.529
R1755 B.n606 B.t15 414.529
R1756 B.n164 B.t12 414.529
R1757 B.n607 B.t17 360.18
R1758 B.n605 B.t13 360.18
R1759 B.n163 B.t10 360.18
R1760 B.n160 B.t6 360.18
R1761 B.n1097 B.n1096 256.663
R1762 B.n1097 B.n158 256.663
R1763 B.n1097 B.n157 256.663
R1764 B.n1097 B.n156 256.663
R1765 B.n1097 B.n155 256.663
R1766 B.n1097 B.n154 256.663
R1767 B.n1097 B.n153 256.663
R1768 B.n1097 B.n152 256.663
R1769 B.n1097 B.n151 256.663
R1770 B.n1097 B.n150 256.663
R1771 B.n1097 B.n149 256.663
R1772 B.n1097 B.n148 256.663
R1773 B.n1097 B.n147 256.663
R1774 B.n1097 B.n146 256.663
R1775 B.n1097 B.n145 256.663
R1776 B.n1097 B.n144 256.663
R1777 B.n1097 B.n143 256.663
R1778 B.n1097 B.n142 256.663
R1779 B.n1097 B.n141 256.663
R1780 B.n1097 B.n140 256.663
R1781 B.n1097 B.n139 256.663
R1782 B.n1097 B.n138 256.663
R1783 B.n1097 B.n137 256.663
R1784 B.n1097 B.n136 256.663
R1785 B.n1097 B.n135 256.663
R1786 B.n1097 B.n134 256.663
R1787 B.n1097 B.n133 256.663
R1788 B.n1097 B.n132 256.663
R1789 B.n1097 B.n131 256.663
R1790 B.n1097 B.n130 256.663
R1791 B.n1097 B.n129 256.663
R1792 B.n1097 B.n128 256.663
R1793 B.n1097 B.n127 256.663
R1794 B.n1097 B.n126 256.663
R1795 B.n1097 B.n125 256.663
R1796 B.n1097 B.n124 256.663
R1797 B.n1097 B.n123 256.663
R1798 B.n1097 B.n122 256.663
R1799 B.n1097 B.n121 256.663
R1800 B.n1097 B.n120 256.663
R1801 B.n1097 B.n119 256.663
R1802 B.n1097 B.n118 256.663
R1803 B.n1097 B.n117 256.663
R1804 B.n1097 B.n116 256.663
R1805 B.n1097 B.n115 256.663
R1806 B.n1097 B.n114 256.663
R1807 B.n1097 B.n113 256.663
R1808 B.n1097 B.n112 256.663
R1809 B.n1097 B.n111 256.663
R1810 B.n1097 B.n110 256.663
R1811 B.n1097 B.n109 256.663
R1812 B.n1097 B.n108 256.663
R1813 B.n1097 B.n107 256.663
R1814 B.n1097 B.n106 256.663
R1815 B.n1097 B.n105 256.663
R1816 B.n1097 B.n104 256.663
R1817 B.n1097 B.n103 256.663
R1818 B.n1097 B.n102 256.663
R1819 B.n1097 B.n101 256.663
R1820 B.n1097 B.n100 256.663
R1821 B.n1097 B.n99 256.663
R1822 B.n1097 B.n98 256.663
R1823 B.n1097 B.n97 256.663
R1824 B.n1097 B.n96 256.663
R1825 B.n1097 B.n95 256.663
R1826 B.n1097 B.n94 256.663
R1827 B.n1097 B.n93 256.663
R1828 B.n1097 B.n92 256.663
R1829 B.n1097 B.n91 256.663
R1830 B.n882 B.n881 256.663
R1831 B.n882 B.n536 256.663
R1832 B.n882 B.n537 256.663
R1833 B.n882 B.n538 256.663
R1834 B.n882 B.n539 256.663
R1835 B.n882 B.n540 256.663
R1836 B.n882 B.n541 256.663
R1837 B.n882 B.n542 256.663
R1838 B.n882 B.n543 256.663
R1839 B.n882 B.n544 256.663
R1840 B.n882 B.n545 256.663
R1841 B.n882 B.n546 256.663
R1842 B.n882 B.n547 256.663
R1843 B.n882 B.n548 256.663
R1844 B.n882 B.n549 256.663
R1845 B.n882 B.n550 256.663
R1846 B.n882 B.n551 256.663
R1847 B.n882 B.n552 256.663
R1848 B.n882 B.n553 256.663
R1849 B.n882 B.n554 256.663
R1850 B.n882 B.n555 256.663
R1851 B.n882 B.n556 256.663
R1852 B.n882 B.n557 256.663
R1853 B.n882 B.n558 256.663
R1854 B.n882 B.n559 256.663
R1855 B.n882 B.n560 256.663
R1856 B.n882 B.n561 256.663
R1857 B.n882 B.n562 256.663
R1858 B.n882 B.n563 256.663
R1859 B.n882 B.n564 256.663
R1860 B.n882 B.n565 256.663
R1861 B.n882 B.n566 256.663
R1862 B.n882 B.n567 256.663
R1863 B.n882 B.n568 256.663
R1864 B.n882 B.n569 256.663
R1865 B.n882 B.n570 256.663
R1866 B.n882 B.n571 256.663
R1867 B.n882 B.n572 256.663
R1868 B.n882 B.n573 256.663
R1869 B.n882 B.n574 256.663
R1870 B.n882 B.n575 256.663
R1871 B.n882 B.n576 256.663
R1872 B.n882 B.n577 256.663
R1873 B.n882 B.n578 256.663
R1874 B.n882 B.n579 256.663
R1875 B.n882 B.n580 256.663
R1876 B.n882 B.n581 256.663
R1877 B.n882 B.n582 256.663
R1878 B.n882 B.n583 256.663
R1879 B.n882 B.n584 256.663
R1880 B.n882 B.n585 256.663
R1881 B.n882 B.n586 256.663
R1882 B.n882 B.n587 256.663
R1883 B.n882 B.n588 256.663
R1884 B.n882 B.n589 256.663
R1885 B.n882 B.n590 256.663
R1886 B.n882 B.n591 256.663
R1887 B.n882 B.n592 256.663
R1888 B.n882 B.n593 256.663
R1889 B.n882 B.n594 256.663
R1890 B.n882 B.n595 256.663
R1891 B.n882 B.n596 256.663
R1892 B.n882 B.n597 256.663
R1893 B.n882 B.n598 256.663
R1894 B.n882 B.n599 256.663
R1895 B.n882 B.n600 256.663
R1896 B.n882 B.n601 256.663
R1897 B.n882 B.n602 256.663
R1898 B.n889 B.n531 163.367
R1899 B.n889 B.n529 163.367
R1900 B.n893 B.n529 163.367
R1901 B.n893 B.n523 163.367
R1902 B.n901 B.n523 163.367
R1903 B.n901 B.n521 163.367
R1904 B.n905 B.n521 163.367
R1905 B.n905 B.n515 163.367
R1906 B.n913 B.n515 163.367
R1907 B.n913 B.n513 163.367
R1908 B.n917 B.n513 163.367
R1909 B.n917 B.n507 163.367
R1910 B.n925 B.n507 163.367
R1911 B.n925 B.n505 163.367
R1912 B.n929 B.n505 163.367
R1913 B.n929 B.n499 163.367
R1914 B.n937 B.n499 163.367
R1915 B.n937 B.n497 163.367
R1916 B.n941 B.n497 163.367
R1917 B.n941 B.n491 163.367
R1918 B.n949 B.n491 163.367
R1919 B.n949 B.n489 163.367
R1920 B.n953 B.n489 163.367
R1921 B.n953 B.n483 163.367
R1922 B.n961 B.n483 163.367
R1923 B.n961 B.n481 163.367
R1924 B.n965 B.n481 163.367
R1925 B.n965 B.n475 163.367
R1926 B.n973 B.n475 163.367
R1927 B.n973 B.n473 163.367
R1928 B.n977 B.n473 163.367
R1929 B.n977 B.n467 163.367
R1930 B.n985 B.n467 163.367
R1931 B.n985 B.n465 163.367
R1932 B.n989 B.n465 163.367
R1933 B.n989 B.n459 163.367
R1934 B.n997 B.n459 163.367
R1935 B.n997 B.n457 163.367
R1936 B.n1001 B.n457 163.367
R1937 B.n1001 B.n451 163.367
R1938 B.n1010 B.n451 163.367
R1939 B.n1010 B.n449 163.367
R1940 B.n1014 B.n449 163.367
R1941 B.n1014 B.n444 163.367
R1942 B.n1023 B.n444 163.367
R1943 B.n1023 B.n442 163.367
R1944 B.n1027 B.n442 163.367
R1945 B.n1027 B.n2 163.367
R1946 B.n1196 B.n2 163.367
R1947 B.n1196 B.n3 163.367
R1948 B.n1192 B.n3 163.367
R1949 B.n1192 B.n9 163.367
R1950 B.n1188 B.n9 163.367
R1951 B.n1188 B.n11 163.367
R1952 B.n1184 B.n11 163.367
R1953 B.n1184 B.n15 163.367
R1954 B.n1180 B.n15 163.367
R1955 B.n1180 B.n17 163.367
R1956 B.n1176 B.n17 163.367
R1957 B.n1176 B.n23 163.367
R1958 B.n1172 B.n23 163.367
R1959 B.n1172 B.n25 163.367
R1960 B.n1168 B.n25 163.367
R1961 B.n1168 B.n30 163.367
R1962 B.n1164 B.n30 163.367
R1963 B.n1164 B.n32 163.367
R1964 B.n1160 B.n32 163.367
R1965 B.n1160 B.n37 163.367
R1966 B.n1156 B.n37 163.367
R1967 B.n1156 B.n39 163.367
R1968 B.n1152 B.n39 163.367
R1969 B.n1152 B.n44 163.367
R1970 B.n1148 B.n44 163.367
R1971 B.n1148 B.n46 163.367
R1972 B.n1144 B.n46 163.367
R1973 B.n1144 B.n51 163.367
R1974 B.n1140 B.n51 163.367
R1975 B.n1140 B.n53 163.367
R1976 B.n1136 B.n53 163.367
R1977 B.n1136 B.n58 163.367
R1978 B.n1132 B.n58 163.367
R1979 B.n1132 B.n60 163.367
R1980 B.n1128 B.n60 163.367
R1981 B.n1128 B.n65 163.367
R1982 B.n1124 B.n65 163.367
R1983 B.n1124 B.n67 163.367
R1984 B.n1120 B.n67 163.367
R1985 B.n1120 B.n72 163.367
R1986 B.n1116 B.n72 163.367
R1987 B.n1116 B.n74 163.367
R1988 B.n1112 B.n74 163.367
R1989 B.n1112 B.n79 163.367
R1990 B.n1108 B.n79 163.367
R1991 B.n1108 B.n81 163.367
R1992 B.n1104 B.n81 163.367
R1993 B.n1104 B.n86 163.367
R1994 B.n1100 B.n86 163.367
R1995 B.n1100 B.n88 163.367
R1996 B.n604 B.n603 163.367
R1997 B.n875 B.n603 163.367
R1998 B.n873 B.n872 163.367
R1999 B.n869 B.n868 163.367
R2000 B.n865 B.n864 163.367
R2001 B.n861 B.n860 163.367
R2002 B.n857 B.n856 163.367
R2003 B.n853 B.n852 163.367
R2004 B.n849 B.n848 163.367
R2005 B.n845 B.n844 163.367
R2006 B.n841 B.n840 163.367
R2007 B.n837 B.n836 163.367
R2008 B.n833 B.n832 163.367
R2009 B.n829 B.n828 163.367
R2010 B.n825 B.n824 163.367
R2011 B.n821 B.n820 163.367
R2012 B.n817 B.n816 163.367
R2013 B.n813 B.n812 163.367
R2014 B.n809 B.n808 163.367
R2015 B.n805 B.n804 163.367
R2016 B.n801 B.n800 163.367
R2017 B.n797 B.n796 163.367
R2018 B.n793 B.n792 163.367
R2019 B.n789 B.n788 163.367
R2020 B.n785 B.n784 163.367
R2021 B.n781 B.n780 163.367
R2022 B.n777 B.n776 163.367
R2023 B.n773 B.n772 163.367
R2024 B.n769 B.n768 163.367
R2025 B.n765 B.n764 163.367
R2026 B.n761 B.n760 163.367
R2027 B.n757 B.n756 163.367
R2028 B.n752 B.n751 163.367
R2029 B.n748 B.n747 163.367
R2030 B.n744 B.n743 163.367
R2031 B.n740 B.n739 163.367
R2032 B.n736 B.n735 163.367
R2033 B.n731 B.n730 163.367
R2034 B.n727 B.n726 163.367
R2035 B.n723 B.n722 163.367
R2036 B.n719 B.n718 163.367
R2037 B.n715 B.n714 163.367
R2038 B.n711 B.n710 163.367
R2039 B.n707 B.n706 163.367
R2040 B.n703 B.n702 163.367
R2041 B.n699 B.n698 163.367
R2042 B.n695 B.n694 163.367
R2043 B.n691 B.n690 163.367
R2044 B.n687 B.n686 163.367
R2045 B.n683 B.n682 163.367
R2046 B.n679 B.n678 163.367
R2047 B.n675 B.n674 163.367
R2048 B.n671 B.n670 163.367
R2049 B.n667 B.n666 163.367
R2050 B.n663 B.n662 163.367
R2051 B.n659 B.n658 163.367
R2052 B.n655 B.n654 163.367
R2053 B.n651 B.n650 163.367
R2054 B.n647 B.n646 163.367
R2055 B.n643 B.n642 163.367
R2056 B.n639 B.n638 163.367
R2057 B.n635 B.n634 163.367
R2058 B.n631 B.n630 163.367
R2059 B.n627 B.n626 163.367
R2060 B.n623 B.n622 163.367
R2061 B.n619 B.n618 163.367
R2062 B.n615 B.n614 163.367
R2063 B.n611 B.n610 163.367
R2064 B.n883 B.n535 163.367
R2065 B.n887 B.n533 163.367
R2066 B.n887 B.n527 163.367
R2067 B.n895 B.n527 163.367
R2068 B.n895 B.n525 163.367
R2069 B.n899 B.n525 163.367
R2070 B.n899 B.n518 163.367
R2071 B.n907 B.n518 163.367
R2072 B.n907 B.n516 163.367
R2073 B.n911 B.n516 163.367
R2074 B.n911 B.n511 163.367
R2075 B.n919 B.n511 163.367
R2076 B.n919 B.n509 163.367
R2077 B.n923 B.n509 163.367
R2078 B.n923 B.n503 163.367
R2079 B.n931 B.n503 163.367
R2080 B.n931 B.n501 163.367
R2081 B.n935 B.n501 163.367
R2082 B.n935 B.n495 163.367
R2083 B.n943 B.n495 163.367
R2084 B.n943 B.n493 163.367
R2085 B.n947 B.n493 163.367
R2086 B.n947 B.n487 163.367
R2087 B.n955 B.n487 163.367
R2088 B.n955 B.n485 163.367
R2089 B.n959 B.n485 163.367
R2090 B.n959 B.n479 163.367
R2091 B.n967 B.n479 163.367
R2092 B.n967 B.n477 163.367
R2093 B.n971 B.n477 163.367
R2094 B.n971 B.n470 163.367
R2095 B.n979 B.n470 163.367
R2096 B.n979 B.n468 163.367
R2097 B.n983 B.n468 163.367
R2098 B.n983 B.n463 163.367
R2099 B.n991 B.n463 163.367
R2100 B.n991 B.n461 163.367
R2101 B.n995 B.n461 163.367
R2102 B.n995 B.n455 163.367
R2103 B.n1003 B.n455 163.367
R2104 B.n1003 B.n453 163.367
R2105 B.n1007 B.n453 163.367
R2106 B.n1007 B.n448 163.367
R2107 B.n1016 B.n448 163.367
R2108 B.n1016 B.n446 163.367
R2109 B.n1021 B.n446 163.367
R2110 B.n1021 B.n440 163.367
R2111 B.n1029 B.n440 163.367
R2112 B.n1030 B.n1029 163.367
R2113 B.n1030 B.n5 163.367
R2114 B.n6 B.n5 163.367
R2115 B.n7 B.n6 163.367
R2116 B.n1035 B.n7 163.367
R2117 B.n1035 B.n12 163.367
R2118 B.n13 B.n12 163.367
R2119 B.n14 B.n13 163.367
R2120 B.n1040 B.n14 163.367
R2121 B.n1040 B.n19 163.367
R2122 B.n20 B.n19 163.367
R2123 B.n21 B.n20 163.367
R2124 B.n1045 B.n21 163.367
R2125 B.n1045 B.n26 163.367
R2126 B.n27 B.n26 163.367
R2127 B.n28 B.n27 163.367
R2128 B.n1050 B.n28 163.367
R2129 B.n1050 B.n33 163.367
R2130 B.n34 B.n33 163.367
R2131 B.n35 B.n34 163.367
R2132 B.n1055 B.n35 163.367
R2133 B.n1055 B.n40 163.367
R2134 B.n41 B.n40 163.367
R2135 B.n42 B.n41 163.367
R2136 B.n1060 B.n42 163.367
R2137 B.n1060 B.n47 163.367
R2138 B.n48 B.n47 163.367
R2139 B.n49 B.n48 163.367
R2140 B.n1065 B.n49 163.367
R2141 B.n1065 B.n54 163.367
R2142 B.n55 B.n54 163.367
R2143 B.n56 B.n55 163.367
R2144 B.n1070 B.n56 163.367
R2145 B.n1070 B.n61 163.367
R2146 B.n62 B.n61 163.367
R2147 B.n63 B.n62 163.367
R2148 B.n1075 B.n63 163.367
R2149 B.n1075 B.n68 163.367
R2150 B.n69 B.n68 163.367
R2151 B.n70 B.n69 163.367
R2152 B.n1080 B.n70 163.367
R2153 B.n1080 B.n75 163.367
R2154 B.n76 B.n75 163.367
R2155 B.n77 B.n76 163.367
R2156 B.n1085 B.n77 163.367
R2157 B.n1085 B.n82 163.367
R2158 B.n83 B.n82 163.367
R2159 B.n84 B.n83 163.367
R2160 B.n1090 B.n84 163.367
R2161 B.n1090 B.n89 163.367
R2162 B.n90 B.n89 163.367
R2163 B.n170 B.n169 163.367
R2164 B.n174 B.n173 163.367
R2165 B.n178 B.n177 163.367
R2166 B.n182 B.n181 163.367
R2167 B.n186 B.n185 163.367
R2168 B.n190 B.n189 163.367
R2169 B.n194 B.n193 163.367
R2170 B.n198 B.n197 163.367
R2171 B.n202 B.n201 163.367
R2172 B.n206 B.n205 163.367
R2173 B.n210 B.n209 163.367
R2174 B.n214 B.n213 163.367
R2175 B.n218 B.n217 163.367
R2176 B.n222 B.n221 163.367
R2177 B.n226 B.n225 163.367
R2178 B.n230 B.n229 163.367
R2179 B.n234 B.n233 163.367
R2180 B.n238 B.n237 163.367
R2181 B.n242 B.n241 163.367
R2182 B.n246 B.n245 163.367
R2183 B.n250 B.n249 163.367
R2184 B.n254 B.n253 163.367
R2185 B.n258 B.n257 163.367
R2186 B.n262 B.n261 163.367
R2187 B.n266 B.n265 163.367
R2188 B.n270 B.n269 163.367
R2189 B.n274 B.n273 163.367
R2190 B.n278 B.n277 163.367
R2191 B.n282 B.n281 163.367
R2192 B.n286 B.n285 163.367
R2193 B.n290 B.n289 163.367
R2194 B.n294 B.n293 163.367
R2195 B.n298 B.n297 163.367
R2196 B.n302 B.n301 163.367
R2197 B.n306 B.n305 163.367
R2198 B.n310 B.n309 163.367
R2199 B.n314 B.n313 163.367
R2200 B.n318 B.n317 163.367
R2201 B.n322 B.n321 163.367
R2202 B.n326 B.n325 163.367
R2203 B.n330 B.n329 163.367
R2204 B.n334 B.n333 163.367
R2205 B.n338 B.n337 163.367
R2206 B.n342 B.n341 163.367
R2207 B.n346 B.n345 163.367
R2208 B.n350 B.n349 163.367
R2209 B.n354 B.n353 163.367
R2210 B.n358 B.n357 163.367
R2211 B.n362 B.n361 163.367
R2212 B.n366 B.n365 163.367
R2213 B.n370 B.n369 163.367
R2214 B.n374 B.n373 163.367
R2215 B.n378 B.n377 163.367
R2216 B.n382 B.n381 163.367
R2217 B.n386 B.n385 163.367
R2218 B.n390 B.n389 163.367
R2219 B.n394 B.n393 163.367
R2220 B.n398 B.n397 163.367
R2221 B.n402 B.n401 163.367
R2222 B.n406 B.n405 163.367
R2223 B.n410 B.n409 163.367
R2224 B.n414 B.n413 163.367
R2225 B.n418 B.n417 163.367
R2226 B.n422 B.n421 163.367
R2227 B.n426 B.n425 163.367
R2228 B.n430 B.n429 163.367
R2229 B.n434 B.n433 163.367
R2230 B.n436 B.n159 163.367
R2231 B.n881 B.n880 71.676
R2232 B.n875 B.n536 71.676
R2233 B.n872 B.n537 71.676
R2234 B.n868 B.n538 71.676
R2235 B.n864 B.n539 71.676
R2236 B.n860 B.n540 71.676
R2237 B.n856 B.n541 71.676
R2238 B.n852 B.n542 71.676
R2239 B.n848 B.n543 71.676
R2240 B.n844 B.n544 71.676
R2241 B.n840 B.n545 71.676
R2242 B.n836 B.n546 71.676
R2243 B.n832 B.n547 71.676
R2244 B.n828 B.n548 71.676
R2245 B.n824 B.n549 71.676
R2246 B.n820 B.n550 71.676
R2247 B.n816 B.n551 71.676
R2248 B.n812 B.n552 71.676
R2249 B.n808 B.n553 71.676
R2250 B.n804 B.n554 71.676
R2251 B.n800 B.n555 71.676
R2252 B.n796 B.n556 71.676
R2253 B.n792 B.n557 71.676
R2254 B.n788 B.n558 71.676
R2255 B.n784 B.n559 71.676
R2256 B.n780 B.n560 71.676
R2257 B.n776 B.n561 71.676
R2258 B.n772 B.n562 71.676
R2259 B.n768 B.n563 71.676
R2260 B.n764 B.n564 71.676
R2261 B.n760 B.n565 71.676
R2262 B.n756 B.n566 71.676
R2263 B.n751 B.n567 71.676
R2264 B.n747 B.n568 71.676
R2265 B.n743 B.n569 71.676
R2266 B.n739 B.n570 71.676
R2267 B.n735 B.n571 71.676
R2268 B.n730 B.n572 71.676
R2269 B.n726 B.n573 71.676
R2270 B.n722 B.n574 71.676
R2271 B.n718 B.n575 71.676
R2272 B.n714 B.n576 71.676
R2273 B.n710 B.n577 71.676
R2274 B.n706 B.n578 71.676
R2275 B.n702 B.n579 71.676
R2276 B.n698 B.n580 71.676
R2277 B.n694 B.n581 71.676
R2278 B.n690 B.n582 71.676
R2279 B.n686 B.n583 71.676
R2280 B.n682 B.n584 71.676
R2281 B.n678 B.n585 71.676
R2282 B.n674 B.n586 71.676
R2283 B.n670 B.n587 71.676
R2284 B.n666 B.n588 71.676
R2285 B.n662 B.n589 71.676
R2286 B.n658 B.n590 71.676
R2287 B.n654 B.n591 71.676
R2288 B.n650 B.n592 71.676
R2289 B.n646 B.n593 71.676
R2290 B.n642 B.n594 71.676
R2291 B.n638 B.n595 71.676
R2292 B.n634 B.n596 71.676
R2293 B.n630 B.n597 71.676
R2294 B.n626 B.n598 71.676
R2295 B.n622 B.n599 71.676
R2296 B.n618 B.n600 71.676
R2297 B.n614 B.n601 71.676
R2298 B.n610 B.n602 71.676
R2299 B.n166 B.n91 71.676
R2300 B.n170 B.n92 71.676
R2301 B.n174 B.n93 71.676
R2302 B.n178 B.n94 71.676
R2303 B.n182 B.n95 71.676
R2304 B.n186 B.n96 71.676
R2305 B.n190 B.n97 71.676
R2306 B.n194 B.n98 71.676
R2307 B.n198 B.n99 71.676
R2308 B.n202 B.n100 71.676
R2309 B.n206 B.n101 71.676
R2310 B.n210 B.n102 71.676
R2311 B.n214 B.n103 71.676
R2312 B.n218 B.n104 71.676
R2313 B.n222 B.n105 71.676
R2314 B.n226 B.n106 71.676
R2315 B.n230 B.n107 71.676
R2316 B.n234 B.n108 71.676
R2317 B.n238 B.n109 71.676
R2318 B.n242 B.n110 71.676
R2319 B.n246 B.n111 71.676
R2320 B.n250 B.n112 71.676
R2321 B.n254 B.n113 71.676
R2322 B.n258 B.n114 71.676
R2323 B.n262 B.n115 71.676
R2324 B.n266 B.n116 71.676
R2325 B.n270 B.n117 71.676
R2326 B.n274 B.n118 71.676
R2327 B.n278 B.n119 71.676
R2328 B.n282 B.n120 71.676
R2329 B.n286 B.n121 71.676
R2330 B.n290 B.n122 71.676
R2331 B.n294 B.n123 71.676
R2332 B.n298 B.n124 71.676
R2333 B.n302 B.n125 71.676
R2334 B.n306 B.n126 71.676
R2335 B.n310 B.n127 71.676
R2336 B.n314 B.n128 71.676
R2337 B.n318 B.n129 71.676
R2338 B.n322 B.n130 71.676
R2339 B.n326 B.n131 71.676
R2340 B.n330 B.n132 71.676
R2341 B.n334 B.n133 71.676
R2342 B.n338 B.n134 71.676
R2343 B.n342 B.n135 71.676
R2344 B.n346 B.n136 71.676
R2345 B.n350 B.n137 71.676
R2346 B.n354 B.n138 71.676
R2347 B.n358 B.n139 71.676
R2348 B.n362 B.n140 71.676
R2349 B.n366 B.n141 71.676
R2350 B.n370 B.n142 71.676
R2351 B.n374 B.n143 71.676
R2352 B.n378 B.n144 71.676
R2353 B.n382 B.n145 71.676
R2354 B.n386 B.n146 71.676
R2355 B.n390 B.n147 71.676
R2356 B.n394 B.n148 71.676
R2357 B.n398 B.n149 71.676
R2358 B.n402 B.n150 71.676
R2359 B.n406 B.n151 71.676
R2360 B.n410 B.n152 71.676
R2361 B.n414 B.n153 71.676
R2362 B.n418 B.n154 71.676
R2363 B.n422 B.n155 71.676
R2364 B.n426 B.n156 71.676
R2365 B.n430 B.n157 71.676
R2366 B.n434 B.n158 71.676
R2367 B.n1096 B.n159 71.676
R2368 B.n1096 B.n1095 71.676
R2369 B.n436 B.n158 71.676
R2370 B.n433 B.n157 71.676
R2371 B.n429 B.n156 71.676
R2372 B.n425 B.n155 71.676
R2373 B.n421 B.n154 71.676
R2374 B.n417 B.n153 71.676
R2375 B.n413 B.n152 71.676
R2376 B.n409 B.n151 71.676
R2377 B.n405 B.n150 71.676
R2378 B.n401 B.n149 71.676
R2379 B.n397 B.n148 71.676
R2380 B.n393 B.n147 71.676
R2381 B.n389 B.n146 71.676
R2382 B.n385 B.n145 71.676
R2383 B.n381 B.n144 71.676
R2384 B.n377 B.n143 71.676
R2385 B.n373 B.n142 71.676
R2386 B.n369 B.n141 71.676
R2387 B.n365 B.n140 71.676
R2388 B.n361 B.n139 71.676
R2389 B.n357 B.n138 71.676
R2390 B.n353 B.n137 71.676
R2391 B.n349 B.n136 71.676
R2392 B.n345 B.n135 71.676
R2393 B.n341 B.n134 71.676
R2394 B.n337 B.n133 71.676
R2395 B.n333 B.n132 71.676
R2396 B.n329 B.n131 71.676
R2397 B.n325 B.n130 71.676
R2398 B.n321 B.n129 71.676
R2399 B.n317 B.n128 71.676
R2400 B.n313 B.n127 71.676
R2401 B.n309 B.n126 71.676
R2402 B.n305 B.n125 71.676
R2403 B.n301 B.n124 71.676
R2404 B.n297 B.n123 71.676
R2405 B.n293 B.n122 71.676
R2406 B.n289 B.n121 71.676
R2407 B.n285 B.n120 71.676
R2408 B.n281 B.n119 71.676
R2409 B.n277 B.n118 71.676
R2410 B.n273 B.n117 71.676
R2411 B.n269 B.n116 71.676
R2412 B.n265 B.n115 71.676
R2413 B.n261 B.n114 71.676
R2414 B.n257 B.n113 71.676
R2415 B.n253 B.n112 71.676
R2416 B.n249 B.n111 71.676
R2417 B.n245 B.n110 71.676
R2418 B.n241 B.n109 71.676
R2419 B.n237 B.n108 71.676
R2420 B.n233 B.n107 71.676
R2421 B.n229 B.n106 71.676
R2422 B.n225 B.n105 71.676
R2423 B.n221 B.n104 71.676
R2424 B.n217 B.n103 71.676
R2425 B.n213 B.n102 71.676
R2426 B.n209 B.n101 71.676
R2427 B.n205 B.n100 71.676
R2428 B.n201 B.n99 71.676
R2429 B.n197 B.n98 71.676
R2430 B.n193 B.n97 71.676
R2431 B.n189 B.n96 71.676
R2432 B.n185 B.n95 71.676
R2433 B.n181 B.n94 71.676
R2434 B.n177 B.n93 71.676
R2435 B.n173 B.n92 71.676
R2436 B.n169 B.n91 71.676
R2437 B.n881 B.n604 71.676
R2438 B.n873 B.n536 71.676
R2439 B.n869 B.n537 71.676
R2440 B.n865 B.n538 71.676
R2441 B.n861 B.n539 71.676
R2442 B.n857 B.n540 71.676
R2443 B.n853 B.n541 71.676
R2444 B.n849 B.n542 71.676
R2445 B.n845 B.n543 71.676
R2446 B.n841 B.n544 71.676
R2447 B.n837 B.n545 71.676
R2448 B.n833 B.n546 71.676
R2449 B.n829 B.n547 71.676
R2450 B.n825 B.n548 71.676
R2451 B.n821 B.n549 71.676
R2452 B.n817 B.n550 71.676
R2453 B.n813 B.n551 71.676
R2454 B.n809 B.n552 71.676
R2455 B.n805 B.n553 71.676
R2456 B.n801 B.n554 71.676
R2457 B.n797 B.n555 71.676
R2458 B.n793 B.n556 71.676
R2459 B.n789 B.n557 71.676
R2460 B.n785 B.n558 71.676
R2461 B.n781 B.n559 71.676
R2462 B.n777 B.n560 71.676
R2463 B.n773 B.n561 71.676
R2464 B.n769 B.n562 71.676
R2465 B.n765 B.n563 71.676
R2466 B.n761 B.n564 71.676
R2467 B.n757 B.n565 71.676
R2468 B.n752 B.n566 71.676
R2469 B.n748 B.n567 71.676
R2470 B.n744 B.n568 71.676
R2471 B.n740 B.n569 71.676
R2472 B.n736 B.n570 71.676
R2473 B.n731 B.n571 71.676
R2474 B.n727 B.n572 71.676
R2475 B.n723 B.n573 71.676
R2476 B.n719 B.n574 71.676
R2477 B.n715 B.n575 71.676
R2478 B.n711 B.n576 71.676
R2479 B.n707 B.n577 71.676
R2480 B.n703 B.n578 71.676
R2481 B.n699 B.n579 71.676
R2482 B.n695 B.n580 71.676
R2483 B.n691 B.n581 71.676
R2484 B.n687 B.n582 71.676
R2485 B.n683 B.n583 71.676
R2486 B.n679 B.n584 71.676
R2487 B.n675 B.n585 71.676
R2488 B.n671 B.n586 71.676
R2489 B.n667 B.n587 71.676
R2490 B.n663 B.n588 71.676
R2491 B.n659 B.n589 71.676
R2492 B.n655 B.n590 71.676
R2493 B.n651 B.n591 71.676
R2494 B.n647 B.n592 71.676
R2495 B.n643 B.n593 71.676
R2496 B.n639 B.n594 71.676
R2497 B.n635 B.n595 71.676
R2498 B.n631 B.n596 71.676
R2499 B.n627 B.n597 71.676
R2500 B.n623 B.n598 71.676
R2501 B.n619 B.n599 71.676
R2502 B.n615 B.n600 71.676
R2503 B.n611 B.n601 71.676
R2504 B.n602 B.n535 71.676
R2505 B.n608 B.n607 67.1035
R2506 B.n606 B.n605 67.1035
R2507 B.n164 B.n163 67.1035
R2508 B.n161 B.n160 67.1035
R2509 B.n733 B.n608 59.5399
R2510 B.n754 B.n606 59.5399
R2511 B.n165 B.n164 59.5399
R2512 B.n162 B.n161 59.5399
R2513 B.n882 B.n532 48.9482
R2514 B.n1098 B.n1097 48.9482
R2515 B.n167 B.n87 30.1273
R2516 B.n885 B.n884 30.1273
R2517 B.n879 B.n530 30.1273
R2518 B.n1094 B.n1093 30.1273
R2519 B.n888 B.n532 29.9865
R2520 B.n888 B.n528 29.9865
R2521 B.n894 B.n528 29.9865
R2522 B.n894 B.n524 29.9865
R2523 B.n900 B.n524 29.9865
R2524 B.n900 B.n519 29.9865
R2525 B.n906 B.n519 29.9865
R2526 B.n906 B.n520 29.9865
R2527 B.n912 B.n512 29.9865
R2528 B.n918 B.n512 29.9865
R2529 B.n918 B.n508 29.9865
R2530 B.n924 B.n508 29.9865
R2531 B.n924 B.n504 29.9865
R2532 B.n930 B.n504 29.9865
R2533 B.n930 B.n500 29.9865
R2534 B.n936 B.n500 29.9865
R2535 B.n936 B.n496 29.9865
R2536 B.n942 B.n496 29.9865
R2537 B.n942 B.n492 29.9865
R2538 B.n948 B.n492 29.9865
R2539 B.n954 B.n488 29.9865
R2540 B.n954 B.n484 29.9865
R2541 B.n960 B.n484 29.9865
R2542 B.n960 B.n480 29.9865
R2543 B.n966 B.n480 29.9865
R2544 B.n966 B.n476 29.9865
R2545 B.n972 B.n476 29.9865
R2546 B.n972 B.n471 29.9865
R2547 B.n978 B.n471 29.9865
R2548 B.n978 B.n472 29.9865
R2549 B.n984 B.n464 29.9865
R2550 B.n990 B.n464 29.9865
R2551 B.n990 B.n460 29.9865
R2552 B.n996 B.n460 29.9865
R2553 B.n996 B.n456 29.9865
R2554 B.n1002 B.n456 29.9865
R2555 B.n1002 B.n452 29.9865
R2556 B.n1009 B.n452 29.9865
R2557 B.n1009 B.n1008 29.9865
R2558 B.n1015 B.n445 29.9865
R2559 B.n1022 B.n445 29.9865
R2560 B.n1022 B.n441 29.9865
R2561 B.n1028 B.n441 29.9865
R2562 B.n1028 B.n4 29.9865
R2563 B.n1195 B.n4 29.9865
R2564 B.n1195 B.n1194 29.9865
R2565 B.n1194 B.n1193 29.9865
R2566 B.n1193 B.n8 29.9865
R2567 B.n1187 B.n8 29.9865
R2568 B.n1187 B.n1186 29.9865
R2569 B.n1186 B.n1185 29.9865
R2570 B.n1179 B.n18 29.9865
R2571 B.n1179 B.n1178 29.9865
R2572 B.n1178 B.n1177 29.9865
R2573 B.n1177 B.n22 29.9865
R2574 B.n1171 B.n22 29.9865
R2575 B.n1171 B.n1170 29.9865
R2576 B.n1170 B.n1169 29.9865
R2577 B.n1169 B.n29 29.9865
R2578 B.n1163 B.n29 29.9865
R2579 B.n1162 B.n1161 29.9865
R2580 B.n1161 B.n36 29.9865
R2581 B.n1155 B.n36 29.9865
R2582 B.n1155 B.n1154 29.9865
R2583 B.n1154 B.n1153 29.9865
R2584 B.n1153 B.n43 29.9865
R2585 B.n1147 B.n43 29.9865
R2586 B.n1147 B.n1146 29.9865
R2587 B.n1146 B.n1145 29.9865
R2588 B.n1145 B.n50 29.9865
R2589 B.n1139 B.n1138 29.9865
R2590 B.n1138 B.n1137 29.9865
R2591 B.n1137 B.n57 29.9865
R2592 B.n1131 B.n57 29.9865
R2593 B.n1131 B.n1130 29.9865
R2594 B.n1130 B.n1129 29.9865
R2595 B.n1129 B.n64 29.9865
R2596 B.n1123 B.n64 29.9865
R2597 B.n1123 B.n1122 29.9865
R2598 B.n1122 B.n1121 29.9865
R2599 B.n1121 B.n71 29.9865
R2600 B.n1115 B.n71 29.9865
R2601 B.n1114 B.n1113 29.9865
R2602 B.n1113 B.n78 29.9865
R2603 B.n1107 B.n78 29.9865
R2604 B.n1107 B.n1106 29.9865
R2605 B.n1106 B.n1105 29.9865
R2606 B.n1105 B.n85 29.9865
R2607 B.n1099 B.n85 29.9865
R2608 B.n1099 B.n1098 29.9865
R2609 B.n948 B.t2 28.6636
R2610 B.n1139 B.t5 28.6636
R2611 B.n984 B.t0 26.0177
R2612 B.n1163 B.t1 26.0177
R2613 B.n1015 B.t4 20.7261
R2614 B.n1185 B.t3 20.7261
R2615 B B.n1197 18.0485
R2616 B.n520 B.t14 17.1983
R2617 B.t7 B.n1114 17.1983
R2618 B.n912 B.t14 12.7886
R2619 B.n1115 B.t7 12.7886
R2620 B.n168 B.n167 10.6151
R2621 B.n171 B.n168 10.6151
R2622 B.n172 B.n171 10.6151
R2623 B.n175 B.n172 10.6151
R2624 B.n176 B.n175 10.6151
R2625 B.n179 B.n176 10.6151
R2626 B.n180 B.n179 10.6151
R2627 B.n183 B.n180 10.6151
R2628 B.n184 B.n183 10.6151
R2629 B.n187 B.n184 10.6151
R2630 B.n188 B.n187 10.6151
R2631 B.n191 B.n188 10.6151
R2632 B.n192 B.n191 10.6151
R2633 B.n195 B.n192 10.6151
R2634 B.n196 B.n195 10.6151
R2635 B.n199 B.n196 10.6151
R2636 B.n200 B.n199 10.6151
R2637 B.n203 B.n200 10.6151
R2638 B.n204 B.n203 10.6151
R2639 B.n207 B.n204 10.6151
R2640 B.n208 B.n207 10.6151
R2641 B.n211 B.n208 10.6151
R2642 B.n212 B.n211 10.6151
R2643 B.n215 B.n212 10.6151
R2644 B.n216 B.n215 10.6151
R2645 B.n219 B.n216 10.6151
R2646 B.n220 B.n219 10.6151
R2647 B.n223 B.n220 10.6151
R2648 B.n224 B.n223 10.6151
R2649 B.n227 B.n224 10.6151
R2650 B.n228 B.n227 10.6151
R2651 B.n231 B.n228 10.6151
R2652 B.n232 B.n231 10.6151
R2653 B.n235 B.n232 10.6151
R2654 B.n236 B.n235 10.6151
R2655 B.n239 B.n236 10.6151
R2656 B.n240 B.n239 10.6151
R2657 B.n243 B.n240 10.6151
R2658 B.n244 B.n243 10.6151
R2659 B.n247 B.n244 10.6151
R2660 B.n248 B.n247 10.6151
R2661 B.n251 B.n248 10.6151
R2662 B.n252 B.n251 10.6151
R2663 B.n255 B.n252 10.6151
R2664 B.n256 B.n255 10.6151
R2665 B.n259 B.n256 10.6151
R2666 B.n260 B.n259 10.6151
R2667 B.n263 B.n260 10.6151
R2668 B.n264 B.n263 10.6151
R2669 B.n267 B.n264 10.6151
R2670 B.n268 B.n267 10.6151
R2671 B.n271 B.n268 10.6151
R2672 B.n272 B.n271 10.6151
R2673 B.n275 B.n272 10.6151
R2674 B.n276 B.n275 10.6151
R2675 B.n279 B.n276 10.6151
R2676 B.n280 B.n279 10.6151
R2677 B.n283 B.n280 10.6151
R2678 B.n284 B.n283 10.6151
R2679 B.n287 B.n284 10.6151
R2680 B.n288 B.n287 10.6151
R2681 B.n291 B.n288 10.6151
R2682 B.n292 B.n291 10.6151
R2683 B.n296 B.n295 10.6151
R2684 B.n299 B.n296 10.6151
R2685 B.n300 B.n299 10.6151
R2686 B.n303 B.n300 10.6151
R2687 B.n304 B.n303 10.6151
R2688 B.n307 B.n304 10.6151
R2689 B.n308 B.n307 10.6151
R2690 B.n311 B.n308 10.6151
R2691 B.n312 B.n311 10.6151
R2692 B.n316 B.n315 10.6151
R2693 B.n319 B.n316 10.6151
R2694 B.n320 B.n319 10.6151
R2695 B.n323 B.n320 10.6151
R2696 B.n324 B.n323 10.6151
R2697 B.n327 B.n324 10.6151
R2698 B.n328 B.n327 10.6151
R2699 B.n331 B.n328 10.6151
R2700 B.n332 B.n331 10.6151
R2701 B.n335 B.n332 10.6151
R2702 B.n336 B.n335 10.6151
R2703 B.n339 B.n336 10.6151
R2704 B.n340 B.n339 10.6151
R2705 B.n343 B.n340 10.6151
R2706 B.n344 B.n343 10.6151
R2707 B.n347 B.n344 10.6151
R2708 B.n348 B.n347 10.6151
R2709 B.n351 B.n348 10.6151
R2710 B.n352 B.n351 10.6151
R2711 B.n355 B.n352 10.6151
R2712 B.n356 B.n355 10.6151
R2713 B.n359 B.n356 10.6151
R2714 B.n360 B.n359 10.6151
R2715 B.n363 B.n360 10.6151
R2716 B.n364 B.n363 10.6151
R2717 B.n367 B.n364 10.6151
R2718 B.n368 B.n367 10.6151
R2719 B.n371 B.n368 10.6151
R2720 B.n372 B.n371 10.6151
R2721 B.n375 B.n372 10.6151
R2722 B.n376 B.n375 10.6151
R2723 B.n379 B.n376 10.6151
R2724 B.n380 B.n379 10.6151
R2725 B.n383 B.n380 10.6151
R2726 B.n384 B.n383 10.6151
R2727 B.n387 B.n384 10.6151
R2728 B.n388 B.n387 10.6151
R2729 B.n391 B.n388 10.6151
R2730 B.n392 B.n391 10.6151
R2731 B.n395 B.n392 10.6151
R2732 B.n396 B.n395 10.6151
R2733 B.n399 B.n396 10.6151
R2734 B.n400 B.n399 10.6151
R2735 B.n403 B.n400 10.6151
R2736 B.n404 B.n403 10.6151
R2737 B.n407 B.n404 10.6151
R2738 B.n408 B.n407 10.6151
R2739 B.n411 B.n408 10.6151
R2740 B.n412 B.n411 10.6151
R2741 B.n415 B.n412 10.6151
R2742 B.n416 B.n415 10.6151
R2743 B.n419 B.n416 10.6151
R2744 B.n420 B.n419 10.6151
R2745 B.n423 B.n420 10.6151
R2746 B.n424 B.n423 10.6151
R2747 B.n427 B.n424 10.6151
R2748 B.n428 B.n427 10.6151
R2749 B.n431 B.n428 10.6151
R2750 B.n432 B.n431 10.6151
R2751 B.n435 B.n432 10.6151
R2752 B.n437 B.n435 10.6151
R2753 B.n438 B.n437 10.6151
R2754 B.n1094 B.n438 10.6151
R2755 B.n886 B.n885 10.6151
R2756 B.n886 B.n526 10.6151
R2757 B.n896 B.n526 10.6151
R2758 B.n897 B.n896 10.6151
R2759 B.n898 B.n897 10.6151
R2760 B.n898 B.n517 10.6151
R2761 B.n908 B.n517 10.6151
R2762 B.n909 B.n908 10.6151
R2763 B.n910 B.n909 10.6151
R2764 B.n910 B.n510 10.6151
R2765 B.n920 B.n510 10.6151
R2766 B.n921 B.n920 10.6151
R2767 B.n922 B.n921 10.6151
R2768 B.n922 B.n502 10.6151
R2769 B.n932 B.n502 10.6151
R2770 B.n933 B.n932 10.6151
R2771 B.n934 B.n933 10.6151
R2772 B.n934 B.n494 10.6151
R2773 B.n944 B.n494 10.6151
R2774 B.n945 B.n944 10.6151
R2775 B.n946 B.n945 10.6151
R2776 B.n946 B.n486 10.6151
R2777 B.n956 B.n486 10.6151
R2778 B.n957 B.n956 10.6151
R2779 B.n958 B.n957 10.6151
R2780 B.n958 B.n478 10.6151
R2781 B.n968 B.n478 10.6151
R2782 B.n969 B.n968 10.6151
R2783 B.n970 B.n969 10.6151
R2784 B.n970 B.n469 10.6151
R2785 B.n980 B.n469 10.6151
R2786 B.n981 B.n980 10.6151
R2787 B.n982 B.n981 10.6151
R2788 B.n982 B.n462 10.6151
R2789 B.n992 B.n462 10.6151
R2790 B.n993 B.n992 10.6151
R2791 B.n994 B.n993 10.6151
R2792 B.n994 B.n454 10.6151
R2793 B.n1004 B.n454 10.6151
R2794 B.n1005 B.n1004 10.6151
R2795 B.n1006 B.n1005 10.6151
R2796 B.n1006 B.n447 10.6151
R2797 B.n1017 B.n447 10.6151
R2798 B.n1018 B.n1017 10.6151
R2799 B.n1020 B.n1018 10.6151
R2800 B.n1020 B.n1019 10.6151
R2801 B.n1019 B.n439 10.6151
R2802 B.n1031 B.n439 10.6151
R2803 B.n1032 B.n1031 10.6151
R2804 B.n1033 B.n1032 10.6151
R2805 B.n1034 B.n1033 10.6151
R2806 B.n1036 B.n1034 10.6151
R2807 B.n1037 B.n1036 10.6151
R2808 B.n1038 B.n1037 10.6151
R2809 B.n1039 B.n1038 10.6151
R2810 B.n1041 B.n1039 10.6151
R2811 B.n1042 B.n1041 10.6151
R2812 B.n1043 B.n1042 10.6151
R2813 B.n1044 B.n1043 10.6151
R2814 B.n1046 B.n1044 10.6151
R2815 B.n1047 B.n1046 10.6151
R2816 B.n1048 B.n1047 10.6151
R2817 B.n1049 B.n1048 10.6151
R2818 B.n1051 B.n1049 10.6151
R2819 B.n1052 B.n1051 10.6151
R2820 B.n1053 B.n1052 10.6151
R2821 B.n1054 B.n1053 10.6151
R2822 B.n1056 B.n1054 10.6151
R2823 B.n1057 B.n1056 10.6151
R2824 B.n1058 B.n1057 10.6151
R2825 B.n1059 B.n1058 10.6151
R2826 B.n1061 B.n1059 10.6151
R2827 B.n1062 B.n1061 10.6151
R2828 B.n1063 B.n1062 10.6151
R2829 B.n1064 B.n1063 10.6151
R2830 B.n1066 B.n1064 10.6151
R2831 B.n1067 B.n1066 10.6151
R2832 B.n1068 B.n1067 10.6151
R2833 B.n1069 B.n1068 10.6151
R2834 B.n1071 B.n1069 10.6151
R2835 B.n1072 B.n1071 10.6151
R2836 B.n1073 B.n1072 10.6151
R2837 B.n1074 B.n1073 10.6151
R2838 B.n1076 B.n1074 10.6151
R2839 B.n1077 B.n1076 10.6151
R2840 B.n1078 B.n1077 10.6151
R2841 B.n1079 B.n1078 10.6151
R2842 B.n1081 B.n1079 10.6151
R2843 B.n1082 B.n1081 10.6151
R2844 B.n1083 B.n1082 10.6151
R2845 B.n1084 B.n1083 10.6151
R2846 B.n1086 B.n1084 10.6151
R2847 B.n1087 B.n1086 10.6151
R2848 B.n1088 B.n1087 10.6151
R2849 B.n1089 B.n1088 10.6151
R2850 B.n1091 B.n1089 10.6151
R2851 B.n1092 B.n1091 10.6151
R2852 B.n1093 B.n1092 10.6151
R2853 B.n879 B.n878 10.6151
R2854 B.n878 B.n877 10.6151
R2855 B.n877 B.n876 10.6151
R2856 B.n876 B.n874 10.6151
R2857 B.n874 B.n871 10.6151
R2858 B.n871 B.n870 10.6151
R2859 B.n870 B.n867 10.6151
R2860 B.n867 B.n866 10.6151
R2861 B.n866 B.n863 10.6151
R2862 B.n863 B.n862 10.6151
R2863 B.n862 B.n859 10.6151
R2864 B.n859 B.n858 10.6151
R2865 B.n858 B.n855 10.6151
R2866 B.n855 B.n854 10.6151
R2867 B.n854 B.n851 10.6151
R2868 B.n851 B.n850 10.6151
R2869 B.n850 B.n847 10.6151
R2870 B.n847 B.n846 10.6151
R2871 B.n846 B.n843 10.6151
R2872 B.n843 B.n842 10.6151
R2873 B.n842 B.n839 10.6151
R2874 B.n839 B.n838 10.6151
R2875 B.n838 B.n835 10.6151
R2876 B.n835 B.n834 10.6151
R2877 B.n834 B.n831 10.6151
R2878 B.n831 B.n830 10.6151
R2879 B.n830 B.n827 10.6151
R2880 B.n827 B.n826 10.6151
R2881 B.n826 B.n823 10.6151
R2882 B.n823 B.n822 10.6151
R2883 B.n822 B.n819 10.6151
R2884 B.n819 B.n818 10.6151
R2885 B.n818 B.n815 10.6151
R2886 B.n815 B.n814 10.6151
R2887 B.n814 B.n811 10.6151
R2888 B.n811 B.n810 10.6151
R2889 B.n810 B.n807 10.6151
R2890 B.n807 B.n806 10.6151
R2891 B.n806 B.n803 10.6151
R2892 B.n803 B.n802 10.6151
R2893 B.n802 B.n799 10.6151
R2894 B.n799 B.n798 10.6151
R2895 B.n798 B.n795 10.6151
R2896 B.n795 B.n794 10.6151
R2897 B.n794 B.n791 10.6151
R2898 B.n791 B.n790 10.6151
R2899 B.n790 B.n787 10.6151
R2900 B.n787 B.n786 10.6151
R2901 B.n786 B.n783 10.6151
R2902 B.n783 B.n782 10.6151
R2903 B.n782 B.n779 10.6151
R2904 B.n779 B.n778 10.6151
R2905 B.n778 B.n775 10.6151
R2906 B.n775 B.n774 10.6151
R2907 B.n774 B.n771 10.6151
R2908 B.n771 B.n770 10.6151
R2909 B.n770 B.n767 10.6151
R2910 B.n767 B.n766 10.6151
R2911 B.n766 B.n763 10.6151
R2912 B.n763 B.n762 10.6151
R2913 B.n762 B.n759 10.6151
R2914 B.n759 B.n758 10.6151
R2915 B.n758 B.n755 10.6151
R2916 B.n753 B.n750 10.6151
R2917 B.n750 B.n749 10.6151
R2918 B.n749 B.n746 10.6151
R2919 B.n746 B.n745 10.6151
R2920 B.n745 B.n742 10.6151
R2921 B.n742 B.n741 10.6151
R2922 B.n741 B.n738 10.6151
R2923 B.n738 B.n737 10.6151
R2924 B.n737 B.n734 10.6151
R2925 B.n732 B.n729 10.6151
R2926 B.n729 B.n728 10.6151
R2927 B.n728 B.n725 10.6151
R2928 B.n725 B.n724 10.6151
R2929 B.n724 B.n721 10.6151
R2930 B.n721 B.n720 10.6151
R2931 B.n720 B.n717 10.6151
R2932 B.n717 B.n716 10.6151
R2933 B.n716 B.n713 10.6151
R2934 B.n713 B.n712 10.6151
R2935 B.n712 B.n709 10.6151
R2936 B.n709 B.n708 10.6151
R2937 B.n708 B.n705 10.6151
R2938 B.n705 B.n704 10.6151
R2939 B.n704 B.n701 10.6151
R2940 B.n701 B.n700 10.6151
R2941 B.n700 B.n697 10.6151
R2942 B.n697 B.n696 10.6151
R2943 B.n696 B.n693 10.6151
R2944 B.n693 B.n692 10.6151
R2945 B.n692 B.n689 10.6151
R2946 B.n689 B.n688 10.6151
R2947 B.n688 B.n685 10.6151
R2948 B.n685 B.n684 10.6151
R2949 B.n684 B.n681 10.6151
R2950 B.n681 B.n680 10.6151
R2951 B.n680 B.n677 10.6151
R2952 B.n677 B.n676 10.6151
R2953 B.n676 B.n673 10.6151
R2954 B.n673 B.n672 10.6151
R2955 B.n672 B.n669 10.6151
R2956 B.n669 B.n668 10.6151
R2957 B.n668 B.n665 10.6151
R2958 B.n665 B.n664 10.6151
R2959 B.n664 B.n661 10.6151
R2960 B.n661 B.n660 10.6151
R2961 B.n660 B.n657 10.6151
R2962 B.n657 B.n656 10.6151
R2963 B.n656 B.n653 10.6151
R2964 B.n653 B.n652 10.6151
R2965 B.n652 B.n649 10.6151
R2966 B.n649 B.n648 10.6151
R2967 B.n648 B.n645 10.6151
R2968 B.n645 B.n644 10.6151
R2969 B.n644 B.n641 10.6151
R2970 B.n641 B.n640 10.6151
R2971 B.n640 B.n637 10.6151
R2972 B.n637 B.n636 10.6151
R2973 B.n636 B.n633 10.6151
R2974 B.n633 B.n632 10.6151
R2975 B.n632 B.n629 10.6151
R2976 B.n629 B.n628 10.6151
R2977 B.n628 B.n625 10.6151
R2978 B.n625 B.n624 10.6151
R2979 B.n624 B.n621 10.6151
R2980 B.n621 B.n620 10.6151
R2981 B.n620 B.n617 10.6151
R2982 B.n617 B.n616 10.6151
R2983 B.n616 B.n613 10.6151
R2984 B.n613 B.n612 10.6151
R2985 B.n612 B.n609 10.6151
R2986 B.n609 B.n534 10.6151
R2987 B.n884 B.n534 10.6151
R2988 B.n890 B.n530 10.6151
R2989 B.n891 B.n890 10.6151
R2990 B.n892 B.n891 10.6151
R2991 B.n892 B.n522 10.6151
R2992 B.n902 B.n522 10.6151
R2993 B.n903 B.n902 10.6151
R2994 B.n904 B.n903 10.6151
R2995 B.n904 B.n514 10.6151
R2996 B.n914 B.n514 10.6151
R2997 B.n915 B.n914 10.6151
R2998 B.n916 B.n915 10.6151
R2999 B.n916 B.n506 10.6151
R3000 B.n926 B.n506 10.6151
R3001 B.n927 B.n926 10.6151
R3002 B.n928 B.n927 10.6151
R3003 B.n928 B.n498 10.6151
R3004 B.n938 B.n498 10.6151
R3005 B.n939 B.n938 10.6151
R3006 B.n940 B.n939 10.6151
R3007 B.n940 B.n490 10.6151
R3008 B.n950 B.n490 10.6151
R3009 B.n951 B.n950 10.6151
R3010 B.n952 B.n951 10.6151
R3011 B.n952 B.n482 10.6151
R3012 B.n962 B.n482 10.6151
R3013 B.n963 B.n962 10.6151
R3014 B.n964 B.n963 10.6151
R3015 B.n964 B.n474 10.6151
R3016 B.n974 B.n474 10.6151
R3017 B.n975 B.n974 10.6151
R3018 B.n976 B.n975 10.6151
R3019 B.n976 B.n466 10.6151
R3020 B.n986 B.n466 10.6151
R3021 B.n987 B.n986 10.6151
R3022 B.n988 B.n987 10.6151
R3023 B.n988 B.n458 10.6151
R3024 B.n998 B.n458 10.6151
R3025 B.n999 B.n998 10.6151
R3026 B.n1000 B.n999 10.6151
R3027 B.n1000 B.n450 10.6151
R3028 B.n1011 B.n450 10.6151
R3029 B.n1012 B.n1011 10.6151
R3030 B.n1013 B.n1012 10.6151
R3031 B.n1013 B.n443 10.6151
R3032 B.n1024 B.n443 10.6151
R3033 B.n1025 B.n1024 10.6151
R3034 B.n1026 B.n1025 10.6151
R3035 B.n1026 B.n0 10.6151
R3036 B.n1191 B.n1 10.6151
R3037 B.n1191 B.n1190 10.6151
R3038 B.n1190 B.n1189 10.6151
R3039 B.n1189 B.n10 10.6151
R3040 B.n1183 B.n10 10.6151
R3041 B.n1183 B.n1182 10.6151
R3042 B.n1182 B.n1181 10.6151
R3043 B.n1181 B.n16 10.6151
R3044 B.n1175 B.n16 10.6151
R3045 B.n1175 B.n1174 10.6151
R3046 B.n1174 B.n1173 10.6151
R3047 B.n1173 B.n24 10.6151
R3048 B.n1167 B.n24 10.6151
R3049 B.n1167 B.n1166 10.6151
R3050 B.n1166 B.n1165 10.6151
R3051 B.n1165 B.n31 10.6151
R3052 B.n1159 B.n31 10.6151
R3053 B.n1159 B.n1158 10.6151
R3054 B.n1158 B.n1157 10.6151
R3055 B.n1157 B.n38 10.6151
R3056 B.n1151 B.n38 10.6151
R3057 B.n1151 B.n1150 10.6151
R3058 B.n1150 B.n1149 10.6151
R3059 B.n1149 B.n45 10.6151
R3060 B.n1143 B.n45 10.6151
R3061 B.n1143 B.n1142 10.6151
R3062 B.n1142 B.n1141 10.6151
R3063 B.n1141 B.n52 10.6151
R3064 B.n1135 B.n52 10.6151
R3065 B.n1135 B.n1134 10.6151
R3066 B.n1134 B.n1133 10.6151
R3067 B.n1133 B.n59 10.6151
R3068 B.n1127 B.n59 10.6151
R3069 B.n1127 B.n1126 10.6151
R3070 B.n1126 B.n1125 10.6151
R3071 B.n1125 B.n66 10.6151
R3072 B.n1119 B.n66 10.6151
R3073 B.n1119 B.n1118 10.6151
R3074 B.n1118 B.n1117 10.6151
R3075 B.n1117 B.n73 10.6151
R3076 B.n1111 B.n73 10.6151
R3077 B.n1111 B.n1110 10.6151
R3078 B.n1110 B.n1109 10.6151
R3079 B.n1109 B.n80 10.6151
R3080 B.n1103 B.n80 10.6151
R3081 B.n1103 B.n1102 10.6151
R3082 B.n1102 B.n1101 10.6151
R3083 B.n1101 B.n87 10.6151
R3084 B.n292 B.n165 9.36635
R3085 B.n315 B.n162 9.36635
R3086 B.n755 B.n754 9.36635
R3087 B.n733 B.n732 9.36635
R3088 B.n1008 B.t4 9.26087
R3089 B.n18 B.t3 9.26087
R3090 B.n472 B.t0 3.96923
R3091 B.t1 B.n1162 3.96923
R3092 B.n1197 B.n0 2.81026
R3093 B.n1197 B.n1 2.81026
R3094 B.t2 B.n488 1.32341
R3095 B.t5 B.n50 1.32341
R3096 B.n295 B.n165 1.24928
R3097 B.n312 B.n162 1.24928
R3098 B.n754 B.n753 1.24928
R3099 B.n734 B.n733 1.24928
R3100 VP.n11 VP.t0 184.864
R3101 VP.n13 VP.n10 161.3
R3102 VP.n15 VP.n14 161.3
R3103 VP.n16 VP.n9 161.3
R3104 VP.n18 VP.n17 161.3
R3105 VP.n19 VP.n8 161.3
R3106 VP.n21 VP.n20 161.3
R3107 VP.n44 VP.n43 161.3
R3108 VP.n42 VP.n1 161.3
R3109 VP.n41 VP.n40 161.3
R3110 VP.n39 VP.n2 161.3
R3111 VP.n38 VP.n37 161.3
R3112 VP.n36 VP.n3 161.3
R3113 VP.n35 VP.n34 161.3
R3114 VP.n33 VP.n4 161.3
R3115 VP.n32 VP.n31 161.3
R3116 VP.n30 VP.n5 161.3
R3117 VP.n29 VP.n28 161.3
R3118 VP.n27 VP.n6 161.3
R3119 VP.n26 VP.n25 161.3
R3120 VP.n35 VP.t4 151.453
R3121 VP.n24 VP.t1 151.453
R3122 VP.n0 VP.t3 151.453
R3123 VP.n12 VP.t2 151.453
R3124 VP.n7 VP.t5 151.453
R3125 VP.n24 VP.n23 67.5578
R3126 VP.n45 VP.n0 67.5578
R3127 VP.n22 VP.n7 67.5578
R3128 VP.n23 VP.n22 56.7569
R3129 VP.n30 VP.n29 56.5193
R3130 VP.n41 VP.n2 56.5193
R3131 VP.n18 VP.n9 56.5193
R3132 VP.n12 VP.n11 49.5199
R3133 VP.n25 VP.n6 24.4675
R3134 VP.n29 VP.n6 24.4675
R3135 VP.n31 VP.n30 24.4675
R3136 VP.n31 VP.n4 24.4675
R3137 VP.n35 VP.n4 24.4675
R3138 VP.n36 VP.n35 24.4675
R3139 VP.n37 VP.n36 24.4675
R3140 VP.n37 VP.n2 24.4675
R3141 VP.n42 VP.n41 24.4675
R3142 VP.n43 VP.n42 24.4675
R3143 VP.n19 VP.n18 24.4675
R3144 VP.n20 VP.n19 24.4675
R3145 VP.n13 VP.n12 24.4675
R3146 VP.n14 VP.n13 24.4675
R3147 VP.n14 VP.n9 24.4675
R3148 VP.n25 VP.n24 22.5101
R3149 VP.n43 VP.n0 22.5101
R3150 VP.n20 VP.n7 22.5101
R3151 VP.n11 VP.n10 3.79384
R3152 VP.n22 VP.n21 0.354971
R3153 VP.n26 VP.n23 0.354971
R3154 VP.n45 VP.n44 0.354971
R3155 VP VP.n45 0.26696
R3156 VP.n15 VP.n10 0.189894
R3157 VP.n16 VP.n15 0.189894
R3158 VP.n17 VP.n16 0.189894
R3159 VP.n17 VP.n8 0.189894
R3160 VP.n21 VP.n8 0.189894
R3161 VP.n27 VP.n26 0.189894
R3162 VP.n28 VP.n27 0.189894
R3163 VP.n28 VP.n5 0.189894
R3164 VP.n32 VP.n5 0.189894
R3165 VP.n33 VP.n32 0.189894
R3166 VP.n34 VP.n33 0.189894
R3167 VP.n34 VP.n3 0.189894
R3168 VP.n38 VP.n3 0.189894
R3169 VP.n39 VP.n38 0.189894
R3170 VP.n40 VP.n39 0.189894
R3171 VP.n40 VP.n1 0.189894
R3172 VP.n44 VP.n1 0.189894
R3173 VDD1.n104 VDD1.n0 289.615
R3174 VDD1.n213 VDD1.n109 289.615
R3175 VDD1.n105 VDD1.n104 185
R3176 VDD1.n103 VDD1.n102 185
R3177 VDD1.n4 VDD1.n3 185
R3178 VDD1.n97 VDD1.n96 185
R3179 VDD1.n95 VDD1.n94 185
R3180 VDD1.n8 VDD1.n7 185
R3181 VDD1.n89 VDD1.n88 185
R3182 VDD1.n87 VDD1.n86 185
R3183 VDD1.n12 VDD1.n11 185
R3184 VDD1.n16 VDD1.n14 185
R3185 VDD1.n81 VDD1.n80 185
R3186 VDD1.n79 VDD1.n78 185
R3187 VDD1.n18 VDD1.n17 185
R3188 VDD1.n73 VDD1.n72 185
R3189 VDD1.n71 VDD1.n70 185
R3190 VDD1.n22 VDD1.n21 185
R3191 VDD1.n65 VDD1.n64 185
R3192 VDD1.n63 VDD1.n62 185
R3193 VDD1.n26 VDD1.n25 185
R3194 VDD1.n57 VDD1.n56 185
R3195 VDD1.n55 VDD1.n54 185
R3196 VDD1.n30 VDD1.n29 185
R3197 VDD1.n49 VDD1.n48 185
R3198 VDD1.n47 VDD1.n46 185
R3199 VDD1.n34 VDD1.n33 185
R3200 VDD1.n41 VDD1.n40 185
R3201 VDD1.n39 VDD1.n38 185
R3202 VDD1.n146 VDD1.n145 185
R3203 VDD1.n148 VDD1.n147 185
R3204 VDD1.n141 VDD1.n140 185
R3205 VDD1.n154 VDD1.n153 185
R3206 VDD1.n156 VDD1.n155 185
R3207 VDD1.n137 VDD1.n136 185
R3208 VDD1.n162 VDD1.n161 185
R3209 VDD1.n164 VDD1.n163 185
R3210 VDD1.n133 VDD1.n132 185
R3211 VDD1.n170 VDD1.n169 185
R3212 VDD1.n172 VDD1.n171 185
R3213 VDD1.n129 VDD1.n128 185
R3214 VDD1.n178 VDD1.n177 185
R3215 VDD1.n180 VDD1.n179 185
R3216 VDD1.n125 VDD1.n124 185
R3217 VDD1.n187 VDD1.n186 185
R3218 VDD1.n188 VDD1.n123 185
R3219 VDD1.n190 VDD1.n189 185
R3220 VDD1.n121 VDD1.n120 185
R3221 VDD1.n196 VDD1.n195 185
R3222 VDD1.n198 VDD1.n197 185
R3223 VDD1.n117 VDD1.n116 185
R3224 VDD1.n204 VDD1.n203 185
R3225 VDD1.n206 VDD1.n205 185
R3226 VDD1.n113 VDD1.n112 185
R3227 VDD1.n212 VDD1.n211 185
R3228 VDD1.n214 VDD1.n213 185
R3229 VDD1.n37 VDD1.t5 147.659
R3230 VDD1.n144 VDD1.t4 147.659
R3231 VDD1.n104 VDD1.n103 104.615
R3232 VDD1.n103 VDD1.n3 104.615
R3233 VDD1.n96 VDD1.n3 104.615
R3234 VDD1.n96 VDD1.n95 104.615
R3235 VDD1.n95 VDD1.n7 104.615
R3236 VDD1.n88 VDD1.n7 104.615
R3237 VDD1.n88 VDD1.n87 104.615
R3238 VDD1.n87 VDD1.n11 104.615
R3239 VDD1.n16 VDD1.n11 104.615
R3240 VDD1.n80 VDD1.n16 104.615
R3241 VDD1.n80 VDD1.n79 104.615
R3242 VDD1.n79 VDD1.n17 104.615
R3243 VDD1.n72 VDD1.n17 104.615
R3244 VDD1.n72 VDD1.n71 104.615
R3245 VDD1.n71 VDD1.n21 104.615
R3246 VDD1.n64 VDD1.n21 104.615
R3247 VDD1.n64 VDD1.n63 104.615
R3248 VDD1.n63 VDD1.n25 104.615
R3249 VDD1.n56 VDD1.n25 104.615
R3250 VDD1.n56 VDD1.n55 104.615
R3251 VDD1.n55 VDD1.n29 104.615
R3252 VDD1.n48 VDD1.n29 104.615
R3253 VDD1.n48 VDD1.n47 104.615
R3254 VDD1.n47 VDD1.n33 104.615
R3255 VDD1.n40 VDD1.n33 104.615
R3256 VDD1.n40 VDD1.n39 104.615
R3257 VDD1.n147 VDD1.n146 104.615
R3258 VDD1.n147 VDD1.n140 104.615
R3259 VDD1.n154 VDD1.n140 104.615
R3260 VDD1.n155 VDD1.n154 104.615
R3261 VDD1.n155 VDD1.n136 104.615
R3262 VDD1.n162 VDD1.n136 104.615
R3263 VDD1.n163 VDD1.n162 104.615
R3264 VDD1.n163 VDD1.n132 104.615
R3265 VDD1.n170 VDD1.n132 104.615
R3266 VDD1.n171 VDD1.n170 104.615
R3267 VDD1.n171 VDD1.n128 104.615
R3268 VDD1.n178 VDD1.n128 104.615
R3269 VDD1.n179 VDD1.n178 104.615
R3270 VDD1.n179 VDD1.n124 104.615
R3271 VDD1.n187 VDD1.n124 104.615
R3272 VDD1.n188 VDD1.n187 104.615
R3273 VDD1.n189 VDD1.n188 104.615
R3274 VDD1.n189 VDD1.n120 104.615
R3275 VDD1.n196 VDD1.n120 104.615
R3276 VDD1.n197 VDD1.n196 104.615
R3277 VDD1.n197 VDD1.n116 104.615
R3278 VDD1.n204 VDD1.n116 104.615
R3279 VDD1.n205 VDD1.n204 104.615
R3280 VDD1.n205 VDD1.n112 104.615
R3281 VDD1.n212 VDD1.n112 104.615
R3282 VDD1.n213 VDD1.n212 104.615
R3283 VDD1.n219 VDD1.n218 61.0984
R3284 VDD1.n221 VDD1.n220 60.408
R3285 VDD1.n221 VDD1.n219 52.4405
R3286 VDD1.n39 VDD1.t5 52.3082
R3287 VDD1.n146 VDD1.t4 52.3082
R3288 VDD1 VDD1.n108 50.9655
R3289 VDD1.n219 VDD1.n217 50.8519
R3290 VDD1.n38 VDD1.n37 15.6677
R3291 VDD1.n145 VDD1.n144 15.6677
R3292 VDD1.n14 VDD1.n12 13.1884
R3293 VDD1.n190 VDD1.n121 13.1884
R3294 VDD1.n86 VDD1.n85 12.8005
R3295 VDD1.n82 VDD1.n81 12.8005
R3296 VDD1.n41 VDD1.n36 12.8005
R3297 VDD1.n148 VDD1.n143 12.8005
R3298 VDD1.n191 VDD1.n123 12.8005
R3299 VDD1.n195 VDD1.n194 12.8005
R3300 VDD1.n89 VDD1.n10 12.0247
R3301 VDD1.n78 VDD1.n15 12.0247
R3302 VDD1.n42 VDD1.n34 12.0247
R3303 VDD1.n149 VDD1.n141 12.0247
R3304 VDD1.n186 VDD1.n185 12.0247
R3305 VDD1.n198 VDD1.n119 12.0247
R3306 VDD1.n90 VDD1.n8 11.249
R3307 VDD1.n77 VDD1.n18 11.249
R3308 VDD1.n46 VDD1.n45 11.249
R3309 VDD1.n153 VDD1.n152 11.249
R3310 VDD1.n184 VDD1.n125 11.249
R3311 VDD1.n199 VDD1.n117 11.249
R3312 VDD1.n94 VDD1.n93 10.4732
R3313 VDD1.n74 VDD1.n73 10.4732
R3314 VDD1.n49 VDD1.n32 10.4732
R3315 VDD1.n156 VDD1.n139 10.4732
R3316 VDD1.n181 VDD1.n180 10.4732
R3317 VDD1.n203 VDD1.n202 10.4732
R3318 VDD1.n97 VDD1.n6 9.69747
R3319 VDD1.n70 VDD1.n20 9.69747
R3320 VDD1.n50 VDD1.n30 9.69747
R3321 VDD1.n157 VDD1.n137 9.69747
R3322 VDD1.n177 VDD1.n127 9.69747
R3323 VDD1.n206 VDD1.n115 9.69747
R3324 VDD1.n108 VDD1.n107 9.45567
R3325 VDD1.n217 VDD1.n216 9.45567
R3326 VDD1.n24 VDD1.n23 9.3005
R3327 VDD1.n67 VDD1.n66 9.3005
R3328 VDD1.n69 VDD1.n68 9.3005
R3329 VDD1.n20 VDD1.n19 9.3005
R3330 VDD1.n75 VDD1.n74 9.3005
R3331 VDD1.n77 VDD1.n76 9.3005
R3332 VDD1.n15 VDD1.n13 9.3005
R3333 VDD1.n83 VDD1.n82 9.3005
R3334 VDD1.n107 VDD1.n106 9.3005
R3335 VDD1.n2 VDD1.n1 9.3005
R3336 VDD1.n101 VDD1.n100 9.3005
R3337 VDD1.n99 VDD1.n98 9.3005
R3338 VDD1.n6 VDD1.n5 9.3005
R3339 VDD1.n93 VDD1.n92 9.3005
R3340 VDD1.n91 VDD1.n90 9.3005
R3341 VDD1.n10 VDD1.n9 9.3005
R3342 VDD1.n85 VDD1.n84 9.3005
R3343 VDD1.n61 VDD1.n60 9.3005
R3344 VDD1.n59 VDD1.n58 9.3005
R3345 VDD1.n28 VDD1.n27 9.3005
R3346 VDD1.n53 VDD1.n52 9.3005
R3347 VDD1.n51 VDD1.n50 9.3005
R3348 VDD1.n32 VDD1.n31 9.3005
R3349 VDD1.n45 VDD1.n44 9.3005
R3350 VDD1.n43 VDD1.n42 9.3005
R3351 VDD1.n36 VDD1.n35 9.3005
R3352 VDD1.n216 VDD1.n215 9.3005
R3353 VDD1.n210 VDD1.n209 9.3005
R3354 VDD1.n208 VDD1.n207 9.3005
R3355 VDD1.n115 VDD1.n114 9.3005
R3356 VDD1.n202 VDD1.n201 9.3005
R3357 VDD1.n200 VDD1.n199 9.3005
R3358 VDD1.n119 VDD1.n118 9.3005
R3359 VDD1.n194 VDD1.n193 9.3005
R3360 VDD1.n166 VDD1.n165 9.3005
R3361 VDD1.n135 VDD1.n134 9.3005
R3362 VDD1.n160 VDD1.n159 9.3005
R3363 VDD1.n158 VDD1.n157 9.3005
R3364 VDD1.n139 VDD1.n138 9.3005
R3365 VDD1.n152 VDD1.n151 9.3005
R3366 VDD1.n150 VDD1.n149 9.3005
R3367 VDD1.n143 VDD1.n142 9.3005
R3368 VDD1.n168 VDD1.n167 9.3005
R3369 VDD1.n131 VDD1.n130 9.3005
R3370 VDD1.n174 VDD1.n173 9.3005
R3371 VDD1.n176 VDD1.n175 9.3005
R3372 VDD1.n127 VDD1.n126 9.3005
R3373 VDD1.n182 VDD1.n181 9.3005
R3374 VDD1.n184 VDD1.n183 9.3005
R3375 VDD1.n185 VDD1.n122 9.3005
R3376 VDD1.n192 VDD1.n191 9.3005
R3377 VDD1.n111 VDD1.n110 9.3005
R3378 VDD1.n98 VDD1.n4 8.92171
R3379 VDD1.n69 VDD1.n22 8.92171
R3380 VDD1.n54 VDD1.n53 8.92171
R3381 VDD1.n161 VDD1.n160 8.92171
R3382 VDD1.n176 VDD1.n129 8.92171
R3383 VDD1.n207 VDD1.n113 8.92171
R3384 VDD1.n102 VDD1.n101 8.14595
R3385 VDD1.n66 VDD1.n65 8.14595
R3386 VDD1.n57 VDD1.n28 8.14595
R3387 VDD1.n164 VDD1.n135 8.14595
R3388 VDD1.n173 VDD1.n172 8.14595
R3389 VDD1.n211 VDD1.n210 8.14595
R3390 VDD1.n108 VDD1.n0 7.3702
R3391 VDD1.n105 VDD1.n2 7.3702
R3392 VDD1.n62 VDD1.n24 7.3702
R3393 VDD1.n58 VDD1.n26 7.3702
R3394 VDD1.n165 VDD1.n133 7.3702
R3395 VDD1.n169 VDD1.n131 7.3702
R3396 VDD1.n214 VDD1.n111 7.3702
R3397 VDD1.n217 VDD1.n109 7.3702
R3398 VDD1.n106 VDD1.n0 6.59444
R3399 VDD1.n106 VDD1.n105 6.59444
R3400 VDD1.n62 VDD1.n61 6.59444
R3401 VDD1.n61 VDD1.n26 6.59444
R3402 VDD1.n168 VDD1.n133 6.59444
R3403 VDD1.n169 VDD1.n168 6.59444
R3404 VDD1.n215 VDD1.n214 6.59444
R3405 VDD1.n215 VDD1.n109 6.59444
R3406 VDD1.n102 VDD1.n2 5.81868
R3407 VDD1.n65 VDD1.n24 5.81868
R3408 VDD1.n58 VDD1.n57 5.81868
R3409 VDD1.n165 VDD1.n164 5.81868
R3410 VDD1.n172 VDD1.n131 5.81868
R3411 VDD1.n211 VDD1.n111 5.81868
R3412 VDD1.n101 VDD1.n4 5.04292
R3413 VDD1.n66 VDD1.n22 5.04292
R3414 VDD1.n54 VDD1.n28 5.04292
R3415 VDD1.n161 VDD1.n135 5.04292
R3416 VDD1.n173 VDD1.n129 5.04292
R3417 VDD1.n210 VDD1.n113 5.04292
R3418 VDD1.n37 VDD1.n35 4.38563
R3419 VDD1.n144 VDD1.n142 4.38563
R3420 VDD1.n98 VDD1.n97 4.26717
R3421 VDD1.n70 VDD1.n69 4.26717
R3422 VDD1.n53 VDD1.n30 4.26717
R3423 VDD1.n160 VDD1.n137 4.26717
R3424 VDD1.n177 VDD1.n176 4.26717
R3425 VDD1.n207 VDD1.n206 4.26717
R3426 VDD1.n94 VDD1.n6 3.49141
R3427 VDD1.n73 VDD1.n20 3.49141
R3428 VDD1.n50 VDD1.n49 3.49141
R3429 VDD1.n157 VDD1.n156 3.49141
R3430 VDD1.n180 VDD1.n127 3.49141
R3431 VDD1.n203 VDD1.n115 3.49141
R3432 VDD1.n93 VDD1.n8 2.71565
R3433 VDD1.n74 VDD1.n18 2.71565
R3434 VDD1.n46 VDD1.n32 2.71565
R3435 VDD1.n153 VDD1.n139 2.71565
R3436 VDD1.n181 VDD1.n125 2.71565
R3437 VDD1.n202 VDD1.n117 2.71565
R3438 VDD1.n90 VDD1.n89 1.93989
R3439 VDD1.n78 VDD1.n77 1.93989
R3440 VDD1.n45 VDD1.n34 1.93989
R3441 VDD1.n152 VDD1.n141 1.93989
R3442 VDD1.n186 VDD1.n184 1.93989
R3443 VDD1.n199 VDD1.n198 1.93989
R3444 VDD1.n86 VDD1.n10 1.16414
R3445 VDD1.n81 VDD1.n15 1.16414
R3446 VDD1.n42 VDD1.n41 1.16414
R3447 VDD1.n149 VDD1.n148 1.16414
R3448 VDD1.n185 VDD1.n123 1.16414
R3449 VDD1.n195 VDD1.n119 1.16414
R3450 VDD1.n220 VDD1.t3 1.00711
R3451 VDD1.n220 VDD1.t0 1.00711
R3452 VDD1.n218 VDD1.t1 1.00711
R3453 VDD1.n218 VDD1.t2 1.00711
R3454 VDD1 VDD1.n221 0.688
R3455 VDD1.n85 VDD1.n12 0.388379
R3456 VDD1.n82 VDD1.n14 0.388379
R3457 VDD1.n38 VDD1.n36 0.388379
R3458 VDD1.n145 VDD1.n143 0.388379
R3459 VDD1.n191 VDD1.n190 0.388379
R3460 VDD1.n194 VDD1.n121 0.388379
R3461 VDD1.n107 VDD1.n1 0.155672
R3462 VDD1.n100 VDD1.n1 0.155672
R3463 VDD1.n100 VDD1.n99 0.155672
R3464 VDD1.n99 VDD1.n5 0.155672
R3465 VDD1.n92 VDD1.n5 0.155672
R3466 VDD1.n92 VDD1.n91 0.155672
R3467 VDD1.n91 VDD1.n9 0.155672
R3468 VDD1.n84 VDD1.n9 0.155672
R3469 VDD1.n84 VDD1.n83 0.155672
R3470 VDD1.n83 VDD1.n13 0.155672
R3471 VDD1.n76 VDD1.n13 0.155672
R3472 VDD1.n76 VDD1.n75 0.155672
R3473 VDD1.n75 VDD1.n19 0.155672
R3474 VDD1.n68 VDD1.n19 0.155672
R3475 VDD1.n68 VDD1.n67 0.155672
R3476 VDD1.n67 VDD1.n23 0.155672
R3477 VDD1.n60 VDD1.n23 0.155672
R3478 VDD1.n60 VDD1.n59 0.155672
R3479 VDD1.n59 VDD1.n27 0.155672
R3480 VDD1.n52 VDD1.n27 0.155672
R3481 VDD1.n52 VDD1.n51 0.155672
R3482 VDD1.n51 VDD1.n31 0.155672
R3483 VDD1.n44 VDD1.n31 0.155672
R3484 VDD1.n44 VDD1.n43 0.155672
R3485 VDD1.n43 VDD1.n35 0.155672
R3486 VDD1.n150 VDD1.n142 0.155672
R3487 VDD1.n151 VDD1.n150 0.155672
R3488 VDD1.n151 VDD1.n138 0.155672
R3489 VDD1.n158 VDD1.n138 0.155672
R3490 VDD1.n159 VDD1.n158 0.155672
R3491 VDD1.n159 VDD1.n134 0.155672
R3492 VDD1.n166 VDD1.n134 0.155672
R3493 VDD1.n167 VDD1.n166 0.155672
R3494 VDD1.n167 VDD1.n130 0.155672
R3495 VDD1.n174 VDD1.n130 0.155672
R3496 VDD1.n175 VDD1.n174 0.155672
R3497 VDD1.n175 VDD1.n126 0.155672
R3498 VDD1.n182 VDD1.n126 0.155672
R3499 VDD1.n183 VDD1.n182 0.155672
R3500 VDD1.n183 VDD1.n122 0.155672
R3501 VDD1.n192 VDD1.n122 0.155672
R3502 VDD1.n193 VDD1.n192 0.155672
R3503 VDD1.n193 VDD1.n118 0.155672
R3504 VDD1.n200 VDD1.n118 0.155672
R3505 VDD1.n201 VDD1.n200 0.155672
R3506 VDD1.n201 VDD1.n114 0.155672
R3507 VDD1.n208 VDD1.n114 0.155672
R3508 VDD1.n209 VDD1.n208 0.155672
R3509 VDD1.n209 VDD1.n110 0.155672
R3510 VDD1.n216 VDD1.n110 0.155672
C0 VDD1 VDD2 1.61505f
C1 VN VTAIL 11.0683f
C2 VP VDD1 11.4818f
C3 VP VDD2 0.503873f
C4 VN VDD1 0.151553f
C5 VN VDD2 11.1337f
C6 VTAIL VDD1 10.4728f
C7 VTAIL VDD2 10.5262f
C8 VN VP 8.86057f
C9 VTAIL VP 11.0826f
C10 VDD2 B 7.753998f
C11 VDD1 B 7.907286f
C12 VTAIL B 11.277824f
C13 VN B 15.06955f
C14 VP B 13.636726f
C15 VDD1.n0 B 0.031009f
C16 VDD1.n1 B 0.021344f
C17 VDD1.n2 B 0.011469f
C18 VDD1.n3 B 0.027109f
C19 VDD1.n4 B 0.012144f
C20 VDD1.n5 B 0.021344f
C21 VDD1.n6 B 0.011469f
C22 VDD1.n7 B 0.027109f
C23 VDD1.n8 B 0.012144f
C24 VDD1.n9 B 0.021344f
C25 VDD1.n10 B 0.011469f
C26 VDD1.n11 B 0.027109f
C27 VDD1.n12 B 0.011807f
C28 VDD1.n13 B 0.021344f
C29 VDD1.n14 B 0.011807f
C30 VDD1.n15 B 0.011469f
C31 VDD1.n16 B 0.027109f
C32 VDD1.n17 B 0.027109f
C33 VDD1.n18 B 0.012144f
C34 VDD1.n19 B 0.021344f
C35 VDD1.n20 B 0.011469f
C36 VDD1.n21 B 0.027109f
C37 VDD1.n22 B 0.012144f
C38 VDD1.n23 B 0.021344f
C39 VDD1.n24 B 0.011469f
C40 VDD1.n25 B 0.027109f
C41 VDD1.n26 B 0.012144f
C42 VDD1.n27 B 0.021344f
C43 VDD1.n28 B 0.011469f
C44 VDD1.n29 B 0.027109f
C45 VDD1.n30 B 0.012144f
C46 VDD1.n31 B 0.021344f
C47 VDD1.n32 B 0.011469f
C48 VDD1.n33 B 0.027109f
C49 VDD1.n34 B 0.012144f
C50 VDD1.n35 B 1.84549f
C51 VDD1.n36 B 0.011469f
C52 VDD1.t5 B 0.045042f
C53 VDD1.n37 B 0.164201f
C54 VDD1.n38 B 0.016014f
C55 VDD1.n39 B 0.020332f
C56 VDD1.n40 B 0.027109f
C57 VDD1.n41 B 0.012144f
C58 VDD1.n42 B 0.011469f
C59 VDD1.n43 B 0.021344f
C60 VDD1.n44 B 0.021344f
C61 VDD1.n45 B 0.011469f
C62 VDD1.n46 B 0.012144f
C63 VDD1.n47 B 0.027109f
C64 VDD1.n48 B 0.027109f
C65 VDD1.n49 B 0.012144f
C66 VDD1.n50 B 0.011469f
C67 VDD1.n51 B 0.021344f
C68 VDD1.n52 B 0.021344f
C69 VDD1.n53 B 0.011469f
C70 VDD1.n54 B 0.012144f
C71 VDD1.n55 B 0.027109f
C72 VDD1.n56 B 0.027109f
C73 VDD1.n57 B 0.012144f
C74 VDD1.n58 B 0.011469f
C75 VDD1.n59 B 0.021344f
C76 VDD1.n60 B 0.021344f
C77 VDD1.n61 B 0.011469f
C78 VDD1.n62 B 0.012144f
C79 VDD1.n63 B 0.027109f
C80 VDD1.n64 B 0.027109f
C81 VDD1.n65 B 0.012144f
C82 VDD1.n66 B 0.011469f
C83 VDD1.n67 B 0.021344f
C84 VDD1.n68 B 0.021344f
C85 VDD1.n69 B 0.011469f
C86 VDD1.n70 B 0.012144f
C87 VDD1.n71 B 0.027109f
C88 VDD1.n72 B 0.027109f
C89 VDD1.n73 B 0.012144f
C90 VDD1.n74 B 0.011469f
C91 VDD1.n75 B 0.021344f
C92 VDD1.n76 B 0.021344f
C93 VDD1.n77 B 0.011469f
C94 VDD1.n78 B 0.012144f
C95 VDD1.n79 B 0.027109f
C96 VDD1.n80 B 0.027109f
C97 VDD1.n81 B 0.012144f
C98 VDD1.n82 B 0.011469f
C99 VDD1.n83 B 0.021344f
C100 VDD1.n84 B 0.021344f
C101 VDD1.n85 B 0.011469f
C102 VDD1.n86 B 0.012144f
C103 VDD1.n87 B 0.027109f
C104 VDD1.n88 B 0.027109f
C105 VDD1.n89 B 0.012144f
C106 VDD1.n90 B 0.011469f
C107 VDD1.n91 B 0.021344f
C108 VDD1.n92 B 0.021344f
C109 VDD1.n93 B 0.011469f
C110 VDD1.n94 B 0.012144f
C111 VDD1.n95 B 0.027109f
C112 VDD1.n96 B 0.027109f
C113 VDD1.n97 B 0.012144f
C114 VDD1.n98 B 0.011469f
C115 VDD1.n99 B 0.021344f
C116 VDD1.n100 B 0.021344f
C117 VDD1.n101 B 0.011469f
C118 VDD1.n102 B 0.012144f
C119 VDD1.n103 B 0.027109f
C120 VDD1.n104 B 0.06047f
C121 VDD1.n105 B 0.012144f
C122 VDD1.n106 B 0.011469f
C123 VDD1.n107 B 0.049044f
C124 VDD1.n108 B 0.057702f
C125 VDD1.n109 B 0.031009f
C126 VDD1.n110 B 0.021344f
C127 VDD1.n111 B 0.011469f
C128 VDD1.n112 B 0.027109f
C129 VDD1.n113 B 0.012144f
C130 VDD1.n114 B 0.021344f
C131 VDD1.n115 B 0.011469f
C132 VDD1.n116 B 0.027109f
C133 VDD1.n117 B 0.012144f
C134 VDD1.n118 B 0.021344f
C135 VDD1.n119 B 0.011469f
C136 VDD1.n120 B 0.027109f
C137 VDD1.n121 B 0.011807f
C138 VDD1.n122 B 0.021344f
C139 VDD1.n123 B 0.012144f
C140 VDD1.n124 B 0.027109f
C141 VDD1.n125 B 0.012144f
C142 VDD1.n126 B 0.021344f
C143 VDD1.n127 B 0.011469f
C144 VDD1.n128 B 0.027109f
C145 VDD1.n129 B 0.012144f
C146 VDD1.n130 B 0.021344f
C147 VDD1.n131 B 0.011469f
C148 VDD1.n132 B 0.027109f
C149 VDD1.n133 B 0.012144f
C150 VDD1.n134 B 0.021344f
C151 VDD1.n135 B 0.011469f
C152 VDD1.n136 B 0.027109f
C153 VDD1.n137 B 0.012144f
C154 VDD1.n138 B 0.021344f
C155 VDD1.n139 B 0.011469f
C156 VDD1.n140 B 0.027109f
C157 VDD1.n141 B 0.012144f
C158 VDD1.n142 B 1.84549f
C159 VDD1.n143 B 0.011469f
C160 VDD1.t4 B 0.045042f
C161 VDD1.n144 B 0.164201f
C162 VDD1.n145 B 0.016014f
C163 VDD1.n146 B 0.020332f
C164 VDD1.n147 B 0.027109f
C165 VDD1.n148 B 0.012144f
C166 VDD1.n149 B 0.011469f
C167 VDD1.n150 B 0.021344f
C168 VDD1.n151 B 0.021344f
C169 VDD1.n152 B 0.011469f
C170 VDD1.n153 B 0.012144f
C171 VDD1.n154 B 0.027109f
C172 VDD1.n155 B 0.027109f
C173 VDD1.n156 B 0.012144f
C174 VDD1.n157 B 0.011469f
C175 VDD1.n158 B 0.021344f
C176 VDD1.n159 B 0.021344f
C177 VDD1.n160 B 0.011469f
C178 VDD1.n161 B 0.012144f
C179 VDD1.n162 B 0.027109f
C180 VDD1.n163 B 0.027109f
C181 VDD1.n164 B 0.012144f
C182 VDD1.n165 B 0.011469f
C183 VDD1.n166 B 0.021344f
C184 VDD1.n167 B 0.021344f
C185 VDD1.n168 B 0.011469f
C186 VDD1.n169 B 0.012144f
C187 VDD1.n170 B 0.027109f
C188 VDD1.n171 B 0.027109f
C189 VDD1.n172 B 0.012144f
C190 VDD1.n173 B 0.011469f
C191 VDD1.n174 B 0.021344f
C192 VDD1.n175 B 0.021344f
C193 VDD1.n176 B 0.011469f
C194 VDD1.n177 B 0.012144f
C195 VDD1.n178 B 0.027109f
C196 VDD1.n179 B 0.027109f
C197 VDD1.n180 B 0.012144f
C198 VDD1.n181 B 0.011469f
C199 VDD1.n182 B 0.021344f
C200 VDD1.n183 B 0.021344f
C201 VDD1.n184 B 0.011469f
C202 VDD1.n185 B 0.011469f
C203 VDD1.n186 B 0.012144f
C204 VDD1.n187 B 0.027109f
C205 VDD1.n188 B 0.027109f
C206 VDD1.n189 B 0.027109f
C207 VDD1.n190 B 0.011807f
C208 VDD1.n191 B 0.011469f
C209 VDD1.n192 B 0.021344f
C210 VDD1.n193 B 0.021344f
C211 VDD1.n194 B 0.011469f
C212 VDD1.n195 B 0.012144f
C213 VDD1.n196 B 0.027109f
C214 VDD1.n197 B 0.027109f
C215 VDD1.n198 B 0.012144f
C216 VDD1.n199 B 0.011469f
C217 VDD1.n200 B 0.021344f
C218 VDD1.n201 B 0.021344f
C219 VDD1.n202 B 0.011469f
C220 VDD1.n203 B 0.012144f
C221 VDD1.n204 B 0.027109f
C222 VDD1.n205 B 0.027109f
C223 VDD1.n206 B 0.012144f
C224 VDD1.n207 B 0.011469f
C225 VDD1.n208 B 0.021344f
C226 VDD1.n209 B 0.021344f
C227 VDD1.n210 B 0.011469f
C228 VDD1.n211 B 0.012144f
C229 VDD1.n212 B 0.027109f
C230 VDD1.n213 B 0.06047f
C231 VDD1.n214 B 0.012144f
C232 VDD1.n215 B 0.011469f
C233 VDD1.n216 B 0.049044f
C234 VDD1.n217 B 0.056953f
C235 VDD1.t1 B 0.331767f
C236 VDD1.t2 B 0.331767f
C237 VDD1.n218 B 3.03694f
C238 VDD1.n219 B 3.01888f
C239 VDD1.t3 B 0.331767f
C240 VDD1.t0 B 0.331767f
C241 VDD1.n220 B 3.03195f
C242 VDD1.n221 B 3.00581f
C243 VP.t3 B 3.33694f
C244 VP.n0 B 1.23393f
C245 VP.n1 B 0.019674f
C246 VP.n2 B 0.027623f
C247 VP.n3 B 0.019674f
C248 VP.t4 B 3.33694f
C249 VP.n4 B 0.036666f
C250 VP.n5 B 0.019674f
C251 VP.n6 B 0.036666f
C252 VP.t5 B 3.33694f
C253 VP.n7 B 1.23393f
C254 VP.n8 B 0.019674f
C255 VP.n9 B 0.027623f
C256 VP.n10 B 0.223676f
C257 VP.t2 B 3.33694f
C258 VP.t0 B 3.5706f
C259 VP.n11 B 1.17536f
C260 VP.n12 B 1.22404f
C261 VP.n13 B 0.036666f
C262 VP.n14 B 0.036666f
C263 VP.n15 B 0.019674f
C264 VP.n16 B 0.019674f
C265 VP.n17 B 0.019674f
C266 VP.n18 B 0.029816f
C267 VP.n19 B 0.036666f
C268 VP.n20 B 0.035218f
C269 VP.n21 B 0.031753f
C270 VP.n22 B 1.32919f
C271 VP.n23 B 1.34165f
C272 VP.t1 B 3.33694f
C273 VP.n24 B 1.23393f
C274 VP.n25 B 0.035218f
C275 VP.n26 B 0.031753f
C276 VP.n27 B 0.019674f
C277 VP.n28 B 0.019674f
C278 VP.n29 B 0.029816f
C279 VP.n30 B 0.027623f
C280 VP.n31 B 0.036666f
C281 VP.n32 B 0.019674f
C282 VP.n33 B 0.019674f
C283 VP.n34 B 0.019674f
C284 VP.n35 B 1.16815f
C285 VP.n36 B 0.036666f
C286 VP.n37 B 0.036666f
C287 VP.n38 B 0.019674f
C288 VP.n39 B 0.019674f
C289 VP.n40 B 0.019674f
C290 VP.n41 B 0.029816f
C291 VP.n42 B 0.036666f
C292 VP.n43 B 0.035218f
C293 VP.n44 B 0.031753f
C294 VP.n45 B 0.039307f
C295 VTAIL.t9 B 0.349856f
C296 VTAIL.t10 B 0.349856f
C297 VTAIL.n0 B 3.12683f
C298 VTAIL.n1 B 0.429321f
C299 VTAIL.n2 B 0.0327f
C300 VTAIL.n3 B 0.022508f
C301 VTAIL.n4 B 0.012095f
C302 VTAIL.n5 B 0.028587f
C303 VTAIL.n6 B 0.012806f
C304 VTAIL.n7 B 0.022508f
C305 VTAIL.n8 B 0.012095f
C306 VTAIL.n9 B 0.028587f
C307 VTAIL.n10 B 0.012806f
C308 VTAIL.n11 B 0.022508f
C309 VTAIL.n12 B 0.012095f
C310 VTAIL.n13 B 0.028587f
C311 VTAIL.n14 B 0.01245f
C312 VTAIL.n15 B 0.022508f
C313 VTAIL.n16 B 0.012806f
C314 VTAIL.n17 B 0.028587f
C315 VTAIL.n18 B 0.012806f
C316 VTAIL.n19 B 0.022508f
C317 VTAIL.n20 B 0.012095f
C318 VTAIL.n21 B 0.028587f
C319 VTAIL.n22 B 0.012806f
C320 VTAIL.n23 B 0.022508f
C321 VTAIL.n24 B 0.012095f
C322 VTAIL.n25 B 0.028587f
C323 VTAIL.n26 B 0.012806f
C324 VTAIL.n27 B 0.022508f
C325 VTAIL.n28 B 0.012095f
C326 VTAIL.n29 B 0.028587f
C327 VTAIL.n30 B 0.012806f
C328 VTAIL.n31 B 0.022508f
C329 VTAIL.n32 B 0.012095f
C330 VTAIL.n33 B 0.028587f
C331 VTAIL.n34 B 0.012806f
C332 VTAIL.n35 B 1.94611f
C333 VTAIL.n36 B 0.012095f
C334 VTAIL.t4 B 0.047498f
C335 VTAIL.n37 B 0.173154f
C336 VTAIL.n38 B 0.016887f
C337 VTAIL.n39 B 0.021441f
C338 VTAIL.n40 B 0.028587f
C339 VTAIL.n41 B 0.012806f
C340 VTAIL.n42 B 0.012095f
C341 VTAIL.n43 B 0.022508f
C342 VTAIL.n44 B 0.022508f
C343 VTAIL.n45 B 0.012095f
C344 VTAIL.n46 B 0.012806f
C345 VTAIL.n47 B 0.028587f
C346 VTAIL.n48 B 0.028587f
C347 VTAIL.n49 B 0.012806f
C348 VTAIL.n50 B 0.012095f
C349 VTAIL.n51 B 0.022508f
C350 VTAIL.n52 B 0.022508f
C351 VTAIL.n53 B 0.012095f
C352 VTAIL.n54 B 0.012806f
C353 VTAIL.n55 B 0.028587f
C354 VTAIL.n56 B 0.028587f
C355 VTAIL.n57 B 0.012806f
C356 VTAIL.n58 B 0.012095f
C357 VTAIL.n59 B 0.022508f
C358 VTAIL.n60 B 0.022508f
C359 VTAIL.n61 B 0.012095f
C360 VTAIL.n62 B 0.012806f
C361 VTAIL.n63 B 0.028587f
C362 VTAIL.n64 B 0.028587f
C363 VTAIL.n65 B 0.012806f
C364 VTAIL.n66 B 0.012095f
C365 VTAIL.n67 B 0.022508f
C366 VTAIL.n68 B 0.022508f
C367 VTAIL.n69 B 0.012095f
C368 VTAIL.n70 B 0.012806f
C369 VTAIL.n71 B 0.028587f
C370 VTAIL.n72 B 0.028587f
C371 VTAIL.n73 B 0.012806f
C372 VTAIL.n74 B 0.012095f
C373 VTAIL.n75 B 0.022508f
C374 VTAIL.n76 B 0.022508f
C375 VTAIL.n77 B 0.012095f
C376 VTAIL.n78 B 0.012095f
C377 VTAIL.n79 B 0.012806f
C378 VTAIL.n80 B 0.028587f
C379 VTAIL.n81 B 0.028587f
C380 VTAIL.n82 B 0.028587f
C381 VTAIL.n83 B 0.01245f
C382 VTAIL.n84 B 0.012095f
C383 VTAIL.n85 B 0.022508f
C384 VTAIL.n86 B 0.022508f
C385 VTAIL.n87 B 0.012095f
C386 VTAIL.n88 B 0.012806f
C387 VTAIL.n89 B 0.028587f
C388 VTAIL.n90 B 0.028587f
C389 VTAIL.n91 B 0.012806f
C390 VTAIL.n92 B 0.012095f
C391 VTAIL.n93 B 0.022508f
C392 VTAIL.n94 B 0.022508f
C393 VTAIL.n95 B 0.012095f
C394 VTAIL.n96 B 0.012806f
C395 VTAIL.n97 B 0.028587f
C396 VTAIL.n98 B 0.028587f
C397 VTAIL.n99 B 0.012806f
C398 VTAIL.n100 B 0.012095f
C399 VTAIL.n101 B 0.022508f
C400 VTAIL.n102 B 0.022508f
C401 VTAIL.n103 B 0.012095f
C402 VTAIL.n104 B 0.012806f
C403 VTAIL.n105 B 0.028587f
C404 VTAIL.n106 B 0.063767f
C405 VTAIL.n107 B 0.012806f
C406 VTAIL.n108 B 0.012095f
C407 VTAIL.n109 B 0.051718f
C408 VTAIL.n110 B 0.035864f
C409 VTAIL.n111 B 0.37761f
C410 VTAIL.t2 B 0.349856f
C411 VTAIL.t0 B 0.349856f
C412 VTAIL.n112 B 3.12683f
C413 VTAIL.n113 B 2.41329f
C414 VTAIL.t7 B 0.349856f
C415 VTAIL.t11 B 0.349856f
C416 VTAIL.n114 B 3.12684f
C417 VTAIL.n115 B 2.41328f
C418 VTAIL.n116 B 0.0327f
C419 VTAIL.n117 B 0.022508f
C420 VTAIL.n118 B 0.012095f
C421 VTAIL.n119 B 0.028587f
C422 VTAIL.n120 B 0.012806f
C423 VTAIL.n121 B 0.022508f
C424 VTAIL.n122 B 0.012095f
C425 VTAIL.n123 B 0.028587f
C426 VTAIL.n124 B 0.012806f
C427 VTAIL.n125 B 0.022508f
C428 VTAIL.n126 B 0.012095f
C429 VTAIL.n127 B 0.028587f
C430 VTAIL.n128 B 0.01245f
C431 VTAIL.n129 B 0.022508f
C432 VTAIL.n130 B 0.01245f
C433 VTAIL.n131 B 0.012095f
C434 VTAIL.n132 B 0.028587f
C435 VTAIL.n133 B 0.028587f
C436 VTAIL.n134 B 0.012806f
C437 VTAIL.n135 B 0.022508f
C438 VTAIL.n136 B 0.012095f
C439 VTAIL.n137 B 0.028587f
C440 VTAIL.n138 B 0.012806f
C441 VTAIL.n139 B 0.022508f
C442 VTAIL.n140 B 0.012095f
C443 VTAIL.n141 B 0.028587f
C444 VTAIL.n142 B 0.012806f
C445 VTAIL.n143 B 0.022508f
C446 VTAIL.n144 B 0.012095f
C447 VTAIL.n145 B 0.028587f
C448 VTAIL.n146 B 0.012806f
C449 VTAIL.n147 B 0.022508f
C450 VTAIL.n148 B 0.012095f
C451 VTAIL.n149 B 0.028587f
C452 VTAIL.n150 B 0.012806f
C453 VTAIL.n151 B 1.94611f
C454 VTAIL.n152 B 0.012095f
C455 VTAIL.t8 B 0.047498f
C456 VTAIL.n153 B 0.173154f
C457 VTAIL.n154 B 0.016887f
C458 VTAIL.n155 B 0.021441f
C459 VTAIL.n156 B 0.028587f
C460 VTAIL.n157 B 0.012806f
C461 VTAIL.n158 B 0.012095f
C462 VTAIL.n159 B 0.022508f
C463 VTAIL.n160 B 0.022508f
C464 VTAIL.n161 B 0.012095f
C465 VTAIL.n162 B 0.012806f
C466 VTAIL.n163 B 0.028587f
C467 VTAIL.n164 B 0.028587f
C468 VTAIL.n165 B 0.012806f
C469 VTAIL.n166 B 0.012095f
C470 VTAIL.n167 B 0.022508f
C471 VTAIL.n168 B 0.022508f
C472 VTAIL.n169 B 0.012095f
C473 VTAIL.n170 B 0.012806f
C474 VTAIL.n171 B 0.028587f
C475 VTAIL.n172 B 0.028587f
C476 VTAIL.n173 B 0.012806f
C477 VTAIL.n174 B 0.012095f
C478 VTAIL.n175 B 0.022508f
C479 VTAIL.n176 B 0.022508f
C480 VTAIL.n177 B 0.012095f
C481 VTAIL.n178 B 0.012806f
C482 VTAIL.n179 B 0.028587f
C483 VTAIL.n180 B 0.028587f
C484 VTAIL.n181 B 0.012806f
C485 VTAIL.n182 B 0.012095f
C486 VTAIL.n183 B 0.022508f
C487 VTAIL.n184 B 0.022508f
C488 VTAIL.n185 B 0.012095f
C489 VTAIL.n186 B 0.012806f
C490 VTAIL.n187 B 0.028587f
C491 VTAIL.n188 B 0.028587f
C492 VTAIL.n189 B 0.012806f
C493 VTAIL.n190 B 0.012095f
C494 VTAIL.n191 B 0.022508f
C495 VTAIL.n192 B 0.022508f
C496 VTAIL.n193 B 0.012095f
C497 VTAIL.n194 B 0.012806f
C498 VTAIL.n195 B 0.028587f
C499 VTAIL.n196 B 0.028587f
C500 VTAIL.n197 B 0.012806f
C501 VTAIL.n198 B 0.012095f
C502 VTAIL.n199 B 0.022508f
C503 VTAIL.n200 B 0.022508f
C504 VTAIL.n201 B 0.012095f
C505 VTAIL.n202 B 0.012806f
C506 VTAIL.n203 B 0.028587f
C507 VTAIL.n204 B 0.028587f
C508 VTAIL.n205 B 0.012806f
C509 VTAIL.n206 B 0.012095f
C510 VTAIL.n207 B 0.022508f
C511 VTAIL.n208 B 0.022508f
C512 VTAIL.n209 B 0.012095f
C513 VTAIL.n210 B 0.012806f
C514 VTAIL.n211 B 0.028587f
C515 VTAIL.n212 B 0.028587f
C516 VTAIL.n213 B 0.012806f
C517 VTAIL.n214 B 0.012095f
C518 VTAIL.n215 B 0.022508f
C519 VTAIL.n216 B 0.022508f
C520 VTAIL.n217 B 0.012095f
C521 VTAIL.n218 B 0.012806f
C522 VTAIL.n219 B 0.028587f
C523 VTAIL.n220 B 0.063767f
C524 VTAIL.n221 B 0.012806f
C525 VTAIL.n222 B 0.012095f
C526 VTAIL.n223 B 0.051718f
C527 VTAIL.n224 B 0.035864f
C528 VTAIL.n225 B 0.37761f
C529 VTAIL.t3 B 0.349856f
C530 VTAIL.t1 B 0.349856f
C531 VTAIL.n226 B 3.12684f
C532 VTAIL.n227 B 0.587331f
C533 VTAIL.n228 B 0.0327f
C534 VTAIL.n229 B 0.022508f
C535 VTAIL.n230 B 0.012095f
C536 VTAIL.n231 B 0.028587f
C537 VTAIL.n232 B 0.012806f
C538 VTAIL.n233 B 0.022508f
C539 VTAIL.n234 B 0.012095f
C540 VTAIL.n235 B 0.028587f
C541 VTAIL.n236 B 0.012806f
C542 VTAIL.n237 B 0.022508f
C543 VTAIL.n238 B 0.012095f
C544 VTAIL.n239 B 0.028587f
C545 VTAIL.n240 B 0.01245f
C546 VTAIL.n241 B 0.022508f
C547 VTAIL.n242 B 0.01245f
C548 VTAIL.n243 B 0.012095f
C549 VTAIL.n244 B 0.028587f
C550 VTAIL.n245 B 0.028587f
C551 VTAIL.n246 B 0.012806f
C552 VTAIL.n247 B 0.022508f
C553 VTAIL.n248 B 0.012095f
C554 VTAIL.n249 B 0.028587f
C555 VTAIL.n250 B 0.012806f
C556 VTAIL.n251 B 0.022508f
C557 VTAIL.n252 B 0.012095f
C558 VTAIL.n253 B 0.028587f
C559 VTAIL.n254 B 0.012806f
C560 VTAIL.n255 B 0.022508f
C561 VTAIL.n256 B 0.012095f
C562 VTAIL.n257 B 0.028587f
C563 VTAIL.n258 B 0.012806f
C564 VTAIL.n259 B 0.022508f
C565 VTAIL.n260 B 0.012095f
C566 VTAIL.n261 B 0.028587f
C567 VTAIL.n262 B 0.012806f
C568 VTAIL.n263 B 1.94611f
C569 VTAIL.n264 B 0.012095f
C570 VTAIL.t5 B 0.047498f
C571 VTAIL.n265 B 0.173154f
C572 VTAIL.n266 B 0.016887f
C573 VTAIL.n267 B 0.021441f
C574 VTAIL.n268 B 0.028587f
C575 VTAIL.n269 B 0.012806f
C576 VTAIL.n270 B 0.012095f
C577 VTAIL.n271 B 0.022508f
C578 VTAIL.n272 B 0.022508f
C579 VTAIL.n273 B 0.012095f
C580 VTAIL.n274 B 0.012806f
C581 VTAIL.n275 B 0.028587f
C582 VTAIL.n276 B 0.028587f
C583 VTAIL.n277 B 0.012806f
C584 VTAIL.n278 B 0.012095f
C585 VTAIL.n279 B 0.022508f
C586 VTAIL.n280 B 0.022508f
C587 VTAIL.n281 B 0.012095f
C588 VTAIL.n282 B 0.012806f
C589 VTAIL.n283 B 0.028587f
C590 VTAIL.n284 B 0.028587f
C591 VTAIL.n285 B 0.012806f
C592 VTAIL.n286 B 0.012095f
C593 VTAIL.n287 B 0.022508f
C594 VTAIL.n288 B 0.022508f
C595 VTAIL.n289 B 0.012095f
C596 VTAIL.n290 B 0.012806f
C597 VTAIL.n291 B 0.028587f
C598 VTAIL.n292 B 0.028587f
C599 VTAIL.n293 B 0.012806f
C600 VTAIL.n294 B 0.012095f
C601 VTAIL.n295 B 0.022508f
C602 VTAIL.n296 B 0.022508f
C603 VTAIL.n297 B 0.012095f
C604 VTAIL.n298 B 0.012806f
C605 VTAIL.n299 B 0.028587f
C606 VTAIL.n300 B 0.028587f
C607 VTAIL.n301 B 0.012806f
C608 VTAIL.n302 B 0.012095f
C609 VTAIL.n303 B 0.022508f
C610 VTAIL.n304 B 0.022508f
C611 VTAIL.n305 B 0.012095f
C612 VTAIL.n306 B 0.012806f
C613 VTAIL.n307 B 0.028587f
C614 VTAIL.n308 B 0.028587f
C615 VTAIL.n309 B 0.012806f
C616 VTAIL.n310 B 0.012095f
C617 VTAIL.n311 B 0.022508f
C618 VTAIL.n312 B 0.022508f
C619 VTAIL.n313 B 0.012095f
C620 VTAIL.n314 B 0.012806f
C621 VTAIL.n315 B 0.028587f
C622 VTAIL.n316 B 0.028587f
C623 VTAIL.n317 B 0.012806f
C624 VTAIL.n318 B 0.012095f
C625 VTAIL.n319 B 0.022508f
C626 VTAIL.n320 B 0.022508f
C627 VTAIL.n321 B 0.012095f
C628 VTAIL.n322 B 0.012806f
C629 VTAIL.n323 B 0.028587f
C630 VTAIL.n324 B 0.028587f
C631 VTAIL.n325 B 0.012806f
C632 VTAIL.n326 B 0.012095f
C633 VTAIL.n327 B 0.022508f
C634 VTAIL.n328 B 0.022508f
C635 VTAIL.n329 B 0.012095f
C636 VTAIL.n330 B 0.012806f
C637 VTAIL.n331 B 0.028587f
C638 VTAIL.n332 B 0.063767f
C639 VTAIL.n333 B 0.012806f
C640 VTAIL.n334 B 0.012095f
C641 VTAIL.n335 B 0.051718f
C642 VTAIL.n336 B 0.035864f
C643 VTAIL.n337 B 1.98724f
C644 VTAIL.n338 B 0.0327f
C645 VTAIL.n339 B 0.022508f
C646 VTAIL.n340 B 0.012095f
C647 VTAIL.n341 B 0.028587f
C648 VTAIL.n342 B 0.012806f
C649 VTAIL.n343 B 0.022508f
C650 VTAIL.n344 B 0.012095f
C651 VTAIL.n345 B 0.028587f
C652 VTAIL.n346 B 0.012806f
C653 VTAIL.n347 B 0.022508f
C654 VTAIL.n348 B 0.012095f
C655 VTAIL.n349 B 0.028587f
C656 VTAIL.n350 B 0.01245f
C657 VTAIL.n351 B 0.022508f
C658 VTAIL.n352 B 0.012806f
C659 VTAIL.n353 B 0.028587f
C660 VTAIL.n354 B 0.012806f
C661 VTAIL.n355 B 0.022508f
C662 VTAIL.n356 B 0.012095f
C663 VTAIL.n357 B 0.028587f
C664 VTAIL.n358 B 0.012806f
C665 VTAIL.n359 B 0.022508f
C666 VTAIL.n360 B 0.012095f
C667 VTAIL.n361 B 0.028587f
C668 VTAIL.n362 B 0.012806f
C669 VTAIL.n363 B 0.022508f
C670 VTAIL.n364 B 0.012095f
C671 VTAIL.n365 B 0.028587f
C672 VTAIL.n366 B 0.012806f
C673 VTAIL.n367 B 0.022508f
C674 VTAIL.n368 B 0.012095f
C675 VTAIL.n369 B 0.028587f
C676 VTAIL.n370 B 0.012806f
C677 VTAIL.n371 B 1.94611f
C678 VTAIL.n372 B 0.012095f
C679 VTAIL.t6 B 0.047498f
C680 VTAIL.n373 B 0.173154f
C681 VTAIL.n374 B 0.016887f
C682 VTAIL.n375 B 0.021441f
C683 VTAIL.n376 B 0.028587f
C684 VTAIL.n377 B 0.012806f
C685 VTAIL.n378 B 0.012095f
C686 VTAIL.n379 B 0.022508f
C687 VTAIL.n380 B 0.022508f
C688 VTAIL.n381 B 0.012095f
C689 VTAIL.n382 B 0.012806f
C690 VTAIL.n383 B 0.028587f
C691 VTAIL.n384 B 0.028587f
C692 VTAIL.n385 B 0.012806f
C693 VTAIL.n386 B 0.012095f
C694 VTAIL.n387 B 0.022508f
C695 VTAIL.n388 B 0.022508f
C696 VTAIL.n389 B 0.012095f
C697 VTAIL.n390 B 0.012806f
C698 VTAIL.n391 B 0.028587f
C699 VTAIL.n392 B 0.028587f
C700 VTAIL.n393 B 0.012806f
C701 VTAIL.n394 B 0.012095f
C702 VTAIL.n395 B 0.022508f
C703 VTAIL.n396 B 0.022508f
C704 VTAIL.n397 B 0.012095f
C705 VTAIL.n398 B 0.012806f
C706 VTAIL.n399 B 0.028587f
C707 VTAIL.n400 B 0.028587f
C708 VTAIL.n401 B 0.012806f
C709 VTAIL.n402 B 0.012095f
C710 VTAIL.n403 B 0.022508f
C711 VTAIL.n404 B 0.022508f
C712 VTAIL.n405 B 0.012095f
C713 VTAIL.n406 B 0.012806f
C714 VTAIL.n407 B 0.028587f
C715 VTAIL.n408 B 0.028587f
C716 VTAIL.n409 B 0.012806f
C717 VTAIL.n410 B 0.012095f
C718 VTAIL.n411 B 0.022508f
C719 VTAIL.n412 B 0.022508f
C720 VTAIL.n413 B 0.012095f
C721 VTAIL.n414 B 0.012095f
C722 VTAIL.n415 B 0.012806f
C723 VTAIL.n416 B 0.028587f
C724 VTAIL.n417 B 0.028587f
C725 VTAIL.n418 B 0.028587f
C726 VTAIL.n419 B 0.01245f
C727 VTAIL.n420 B 0.012095f
C728 VTAIL.n421 B 0.022508f
C729 VTAIL.n422 B 0.022508f
C730 VTAIL.n423 B 0.012095f
C731 VTAIL.n424 B 0.012806f
C732 VTAIL.n425 B 0.028587f
C733 VTAIL.n426 B 0.028587f
C734 VTAIL.n427 B 0.012806f
C735 VTAIL.n428 B 0.012095f
C736 VTAIL.n429 B 0.022508f
C737 VTAIL.n430 B 0.022508f
C738 VTAIL.n431 B 0.012095f
C739 VTAIL.n432 B 0.012806f
C740 VTAIL.n433 B 0.028587f
C741 VTAIL.n434 B 0.028587f
C742 VTAIL.n435 B 0.012806f
C743 VTAIL.n436 B 0.012095f
C744 VTAIL.n437 B 0.022508f
C745 VTAIL.n438 B 0.022508f
C746 VTAIL.n439 B 0.012095f
C747 VTAIL.n440 B 0.012806f
C748 VTAIL.n441 B 0.028587f
C749 VTAIL.n442 B 0.063767f
C750 VTAIL.n443 B 0.012806f
C751 VTAIL.n444 B 0.012095f
C752 VTAIL.n445 B 0.051718f
C753 VTAIL.n446 B 0.035864f
C754 VTAIL.n447 B 1.92893f
C755 VDD2.n0 B 0.030555f
C756 VDD2.n1 B 0.021031f
C757 VDD2.n2 B 0.011301f
C758 VDD2.n3 B 0.026712f
C759 VDD2.n4 B 0.011966f
C760 VDD2.n5 B 0.021031f
C761 VDD2.n6 B 0.011301f
C762 VDD2.n7 B 0.026712f
C763 VDD2.n8 B 0.011966f
C764 VDD2.n9 B 0.021031f
C765 VDD2.n10 B 0.011301f
C766 VDD2.n11 B 0.026712f
C767 VDD2.n12 B 0.011634f
C768 VDD2.n13 B 0.021031f
C769 VDD2.n14 B 0.011966f
C770 VDD2.n15 B 0.026712f
C771 VDD2.n16 B 0.011966f
C772 VDD2.n17 B 0.021031f
C773 VDD2.n18 B 0.011301f
C774 VDD2.n19 B 0.026712f
C775 VDD2.n20 B 0.011966f
C776 VDD2.n21 B 0.021031f
C777 VDD2.n22 B 0.011301f
C778 VDD2.n23 B 0.026712f
C779 VDD2.n24 B 0.011966f
C780 VDD2.n25 B 0.021031f
C781 VDD2.n26 B 0.011301f
C782 VDD2.n27 B 0.026712f
C783 VDD2.n28 B 0.011966f
C784 VDD2.n29 B 0.021031f
C785 VDD2.n30 B 0.011301f
C786 VDD2.n31 B 0.026712f
C787 VDD2.n32 B 0.011966f
C788 VDD2.n33 B 1.81845f
C789 VDD2.n34 B 0.011301f
C790 VDD2.t3 B 0.044382f
C791 VDD2.n35 B 0.161796f
C792 VDD2.n36 B 0.01578f
C793 VDD2.n37 B 0.020034f
C794 VDD2.n38 B 0.026712f
C795 VDD2.n39 B 0.011966f
C796 VDD2.n40 B 0.011301f
C797 VDD2.n41 B 0.021031f
C798 VDD2.n42 B 0.021031f
C799 VDD2.n43 B 0.011301f
C800 VDD2.n44 B 0.011966f
C801 VDD2.n45 B 0.026712f
C802 VDD2.n46 B 0.026712f
C803 VDD2.n47 B 0.011966f
C804 VDD2.n48 B 0.011301f
C805 VDD2.n49 B 0.021031f
C806 VDD2.n50 B 0.021031f
C807 VDD2.n51 B 0.011301f
C808 VDD2.n52 B 0.011966f
C809 VDD2.n53 B 0.026712f
C810 VDD2.n54 B 0.026712f
C811 VDD2.n55 B 0.011966f
C812 VDD2.n56 B 0.011301f
C813 VDD2.n57 B 0.021031f
C814 VDD2.n58 B 0.021031f
C815 VDD2.n59 B 0.011301f
C816 VDD2.n60 B 0.011966f
C817 VDD2.n61 B 0.026712f
C818 VDD2.n62 B 0.026712f
C819 VDD2.n63 B 0.011966f
C820 VDD2.n64 B 0.011301f
C821 VDD2.n65 B 0.021031f
C822 VDD2.n66 B 0.021031f
C823 VDD2.n67 B 0.011301f
C824 VDD2.n68 B 0.011966f
C825 VDD2.n69 B 0.026712f
C826 VDD2.n70 B 0.026712f
C827 VDD2.n71 B 0.011966f
C828 VDD2.n72 B 0.011301f
C829 VDD2.n73 B 0.021031f
C830 VDD2.n74 B 0.021031f
C831 VDD2.n75 B 0.011301f
C832 VDD2.n76 B 0.011301f
C833 VDD2.n77 B 0.011966f
C834 VDD2.n78 B 0.026712f
C835 VDD2.n79 B 0.026712f
C836 VDD2.n80 B 0.026712f
C837 VDD2.n81 B 0.011634f
C838 VDD2.n82 B 0.011301f
C839 VDD2.n83 B 0.021031f
C840 VDD2.n84 B 0.021031f
C841 VDD2.n85 B 0.011301f
C842 VDD2.n86 B 0.011966f
C843 VDD2.n87 B 0.026712f
C844 VDD2.n88 B 0.026712f
C845 VDD2.n89 B 0.011966f
C846 VDD2.n90 B 0.011301f
C847 VDD2.n91 B 0.021031f
C848 VDD2.n92 B 0.021031f
C849 VDD2.n93 B 0.011301f
C850 VDD2.n94 B 0.011966f
C851 VDD2.n95 B 0.026712f
C852 VDD2.n96 B 0.026712f
C853 VDD2.n97 B 0.011966f
C854 VDD2.n98 B 0.011301f
C855 VDD2.n99 B 0.021031f
C856 VDD2.n100 B 0.021031f
C857 VDD2.n101 B 0.011301f
C858 VDD2.n102 B 0.011966f
C859 VDD2.n103 B 0.026712f
C860 VDD2.n104 B 0.059584f
C861 VDD2.n105 B 0.011966f
C862 VDD2.n106 B 0.011301f
C863 VDD2.n107 B 0.048325f
C864 VDD2.n108 B 0.056118f
C865 VDD2.t1 B 0.326907f
C866 VDD2.t2 B 0.326907f
C867 VDD2.n109 B 2.99244f
C868 VDD2.n110 B 2.85389f
C869 VDD2.n111 B 0.030555f
C870 VDD2.n112 B 0.021031f
C871 VDD2.n113 B 0.011301f
C872 VDD2.n114 B 0.026712f
C873 VDD2.n115 B 0.011966f
C874 VDD2.n116 B 0.021031f
C875 VDD2.n117 B 0.011301f
C876 VDD2.n118 B 0.026712f
C877 VDD2.n119 B 0.011966f
C878 VDD2.n120 B 0.021031f
C879 VDD2.n121 B 0.011301f
C880 VDD2.n122 B 0.026712f
C881 VDD2.n123 B 0.011634f
C882 VDD2.n124 B 0.021031f
C883 VDD2.n125 B 0.011634f
C884 VDD2.n126 B 0.011301f
C885 VDD2.n127 B 0.026712f
C886 VDD2.n128 B 0.026712f
C887 VDD2.n129 B 0.011966f
C888 VDD2.n130 B 0.021031f
C889 VDD2.n131 B 0.011301f
C890 VDD2.n132 B 0.026712f
C891 VDD2.n133 B 0.011966f
C892 VDD2.n134 B 0.021031f
C893 VDD2.n135 B 0.011301f
C894 VDD2.n136 B 0.026712f
C895 VDD2.n137 B 0.011966f
C896 VDD2.n138 B 0.021031f
C897 VDD2.n139 B 0.011301f
C898 VDD2.n140 B 0.026712f
C899 VDD2.n141 B 0.011966f
C900 VDD2.n142 B 0.021031f
C901 VDD2.n143 B 0.011301f
C902 VDD2.n144 B 0.026712f
C903 VDD2.n145 B 0.011966f
C904 VDD2.n146 B 1.81845f
C905 VDD2.n147 B 0.011301f
C906 VDD2.t0 B 0.044382f
C907 VDD2.n148 B 0.161796f
C908 VDD2.n149 B 0.01578f
C909 VDD2.n150 B 0.020034f
C910 VDD2.n151 B 0.026712f
C911 VDD2.n152 B 0.011966f
C912 VDD2.n153 B 0.011301f
C913 VDD2.n154 B 0.021031f
C914 VDD2.n155 B 0.021031f
C915 VDD2.n156 B 0.011301f
C916 VDD2.n157 B 0.011966f
C917 VDD2.n158 B 0.026712f
C918 VDD2.n159 B 0.026712f
C919 VDD2.n160 B 0.011966f
C920 VDD2.n161 B 0.011301f
C921 VDD2.n162 B 0.021031f
C922 VDD2.n163 B 0.021031f
C923 VDD2.n164 B 0.011301f
C924 VDD2.n165 B 0.011966f
C925 VDD2.n166 B 0.026712f
C926 VDD2.n167 B 0.026712f
C927 VDD2.n168 B 0.011966f
C928 VDD2.n169 B 0.011301f
C929 VDD2.n170 B 0.021031f
C930 VDD2.n171 B 0.021031f
C931 VDD2.n172 B 0.011301f
C932 VDD2.n173 B 0.011966f
C933 VDD2.n174 B 0.026712f
C934 VDD2.n175 B 0.026712f
C935 VDD2.n176 B 0.011966f
C936 VDD2.n177 B 0.011301f
C937 VDD2.n178 B 0.021031f
C938 VDD2.n179 B 0.021031f
C939 VDD2.n180 B 0.011301f
C940 VDD2.n181 B 0.011966f
C941 VDD2.n182 B 0.026712f
C942 VDD2.n183 B 0.026712f
C943 VDD2.n184 B 0.011966f
C944 VDD2.n185 B 0.011301f
C945 VDD2.n186 B 0.021031f
C946 VDD2.n187 B 0.021031f
C947 VDD2.n188 B 0.011301f
C948 VDD2.n189 B 0.011966f
C949 VDD2.n190 B 0.026712f
C950 VDD2.n191 B 0.026712f
C951 VDD2.n192 B 0.011966f
C952 VDD2.n193 B 0.011301f
C953 VDD2.n194 B 0.021031f
C954 VDD2.n195 B 0.021031f
C955 VDD2.n196 B 0.011301f
C956 VDD2.n197 B 0.011966f
C957 VDD2.n198 B 0.026712f
C958 VDD2.n199 B 0.026712f
C959 VDD2.n200 B 0.011966f
C960 VDD2.n201 B 0.011301f
C961 VDD2.n202 B 0.021031f
C962 VDD2.n203 B 0.021031f
C963 VDD2.n204 B 0.011301f
C964 VDD2.n205 B 0.011966f
C965 VDD2.n206 B 0.026712f
C966 VDD2.n207 B 0.026712f
C967 VDD2.n208 B 0.011966f
C968 VDD2.n209 B 0.011301f
C969 VDD2.n210 B 0.021031f
C970 VDD2.n211 B 0.021031f
C971 VDD2.n212 B 0.011301f
C972 VDD2.n213 B 0.011966f
C973 VDD2.n214 B 0.026712f
C974 VDD2.n215 B 0.059584f
C975 VDD2.n216 B 0.011966f
C976 VDD2.n217 B 0.011301f
C977 VDD2.n218 B 0.048325f
C978 VDD2.n219 B 0.048035f
C979 VDD2.n220 B 2.76699f
C980 VDD2.t5 B 0.326907f
C981 VDD2.t4 B 0.326907f
C982 VDD2.n221 B 2.99241f
C983 VN.t5 B 3.29167f
C984 VN.n0 B 1.21719f
C985 VN.n1 B 0.019407f
C986 VN.n2 B 0.027249f
C987 VN.n3 B 0.220641f
C988 VN.t1 B 3.29167f
C989 VN.t2 B 3.52216f
C990 VN.n4 B 1.15942f
C991 VN.n5 B 1.20743f
C992 VN.n6 B 0.036169f
C993 VN.n7 B 0.036169f
C994 VN.n8 B 0.019407f
C995 VN.n9 B 0.019407f
C996 VN.n10 B 0.019407f
C997 VN.n11 B 0.029412f
C998 VN.n12 B 0.036169f
C999 VN.n13 B 0.034741f
C1000 VN.n14 B 0.031322f
C1001 VN.n15 B 0.038774f
C1002 VN.t4 B 3.29167f
C1003 VN.n16 B 1.21719f
C1004 VN.n17 B 0.019407f
C1005 VN.n18 B 0.027249f
C1006 VN.n19 B 0.220641f
C1007 VN.t0 B 3.29167f
C1008 VN.t3 B 3.52216f
C1009 VN.n20 B 1.15942f
C1010 VN.n21 B 1.20743f
C1011 VN.n22 B 0.036169f
C1012 VN.n23 B 0.036169f
C1013 VN.n24 B 0.019407f
C1014 VN.n25 B 0.019407f
C1015 VN.n26 B 0.019407f
C1016 VN.n27 B 0.029412f
C1017 VN.n28 B 0.036169f
C1018 VN.n29 B 0.034741f
C1019 VN.n30 B 0.031322f
C1020 VN.n31 B 1.31877f
.ends

