* NGSPICE file created from diff_pair_sample_0242.ext - technology: sky130A

.subckt diff_pair_sample_0242 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t3 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=2.2308 ps=12.22 w=5.72 l=1.76
X1 B.t21 B.t19 B.t20 B.t16 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0 ps=0 w=5.72 l=1.76
X2 VDD2.t7 VN.t0 VTAIL.t12 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=2.2308 ps=12.22 w=5.72 l=1.76
X3 VTAIL.t11 VN.t1 VDD2.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0.9438 ps=6.05 w=5.72 l=1.76
X4 B.t18 B.t15 B.t17 B.t16 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0 ps=0 w=5.72 l=1.76
X5 VTAIL.t13 VN.t2 VDD2.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X6 VDD2.t4 VN.t3 VTAIL.t15 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X7 VTAIL.t7 VP.t1 VDD1.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0.9438 ps=6.05 w=5.72 l=1.76
X8 VDD2.t3 VN.t4 VTAIL.t14 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X9 VTAIL.t10 VN.t5 VDD2.t2 B.t6 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0.9438 ps=6.05 w=5.72 l=1.76
X10 VTAIL.t8 VN.t6 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X11 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0 ps=0 w=5.72 l=1.76
X12 VDD2.t0 VN.t7 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=2.2308 ps=12.22 w=5.72 l=1.76
X13 VTAIL.t5 VP.t2 VDD1.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0.9438 ps=6.05 w=5.72 l=1.76
X14 VDD1.t4 VP.t3 VTAIL.t0 B.t4 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=2.2308 ps=12.22 w=5.72 l=1.76
X15 VTAIL.t6 VP.t4 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X16 VDD1.t2 VP.t5 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X17 VTAIL.t2 VP.t6 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X18 VDD1.t0 VP.t7 VTAIL.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=0.9438 pd=6.05 as=0.9438 ps=6.05 w=5.72 l=1.76
X19 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=2.2308 pd=12.22 as=0 ps=0 w=5.72 l=1.76
R0 VP.n31 VP.n30 179.252
R1 VP.n54 VP.n53 179.252
R2 VP.n29 VP.n28 179.252
R3 VP.n14 VP.n11 161.3
R4 VP.n16 VP.n15 161.3
R5 VP.n17 VP.n10 161.3
R6 VP.n19 VP.n18 161.3
R7 VP.n20 VP.n9 161.3
R8 VP.n23 VP.n22 161.3
R9 VP.n24 VP.n8 161.3
R10 VP.n26 VP.n25 161.3
R11 VP.n27 VP.n7 161.3
R12 VP.n52 VP.n0 161.3
R13 VP.n51 VP.n50 161.3
R14 VP.n49 VP.n1 161.3
R15 VP.n48 VP.n47 161.3
R16 VP.n45 VP.n2 161.3
R17 VP.n44 VP.n43 161.3
R18 VP.n42 VP.n3 161.3
R19 VP.n41 VP.n40 161.3
R20 VP.n39 VP.n4 161.3
R21 VP.n37 VP.n36 161.3
R22 VP.n35 VP.n5 161.3
R23 VP.n34 VP.n33 161.3
R24 VP.n32 VP.n6 161.3
R25 VP.n12 VP.t2 109.865
R26 VP.n31 VP.t1 78.3255
R27 VP.n38 VP.t5 78.3255
R28 VP.n46 VP.t4 78.3255
R29 VP.n53 VP.t0 78.3255
R30 VP.n28 VP.t3 78.3255
R31 VP.n21 VP.t6 78.3255
R32 VP.n13 VP.t7 78.3255
R33 VP.n13 VP.n12 65.8068
R34 VP.n33 VP.n5 49.296
R35 VP.n51 VP.n1 49.296
R36 VP.n26 VP.n8 49.296
R37 VP.n30 VP.n29 42.1444
R38 VP.n40 VP.n3 40.577
R39 VP.n44 VP.n3 40.577
R40 VP.n19 VP.n10 40.577
R41 VP.n15 VP.n10 40.577
R42 VP.n37 VP.n5 31.8581
R43 VP.n47 VP.n1 31.8581
R44 VP.n22 VP.n8 31.8581
R45 VP.n33 VP.n32 24.5923
R46 VP.n40 VP.n39 24.5923
R47 VP.n45 VP.n44 24.5923
R48 VP.n52 VP.n51 24.5923
R49 VP.n27 VP.n26 24.5923
R50 VP.n20 VP.n19 24.5923
R51 VP.n15 VP.n14 24.5923
R52 VP.n38 VP.n37 22.3791
R53 VP.n47 VP.n46 22.3791
R54 VP.n22 VP.n21 22.3791
R55 VP.n12 VP.n11 18.2204
R56 VP.n32 VP.n31 6.6403
R57 VP.n53 VP.n52 6.6403
R58 VP.n28 VP.n27 6.6403
R59 VP.n39 VP.n38 2.21377
R60 VP.n46 VP.n45 2.21377
R61 VP.n21 VP.n20 2.21377
R62 VP.n14 VP.n13 2.21377
R63 VP.n16 VP.n11 0.189894
R64 VP.n17 VP.n16 0.189894
R65 VP.n18 VP.n17 0.189894
R66 VP.n18 VP.n9 0.189894
R67 VP.n23 VP.n9 0.189894
R68 VP.n24 VP.n23 0.189894
R69 VP.n25 VP.n24 0.189894
R70 VP.n25 VP.n7 0.189894
R71 VP.n29 VP.n7 0.189894
R72 VP.n30 VP.n6 0.189894
R73 VP.n34 VP.n6 0.189894
R74 VP.n35 VP.n34 0.189894
R75 VP.n36 VP.n35 0.189894
R76 VP.n36 VP.n4 0.189894
R77 VP.n41 VP.n4 0.189894
R78 VP.n42 VP.n41 0.189894
R79 VP.n43 VP.n42 0.189894
R80 VP.n43 VP.n2 0.189894
R81 VP.n48 VP.n2 0.189894
R82 VP.n49 VP.n48 0.189894
R83 VP.n50 VP.n49 0.189894
R84 VP.n50 VP.n0 0.189894
R85 VP.n54 VP.n0 0.189894
R86 VP VP.n54 0.0516364
R87 VTAIL.n11 VTAIL.t5 56.2043
R88 VTAIL.n10 VTAIL.t9 56.2043
R89 VTAIL.n7 VTAIL.t10 56.2043
R90 VTAIL.n15 VTAIL.t12 56.2041
R91 VTAIL.n2 VTAIL.t11 56.2041
R92 VTAIL.n3 VTAIL.t3 56.2041
R93 VTAIL.n6 VTAIL.t7 56.2041
R94 VTAIL.n14 VTAIL.t0 56.2041
R95 VTAIL.n13 VTAIL.n12 52.7427
R96 VTAIL.n9 VTAIL.n8 52.7427
R97 VTAIL.n1 VTAIL.n0 52.7425
R98 VTAIL.n5 VTAIL.n4 52.7425
R99 VTAIL.n15 VTAIL.n14 19.0996
R100 VTAIL.n7 VTAIL.n6 19.0996
R101 VTAIL.n0 VTAIL.t15 3.46204
R102 VTAIL.n0 VTAIL.t13 3.46204
R103 VTAIL.n4 VTAIL.t4 3.46204
R104 VTAIL.n4 VTAIL.t6 3.46204
R105 VTAIL.n12 VTAIL.t1 3.46204
R106 VTAIL.n12 VTAIL.t2 3.46204
R107 VTAIL.n8 VTAIL.t14 3.46204
R108 VTAIL.n8 VTAIL.t8 3.46204
R109 VTAIL.n9 VTAIL.n7 1.80222
R110 VTAIL.n10 VTAIL.n9 1.80222
R111 VTAIL.n13 VTAIL.n11 1.80222
R112 VTAIL.n14 VTAIL.n13 1.80222
R113 VTAIL.n6 VTAIL.n5 1.80222
R114 VTAIL.n5 VTAIL.n3 1.80222
R115 VTAIL.n2 VTAIL.n1 1.80222
R116 VTAIL VTAIL.n15 1.74403
R117 VTAIL.n11 VTAIL.n10 0.470328
R118 VTAIL.n3 VTAIL.n2 0.470328
R119 VTAIL VTAIL.n1 0.0586897
R120 VDD1 VDD1.n0 70.3806
R121 VDD1.n3 VDD1.n2 70.2668
R122 VDD1.n3 VDD1.n1 70.2668
R123 VDD1.n5 VDD1.n4 69.4214
R124 VDD1.n5 VDD1.n3 37.3371
R125 VDD1.n4 VDD1.t1 3.46204
R126 VDD1.n4 VDD1.t4 3.46204
R127 VDD1.n0 VDD1.t5 3.46204
R128 VDD1.n0 VDD1.t0 3.46204
R129 VDD1.n2 VDD1.t3 3.46204
R130 VDD1.n2 VDD1.t7 3.46204
R131 VDD1.n1 VDD1.t6 3.46204
R132 VDD1.n1 VDD1.t2 3.46204
R133 VDD1 VDD1.n5 0.843172
R134 B.n602 B.n601 585
R135 B.n213 B.n101 585
R136 B.n212 B.n211 585
R137 B.n210 B.n209 585
R138 B.n208 B.n207 585
R139 B.n206 B.n205 585
R140 B.n204 B.n203 585
R141 B.n202 B.n201 585
R142 B.n200 B.n199 585
R143 B.n198 B.n197 585
R144 B.n196 B.n195 585
R145 B.n194 B.n193 585
R146 B.n192 B.n191 585
R147 B.n190 B.n189 585
R148 B.n188 B.n187 585
R149 B.n186 B.n185 585
R150 B.n184 B.n183 585
R151 B.n182 B.n181 585
R152 B.n180 B.n179 585
R153 B.n178 B.n177 585
R154 B.n176 B.n175 585
R155 B.n174 B.n173 585
R156 B.n172 B.n171 585
R157 B.n169 B.n168 585
R158 B.n167 B.n166 585
R159 B.n165 B.n164 585
R160 B.n163 B.n162 585
R161 B.n161 B.n160 585
R162 B.n159 B.n158 585
R163 B.n157 B.n156 585
R164 B.n155 B.n154 585
R165 B.n153 B.n152 585
R166 B.n151 B.n150 585
R167 B.n148 B.n147 585
R168 B.n146 B.n145 585
R169 B.n144 B.n143 585
R170 B.n142 B.n141 585
R171 B.n140 B.n139 585
R172 B.n138 B.n137 585
R173 B.n136 B.n135 585
R174 B.n134 B.n133 585
R175 B.n132 B.n131 585
R176 B.n130 B.n129 585
R177 B.n128 B.n127 585
R178 B.n126 B.n125 585
R179 B.n124 B.n123 585
R180 B.n122 B.n121 585
R181 B.n120 B.n119 585
R182 B.n118 B.n117 585
R183 B.n116 B.n115 585
R184 B.n114 B.n113 585
R185 B.n112 B.n111 585
R186 B.n110 B.n109 585
R187 B.n108 B.n107 585
R188 B.n74 B.n73 585
R189 B.n607 B.n606 585
R190 B.n600 B.n102 585
R191 B.n102 B.n71 585
R192 B.n599 B.n70 585
R193 B.n611 B.n70 585
R194 B.n598 B.n69 585
R195 B.n612 B.n69 585
R196 B.n597 B.n68 585
R197 B.n613 B.n68 585
R198 B.n596 B.n595 585
R199 B.n595 B.n64 585
R200 B.n594 B.n63 585
R201 B.n619 B.n63 585
R202 B.n593 B.n62 585
R203 B.n620 B.n62 585
R204 B.n592 B.n61 585
R205 B.n621 B.n61 585
R206 B.n591 B.n590 585
R207 B.n590 B.n57 585
R208 B.n589 B.n56 585
R209 B.n627 B.n56 585
R210 B.n588 B.n55 585
R211 B.n628 B.n55 585
R212 B.n587 B.n54 585
R213 B.n629 B.n54 585
R214 B.n586 B.n585 585
R215 B.n585 B.n50 585
R216 B.n584 B.n49 585
R217 B.n635 B.n49 585
R218 B.n583 B.n48 585
R219 B.n636 B.n48 585
R220 B.n582 B.n47 585
R221 B.n637 B.n47 585
R222 B.n581 B.n580 585
R223 B.n580 B.n43 585
R224 B.n579 B.n42 585
R225 B.n643 B.n42 585
R226 B.n578 B.n41 585
R227 B.n644 B.n41 585
R228 B.n577 B.n40 585
R229 B.n645 B.n40 585
R230 B.n576 B.n575 585
R231 B.n575 B.n36 585
R232 B.n574 B.n35 585
R233 B.n651 B.n35 585
R234 B.n573 B.n34 585
R235 B.n652 B.n34 585
R236 B.n572 B.n33 585
R237 B.n653 B.n33 585
R238 B.n571 B.n570 585
R239 B.n570 B.n29 585
R240 B.n569 B.n28 585
R241 B.n659 B.n28 585
R242 B.n568 B.n27 585
R243 B.n660 B.n27 585
R244 B.n567 B.n26 585
R245 B.n661 B.n26 585
R246 B.n566 B.n565 585
R247 B.n565 B.n25 585
R248 B.n564 B.n21 585
R249 B.n667 B.n21 585
R250 B.n563 B.n20 585
R251 B.n668 B.n20 585
R252 B.n562 B.n19 585
R253 B.n669 B.n19 585
R254 B.n561 B.n560 585
R255 B.n560 B.n15 585
R256 B.n559 B.n14 585
R257 B.n675 B.n14 585
R258 B.n558 B.n13 585
R259 B.n676 B.n13 585
R260 B.n557 B.n12 585
R261 B.n677 B.n12 585
R262 B.n556 B.n555 585
R263 B.n555 B.n8 585
R264 B.n554 B.n7 585
R265 B.n683 B.n7 585
R266 B.n553 B.n6 585
R267 B.n684 B.n6 585
R268 B.n552 B.n5 585
R269 B.n685 B.n5 585
R270 B.n551 B.n550 585
R271 B.n550 B.n4 585
R272 B.n549 B.n214 585
R273 B.n549 B.n548 585
R274 B.n539 B.n215 585
R275 B.n216 B.n215 585
R276 B.n541 B.n540 585
R277 B.n542 B.n541 585
R278 B.n538 B.n220 585
R279 B.n224 B.n220 585
R280 B.n537 B.n536 585
R281 B.n536 B.n535 585
R282 B.n222 B.n221 585
R283 B.n223 B.n222 585
R284 B.n528 B.n527 585
R285 B.n529 B.n528 585
R286 B.n526 B.n229 585
R287 B.n229 B.n228 585
R288 B.n525 B.n524 585
R289 B.n524 B.n523 585
R290 B.n231 B.n230 585
R291 B.n516 B.n231 585
R292 B.n515 B.n514 585
R293 B.n517 B.n515 585
R294 B.n513 B.n236 585
R295 B.n236 B.n235 585
R296 B.n512 B.n511 585
R297 B.n511 B.n510 585
R298 B.n238 B.n237 585
R299 B.n239 B.n238 585
R300 B.n503 B.n502 585
R301 B.n504 B.n503 585
R302 B.n501 B.n243 585
R303 B.n247 B.n243 585
R304 B.n500 B.n499 585
R305 B.n499 B.n498 585
R306 B.n245 B.n244 585
R307 B.n246 B.n245 585
R308 B.n491 B.n490 585
R309 B.n492 B.n491 585
R310 B.n489 B.n252 585
R311 B.n252 B.n251 585
R312 B.n488 B.n487 585
R313 B.n487 B.n486 585
R314 B.n254 B.n253 585
R315 B.n255 B.n254 585
R316 B.n479 B.n478 585
R317 B.n480 B.n479 585
R318 B.n477 B.n260 585
R319 B.n260 B.n259 585
R320 B.n476 B.n475 585
R321 B.n475 B.n474 585
R322 B.n262 B.n261 585
R323 B.n263 B.n262 585
R324 B.n467 B.n466 585
R325 B.n468 B.n467 585
R326 B.n465 B.n268 585
R327 B.n268 B.n267 585
R328 B.n464 B.n463 585
R329 B.n463 B.n462 585
R330 B.n270 B.n269 585
R331 B.n271 B.n270 585
R332 B.n455 B.n454 585
R333 B.n456 B.n455 585
R334 B.n453 B.n275 585
R335 B.n279 B.n275 585
R336 B.n452 B.n451 585
R337 B.n451 B.n450 585
R338 B.n277 B.n276 585
R339 B.n278 B.n277 585
R340 B.n443 B.n442 585
R341 B.n444 B.n443 585
R342 B.n441 B.n284 585
R343 B.n284 B.n283 585
R344 B.n440 B.n439 585
R345 B.n439 B.n438 585
R346 B.n286 B.n285 585
R347 B.n287 B.n286 585
R348 B.n434 B.n433 585
R349 B.n290 B.n289 585
R350 B.n430 B.n429 585
R351 B.n431 B.n430 585
R352 B.n428 B.n318 585
R353 B.n427 B.n426 585
R354 B.n425 B.n424 585
R355 B.n423 B.n422 585
R356 B.n421 B.n420 585
R357 B.n419 B.n418 585
R358 B.n417 B.n416 585
R359 B.n415 B.n414 585
R360 B.n413 B.n412 585
R361 B.n411 B.n410 585
R362 B.n409 B.n408 585
R363 B.n407 B.n406 585
R364 B.n405 B.n404 585
R365 B.n403 B.n402 585
R366 B.n401 B.n400 585
R367 B.n399 B.n398 585
R368 B.n397 B.n396 585
R369 B.n395 B.n394 585
R370 B.n393 B.n392 585
R371 B.n391 B.n390 585
R372 B.n389 B.n388 585
R373 B.n387 B.n386 585
R374 B.n385 B.n384 585
R375 B.n383 B.n382 585
R376 B.n381 B.n380 585
R377 B.n379 B.n378 585
R378 B.n377 B.n376 585
R379 B.n375 B.n374 585
R380 B.n373 B.n372 585
R381 B.n371 B.n370 585
R382 B.n369 B.n368 585
R383 B.n367 B.n366 585
R384 B.n365 B.n364 585
R385 B.n363 B.n362 585
R386 B.n361 B.n360 585
R387 B.n359 B.n358 585
R388 B.n357 B.n356 585
R389 B.n355 B.n354 585
R390 B.n353 B.n352 585
R391 B.n351 B.n350 585
R392 B.n349 B.n348 585
R393 B.n347 B.n346 585
R394 B.n345 B.n344 585
R395 B.n343 B.n342 585
R396 B.n341 B.n340 585
R397 B.n339 B.n338 585
R398 B.n337 B.n336 585
R399 B.n335 B.n334 585
R400 B.n333 B.n332 585
R401 B.n331 B.n330 585
R402 B.n329 B.n328 585
R403 B.n327 B.n326 585
R404 B.n325 B.n317 585
R405 B.n431 B.n317 585
R406 B.n435 B.n288 585
R407 B.n288 B.n287 585
R408 B.n437 B.n436 585
R409 B.n438 B.n437 585
R410 B.n282 B.n281 585
R411 B.n283 B.n282 585
R412 B.n446 B.n445 585
R413 B.n445 B.n444 585
R414 B.n447 B.n280 585
R415 B.n280 B.n278 585
R416 B.n449 B.n448 585
R417 B.n450 B.n449 585
R418 B.n274 B.n273 585
R419 B.n279 B.n274 585
R420 B.n458 B.n457 585
R421 B.n457 B.n456 585
R422 B.n459 B.n272 585
R423 B.n272 B.n271 585
R424 B.n461 B.n460 585
R425 B.n462 B.n461 585
R426 B.n266 B.n265 585
R427 B.n267 B.n266 585
R428 B.n470 B.n469 585
R429 B.n469 B.n468 585
R430 B.n471 B.n264 585
R431 B.n264 B.n263 585
R432 B.n473 B.n472 585
R433 B.n474 B.n473 585
R434 B.n258 B.n257 585
R435 B.n259 B.n258 585
R436 B.n482 B.n481 585
R437 B.n481 B.n480 585
R438 B.n483 B.n256 585
R439 B.n256 B.n255 585
R440 B.n485 B.n484 585
R441 B.n486 B.n485 585
R442 B.n250 B.n249 585
R443 B.n251 B.n250 585
R444 B.n494 B.n493 585
R445 B.n493 B.n492 585
R446 B.n495 B.n248 585
R447 B.n248 B.n246 585
R448 B.n497 B.n496 585
R449 B.n498 B.n497 585
R450 B.n242 B.n241 585
R451 B.n247 B.n242 585
R452 B.n506 B.n505 585
R453 B.n505 B.n504 585
R454 B.n507 B.n240 585
R455 B.n240 B.n239 585
R456 B.n509 B.n508 585
R457 B.n510 B.n509 585
R458 B.n234 B.n233 585
R459 B.n235 B.n234 585
R460 B.n519 B.n518 585
R461 B.n518 B.n517 585
R462 B.n520 B.n232 585
R463 B.n516 B.n232 585
R464 B.n522 B.n521 585
R465 B.n523 B.n522 585
R466 B.n227 B.n226 585
R467 B.n228 B.n227 585
R468 B.n531 B.n530 585
R469 B.n530 B.n529 585
R470 B.n532 B.n225 585
R471 B.n225 B.n223 585
R472 B.n534 B.n533 585
R473 B.n535 B.n534 585
R474 B.n219 B.n218 585
R475 B.n224 B.n219 585
R476 B.n544 B.n543 585
R477 B.n543 B.n542 585
R478 B.n545 B.n217 585
R479 B.n217 B.n216 585
R480 B.n547 B.n546 585
R481 B.n548 B.n547 585
R482 B.n2 B.n0 585
R483 B.n4 B.n2 585
R484 B.n3 B.n1 585
R485 B.n684 B.n3 585
R486 B.n682 B.n681 585
R487 B.n683 B.n682 585
R488 B.n680 B.n9 585
R489 B.n9 B.n8 585
R490 B.n679 B.n678 585
R491 B.n678 B.n677 585
R492 B.n11 B.n10 585
R493 B.n676 B.n11 585
R494 B.n674 B.n673 585
R495 B.n675 B.n674 585
R496 B.n672 B.n16 585
R497 B.n16 B.n15 585
R498 B.n671 B.n670 585
R499 B.n670 B.n669 585
R500 B.n18 B.n17 585
R501 B.n668 B.n18 585
R502 B.n666 B.n665 585
R503 B.n667 B.n666 585
R504 B.n664 B.n22 585
R505 B.n25 B.n22 585
R506 B.n663 B.n662 585
R507 B.n662 B.n661 585
R508 B.n24 B.n23 585
R509 B.n660 B.n24 585
R510 B.n658 B.n657 585
R511 B.n659 B.n658 585
R512 B.n656 B.n30 585
R513 B.n30 B.n29 585
R514 B.n655 B.n654 585
R515 B.n654 B.n653 585
R516 B.n32 B.n31 585
R517 B.n652 B.n32 585
R518 B.n650 B.n649 585
R519 B.n651 B.n650 585
R520 B.n648 B.n37 585
R521 B.n37 B.n36 585
R522 B.n647 B.n646 585
R523 B.n646 B.n645 585
R524 B.n39 B.n38 585
R525 B.n644 B.n39 585
R526 B.n642 B.n641 585
R527 B.n643 B.n642 585
R528 B.n640 B.n44 585
R529 B.n44 B.n43 585
R530 B.n639 B.n638 585
R531 B.n638 B.n637 585
R532 B.n46 B.n45 585
R533 B.n636 B.n46 585
R534 B.n634 B.n633 585
R535 B.n635 B.n634 585
R536 B.n632 B.n51 585
R537 B.n51 B.n50 585
R538 B.n631 B.n630 585
R539 B.n630 B.n629 585
R540 B.n53 B.n52 585
R541 B.n628 B.n53 585
R542 B.n626 B.n625 585
R543 B.n627 B.n626 585
R544 B.n624 B.n58 585
R545 B.n58 B.n57 585
R546 B.n623 B.n622 585
R547 B.n622 B.n621 585
R548 B.n60 B.n59 585
R549 B.n620 B.n60 585
R550 B.n618 B.n617 585
R551 B.n619 B.n618 585
R552 B.n616 B.n65 585
R553 B.n65 B.n64 585
R554 B.n615 B.n614 585
R555 B.n614 B.n613 585
R556 B.n67 B.n66 585
R557 B.n612 B.n67 585
R558 B.n610 B.n609 585
R559 B.n611 B.n610 585
R560 B.n608 B.n72 585
R561 B.n72 B.n71 585
R562 B.n687 B.n686 585
R563 B.n686 B.n685 585
R564 B.n433 B.n288 463.671
R565 B.n606 B.n72 463.671
R566 B.n317 B.n286 463.671
R567 B.n602 B.n102 463.671
R568 B.n322 B.t15 284.618
R569 B.n319 B.t19 284.618
R570 B.n105 B.t8 284.618
R571 B.n103 B.t12 284.618
R572 B.n604 B.n603 256.663
R573 B.n604 B.n100 256.663
R574 B.n604 B.n99 256.663
R575 B.n604 B.n98 256.663
R576 B.n604 B.n97 256.663
R577 B.n604 B.n96 256.663
R578 B.n604 B.n95 256.663
R579 B.n604 B.n94 256.663
R580 B.n604 B.n93 256.663
R581 B.n604 B.n92 256.663
R582 B.n604 B.n91 256.663
R583 B.n604 B.n90 256.663
R584 B.n604 B.n89 256.663
R585 B.n604 B.n88 256.663
R586 B.n604 B.n87 256.663
R587 B.n604 B.n86 256.663
R588 B.n604 B.n85 256.663
R589 B.n604 B.n84 256.663
R590 B.n604 B.n83 256.663
R591 B.n604 B.n82 256.663
R592 B.n604 B.n81 256.663
R593 B.n604 B.n80 256.663
R594 B.n604 B.n79 256.663
R595 B.n604 B.n78 256.663
R596 B.n604 B.n77 256.663
R597 B.n604 B.n76 256.663
R598 B.n604 B.n75 256.663
R599 B.n605 B.n604 256.663
R600 B.n432 B.n431 256.663
R601 B.n431 B.n291 256.663
R602 B.n431 B.n292 256.663
R603 B.n431 B.n293 256.663
R604 B.n431 B.n294 256.663
R605 B.n431 B.n295 256.663
R606 B.n431 B.n296 256.663
R607 B.n431 B.n297 256.663
R608 B.n431 B.n298 256.663
R609 B.n431 B.n299 256.663
R610 B.n431 B.n300 256.663
R611 B.n431 B.n301 256.663
R612 B.n431 B.n302 256.663
R613 B.n431 B.n303 256.663
R614 B.n431 B.n304 256.663
R615 B.n431 B.n305 256.663
R616 B.n431 B.n306 256.663
R617 B.n431 B.n307 256.663
R618 B.n431 B.n308 256.663
R619 B.n431 B.n309 256.663
R620 B.n431 B.n310 256.663
R621 B.n431 B.n311 256.663
R622 B.n431 B.n312 256.663
R623 B.n431 B.n313 256.663
R624 B.n431 B.n314 256.663
R625 B.n431 B.n315 256.663
R626 B.n431 B.n316 256.663
R627 B.n437 B.n288 163.367
R628 B.n437 B.n282 163.367
R629 B.n445 B.n282 163.367
R630 B.n445 B.n280 163.367
R631 B.n449 B.n280 163.367
R632 B.n449 B.n274 163.367
R633 B.n457 B.n274 163.367
R634 B.n457 B.n272 163.367
R635 B.n461 B.n272 163.367
R636 B.n461 B.n266 163.367
R637 B.n469 B.n266 163.367
R638 B.n469 B.n264 163.367
R639 B.n473 B.n264 163.367
R640 B.n473 B.n258 163.367
R641 B.n481 B.n258 163.367
R642 B.n481 B.n256 163.367
R643 B.n485 B.n256 163.367
R644 B.n485 B.n250 163.367
R645 B.n493 B.n250 163.367
R646 B.n493 B.n248 163.367
R647 B.n497 B.n248 163.367
R648 B.n497 B.n242 163.367
R649 B.n505 B.n242 163.367
R650 B.n505 B.n240 163.367
R651 B.n509 B.n240 163.367
R652 B.n509 B.n234 163.367
R653 B.n518 B.n234 163.367
R654 B.n518 B.n232 163.367
R655 B.n522 B.n232 163.367
R656 B.n522 B.n227 163.367
R657 B.n530 B.n227 163.367
R658 B.n530 B.n225 163.367
R659 B.n534 B.n225 163.367
R660 B.n534 B.n219 163.367
R661 B.n543 B.n219 163.367
R662 B.n543 B.n217 163.367
R663 B.n547 B.n217 163.367
R664 B.n547 B.n2 163.367
R665 B.n686 B.n2 163.367
R666 B.n686 B.n3 163.367
R667 B.n682 B.n3 163.367
R668 B.n682 B.n9 163.367
R669 B.n678 B.n9 163.367
R670 B.n678 B.n11 163.367
R671 B.n674 B.n11 163.367
R672 B.n674 B.n16 163.367
R673 B.n670 B.n16 163.367
R674 B.n670 B.n18 163.367
R675 B.n666 B.n18 163.367
R676 B.n666 B.n22 163.367
R677 B.n662 B.n22 163.367
R678 B.n662 B.n24 163.367
R679 B.n658 B.n24 163.367
R680 B.n658 B.n30 163.367
R681 B.n654 B.n30 163.367
R682 B.n654 B.n32 163.367
R683 B.n650 B.n32 163.367
R684 B.n650 B.n37 163.367
R685 B.n646 B.n37 163.367
R686 B.n646 B.n39 163.367
R687 B.n642 B.n39 163.367
R688 B.n642 B.n44 163.367
R689 B.n638 B.n44 163.367
R690 B.n638 B.n46 163.367
R691 B.n634 B.n46 163.367
R692 B.n634 B.n51 163.367
R693 B.n630 B.n51 163.367
R694 B.n630 B.n53 163.367
R695 B.n626 B.n53 163.367
R696 B.n626 B.n58 163.367
R697 B.n622 B.n58 163.367
R698 B.n622 B.n60 163.367
R699 B.n618 B.n60 163.367
R700 B.n618 B.n65 163.367
R701 B.n614 B.n65 163.367
R702 B.n614 B.n67 163.367
R703 B.n610 B.n67 163.367
R704 B.n610 B.n72 163.367
R705 B.n430 B.n290 163.367
R706 B.n430 B.n318 163.367
R707 B.n426 B.n425 163.367
R708 B.n422 B.n421 163.367
R709 B.n418 B.n417 163.367
R710 B.n414 B.n413 163.367
R711 B.n410 B.n409 163.367
R712 B.n406 B.n405 163.367
R713 B.n402 B.n401 163.367
R714 B.n398 B.n397 163.367
R715 B.n394 B.n393 163.367
R716 B.n390 B.n389 163.367
R717 B.n386 B.n385 163.367
R718 B.n382 B.n381 163.367
R719 B.n378 B.n377 163.367
R720 B.n374 B.n373 163.367
R721 B.n370 B.n369 163.367
R722 B.n366 B.n365 163.367
R723 B.n362 B.n361 163.367
R724 B.n358 B.n357 163.367
R725 B.n354 B.n353 163.367
R726 B.n350 B.n349 163.367
R727 B.n346 B.n345 163.367
R728 B.n342 B.n341 163.367
R729 B.n338 B.n337 163.367
R730 B.n334 B.n333 163.367
R731 B.n330 B.n329 163.367
R732 B.n326 B.n317 163.367
R733 B.n439 B.n286 163.367
R734 B.n439 B.n284 163.367
R735 B.n443 B.n284 163.367
R736 B.n443 B.n277 163.367
R737 B.n451 B.n277 163.367
R738 B.n451 B.n275 163.367
R739 B.n455 B.n275 163.367
R740 B.n455 B.n270 163.367
R741 B.n463 B.n270 163.367
R742 B.n463 B.n268 163.367
R743 B.n467 B.n268 163.367
R744 B.n467 B.n262 163.367
R745 B.n475 B.n262 163.367
R746 B.n475 B.n260 163.367
R747 B.n479 B.n260 163.367
R748 B.n479 B.n254 163.367
R749 B.n487 B.n254 163.367
R750 B.n487 B.n252 163.367
R751 B.n491 B.n252 163.367
R752 B.n491 B.n245 163.367
R753 B.n499 B.n245 163.367
R754 B.n499 B.n243 163.367
R755 B.n503 B.n243 163.367
R756 B.n503 B.n238 163.367
R757 B.n511 B.n238 163.367
R758 B.n511 B.n236 163.367
R759 B.n515 B.n236 163.367
R760 B.n515 B.n231 163.367
R761 B.n524 B.n231 163.367
R762 B.n524 B.n229 163.367
R763 B.n528 B.n229 163.367
R764 B.n528 B.n222 163.367
R765 B.n536 B.n222 163.367
R766 B.n536 B.n220 163.367
R767 B.n541 B.n220 163.367
R768 B.n541 B.n215 163.367
R769 B.n549 B.n215 163.367
R770 B.n550 B.n549 163.367
R771 B.n550 B.n5 163.367
R772 B.n6 B.n5 163.367
R773 B.n7 B.n6 163.367
R774 B.n555 B.n7 163.367
R775 B.n555 B.n12 163.367
R776 B.n13 B.n12 163.367
R777 B.n14 B.n13 163.367
R778 B.n560 B.n14 163.367
R779 B.n560 B.n19 163.367
R780 B.n20 B.n19 163.367
R781 B.n21 B.n20 163.367
R782 B.n565 B.n21 163.367
R783 B.n565 B.n26 163.367
R784 B.n27 B.n26 163.367
R785 B.n28 B.n27 163.367
R786 B.n570 B.n28 163.367
R787 B.n570 B.n33 163.367
R788 B.n34 B.n33 163.367
R789 B.n35 B.n34 163.367
R790 B.n575 B.n35 163.367
R791 B.n575 B.n40 163.367
R792 B.n41 B.n40 163.367
R793 B.n42 B.n41 163.367
R794 B.n580 B.n42 163.367
R795 B.n580 B.n47 163.367
R796 B.n48 B.n47 163.367
R797 B.n49 B.n48 163.367
R798 B.n585 B.n49 163.367
R799 B.n585 B.n54 163.367
R800 B.n55 B.n54 163.367
R801 B.n56 B.n55 163.367
R802 B.n590 B.n56 163.367
R803 B.n590 B.n61 163.367
R804 B.n62 B.n61 163.367
R805 B.n63 B.n62 163.367
R806 B.n595 B.n63 163.367
R807 B.n595 B.n68 163.367
R808 B.n69 B.n68 163.367
R809 B.n70 B.n69 163.367
R810 B.n102 B.n70 163.367
R811 B.n107 B.n74 163.367
R812 B.n111 B.n110 163.367
R813 B.n115 B.n114 163.367
R814 B.n119 B.n118 163.367
R815 B.n123 B.n122 163.367
R816 B.n127 B.n126 163.367
R817 B.n131 B.n130 163.367
R818 B.n135 B.n134 163.367
R819 B.n139 B.n138 163.367
R820 B.n143 B.n142 163.367
R821 B.n147 B.n146 163.367
R822 B.n152 B.n151 163.367
R823 B.n156 B.n155 163.367
R824 B.n160 B.n159 163.367
R825 B.n164 B.n163 163.367
R826 B.n168 B.n167 163.367
R827 B.n173 B.n172 163.367
R828 B.n177 B.n176 163.367
R829 B.n181 B.n180 163.367
R830 B.n185 B.n184 163.367
R831 B.n189 B.n188 163.367
R832 B.n193 B.n192 163.367
R833 B.n197 B.n196 163.367
R834 B.n201 B.n200 163.367
R835 B.n205 B.n204 163.367
R836 B.n209 B.n208 163.367
R837 B.n211 B.n101 163.367
R838 B.n322 B.t18 115.59
R839 B.n103 B.t13 115.59
R840 B.n319 B.t21 115.584
R841 B.n105 B.t10 115.584
R842 B.n431 B.n287 113.052
R843 B.n604 B.n71 113.052
R844 B.n323 B.t17 75.0562
R845 B.n104 B.t14 75.0562
R846 B.n320 B.t20 75.0504
R847 B.n106 B.t11 75.0504
R848 B.n433 B.n432 71.676
R849 B.n318 B.n291 71.676
R850 B.n425 B.n292 71.676
R851 B.n421 B.n293 71.676
R852 B.n417 B.n294 71.676
R853 B.n413 B.n295 71.676
R854 B.n409 B.n296 71.676
R855 B.n405 B.n297 71.676
R856 B.n401 B.n298 71.676
R857 B.n397 B.n299 71.676
R858 B.n393 B.n300 71.676
R859 B.n389 B.n301 71.676
R860 B.n385 B.n302 71.676
R861 B.n381 B.n303 71.676
R862 B.n377 B.n304 71.676
R863 B.n373 B.n305 71.676
R864 B.n369 B.n306 71.676
R865 B.n365 B.n307 71.676
R866 B.n361 B.n308 71.676
R867 B.n357 B.n309 71.676
R868 B.n353 B.n310 71.676
R869 B.n349 B.n311 71.676
R870 B.n345 B.n312 71.676
R871 B.n341 B.n313 71.676
R872 B.n337 B.n314 71.676
R873 B.n333 B.n315 71.676
R874 B.n329 B.n316 71.676
R875 B.n606 B.n605 71.676
R876 B.n107 B.n75 71.676
R877 B.n111 B.n76 71.676
R878 B.n115 B.n77 71.676
R879 B.n119 B.n78 71.676
R880 B.n123 B.n79 71.676
R881 B.n127 B.n80 71.676
R882 B.n131 B.n81 71.676
R883 B.n135 B.n82 71.676
R884 B.n139 B.n83 71.676
R885 B.n143 B.n84 71.676
R886 B.n147 B.n85 71.676
R887 B.n152 B.n86 71.676
R888 B.n156 B.n87 71.676
R889 B.n160 B.n88 71.676
R890 B.n164 B.n89 71.676
R891 B.n168 B.n90 71.676
R892 B.n173 B.n91 71.676
R893 B.n177 B.n92 71.676
R894 B.n181 B.n93 71.676
R895 B.n185 B.n94 71.676
R896 B.n189 B.n95 71.676
R897 B.n193 B.n96 71.676
R898 B.n197 B.n97 71.676
R899 B.n201 B.n98 71.676
R900 B.n205 B.n99 71.676
R901 B.n209 B.n100 71.676
R902 B.n603 B.n101 71.676
R903 B.n603 B.n602 71.676
R904 B.n211 B.n100 71.676
R905 B.n208 B.n99 71.676
R906 B.n204 B.n98 71.676
R907 B.n200 B.n97 71.676
R908 B.n196 B.n96 71.676
R909 B.n192 B.n95 71.676
R910 B.n188 B.n94 71.676
R911 B.n184 B.n93 71.676
R912 B.n180 B.n92 71.676
R913 B.n176 B.n91 71.676
R914 B.n172 B.n90 71.676
R915 B.n167 B.n89 71.676
R916 B.n163 B.n88 71.676
R917 B.n159 B.n87 71.676
R918 B.n155 B.n86 71.676
R919 B.n151 B.n85 71.676
R920 B.n146 B.n84 71.676
R921 B.n142 B.n83 71.676
R922 B.n138 B.n82 71.676
R923 B.n134 B.n81 71.676
R924 B.n130 B.n80 71.676
R925 B.n126 B.n79 71.676
R926 B.n122 B.n78 71.676
R927 B.n118 B.n77 71.676
R928 B.n114 B.n76 71.676
R929 B.n110 B.n75 71.676
R930 B.n605 B.n74 71.676
R931 B.n432 B.n290 71.676
R932 B.n426 B.n291 71.676
R933 B.n422 B.n292 71.676
R934 B.n418 B.n293 71.676
R935 B.n414 B.n294 71.676
R936 B.n410 B.n295 71.676
R937 B.n406 B.n296 71.676
R938 B.n402 B.n297 71.676
R939 B.n398 B.n298 71.676
R940 B.n394 B.n299 71.676
R941 B.n390 B.n300 71.676
R942 B.n386 B.n301 71.676
R943 B.n382 B.n302 71.676
R944 B.n378 B.n303 71.676
R945 B.n374 B.n304 71.676
R946 B.n370 B.n305 71.676
R947 B.n366 B.n306 71.676
R948 B.n362 B.n307 71.676
R949 B.n358 B.n308 71.676
R950 B.n354 B.n309 71.676
R951 B.n350 B.n310 71.676
R952 B.n346 B.n311 71.676
R953 B.n342 B.n312 71.676
R954 B.n338 B.n313 71.676
R955 B.n334 B.n314 71.676
R956 B.n330 B.n315 71.676
R957 B.n326 B.n316 71.676
R958 B.n438 B.n287 68.0314
R959 B.n438 B.n283 68.0314
R960 B.n444 B.n283 68.0314
R961 B.n444 B.n278 68.0314
R962 B.n450 B.n278 68.0314
R963 B.n450 B.n279 68.0314
R964 B.n456 B.n271 68.0314
R965 B.n462 B.n271 68.0314
R966 B.n462 B.n267 68.0314
R967 B.n468 B.n267 68.0314
R968 B.n468 B.n263 68.0314
R969 B.n474 B.n263 68.0314
R970 B.n474 B.n259 68.0314
R971 B.n480 B.n259 68.0314
R972 B.n486 B.n255 68.0314
R973 B.n486 B.n251 68.0314
R974 B.n492 B.n251 68.0314
R975 B.n492 B.n246 68.0314
R976 B.n498 B.n246 68.0314
R977 B.n498 B.n247 68.0314
R978 B.n504 B.n239 68.0314
R979 B.n510 B.n239 68.0314
R980 B.n510 B.n235 68.0314
R981 B.n517 B.n235 68.0314
R982 B.n517 B.n516 68.0314
R983 B.n523 B.n228 68.0314
R984 B.n529 B.n228 68.0314
R985 B.n529 B.n223 68.0314
R986 B.n535 B.n223 68.0314
R987 B.n535 B.n224 68.0314
R988 B.n542 B.n216 68.0314
R989 B.n548 B.n216 68.0314
R990 B.n548 B.n4 68.0314
R991 B.n685 B.n4 68.0314
R992 B.n685 B.n684 68.0314
R993 B.n684 B.n683 68.0314
R994 B.n683 B.n8 68.0314
R995 B.n677 B.n8 68.0314
R996 B.n676 B.n675 68.0314
R997 B.n675 B.n15 68.0314
R998 B.n669 B.n15 68.0314
R999 B.n669 B.n668 68.0314
R1000 B.n668 B.n667 68.0314
R1001 B.n661 B.n25 68.0314
R1002 B.n661 B.n660 68.0314
R1003 B.n660 B.n659 68.0314
R1004 B.n659 B.n29 68.0314
R1005 B.n653 B.n29 68.0314
R1006 B.n652 B.n651 68.0314
R1007 B.n651 B.n36 68.0314
R1008 B.n645 B.n36 68.0314
R1009 B.n645 B.n644 68.0314
R1010 B.n644 B.n643 68.0314
R1011 B.n643 B.n43 68.0314
R1012 B.n637 B.n636 68.0314
R1013 B.n636 B.n635 68.0314
R1014 B.n635 B.n50 68.0314
R1015 B.n629 B.n50 68.0314
R1016 B.n629 B.n628 68.0314
R1017 B.n628 B.n627 68.0314
R1018 B.n627 B.n57 68.0314
R1019 B.n621 B.n57 68.0314
R1020 B.n620 B.n619 68.0314
R1021 B.n619 B.n64 68.0314
R1022 B.n613 B.n64 68.0314
R1023 B.n613 B.n612 68.0314
R1024 B.n612 B.n611 68.0314
R1025 B.n611 B.n71 68.0314
R1026 B.n504 B.t2 66.0305
R1027 B.n653 B.t1 66.0305
R1028 B.n480 B.t6 60.0278
R1029 B.n637 B.t4 60.0278
R1030 B.n324 B.n323 59.5399
R1031 B.n321 B.n320 59.5399
R1032 B.n149 B.n106 59.5399
R1033 B.n170 B.n104 59.5399
R1034 B.n523 B.t3 56.026
R1035 B.n667 B.t0 56.026
R1036 B.n542 B.t7 46.0214
R1037 B.n677 B.t5 46.0214
R1038 B.n323 B.n322 40.5338
R1039 B.n320 B.n319 40.5338
R1040 B.n106 B.n105 40.5338
R1041 B.n104 B.n103 40.5338
R1042 B.n279 B.t16 36.0169
R1043 B.t9 B.n620 36.0169
R1044 B.n456 B.t16 32.0151
R1045 B.n621 B.t9 32.0151
R1046 B.n608 B.n607 30.1273
R1047 B.n601 B.n600 30.1273
R1048 B.n325 B.n285 30.1273
R1049 B.n435 B.n434 30.1273
R1050 B.n224 B.t7 22.0105
R1051 B.t5 B.n676 22.0105
R1052 B B.n687 18.0485
R1053 B.n516 B.t3 12.006
R1054 B.n25 B.t0 12.006
R1055 B.n607 B.n73 10.6151
R1056 B.n108 B.n73 10.6151
R1057 B.n109 B.n108 10.6151
R1058 B.n112 B.n109 10.6151
R1059 B.n113 B.n112 10.6151
R1060 B.n116 B.n113 10.6151
R1061 B.n117 B.n116 10.6151
R1062 B.n120 B.n117 10.6151
R1063 B.n121 B.n120 10.6151
R1064 B.n124 B.n121 10.6151
R1065 B.n125 B.n124 10.6151
R1066 B.n128 B.n125 10.6151
R1067 B.n129 B.n128 10.6151
R1068 B.n132 B.n129 10.6151
R1069 B.n133 B.n132 10.6151
R1070 B.n136 B.n133 10.6151
R1071 B.n137 B.n136 10.6151
R1072 B.n140 B.n137 10.6151
R1073 B.n141 B.n140 10.6151
R1074 B.n144 B.n141 10.6151
R1075 B.n145 B.n144 10.6151
R1076 B.n148 B.n145 10.6151
R1077 B.n153 B.n150 10.6151
R1078 B.n154 B.n153 10.6151
R1079 B.n157 B.n154 10.6151
R1080 B.n158 B.n157 10.6151
R1081 B.n161 B.n158 10.6151
R1082 B.n162 B.n161 10.6151
R1083 B.n165 B.n162 10.6151
R1084 B.n166 B.n165 10.6151
R1085 B.n169 B.n166 10.6151
R1086 B.n174 B.n171 10.6151
R1087 B.n175 B.n174 10.6151
R1088 B.n178 B.n175 10.6151
R1089 B.n179 B.n178 10.6151
R1090 B.n182 B.n179 10.6151
R1091 B.n183 B.n182 10.6151
R1092 B.n186 B.n183 10.6151
R1093 B.n187 B.n186 10.6151
R1094 B.n190 B.n187 10.6151
R1095 B.n191 B.n190 10.6151
R1096 B.n194 B.n191 10.6151
R1097 B.n195 B.n194 10.6151
R1098 B.n198 B.n195 10.6151
R1099 B.n199 B.n198 10.6151
R1100 B.n202 B.n199 10.6151
R1101 B.n203 B.n202 10.6151
R1102 B.n206 B.n203 10.6151
R1103 B.n207 B.n206 10.6151
R1104 B.n210 B.n207 10.6151
R1105 B.n212 B.n210 10.6151
R1106 B.n213 B.n212 10.6151
R1107 B.n601 B.n213 10.6151
R1108 B.n440 B.n285 10.6151
R1109 B.n441 B.n440 10.6151
R1110 B.n442 B.n441 10.6151
R1111 B.n442 B.n276 10.6151
R1112 B.n452 B.n276 10.6151
R1113 B.n453 B.n452 10.6151
R1114 B.n454 B.n453 10.6151
R1115 B.n454 B.n269 10.6151
R1116 B.n464 B.n269 10.6151
R1117 B.n465 B.n464 10.6151
R1118 B.n466 B.n465 10.6151
R1119 B.n466 B.n261 10.6151
R1120 B.n476 B.n261 10.6151
R1121 B.n477 B.n476 10.6151
R1122 B.n478 B.n477 10.6151
R1123 B.n478 B.n253 10.6151
R1124 B.n488 B.n253 10.6151
R1125 B.n489 B.n488 10.6151
R1126 B.n490 B.n489 10.6151
R1127 B.n490 B.n244 10.6151
R1128 B.n500 B.n244 10.6151
R1129 B.n501 B.n500 10.6151
R1130 B.n502 B.n501 10.6151
R1131 B.n502 B.n237 10.6151
R1132 B.n512 B.n237 10.6151
R1133 B.n513 B.n512 10.6151
R1134 B.n514 B.n513 10.6151
R1135 B.n514 B.n230 10.6151
R1136 B.n525 B.n230 10.6151
R1137 B.n526 B.n525 10.6151
R1138 B.n527 B.n526 10.6151
R1139 B.n527 B.n221 10.6151
R1140 B.n537 B.n221 10.6151
R1141 B.n538 B.n537 10.6151
R1142 B.n540 B.n538 10.6151
R1143 B.n540 B.n539 10.6151
R1144 B.n539 B.n214 10.6151
R1145 B.n551 B.n214 10.6151
R1146 B.n552 B.n551 10.6151
R1147 B.n553 B.n552 10.6151
R1148 B.n554 B.n553 10.6151
R1149 B.n556 B.n554 10.6151
R1150 B.n557 B.n556 10.6151
R1151 B.n558 B.n557 10.6151
R1152 B.n559 B.n558 10.6151
R1153 B.n561 B.n559 10.6151
R1154 B.n562 B.n561 10.6151
R1155 B.n563 B.n562 10.6151
R1156 B.n564 B.n563 10.6151
R1157 B.n566 B.n564 10.6151
R1158 B.n567 B.n566 10.6151
R1159 B.n568 B.n567 10.6151
R1160 B.n569 B.n568 10.6151
R1161 B.n571 B.n569 10.6151
R1162 B.n572 B.n571 10.6151
R1163 B.n573 B.n572 10.6151
R1164 B.n574 B.n573 10.6151
R1165 B.n576 B.n574 10.6151
R1166 B.n577 B.n576 10.6151
R1167 B.n578 B.n577 10.6151
R1168 B.n579 B.n578 10.6151
R1169 B.n581 B.n579 10.6151
R1170 B.n582 B.n581 10.6151
R1171 B.n583 B.n582 10.6151
R1172 B.n584 B.n583 10.6151
R1173 B.n586 B.n584 10.6151
R1174 B.n587 B.n586 10.6151
R1175 B.n588 B.n587 10.6151
R1176 B.n589 B.n588 10.6151
R1177 B.n591 B.n589 10.6151
R1178 B.n592 B.n591 10.6151
R1179 B.n593 B.n592 10.6151
R1180 B.n594 B.n593 10.6151
R1181 B.n596 B.n594 10.6151
R1182 B.n597 B.n596 10.6151
R1183 B.n598 B.n597 10.6151
R1184 B.n599 B.n598 10.6151
R1185 B.n600 B.n599 10.6151
R1186 B.n434 B.n289 10.6151
R1187 B.n429 B.n289 10.6151
R1188 B.n429 B.n428 10.6151
R1189 B.n428 B.n427 10.6151
R1190 B.n427 B.n424 10.6151
R1191 B.n424 B.n423 10.6151
R1192 B.n423 B.n420 10.6151
R1193 B.n420 B.n419 10.6151
R1194 B.n419 B.n416 10.6151
R1195 B.n416 B.n415 10.6151
R1196 B.n415 B.n412 10.6151
R1197 B.n412 B.n411 10.6151
R1198 B.n411 B.n408 10.6151
R1199 B.n408 B.n407 10.6151
R1200 B.n407 B.n404 10.6151
R1201 B.n404 B.n403 10.6151
R1202 B.n403 B.n400 10.6151
R1203 B.n400 B.n399 10.6151
R1204 B.n399 B.n396 10.6151
R1205 B.n396 B.n395 10.6151
R1206 B.n395 B.n392 10.6151
R1207 B.n392 B.n391 10.6151
R1208 B.n388 B.n387 10.6151
R1209 B.n387 B.n384 10.6151
R1210 B.n384 B.n383 10.6151
R1211 B.n383 B.n380 10.6151
R1212 B.n380 B.n379 10.6151
R1213 B.n379 B.n376 10.6151
R1214 B.n376 B.n375 10.6151
R1215 B.n375 B.n372 10.6151
R1216 B.n372 B.n371 10.6151
R1217 B.n368 B.n367 10.6151
R1218 B.n367 B.n364 10.6151
R1219 B.n364 B.n363 10.6151
R1220 B.n363 B.n360 10.6151
R1221 B.n360 B.n359 10.6151
R1222 B.n359 B.n356 10.6151
R1223 B.n356 B.n355 10.6151
R1224 B.n355 B.n352 10.6151
R1225 B.n352 B.n351 10.6151
R1226 B.n351 B.n348 10.6151
R1227 B.n348 B.n347 10.6151
R1228 B.n347 B.n344 10.6151
R1229 B.n344 B.n343 10.6151
R1230 B.n343 B.n340 10.6151
R1231 B.n340 B.n339 10.6151
R1232 B.n339 B.n336 10.6151
R1233 B.n336 B.n335 10.6151
R1234 B.n335 B.n332 10.6151
R1235 B.n332 B.n331 10.6151
R1236 B.n331 B.n328 10.6151
R1237 B.n328 B.n327 10.6151
R1238 B.n327 B.n325 10.6151
R1239 B.n436 B.n435 10.6151
R1240 B.n436 B.n281 10.6151
R1241 B.n446 B.n281 10.6151
R1242 B.n447 B.n446 10.6151
R1243 B.n448 B.n447 10.6151
R1244 B.n448 B.n273 10.6151
R1245 B.n458 B.n273 10.6151
R1246 B.n459 B.n458 10.6151
R1247 B.n460 B.n459 10.6151
R1248 B.n460 B.n265 10.6151
R1249 B.n470 B.n265 10.6151
R1250 B.n471 B.n470 10.6151
R1251 B.n472 B.n471 10.6151
R1252 B.n472 B.n257 10.6151
R1253 B.n482 B.n257 10.6151
R1254 B.n483 B.n482 10.6151
R1255 B.n484 B.n483 10.6151
R1256 B.n484 B.n249 10.6151
R1257 B.n494 B.n249 10.6151
R1258 B.n495 B.n494 10.6151
R1259 B.n496 B.n495 10.6151
R1260 B.n496 B.n241 10.6151
R1261 B.n506 B.n241 10.6151
R1262 B.n507 B.n506 10.6151
R1263 B.n508 B.n507 10.6151
R1264 B.n508 B.n233 10.6151
R1265 B.n519 B.n233 10.6151
R1266 B.n520 B.n519 10.6151
R1267 B.n521 B.n520 10.6151
R1268 B.n521 B.n226 10.6151
R1269 B.n531 B.n226 10.6151
R1270 B.n532 B.n531 10.6151
R1271 B.n533 B.n532 10.6151
R1272 B.n533 B.n218 10.6151
R1273 B.n544 B.n218 10.6151
R1274 B.n545 B.n544 10.6151
R1275 B.n546 B.n545 10.6151
R1276 B.n546 B.n0 10.6151
R1277 B.n681 B.n1 10.6151
R1278 B.n681 B.n680 10.6151
R1279 B.n680 B.n679 10.6151
R1280 B.n679 B.n10 10.6151
R1281 B.n673 B.n10 10.6151
R1282 B.n673 B.n672 10.6151
R1283 B.n672 B.n671 10.6151
R1284 B.n671 B.n17 10.6151
R1285 B.n665 B.n17 10.6151
R1286 B.n665 B.n664 10.6151
R1287 B.n664 B.n663 10.6151
R1288 B.n663 B.n23 10.6151
R1289 B.n657 B.n23 10.6151
R1290 B.n657 B.n656 10.6151
R1291 B.n656 B.n655 10.6151
R1292 B.n655 B.n31 10.6151
R1293 B.n649 B.n31 10.6151
R1294 B.n649 B.n648 10.6151
R1295 B.n648 B.n647 10.6151
R1296 B.n647 B.n38 10.6151
R1297 B.n641 B.n38 10.6151
R1298 B.n641 B.n640 10.6151
R1299 B.n640 B.n639 10.6151
R1300 B.n639 B.n45 10.6151
R1301 B.n633 B.n45 10.6151
R1302 B.n633 B.n632 10.6151
R1303 B.n632 B.n631 10.6151
R1304 B.n631 B.n52 10.6151
R1305 B.n625 B.n52 10.6151
R1306 B.n625 B.n624 10.6151
R1307 B.n624 B.n623 10.6151
R1308 B.n623 B.n59 10.6151
R1309 B.n617 B.n59 10.6151
R1310 B.n617 B.n616 10.6151
R1311 B.n616 B.n615 10.6151
R1312 B.n615 B.n66 10.6151
R1313 B.n609 B.n66 10.6151
R1314 B.n609 B.n608 10.6151
R1315 B.n149 B.n148 9.36635
R1316 B.n171 B.n170 9.36635
R1317 B.n391 B.n321 9.36635
R1318 B.n368 B.n324 9.36635
R1319 B.t6 B.n255 8.00414
R1320 B.t4 B.n43 8.00414
R1321 B.n687 B.n0 2.81026
R1322 B.n687 B.n1 2.81026
R1323 B.n247 B.t2 2.00141
R1324 B.t1 B.n652 2.00141
R1325 B.n150 B.n149 1.24928
R1326 B.n170 B.n169 1.24928
R1327 B.n388 B.n321 1.24928
R1328 B.n371 B.n324 1.24928
R1329 VN.n22 VN.n21 179.252
R1330 VN.n45 VN.n44 179.252
R1331 VN.n43 VN.n23 161.3
R1332 VN.n42 VN.n41 161.3
R1333 VN.n40 VN.n24 161.3
R1334 VN.n39 VN.n38 161.3
R1335 VN.n36 VN.n25 161.3
R1336 VN.n35 VN.n34 161.3
R1337 VN.n33 VN.n26 161.3
R1338 VN.n32 VN.n31 161.3
R1339 VN.n30 VN.n27 161.3
R1340 VN.n20 VN.n0 161.3
R1341 VN.n19 VN.n18 161.3
R1342 VN.n17 VN.n1 161.3
R1343 VN.n16 VN.n15 161.3
R1344 VN.n13 VN.n2 161.3
R1345 VN.n12 VN.n11 161.3
R1346 VN.n10 VN.n3 161.3
R1347 VN.n9 VN.n8 161.3
R1348 VN.n7 VN.n4 161.3
R1349 VN.n5 VN.t1 109.865
R1350 VN.n28 VN.t7 109.865
R1351 VN.n6 VN.t3 78.3255
R1352 VN.n14 VN.t2 78.3255
R1353 VN.n21 VN.t0 78.3255
R1354 VN.n29 VN.t6 78.3255
R1355 VN.n37 VN.t4 78.3255
R1356 VN.n44 VN.t5 78.3255
R1357 VN.n6 VN.n5 65.8068
R1358 VN.n29 VN.n28 65.8068
R1359 VN.n19 VN.n1 49.296
R1360 VN.n42 VN.n24 49.296
R1361 VN VN.n45 42.5251
R1362 VN.n8 VN.n3 40.577
R1363 VN.n12 VN.n3 40.577
R1364 VN.n31 VN.n26 40.577
R1365 VN.n35 VN.n26 40.577
R1366 VN.n15 VN.n1 31.8581
R1367 VN.n38 VN.n24 31.8581
R1368 VN.n8 VN.n7 24.5923
R1369 VN.n13 VN.n12 24.5923
R1370 VN.n20 VN.n19 24.5923
R1371 VN.n31 VN.n30 24.5923
R1372 VN.n36 VN.n35 24.5923
R1373 VN.n43 VN.n42 24.5923
R1374 VN.n15 VN.n14 22.3791
R1375 VN.n38 VN.n37 22.3791
R1376 VN.n28 VN.n27 18.2204
R1377 VN.n5 VN.n4 18.2204
R1378 VN.n21 VN.n20 6.6403
R1379 VN.n44 VN.n43 6.6403
R1380 VN.n7 VN.n6 2.21377
R1381 VN.n14 VN.n13 2.21377
R1382 VN.n30 VN.n29 2.21377
R1383 VN.n37 VN.n36 2.21377
R1384 VN.n45 VN.n23 0.189894
R1385 VN.n41 VN.n23 0.189894
R1386 VN.n41 VN.n40 0.189894
R1387 VN.n40 VN.n39 0.189894
R1388 VN.n39 VN.n25 0.189894
R1389 VN.n34 VN.n25 0.189894
R1390 VN.n34 VN.n33 0.189894
R1391 VN.n33 VN.n32 0.189894
R1392 VN.n32 VN.n27 0.189894
R1393 VN.n9 VN.n4 0.189894
R1394 VN.n10 VN.n9 0.189894
R1395 VN.n11 VN.n10 0.189894
R1396 VN.n11 VN.n2 0.189894
R1397 VN.n16 VN.n2 0.189894
R1398 VN.n17 VN.n16 0.189894
R1399 VN.n18 VN.n17 0.189894
R1400 VN.n18 VN.n0 0.189894
R1401 VN.n22 VN.n0 0.189894
R1402 VN VN.n22 0.0516364
R1403 VDD2.n2 VDD2.n1 70.2668
R1404 VDD2.n2 VDD2.n0 70.2668
R1405 VDD2 VDD2.n5 70.264
R1406 VDD2.n4 VDD2.n3 69.4215
R1407 VDD2.n4 VDD2.n2 36.7541
R1408 VDD2.n5 VDD2.t1 3.46204
R1409 VDD2.n5 VDD2.t0 3.46204
R1410 VDD2.n3 VDD2.t2 3.46204
R1411 VDD2.n3 VDD2.t3 3.46204
R1412 VDD2.n1 VDD2.t5 3.46204
R1413 VDD2.n1 VDD2.t7 3.46204
R1414 VDD2.n0 VDD2.t6 3.46204
R1415 VDD2.n0 VDD2.t4 3.46204
R1416 VDD2 VDD2.n4 0.959552
C0 VTAIL VDD1 5.58507f
C1 VTAIL VN 4.5216f
C2 VP VDD2 0.430413f
C3 VTAIL VP 4.5357f
C4 VN VDD1 0.150337f
C5 VTAIL VDD2 5.63385f
C6 VP VDD1 4.28789f
C7 VN VP 5.46551f
C8 VDD1 VDD2 1.33895f
C9 VN VDD2 4.00879f
C10 VDD2 B 4.042892f
C11 VDD1 B 4.396973f
C12 VTAIL B 5.886528f
C13 VN B 11.64085f
C14 VP B 10.209142f
C15 VDD2.t6 B 0.110718f
C16 VDD2.t4 B 0.110718f
C17 VDD2.n0 B 0.923341f
C18 VDD2.t5 B 0.110718f
C19 VDD2.t7 B 0.110718f
C20 VDD2.n1 B 0.923341f
C21 VDD2.n2 B 2.3521f
C22 VDD2.t2 B 0.110718f
C23 VDD2.t3 B 0.110718f
C24 VDD2.n3 B 0.918327f
C25 VDD2.n4 B 2.12053f
C26 VDD2.t1 B 0.110718f
C27 VDD2.t0 B 0.110718f
C28 VDD2.n5 B 0.923312f
C29 VN.n0 B 0.030673f
C30 VN.t0 B 0.814944f
C31 VN.n1 B 0.028094f
C32 VN.n2 B 0.030673f
C33 VN.t2 B 0.814944f
C34 VN.n3 B 0.024773f
C35 VN.n4 B 0.198654f
C36 VN.t3 B 0.814944f
C37 VN.t1 B 0.944242f
C38 VN.n5 B 0.387219f
C39 VN.n6 B 0.370938f
C40 VN.n7 B 0.031327f
C41 VN.n8 B 0.060641f
C42 VN.n9 B 0.030673f
C43 VN.n10 B 0.030673f
C44 VN.n11 B 0.030673f
C45 VN.n12 B 0.060641f
C46 VN.n13 B 0.031327f
C47 VN.n14 B 0.316538f
C48 VN.n15 B 0.058836f
C49 VN.n16 B 0.030673f
C50 VN.n17 B 0.030673f
C51 VN.n18 B 0.030673f
C52 VN.n19 B 0.056598f
C53 VN.n20 B 0.036381f
C54 VN.n21 B 0.387683f
C55 VN.n22 B 0.031688f
C56 VN.n23 B 0.030673f
C57 VN.t5 B 0.814944f
C58 VN.n24 B 0.028094f
C59 VN.n25 B 0.030673f
C60 VN.t4 B 0.814944f
C61 VN.n26 B 0.024773f
C62 VN.n27 B 0.198654f
C63 VN.t6 B 0.814944f
C64 VN.t7 B 0.944242f
C65 VN.n28 B 0.387219f
C66 VN.n29 B 0.370938f
C67 VN.n30 B 0.031327f
C68 VN.n31 B 0.060641f
C69 VN.n32 B 0.030673f
C70 VN.n33 B 0.030673f
C71 VN.n34 B 0.030673f
C72 VN.n35 B 0.060641f
C73 VN.n36 B 0.031327f
C74 VN.n37 B 0.316538f
C75 VN.n38 B 0.058836f
C76 VN.n39 B 0.030673f
C77 VN.n40 B 0.030673f
C78 VN.n41 B 0.030673f
C79 VN.n42 B 0.056598f
C80 VN.n43 B 0.036381f
C81 VN.n44 B 0.387683f
C82 VN.n45 B 1.30135f
C83 VDD1.t5 B 0.113112f
C84 VDD1.t0 B 0.113112f
C85 VDD1.n0 B 0.944103f
C86 VDD1.t6 B 0.113112f
C87 VDD1.t2 B 0.113112f
C88 VDD1.n1 B 0.943306f
C89 VDD1.t3 B 0.113112f
C90 VDD1.t7 B 0.113112f
C91 VDD1.n2 B 0.943306f
C92 VDD1.n3 B 2.4558f
C93 VDD1.t1 B 0.113112f
C94 VDD1.t4 B 0.113112f
C95 VDD1.n4 B 0.938179f
C96 VDD1.n5 B 2.19659f
C97 VTAIL.t15 B 0.100871f
C98 VTAIL.t13 B 0.100871f
C99 VTAIL.n0 B 0.781089f
C100 VTAIL.n1 B 0.338909f
C101 VTAIL.t11 B 0.997354f
C102 VTAIL.n2 B 0.427346f
C103 VTAIL.t3 B 0.997354f
C104 VTAIL.n3 B 0.427346f
C105 VTAIL.t4 B 0.100871f
C106 VTAIL.t6 B 0.100871f
C107 VTAIL.n4 B 0.781089f
C108 VTAIL.n5 B 0.464281f
C109 VTAIL.t7 B 0.997354f
C110 VTAIL.n6 B 1.18083f
C111 VTAIL.t10 B 0.997358f
C112 VTAIL.n7 B 1.18083f
C113 VTAIL.t14 B 0.100871f
C114 VTAIL.t8 B 0.100871f
C115 VTAIL.n8 B 0.781093f
C116 VTAIL.n9 B 0.464277f
C117 VTAIL.t9 B 0.997358f
C118 VTAIL.n10 B 0.427342f
C119 VTAIL.t5 B 0.997358f
C120 VTAIL.n11 B 0.427342f
C121 VTAIL.t1 B 0.100871f
C122 VTAIL.t2 B 0.100871f
C123 VTAIL.n12 B 0.781093f
C124 VTAIL.n13 B 0.464277f
C125 VTAIL.t0 B 0.997354f
C126 VTAIL.n14 B 1.18083f
C127 VTAIL.t12 B 0.997354f
C128 VTAIL.n15 B 1.17665f
C129 VP.n0 B 0.031427f
C130 VP.t0 B 0.834978f
C131 VP.n1 B 0.028785f
C132 VP.n2 B 0.031427f
C133 VP.t4 B 0.834978f
C134 VP.n3 B 0.025382f
C135 VP.n4 B 0.031427f
C136 VP.t5 B 0.834978f
C137 VP.n5 B 0.028785f
C138 VP.n6 B 0.031427f
C139 VP.t1 B 0.834978f
C140 VP.n7 B 0.031427f
C141 VP.t3 B 0.834978f
C142 VP.n8 B 0.028785f
C143 VP.n9 B 0.031427f
C144 VP.t6 B 0.834978f
C145 VP.n10 B 0.025382f
C146 VP.n11 B 0.203537f
C147 VP.t7 B 0.834978f
C148 VP.t2 B 0.967456f
C149 VP.n12 B 0.396738f
C150 VP.n13 B 0.380057f
C151 VP.n14 B 0.032097f
C152 VP.n15 B 0.062132f
C153 VP.n16 B 0.031427f
C154 VP.n17 B 0.031427f
C155 VP.n18 B 0.031427f
C156 VP.n19 B 0.062132f
C157 VP.n20 B 0.032097f
C158 VP.n21 B 0.32432f
C159 VP.n22 B 0.060282f
C160 VP.n23 B 0.031427f
C161 VP.n24 B 0.031427f
C162 VP.n25 B 0.031427f
C163 VP.n26 B 0.05799f
C164 VP.n27 B 0.037276f
C165 VP.n28 B 0.397214f
C166 VP.n29 B 1.31271f
C167 VP.n30 B 1.3396f
C168 VP.n31 B 0.397214f
C169 VP.n32 B 0.037276f
C170 VP.n33 B 0.05799f
C171 VP.n34 B 0.031427f
C172 VP.n35 B 0.031427f
C173 VP.n36 B 0.031427f
C174 VP.n37 B 0.060282f
C175 VP.n38 B 0.32432f
C176 VP.n39 B 0.032097f
C177 VP.n40 B 0.062132f
C178 VP.n41 B 0.031427f
C179 VP.n42 B 0.031427f
C180 VP.n43 B 0.031427f
C181 VP.n44 B 0.062132f
C182 VP.n45 B 0.032097f
C183 VP.n46 B 0.32432f
C184 VP.n47 B 0.060282f
C185 VP.n48 B 0.031427f
C186 VP.n49 B 0.031427f
C187 VP.n50 B 0.031427f
C188 VP.n51 B 0.05799f
C189 VP.n52 B 0.037276f
C190 VP.n53 B 0.397214f
C191 VP.n54 B 0.032467f
.ends

