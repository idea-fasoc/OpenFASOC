* NGSPICE file created from diff_pair_sample_0042.ext - technology: sky130A

.subckt diff_pair_sample_0042 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=0.59
X1 VTAIL.t11 VN.t0 VDD2.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=0.59
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=0.59
X3 VDD2.t0 VN.t1 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=0.59
X4 VTAIL.t9 VN.t2 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=0.59
X5 VDD2.t1 VN.t3 VTAIL.t8 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=0.59
X6 VDD1.t5 VP.t0 VTAIL.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=0.59
X7 VDD1.t4 VP.t1 VTAIL.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=0.59
X8 VDD2.t3 VN.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=0.59
X9 VDD1.t3 VP.t2 VTAIL.t4 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=0.59
X10 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=0.59
X11 VDD1.t2 VP.t3 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=4.7385 ps=25.08 w=12.15 l=0.59
X12 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=0 ps=0 w=12.15 l=0.59
X13 VTAIL.t1 VP.t4 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=0.59
X14 VDD2.t5 VN.t5 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=4.7385 pd=25.08 as=2.00475 ps=12.48 w=12.15 l=0.59
X15 VTAIL.t0 VP.t5 VDD1.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.00475 pd=12.48 as=2.00475 ps=12.48 w=12.15 l=0.59
R0 B.n359 B.t6 700.866
R1 B.n357 B.t17 700.866
R2 B.n90 B.t10 700.866
R3 B.n87 B.t14 700.866
R4 B.n632 B.n631 585
R5 B.n273 B.n85 585
R6 B.n272 B.n271 585
R7 B.n270 B.n269 585
R8 B.n268 B.n267 585
R9 B.n266 B.n265 585
R10 B.n264 B.n263 585
R11 B.n262 B.n261 585
R12 B.n260 B.n259 585
R13 B.n258 B.n257 585
R14 B.n256 B.n255 585
R15 B.n254 B.n253 585
R16 B.n252 B.n251 585
R17 B.n250 B.n249 585
R18 B.n248 B.n247 585
R19 B.n246 B.n245 585
R20 B.n244 B.n243 585
R21 B.n242 B.n241 585
R22 B.n240 B.n239 585
R23 B.n238 B.n237 585
R24 B.n236 B.n235 585
R25 B.n234 B.n233 585
R26 B.n232 B.n231 585
R27 B.n230 B.n229 585
R28 B.n228 B.n227 585
R29 B.n226 B.n225 585
R30 B.n224 B.n223 585
R31 B.n222 B.n221 585
R32 B.n220 B.n219 585
R33 B.n218 B.n217 585
R34 B.n216 B.n215 585
R35 B.n214 B.n213 585
R36 B.n212 B.n211 585
R37 B.n210 B.n209 585
R38 B.n208 B.n207 585
R39 B.n206 B.n205 585
R40 B.n204 B.n203 585
R41 B.n202 B.n201 585
R42 B.n200 B.n199 585
R43 B.n198 B.n197 585
R44 B.n196 B.n195 585
R45 B.n194 B.n193 585
R46 B.n192 B.n191 585
R47 B.n190 B.n189 585
R48 B.n188 B.n187 585
R49 B.n186 B.n185 585
R50 B.n184 B.n183 585
R51 B.n182 B.n181 585
R52 B.n180 B.n179 585
R53 B.n178 B.n177 585
R54 B.n176 B.n175 585
R55 B.n174 B.n173 585
R56 B.n172 B.n171 585
R57 B.n170 B.n169 585
R58 B.n168 B.n167 585
R59 B.n166 B.n165 585
R60 B.n164 B.n163 585
R61 B.n162 B.n161 585
R62 B.n160 B.n159 585
R63 B.n158 B.n157 585
R64 B.n156 B.n155 585
R65 B.n154 B.n153 585
R66 B.n152 B.n151 585
R67 B.n150 B.n149 585
R68 B.n148 B.n147 585
R69 B.n146 B.n145 585
R70 B.n144 B.n143 585
R71 B.n142 B.n141 585
R72 B.n140 B.n139 585
R73 B.n138 B.n137 585
R74 B.n136 B.n135 585
R75 B.n134 B.n133 585
R76 B.n132 B.n131 585
R77 B.n130 B.n129 585
R78 B.n128 B.n127 585
R79 B.n126 B.n125 585
R80 B.n124 B.n123 585
R81 B.n122 B.n121 585
R82 B.n120 B.n119 585
R83 B.n118 B.n117 585
R84 B.n116 B.n115 585
R85 B.n114 B.n113 585
R86 B.n112 B.n111 585
R87 B.n110 B.n109 585
R88 B.n108 B.n107 585
R89 B.n106 B.n105 585
R90 B.n104 B.n103 585
R91 B.n102 B.n101 585
R92 B.n100 B.n99 585
R93 B.n98 B.n97 585
R94 B.n96 B.n95 585
R95 B.n94 B.n93 585
R96 B.n39 B.n38 585
R97 B.n637 B.n636 585
R98 B.n630 B.n86 585
R99 B.n86 B.n36 585
R100 B.n629 B.n35 585
R101 B.n641 B.n35 585
R102 B.n628 B.n34 585
R103 B.n642 B.n34 585
R104 B.n627 B.n33 585
R105 B.n643 B.n33 585
R106 B.n626 B.n625 585
R107 B.n625 B.n32 585
R108 B.n624 B.n28 585
R109 B.n649 B.n28 585
R110 B.n623 B.n27 585
R111 B.n650 B.n27 585
R112 B.n622 B.n26 585
R113 B.n651 B.n26 585
R114 B.n621 B.n620 585
R115 B.n620 B.n22 585
R116 B.n619 B.n21 585
R117 B.n657 B.n21 585
R118 B.n618 B.n20 585
R119 B.n658 B.n20 585
R120 B.n617 B.n19 585
R121 B.n659 B.n19 585
R122 B.n616 B.n615 585
R123 B.n615 B.n15 585
R124 B.n614 B.n14 585
R125 B.n665 B.n14 585
R126 B.n613 B.n13 585
R127 B.n666 B.n13 585
R128 B.n612 B.n12 585
R129 B.n667 B.n12 585
R130 B.n611 B.n610 585
R131 B.n610 B.n11 585
R132 B.n609 B.n7 585
R133 B.n673 B.n7 585
R134 B.n608 B.n6 585
R135 B.n674 B.n6 585
R136 B.n607 B.n5 585
R137 B.n675 B.n5 585
R138 B.n606 B.n605 585
R139 B.n605 B.n4 585
R140 B.n604 B.n274 585
R141 B.n604 B.n603 585
R142 B.n593 B.n275 585
R143 B.n596 B.n275 585
R144 B.n595 B.n594 585
R145 B.n597 B.n595 585
R146 B.n592 B.n280 585
R147 B.n280 B.n279 585
R148 B.n591 B.n590 585
R149 B.n590 B.n589 585
R150 B.n282 B.n281 585
R151 B.n283 B.n282 585
R152 B.n582 B.n581 585
R153 B.n583 B.n582 585
R154 B.n580 B.n287 585
R155 B.n291 B.n287 585
R156 B.n579 B.n578 585
R157 B.n578 B.n577 585
R158 B.n289 B.n288 585
R159 B.n290 B.n289 585
R160 B.n570 B.n569 585
R161 B.n571 B.n570 585
R162 B.n568 B.n296 585
R163 B.n296 B.n295 585
R164 B.n567 B.n566 585
R165 B.n566 B.n565 585
R166 B.n298 B.n297 585
R167 B.n558 B.n298 585
R168 B.n557 B.n556 585
R169 B.n559 B.n557 585
R170 B.n555 B.n303 585
R171 B.n303 B.n302 585
R172 B.n554 B.n553 585
R173 B.n553 B.n552 585
R174 B.n305 B.n304 585
R175 B.n306 B.n305 585
R176 B.n548 B.n547 585
R177 B.n309 B.n308 585
R178 B.n544 B.n543 585
R179 B.n545 B.n544 585
R180 B.n542 B.n356 585
R181 B.n541 B.n540 585
R182 B.n539 B.n538 585
R183 B.n537 B.n536 585
R184 B.n535 B.n534 585
R185 B.n533 B.n532 585
R186 B.n531 B.n530 585
R187 B.n529 B.n528 585
R188 B.n527 B.n526 585
R189 B.n525 B.n524 585
R190 B.n523 B.n522 585
R191 B.n521 B.n520 585
R192 B.n519 B.n518 585
R193 B.n517 B.n516 585
R194 B.n515 B.n514 585
R195 B.n513 B.n512 585
R196 B.n511 B.n510 585
R197 B.n509 B.n508 585
R198 B.n507 B.n506 585
R199 B.n505 B.n504 585
R200 B.n503 B.n502 585
R201 B.n501 B.n500 585
R202 B.n499 B.n498 585
R203 B.n497 B.n496 585
R204 B.n495 B.n494 585
R205 B.n493 B.n492 585
R206 B.n491 B.n490 585
R207 B.n489 B.n488 585
R208 B.n487 B.n486 585
R209 B.n485 B.n484 585
R210 B.n483 B.n482 585
R211 B.n481 B.n480 585
R212 B.n479 B.n478 585
R213 B.n477 B.n476 585
R214 B.n475 B.n474 585
R215 B.n473 B.n472 585
R216 B.n471 B.n470 585
R217 B.n469 B.n468 585
R218 B.n467 B.n466 585
R219 B.n464 B.n463 585
R220 B.n462 B.n461 585
R221 B.n460 B.n459 585
R222 B.n458 B.n457 585
R223 B.n456 B.n455 585
R224 B.n454 B.n453 585
R225 B.n452 B.n451 585
R226 B.n450 B.n449 585
R227 B.n448 B.n447 585
R228 B.n446 B.n445 585
R229 B.n443 B.n442 585
R230 B.n441 B.n440 585
R231 B.n439 B.n438 585
R232 B.n437 B.n436 585
R233 B.n435 B.n434 585
R234 B.n433 B.n432 585
R235 B.n431 B.n430 585
R236 B.n429 B.n428 585
R237 B.n427 B.n426 585
R238 B.n425 B.n424 585
R239 B.n423 B.n422 585
R240 B.n421 B.n420 585
R241 B.n419 B.n418 585
R242 B.n417 B.n416 585
R243 B.n415 B.n414 585
R244 B.n413 B.n412 585
R245 B.n411 B.n410 585
R246 B.n409 B.n408 585
R247 B.n407 B.n406 585
R248 B.n405 B.n404 585
R249 B.n403 B.n402 585
R250 B.n401 B.n400 585
R251 B.n399 B.n398 585
R252 B.n397 B.n396 585
R253 B.n395 B.n394 585
R254 B.n393 B.n392 585
R255 B.n391 B.n390 585
R256 B.n389 B.n388 585
R257 B.n387 B.n386 585
R258 B.n385 B.n384 585
R259 B.n383 B.n382 585
R260 B.n381 B.n380 585
R261 B.n379 B.n378 585
R262 B.n377 B.n376 585
R263 B.n375 B.n374 585
R264 B.n373 B.n372 585
R265 B.n371 B.n370 585
R266 B.n369 B.n368 585
R267 B.n367 B.n366 585
R268 B.n365 B.n364 585
R269 B.n363 B.n362 585
R270 B.n361 B.n355 585
R271 B.n545 B.n355 585
R272 B.n549 B.n307 585
R273 B.n307 B.n306 585
R274 B.n551 B.n550 585
R275 B.n552 B.n551 585
R276 B.n301 B.n300 585
R277 B.n302 B.n301 585
R278 B.n561 B.n560 585
R279 B.n560 B.n559 585
R280 B.n562 B.n299 585
R281 B.n558 B.n299 585
R282 B.n564 B.n563 585
R283 B.n565 B.n564 585
R284 B.n294 B.n293 585
R285 B.n295 B.n294 585
R286 B.n573 B.n572 585
R287 B.n572 B.n571 585
R288 B.n574 B.n292 585
R289 B.n292 B.n290 585
R290 B.n576 B.n575 585
R291 B.n577 B.n576 585
R292 B.n286 B.n285 585
R293 B.n291 B.n286 585
R294 B.n585 B.n584 585
R295 B.n584 B.n583 585
R296 B.n586 B.n284 585
R297 B.n284 B.n283 585
R298 B.n588 B.n587 585
R299 B.n589 B.n588 585
R300 B.n278 B.n277 585
R301 B.n279 B.n278 585
R302 B.n599 B.n598 585
R303 B.n598 B.n597 585
R304 B.n600 B.n276 585
R305 B.n596 B.n276 585
R306 B.n602 B.n601 585
R307 B.n603 B.n602 585
R308 B.n2 B.n0 585
R309 B.n4 B.n2 585
R310 B.n3 B.n1 585
R311 B.n674 B.n3 585
R312 B.n672 B.n671 585
R313 B.n673 B.n672 585
R314 B.n670 B.n8 585
R315 B.n11 B.n8 585
R316 B.n669 B.n668 585
R317 B.n668 B.n667 585
R318 B.n10 B.n9 585
R319 B.n666 B.n10 585
R320 B.n664 B.n663 585
R321 B.n665 B.n664 585
R322 B.n662 B.n16 585
R323 B.n16 B.n15 585
R324 B.n661 B.n660 585
R325 B.n660 B.n659 585
R326 B.n18 B.n17 585
R327 B.n658 B.n18 585
R328 B.n656 B.n655 585
R329 B.n657 B.n656 585
R330 B.n654 B.n23 585
R331 B.n23 B.n22 585
R332 B.n653 B.n652 585
R333 B.n652 B.n651 585
R334 B.n25 B.n24 585
R335 B.n650 B.n25 585
R336 B.n648 B.n647 585
R337 B.n649 B.n648 585
R338 B.n646 B.n29 585
R339 B.n32 B.n29 585
R340 B.n645 B.n644 585
R341 B.n644 B.n643 585
R342 B.n31 B.n30 585
R343 B.n642 B.n31 585
R344 B.n640 B.n639 585
R345 B.n641 B.n640 585
R346 B.n638 B.n37 585
R347 B.n37 B.n36 585
R348 B.n677 B.n676 585
R349 B.n676 B.n675 585
R350 B.n547 B.n307 463.671
R351 B.n636 B.n37 463.671
R352 B.n355 B.n305 463.671
R353 B.n632 B.n86 463.671
R354 B.n359 B.t9 302.76
R355 B.n87 B.t15 302.76
R356 B.n357 B.t19 302.76
R357 B.n90 B.t12 302.76
R358 B.n360 B.t8 284.918
R359 B.n88 B.t16 284.918
R360 B.n358 B.t18 284.918
R361 B.n91 B.t13 284.918
R362 B.n634 B.n633 256.663
R363 B.n634 B.n84 256.663
R364 B.n634 B.n83 256.663
R365 B.n634 B.n82 256.663
R366 B.n634 B.n81 256.663
R367 B.n634 B.n80 256.663
R368 B.n634 B.n79 256.663
R369 B.n634 B.n78 256.663
R370 B.n634 B.n77 256.663
R371 B.n634 B.n76 256.663
R372 B.n634 B.n75 256.663
R373 B.n634 B.n74 256.663
R374 B.n634 B.n73 256.663
R375 B.n634 B.n72 256.663
R376 B.n634 B.n71 256.663
R377 B.n634 B.n70 256.663
R378 B.n634 B.n69 256.663
R379 B.n634 B.n68 256.663
R380 B.n634 B.n67 256.663
R381 B.n634 B.n66 256.663
R382 B.n634 B.n65 256.663
R383 B.n634 B.n64 256.663
R384 B.n634 B.n63 256.663
R385 B.n634 B.n62 256.663
R386 B.n634 B.n61 256.663
R387 B.n634 B.n60 256.663
R388 B.n634 B.n59 256.663
R389 B.n634 B.n58 256.663
R390 B.n634 B.n57 256.663
R391 B.n634 B.n56 256.663
R392 B.n634 B.n55 256.663
R393 B.n634 B.n54 256.663
R394 B.n634 B.n53 256.663
R395 B.n634 B.n52 256.663
R396 B.n634 B.n51 256.663
R397 B.n634 B.n50 256.663
R398 B.n634 B.n49 256.663
R399 B.n634 B.n48 256.663
R400 B.n634 B.n47 256.663
R401 B.n634 B.n46 256.663
R402 B.n634 B.n45 256.663
R403 B.n634 B.n44 256.663
R404 B.n634 B.n43 256.663
R405 B.n634 B.n42 256.663
R406 B.n634 B.n41 256.663
R407 B.n634 B.n40 256.663
R408 B.n635 B.n634 256.663
R409 B.n546 B.n545 256.663
R410 B.n545 B.n310 256.663
R411 B.n545 B.n311 256.663
R412 B.n545 B.n312 256.663
R413 B.n545 B.n313 256.663
R414 B.n545 B.n314 256.663
R415 B.n545 B.n315 256.663
R416 B.n545 B.n316 256.663
R417 B.n545 B.n317 256.663
R418 B.n545 B.n318 256.663
R419 B.n545 B.n319 256.663
R420 B.n545 B.n320 256.663
R421 B.n545 B.n321 256.663
R422 B.n545 B.n322 256.663
R423 B.n545 B.n323 256.663
R424 B.n545 B.n324 256.663
R425 B.n545 B.n325 256.663
R426 B.n545 B.n326 256.663
R427 B.n545 B.n327 256.663
R428 B.n545 B.n328 256.663
R429 B.n545 B.n329 256.663
R430 B.n545 B.n330 256.663
R431 B.n545 B.n331 256.663
R432 B.n545 B.n332 256.663
R433 B.n545 B.n333 256.663
R434 B.n545 B.n334 256.663
R435 B.n545 B.n335 256.663
R436 B.n545 B.n336 256.663
R437 B.n545 B.n337 256.663
R438 B.n545 B.n338 256.663
R439 B.n545 B.n339 256.663
R440 B.n545 B.n340 256.663
R441 B.n545 B.n341 256.663
R442 B.n545 B.n342 256.663
R443 B.n545 B.n343 256.663
R444 B.n545 B.n344 256.663
R445 B.n545 B.n345 256.663
R446 B.n545 B.n346 256.663
R447 B.n545 B.n347 256.663
R448 B.n545 B.n348 256.663
R449 B.n545 B.n349 256.663
R450 B.n545 B.n350 256.663
R451 B.n545 B.n351 256.663
R452 B.n545 B.n352 256.663
R453 B.n545 B.n353 256.663
R454 B.n545 B.n354 256.663
R455 B.n551 B.n307 163.367
R456 B.n551 B.n301 163.367
R457 B.n560 B.n301 163.367
R458 B.n560 B.n299 163.367
R459 B.n564 B.n299 163.367
R460 B.n564 B.n294 163.367
R461 B.n572 B.n294 163.367
R462 B.n572 B.n292 163.367
R463 B.n576 B.n292 163.367
R464 B.n576 B.n286 163.367
R465 B.n584 B.n286 163.367
R466 B.n584 B.n284 163.367
R467 B.n588 B.n284 163.367
R468 B.n588 B.n278 163.367
R469 B.n598 B.n278 163.367
R470 B.n598 B.n276 163.367
R471 B.n602 B.n276 163.367
R472 B.n602 B.n2 163.367
R473 B.n676 B.n2 163.367
R474 B.n676 B.n3 163.367
R475 B.n672 B.n3 163.367
R476 B.n672 B.n8 163.367
R477 B.n668 B.n8 163.367
R478 B.n668 B.n10 163.367
R479 B.n664 B.n10 163.367
R480 B.n664 B.n16 163.367
R481 B.n660 B.n16 163.367
R482 B.n660 B.n18 163.367
R483 B.n656 B.n18 163.367
R484 B.n656 B.n23 163.367
R485 B.n652 B.n23 163.367
R486 B.n652 B.n25 163.367
R487 B.n648 B.n25 163.367
R488 B.n648 B.n29 163.367
R489 B.n644 B.n29 163.367
R490 B.n644 B.n31 163.367
R491 B.n640 B.n31 163.367
R492 B.n640 B.n37 163.367
R493 B.n544 B.n309 163.367
R494 B.n544 B.n356 163.367
R495 B.n540 B.n539 163.367
R496 B.n536 B.n535 163.367
R497 B.n532 B.n531 163.367
R498 B.n528 B.n527 163.367
R499 B.n524 B.n523 163.367
R500 B.n520 B.n519 163.367
R501 B.n516 B.n515 163.367
R502 B.n512 B.n511 163.367
R503 B.n508 B.n507 163.367
R504 B.n504 B.n503 163.367
R505 B.n500 B.n499 163.367
R506 B.n496 B.n495 163.367
R507 B.n492 B.n491 163.367
R508 B.n488 B.n487 163.367
R509 B.n484 B.n483 163.367
R510 B.n480 B.n479 163.367
R511 B.n476 B.n475 163.367
R512 B.n472 B.n471 163.367
R513 B.n468 B.n467 163.367
R514 B.n463 B.n462 163.367
R515 B.n459 B.n458 163.367
R516 B.n455 B.n454 163.367
R517 B.n451 B.n450 163.367
R518 B.n447 B.n446 163.367
R519 B.n442 B.n441 163.367
R520 B.n438 B.n437 163.367
R521 B.n434 B.n433 163.367
R522 B.n430 B.n429 163.367
R523 B.n426 B.n425 163.367
R524 B.n422 B.n421 163.367
R525 B.n418 B.n417 163.367
R526 B.n414 B.n413 163.367
R527 B.n410 B.n409 163.367
R528 B.n406 B.n405 163.367
R529 B.n402 B.n401 163.367
R530 B.n398 B.n397 163.367
R531 B.n394 B.n393 163.367
R532 B.n390 B.n389 163.367
R533 B.n386 B.n385 163.367
R534 B.n382 B.n381 163.367
R535 B.n378 B.n377 163.367
R536 B.n374 B.n373 163.367
R537 B.n370 B.n369 163.367
R538 B.n366 B.n365 163.367
R539 B.n362 B.n355 163.367
R540 B.n553 B.n305 163.367
R541 B.n553 B.n303 163.367
R542 B.n557 B.n303 163.367
R543 B.n557 B.n298 163.367
R544 B.n566 B.n298 163.367
R545 B.n566 B.n296 163.367
R546 B.n570 B.n296 163.367
R547 B.n570 B.n289 163.367
R548 B.n578 B.n289 163.367
R549 B.n578 B.n287 163.367
R550 B.n582 B.n287 163.367
R551 B.n582 B.n282 163.367
R552 B.n590 B.n282 163.367
R553 B.n590 B.n280 163.367
R554 B.n595 B.n280 163.367
R555 B.n595 B.n275 163.367
R556 B.n604 B.n275 163.367
R557 B.n605 B.n604 163.367
R558 B.n605 B.n5 163.367
R559 B.n6 B.n5 163.367
R560 B.n7 B.n6 163.367
R561 B.n610 B.n7 163.367
R562 B.n610 B.n12 163.367
R563 B.n13 B.n12 163.367
R564 B.n14 B.n13 163.367
R565 B.n615 B.n14 163.367
R566 B.n615 B.n19 163.367
R567 B.n20 B.n19 163.367
R568 B.n21 B.n20 163.367
R569 B.n620 B.n21 163.367
R570 B.n620 B.n26 163.367
R571 B.n27 B.n26 163.367
R572 B.n28 B.n27 163.367
R573 B.n625 B.n28 163.367
R574 B.n625 B.n33 163.367
R575 B.n34 B.n33 163.367
R576 B.n35 B.n34 163.367
R577 B.n86 B.n35 163.367
R578 B.n93 B.n39 163.367
R579 B.n97 B.n96 163.367
R580 B.n101 B.n100 163.367
R581 B.n105 B.n104 163.367
R582 B.n109 B.n108 163.367
R583 B.n113 B.n112 163.367
R584 B.n117 B.n116 163.367
R585 B.n121 B.n120 163.367
R586 B.n125 B.n124 163.367
R587 B.n129 B.n128 163.367
R588 B.n133 B.n132 163.367
R589 B.n137 B.n136 163.367
R590 B.n141 B.n140 163.367
R591 B.n145 B.n144 163.367
R592 B.n149 B.n148 163.367
R593 B.n153 B.n152 163.367
R594 B.n157 B.n156 163.367
R595 B.n161 B.n160 163.367
R596 B.n165 B.n164 163.367
R597 B.n169 B.n168 163.367
R598 B.n173 B.n172 163.367
R599 B.n177 B.n176 163.367
R600 B.n181 B.n180 163.367
R601 B.n185 B.n184 163.367
R602 B.n189 B.n188 163.367
R603 B.n193 B.n192 163.367
R604 B.n197 B.n196 163.367
R605 B.n201 B.n200 163.367
R606 B.n205 B.n204 163.367
R607 B.n209 B.n208 163.367
R608 B.n213 B.n212 163.367
R609 B.n217 B.n216 163.367
R610 B.n221 B.n220 163.367
R611 B.n225 B.n224 163.367
R612 B.n229 B.n228 163.367
R613 B.n233 B.n232 163.367
R614 B.n237 B.n236 163.367
R615 B.n241 B.n240 163.367
R616 B.n245 B.n244 163.367
R617 B.n249 B.n248 163.367
R618 B.n253 B.n252 163.367
R619 B.n257 B.n256 163.367
R620 B.n261 B.n260 163.367
R621 B.n265 B.n264 163.367
R622 B.n269 B.n268 163.367
R623 B.n271 B.n85 163.367
R624 B.n545 B.n306 75.1225
R625 B.n634 B.n36 75.1225
R626 B.n547 B.n546 71.676
R627 B.n356 B.n310 71.676
R628 B.n539 B.n311 71.676
R629 B.n535 B.n312 71.676
R630 B.n531 B.n313 71.676
R631 B.n527 B.n314 71.676
R632 B.n523 B.n315 71.676
R633 B.n519 B.n316 71.676
R634 B.n515 B.n317 71.676
R635 B.n511 B.n318 71.676
R636 B.n507 B.n319 71.676
R637 B.n503 B.n320 71.676
R638 B.n499 B.n321 71.676
R639 B.n495 B.n322 71.676
R640 B.n491 B.n323 71.676
R641 B.n487 B.n324 71.676
R642 B.n483 B.n325 71.676
R643 B.n479 B.n326 71.676
R644 B.n475 B.n327 71.676
R645 B.n471 B.n328 71.676
R646 B.n467 B.n329 71.676
R647 B.n462 B.n330 71.676
R648 B.n458 B.n331 71.676
R649 B.n454 B.n332 71.676
R650 B.n450 B.n333 71.676
R651 B.n446 B.n334 71.676
R652 B.n441 B.n335 71.676
R653 B.n437 B.n336 71.676
R654 B.n433 B.n337 71.676
R655 B.n429 B.n338 71.676
R656 B.n425 B.n339 71.676
R657 B.n421 B.n340 71.676
R658 B.n417 B.n341 71.676
R659 B.n413 B.n342 71.676
R660 B.n409 B.n343 71.676
R661 B.n405 B.n344 71.676
R662 B.n401 B.n345 71.676
R663 B.n397 B.n346 71.676
R664 B.n393 B.n347 71.676
R665 B.n389 B.n348 71.676
R666 B.n385 B.n349 71.676
R667 B.n381 B.n350 71.676
R668 B.n377 B.n351 71.676
R669 B.n373 B.n352 71.676
R670 B.n369 B.n353 71.676
R671 B.n365 B.n354 71.676
R672 B.n636 B.n635 71.676
R673 B.n93 B.n40 71.676
R674 B.n97 B.n41 71.676
R675 B.n101 B.n42 71.676
R676 B.n105 B.n43 71.676
R677 B.n109 B.n44 71.676
R678 B.n113 B.n45 71.676
R679 B.n117 B.n46 71.676
R680 B.n121 B.n47 71.676
R681 B.n125 B.n48 71.676
R682 B.n129 B.n49 71.676
R683 B.n133 B.n50 71.676
R684 B.n137 B.n51 71.676
R685 B.n141 B.n52 71.676
R686 B.n145 B.n53 71.676
R687 B.n149 B.n54 71.676
R688 B.n153 B.n55 71.676
R689 B.n157 B.n56 71.676
R690 B.n161 B.n57 71.676
R691 B.n165 B.n58 71.676
R692 B.n169 B.n59 71.676
R693 B.n173 B.n60 71.676
R694 B.n177 B.n61 71.676
R695 B.n181 B.n62 71.676
R696 B.n185 B.n63 71.676
R697 B.n189 B.n64 71.676
R698 B.n193 B.n65 71.676
R699 B.n197 B.n66 71.676
R700 B.n201 B.n67 71.676
R701 B.n205 B.n68 71.676
R702 B.n209 B.n69 71.676
R703 B.n213 B.n70 71.676
R704 B.n217 B.n71 71.676
R705 B.n221 B.n72 71.676
R706 B.n225 B.n73 71.676
R707 B.n229 B.n74 71.676
R708 B.n233 B.n75 71.676
R709 B.n237 B.n76 71.676
R710 B.n241 B.n77 71.676
R711 B.n245 B.n78 71.676
R712 B.n249 B.n79 71.676
R713 B.n253 B.n80 71.676
R714 B.n257 B.n81 71.676
R715 B.n261 B.n82 71.676
R716 B.n265 B.n83 71.676
R717 B.n269 B.n84 71.676
R718 B.n633 B.n85 71.676
R719 B.n633 B.n632 71.676
R720 B.n271 B.n84 71.676
R721 B.n268 B.n83 71.676
R722 B.n264 B.n82 71.676
R723 B.n260 B.n81 71.676
R724 B.n256 B.n80 71.676
R725 B.n252 B.n79 71.676
R726 B.n248 B.n78 71.676
R727 B.n244 B.n77 71.676
R728 B.n240 B.n76 71.676
R729 B.n236 B.n75 71.676
R730 B.n232 B.n74 71.676
R731 B.n228 B.n73 71.676
R732 B.n224 B.n72 71.676
R733 B.n220 B.n71 71.676
R734 B.n216 B.n70 71.676
R735 B.n212 B.n69 71.676
R736 B.n208 B.n68 71.676
R737 B.n204 B.n67 71.676
R738 B.n200 B.n66 71.676
R739 B.n196 B.n65 71.676
R740 B.n192 B.n64 71.676
R741 B.n188 B.n63 71.676
R742 B.n184 B.n62 71.676
R743 B.n180 B.n61 71.676
R744 B.n176 B.n60 71.676
R745 B.n172 B.n59 71.676
R746 B.n168 B.n58 71.676
R747 B.n164 B.n57 71.676
R748 B.n160 B.n56 71.676
R749 B.n156 B.n55 71.676
R750 B.n152 B.n54 71.676
R751 B.n148 B.n53 71.676
R752 B.n144 B.n52 71.676
R753 B.n140 B.n51 71.676
R754 B.n136 B.n50 71.676
R755 B.n132 B.n49 71.676
R756 B.n128 B.n48 71.676
R757 B.n124 B.n47 71.676
R758 B.n120 B.n46 71.676
R759 B.n116 B.n45 71.676
R760 B.n112 B.n44 71.676
R761 B.n108 B.n43 71.676
R762 B.n104 B.n42 71.676
R763 B.n100 B.n41 71.676
R764 B.n96 B.n40 71.676
R765 B.n635 B.n39 71.676
R766 B.n546 B.n309 71.676
R767 B.n540 B.n310 71.676
R768 B.n536 B.n311 71.676
R769 B.n532 B.n312 71.676
R770 B.n528 B.n313 71.676
R771 B.n524 B.n314 71.676
R772 B.n520 B.n315 71.676
R773 B.n516 B.n316 71.676
R774 B.n512 B.n317 71.676
R775 B.n508 B.n318 71.676
R776 B.n504 B.n319 71.676
R777 B.n500 B.n320 71.676
R778 B.n496 B.n321 71.676
R779 B.n492 B.n322 71.676
R780 B.n488 B.n323 71.676
R781 B.n484 B.n324 71.676
R782 B.n480 B.n325 71.676
R783 B.n476 B.n326 71.676
R784 B.n472 B.n327 71.676
R785 B.n468 B.n328 71.676
R786 B.n463 B.n329 71.676
R787 B.n459 B.n330 71.676
R788 B.n455 B.n331 71.676
R789 B.n451 B.n332 71.676
R790 B.n447 B.n333 71.676
R791 B.n442 B.n334 71.676
R792 B.n438 B.n335 71.676
R793 B.n434 B.n336 71.676
R794 B.n430 B.n337 71.676
R795 B.n426 B.n338 71.676
R796 B.n422 B.n339 71.676
R797 B.n418 B.n340 71.676
R798 B.n414 B.n341 71.676
R799 B.n410 B.n342 71.676
R800 B.n406 B.n343 71.676
R801 B.n402 B.n344 71.676
R802 B.n398 B.n345 71.676
R803 B.n394 B.n346 71.676
R804 B.n390 B.n347 71.676
R805 B.n386 B.n348 71.676
R806 B.n382 B.n349 71.676
R807 B.n378 B.n350 71.676
R808 B.n374 B.n351 71.676
R809 B.n370 B.n352 71.676
R810 B.n366 B.n353 71.676
R811 B.n362 B.n354 71.676
R812 B.n444 B.n360 59.5399
R813 B.n465 B.n358 59.5399
R814 B.n92 B.n91 59.5399
R815 B.n89 B.n88 59.5399
R816 B.n552 B.n306 42.9273
R817 B.n552 B.n302 42.9273
R818 B.n559 B.n302 42.9273
R819 B.n559 B.n558 42.9273
R820 B.n565 B.n295 42.9273
R821 B.n571 B.n295 42.9273
R822 B.n571 B.n290 42.9273
R823 B.n577 B.n290 42.9273
R824 B.n577 B.n291 42.9273
R825 B.n583 B.n283 42.9273
R826 B.n589 B.n283 42.9273
R827 B.n597 B.n279 42.9273
R828 B.n597 B.n596 42.9273
R829 B.n603 B.n4 42.9273
R830 B.n675 B.n4 42.9273
R831 B.n675 B.n674 42.9273
R832 B.n674 B.n673 42.9273
R833 B.n667 B.n11 42.9273
R834 B.n667 B.n666 42.9273
R835 B.n665 B.n15 42.9273
R836 B.n659 B.n15 42.9273
R837 B.n658 B.n657 42.9273
R838 B.n657 B.n22 42.9273
R839 B.n651 B.n22 42.9273
R840 B.n651 B.n650 42.9273
R841 B.n650 B.n649 42.9273
R842 B.n643 B.n32 42.9273
R843 B.n643 B.n642 42.9273
R844 B.n642 B.n641 42.9273
R845 B.n641 B.n36 42.9273
R846 B.n603 B.t1 41.0335
R847 B.n673 B.t3 41.0335
R848 B.n558 B.t7 30.9331
R849 B.n32 B.t11 30.9331
R850 B.n638 B.n637 30.1273
R851 B.n631 B.n630 30.1273
R852 B.n361 B.n304 30.1273
R853 B.n549 B.n548 30.1273
R854 B.t2 B.n279 28.408
R855 B.n666 B.t0 28.408
R856 B.n291 B.t5 27.1454
R857 B.t4 B.n658 27.1454
R858 B B.n677 18.0485
R859 B.n360 B.n359 17.8429
R860 B.n358 B.n357 17.8429
R861 B.n91 B.n90 17.8429
R862 B.n88 B.n87 17.8429
R863 B.n583 B.t5 15.7824
R864 B.n659 B.t4 15.7824
R865 B.n589 B.t2 14.5199
R866 B.t0 B.n665 14.5199
R867 B.n565 B.t7 11.9948
R868 B.n649 B.t11 11.9948
R869 B.n637 B.n38 10.6151
R870 B.n94 B.n38 10.6151
R871 B.n95 B.n94 10.6151
R872 B.n98 B.n95 10.6151
R873 B.n99 B.n98 10.6151
R874 B.n102 B.n99 10.6151
R875 B.n103 B.n102 10.6151
R876 B.n106 B.n103 10.6151
R877 B.n107 B.n106 10.6151
R878 B.n110 B.n107 10.6151
R879 B.n111 B.n110 10.6151
R880 B.n114 B.n111 10.6151
R881 B.n115 B.n114 10.6151
R882 B.n118 B.n115 10.6151
R883 B.n119 B.n118 10.6151
R884 B.n122 B.n119 10.6151
R885 B.n123 B.n122 10.6151
R886 B.n126 B.n123 10.6151
R887 B.n127 B.n126 10.6151
R888 B.n130 B.n127 10.6151
R889 B.n131 B.n130 10.6151
R890 B.n134 B.n131 10.6151
R891 B.n135 B.n134 10.6151
R892 B.n138 B.n135 10.6151
R893 B.n139 B.n138 10.6151
R894 B.n142 B.n139 10.6151
R895 B.n143 B.n142 10.6151
R896 B.n146 B.n143 10.6151
R897 B.n147 B.n146 10.6151
R898 B.n150 B.n147 10.6151
R899 B.n151 B.n150 10.6151
R900 B.n154 B.n151 10.6151
R901 B.n155 B.n154 10.6151
R902 B.n158 B.n155 10.6151
R903 B.n159 B.n158 10.6151
R904 B.n162 B.n159 10.6151
R905 B.n163 B.n162 10.6151
R906 B.n166 B.n163 10.6151
R907 B.n167 B.n166 10.6151
R908 B.n170 B.n167 10.6151
R909 B.n171 B.n170 10.6151
R910 B.n175 B.n174 10.6151
R911 B.n178 B.n175 10.6151
R912 B.n179 B.n178 10.6151
R913 B.n182 B.n179 10.6151
R914 B.n183 B.n182 10.6151
R915 B.n186 B.n183 10.6151
R916 B.n187 B.n186 10.6151
R917 B.n190 B.n187 10.6151
R918 B.n191 B.n190 10.6151
R919 B.n195 B.n194 10.6151
R920 B.n198 B.n195 10.6151
R921 B.n199 B.n198 10.6151
R922 B.n202 B.n199 10.6151
R923 B.n203 B.n202 10.6151
R924 B.n206 B.n203 10.6151
R925 B.n207 B.n206 10.6151
R926 B.n210 B.n207 10.6151
R927 B.n211 B.n210 10.6151
R928 B.n214 B.n211 10.6151
R929 B.n215 B.n214 10.6151
R930 B.n218 B.n215 10.6151
R931 B.n219 B.n218 10.6151
R932 B.n222 B.n219 10.6151
R933 B.n223 B.n222 10.6151
R934 B.n226 B.n223 10.6151
R935 B.n227 B.n226 10.6151
R936 B.n230 B.n227 10.6151
R937 B.n231 B.n230 10.6151
R938 B.n234 B.n231 10.6151
R939 B.n235 B.n234 10.6151
R940 B.n238 B.n235 10.6151
R941 B.n239 B.n238 10.6151
R942 B.n242 B.n239 10.6151
R943 B.n243 B.n242 10.6151
R944 B.n246 B.n243 10.6151
R945 B.n247 B.n246 10.6151
R946 B.n250 B.n247 10.6151
R947 B.n251 B.n250 10.6151
R948 B.n254 B.n251 10.6151
R949 B.n255 B.n254 10.6151
R950 B.n258 B.n255 10.6151
R951 B.n259 B.n258 10.6151
R952 B.n262 B.n259 10.6151
R953 B.n263 B.n262 10.6151
R954 B.n266 B.n263 10.6151
R955 B.n267 B.n266 10.6151
R956 B.n270 B.n267 10.6151
R957 B.n272 B.n270 10.6151
R958 B.n273 B.n272 10.6151
R959 B.n631 B.n273 10.6151
R960 B.n554 B.n304 10.6151
R961 B.n555 B.n554 10.6151
R962 B.n556 B.n555 10.6151
R963 B.n556 B.n297 10.6151
R964 B.n567 B.n297 10.6151
R965 B.n568 B.n567 10.6151
R966 B.n569 B.n568 10.6151
R967 B.n569 B.n288 10.6151
R968 B.n579 B.n288 10.6151
R969 B.n580 B.n579 10.6151
R970 B.n581 B.n580 10.6151
R971 B.n581 B.n281 10.6151
R972 B.n591 B.n281 10.6151
R973 B.n592 B.n591 10.6151
R974 B.n594 B.n592 10.6151
R975 B.n594 B.n593 10.6151
R976 B.n593 B.n274 10.6151
R977 B.n606 B.n274 10.6151
R978 B.n607 B.n606 10.6151
R979 B.n608 B.n607 10.6151
R980 B.n609 B.n608 10.6151
R981 B.n611 B.n609 10.6151
R982 B.n612 B.n611 10.6151
R983 B.n613 B.n612 10.6151
R984 B.n614 B.n613 10.6151
R985 B.n616 B.n614 10.6151
R986 B.n617 B.n616 10.6151
R987 B.n618 B.n617 10.6151
R988 B.n619 B.n618 10.6151
R989 B.n621 B.n619 10.6151
R990 B.n622 B.n621 10.6151
R991 B.n623 B.n622 10.6151
R992 B.n624 B.n623 10.6151
R993 B.n626 B.n624 10.6151
R994 B.n627 B.n626 10.6151
R995 B.n628 B.n627 10.6151
R996 B.n629 B.n628 10.6151
R997 B.n630 B.n629 10.6151
R998 B.n548 B.n308 10.6151
R999 B.n543 B.n308 10.6151
R1000 B.n543 B.n542 10.6151
R1001 B.n542 B.n541 10.6151
R1002 B.n541 B.n538 10.6151
R1003 B.n538 B.n537 10.6151
R1004 B.n537 B.n534 10.6151
R1005 B.n534 B.n533 10.6151
R1006 B.n533 B.n530 10.6151
R1007 B.n530 B.n529 10.6151
R1008 B.n529 B.n526 10.6151
R1009 B.n526 B.n525 10.6151
R1010 B.n525 B.n522 10.6151
R1011 B.n522 B.n521 10.6151
R1012 B.n521 B.n518 10.6151
R1013 B.n518 B.n517 10.6151
R1014 B.n517 B.n514 10.6151
R1015 B.n514 B.n513 10.6151
R1016 B.n513 B.n510 10.6151
R1017 B.n510 B.n509 10.6151
R1018 B.n509 B.n506 10.6151
R1019 B.n506 B.n505 10.6151
R1020 B.n505 B.n502 10.6151
R1021 B.n502 B.n501 10.6151
R1022 B.n501 B.n498 10.6151
R1023 B.n498 B.n497 10.6151
R1024 B.n497 B.n494 10.6151
R1025 B.n494 B.n493 10.6151
R1026 B.n493 B.n490 10.6151
R1027 B.n490 B.n489 10.6151
R1028 B.n489 B.n486 10.6151
R1029 B.n486 B.n485 10.6151
R1030 B.n485 B.n482 10.6151
R1031 B.n482 B.n481 10.6151
R1032 B.n481 B.n478 10.6151
R1033 B.n478 B.n477 10.6151
R1034 B.n477 B.n474 10.6151
R1035 B.n474 B.n473 10.6151
R1036 B.n473 B.n470 10.6151
R1037 B.n470 B.n469 10.6151
R1038 B.n469 B.n466 10.6151
R1039 B.n464 B.n461 10.6151
R1040 B.n461 B.n460 10.6151
R1041 B.n460 B.n457 10.6151
R1042 B.n457 B.n456 10.6151
R1043 B.n456 B.n453 10.6151
R1044 B.n453 B.n452 10.6151
R1045 B.n452 B.n449 10.6151
R1046 B.n449 B.n448 10.6151
R1047 B.n448 B.n445 10.6151
R1048 B.n443 B.n440 10.6151
R1049 B.n440 B.n439 10.6151
R1050 B.n439 B.n436 10.6151
R1051 B.n436 B.n435 10.6151
R1052 B.n435 B.n432 10.6151
R1053 B.n432 B.n431 10.6151
R1054 B.n431 B.n428 10.6151
R1055 B.n428 B.n427 10.6151
R1056 B.n427 B.n424 10.6151
R1057 B.n424 B.n423 10.6151
R1058 B.n423 B.n420 10.6151
R1059 B.n420 B.n419 10.6151
R1060 B.n419 B.n416 10.6151
R1061 B.n416 B.n415 10.6151
R1062 B.n415 B.n412 10.6151
R1063 B.n412 B.n411 10.6151
R1064 B.n411 B.n408 10.6151
R1065 B.n408 B.n407 10.6151
R1066 B.n407 B.n404 10.6151
R1067 B.n404 B.n403 10.6151
R1068 B.n403 B.n400 10.6151
R1069 B.n400 B.n399 10.6151
R1070 B.n399 B.n396 10.6151
R1071 B.n396 B.n395 10.6151
R1072 B.n395 B.n392 10.6151
R1073 B.n392 B.n391 10.6151
R1074 B.n391 B.n388 10.6151
R1075 B.n388 B.n387 10.6151
R1076 B.n387 B.n384 10.6151
R1077 B.n384 B.n383 10.6151
R1078 B.n383 B.n380 10.6151
R1079 B.n380 B.n379 10.6151
R1080 B.n379 B.n376 10.6151
R1081 B.n376 B.n375 10.6151
R1082 B.n375 B.n372 10.6151
R1083 B.n372 B.n371 10.6151
R1084 B.n371 B.n368 10.6151
R1085 B.n368 B.n367 10.6151
R1086 B.n367 B.n364 10.6151
R1087 B.n364 B.n363 10.6151
R1088 B.n363 B.n361 10.6151
R1089 B.n550 B.n549 10.6151
R1090 B.n550 B.n300 10.6151
R1091 B.n561 B.n300 10.6151
R1092 B.n562 B.n561 10.6151
R1093 B.n563 B.n562 10.6151
R1094 B.n563 B.n293 10.6151
R1095 B.n573 B.n293 10.6151
R1096 B.n574 B.n573 10.6151
R1097 B.n575 B.n574 10.6151
R1098 B.n575 B.n285 10.6151
R1099 B.n585 B.n285 10.6151
R1100 B.n586 B.n585 10.6151
R1101 B.n587 B.n586 10.6151
R1102 B.n587 B.n277 10.6151
R1103 B.n599 B.n277 10.6151
R1104 B.n600 B.n599 10.6151
R1105 B.n601 B.n600 10.6151
R1106 B.n601 B.n0 10.6151
R1107 B.n671 B.n1 10.6151
R1108 B.n671 B.n670 10.6151
R1109 B.n670 B.n669 10.6151
R1110 B.n669 B.n9 10.6151
R1111 B.n663 B.n9 10.6151
R1112 B.n663 B.n662 10.6151
R1113 B.n662 B.n661 10.6151
R1114 B.n661 B.n17 10.6151
R1115 B.n655 B.n17 10.6151
R1116 B.n655 B.n654 10.6151
R1117 B.n654 B.n653 10.6151
R1118 B.n653 B.n24 10.6151
R1119 B.n647 B.n24 10.6151
R1120 B.n647 B.n646 10.6151
R1121 B.n646 B.n645 10.6151
R1122 B.n645 B.n30 10.6151
R1123 B.n639 B.n30 10.6151
R1124 B.n639 B.n638 10.6151
R1125 B.n171 B.n92 9.36635
R1126 B.n194 B.n89 9.36635
R1127 B.n466 B.n465 9.36635
R1128 B.n444 B.n443 9.36635
R1129 B.n677 B.n0 2.81026
R1130 B.n677 B.n1 2.81026
R1131 B.n596 B.t1 1.89433
R1132 B.n11 B.t3 1.89433
R1133 B.n174 B.n92 1.24928
R1134 B.n191 B.n89 1.24928
R1135 B.n465 B.n464 1.24928
R1136 B.n445 B.n444 1.24928
R1137 VN.n0 VN.t3 590.109
R1138 VN.n4 VN.t4 590.109
R1139 VN.n1 VN.t0 563.287
R1140 VN.n2 VN.t1 563.287
R1141 VN.n5 VN.t2 563.287
R1142 VN.n6 VN.t5 563.287
R1143 VN.n3 VN.n2 161.3
R1144 VN.n7 VN.n6 161.3
R1145 VN.n2 VN.n1 48.2005
R1146 VN.n6 VN.n5 48.2005
R1147 VN.n7 VN.n4 45.1367
R1148 VN.n3 VN.n0 45.1367
R1149 VN VN.n7 41.3433
R1150 VN.n5 VN.n4 13.3799
R1151 VN.n1 VN.n0 13.3799
R1152 VN VN.n3 0.0516364
R1153 VDD2.n127 VDD2.n67 289.615
R1154 VDD2.n60 VDD2.n0 289.615
R1155 VDD2.n128 VDD2.n127 185
R1156 VDD2.n126 VDD2.n125 185
R1157 VDD2.n71 VDD2.n70 185
R1158 VDD2.n120 VDD2.n119 185
R1159 VDD2.n118 VDD2.n117 185
R1160 VDD2.n75 VDD2.n74 185
R1161 VDD2.n112 VDD2.n111 185
R1162 VDD2.n110 VDD2.n77 185
R1163 VDD2.n109 VDD2.n108 185
R1164 VDD2.n80 VDD2.n78 185
R1165 VDD2.n103 VDD2.n102 185
R1166 VDD2.n101 VDD2.n100 185
R1167 VDD2.n84 VDD2.n83 185
R1168 VDD2.n95 VDD2.n94 185
R1169 VDD2.n93 VDD2.n92 185
R1170 VDD2.n88 VDD2.n87 185
R1171 VDD2.n20 VDD2.n19 185
R1172 VDD2.n25 VDD2.n24 185
R1173 VDD2.n27 VDD2.n26 185
R1174 VDD2.n16 VDD2.n15 185
R1175 VDD2.n33 VDD2.n32 185
R1176 VDD2.n35 VDD2.n34 185
R1177 VDD2.n12 VDD2.n11 185
R1178 VDD2.n42 VDD2.n41 185
R1179 VDD2.n43 VDD2.n10 185
R1180 VDD2.n45 VDD2.n44 185
R1181 VDD2.n8 VDD2.n7 185
R1182 VDD2.n51 VDD2.n50 185
R1183 VDD2.n53 VDD2.n52 185
R1184 VDD2.n4 VDD2.n3 185
R1185 VDD2.n59 VDD2.n58 185
R1186 VDD2.n61 VDD2.n60 185
R1187 VDD2.n89 VDD2.t5 149.524
R1188 VDD2.n21 VDD2.t1 149.524
R1189 VDD2.n127 VDD2.n126 104.615
R1190 VDD2.n126 VDD2.n70 104.615
R1191 VDD2.n119 VDD2.n70 104.615
R1192 VDD2.n119 VDD2.n118 104.615
R1193 VDD2.n118 VDD2.n74 104.615
R1194 VDD2.n111 VDD2.n74 104.615
R1195 VDD2.n111 VDD2.n110 104.615
R1196 VDD2.n110 VDD2.n109 104.615
R1197 VDD2.n109 VDD2.n78 104.615
R1198 VDD2.n102 VDD2.n78 104.615
R1199 VDD2.n102 VDD2.n101 104.615
R1200 VDD2.n101 VDD2.n83 104.615
R1201 VDD2.n94 VDD2.n83 104.615
R1202 VDD2.n94 VDD2.n93 104.615
R1203 VDD2.n93 VDD2.n87 104.615
R1204 VDD2.n25 VDD2.n19 104.615
R1205 VDD2.n26 VDD2.n25 104.615
R1206 VDD2.n26 VDD2.n15 104.615
R1207 VDD2.n33 VDD2.n15 104.615
R1208 VDD2.n34 VDD2.n33 104.615
R1209 VDD2.n34 VDD2.n11 104.615
R1210 VDD2.n42 VDD2.n11 104.615
R1211 VDD2.n43 VDD2.n42 104.615
R1212 VDD2.n44 VDD2.n43 104.615
R1213 VDD2.n44 VDD2.n7 104.615
R1214 VDD2.n51 VDD2.n7 104.615
R1215 VDD2.n52 VDD2.n51 104.615
R1216 VDD2.n52 VDD2.n3 104.615
R1217 VDD2.n59 VDD2.n3 104.615
R1218 VDD2.n60 VDD2.n59 104.615
R1219 VDD2.n66 VDD2.n65 62.6045
R1220 VDD2 VDD2.n133 62.6017
R1221 VDD2.t5 VDD2.n87 52.3082
R1222 VDD2.t1 VDD2.n19 52.3082
R1223 VDD2.n66 VDD2.n64 49.9854
R1224 VDD2.n132 VDD2.n131 49.446
R1225 VDD2.n132 VDD2.n66 36.767
R1226 VDD2.n112 VDD2.n77 13.1884
R1227 VDD2.n45 VDD2.n10 13.1884
R1228 VDD2.n113 VDD2.n75 12.8005
R1229 VDD2.n108 VDD2.n79 12.8005
R1230 VDD2.n41 VDD2.n40 12.8005
R1231 VDD2.n46 VDD2.n8 12.8005
R1232 VDD2.n117 VDD2.n116 12.0247
R1233 VDD2.n107 VDD2.n80 12.0247
R1234 VDD2.n39 VDD2.n12 12.0247
R1235 VDD2.n50 VDD2.n49 12.0247
R1236 VDD2.n120 VDD2.n73 11.249
R1237 VDD2.n104 VDD2.n103 11.249
R1238 VDD2.n36 VDD2.n35 11.249
R1239 VDD2.n53 VDD2.n6 11.249
R1240 VDD2.n121 VDD2.n71 10.4732
R1241 VDD2.n100 VDD2.n82 10.4732
R1242 VDD2.n32 VDD2.n14 10.4732
R1243 VDD2.n54 VDD2.n4 10.4732
R1244 VDD2.n89 VDD2.n88 10.2747
R1245 VDD2.n21 VDD2.n20 10.2747
R1246 VDD2.n125 VDD2.n124 9.69747
R1247 VDD2.n99 VDD2.n84 9.69747
R1248 VDD2.n31 VDD2.n16 9.69747
R1249 VDD2.n58 VDD2.n57 9.69747
R1250 VDD2.n131 VDD2.n130 9.45567
R1251 VDD2.n64 VDD2.n63 9.45567
R1252 VDD2.n91 VDD2.n90 9.3005
R1253 VDD2.n86 VDD2.n85 9.3005
R1254 VDD2.n97 VDD2.n96 9.3005
R1255 VDD2.n99 VDD2.n98 9.3005
R1256 VDD2.n82 VDD2.n81 9.3005
R1257 VDD2.n105 VDD2.n104 9.3005
R1258 VDD2.n107 VDD2.n106 9.3005
R1259 VDD2.n79 VDD2.n76 9.3005
R1260 VDD2.n130 VDD2.n129 9.3005
R1261 VDD2.n69 VDD2.n68 9.3005
R1262 VDD2.n124 VDD2.n123 9.3005
R1263 VDD2.n122 VDD2.n121 9.3005
R1264 VDD2.n73 VDD2.n72 9.3005
R1265 VDD2.n116 VDD2.n115 9.3005
R1266 VDD2.n114 VDD2.n113 9.3005
R1267 VDD2.n63 VDD2.n62 9.3005
R1268 VDD2.n2 VDD2.n1 9.3005
R1269 VDD2.n57 VDD2.n56 9.3005
R1270 VDD2.n55 VDD2.n54 9.3005
R1271 VDD2.n6 VDD2.n5 9.3005
R1272 VDD2.n49 VDD2.n48 9.3005
R1273 VDD2.n47 VDD2.n46 9.3005
R1274 VDD2.n23 VDD2.n22 9.3005
R1275 VDD2.n18 VDD2.n17 9.3005
R1276 VDD2.n29 VDD2.n28 9.3005
R1277 VDD2.n31 VDD2.n30 9.3005
R1278 VDD2.n14 VDD2.n13 9.3005
R1279 VDD2.n37 VDD2.n36 9.3005
R1280 VDD2.n39 VDD2.n38 9.3005
R1281 VDD2.n40 VDD2.n9 9.3005
R1282 VDD2.n128 VDD2.n69 8.92171
R1283 VDD2.n96 VDD2.n95 8.92171
R1284 VDD2.n28 VDD2.n27 8.92171
R1285 VDD2.n61 VDD2.n2 8.92171
R1286 VDD2.n129 VDD2.n67 8.14595
R1287 VDD2.n92 VDD2.n86 8.14595
R1288 VDD2.n24 VDD2.n18 8.14595
R1289 VDD2.n62 VDD2.n0 8.14595
R1290 VDD2.n91 VDD2.n88 7.3702
R1291 VDD2.n23 VDD2.n20 7.3702
R1292 VDD2.n131 VDD2.n67 5.81868
R1293 VDD2.n92 VDD2.n91 5.81868
R1294 VDD2.n24 VDD2.n23 5.81868
R1295 VDD2.n64 VDD2.n0 5.81868
R1296 VDD2.n129 VDD2.n128 5.04292
R1297 VDD2.n95 VDD2.n86 5.04292
R1298 VDD2.n27 VDD2.n18 5.04292
R1299 VDD2.n62 VDD2.n61 5.04292
R1300 VDD2.n125 VDD2.n69 4.26717
R1301 VDD2.n96 VDD2.n84 4.26717
R1302 VDD2.n28 VDD2.n16 4.26717
R1303 VDD2.n58 VDD2.n2 4.26717
R1304 VDD2.n124 VDD2.n71 3.49141
R1305 VDD2.n100 VDD2.n99 3.49141
R1306 VDD2.n32 VDD2.n31 3.49141
R1307 VDD2.n57 VDD2.n4 3.49141
R1308 VDD2.n90 VDD2.n89 2.84303
R1309 VDD2.n22 VDD2.n21 2.84303
R1310 VDD2.n121 VDD2.n120 2.71565
R1311 VDD2.n103 VDD2.n82 2.71565
R1312 VDD2.n35 VDD2.n14 2.71565
R1313 VDD2.n54 VDD2.n53 2.71565
R1314 VDD2.n117 VDD2.n73 1.93989
R1315 VDD2.n104 VDD2.n80 1.93989
R1316 VDD2.n36 VDD2.n12 1.93989
R1317 VDD2.n50 VDD2.n6 1.93989
R1318 VDD2.n133 VDD2.t2 1.63013
R1319 VDD2.n133 VDD2.t3 1.63013
R1320 VDD2.n65 VDD2.t4 1.63013
R1321 VDD2.n65 VDD2.t0 1.63013
R1322 VDD2.n116 VDD2.n75 1.16414
R1323 VDD2.n108 VDD2.n107 1.16414
R1324 VDD2.n41 VDD2.n39 1.16414
R1325 VDD2.n49 VDD2.n8 1.16414
R1326 VDD2 VDD2.n132 0.653517
R1327 VDD2.n113 VDD2.n112 0.388379
R1328 VDD2.n79 VDD2.n77 0.388379
R1329 VDD2.n40 VDD2.n10 0.388379
R1330 VDD2.n46 VDD2.n45 0.388379
R1331 VDD2.n130 VDD2.n68 0.155672
R1332 VDD2.n123 VDD2.n68 0.155672
R1333 VDD2.n123 VDD2.n122 0.155672
R1334 VDD2.n122 VDD2.n72 0.155672
R1335 VDD2.n115 VDD2.n72 0.155672
R1336 VDD2.n115 VDD2.n114 0.155672
R1337 VDD2.n114 VDD2.n76 0.155672
R1338 VDD2.n106 VDD2.n76 0.155672
R1339 VDD2.n106 VDD2.n105 0.155672
R1340 VDD2.n105 VDD2.n81 0.155672
R1341 VDD2.n98 VDD2.n81 0.155672
R1342 VDD2.n98 VDD2.n97 0.155672
R1343 VDD2.n97 VDD2.n85 0.155672
R1344 VDD2.n90 VDD2.n85 0.155672
R1345 VDD2.n22 VDD2.n17 0.155672
R1346 VDD2.n29 VDD2.n17 0.155672
R1347 VDD2.n30 VDD2.n29 0.155672
R1348 VDD2.n30 VDD2.n13 0.155672
R1349 VDD2.n37 VDD2.n13 0.155672
R1350 VDD2.n38 VDD2.n37 0.155672
R1351 VDD2.n38 VDD2.n9 0.155672
R1352 VDD2.n47 VDD2.n9 0.155672
R1353 VDD2.n48 VDD2.n47 0.155672
R1354 VDD2.n48 VDD2.n5 0.155672
R1355 VDD2.n55 VDD2.n5 0.155672
R1356 VDD2.n56 VDD2.n55 0.155672
R1357 VDD2.n56 VDD2.n1 0.155672
R1358 VDD2.n63 VDD2.n1 0.155672
R1359 VTAIL.n266 VTAIL.n206 289.615
R1360 VTAIL.n62 VTAIL.n2 289.615
R1361 VTAIL.n200 VTAIL.n140 289.615
R1362 VTAIL.n132 VTAIL.n72 289.615
R1363 VTAIL.n226 VTAIL.n225 185
R1364 VTAIL.n231 VTAIL.n230 185
R1365 VTAIL.n233 VTAIL.n232 185
R1366 VTAIL.n222 VTAIL.n221 185
R1367 VTAIL.n239 VTAIL.n238 185
R1368 VTAIL.n241 VTAIL.n240 185
R1369 VTAIL.n218 VTAIL.n217 185
R1370 VTAIL.n248 VTAIL.n247 185
R1371 VTAIL.n249 VTAIL.n216 185
R1372 VTAIL.n251 VTAIL.n250 185
R1373 VTAIL.n214 VTAIL.n213 185
R1374 VTAIL.n257 VTAIL.n256 185
R1375 VTAIL.n259 VTAIL.n258 185
R1376 VTAIL.n210 VTAIL.n209 185
R1377 VTAIL.n265 VTAIL.n264 185
R1378 VTAIL.n267 VTAIL.n266 185
R1379 VTAIL.n22 VTAIL.n21 185
R1380 VTAIL.n27 VTAIL.n26 185
R1381 VTAIL.n29 VTAIL.n28 185
R1382 VTAIL.n18 VTAIL.n17 185
R1383 VTAIL.n35 VTAIL.n34 185
R1384 VTAIL.n37 VTAIL.n36 185
R1385 VTAIL.n14 VTAIL.n13 185
R1386 VTAIL.n44 VTAIL.n43 185
R1387 VTAIL.n45 VTAIL.n12 185
R1388 VTAIL.n47 VTAIL.n46 185
R1389 VTAIL.n10 VTAIL.n9 185
R1390 VTAIL.n53 VTAIL.n52 185
R1391 VTAIL.n55 VTAIL.n54 185
R1392 VTAIL.n6 VTAIL.n5 185
R1393 VTAIL.n61 VTAIL.n60 185
R1394 VTAIL.n63 VTAIL.n62 185
R1395 VTAIL.n201 VTAIL.n200 185
R1396 VTAIL.n199 VTAIL.n198 185
R1397 VTAIL.n144 VTAIL.n143 185
R1398 VTAIL.n193 VTAIL.n192 185
R1399 VTAIL.n191 VTAIL.n190 185
R1400 VTAIL.n148 VTAIL.n147 185
R1401 VTAIL.n185 VTAIL.n184 185
R1402 VTAIL.n183 VTAIL.n150 185
R1403 VTAIL.n182 VTAIL.n181 185
R1404 VTAIL.n153 VTAIL.n151 185
R1405 VTAIL.n176 VTAIL.n175 185
R1406 VTAIL.n174 VTAIL.n173 185
R1407 VTAIL.n157 VTAIL.n156 185
R1408 VTAIL.n168 VTAIL.n167 185
R1409 VTAIL.n166 VTAIL.n165 185
R1410 VTAIL.n161 VTAIL.n160 185
R1411 VTAIL.n133 VTAIL.n132 185
R1412 VTAIL.n131 VTAIL.n130 185
R1413 VTAIL.n76 VTAIL.n75 185
R1414 VTAIL.n125 VTAIL.n124 185
R1415 VTAIL.n123 VTAIL.n122 185
R1416 VTAIL.n80 VTAIL.n79 185
R1417 VTAIL.n117 VTAIL.n116 185
R1418 VTAIL.n115 VTAIL.n82 185
R1419 VTAIL.n114 VTAIL.n113 185
R1420 VTAIL.n85 VTAIL.n83 185
R1421 VTAIL.n108 VTAIL.n107 185
R1422 VTAIL.n106 VTAIL.n105 185
R1423 VTAIL.n89 VTAIL.n88 185
R1424 VTAIL.n100 VTAIL.n99 185
R1425 VTAIL.n98 VTAIL.n97 185
R1426 VTAIL.n93 VTAIL.n92 185
R1427 VTAIL.n227 VTAIL.t10 149.524
R1428 VTAIL.n23 VTAIL.t2 149.524
R1429 VTAIL.n162 VTAIL.t3 149.524
R1430 VTAIL.n94 VTAIL.t7 149.524
R1431 VTAIL.n231 VTAIL.n225 104.615
R1432 VTAIL.n232 VTAIL.n231 104.615
R1433 VTAIL.n232 VTAIL.n221 104.615
R1434 VTAIL.n239 VTAIL.n221 104.615
R1435 VTAIL.n240 VTAIL.n239 104.615
R1436 VTAIL.n240 VTAIL.n217 104.615
R1437 VTAIL.n248 VTAIL.n217 104.615
R1438 VTAIL.n249 VTAIL.n248 104.615
R1439 VTAIL.n250 VTAIL.n249 104.615
R1440 VTAIL.n250 VTAIL.n213 104.615
R1441 VTAIL.n257 VTAIL.n213 104.615
R1442 VTAIL.n258 VTAIL.n257 104.615
R1443 VTAIL.n258 VTAIL.n209 104.615
R1444 VTAIL.n265 VTAIL.n209 104.615
R1445 VTAIL.n266 VTAIL.n265 104.615
R1446 VTAIL.n27 VTAIL.n21 104.615
R1447 VTAIL.n28 VTAIL.n27 104.615
R1448 VTAIL.n28 VTAIL.n17 104.615
R1449 VTAIL.n35 VTAIL.n17 104.615
R1450 VTAIL.n36 VTAIL.n35 104.615
R1451 VTAIL.n36 VTAIL.n13 104.615
R1452 VTAIL.n44 VTAIL.n13 104.615
R1453 VTAIL.n45 VTAIL.n44 104.615
R1454 VTAIL.n46 VTAIL.n45 104.615
R1455 VTAIL.n46 VTAIL.n9 104.615
R1456 VTAIL.n53 VTAIL.n9 104.615
R1457 VTAIL.n54 VTAIL.n53 104.615
R1458 VTAIL.n54 VTAIL.n5 104.615
R1459 VTAIL.n61 VTAIL.n5 104.615
R1460 VTAIL.n62 VTAIL.n61 104.615
R1461 VTAIL.n200 VTAIL.n199 104.615
R1462 VTAIL.n199 VTAIL.n143 104.615
R1463 VTAIL.n192 VTAIL.n143 104.615
R1464 VTAIL.n192 VTAIL.n191 104.615
R1465 VTAIL.n191 VTAIL.n147 104.615
R1466 VTAIL.n184 VTAIL.n147 104.615
R1467 VTAIL.n184 VTAIL.n183 104.615
R1468 VTAIL.n183 VTAIL.n182 104.615
R1469 VTAIL.n182 VTAIL.n151 104.615
R1470 VTAIL.n175 VTAIL.n151 104.615
R1471 VTAIL.n175 VTAIL.n174 104.615
R1472 VTAIL.n174 VTAIL.n156 104.615
R1473 VTAIL.n167 VTAIL.n156 104.615
R1474 VTAIL.n167 VTAIL.n166 104.615
R1475 VTAIL.n166 VTAIL.n160 104.615
R1476 VTAIL.n132 VTAIL.n131 104.615
R1477 VTAIL.n131 VTAIL.n75 104.615
R1478 VTAIL.n124 VTAIL.n75 104.615
R1479 VTAIL.n124 VTAIL.n123 104.615
R1480 VTAIL.n123 VTAIL.n79 104.615
R1481 VTAIL.n116 VTAIL.n79 104.615
R1482 VTAIL.n116 VTAIL.n115 104.615
R1483 VTAIL.n115 VTAIL.n114 104.615
R1484 VTAIL.n114 VTAIL.n83 104.615
R1485 VTAIL.n107 VTAIL.n83 104.615
R1486 VTAIL.n107 VTAIL.n106 104.615
R1487 VTAIL.n106 VTAIL.n88 104.615
R1488 VTAIL.n99 VTAIL.n88 104.615
R1489 VTAIL.n99 VTAIL.n98 104.615
R1490 VTAIL.n98 VTAIL.n92 104.615
R1491 VTAIL.t10 VTAIL.n225 52.3082
R1492 VTAIL.t2 VTAIL.n21 52.3082
R1493 VTAIL.t3 VTAIL.n160 52.3082
R1494 VTAIL.t7 VTAIL.n92 52.3082
R1495 VTAIL.n139 VTAIL.n138 45.783
R1496 VTAIL.n71 VTAIL.n70 45.783
R1497 VTAIL.n1 VTAIL.n0 45.7828
R1498 VTAIL.n69 VTAIL.n68 45.7828
R1499 VTAIL.n271 VTAIL.n270 32.7672
R1500 VTAIL.n67 VTAIL.n66 32.7672
R1501 VTAIL.n205 VTAIL.n204 32.7672
R1502 VTAIL.n137 VTAIL.n136 32.7672
R1503 VTAIL.n71 VTAIL.n69 24.4272
R1504 VTAIL.n271 VTAIL.n205 23.6341
R1505 VTAIL.n251 VTAIL.n216 13.1884
R1506 VTAIL.n47 VTAIL.n12 13.1884
R1507 VTAIL.n185 VTAIL.n150 13.1884
R1508 VTAIL.n117 VTAIL.n82 13.1884
R1509 VTAIL.n247 VTAIL.n246 12.8005
R1510 VTAIL.n252 VTAIL.n214 12.8005
R1511 VTAIL.n43 VTAIL.n42 12.8005
R1512 VTAIL.n48 VTAIL.n10 12.8005
R1513 VTAIL.n186 VTAIL.n148 12.8005
R1514 VTAIL.n181 VTAIL.n152 12.8005
R1515 VTAIL.n118 VTAIL.n80 12.8005
R1516 VTAIL.n113 VTAIL.n84 12.8005
R1517 VTAIL.n245 VTAIL.n218 12.0247
R1518 VTAIL.n256 VTAIL.n255 12.0247
R1519 VTAIL.n41 VTAIL.n14 12.0247
R1520 VTAIL.n52 VTAIL.n51 12.0247
R1521 VTAIL.n190 VTAIL.n189 12.0247
R1522 VTAIL.n180 VTAIL.n153 12.0247
R1523 VTAIL.n122 VTAIL.n121 12.0247
R1524 VTAIL.n112 VTAIL.n85 12.0247
R1525 VTAIL.n242 VTAIL.n241 11.249
R1526 VTAIL.n259 VTAIL.n212 11.249
R1527 VTAIL.n38 VTAIL.n37 11.249
R1528 VTAIL.n55 VTAIL.n8 11.249
R1529 VTAIL.n193 VTAIL.n146 11.249
R1530 VTAIL.n177 VTAIL.n176 11.249
R1531 VTAIL.n125 VTAIL.n78 11.249
R1532 VTAIL.n109 VTAIL.n108 11.249
R1533 VTAIL.n238 VTAIL.n220 10.4732
R1534 VTAIL.n260 VTAIL.n210 10.4732
R1535 VTAIL.n34 VTAIL.n16 10.4732
R1536 VTAIL.n56 VTAIL.n6 10.4732
R1537 VTAIL.n194 VTAIL.n144 10.4732
R1538 VTAIL.n173 VTAIL.n155 10.4732
R1539 VTAIL.n126 VTAIL.n76 10.4732
R1540 VTAIL.n105 VTAIL.n87 10.4732
R1541 VTAIL.n227 VTAIL.n226 10.2747
R1542 VTAIL.n23 VTAIL.n22 10.2747
R1543 VTAIL.n162 VTAIL.n161 10.2747
R1544 VTAIL.n94 VTAIL.n93 10.2747
R1545 VTAIL.n237 VTAIL.n222 9.69747
R1546 VTAIL.n264 VTAIL.n263 9.69747
R1547 VTAIL.n33 VTAIL.n18 9.69747
R1548 VTAIL.n60 VTAIL.n59 9.69747
R1549 VTAIL.n198 VTAIL.n197 9.69747
R1550 VTAIL.n172 VTAIL.n157 9.69747
R1551 VTAIL.n130 VTAIL.n129 9.69747
R1552 VTAIL.n104 VTAIL.n89 9.69747
R1553 VTAIL.n270 VTAIL.n269 9.45567
R1554 VTAIL.n66 VTAIL.n65 9.45567
R1555 VTAIL.n204 VTAIL.n203 9.45567
R1556 VTAIL.n136 VTAIL.n135 9.45567
R1557 VTAIL.n269 VTAIL.n268 9.3005
R1558 VTAIL.n208 VTAIL.n207 9.3005
R1559 VTAIL.n263 VTAIL.n262 9.3005
R1560 VTAIL.n261 VTAIL.n260 9.3005
R1561 VTAIL.n212 VTAIL.n211 9.3005
R1562 VTAIL.n255 VTAIL.n254 9.3005
R1563 VTAIL.n253 VTAIL.n252 9.3005
R1564 VTAIL.n229 VTAIL.n228 9.3005
R1565 VTAIL.n224 VTAIL.n223 9.3005
R1566 VTAIL.n235 VTAIL.n234 9.3005
R1567 VTAIL.n237 VTAIL.n236 9.3005
R1568 VTAIL.n220 VTAIL.n219 9.3005
R1569 VTAIL.n243 VTAIL.n242 9.3005
R1570 VTAIL.n245 VTAIL.n244 9.3005
R1571 VTAIL.n246 VTAIL.n215 9.3005
R1572 VTAIL.n65 VTAIL.n64 9.3005
R1573 VTAIL.n4 VTAIL.n3 9.3005
R1574 VTAIL.n59 VTAIL.n58 9.3005
R1575 VTAIL.n57 VTAIL.n56 9.3005
R1576 VTAIL.n8 VTAIL.n7 9.3005
R1577 VTAIL.n51 VTAIL.n50 9.3005
R1578 VTAIL.n49 VTAIL.n48 9.3005
R1579 VTAIL.n25 VTAIL.n24 9.3005
R1580 VTAIL.n20 VTAIL.n19 9.3005
R1581 VTAIL.n31 VTAIL.n30 9.3005
R1582 VTAIL.n33 VTAIL.n32 9.3005
R1583 VTAIL.n16 VTAIL.n15 9.3005
R1584 VTAIL.n39 VTAIL.n38 9.3005
R1585 VTAIL.n41 VTAIL.n40 9.3005
R1586 VTAIL.n42 VTAIL.n11 9.3005
R1587 VTAIL.n164 VTAIL.n163 9.3005
R1588 VTAIL.n159 VTAIL.n158 9.3005
R1589 VTAIL.n170 VTAIL.n169 9.3005
R1590 VTAIL.n172 VTAIL.n171 9.3005
R1591 VTAIL.n155 VTAIL.n154 9.3005
R1592 VTAIL.n178 VTAIL.n177 9.3005
R1593 VTAIL.n180 VTAIL.n179 9.3005
R1594 VTAIL.n152 VTAIL.n149 9.3005
R1595 VTAIL.n203 VTAIL.n202 9.3005
R1596 VTAIL.n142 VTAIL.n141 9.3005
R1597 VTAIL.n197 VTAIL.n196 9.3005
R1598 VTAIL.n195 VTAIL.n194 9.3005
R1599 VTAIL.n146 VTAIL.n145 9.3005
R1600 VTAIL.n189 VTAIL.n188 9.3005
R1601 VTAIL.n187 VTAIL.n186 9.3005
R1602 VTAIL.n96 VTAIL.n95 9.3005
R1603 VTAIL.n91 VTAIL.n90 9.3005
R1604 VTAIL.n102 VTAIL.n101 9.3005
R1605 VTAIL.n104 VTAIL.n103 9.3005
R1606 VTAIL.n87 VTAIL.n86 9.3005
R1607 VTAIL.n110 VTAIL.n109 9.3005
R1608 VTAIL.n112 VTAIL.n111 9.3005
R1609 VTAIL.n84 VTAIL.n81 9.3005
R1610 VTAIL.n135 VTAIL.n134 9.3005
R1611 VTAIL.n74 VTAIL.n73 9.3005
R1612 VTAIL.n129 VTAIL.n128 9.3005
R1613 VTAIL.n127 VTAIL.n126 9.3005
R1614 VTAIL.n78 VTAIL.n77 9.3005
R1615 VTAIL.n121 VTAIL.n120 9.3005
R1616 VTAIL.n119 VTAIL.n118 9.3005
R1617 VTAIL.n234 VTAIL.n233 8.92171
R1618 VTAIL.n267 VTAIL.n208 8.92171
R1619 VTAIL.n30 VTAIL.n29 8.92171
R1620 VTAIL.n63 VTAIL.n4 8.92171
R1621 VTAIL.n201 VTAIL.n142 8.92171
R1622 VTAIL.n169 VTAIL.n168 8.92171
R1623 VTAIL.n133 VTAIL.n74 8.92171
R1624 VTAIL.n101 VTAIL.n100 8.92171
R1625 VTAIL.n230 VTAIL.n224 8.14595
R1626 VTAIL.n268 VTAIL.n206 8.14595
R1627 VTAIL.n26 VTAIL.n20 8.14595
R1628 VTAIL.n64 VTAIL.n2 8.14595
R1629 VTAIL.n202 VTAIL.n140 8.14595
R1630 VTAIL.n165 VTAIL.n159 8.14595
R1631 VTAIL.n134 VTAIL.n72 8.14595
R1632 VTAIL.n97 VTAIL.n91 8.14595
R1633 VTAIL.n229 VTAIL.n226 7.3702
R1634 VTAIL.n25 VTAIL.n22 7.3702
R1635 VTAIL.n164 VTAIL.n161 7.3702
R1636 VTAIL.n96 VTAIL.n93 7.3702
R1637 VTAIL.n230 VTAIL.n229 5.81868
R1638 VTAIL.n270 VTAIL.n206 5.81868
R1639 VTAIL.n26 VTAIL.n25 5.81868
R1640 VTAIL.n66 VTAIL.n2 5.81868
R1641 VTAIL.n204 VTAIL.n140 5.81868
R1642 VTAIL.n165 VTAIL.n164 5.81868
R1643 VTAIL.n136 VTAIL.n72 5.81868
R1644 VTAIL.n97 VTAIL.n96 5.81868
R1645 VTAIL.n233 VTAIL.n224 5.04292
R1646 VTAIL.n268 VTAIL.n267 5.04292
R1647 VTAIL.n29 VTAIL.n20 5.04292
R1648 VTAIL.n64 VTAIL.n63 5.04292
R1649 VTAIL.n202 VTAIL.n201 5.04292
R1650 VTAIL.n168 VTAIL.n159 5.04292
R1651 VTAIL.n134 VTAIL.n133 5.04292
R1652 VTAIL.n100 VTAIL.n91 5.04292
R1653 VTAIL.n234 VTAIL.n222 4.26717
R1654 VTAIL.n264 VTAIL.n208 4.26717
R1655 VTAIL.n30 VTAIL.n18 4.26717
R1656 VTAIL.n60 VTAIL.n4 4.26717
R1657 VTAIL.n198 VTAIL.n142 4.26717
R1658 VTAIL.n169 VTAIL.n157 4.26717
R1659 VTAIL.n130 VTAIL.n74 4.26717
R1660 VTAIL.n101 VTAIL.n89 4.26717
R1661 VTAIL.n238 VTAIL.n237 3.49141
R1662 VTAIL.n263 VTAIL.n210 3.49141
R1663 VTAIL.n34 VTAIL.n33 3.49141
R1664 VTAIL.n59 VTAIL.n6 3.49141
R1665 VTAIL.n197 VTAIL.n144 3.49141
R1666 VTAIL.n173 VTAIL.n172 3.49141
R1667 VTAIL.n129 VTAIL.n76 3.49141
R1668 VTAIL.n105 VTAIL.n104 3.49141
R1669 VTAIL.n228 VTAIL.n227 2.84303
R1670 VTAIL.n24 VTAIL.n23 2.84303
R1671 VTAIL.n163 VTAIL.n162 2.84303
R1672 VTAIL.n95 VTAIL.n94 2.84303
R1673 VTAIL.n241 VTAIL.n220 2.71565
R1674 VTAIL.n260 VTAIL.n259 2.71565
R1675 VTAIL.n37 VTAIL.n16 2.71565
R1676 VTAIL.n56 VTAIL.n55 2.71565
R1677 VTAIL.n194 VTAIL.n193 2.71565
R1678 VTAIL.n176 VTAIL.n155 2.71565
R1679 VTAIL.n126 VTAIL.n125 2.71565
R1680 VTAIL.n108 VTAIL.n87 2.71565
R1681 VTAIL.n242 VTAIL.n218 1.93989
R1682 VTAIL.n256 VTAIL.n212 1.93989
R1683 VTAIL.n38 VTAIL.n14 1.93989
R1684 VTAIL.n52 VTAIL.n8 1.93989
R1685 VTAIL.n190 VTAIL.n146 1.93989
R1686 VTAIL.n177 VTAIL.n153 1.93989
R1687 VTAIL.n122 VTAIL.n78 1.93989
R1688 VTAIL.n109 VTAIL.n85 1.93989
R1689 VTAIL.n0 VTAIL.t8 1.63013
R1690 VTAIL.n0 VTAIL.t11 1.63013
R1691 VTAIL.n68 VTAIL.t4 1.63013
R1692 VTAIL.n68 VTAIL.t1 1.63013
R1693 VTAIL.n138 VTAIL.t5 1.63013
R1694 VTAIL.n138 VTAIL.t0 1.63013
R1695 VTAIL.n70 VTAIL.t6 1.63013
R1696 VTAIL.n70 VTAIL.t9 1.63013
R1697 VTAIL.n247 VTAIL.n245 1.16414
R1698 VTAIL.n255 VTAIL.n214 1.16414
R1699 VTAIL.n43 VTAIL.n41 1.16414
R1700 VTAIL.n51 VTAIL.n10 1.16414
R1701 VTAIL.n189 VTAIL.n148 1.16414
R1702 VTAIL.n181 VTAIL.n180 1.16414
R1703 VTAIL.n121 VTAIL.n80 1.16414
R1704 VTAIL.n113 VTAIL.n112 1.16414
R1705 VTAIL.n139 VTAIL.n137 0.866879
R1706 VTAIL.n67 VTAIL.n1 0.866879
R1707 VTAIL.n137 VTAIL.n71 0.793603
R1708 VTAIL.n205 VTAIL.n139 0.793603
R1709 VTAIL.n69 VTAIL.n67 0.793603
R1710 VTAIL VTAIL.n271 0.537138
R1711 VTAIL.n246 VTAIL.n216 0.388379
R1712 VTAIL.n252 VTAIL.n251 0.388379
R1713 VTAIL.n42 VTAIL.n12 0.388379
R1714 VTAIL.n48 VTAIL.n47 0.388379
R1715 VTAIL.n186 VTAIL.n185 0.388379
R1716 VTAIL.n152 VTAIL.n150 0.388379
R1717 VTAIL.n118 VTAIL.n117 0.388379
R1718 VTAIL.n84 VTAIL.n82 0.388379
R1719 VTAIL VTAIL.n1 0.256966
R1720 VTAIL.n228 VTAIL.n223 0.155672
R1721 VTAIL.n235 VTAIL.n223 0.155672
R1722 VTAIL.n236 VTAIL.n235 0.155672
R1723 VTAIL.n236 VTAIL.n219 0.155672
R1724 VTAIL.n243 VTAIL.n219 0.155672
R1725 VTAIL.n244 VTAIL.n243 0.155672
R1726 VTAIL.n244 VTAIL.n215 0.155672
R1727 VTAIL.n253 VTAIL.n215 0.155672
R1728 VTAIL.n254 VTAIL.n253 0.155672
R1729 VTAIL.n254 VTAIL.n211 0.155672
R1730 VTAIL.n261 VTAIL.n211 0.155672
R1731 VTAIL.n262 VTAIL.n261 0.155672
R1732 VTAIL.n262 VTAIL.n207 0.155672
R1733 VTAIL.n269 VTAIL.n207 0.155672
R1734 VTAIL.n24 VTAIL.n19 0.155672
R1735 VTAIL.n31 VTAIL.n19 0.155672
R1736 VTAIL.n32 VTAIL.n31 0.155672
R1737 VTAIL.n32 VTAIL.n15 0.155672
R1738 VTAIL.n39 VTAIL.n15 0.155672
R1739 VTAIL.n40 VTAIL.n39 0.155672
R1740 VTAIL.n40 VTAIL.n11 0.155672
R1741 VTAIL.n49 VTAIL.n11 0.155672
R1742 VTAIL.n50 VTAIL.n49 0.155672
R1743 VTAIL.n50 VTAIL.n7 0.155672
R1744 VTAIL.n57 VTAIL.n7 0.155672
R1745 VTAIL.n58 VTAIL.n57 0.155672
R1746 VTAIL.n58 VTAIL.n3 0.155672
R1747 VTAIL.n65 VTAIL.n3 0.155672
R1748 VTAIL.n203 VTAIL.n141 0.155672
R1749 VTAIL.n196 VTAIL.n141 0.155672
R1750 VTAIL.n196 VTAIL.n195 0.155672
R1751 VTAIL.n195 VTAIL.n145 0.155672
R1752 VTAIL.n188 VTAIL.n145 0.155672
R1753 VTAIL.n188 VTAIL.n187 0.155672
R1754 VTAIL.n187 VTAIL.n149 0.155672
R1755 VTAIL.n179 VTAIL.n149 0.155672
R1756 VTAIL.n179 VTAIL.n178 0.155672
R1757 VTAIL.n178 VTAIL.n154 0.155672
R1758 VTAIL.n171 VTAIL.n154 0.155672
R1759 VTAIL.n171 VTAIL.n170 0.155672
R1760 VTAIL.n170 VTAIL.n158 0.155672
R1761 VTAIL.n163 VTAIL.n158 0.155672
R1762 VTAIL.n135 VTAIL.n73 0.155672
R1763 VTAIL.n128 VTAIL.n73 0.155672
R1764 VTAIL.n128 VTAIL.n127 0.155672
R1765 VTAIL.n127 VTAIL.n77 0.155672
R1766 VTAIL.n120 VTAIL.n77 0.155672
R1767 VTAIL.n120 VTAIL.n119 0.155672
R1768 VTAIL.n119 VTAIL.n81 0.155672
R1769 VTAIL.n111 VTAIL.n81 0.155672
R1770 VTAIL.n111 VTAIL.n110 0.155672
R1771 VTAIL.n110 VTAIL.n86 0.155672
R1772 VTAIL.n103 VTAIL.n86 0.155672
R1773 VTAIL.n103 VTAIL.n102 0.155672
R1774 VTAIL.n102 VTAIL.n90 0.155672
R1775 VTAIL.n95 VTAIL.n90 0.155672
R1776 VP.n1 VP.t0 590.109
R1777 VP.n6 VP.t2 563.287
R1778 VP.n7 VP.t4 563.287
R1779 VP.n8 VP.t3 563.287
R1780 VP.n3 VP.t1 563.287
R1781 VP.n2 VP.t5 563.287
R1782 VP.n9 VP.n8 161.3
R1783 VP.n4 VP.n3 161.3
R1784 VP.n6 VP.n5 161.3
R1785 VP.n7 VP.n0 80.6037
R1786 VP.n7 VP.n6 48.2005
R1787 VP.n8 VP.n7 48.2005
R1788 VP.n3 VP.n2 48.2005
R1789 VP.n4 VP.n1 45.1367
R1790 VP.n5 VP.n4 40.9626
R1791 VP.n2 VP.n1 13.3799
R1792 VP.n5 VP.n0 0.285035
R1793 VP.n9 VP.n0 0.285035
R1794 VP VP.n9 0.0516364
R1795 VDD1.n60 VDD1.n0 289.615
R1796 VDD1.n125 VDD1.n65 289.615
R1797 VDD1.n61 VDD1.n60 185
R1798 VDD1.n59 VDD1.n58 185
R1799 VDD1.n4 VDD1.n3 185
R1800 VDD1.n53 VDD1.n52 185
R1801 VDD1.n51 VDD1.n50 185
R1802 VDD1.n8 VDD1.n7 185
R1803 VDD1.n45 VDD1.n44 185
R1804 VDD1.n43 VDD1.n10 185
R1805 VDD1.n42 VDD1.n41 185
R1806 VDD1.n13 VDD1.n11 185
R1807 VDD1.n36 VDD1.n35 185
R1808 VDD1.n34 VDD1.n33 185
R1809 VDD1.n17 VDD1.n16 185
R1810 VDD1.n28 VDD1.n27 185
R1811 VDD1.n26 VDD1.n25 185
R1812 VDD1.n21 VDD1.n20 185
R1813 VDD1.n85 VDD1.n84 185
R1814 VDD1.n90 VDD1.n89 185
R1815 VDD1.n92 VDD1.n91 185
R1816 VDD1.n81 VDD1.n80 185
R1817 VDD1.n98 VDD1.n97 185
R1818 VDD1.n100 VDD1.n99 185
R1819 VDD1.n77 VDD1.n76 185
R1820 VDD1.n107 VDD1.n106 185
R1821 VDD1.n108 VDD1.n75 185
R1822 VDD1.n110 VDD1.n109 185
R1823 VDD1.n73 VDD1.n72 185
R1824 VDD1.n116 VDD1.n115 185
R1825 VDD1.n118 VDD1.n117 185
R1826 VDD1.n69 VDD1.n68 185
R1827 VDD1.n124 VDD1.n123 185
R1828 VDD1.n126 VDD1.n125 185
R1829 VDD1.n22 VDD1.t5 149.524
R1830 VDD1.n86 VDD1.t3 149.524
R1831 VDD1.n60 VDD1.n59 104.615
R1832 VDD1.n59 VDD1.n3 104.615
R1833 VDD1.n52 VDD1.n3 104.615
R1834 VDD1.n52 VDD1.n51 104.615
R1835 VDD1.n51 VDD1.n7 104.615
R1836 VDD1.n44 VDD1.n7 104.615
R1837 VDD1.n44 VDD1.n43 104.615
R1838 VDD1.n43 VDD1.n42 104.615
R1839 VDD1.n42 VDD1.n11 104.615
R1840 VDD1.n35 VDD1.n11 104.615
R1841 VDD1.n35 VDD1.n34 104.615
R1842 VDD1.n34 VDD1.n16 104.615
R1843 VDD1.n27 VDD1.n16 104.615
R1844 VDD1.n27 VDD1.n26 104.615
R1845 VDD1.n26 VDD1.n20 104.615
R1846 VDD1.n90 VDD1.n84 104.615
R1847 VDD1.n91 VDD1.n90 104.615
R1848 VDD1.n91 VDD1.n80 104.615
R1849 VDD1.n98 VDD1.n80 104.615
R1850 VDD1.n99 VDD1.n98 104.615
R1851 VDD1.n99 VDD1.n76 104.615
R1852 VDD1.n107 VDD1.n76 104.615
R1853 VDD1.n108 VDD1.n107 104.615
R1854 VDD1.n109 VDD1.n108 104.615
R1855 VDD1.n109 VDD1.n72 104.615
R1856 VDD1.n116 VDD1.n72 104.615
R1857 VDD1.n117 VDD1.n116 104.615
R1858 VDD1.n117 VDD1.n68 104.615
R1859 VDD1.n124 VDD1.n68 104.615
R1860 VDD1.n125 VDD1.n124 104.615
R1861 VDD1.n131 VDD1.n130 62.6045
R1862 VDD1.n133 VDD1.n132 62.4616
R1863 VDD1.t5 VDD1.n20 52.3082
R1864 VDD1.t3 VDD1.n84 52.3082
R1865 VDD1 VDD1.n64 50.099
R1866 VDD1.n131 VDD1.n129 49.9854
R1867 VDD1.n133 VDD1.n131 37.7466
R1868 VDD1.n45 VDD1.n10 13.1884
R1869 VDD1.n110 VDD1.n75 13.1884
R1870 VDD1.n46 VDD1.n8 12.8005
R1871 VDD1.n41 VDD1.n12 12.8005
R1872 VDD1.n106 VDD1.n105 12.8005
R1873 VDD1.n111 VDD1.n73 12.8005
R1874 VDD1.n50 VDD1.n49 12.0247
R1875 VDD1.n40 VDD1.n13 12.0247
R1876 VDD1.n104 VDD1.n77 12.0247
R1877 VDD1.n115 VDD1.n114 12.0247
R1878 VDD1.n53 VDD1.n6 11.249
R1879 VDD1.n37 VDD1.n36 11.249
R1880 VDD1.n101 VDD1.n100 11.249
R1881 VDD1.n118 VDD1.n71 11.249
R1882 VDD1.n54 VDD1.n4 10.4732
R1883 VDD1.n33 VDD1.n15 10.4732
R1884 VDD1.n97 VDD1.n79 10.4732
R1885 VDD1.n119 VDD1.n69 10.4732
R1886 VDD1.n22 VDD1.n21 10.2747
R1887 VDD1.n86 VDD1.n85 10.2747
R1888 VDD1.n58 VDD1.n57 9.69747
R1889 VDD1.n32 VDD1.n17 9.69747
R1890 VDD1.n96 VDD1.n81 9.69747
R1891 VDD1.n123 VDD1.n122 9.69747
R1892 VDD1.n64 VDD1.n63 9.45567
R1893 VDD1.n129 VDD1.n128 9.45567
R1894 VDD1.n24 VDD1.n23 9.3005
R1895 VDD1.n19 VDD1.n18 9.3005
R1896 VDD1.n30 VDD1.n29 9.3005
R1897 VDD1.n32 VDD1.n31 9.3005
R1898 VDD1.n15 VDD1.n14 9.3005
R1899 VDD1.n38 VDD1.n37 9.3005
R1900 VDD1.n40 VDD1.n39 9.3005
R1901 VDD1.n12 VDD1.n9 9.3005
R1902 VDD1.n63 VDD1.n62 9.3005
R1903 VDD1.n2 VDD1.n1 9.3005
R1904 VDD1.n57 VDD1.n56 9.3005
R1905 VDD1.n55 VDD1.n54 9.3005
R1906 VDD1.n6 VDD1.n5 9.3005
R1907 VDD1.n49 VDD1.n48 9.3005
R1908 VDD1.n47 VDD1.n46 9.3005
R1909 VDD1.n128 VDD1.n127 9.3005
R1910 VDD1.n67 VDD1.n66 9.3005
R1911 VDD1.n122 VDD1.n121 9.3005
R1912 VDD1.n120 VDD1.n119 9.3005
R1913 VDD1.n71 VDD1.n70 9.3005
R1914 VDD1.n114 VDD1.n113 9.3005
R1915 VDD1.n112 VDD1.n111 9.3005
R1916 VDD1.n88 VDD1.n87 9.3005
R1917 VDD1.n83 VDD1.n82 9.3005
R1918 VDD1.n94 VDD1.n93 9.3005
R1919 VDD1.n96 VDD1.n95 9.3005
R1920 VDD1.n79 VDD1.n78 9.3005
R1921 VDD1.n102 VDD1.n101 9.3005
R1922 VDD1.n104 VDD1.n103 9.3005
R1923 VDD1.n105 VDD1.n74 9.3005
R1924 VDD1.n61 VDD1.n2 8.92171
R1925 VDD1.n29 VDD1.n28 8.92171
R1926 VDD1.n93 VDD1.n92 8.92171
R1927 VDD1.n126 VDD1.n67 8.92171
R1928 VDD1.n62 VDD1.n0 8.14595
R1929 VDD1.n25 VDD1.n19 8.14595
R1930 VDD1.n89 VDD1.n83 8.14595
R1931 VDD1.n127 VDD1.n65 8.14595
R1932 VDD1.n24 VDD1.n21 7.3702
R1933 VDD1.n88 VDD1.n85 7.3702
R1934 VDD1.n64 VDD1.n0 5.81868
R1935 VDD1.n25 VDD1.n24 5.81868
R1936 VDD1.n89 VDD1.n88 5.81868
R1937 VDD1.n129 VDD1.n65 5.81868
R1938 VDD1.n62 VDD1.n61 5.04292
R1939 VDD1.n28 VDD1.n19 5.04292
R1940 VDD1.n92 VDD1.n83 5.04292
R1941 VDD1.n127 VDD1.n126 5.04292
R1942 VDD1.n58 VDD1.n2 4.26717
R1943 VDD1.n29 VDD1.n17 4.26717
R1944 VDD1.n93 VDD1.n81 4.26717
R1945 VDD1.n123 VDD1.n67 4.26717
R1946 VDD1.n57 VDD1.n4 3.49141
R1947 VDD1.n33 VDD1.n32 3.49141
R1948 VDD1.n97 VDD1.n96 3.49141
R1949 VDD1.n122 VDD1.n69 3.49141
R1950 VDD1.n23 VDD1.n22 2.84303
R1951 VDD1.n87 VDD1.n86 2.84303
R1952 VDD1.n54 VDD1.n53 2.71565
R1953 VDD1.n36 VDD1.n15 2.71565
R1954 VDD1.n100 VDD1.n79 2.71565
R1955 VDD1.n119 VDD1.n118 2.71565
R1956 VDD1.n50 VDD1.n6 1.93989
R1957 VDD1.n37 VDD1.n13 1.93989
R1958 VDD1.n101 VDD1.n77 1.93989
R1959 VDD1.n115 VDD1.n71 1.93989
R1960 VDD1.n132 VDD1.t0 1.63013
R1961 VDD1.n132 VDD1.t4 1.63013
R1962 VDD1.n130 VDD1.t1 1.63013
R1963 VDD1.n130 VDD1.t2 1.63013
R1964 VDD1.n49 VDD1.n8 1.16414
R1965 VDD1.n41 VDD1.n40 1.16414
R1966 VDD1.n106 VDD1.n104 1.16414
R1967 VDD1.n114 VDD1.n73 1.16414
R1968 VDD1.n46 VDD1.n45 0.388379
R1969 VDD1.n12 VDD1.n10 0.388379
R1970 VDD1.n105 VDD1.n75 0.388379
R1971 VDD1.n111 VDD1.n110 0.388379
R1972 VDD1.n63 VDD1.n1 0.155672
R1973 VDD1.n56 VDD1.n1 0.155672
R1974 VDD1.n56 VDD1.n55 0.155672
R1975 VDD1.n55 VDD1.n5 0.155672
R1976 VDD1.n48 VDD1.n5 0.155672
R1977 VDD1.n48 VDD1.n47 0.155672
R1978 VDD1.n47 VDD1.n9 0.155672
R1979 VDD1.n39 VDD1.n9 0.155672
R1980 VDD1.n39 VDD1.n38 0.155672
R1981 VDD1.n38 VDD1.n14 0.155672
R1982 VDD1.n31 VDD1.n14 0.155672
R1983 VDD1.n31 VDD1.n30 0.155672
R1984 VDD1.n30 VDD1.n18 0.155672
R1985 VDD1.n23 VDD1.n18 0.155672
R1986 VDD1.n87 VDD1.n82 0.155672
R1987 VDD1.n94 VDD1.n82 0.155672
R1988 VDD1.n95 VDD1.n94 0.155672
R1989 VDD1.n95 VDD1.n78 0.155672
R1990 VDD1.n102 VDD1.n78 0.155672
R1991 VDD1.n103 VDD1.n102 0.155672
R1992 VDD1.n103 VDD1.n74 0.155672
R1993 VDD1.n112 VDD1.n74 0.155672
R1994 VDD1.n113 VDD1.n112 0.155672
R1995 VDD1.n113 VDD1.n70 0.155672
R1996 VDD1.n120 VDD1.n70 0.155672
R1997 VDD1.n121 VDD1.n120 0.155672
R1998 VDD1.n121 VDD1.n66 0.155672
R1999 VDD1.n128 VDD1.n66 0.155672
R2000 VDD1 VDD1.n133 0.140586
C0 VTAIL VN 3.66596f
C1 VP VN 5.00003f
C2 VDD1 VDD2 0.671878f
C3 VTAIL VP 3.68061f
C4 VDD2 VN 4.01913f
C5 VTAIL VDD2 10.7459f
C6 VDD1 VN 0.148047f
C7 VP VDD2 0.288436f
C8 VTAIL VDD1 10.713099f
C9 VP VDD1 4.154779f
C10 VDD2 B 4.437539f
C11 VDD1 B 4.446931f
C12 VTAIL B 6.344298f
C13 VN B 7.49455f
C14 VP B 5.43858f
C15 VDD1.n0 B 0.034354f
C16 VDD1.n1 B 0.024094f
C17 VDD1.n2 B 0.012947f
C18 VDD1.n3 B 0.030603f
C19 VDD1.n4 B 0.013709f
C20 VDD1.n5 B 0.024094f
C21 VDD1.n6 B 0.012947f
C22 VDD1.n7 B 0.030603f
C23 VDD1.n8 B 0.013709f
C24 VDD1.n9 B 0.024094f
C25 VDD1.n10 B 0.013328f
C26 VDD1.n11 B 0.030603f
C27 VDD1.n12 B 0.012947f
C28 VDD1.n13 B 0.013709f
C29 VDD1.n14 B 0.024094f
C30 VDD1.n15 B 0.012947f
C31 VDD1.n16 B 0.030603f
C32 VDD1.n17 B 0.013709f
C33 VDD1.n18 B 0.024094f
C34 VDD1.n19 B 0.012947f
C35 VDD1.n20 B 0.022952f
C36 VDD1.n21 B 0.021634f
C37 VDD1.t5 B 0.051705f
C38 VDD1.n22 B 0.175105f
C39 VDD1.n23 B 1.23159f
C40 VDD1.n24 B 0.012947f
C41 VDD1.n25 B 0.013709f
C42 VDD1.n26 B 0.030603f
C43 VDD1.n27 B 0.030603f
C44 VDD1.n28 B 0.013709f
C45 VDD1.n29 B 0.012947f
C46 VDD1.n30 B 0.024094f
C47 VDD1.n31 B 0.024094f
C48 VDD1.n32 B 0.012947f
C49 VDD1.n33 B 0.013709f
C50 VDD1.n34 B 0.030603f
C51 VDD1.n35 B 0.030603f
C52 VDD1.n36 B 0.013709f
C53 VDD1.n37 B 0.012947f
C54 VDD1.n38 B 0.024094f
C55 VDD1.n39 B 0.024094f
C56 VDD1.n40 B 0.012947f
C57 VDD1.n41 B 0.013709f
C58 VDD1.n42 B 0.030603f
C59 VDD1.n43 B 0.030603f
C60 VDD1.n44 B 0.030603f
C61 VDD1.n45 B 0.013328f
C62 VDD1.n46 B 0.012947f
C63 VDD1.n47 B 0.024094f
C64 VDD1.n48 B 0.024094f
C65 VDD1.n49 B 0.012947f
C66 VDD1.n50 B 0.013709f
C67 VDD1.n51 B 0.030603f
C68 VDD1.n52 B 0.030603f
C69 VDD1.n53 B 0.013709f
C70 VDD1.n54 B 0.012947f
C71 VDD1.n55 B 0.024094f
C72 VDD1.n56 B 0.024094f
C73 VDD1.n57 B 0.012947f
C74 VDD1.n58 B 0.013709f
C75 VDD1.n59 B 0.030603f
C76 VDD1.n60 B 0.067112f
C77 VDD1.n61 B 0.013709f
C78 VDD1.n62 B 0.012947f
C79 VDD1.n63 B 0.05668f
C80 VDD1.n64 B 0.055572f
C81 VDD1.n65 B 0.034354f
C82 VDD1.n66 B 0.024094f
C83 VDD1.n67 B 0.012947f
C84 VDD1.n68 B 0.030603f
C85 VDD1.n69 B 0.013709f
C86 VDD1.n70 B 0.024094f
C87 VDD1.n71 B 0.012947f
C88 VDD1.n72 B 0.030603f
C89 VDD1.n73 B 0.013709f
C90 VDD1.n74 B 0.024094f
C91 VDD1.n75 B 0.013328f
C92 VDD1.n76 B 0.030603f
C93 VDD1.n77 B 0.013709f
C94 VDD1.n78 B 0.024094f
C95 VDD1.n79 B 0.012947f
C96 VDD1.n80 B 0.030603f
C97 VDD1.n81 B 0.013709f
C98 VDD1.n82 B 0.024094f
C99 VDD1.n83 B 0.012947f
C100 VDD1.n84 B 0.022952f
C101 VDD1.n85 B 0.021634f
C102 VDD1.t3 B 0.051705f
C103 VDD1.n86 B 0.175105f
C104 VDD1.n87 B 1.23159f
C105 VDD1.n88 B 0.012947f
C106 VDD1.n89 B 0.013709f
C107 VDD1.n90 B 0.030603f
C108 VDD1.n91 B 0.030603f
C109 VDD1.n92 B 0.013709f
C110 VDD1.n93 B 0.012947f
C111 VDD1.n94 B 0.024094f
C112 VDD1.n95 B 0.024094f
C113 VDD1.n96 B 0.012947f
C114 VDD1.n97 B 0.013709f
C115 VDD1.n98 B 0.030603f
C116 VDD1.n99 B 0.030603f
C117 VDD1.n100 B 0.013709f
C118 VDD1.n101 B 0.012947f
C119 VDD1.n102 B 0.024094f
C120 VDD1.n103 B 0.024094f
C121 VDD1.n104 B 0.012947f
C122 VDD1.n105 B 0.012947f
C123 VDD1.n106 B 0.013709f
C124 VDD1.n107 B 0.030603f
C125 VDD1.n108 B 0.030603f
C126 VDD1.n109 B 0.030603f
C127 VDD1.n110 B 0.013328f
C128 VDD1.n111 B 0.012947f
C129 VDD1.n112 B 0.024094f
C130 VDD1.n113 B 0.024094f
C131 VDD1.n114 B 0.012947f
C132 VDD1.n115 B 0.013709f
C133 VDD1.n116 B 0.030603f
C134 VDD1.n117 B 0.030603f
C135 VDD1.n118 B 0.013709f
C136 VDD1.n119 B 0.012947f
C137 VDD1.n120 B 0.024094f
C138 VDD1.n121 B 0.024094f
C139 VDD1.n122 B 0.012947f
C140 VDD1.n123 B 0.013709f
C141 VDD1.n124 B 0.030603f
C142 VDD1.n125 B 0.067112f
C143 VDD1.n126 B 0.013709f
C144 VDD1.n127 B 0.012947f
C145 VDD1.n128 B 0.05668f
C146 VDD1.n129 B 0.055269f
C147 VDD1.t1 B 0.231337f
C148 VDD1.t2 B 0.231337f
C149 VDD1.n130 B 2.06395f
C150 VDD1.n131 B 1.821f
C151 VDD1.t0 B 0.231337f
C152 VDD1.t4 B 0.231337f
C153 VDD1.n132 B 2.0633f
C154 VDD1.n133 B 2.15384f
C155 VP.n0 B 0.066353f
C156 VP.t0 B 1.03745f
C157 VP.n1 B 0.390759f
C158 VP.t1 B 1.01889f
C159 VP.t5 B 1.01889f
C160 VP.n2 B 0.419572f
C161 VP.n3 B 0.408261f
C162 VP.n4 B 2.13431f
C163 VP.n5 B 2.03304f
C164 VP.t2 B 1.01889f
C165 VP.n6 B 0.408261f
C166 VP.t4 B 1.01889f
C167 VP.n7 B 0.419572f
C168 VP.t3 B 1.01889f
C169 VP.n8 B 0.408261f
C170 VP.n9 B 0.055292f
C171 VTAIL.t8 B 0.238752f
C172 VTAIL.t11 B 0.238752f
C173 VTAIL.n0 B 2.05626f
C174 VTAIL.n1 B 0.334948f
C175 VTAIL.n2 B 0.035456f
C176 VTAIL.n3 B 0.024867f
C177 VTAIL.n4 B 0.013362f
C178 VTAIL.n5 B 0.031583f
C179 VTAIL.n6 B 0.014148f
C180 VTAIL.n7 B 0.024867f
C181 VTAIL.n8 B 0.013362f
C182 VTAIL.n9 B 0.031583f
C183 VTAIL.n10 B 0.014148f
C184 VTAIL.n11 B 0.024867f
C185 VTAIL.n12 B 0.013755f
C186 VTAIL.n13 B 0.031583f
C187 VTAIL.n14 B 0.014148f
C188 VTAIL.n15 B 0.024867f
C189 VTAIL.n16 B 0.013362f
C190 VTAIL.n17 B 0.031583f
C191 VTAIL.n18 B 0.014148f
C192 VTAIL.n19 B 0.024867f
C193 VTAIL.n20 B 0.013362f
C194 VTAIL.n21 B 0.023688f
C195 VTAIL.n22 B 0.022327f
C196 VTAIL.t2 B 0.053363f
C197 VTAIL.n23 B 0.180718f
C198 VTAIL.n24 B 1.27107f
C199 VTAIL.n25 B 0.013362f
C200 VTAIL.n26 B 0.014148f
C201 VTAIL.n27 B 0.031583f
C202 VTAIL.n28 B 0.031583f
C203 VTAIL.n29 B 0.014148f
C204 VTAIL.n30 B 0.013362f
C205 VTAIL.n31 B 0.024867f
C206 VTAIL.n32 B 0.024867f
C207 VTAIL.n33 B 0.013362f
C208 VTAIL.n34 B 0.014148f
C209 VTAIL.n35 B 0.031583f
C210 VTAIL.n36 B 0.031583f
C211 VTAIL.n37 B 0.014148f
C212 VTAIL.n38 B 0.013362f
C213 VTAIL.n39 B 0.024867f
C214 VTAIL.n40 B 0.024867f
C215 VTAIL.n41 B 0.013362f
C216 VTAIL.n42 B 0.013362f
C217 VTAIL.n43 B 0.014148f
C218 VTAIL.n44 B 0.031583f
C219 VTAIL.n45 B 0.031583f
C220 VTAIL.n46 B 0.031583f
C221 VTAIL.n47 B 0.013755f
C222 VTAIL.n48 B 0.013362f
C223 VTAIL.n49 B 0.024867f
C224 VTAIL.n50 B 0.024867f
C225 VTAIL.n51 B 0.013362f
C226 VTAIL.n52 B 0.014148f
C227 VTAIL.n53 B 0.031583f
C228 VTAIL.n54 B 0.031583f
C229 VTAIL.n55 B 0.014148f
C230 VTAIL.n56 B 0.013362f
C231 VTAIL.n57 B 0.024867f
C232 VTAIL.n58 B 0.024867f
C233 VTAIL.n59 B 0.013362f
C234 VTAIL.n60 B 0.014148f
C235 VTAIL.n61 B 0.031583f
C236 VTAIL.n62 B 0.069263f
C237 VTAIL.n63 B 0.014148f
C238 VTAIL.n64 B 0.013362f
C239 VTAIL.n65 B 0.058497f
C240 VTAIL.n66 B 0.038878f
C241 VTAIL.n67 B 0.154781f
C242 VTAIL.t4 B 0.238752f
C243 VTAIL.t1 B 0.238752f
C244 VTAIL.n68 B 2.05626f
C245 VTAIL.n69 B 1.61266f
C246 VTAIL.t6 B 0.238752f
C247 VTAIL.t9 B 0.238752f
C248 VTAIL.n70 B 2.05627f
C249 VTAIL.n71 B 1.61265f
C250 VTAIL.n72 B 0.035456f
C251 VTAIL.n73 B 0.024867f
C252 VTAIL.n74 B 0.013362f
C253 VTAIL.n75 B 0.031583f
C254 VTAIL.n76 B 0.014148f
C255 VTAIL.n77 B 0.024867f
C256 VTAIL.n78 B 0.013362f
C257 VTAIL.n79 B 0.031583f
C258 VTAIL.n80 B 0.014148f
C259 VTAIL.n81 B 0.024867f
C260 VTAIL.n82 B 0.013755f
C261 VTAIL.n83 B 0.031583f
C262 VTAIL.n84 B 0.013362f
C263 VTAIL.n85 B 0.014148f
C264 VTAIL.n86 B 0.024867f
C265 VTAIL.n87 B 0.013362f
C266 VTAIL.n88 B 0.031583f
C267 VTAIL.n89 B 0.014148f
C268 VTAIL.n90 B 0.024867f
C269 VTAIL.n91 B 0.013362f
C270 VTAIL.n92 B 0.023688f
C271 VTAIL.n93 B 0.022327f
C272 VTAIL.t7 B 0.053363f
C273 VTAIL.n94 B 0.180718f
C274 VTAIL.n95 B 1.27107f
C275 VTAIL.n96 B 0.013362f
C276 VTAIL.n97 B 0.014148f
C277 VTAIL.n98 B 0.031583f
C278 VTAIL.n99 B 0.031583f
C279 VTAIL.n100 B 0.014148f
C280 VTAIL.n101 B 0.013362f
C281 VTAIL.n102 B 0.024867f
C282 VTAIL.n103 B 0.024867f
C283 VTAIL.n104 B 0.013362f
C284 VTAIL.n105 B 0.014148f
C285 VTAIL.n106 B 0.031583f
C286 VTAIL.n107 B 0.031583f
C287 VTAIL.n108 B 0.014148f
C288 VTAIL.n109 B 0.013362f
C289 VTAIL.n110 B 0.024867f
C290 VTAIL.n111 B 0.024867f
C291 VTAIL.n112 B 0.013362f
C292 VTAIL.n113 B 0.014148f
C293 VTAIL.n114 B 0.031583f
C294 VTAIL.n115 B 0.031583f
C295 VTAIL.n116 B 0.031583f
C296 VTAIL.n117 B 0.013755f
C297 VTAIL.n118 B 0.013362f
C298 VTAIL.n119 B 0.024867f
C299 VTAIL.n120 B 0.024867f
C300 VTAIL.n121 B 0.013362f
C301 VTAIL.n122 B 0.014148f
C302 VTAIL.n123 B 0.031583f
C303 VTAIL.n124 B 0.031583f
C304 VTAIL.n125 B 0.014148f
C305 VTAIL.n126 B 0.013362f
C306 VTAIL.n127 B 0.024867f
C307 VTAIL.n128 B 0.024867f
C308 VTAIL.n129 B 0.013362f
C309 VTAIL.n130 B 0.014148f
C310 VTAIL.n131 B 0.031583f
C311 VTAIL.n132 B 0.069263f
C312 VTAIL.n133 B 0.014148f
C313 VTAIL.n134 B 0.013362f
C314 VTAIL.n135 B 0.058497f
C315 VTAIL.n136 B 0.038878f
C316 VTAIL.n137 B 0.154781f
C317 VTAIL.t5 B 0.238752f
C318 VTAIL.t0 B 0.238752f
C319 VTAIL.n138 B 2.05627f
C320 VTAIL.n139 B 0.377935f
C321 VTAIL.n140 B 0.035456f
C322 VTAIL.n141 B 0.024867f
C323 VTAIL.n142 B 0.013362f
C324 VTAIL.n143 B 0.031583f
C325 VTAIL.n144 B 0.014148f
C326 VTAIL.n145 B 0.024867f
C327 VTAIL.n146 B 0.013362f
C328 VTAIL.n147 B 0.031583f
C329 VTAIL.n148 B 0.014148f
C330 VTAIL.n149 B 0.024867f
C331 VTAIL.n150 B 0.013755f
C332 VTAIL.n151 B 0.031583f
C333 VTAIL.n152 B 0.013362f
C334 VTAIL.n153 B 0.014148f
C335 VTAIL.n154 B 0.024867f
C336 VTAIL.n155 B 0.013362f
C337 VTAIL.n156 B 0.031583f
C338 VTAIL.n157 B 0.014148f
C339 VTAIL.n158 B 0.024867f
C340 VTAIL.n159 B 0.013362f
C341 VTAIL.n160 B 0.023688f
C342 VTAIL.n161 B 0.022327f
C343 VTAIL.t3 B 0.053363f
C344 VTAIL.n162 B 0.180718f
C345 VTAIL.n163 B 1.27107f
C346 VTAIL.n164 B 0.013362f
C347 VTAIL.n165 B 0.014148f
C348 VTAIL.n166 B 0.031583f
C349 VTAIL.n167 B 0.031583f
C350 VTAIL.n168 B 0.014148f
C351 VTAIL.n169 B 0.013362f
C352 VTAIL.n170 B 0.024867f
C353 VTAIL.n171 B 0.024867f
C354 VTAIL.n172 B 0.013362f
C355 VTAIL.n173 B 0.014148f
C356 VTAIL.n174 B 0.031583f
C357 VTAIL.n175 B 0.031583f
C358 VTAIL.n176 B 0.014148f
C359 VTAIL.n177 B 0.013362f
C360 VTAIL.n178 B 0.024867f
C361 VTAIL.n179 B 0.024867f
C362 VTAIL.n180 B 0.013362f
C363 VTAIL.n181 B 0.014148f
C364 VTAIL.n182 B 0.031583f
C365 VTAIL.n183 B 0.031583f
C366 VTAIL.n184 B 0.031583f
C367 VTAIL.n185 B 0.013755f
C368 VTAIL.n186 B 0.013362f
C369 VTAIL.n187 B 0.024867f
C370 VTAIL.n188 B 0.024867f
C371 VTAIL.n189 B 0.013362f
C372 VTAIL.n190 B 0.014148f
C373 VTAIL.n191 B 0.031583f
C374 VTAIL.n192 B 0.031583f
C375 VTAIL.n193 B 0.014148f
C376 VTAIL.n194 B 0.013362f
C377 VTAIL.n195 B 0.024867f
C378 VTAIL.n196 B 0.024867f
C379 VTAIL.n197 B 0.013362f
C380 VTAIL.n198 B 0.014148f
C381 VTAIL.n199 B 0.031583f
C382 VTAIL.n200 B 0.069263f
C383 VTAIL.n201 B 0.014148f
C384 VTAIL.n202 B 0.013362f
C385 VTAIL.n203 B 0.058497f
C386 VTAIL.n204 B 0.038878f
C387 VTAIL.n205 B 1.32594f
C388 VTAIL.n206 B 0.035456f
C389 VTAIL.n207 B 0.024867f
C390 VTAIL.n208 B 0.013362f
C391 VTAIL.n209 B 0.031583f
C392 VTAIL.n210 B 0.014148f
C393 VTAIL.n211 B 0.024867f
C394 VTAIL.n212 B 0.013362f
C395 VTAIL.n213 B 0.031583f
C396 VTAIL.n214 B 0.014148f
C397 VTAIL.n215 B 0.024867f
C398 VTAIL.n216 B 0.013755f
C399 VTAIL.n217 B 0.031583f
C400 VTAIL.n218 B 0.014148f
C401 VTAIL.n219 B 0.024867f
C402 VTAIL.n220 B 0.013362f
C403 VTAIL.n221 B 0.031583f
C404 VTAIL.n222 B 0.014148f
C405 VTAIL.n223 B 0.024867f
C406 VTAIL.n224 B 0.013362f
C407 VTAIL.n225 B 0.023688f
C408 VTAIL.n226 B 0.022327f
C409 VTAIL.t10 B 0.053363f
C410 VTAIL.n227 B 0.180718f
C411 VTAIL.n228 B 1.27107f
C412 VTAIL.n229 B 0.013362f
C413 VTAIL.n230 B 0.014148f
C414 VTAIL.n231 B 0.031583f
C415 VTAIL.n232 B 0.031583f
C416 VTAIL.n233 B 0.014148f
C417 VTAIL.n234 B 0.013362f
C418 VTAIL.n235 B 0.024867f
C419 VTAIL.n236 B 0.024867f
C420 VTAIL.n237 B 0.013362f
C421 VTAIL.n238 B 0.014148f
C422 VTAIL.n239 B 0.031583f
C423 VTAIL.n240 B 0.031583f
C424 VTAIL.n241 B 0.014148f
C425 VTAIL.n242 B 0.013362f
C426 VTAIL.n243 B 0.024867f
C427 VTAIL.n244 B 0.024867f
C428 VTAIL.n245 B 0.013362f
C429 VTAIL.n246 B 0.013362f
C430 VTAIL.n247 B 0.014148f
C431 VTAIL.n248 B 0.031583f
C432 VTAIL.n249 B 0.031583f
C433 VTAIL.n250 B 0.031583f
C434 VTAIL.n251 B 0.013755f
C435 VTAIL.n252 B 0.013362f
C436 VTAIL.n253 B 0.024867f
C437 VTAIL.n254 B 0.024867f
C438 VTAIL.n255 B 0.013362f
C439 VTAIL.n256 B 0.014148f
C440 VTAIL.n257 B 0.031583f
C441 VTAIL.n258 B 0.031583f
C442 VTAIL.n259 B 0.014148f
C443 VTAIL.n260 B 0.013362f
C444 VTAIL.n261 B 0.024867f
C445 VTAIL.n262 B 0.024867f
C446 VTAIL.n263 B 0.013362f
C447 VTAIL.n264 B 0.014148f
C448 VTAIL.n265 B 0.031583f
C449 VTAIL.n266 B 0.069263f
C450 VTAIL.n267 B 0.014148f
C451 VTAIL.n268 B 0.013362f
C452 VTAIL.n269 B 0.058497f
C453 VTAIL.n270 B 0.038878f
C454 VTAIL.n271 B 1.3054f
C455 VDD2.n0 B 0.034097f
C456 VDD2.n1 B 0.023914f
C457 VDD2.n2 B 0.01285f
C458 VDD2.n3 B 0.030373f
C459 VDD2.n4 B 0.013606f
C460 VDD2.n5 B 0.023914f
C461 VDD2.n6 B 0.01285f
C462 VDD2.n7 B 0.030373f
C463 VDD2.n8 B 0.013606f
C464 VDD2.n9 B 0.023914f
C465 VDD2.n10 B 0.013228f
C466 VDD2.n11 B 0.030373f
C467 VDD2.n12 B 0.013606f
C468 VDD2.n13 B 0.023914f
C469 VDD2.n14 B 0.01285f
C470 VDD2.n15 B 0.030373f
C471 VDD2.n16 B 0.013606f
C472 VDD2.n17 B 0.023914f
C473 VDD2.n18 B 0.01285f
C474 VDD2.n19 B 0.02278f
C475 VDD2.n20 B 0.021472f
C476 VDD2.t1 B 0.051318f
C477 VDD2.n21 B 0.173793f
C478 VDD2.n22 B 1.22236f
C479 VDD2.n23 B 0.01285f
C480 VDD2.n24 B 0.013606f
C481 VDD2.n25 B 0.030373f
C482 VDD2.n26 B 0.030373f
C483 VDD2.n27 B 0.013606f
C484 VDD2.n28 B 0.01285f
C485 VDD2.n29 B 0.023914f
C486 VDD2.n30 B 0.023914f
C487 VDD2.n31 B 0.01285f
C488 VDD2.n32 B 0.013606f
C489 VDD2.n33 B 0.030373f
C490 VDD2.n34 B 0.030373f
C491 VDD2.n35 B 0.013606f
C492 VDD2.n36 B 0.01285f
C493 VDD2.n37 B 0.023914f
C494 VDD2.n38 B 0.023914f
C495 VDD2.n39 B 0.01285f
C496 VDD2.n40 B 0.01285f
C497 VDD2.n41 B 0.013606f
C498 VDD2.n42 B 0.030373f
C499 VDD2.n43 B 0.030373f
C500 VDD2.n44 B 0.030373f
C501 VDD2.n45 B 0.013228f
C502 VDD2.n46 B 0.01285f
C503 VDD2.n47 B 0.023914f
C504 VDD2.n48 B 0.023914f
C505 VDD2.n49 B 0.01285f
C506 VDD2.n50 B 0.013606f
C507 VDD2.n51 B 0.030373f
C508 VDD2.n52 B 0.030373f
C509 VDD2.n53 B 0.013606f
C510 VDD2.n54 B 0.01285f
C511 VDD2.n55 B 0.023914f
C512 VDD2.n56 B 0.023914f
C513 VDD2.n57 B 0.01285f
C514 VDD2.n58 B 0.013606f
C515 VDD2.n59 B 0.030373f
C516 VDD2.n60 B 0.066609f
C517 VDD2.n61 B 0.013606f
C518 VDD2.n62 B 0.01285f
C519 VDD2.n63 B 0.056256f
C520 VDD2.n64 B 0.054855f
C521 VDD2.t4 B 0.229603f
C522 VDD2.t0 B 0.229603f
C523 VDD2.n65 B 2.04848f
C524 VDD2.n66 B 1.73597f
C525 VDD2.n67 B 0.034097f
C526 VDD2.n68 B 0.023914f
C527 VDD2.n69 B 0.01285f
C528 VDD2.n70 B 0.030373f
C529 VDD2.n71 B 0.013606f
C530 VDD2.n72 B 0.023914f
C531 VDD2.n73 B 0.01285f
C532 VDD2.n74 B 0.030373f
C533 VDD2.n75 B 0.013606f
C534 VDD2.n76 B 0.023914f
C535 VDD2.n77 B 0.013228f
C536 VDD2.n78 B 0.030373f
C537 VDD2.n79 B 0.01285f
C538 VDD2.n80 B 0.013606f
C539 VDD2.n81 B 0.023914f
C540 VDD2.n82 B 0.01285f
C541 VDD2.n83 B 0.030373f
C542 VDD2.n84 B 0.013606f
C543 VDD2.n85 B 0.023914f
C544 VDD2.n86 B 0.01285f
C545 VDD2.n87 B 0.02278f
C546 VDD2.n88 B 0.021472f
C547 VDD2.t5 B 0.051318f
C548 VDD2.n89 B 0.173793f
C549 VDD2.n90 B 1.22236f
C550 VDD2.n91 B 0.01285f
C551 VDD2.n92 B 0.013606f
C552 VDD2.n93 B 0.030373f
C553 VDD2.n94 B 0.030373f
C554 VDD2.n95 B 0.013606f
C555 VDD2.n96 B 0.01285f
C556 VDD2.n97 B 0.023914f
C557 VDD2.n98 B 0.023914f
C558 VDD2.n99 B 0.01285f
C559 VDD2.n100 B 0.013606f
C560 VDD2.n101 B 0.030373f
C561 VDD2.n102 B 0.030373f
C562 VDD2.n103 B 0.013606f
C563 VDD2.n104 B 0.01285f
C564 VDD2.n105 B 0.023914f
C565 VDD2.n106 B 0.023914f
C566 VDD2.n107 B 0.01285f
C567 VDD2.n108 B 0.013606f
C568 VDD2.n109 B 0.030373f
C569 VDD2.n110 B 0.030373f
C570 VDD2.n111 B 0.030373f
C571 VDD2.n112 B 0.013228f
C572 VDD2.n113 B 0.01285f
C573 VDD2.n114 B 0.023914f
C574 VDD2.n115 B 0.023914f
C575 VDD2.n116 B 0.01285f
C576 VDD2.n117 B 0.013606f
C577 VDD2.n118 B 0.030373f
C578 VDD2.n119 B 0.030373f
C579 VDD2.n120 B 0.013606f
C580 VDD2.n121 B 0.01285f
C581 VDD2.n122 B 0.023914f
C582 VDD2.n123 B 0.023914f
C583 VDD2.n124 B 0.01285f
C584 VDD2.n125 B 0.013606f
C585 VDD2.n126 B 0.030373f
C586 VDD2.n127 B 0.066609f
C587 VDD2.n128 B 0.013606f
C588 VDD2.n129 B 0.01285f
C589 VDD2.n130 B 0.056256f
C590 VDD2.n131 B 0.053892f
C591 VDD2.n132 B 1.93842f
C592 VDD2.t2 B 0.229603f
C593 VDD2.t3 B 0.229603f
C594 VDD2.n133 B 2.04846f
C595 VN.t3 B 1.01585f
C596 VN.n0 B 0.382623f
C597 VN.t0 B 0.997672f
C598 VN.n1 B 0.410835f
C599 VN.t1 B 0.997672f
C600 VN.n2 B 0.39976f
C601 VN.n3 B 0.196135f
C602 VN.t4 B 1.01585f
C603 VN.n4 B 0.382623f
C604 VN.t2 B 0.997672f
C605 VN.n5 B 0.410835f
C606 VN.t5 B 0.997672f
C607 VN.n6 B 0.39976f
C608 VN.n7 B 2.12196f
.ends

