* NGSPICE file created from diff_pair_sample_0284.ext - technology: sky130A

.subckt diff_pair_sample_0284 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=0.79
X1 VTAIL.t3 VN.t0 VDD2.t3 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=0.79
X2 B.t11 B.t9 B.t10 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=0.79
X3 VTAIL.t5 VP.t1 VDD1.t2 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=0.79
X4 VTAIL.t7 VP.t2 VDD1.t1 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=0.79
X5 VDD2.t2 VN.t1 VTAIL.t0 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=0.79
X6 B.t8 B.t6 B.t7 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=0.79
X7 B.t5 B.t3 B.t4 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=0.79
X8 VTAIL.t1 VN.t2 VDD2.t1 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0.99165 ps=6.34 w=6.01 l=0.79
X9 VDD2.t0 VN.t3 VTAIL.t2 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=0.79
X10 B.t2 B.t0 B.t1 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=2.3439 pd=12.8 as=0 ps=0 w=6.01 l=0.79
X11 VDD1.t0 VP.t3 VTAIL.t6 w_n1642_n2170# sky130_fd_pr__pfet_01v8 ad=0.99165 pd=6.34 as=2.3439 ps=12.8 w=6.01 l=0.79
R0 VP.n1 VP.t2 254.37
R1 VP.n1 VP.t3 254.321
R2 VP.n3 VP.t1 233.374
R3 VP.n5 VP.t0 233.374
R4 VP.n6 VP.n5 161.3
R5 VP.n4 VP.n0 161.3
R6 VP.n3 VP.n2 161.3
R7 VP.n2 VP.n1 80.8742
R8 VP.n4 VP.n3 24.1005
R9 VP.n5 VP.n4 24.1005
R10 VP.n2 VP.n0 0.189894
R11 VP.n6 VP.n0 0.189894
R12 VP VP.n6 0.0516364
R13 VTAIL.n250 VTAIL.n224 756.745
R14 VTAIL.n26 VTAIL.n0 756.745
R15 VTAIL.n58 VTAIL.n32 756.745
R16 VTAIL.n90 VTAIL.n64 756.745
R17 VTAIL.n218 VTAIL.n192 756.745
R18 VTAIL.n186 VTAIL.n160 756.745
R19 VTAIL.n154 VTAIL.n128 756.745
R20 VTAIL.n122 VTAIL.n96 756.745
R21 VTAIL.n235 VTAIL.n234 585
R22 VTAIL.n232 VTAIL.n231 585
R23 VTAIL.n241 VTAIL.n240 585
R24 VTAIL.n243 VTAIL.n242 585
R25 VTAIL.n228 VTAIL.n227 585
R26 VTAIL.n249 VTAIL.n248 585
R27 VTAIL.n251 VTAIL.n250 585
R28 VTAIL.n11 VTAIL.n10 585
R29 VTAIL.n8 VTAIL.n7 585
R30 VTAIL.n17 VTAIL.n16 585
R31 VTAIL.n19 VTAIL.n18 585
R32 VTAIL.n4 VTAIL.n3 585
R33 VTAIL.n25 VTAIL.n24 585
R34 VTAIL.n27 VTAIL.n26 585
R35 VTAIL.n43 VTAIL.n42 585
R36 VTAIL.n40 VTAIL.n39 585
R37 VTAIL.n49 VTAIL.n48 585
R38 VTAIL.n51 VTAIL.n50 585
R39 VTAIL.n36 VTAIL.n35 585
R40 VTAIL.n57 VTAIL.n56 585
R41 VTAIL.n59 VTAIL.n58 585
R42 VTAIL.n75 VTAIL.n74 585
R43 VTAIL.n72 VTAIL.n71 585
R44 VTAIL.n81 VTAIL.n80 585
R45 VTAIL.n83 VTAIL.n82 585
R46 VTAIL.n68 VTAIL.n67 585
R47 VTAIL.n89 VTAIL.n88 585
R48 VTAIL.n91 VTAIL.n90 585
R49 VTAIL.n219 VTAIL.n218 585
R50 VTAIL.n217 VTAIL.n216 585
R51 VTAIL.n196 VTAIL.n195 585
R52 VTAIL.n211 VTAIL.n210 585
R53 VTAIL.n209 VTAIL.n208 585
R54 VTAIL.n200 VTAIL.n199 585
R55 VTAIL.n203 VTAIL.n202 585
R56 VTAIL.n187 VTAIL.n186 585
R57 VTAIL.n185 VTAIL.n184 585
R58 VTAIL.n164 VTAIL.n163 585
R59 VTAIL.n179 VTAIL.n178 585
R60 VTAIL.n177 VTAIL.n176 585
R61 VTAIL.n168 VTAIL.n167 585
R62 VTAIL.n171 VTAIL.n170 585
R63 VTAIL.n155 VTAIL.n154 585
R64 VTAIL.n153 VTAIL.n152 585
R65 VTAIL.n132 VTAIL.n131 585
R66 VTAIL.n147 VTAIL.n146 585
R67 VTAIL.n145 VTAIL.n144 585
R68 VTAIL.n136 VTAIL.n135 585
R69 VTAIL.n139 VTAIL.n138 585
R70 VTAIL.n123 VTAIL.n122 585
R71 VTAIL.n121 VTAIL.n120 585
R72 VTAIL.n100 VTAIL.n99 585
R73 VTAIL.n115 VTAIL.n114 585
R74 VTAIL.n113 VTAIL.n112 585
R75 VTAIL.n104 VTAIL.n103 585
R76 VTAIL.n107 VTAIL.n106 585
R77 VTAIL.t2 VTAIL.n233 327.601
R78 VTAIL.t1 VTAIL.n9 327.601
R79 VTAIL.t4 VTAIL.n41 327.601
R80 VTAIL.t5 VTAIL.n73 327.601
R81 VTAIL.t6 VTAIL.n201 327.601
R82 VTAIL.t7 VTAIL.n169 327.601
R83 VTAIL.t0 VTAIL.n137 327.601
R84 VTAIL.t3 VTAIL.n105 327.601
R85 VTAIL.n234 VTAIL.n231 171.744
R86 VTAIL.n241 VTAIL.n231 171.744
R87 VTAIL.n242 VTAIL.n241 171.744
R88 VTAIL.n242 VTAIL.n227 171.744
R89 VTAIL.n249 VTAIL.n227 171.744
R90 VTAIL.n250 VTAIL.n249 171.744
R91 VTAIL.n10 VTAIL.n7 171.744
R92 VTAIL.n17 VTAIL.n7 171.744
R93 VTAIL.n18 VTAIL.n17 171.744
R94 VTAIL.n18 VTAIL.n3 171.744
R95 VTAIL.n25 VTAIL.n3 171.744
R96 VTAIL.n26 VTAIL.n25 171.744
R97 VTAIL.n42 VTAIL.n39 171.744
R98 VTAIL.n49 VTAIL.n39 171.744
R99 VTAIL.n50 VTAIL.n49 171.744
R100 VTAIL.n50 VTAIL.n35 171.744
R101 VTAIL.n57 VTAIL.n35 171.744
R102 VTAIL.n58 VTAIL.n57 171.744
R103 VTAIL.n74 VTAIL.n71 171.744
R104 VTAIL.n81 VTAIL.n71 171.744
R105 VTAIL.n82 VTAIL.n81 171.744
R106 VTAIL.n82 VTAIL.n67 171.744
R107 VTAIL.n89 VTAIL.n67 171.744
R108 VTAIL.n90 VTAIL.n89 171.744
R109 VTAIL.n218 VTAIL.n217 171.744
R110 VTAIL.n217 VTAIL.n195 171.744
R111 VTAIL.n210 VTAIL.n195 171.744
R112 VTAIL.n210 VTAIL.n209 171.744
R113 VTAIL.n209 VTAIL.n199 171.744
R114 VTAIL.n202 VTAIL.n199 171.744
R115 VTAIL.n186 VTAIL.n185 171.744
R116 VTAIL.n185 VTAIL.n163 171.744
R117 VTAIL.n178 VTAIL.n163 171.744
R118 VTAIL.n178 VTAIL.n177 171.744
R119 VTAIL.n177 VTAIL.n167 171.744
R120 VTAIL.n170 VTAIL.n167 171.744
R121 VTAIL.n154 VTAIL.n153 171.744
R122 VTAIL.n153 VTAIL.n131 171.744
R123 VTAIL.n146 VTAIL.n131 171.744
R124 VTAIL.n146 VTAIL.n145 171.744
R125 VTAIL.n145 VTAIL.n135 171.744
R126 VTAIL.n138 VTAIL.n135 171.744
R127 VTAIL.n122 VTAIL.n121 171.744
R128 VTAIL.n121 VTAIL.n99 171.744
R129 VTAIL.n114 VTAIL.n99 171.744
R130 VTAIL.n114 VTAIL.n113 171.744
R131 VTAIL.n113 VTAIL.n103 171.744
R132 VTAIL.n106 VTAIL.n103 171.744
R133 VTAIL.n234 VTAIL.t2 85.8723
R134 VTAIL.n10 VTAIL.t1 85.8723
R135 VTAIL.n42 VTAIL.t4 85.8723
R136 VTAIL.n74 VTAIL.t5 85.8723
R137 VTAIL.n202 VTAIL.t6 85.8723
R138 VTAIL.n170 VTAIL.t7 85.8723
R139 VTAIL.n138 VTAIL.t0 85.8723
R140 VTAIL.n106 VTAIL.t3 85.8723
R141 VTAIL.n255 VTAIL.n254 32.3793
R142 VTAIL.n31 VTAIL.n30 32.3793
R143 VTAIL.n63 VTAIL.n62 32.3793
R144 VTAIL.n95 VTAIL.n94 32.3793
R145 VTAIL.n223 VTAIL.n222 32.3793
R146 VTAIL.n191 VTAIL.n190 32.3793
R147 VTAIL.n159 VTAIL.n158 32.3793
R148 VTAIL.n127 VTAIL.n126 32.3793
R149 VTAIL.n255 VTAIL.n223 18.5134
R150 VTAIL.n127 VTAIL.n95 18.5134
R151 VTAIL.n235 VTAIL.n233 16.3865
R152 VTAIL.n11 VTAIL.n9 16.3865
R153 VTAIL.n43 VTAIL.n41 16.3865
R154 VTAIL.n75 VTAIL.n73 16.3865
R155 VTAIL.n203 VTAIL.n201 16.3865
R156 VTAIL.n171 VTAIL.n169 16.3865
R157 VTAIL.n139 VTAIL.n137 16.3865
R158 VTAIL.n107 VTAIL.n105 16.3865
R159 VTAIL.n236 VTAIL.n232 12.8005
R160 VTAIL.n12 VTAIL.n8 12.8005
R161 VTAIL.n44 VTAIL.n40 12.8005
R162 VTAIL.n76 VTAIL.n72 12.8005
R163 VTAIL.n204 VTAIL.n200 12.8005
R164 VTAIL.n172 VTAIL.n168 12.8005
R165 VTAIL.n140 VTAIL.n136 12.8005
R166 VTAIL.n108 VTAIL.n104 12.8005
R167 VTAIL.n240 VTAIL.n239 12.0247
R168 VTAIL.n16 VTAIL.n15 12.0247
R169 VTAIL.n48 VTAIL.n47 12.0247
R170 VTAIL.n80 VTAIL.n79 12.0247
R171 VTAIL.n208 VTAIL.n207 12.0247
R172 VTAIL.n176 VTAIL.n175 12.0247
R173 VTAIL.n144 VTAIL.n143 12.0247
R174 VTAIL.n112 VTAIL.n111 12.0247
R175 VTAIL.n243 VTAIL.n230 11.249
R176 VTAIL.n19 VTAIL.n6 11.249
R177 VTAIL.n51 VTAIL.n38 11.249
R178 VTAIL.n83 VTAIL.n70 11.249
R179 VTAIL.n211 VTAIL.n198 11.249
R180 VTAIL.n179 VTAIL.n166 11.249
R181 VTAIL.n147 VTAIL.n134 11.249
R182 VTAIL.n115 VTAIL.n102 11.249
R183 VTAIL.n244 VTAIL.n228 10.4732
R184 VTAIL.n20 VTAIL.n4 10.4732
R185 VTAIL.n52 VTAIL.n36 10.4732
R186 VTAIL.n84 VTAIL.n68 10.4732
R187 VTAIL.n212 VTAIL.n196 10.4732
R188 VTAIL.n180 VTAIL.n164 10.4732
R189 VTAIL.n148 VTAIL.n132 10.4732
R190 VTAIL.n116 VTAIL.n100 10.4732
R191 VTAIL.n248 VTAIL.n247 9.69747
R192 VTAIL.n24 VTAIL.n23 9.69747
R193 VTAIL.n56 VTAIL.n55 9.69747
R194 VTAIL.n88 VTAIL.n87 9.69747
R195 VTAIL.n216 VTAIL.n215 9.69747
R196 VTAIL.n184 VTAIL.n183 9.69747
R197 VTAIL.n152 VTAIL.n151 9.69747
R198 VTAIL.n120 VTAIL.n119 9.69747
R199 VTAIL.n254 VTAIL.n253 9.45567
R200 VTAIL.n30 VTAIL.n29 9.45567
R201 VTAIL.n62 VTAIL.n61 9.45567
R202 VTAIL.n94 VTAIL.n93 9.45567
R203 VTAIL.n222 VTAIL.n221 9.45567
R204 VTAIL.n190 VTAIL.n189 9.45567
R205 VTAIL.n158 VTAIL.n157 9.45567
R206 VTAIL.n126 VTAIL.n125 9.45567
R207 VTAIL.n253 VTAIL.n252 9.3005
R208 VTAIL.n226 VTAIL.n225 9.3005
R209 VTAIL.n247 VTAIL.n246 9.3005
R210 VTAIL.n245 VTAIL.n244 9.3005
R211 VTAIL.n230 VTAIL.n229 9.3005
R212 VTAIL.n239 VTAIL.n238 9.3005
R213 VTAIL.n237 VTAIL.n236 9.3005
R214 VTAIL.n29 VTAIL.n28 9.3005
R215 VTAIL.n2 VTAIL.n1 9.3005
R216 VTAIL.n23 VTAIL.n22 9.3005
R217 VTAIL.n21 VTAIL.n20 9.3005
R218 VTAIL.n6 VTAIL.n5 9.3005
R219 VTAIL.n15 VTAIL.n14 9.3005
R220 VTAIL.n13 VTAIL.n12 9.3005
R221 VTAIL.n61 VTAIL.n60 9.3005
R222 VTAIL.n34 VTAIL.n33 9.3005
R223 VTAIL.n55 VTAIL.n54 9.3005
R224 VTAIL.n53 VTAIL.n52 9.3005
R225 VTAIL.n38 VTAIL.n37 9.3005
R226 VTAIL.n47 VTAIL.n46 9.3005
R227 VTAIL.n45 VTAIL.n44 9.3005
R228 VTAIL.n93 VTAIL.n92 9.3005
R229 VTAIL.n66 VTAIL.n65 9.3005
R230 VTAIL.n87 VTAIL.n86 9.3005
R231 VTAIL.n85 VTAIL.n84 9.3005
R232 VTAIL.n70 VTAIL.n69 9.3005
R233 VTAIL.n79 VTAIL.n78 9.3005
R234 VTAIL.n77 VTAIL.n76 9.3005
R235 VTAIL.n221 VTAIL.n220 9.3005
R236 VTAIL.n194 VTAIL.n193 9.3005
R237 VTAIL.n215 VTAIL.n214 9.3005
R238 VTAIL.n213 VTAIL.n212 9.3005
R239 VTAIL.n198 VTAIL.n197 9.3005
R240 VTAIL.n207 VTAIL.n206 9.3005
R241 VTAIL.n205 VTAIL.n204 9.3005
R242 VTAIL.n189 VTAIL.n188 9.3005
R243 VTAIL.n162 VTAIL.n161 9.3005
R244 VTAIL.n183 VTAIL.n182 9.3005
R245 VTAIL.n181 VTAIL.n180 9.3005
R246 VTAIL.n166 VTAIL.n165 9.3005
R247 VTAIL.n175 VTAIL.n174 9.3005
R248 VTAIL.n173 VTAIL.n172 9.3005
R249 VTAIL.n157 VTAIL.n156 9.3005
R250 VTAIL.n130 VTAIL.n129 9.3005
R251 VTAIL.n151 VTAIL.n150 9.3005
R252 VTAIL.n149 VTAIL.n148 9.3005
R253 VTAIL.n134 VTAIL.n133 9.3005
R254 VTAIL.n143 VTAIL.n142 9.3005
R255 VTAIL.n141 VTAIL.n140 9.3005
R256 VTAIL.n125 VTAIL.n124 9.3005
R257 VTAIL.n98 VTAIL.n97 9.3005
R258 VTAIL.n119 VTAIL.n118 9.3005
R259 VTAIL.n117 VTAIL.n116 9.3005
R260 VTAIL.n102 VTAIL.n101 9.3005
R261 VTAIL.n111 VTAIL.n110 9.3005
R262 VTAIL.n109 VTAIL.n108 9.3005
R263 VTAIL.n251 VTAIL.n226 8.92171
R264 VTAIL.n27 VTAIL.n2 8.92171
R265 VTAIL.n59 VTAIL.n34 8.92171
R266 VTAIL.n91 VTAIL.n66 8.92171
R267 VTAIL.n219 VTAIL.n194 8.92171
R268 VTAIL.n187 VTAIL.n162 8.92171
R269 VTAIL.n155 VTAIL.n130 8.92171
R270 VTAIL.n123 VTAIL.n98 8.92171
R271 VTAIL.n252 VTAIL.n224 8.14595
R272 VTAIL.n28 VTAIL.n0 8.14595
R273 VTAIL.n60 VTAIL.n32 8.14595
R274 VTAIL.n92 VTAIL.n64 8.14595
R275 VTAIL.n220 VTAIL.n192 8.14595
R276 VTAIL.n188 VTAIL.n160 8.14595
R277 VTAIL.n156 VTAIL.n128 8.14595
R278 VTAIL.n124 VTAIL.n96 8.14595
R279 VTAIL.n254 VTAIL.n224 5.81868
R280 VTAIL.n30 VTAIL.n0 5.81868
R281 VTAIL.n62 VTAIL.n32 5.81868
R282 VTAIL.n94 VTAIL.n64 5.81868
R283 VTAIL.n222 VTAIL.n192 5.81868
R284 VTAIL.n190 VTAIL.n160 5.81868
R285 VTAIL.n158 VTAIL.n128 5.81868
R286 VTAIL.n126 VTAIL.n96 5.81868
R287 VTAIL.n252 VTAIL.n251 5.04292
R288 VTAIL.n28 VTAIL.n27 5.04292
R289 VTAIL.n60 VTAIL.n59 5.04292
R290 VTAIL.n92 VTAIL.n91 5.04292
R291 VTAIL.n220 VTAIL.n219 5.04292
R292 VTAIL.n188 VTAIL.n187 5.04292
R293 VTAIL.n156 VTAIL.n155 5.04292
R294 VTAIL.n124 VTAIL.n123 5.04292
R295 VTAIL.n248 VTAIL.n226 4.26717
R296 VTAIL.n24 VTAIL.n2 4.26717
R297 VTAIL.n56 VTAIL.n34 4.26717
R298 VTAIL.n88 VTAIL.n66 4.26717
R299 VTAIL.n216 VTAIL.n194 4.26717
R300 VTAIL.n184 VTAIL.n162 4.26717
R301 VTAIL.n152 VTAIL.n130 4.26717
R302 VTAIL.n120 VTAIL.n98 4.26717
R303 VTAIL.n205 VTAIL.n201 3.71286
R304 VTAIL.n173 VTAIL.n169 3.71286
R305 VTAIL.n141 VTAIL.n137 3.71286
R306 VTAIL.n109 VTAIL.n105 3.71286
R307 VTAIL.n237 VTAIL.n233 3.71286
R308 VTAIL.n13 VTAIL.n9 3.71286
R309 VTAIL.n45 VTAIL.n41 3.71286
R310 VTAIL.n77 VTAIL.n73 3.71286
R311 VTAIL.n247 VTAIL.n228 3.49141
R312 VTAIL.n23 VTAIL.n4 3.49141
R313 VTAIL.n55 VTAIL.n36 3.49141
R314 VTAIL.n87 VTAIL.n68 3.49141
R315 VTAIL.n215 VTAIL.n196 3.49141
R316 VTAIL.n183 VTAIL.n164 3.49141
R317 VTAIL.n151 VTAIL.n132 3.49141
R318 VTAIL.n119 VTAIL.n100 3.49141
R319 VTAIL.n244 VTAIL.n243 2.71565
R320 VTAIL.n20 VTAIL.n19 2.71565
R321 VTAIL.n52 VTAIL.n51 2.71565
R322 VTAIL.n84 VTAIL.n83 2.71565
R323 VTAIL.n212 VTAIL.n211 2.71565
R324 VTAIL.n180 VTAIL.n179 2.71565
R325 VTAIL.n148 VTAIL.n147 2.71565
R326 VTAIL.n116 VTAIL.n115 2.71565
R327 VTAIL.n240 VTAIL.n230 1.93989
R328 VTAIL.n16 VTAIL.n6 1.93989
R329 VTAIL.n48 VTAIL.n38 1.93989
R330 VTAIL.n80 VTAIL.n70 1.93989
R331 VTAIL.n208 VTAIL.n198 1.93989
R332 VTAIL.n176 VTAIL.n166 1.93989
R333 VTAIL.n144 VTAIL.n134 1.93989
R334 VTAIL.n112 VTAIL.n102 1.93989
R335 VTAIL.n239 VTAIL.n232 1.16414
R336 VTAIL.n15 VTAIL.n8 1.16414
R337 VTAIL.n47 VTAIL.n40 1.16414
R338 VTAIL.n79 VTAIL.n72 1.16414
R339 VTAIL.n207 VTAIL.n200 1.16414
R340 VTAIL.n175 VTAIL.n168 1.16414
R341 VTAIL.n143 VTAIL.n136 1.16414
R342 VTAIL.n111 VTAIL.n104 1.16414
R343 VTAIL.n159 VTAIL.n127 0.966017
R344 VTAIL.n223 VTAIL.n191 0.966017
R345 VTAIL.n95 VTAIL.n63 0.966017
R346 VTAIL VTAIL.n31 0.541448
R347 VTAIL.n191 VTAIL.n159 0.470328
R348 VTAIL.n63 VTAIL.n31 0.470328
R349 VTAIL VTAIL.n255 0.425069
R350 VTAIL.n236 VTAIL.n235 0.388379
R351 VTAIL.n12 VTAIL.n11 0.388379
R352 VTAIL.n44 VTAIL.n43 0.388379
R353 VTAIL.n76 VTAIL.n75 0.388379
R354 VTAIL.n204 VTAIL.n203 0.388379
R355 VTAIL.n172 VTAIL.n171 0.388379
R356 VTAIL.n140 VTAIL.n139 0.388379
R357 VTAIL.n108 VTAIL.n107 0.388379
R358 VTAIL.n238 VTAIL.n237 0.155672
R359 VTAIL.n238 VTAIL.n229 0.155672
R360 VTAIL.n245 VTAIL.n229 0.155672
R361 VTAIL.n246 VTAIL.n245 0.155672
R362 VTAIL.n246 VTAIL.n225 0.155672
R363 VTAIL.n253 VTAIL.n225 0.155672
R364 VTAIL.n14 VTAIL.n13 0.155672
R365 VTAIL.n14 VTAIL.n5 0.155672
R366 VTAIL.n21 VTAIL.n5 0.155672
R367 VTAIL.n22 VTAIL.n21 0.155672
R368 VTAIL.n22 VTAIL.n1 0.155672
R369 VTAIL.n29 VTAIL.n1 0.155672
R370 VTAIL.n46 VTAIL.n45 0.155672
R371 VTAIL.n46 VTAIL.n37 0.155672
R372 VTAIL.n53 VTAIL.n37 0.155672
R373 VTAIL.n54 VTAIL.n53 0.155672
R374 VTAIL.n54 VTAIL.n33 0.155672
R375 VTAIL.n61 VTAIL.n33 0.155672
R376 VTAIL.n78 VTAIL.n77 0.155672
R377 VTAIL.n78 VTAIL.n69 0.155672
R378 VTAIL.n85 VTAIL.n69 0.155672
R379 VTAIL.n86 VTAIL.n85 0.155672
R380 VTAIL.n86 VTAIL.n65 0.155672
R381 VTAIL.n93 VTAIL.n65 0.155672
R382 VTAIL.n221 VTAIL.n193 0.155672
R383 VTAIL.n214 VTAIL.n193 0.155672
R384 VTAIL.n214 VTAIL.n213 0.155672
R385 VTAIL.n213 VTAIL.n197 0.155672
R386 VTAIL.n206 VTAIL.n197 0.155672
R387 VTAIL.n206 VTAIL.n205 0.155672
R388 VTAIL.n189 VTAIL.n161 0.155672
R389 VTAIL.n182 VTAIL.n161 0.155672
R390 VTAIL.n182 VTAIL.n181 0.155672
R391 VTAIL.n181 VTAIL.n165 0.155672
R392 VTAIL.n174 VTAIL.n165 0.155672
R393 VTAIL.n174 VTAIL.n173 0.155672
R394 VTAIL.n157 VTAIL.n129 0.155672
R395 VTAIL.n150 VTAIL.n129 0.155672
R396 VTAIL.n150 VTAIL.n149 0.155672
R397 VTAIL.n149 VTAIL.n133 0.155672
R398 VTAIL.n142 VTAIL.n133 0.155672
R399 VTAIL.n142 VTAIL.n141 0.155672
R400 VTAIL.n125 VTAIL.n97 0.155672
R401 VTAIL.n118 VTAIL.n97 0.155672
R402 VTAIL.n118 VTAIL.n117 0.155672
R403 VTAIL.n117 VTAIL.n101 0.155672
R404 VTAIL.n110 VTAIL.n101 0.155672
R405 VTAIL.n110 VTAIL.n109 0.155672
R406 VDD1 VDD1.n1 124.805
R407 VDD1 VDD1.n0 92.5462
R408 VDD1.n0 VDD1.t1 5.40899
R409 VDD1.n0 VDD1.t0 5.40899
R410 VDD1.n1 VDD1.t2 5.40899
R411 VDD1.n1 VDD1.t3 5.40899
R412 VN.n0 VN.t2 254.37
R413 VN.n1 VN.t1 254.37
R414 VN.n0 VN.t3 254.321
R415 VN.n1 VN.t0 254.321
R416 VN VN.n1 81.2549
R417 VN VN.n0 44.7132
R418 VDD2.n2 VDD2.n0 124.281
R419 VDD2.n2 VDD2.n1 92.488
R420 VDD2.n1 VDD2.t3 5.40899
R421 VDD2.n1 VDD2.t2 5.40899
R422 VDD2.n0 VDD2.t1 5.40899
R423 VDD2.n0 VDD2.t0 5.40899
R424 VDD2 VDD2.n2 0.0586897
R425 B.n275 B.n44 585
R426 B.n277 B.n276 585
R427 B.n278 B.n43 585
R428 B.n280 B.n279 585
R429 B.n281 B.n42 585
R430 B.n283 B.n282 585
R431 B.n284 B.n41 585
R432 B.n286 B.n285 585
R433 B.n287 B.n40 585
R434 B.n289 B.n288 585
R435 B.n290 B.n39 585
R436 B.n292 B.n291 585
R437 B.n293 B.n38 585
R438 B.n295 B.n294 585
R439 B.n296 B.n37 585
R440 B.n298 B.n297 585
R441 B.n299 B.n36 585
R442 B.n301 B.n300 585
R443 B.n302 B.n35 585
R444 B.n304 B.n303 585
R445 B.n305 B.n34 585
R446 B.n307 B.n306 585
R447 B.n308 B.n33 585
R448 B.n310 B.n309 585
R449 B.n312 B.n311 585
R450 B.n313 B.n29 585
R451 B.n315 B.n314 585
R452 B.n316 B.n28 585
R453 B.n318 B.n317 585
R454 B.n319 B.n27 585
R455 B.n321 B.n320 585
R456 B.n322 B.n26 585
R457 B.n324 B.n323 585
R458 B.n325 B.n23 585
R459 B.n328 B.n327 585
R460 B.n329 B.n22 585
R461 B.n331 B.n330 585
R462 B.n332 B.n21 585
R463 B.n334 B.n333 585
R464 B.n335 B.n20 585
R465 B.n337 B.n336 585
R466 B.n338 B.n19 585
R467 B.n340 B.n339 585
R468 B.n341 B.n18 585
R469 B.n343 B.n342 585
R470 B.n344 B.n17 585
R471 B.n346 B.n345 585
R472 B.n347 B.n16 585
R473 B.n349 B.n348 585
R474 B.n350 B.n15 585
R475 B.n352 B.n351 585
R476 B.n353 B.n14 585
R477 B.n355 B.n354 585
R478 B.n356 B.n13 585
R479 B.n358 B.n357 585
R480 B.n359 B.n12 585
R481 B.n361 B.n360 585
R482 B.n362 B.n11 585
R483 B.n274 B.n273 585
R484 B.n272 B.n45 585
R485 B.n271 B.n270 585
R486 B.n269 B.n46 585
R487 B.n268 B.n267 585
R488 B.n266 B.n47 585
R489 B.n265 B.n264 585
R490 B.n263 B.n48 585
R491 B.n262 B.n261 585
R492 B.n260 B.n49 585
R493 B.n259 B.n258 585
R494 B.n257 B.n50 585
R495 B.n256 B.n255 585
R496 B.n254 B.n51 585
R497 B.n253 B.n252 585
R498 B.n251 B.n52 585
R499 B.n250 B.n249 585
R500 B.n248 B.n53 585
R501 B.n247 B.n246 585
R502 B.n245 B.n54 585
R503 B.n244 B.n243 585
R504 B.n242 B.n55 585
R505 B.n241 B.n240 585
R506 B.n239 B.n56 585
R507 B.n238 B.n237 585
R508 B.n236 B.n57 585
R509 B.n235 B.n234 585
R510 B.n233 B.n58 585
R511 B.n232 B.n231 585
R512 B.n230 B.n59 585
R513 B.n229 B.n228 585
R514 B.n227 B.n60 585
R515 B.n226 B.n225 585
R516 B.n224 B.n61 585
R517 B.n223 B.n222 585
R518 B.n221 B.n62 585
R519 B.n220 B.n219 585
R520 B.n131 B.n96 585
R521 B.n133 B.n132 585
R522 B.n134 B.n95 585
R523 B.n136 B.n135 585
R524 B.n137 B.n94 585
R525 B.n139 B.n138 585
R526 B.n140 B.n93 585
R527 B.n142 B.n141 585
R528 B.n143 B.n92 585
R529 B.n145 B.n144 585
R530 B.n146 B.n91 585
R531 B.n148 B.n147 585
R532 B.n149 B.n90 585
R533 B.n151 B.n150 585
R534 B.n152 B.n89 585
R535 B.n154 B.n153 585
R536 B.n155 B.n88 585
R537 B.n157 B.n156 585
R538 B.n158 B.n87 585
R539 B.n160 B.n159 585
R540 B.n161 B.n86 585
R541 B.n163 B.n162 585
R542 B.n164 B.n85 585
R543 B.n166 B.n165 585
R544 B.n168 B.n167 585
R545 B.n169 B.n81 585
R546 B.n171 B.n170 585
R547 B.n172 B.n80 585
R548 B.n174 B.n173 585
R549 B.n175 B.n79 585
R550 B.n177 B.n176 585
R551 B.n178 B.n78 585
R552 B.n180 B.n179 585
R553 B.n181 B.n75 585
R554 B.n184 B.n183 585
R555 B.n185 B.n74 585
R556 B.n187 B.n186 585
R557 B.n188 B.n73 585
R558 B.n190 B.n189 585
R559 B.n191 B.n72 585
R560 B.n193 B.n192 585
R561 B.n194 B.n71 585
R562 B.n196 B.n195 585
R563 B.n197 B.n70 585
R564 B.n199 B.n198 585
R565 B.n200 B.n69 585
R566 B.n202 B.n201 585
R567 B.n203 B.n68 585
R568 B.n205 B.n204 585
R569 B.n206 B.n67 585
R570 B.n208 B.n207 585
R571 B.n209 B.n66 585
R572 B.n211 B.n210 585
R573 B.n212 B.n65 585
R574 B.n214 B.n213 585
R575 B.n215 B.n64 585
R576 B.n217 B.n216 585
R577 B.n218 B.n63 585
R578 B.n130 B.n129 585
R579 B.n128 B.n97 585
R580 B.n127 B.n126 585
R581 B.n125 B.n98 585
R582 B.n124 B.n123 585
R583 B.n122 B.n99 585
R584 B.n121 B.n120 585
R585 B.n119 B.n100 585
R586 B.n118 B.n117 585
R587 B.n116 B.n101 585
R588 B.n115 B.n114 585
R589 B.n113 B.n102 585
R590 B.n112 B.n111 585
R591 B.n110 B.n103 585
R592 B.n109 B.n108 585
R593 B.n107 B.n104 585
R594 B.n106 B.n105 585
R595 B.n2 B.n0 585
R596 B.n389 B.n1 585
R597 B.n388 B.n387 585
R598 B.n386 B.n3 585
R599 B.n385 B.n384 585
R600 B.n383 B.n4 585
R601 B.n382 B.n381 585
R602 B.n380 B.n5 585
R603 B.n379 B.n378 585
R604 B.n377 B.n6 585
R605 B.n376 B.n375 585
R606 B.n374 B.n7 585
R607 B.n373 B.n372 585
R608 B.n371 B.n8 585
R609 B.n370 B.n369 585
R610 B.n368 B.n9 585
R611 B.n367 B.n366 585
R612 B.n365 B.n10 585
R613 B.n364 B.n363 585
R614 B.n391 B.n390 585
R615 B.n131 B.n130 463.671
R616 B.n364 B.n11 463.671
R617 B.n220 B.n63 463.671
R618 B.n275 B.n274 463.671
R619 B.n76 B.t3 385.327
R620 B.n82 B.t6 385.327
R621 B.n24 B.t9 385.327
R622 B.n30 B.t0 385.327
R623 B.n76 B.t5 290.108
R624 B.n30 B.t1 290.108
R625 B.n82 B.t8 290.108
R626 B.n24 B.t10 290.108
R627 B.n77 B.t4 268.387
R628 B.n31 B.t2 268.387
R629 B.n83 B.t7 268.387
R630 B.n25 B.t11 268.387
R631 B.n130 B.n97 163.367
R632 B.n126 B.n97 163.367
R633 B.n126 B.n125 163.367
R634 B.n125 B.n124 163.367
R635 B.n124 B.n99 163.367
R636 B.n120 B.n99 163.367
R637 B.n120 B.n119 163.367
R638 B.n119 B.n118 163.367
R639 B.n118 B.n101 163.367
R640 B.n114 B.n101 163.367
R641 B.n114 B.n113 163.367
R642 B.n113 B.n112 163.367
R643 B.n112 B.n103 163.367
R644 B.n108 B.n103 163.367
R645 B.n108 B.n107 163.367
R646 B.n107 B.n106 163.367
R647 B.n106 B.n2 163.367
R648 B.n390 B.n2 163.367
R649 B.n390 B.n389 163.367
R650 B.n389 B.n388 163.367
R651 B.n388 B.n3 163.367
R652 B.n384 B.n3 163.367
R653 B.n384 B.n383 163.367
R654 B.n383 B.n382 163.367
R655 B.n382 B.n5 163.367
R656 B.n378 B.n5 163.367
R657 B.n378 B.n377 163.367
R658 B.n377 B.n376 163.367
R659 B.n376 B.n7 163.367
R660 B.n372 B.n7 163.367
R661 B.n372 B.n371 163.367
R662 B.n371 B.n370 163.367
R663 B.n370 B.n9 163.367
R664 B.n366 B.n9 163.367
R665 B.n366 B.n365 163.367
R666 B.n365 B.n364 163.367
R667 B.n132 B.n131 163.367
R668 B.n132 B.n95 163.367
R669 B.n136 B.n95 163.367
R670 B.n137 B.n136 163.367
R671 B.n138 B.n137 163.367
R672 B.n138 B.n93 163.367
R673 B.n142 B.n93 163.367
R674 B.n143 B.n142 163.367
R675 B.n144 B.n143 163.367
R676 B.n144 B.n91 163.367
R677 B.n148 B.n91 163.367
R678 B.n149 B.n148 163.367
R679 B.n150 B.n149 163.367
R680 B.n150 B.n89 163.367
R681 B.n154 B.n89 163.367
R682 B.n155 B.n154 163.367
R683 B.n156 B.n155 163.367
R684 B.n156 B.n87 163.367
R685 B.n160 B.n87 163.367
R686 B.n161 B.n160 163.367
R687 B.n162 B.n161 163.367
R688 B.n162 B.n85 163.367
R689 B.n166 B.n85 163.367
R690 B.n167 B.n166 163.367
R691 B.n167 B.n81 163.367
R692 B.n171 B.n81 163.367
R693 B.n172 B.n171 163.367
R694 B.n173 B.n172 163.367
R695 B.n173 B.n79 163.367
R696 B.n177 B.n79 163.367
R697 B.n178 B.n177 163.367
R698 B.n179 B.n178 163.367
R699 B.n179 B.n75 163.367
R700 B.n184 B.n75 163.367
R701 B.n185 B.n184 163.367
R702 B.n186 B.n185 163.367
R703 B.n186 B.n73 163.367
R704 B.n190 B.n73 163.367
R705 B.n191 B.n190 163.367
R706 B.n192 B.n191 163.367
R707 B.n192 B.n71 163.367
R708 B.n196 B.n71 163.367
R709 B.n197 B.n196 163.367
R710 B.n198 B.n197 163.367
R711 B.n198 B.n69 163.367
R712 B.n202 B.n69 163.367
R713 B.n203 B.n202 163.367
R714 B.n204 B.n203 163.367
R715 B.n204 B.n67 163.367
R716 B.n208 B.n67 163.367
R717 B.n209 B.n208 163.367
R718 B.n210 B.n209 163.367
R719 B.n210 B.n65 163.367
R720 B.n214 B.n65 163.367
R721 B.n215 B.n214 163.367
R722 B.n216 B.n215 163.367
R723 B.n216 B.n63 163.367
R724 B.n221 B.n220 163.367
R725 B.n222 B.n221 163.367
R726 B.n222 B.n61 163.367
R727 B.n226 B.n61 163.367
R728 B.n227 B.n226 163.367
R729 B.n228 B.n227 163.367
R730 B.n228 B.n59 163.367
R731 B.n232 B.n59 163.367
R732 B.n233 B.n232 163.367
R733 B.n234 B.n233 163.367
R734 B.n234 B.n57 163.367
R735 B.n238 B.n57 163.367
R736 B.n239 B.n238 163.367
R737 B.n240 B.n239 163.367
R738 B.n240 B.n55 163.367
R739 B.n244 B.n55 163.367
R740 B.n245 B.n244 163.367
R741 B.n246 B.n245 163.367
R742 B.n246 B.n53 163.367
R743 B.n250 B.n53 163.367
R744 B.n251 B.n250 163.367
R745 B.n252 B.n251 163.367
R746 B.n252 B.n51 163.367
R747 B.n256 B.n51 163.367
R748 B.n257 B.n256 163.367
R749 B.n258 B.n257 163.367
R750 B.n258 B.n49 163.367
R751 B.n262 B.n49 163.367
R752 B.n263 B.n262 163.367
R753 B.n264 B.n263 163.367
R754 B.n264 B.n47 163.367
R755 B.n268 B.n47 163.367
R756 B.n269 B.n268 163.367
R757 B.n270 B.n269 163.367
R758 B.n270 B.n45 163.367
R759 B.n274 B.n45 163.367
R760 B.n360 B.n11 163.367
R761 B.n360 B.n359 163.367
R762 B.n359 B.n358 163.367
R763 B.n358 B.n13 163.367
R764 B.n354 B.n13 163.367
R765 B.n354 B.n353 163.367
R766 B.n353 B.n352 163.367
R767 B.n352 B.n15 163.367
R768 B.n348 B.n15 163.367
R769 B.n348 B.n347 163.367
R770 B.n347 B.n346 163.367
R771 B.n346 B.n17 163.367
R772 B.n342 B.n17 163.367
R773 B.n342 B.n341 163.367
R774 B.n341 B.n340 163.367
R775 B.n340 B.n19 163.367
R776 B.n336 B.n19 163.367
R777 B.n336 B.n335 163.367
R778 B.n335 B.n334 163.367
R779 B.n334 B.n21 163.367
R780 B.n330 B.n21 163.367
R781 B.n330 B.n329 163.367
R782 B.n329 B.n328 163.367
R783 B.n328 B.n23 163.367
R784 B.n323 B.n23 163.367
R785 B.n323 B.n322 163.367
R786 B.n322 B.n321 163.367
R787 B.n321 B.n27 163.367
R788 B.n317 B.n27 163.367
R789 B.n317 B.n316 163.367
R790 B.n316 B.n315 163.367
R791 B.n315 B.n29 163.367
R792 B.n311 B.n29 163.367
R793 B.n311 B.n310 163.367
R794 B.n310 B.n33 163.367
R795 B.n306 B.n33 163.367
R796 B.n306 B.n305 163.367
R797 B.n305 B.n304 163.367
R798 B.n304 B.n35 163.367
R799 B.n300 B.n35 163.367
R800 B.n300 B.n299 163.367
R801 B.n299 B.n298 163.367
R802 B.n298 B.n37 163.367
R803 B.n294 B.n37 163.367
R804 B.n294 B.n293 163.367
R805 B.n293 B.n292 163.367
R806 B.n292 B.n39 163.367
R807 B.n288 B.n39 163.367
R808 B.n288 B.n287 163.367
R809 B.n287 B.n286 163.367
R810 B.n286 B.n41 163.367
R811 B.n282 B.n41 163.367
R812 B.n282 B.n281 163.367
R813 B.n281 B.n280 163.367
R814 B.n280 B.n43 163.367
R815 B.n276 B.n43 163.367
R816 B.n276 B.n275 163.367
R817 B.n182 B.n77 59.5399
R818 B.n84 B.n83 59.5399
R819 B.n326 B.n25 59.5399
R820 B.n32 B.n31 59.5399
R821 B.n273 B.n44 30.1273
R822 B.n363 B.n362 30.1273
R823 B.n219 B.n218 30.1273
R824 B.n129 B.n96 30.1273
R825 B.n77 B.n76 21.7217
R826 B.n83 B.n82 21.7217
R827 B.n25 B.n24 21.7217
R828 B.n31 B.n30 21.7217
R829 B B.n391 18.0485
R830 B.n362 B.n361 10.6151
R831 B.n361 B.n12 10.6151
R832 B.n357 B.n12 10.6151
R833 B.n357 B.n356 10.6151
R834 B.n356 B.n355 10.6151
R835 B.n355 B.n14 10.6151
R836 B.n351 B.n14 10.6151
R837 B.n351 B.n350 10.6151
R838 B.n350 B.n349 10.6151
R839 B.n349 B.n16 10.6151
R840 B.n345 B.n16 10.6151
R841 B.n345 B.n344 10.6151
R842 B.n344 B.n343 10.6151
R843 B.n343 B.n18 10.6151
R844 B.n339 B.n18 10.6151
R845 B.n339 B.n338 10.6151
R846 B.n338 B.n337 10.6151
R847 B.n337 B.n20 10.6151
R848 B.n333 B.n20 10.6151
R849 B.n333 B.n332 10.6151
R850 B.n332 B.n331 10.6151
R851 B.n331 B.n22 10.6151
R852 B.n327 B.n22 10.6151
R853 B.n325 B.n324 10.6151
R854 B.n324 B.n26 10.6151
R855 B.n320 B.n26 10.6151
R856 B.n320 B.n319 10.6151
R857 B.n319 B.n318 10.6151
R858 B.n318 B.n28 10.6151
R859 B.n314 B.n28 10.6151
R860 B.n314 B.n313 10.6151
R861 B.n313 B.n312 10.6151
R862 B.n309 B.n308 10.6151
R863 B.n308 B.n307 10.6151
R864 B.n307 B.n34 10.6151
R865 B.n303 B.n34 10.6151
R866 B.n303 B.n302 10.6151
R867 B.n302 B.n301 10.6151
R868 B.n301 B.n36 10.6151
R869 B.n297 B.n36 10.6151
R870 B.n297 B.n296 10.6151
R871 B.n296 B.n295 10.6151
R872 B.n295 B.n38 10.6151
R873 B.n291 B.n38 10.6151
R874 B.n291 B.n290 10.6151
R875 B.n290 B.n289 10.6151
R876 B.n289 B.n40 10.6151
R877 B.n285 B.n40 10.6151
R878 B.n285 B.n284 10.6151
R879 B.n284 B.n283 10.6151
R880 B.n283 B.n42 10.6151
R881 B.n279 B.n42 10.6151
R882 B.n279 B.n278 10.6151
R883 B.n278 B.n277 10.6151
R884 B.n277 B.n44 10.6151
R885 B.n219 B.n62 10.6151
R886 B.n223 B.n62 10.6151
R887 B.n224 B.n223 10.6151
R888 B.n225 B.n224 10.6151
R889 B.n225 B.n60 10.6151
R890 B.n229 B.n60 10.6151
R891 B.n230 B.n229 10.6151
R892 B.n231 B.n230 10.6151
R893 B.n231 B.n58 10.6151
R894 B.n235 B.n58 10.6151
R895 B.n236 B.n235 10.6151
R896 B.n237 B.n236 10.6151
R897 B.n237 B.n56 10.6151
R898 B.n241 B.n56 10.6151
R899 B.n242 B.n241 10.6151
R900 B.n243 B.n242 10.6151
R901 B.n243 B.n54 10.6151
R902 B.n247 B.n54 10.6151
R903 B.n248 B.n247 10.6151
R904 B.n249 B.n248 10.6151
R905 B.n249 B.n52 10.6151
R906 B.n253 B.n52 10.6151
R907 B.n254 B.n253 10.6151
R908 B.n255 B.n254 10.6151
R909 B.n255 B.n50 10.6151
R910 B.n259 B.n50 10.6151
R911 B.n260 B.n259 10.6151
R912 B.n261 B.n260 10.6151
R913 B.n261 B.n48 10.6151
R914 B.n265 B.n48 10.6151
R915 B.n266 B.n265 10.6151
R916 B.n267 B.n266 10.6151
R917 B.n267 B.n46 10.6151
R918 B.n271 B.n46 10.6151
R919 B.n272 B.n271 10.6151
R920 B.n273 B.n272 10.6151
R921 B.n133 B.n96 10.6151
R922 B.n134 B.n133 10.6151
R923 B.n135 B.n134 10.6151
R924 B.n135 B.n94 10.6151
R925 B.n139 B.n94 10.6151
R926 B.n140 B.n139 10.6151
R927 B.n141 B.n140 10.6151
R928 B.n141 B.n92 10.6151
R929 B.n145 B.n92 10.6151
R930 B.n146 B.n145 10.6151
R931 B.n147 B.n146 10.6151
R932 B.n147 B.n90 10.6151
R933 B.n151 B.n90 10.6151
R934 B.n152 B.n151 10.6151
R935 B.n153 B.n152 10.6151
R936 B.n153 B.n88 10.6151
R937 B.n157 B.n88 10.6151
R938 B.n158 B.n157 10.6151
R939 B.n159 B.n158 10.6151
R940 B.n159 B.n86 10.6151
R941 B.n163 B.n86 10.6151
R942 B.n164 B.n163 10.6151
R943 B.n165 B.n164 10.6151
R944 B.n169 B.n168 10.6151
R945 B.n170 B.n169 10.6151
R946 B.n170 B.n80 10.6151
R947 B.n174 B.n80 10.6151
R948 B.n175 B.n174 10.6151
R949 B.n176 B.n175 10.6151
R950 B.n176 B.n78 10.6151
R951 B.n180 B.n78 10.6151
R952 B.n181 B.n180 10.6151
R953 B.n183 B.n74 10.6151
R954 B.n187 B.n74 10.6151
R955 B.n188 B.n187 10.6151
R956 B.n189 B.n188 10.6151
R957 B.n189 B.n72 10.6151
R958 B.n193 B.n72 10.6151
R959 B.n194 B.n193 10.6151
R960 B.n195 B.n194 10.6151
R961 B.n195 B.n70 10.6151
R962 B.n199 B.n70 10.6151
R963 B.n200 B.n199 10.6151
R964 B.n201 B.n200 10.6151
R965 B.n201 B.n68 10.6151
R966 B.n205 B.n68 10.6151
R967 B.n206 B.n205 10.6151
R968 B.n207 B.n206 10.6151
R969 B.n207 B.n66 10.6151
R970 B.n211 B.n66 10.6151
R971 B.n212 B.n211 10.6151
R972 B.n213 B.n212 10.6151
R973 B.n213 B.n64 10.6151
R974 B.n217 B.n64 10.6151
R975 B.n218 B.n217 10.6151
R976 B.n129 B.n128 10.6151
R977 B.n128 B.n127 10.6151
R978 B.n127 B.n98 10.6151
R979 B.n123 B.n98 10.6151
R980 B.n123 B.n122 10.6151
R981 B.n122 B.n121 10.6151
R982 B.n121 B.n100 10.6151
R983 B.n117 B.n100 10.6151
R984 B.n117 B.n116 10.6151
R985 B.n116 B.n115 10.6151
R986 B.n115 B.n102 10.6151
R987 B.n111 B.n102 10.6151
R988 B.n111 B.n110 10.6151
R989 B.n110 B.n109 10.6151
R990 B.n109 B.n104 10.6151
R991 B.n105 B.n104 10.6151
R992 B.n105 B.n0 10.6151
R993 B.n387 B.n1 10.6151
R994 B.n387 B.n386 10.6151
R995 B.n386 B.n385 10.6151
R996 B.n385 B.n4 10.6151
R997 B.n381 B.n4 10.6151
R998 B.n381 B.n380 10.6151
R999 B.n380 B.n379 10.6151
R1000 B.n379 B.n6 10.6151
R1001 B.n375 B.n6 10.6151
R1002 B.n375 B.n374 10.6151
R1003 B.n374 B.n373 10.6151
R1004 B.n373 B.n8 10.6151
R1005 B.n369 B.n8 10.6151
R1006 B.n369 B.n368 10.6151
R1007 B.n368 B.n367 10.6151
R1008 B.n367 B.n10 10.6151
R1009 B.n363 B.n10 10.6151
R1010 B.n327 B.n326 9.36635
R1011 B.n309 B.n32 9.36635
R1012 B.n165 B.n84 9.36635
R1013 B.n183 B.n182 9.36635
R1014 B.n391 B.n0 2.81026
R1015 B.n391 B.n1 2.81026
R1016 B.n326 B.n325 1.24928
R1017 B.n312 B.n32 1.24928
R1018 B.n168 B.n84 1.24928
R1019 B.n182 B.n181 1.24928
C0 B VP 1.02585f
C1 VDD2 w_n1642_n2170# 0.936723f
C2 B VDD1 0.780788f
C3 VTAIL VP 1.74623f
C4 B VN 0.691584f
C5 VDD1 VTAIL 4.01805f
C6 VDD1 VP 1.94864f
C7 VN VTAIL 1.73213f
C8 VN VP 3.77667f
C9 VDD1 VN 0.147171f
C10 B VDD2 0.803598f
C11 B w_n1642_n2170# 5.34231f
C12 VDD2 VTAIL 4.06012f
C13 VDD2 VP 0.278939f
C14 VTAIL w_n1642_n2170# 2.59429f
C15 VP w_n1642_n2170# 2.53907f
C16 VDD2 VDD1 0.587163f
C17 VDD2 VN 1.81715f
C18 VDD1 w_n1642_n2170# 0.920381f
C19 VN w_n1642_n2170# 2.33256f
C20 B VTAIL 2.24194f
C21 VDD2 VSUBS 0.509316f
C22 VDD1 VSUBS 2.877959f
C23 VTAIL VSUBS 0.50763f
C24 VN VSUBS 3.88628f
C25 VP VSUBS 1.046312f
C26 B VSUBS 2.191598f
C27 w_n1642_n2170# VSUBS 44.4719f
C28 B.n0 VSUBS 0.00578f
C29 B.n1 VSUBS 0.00578f
C30 B.n2 VSUBS 0.009141f
C31 B.n3 VSUBS 0.009141f
C32 B.n4 VSUBS 0.009141f
C33 B.n5 VSUBS 0.009141f
C34 B.n6 VSUBS 0.009141f
C35 B.n7 VSUBS 0.009141f
C36 B.n8 VSUBS 0.009141f
C37 B.n9 VSUBS 0.009141f
C38 B.n10 VSUBS 0.009141f
C39 B.n11 VSUBS 0.021056f
C40 B.n12 VSUBS 0.009141f
C41 B.n13 VSUBS 0.009141f
C42 B.n14 VSUBS 0.009141f
C43 B.n15 VSUBS 0.009141f
C44 B.n16 VSUBS 0.009141f
C45 B.n17 VSUBS 0.009141f
C46 B.n18 VSUBS 0.009141f
C47 B.n19 VSUBS 0.009141f
C48 B.n20 VSUBS 0.009141f
C49 B.n21 VSUBS 0.009141f
C50 B.n22 VSUBS 0.009141f
C51 B.n23 VSUBS 0.009141f
C52 B.t11 VSUBS 0.11713f
C53 B.t10 VSUBS 0.130732f
C54 B.t9 VSUBS 0.270821f
C55 B.n24 VSUBS 0.227852f
C56 B.n25 VSUBS 0.194707f
C57 B.n26 VSUBS 0.009141f
C58 B.n27 VSUBS 0.009141f
C59 B.n28 VSUBS 0.009141f
C60 B.n29 VSUBS 0.009141f
C61 B.t2 VSUBS 0.117132f
C62 B.t1 VSUBS 0.130734f
C63 B.t0 VSUBS 0.270821f
C64 B.n30 VSUBS 0.22785f
C65 B.n31 VSUBS 0.194705f
C66 B.n32 VSUBS 0.021179f
C67 B.n33 VSUBS 0.009141f
C68 B.n34 VSUBS 0.009141f
C69 B.n35 VSUBS 0.009141f
C70 B.n36 VSUBS 0.009141f
C71 B.n37 VSUBS 0.009141f
C72 B.n38 VSUBS 0.009141f
C73 B.n39 VSUBS 0.009141f
C74 B.n40 VSUBS 0.009141f
C75 B.n41 VSUBS 0.009141f
C76 B.n42 VSUBS 0.009141f
C77 B.n43 VSUBS 0.009141f
C78 B.n44 VSUBS 0.019885f
C79 B.n45 VSUBS 0.009141f
C80 B.n46 VSUBS 0.009141f
C81 B.n47 VSUBS 0.009141f
C82 B.n48 VSUBS 0.009141f
C83 B.n49 VSUBS 0.009141f
C84 B.n50 VSUBS 0.009141f
C85 B.n51 VSUBS 0.009141f
C86 B.n52 VSUBS 0.009141f
C87 B.n53 VSUBS 0.009141f
C88 B.n54 VSUBS 0.009141f
C89 B.n55 VSUBS 0.009141f
C90 B.n56 VSUBS 0.009141f
C91 B.n57 VSUBS 0.009141f
C92 B.n58 VSUBS 0.009141f
C93 B.n59 VSUBS 0.009141f
C94 B.n60 VSUBS 0.009141f
C95 B.n61 VSUBS 0.009141f
C96 B.n62 VSUBS 0.009141f
C97 B.n63 VSUBS 0.021056f
C98 B.n64 VSUBS 0.009141f
C99 B.n65 VSUBS 0.009141f
C100 B.n66 VSUBS 0.009141f
C101 B.n67 VSUBS 0.009141f
C102 B.n68 VSUBS 0.009141f
C103 B.n69 VSUBS 0.009141f
C104 B.n70 VSUBS 0.009141f
C105 B.n71 VSUBS 0.009141f
C106 B.n72 VSUBS 0.009141f
C107 B.n73 VSUBS 0.009141f
C108 B.n74 VSUBS 0.009141f
C109 B.n75 VSUBS 0.009141f
C110 B.t4 VSUBS 0.117132f
C111 B.t5 VSUBS 0.130734f
C112 B.t3 VSUBS 0.270821f
C113 B.n76 VSUBS 0.22785f
C114 B.n77 VSUBS 0.194705f
C115 B.n78 VSUBS 0.009141f
C116 B.n79 VSUBS 0.009141f
C117 B.n80 VSUBS 0.009141f
C118 B.n81 VSUBS 0.009141f
C119 B.t7 VSUBS 0.11713f
C120 B.t8 VSUBS 0.130732f
C121 B.t6 VSUBS 0.270821f
C122 B.n82 VSUBS 0.227852f
C123 B.n83 VSUBS 0.194707f
C124 B.n84 VSUBS 0.021179f
C125 B.n85 VSUBS 0.009141f
C126 B.n86 VSUBS 0.009141f
C127 B.n87 VSUBS 0.009141f
C128 B.n88 VSUBS 0.009141f
C129 B.n89 VSUBS 0.009141f
C130 B.n90 VSUBS 0.009141f
C131 B.n91 VSUBS 0.009141f
C132 B.n92 VSUBS 0.009141f
C133 B.n93 VSUBS 0.009141f
C134 B.n94 VSUBS 0.009141f
C135 B.n95 VSUBS 0.009141f
C136 B.n96 VSUBS 0.021056f
C137 B.n97 VSUBS 0.009141f
C138 B.n98 VSUBS 0.009141f
C139 B.n99 VSUBS 0.009141f
C140 B.n100 VSUBS 0.009141f
C141 B.n101 VSUBS 0.009141f
C142 B.n102 VSUBS 0.009141f
C143 B.n103 VSUBS 0.009141f
C144 B.n104 VSUBS 0.009141f
C145 B.n105 VSUBS 0.009141f
C146 B.n106 VSUBS 0.009141f
C147 B.n107 VSUBS 0.009141f
C148 B.n108 VSUBS 0.009141f
C149 B.n109 VSUBS 0.009141f
C150 B.n110 VSUBS 0.009141f
C151 B.n111 VSUBS 0.009141f
C152 B.n112 VSUBS 0.009141f
C153 B.n113 VSUBS 0.009141f
C154 B.n114 VSUBS 0.009141f
C155 B.n115 VSUBS 0.009141f
C156 B.n116 VSUBS 0.009141f
C157 B.n117 VSUBS 0.009141f
C158 B.n118 VSUBS 0.009141f
C159 B.n119 VSUBS 0.009141f
C160 B.n120 VSUBS 0.009141f
C161 B.n121 VSUBS 0.009141f
C162 B.n122 VSUBS 0.009141f
C163 B.n123 VSUBS 0.009141f
C164 B.n124 VSUBS 0.009141f
C165 B.n125 VSUBS 0.009141f
C166 B.n126 VSUBS 0.009141f
C167 B.n127 VSUBS 0.009141f
C168 B.n128 VSUBS 0.009141f
C169 B.n129 VSUBS 0.019542f
C170 B.n130 VSUBS 0.019542f
C171 B.n131 VSUBS 0.021056f
C172 B.n132 VSUBS 0.009141f
C173 B.n133 VSUBS 0.009141f
C174 B.n134 VSUBS 0.009141f
C175 B.n135 VSUBS 0.009141f
C176 B.n136 VSUBS 0.009141f
C177 B.n137 VSUBS 0.009141f
C178 B.n138 VSUBS 0.009141f
C179 B.n139 VSUBS 0.009141f
C180 B.n140 VSUBS 0.009141f
C181 B.n141 VSUBS 0.009141f
C182 B.n142 VSUBS 0.009141f
C183 B.n143 VSUBS 0.009141f
C184 B.n144 VSUBS 0.009141f
C185 B.n145 VSUBS 0.009141f
C186 B.n146 VSUBS 0.009141f
C187 B.n147 VSUBS 0.009141f
C188 B.n148 VSUBS 0.009141f
C189 B.n149 VSUBS 0.009141f
C190 B.n150 VSUBS 0.009141f
C191 B.n151 VSUBS 0.009141f
C192 B.n152 VSUBS 0.009141f
C193 B.n153 VSUBS 0.009141f
C194 B.n154 VSUBS 0.009141f
C195 B.n155 VSUBS 0.009141f
C196 B.n156 VSUBS 0.009141f
C197 B.n157 VSUBS 0.009141f
C198 B.n158 VSUBS 0.009141f
C199 B.n159 VSUBS 0.009141f
C200 B.n160 VSUBS 0.009141f
C201 B.n161 VSUBS 0.009141f
C202 B.n162 VSUBS 0.009141f
C203 B.n163 VSUBS 0.009141f
C204 B.n164 VSUBS 0.009141f
C205 B.n165 VSUBS 0.008604f
C206 B.n166 VSUBS 0.009141f
C207 B.n167 VSUBS 0.009141f
C208 B.n168 VSUBS 0.005108f
C209 B.n169 VSUBS 0.009141f
C210 B.n170 VSUBS 0.009141f
C211 B.n171 VSUBS 0.009141f
C212 B.n172 VSUBS 0.009141f
C213 B.n173 VSUBS 0.009141f
C214 B.n174 VSUBS 0.009141f
C215 B.n175 VSUBS 0.009141f
C216 B.n176 VSUBS 0.009141f
C217 B.n177 VSUBS 0.009141f
C218 B.n178 VSUBS 0.009141f
C219 B.n179 VSUBS 0.009141f
C220 B.n180 VSUBS 0.009141f
C221 B.n181 VSUBS 0.005108f
C222 B.n182 VSUBS 0.021179f
C223 B.n183 VSUBS 0.008604f
C224 B.n184 VSUBS 0.009141f
C225 B.n185 VSUBS 0.009141f
C226 B.n186 VSUBS 0.009141f
C227 B.n187 VSUBS 0.009141f
C228 B.n188 VSUBS 0.009141f
C229 B.n189 VSUBS 0.009141f
C230 B.n190 VSUBS 0.009141f
C231 B.n191 VSUBS 0.009141f
C232 B.n192 VSUBS 0.009141f
C233 B.n193 VSUBS 0.009141f
C234 B.n194 VSUBS 0.009141f
C235 B.n195 VSUBS 0.009141f
C236 B.n196 VSUBS 0.009141f
C237 B.n197 VSUBS 0.009141f
C238 B.n198 VSUBS 0.009141f
C239 B.n199 VSUBS 0.009141f
C240 B.n200 VSUBS 0.009141f
C241 B.n201 VSUBS 0.009141f
C242 B.n202 VSUBS 0.009141f
C243 B.n203 VSUBS 0.009141f
C244 B.n204 VSUBS 0.009141f
C245 B.n205 VSUBS 0.009141f
C246 B.n206 VSUBS 0.009141f
C247 B.n207 VSUBS 0.009141f
C248 B.n208 VSUBS 0.009141f
C249 B.n209 VSUBS 0.009141f
C250 B.n210 VSUBS 0.009141f
C251 B.n211 VSUBS 0.009141f
C252 B.n212 VSUBS 0.009141f
C253 B.n213 VSUBS 0.009141f
C254 B.n214 VSUBS 0.009141f
C255 B.n215 VSUBS 0.009141f
C256 B.n216 VSUBS 0.009141f
C257 B.n217 VSUBS 0.009141f
C258 B.n218 VSUBS 0.021056f
C259 B.n219 VSUBS 0.019542f
C260 B.n220 VSUBS 0.019542f
C261 B.n221 VSUBS 0.009141f
C262 B.n222 VSUBS 0.009141f
C263 B.n223 VSUBS 0.009141f
C264 B.n224 VSUBS 0.009141f
C265 B.n225 VSUBS 0.009141f
C266 B.n226 VSUBS 0.009141f
C267 B.n227 VSUBS 0.009141f
C268 B.n228 VSUBS 0.009141f
C269 B.n229 VSUBS 0.009141f
C270 B.n230 VSUBS 0.009141f
C271 B.n231 VSUBS 0.009141f
C272 B.n232 VSUBS 0.009141f
C273 B.n233 VSUBS 0.009141f
C274 B.n234 VSUBS 0.009141f
C275 B.n235 VSUBS 0.009141f
C276 B.n236 VSUBS 0.009141f
C277 B.n237 VSUBS 0.009141f
C278 B.n238 VSUBS 0.009141f
C279 B.n239 VSUBS 0.009141f
C280 B.n240 VSUBS 0.009141f
C281 B.n241 VSUBS 0.009141f
C282 B.n242 VSUBS 0.009141f
C283 B.n243 VSUBS 0.009141f
C284 B.n244 VSUBS 0.009141f
C285 B.n245 VSUBS 0.009141f
C286 B.n246 VSUBS 0.009141f
C287 B.n247 VSUBS 0.009141f
C288 B.n248 VSUBS 0.009141f
C289 B.n249 VSUBS 0.009141f
C290 B.n250 VSUBS 0.009141f
C291 B.n251 VSUBS 0.009141f
C292 B.n252 VSUBS 0.009141f
C293 B.n253 VSUBS 0.009141f
C294 B.n254 VSUBS 0.009141f
C295 B.n255 VSUBS 0.009141f
C296 B.n256 VSUBS 0.009141f
C297 B.n257 VSUBS 0.009141f
C298 B.n258 VSUBS 0.009141f
C299 B.n259 VSUBS 0.009141f
C300 B.n260 VSUBS 0.009141f
C301 B.n261 VSUBS 0.009141f
C302 B.n262 VSUBS 0.009141f
C303 B.n263 VSUBS 0.009141f
C304 B.n264 VSUBS 0.009141f
C305 B.n265 VSUBS 0.009141f
C306 B.n266 VSUBS 0.009141f
C307 B.n267 VSUBS 0.009141f
C308 B.n268 VSUBS 0.009141f
C309 B.n269 VSUBS 0.009141f
C310 B.n270 VSUBS 0.009141f
C311 B.n271 VSUBS 0.009141f
C312 B.n272 VSUBS 0.009141f
C313 B.n273 VSUBS 0.020713f
C314 B.n274 VSUBS 0.019542f
C315 B.n275 VSUBS 0.021056f
C316 B.n276 VSUBS 0.009141f
C317 B.n277 VSUBS 0.009141f
C318 B.n278 VSUBS 0.009141f
C319 B.n279 VSUBS 0.009141f
C320 B.n280 VSUBS 0.009141f
C321 B.n281 VSUBS 0.009141f
C322 B.n282 VSUBS 0.009141f
C323 B.n283 VSUBS 0.009141f
C324 B.n284 VSUBS 0.009141f
C325 B.n285 VSUBS 0.009141f
C326 B.n286 VSUBS 0.009141f
C327 B.n287 VSUBS 0.009141f
C328 B.n288 VSUBS 0.009141f
C329 B.n289 VSUBS 0.009141f
C330 B.n290 VSUBS 0.009141f
C331 B.n291 VSUBS 0.009141f
C332 B.n292 VSUBS 0.009141f
C333 B.n293 VSUBS 0.009141f
C334 B.n294 VSUBS 0.009141f
C335 B.n295 VSUBS 0.009141f
C336 B.n296 VSUBS 0.009141f
C337 B.n297 VSUBS 0.009141f
C338 B.n298 VSUBS 0.009141f
C339 B.n299 VSUBS 0.009141f
C340 B.n300 VSUBS 0.009141f
C341 B.n301 VSUBS 0.009141f
C342 B.n302 VSUBS 0.009141f
C343 B.n303 VSUBS 0.009141f
C344 B.n304 VSUBS 0.009141f
C345 B.n305 VSUBS 0.009141f
C346 B.n306 VSUBS 0.009141f
C347 B.n307 VSUBS 0.009141f
C348 B.n308 VSUBS 0.009141f
C349 B.n309 VSUBS 0.008604f
C350 B.n310 VSUBS 0.009141f
C351 B.n311 VSUBS 0.009141f
C352 B.n312 VSUBS 0.005108f
C353 B.n313 VSUBS 0.009141f
C354 B.n314 VSUBS 0.009141f
C355 B.n315 VSUBS 0.009141f
C356 B.n316 VSUBS 0.009141f
C357 B.n317 VSUBS 0.009141f
C358 B.n318 VSUBS 0.009141f
C359 B.n319 VSUBS 0.009141f
C360 B.n320 VSUBS 0.009141f
C361 B.n321 VSUBS 0.009141f
C362 B.n322 VSUBS 0.009141f
C363 B.n323 VSUBS 0.009141f
C364 B.n324 VSUBS 0.009141f
C365 B.n325 VSUBS 0.005108f
C366 B.n326 VSUBS 0.021179f
C367 B.n327 VSUBS 0.008604f
C368 B.n328 VSUBS 0.009141f
C369 B.n329 VSUBS 0.009141f
C370 B.n330 VSUBS 0.009141f
C371 B.n331 VSUBS 0.009141f
C372 B.n332 VSUBS 0.009141f
C373 B.n333 VSUBS 0.009141f
C374 B.n334 VSUBS 0.009141f
C375 B.n335 VSUBS 0.009141f
C376 B.n336 VSUBS 0.009141f
C377 B.n337 VSUBS 0.009141f
C378 B.n338 VSUBS 0.009141f
C379 B.n339 VSUBS 0.009141f
C380 B.n340 VSUBS 0.009141f
C381 B.n341 VSUBS 0.009141f
C382 B.n342 VSUBS 0.009141f
C383 B.n343 VSUBS 0.009141f
C384 B.n344 VSUBS 0.009141f
C385 B.n345 VSUBS 0.009141f
C386 B.n346 VSUBS 0.009141f
C387 B.n347 VSUBS 0.009141f
C388 B.n348 VSUBS 0.009141f
C389 B.n349 VSUBS 0.009141f
C390 B.n350 VSUBS 0.009141f
C391 B.n351 VSUBS 0.009141f
C392 B.n352 VSUBS 0.009141f
C393 B.n353 VSUBS 0.009141f
C394 B.n354 VSUBS 0.009141f
C395 B.n355 VSUBS 0.009141f
C396 B.n356 VSUBS 0.009141f
C397 B.n357 VSUBS 0.009141f
C398 B.n358 VSUBS 0.009141f
C399 B.n359 VSUBS 0.009141f
C400 B.n360 VSUBS 0.009141f
C401 B.n361 VSUBS 0.009141f
C402 B.n362 VSUBS 0.021056f
C403 B.n363 VSUBS 0.019542f
C404 B.n364 VSUBS 0.019542f
C405 B.n365 VSUBS 0.009141f
C406 B.n366 VSUBS 0.009141f
C407 B.n367 VSUBS 0.009141f
C408 B.n368 VSUBS 0.009141f
C409 B.n369 VSUBS 0.009141f
C410 B.n370 VSUBS 0.009141f
C411 B.n371 VSUBS 0.009141f
C412 B.n372 VSUBS 0.009141f
C413 B.n373 VSUBS 0.009141f
C414 B.n374 VSUBS 0.009141f
C415 B.n375 VSUBS 0.009141f
C416 B.n376 VSUBS 0.009141f
C417 B.n377 VSUBS 0.009141f
C418 B.n378 VSUBS 0.009141f
C419 B.n379 VSUBS 0.009141f
C420 B.n380 VSUBS 0.009141f
C421 B.n381 VSUBS 0.009141f
C422 B.n382 VSUBS 0.009141f
C423 B.n383 VSUBS 0.009141f
C424 B.n384 VSUBS 0.009141f
C425 B.n385 VSUBS 0.009141f
C426 B.n386 VSUBS 0.009141f
C427 B.n387 VSUBS 0.009141f
C428 B.n388 VSUBS 0.009141f
C429 B.n389 VSUBS 0.009141f
C430 B.n390 VSUBS 0.009141f
C431 B.n391 VSUBS 0.020699f
C432 VDD2.t1 VSUBS 0.091389f
C433 VDD2.t0 VSUBS 0.091389f
C434 VDD2.n0 VSUBS 0.859809f
C435 VDD2.t3 VSUBS 0.091389f
C436 VDD2.t2 VSUBS 0.091389f
C437 VDD2.n1 VSUBS 0.605821f
C438 VDD2.n2 VSUBS 2.20481f
C439 VN.t2 VSUBS 0.57742f
C440 VN.t3 VSUBS 0.57736f
C441 VN.n0 VSUBS 0.472766f
C442 VN.t1 VSUBS 0.57742f
C443 VN.t0 VSUBS 0.57736f
C444 VN.n1 VSUBS 1.10354f
C445 VDD1.t1 VSUBS 0.087641f
C446 VDD1.t0 VSUBS 0.087641f
C447 VDD1.n0 VSUBS 0.581205f
C448 VDD1.t2 VSUBS 0.087641f
C449 VDD1.t3 VSUBS 0.087641f
C450 VDD1.n1 VSUBS 0.837333f
C451 VTAIL.n0 VSUBS 0.022179f
C452 VTAIL.n1 VSUBS 0.020184f
C453 VTAIL.n2 VSUBS 0.010846f
C454 VTAIL.n3 VSUBS 0.025636f
C455 VTAIL.n4 VSUBS 0.011484f
C456 VTAIL.n5 VSUBS 0.020184f
C457 VTAIL.n6 VSUBS 0.010846f
C458 VTAIL.n7 VSUBS 0.025636f
C459 VTAIL.n8 VSUBS 0.011484f
C460 VTAIL.n9 VSUBS 0.089313f
C461 VTAIL.t1 VSUBS 0.055019f
C462 VTAIL.n10 VSUBS 0.019227f
C463 VTAIL.n11 VSUBS 0.0163f
C464 VTAIL.n12 VSUBS 0.010846f
C465 VTAIL.n13 VSUBS 0.463897f
C466 VTAIL.n14 VSUBS 0.020184f
C467 VTAIL.n15 VSUBS 0.010846f
C468 VTAIL.n16 VSUBS 0.011484f
C469 VTAIL.n17 VSUBS 0.025636f
C470 VTAIL.n18 VSUBS 0.025636f
C471 VTAIL.n19 VSUBS 0.011484f
C472 VTAIL.n20 VSUBS 0.010846f
C473 VTAIL.n21 VSUBS 0.020184f
C474 VTAIL.n22 VSUBS 0.020184f
C475 VTAIL.n23 VSUBS 0.010846f
C476 VTAIL.n24 VSUBS 0.011484f
C477 VTAIL.n25 VSUBS 0.025636f
C478 VTAIL.n26 VSUBS 0.062065f
C479 VTAIL.n27 VSUBS 0.011484f
C480 VTAIL.n28 VSUBS 0.010846f
C481 VTAIL.n29 VSUBS 0.04693f
C482 VTAIL.n30 VSUBS 0.031221f
C483 VTAIL.n31 VSUBS 0.083131f
C484 VTAIL.n32 VSUBS 0.022179f
C485 VTAIL.n33 VSUBS 0.020184f
C486 VTAIL.n34 VSUBS 0.010846f
C487 VTAIL.n35 VSUBS 0.025636f
C488 VTAIL.n36 VSUBS 0.011484f
C489 VTAIL.n37 VSUBS 0.020184f
C490 VTAIL.n38 VSUBS 0.010846f
C491 VTAIL.n39 VSUBS 0.025636f
C492 VTAIL.n40 VSUBS 0.011484f
C493 VTAIL.n41 VSUBS 0.089313f
C494 VTAIL.t4 VSUBS 0.055019f
C495 VTAIL.n42 VSUBS 0.019227f
C496 VTAIL.n43 VSUBS 0.0163f
C497 VTAIL.n44 VSUBS 0.010846f
C498 VTAIL.n45 VSUBS 0.463897f
C499 VTAIL.n46 VSUBS 0.020184f
C500 VTAIL.n47 VSUBS 0.010846f
C501 VTAIL.n48 VSUBS 0.011484f
C502 VTAIL.n49 VSUBS 0.025636f
C503 VTAIL.n50 VSUBS 0.025636f
C504 VTAIL.n51 VSUBS 0.011484f
C505 VTAIL.n52 VSUBS 0.010846f
C506 VTAIL.n53 VSUBS 0.020184f
C507 VTAIL.n54 VSUBS 0.020184f
C508 VTAIL.n55 VSUBS 0.010846f
C509 VTAIL.n56 VSUBS 0.011484f
C510 VTAIL.n57 VSUBS 0.025636f
C511 VTAIL.n58 VSUBS 0.062065f
C512 VTAIL.n59 VSUBS 0.011484f
C513 VTAIL.n60 VSUBS 0.010846f
C514 VTAIL.n61 VSUBS 0.04693f
C515 VTAIL.n62 VSUBS 0.031221f
C516 VTAIL.n63 VSUBS 0.110744f
C517 VTAIL.n64 VSUBS 0.022179f
C518 VTAIL.n65 VSUBS 0.020184f
C519 VTAIL.n66 VSUBS 0.010846f
C520 VTAIL.n67 VSUBS 0.025636f
C521 VTAIL.n68 VSUBS 0.011484f
C522 VTAIL.n69 VSUBS 0.020184f
C523 VTAIL.n70 VSUBS 0.010846f
C524 VTAIL.n71 VSUBS 0.025636f
C525 VTAIL.n72 VSUBS 0.011484f
C526 VTAIL.n73 VSUBS 0.089313f
C527 VTAIL.t5 VSUBS 0.055019f
C528 VTAIL.n74 VSUBS 0.019227f
C529 VTAIL.n75 VSUBS 0.0163f
C530 VTAIL.n76 VSUBS 0.010846f
C531 VTAIL.n77 VSUBS 0.463897f
C532 VTAIL.n78 VSUBS 0.020184f
C533 VTAIL.n79 VSUBS 0.010846f
C534 VTAIL.n80 VSUBS 0.011484f
C535 VTAIL.n81 VSUBS 0.025636f
C536 VTAIL.n82 VSUBS 0.025636f
C537 VTAIL.n83 VSUBS 0.011484f
C538 VTAIL.n84 VSUBS 0.010846f
C539 VTAIL.n85 VSUBS 0.020184f
C540 VTAIL.n86 VSUBS 0.020184f
C541 VTAIL.n87 VSUBS 0.010846f
C542 VTAIL.n88 VSUBS 0.011484f
C543 VTAIL.n89 VSUBS 0.025636f
C544 VTAIL.n90 VSUBS 0.062065f
C545 VTAIL.n91 VSUBS 0.011484f
C546 VTAIL.n92 VSUBS 0.010846f
C547 VTAIL.n93 VSUBS 0.04693f
C548 VTAIL.n94 VSUBS 0.031221f
C549 VTAIL.n95 VSUBS 0.754112f
C550 VTAIL.n96 VSUBS 0.022179f
C551 VTAIL.n97 VSUBS 0.020184f
C552 VTAIL.n98 VSUBS 0.010846f
C553 VTAIL.n99 VSUBS 0.025636f
C554 VTAIL.n100 VSUBS 0.011484f
C555 VTAIL.n101 VSUBS 0.020184f
C556 VTAIL.n102 VSUBS 0.010846f
C557 VTAIL.n103 VSUBS 0.025636f
C558 VTAIL.n104 VSUBS 0.011484f
C559 VTAIL.n105 VSUBS 0.089313f
C560 VTAIL.t3 VSUBS 0.055019f
C561 VTAIL.n106 VSUBS 0.019227f
C562 VTAIL.n107 VSUBS 0.0163f
C563 VTAIL.n108 VSUBS 0.010846f
C564 VTAIL.n109 VSUBS 0.463897f
C565 VTAIL.n110 VSUBS 0.020184f
C566 VTAIL.n111 VSUBS 0.010846f
C567 VTAIL.n112 VSUBS 0.011484f
C568 VTAIL.n113 VSUBS 0.025636f
C569 VTAIL.n114 VSUBS 0.025636f
C570 VTAIL.n115 VSUBS 0.011484f
C571 VTAIL.n116 VSUBS 0.010846f
C572 VTAIL.n117 VSUBS 0.020184f
C573 VTAIL.n118 VSUBS 0.020184f
C574 VTAIL.n119 VSUBS 0.010846f
C575 VTAIL.n120 VSUBS 0.011484f
C576 VTAIL.n121 VSUBS 0.025636f
C577 VTAIL.n122 VSUBS 0.062065f
C578 VTAIL.n123 VSUBS 0.011484f
C579 VTAIL.n124 VSUBS 0.010846f
C580 VTAIL.n125 VSUBS 0.04693f
C581 VTAIL.n126 VSUBS 0.031221f
C582 VTAIL.n127 VSUBS 0.754112f
C583 VTAIL.n128 VSUBS 0.022179f
C584 VTAIL.n129 VSUBS 0.020184f
C585 VTAIL.n130 VSUBS 0.010846f
C586 VTAIL.n131 VSUBS 0.025636f
C587 VTAIL.n132 VSUBS 0.011484f
C588 VTAIL.n133 VSUBS 0.020184f
C589 VTAIL.n134 VSUBS 0.010846f
C590 VTAIL.n135 VSUBS 0.025636f
C591 VTAIL.n136 VSUBS 0.011484f
C592 VTAIL.n137 VSUBS 0.089313f
C593 VTAIL.t0 VSUBS 0.055019f
C594 VTAIL.n138 VSUBS 0.019227f
C595 VTAIL.n139 VSUBS 0.0163f
C596 VTAIL.n140 VSUBS 0.010846f
C597 VTAIL.n141 VSUBS 0.463897f
C598 VTAIL.n142 VSUBS 0.020184f
C599 VTAIL.n143 VSUBS 0.010846f
C600 VTAIL.n144 VSUBS 0.011484f
C601 VTAIL.n145 VSUBS 0.025636f
C602 VTAIL.n146 VSUBS 0.025636f
C603 VTAIL.n147 VSUBS 0.011484f
C604 VTAIL.n148 VSUBS 0.010846f
C605 VTAIL.n149 VSUBS 0.020184f
C606 VTAIL.n150 VSUBS 0.020184f
C607 VTAIL.n151 VSUBS 0.010846f
C608 VTAIL.n152 VSUBS 0.011484f
C609 VTAIL.n153 VSUBS 0.025636f
C610 VTAIL.n154 VSUBS 0.062065f
C611 VTAIL.n155 VSUBS 0.011484f
C612 VTAIL.n156 VSUBS 0.010846f
C613 VTAIL.n157 VSUBS 0.04693f
C614 VTAIL.n158 VSUBS 0.031221f
C615 VTAIL.n159 VSUBS 0.110744f
C616 VTAIL.n160 VSUBS 0.022179f
C617 VTAIL.n161 VSUBS 0.020184f
C618 VTAIL.n162 VSUBS 0.010846f
C619 VTAIL.n163 VSUBS 0.025636f
C620 VTAIL.n164 VSUBS 0.011484f
C621 VTAIL.n165 VSUBS 0.020184f
C622 VTAIL.n166 VSUBS 0.010846f
C623 VTAIL.n167 VSUBS 0.025636f
C624 VTAIL.n168 VSUBS 0.011484f
C625 VTAIL.n169 VSUBS 0.089313f
C626 VTAIL.t7 VSUBS 0.055019f
C627 VTAIL.n170 VSUBS 0.019227f
C628 VTAIL.n171 VSUBS 0.0163f
C629 VTAIL.n172 VSUBS 0.010846f
C630 VTAIL.n173 VSUBS 0.463897f
C631 VTAIL.n174 VSUBS 0.020184f
C632 VTAIL.n175 VSUBS 0.010846f
C633 VTAIL.n176 VSUBS 0.011484f
C634 VTAIL.n177 VSUBS 0.025636f
C635 VTAIL.n178 VSUBS 0.025636f
C636 VTAIL.n179 VSUBS 0.011484f
C637 VTAIL.n180 VSUBS 0.010846f
C638 VTAIL.n181 VSUBS 0.020184f
C639 VTAIL.n182 VSUBS 0.020184f
C640 VTAIL.n183 VSUBS 0.010846f
C641 VTAIL.n184 VSUBS 0.011484f
C642 VTAIL.n185 VSUBS 0.025636f
C643 VTAIL.n186 VSUBS 0.062065f
C644 VTAIL.n187 VSUBS 0.011484f
C645 VTAIL.n188 VSUBS 0.010846f
C646 VTAIL.n189 VSUBS 0.04693f
C647 VTAIL.n190 VSUBS 0.031221f
C648 VTAIL.n191 VSUBS 0.110744f
C649 VTAIL.n192 VSUBS 0.022179f
C650 VTAIL.n193 VSUBS 0.020184f
C651 VTAIL.n194 VSUBS 0.010846f
C652 VTAIL.n195 VSUBS 0.025636f
C653 VTAIL.n196 VSUBS 0.011484f
C654 VTAIL.n197 VSUBS 0.020184f
C655 VTAIL.n198 VSUBS 0.010846f
C656 VTAIL.n199 VSUBS 0.025636f
C657 VTAIL.n200 VSUBS 0.011484f
C658 VTAIL.n201 VSUBS 0.089313f
C659 VTAIL.t6 VSUBS 0.055019f
C660 VTAIL.n202 VSUBS 0.019227f
C661 VTAIL.n203 VSUBS 0.0163f
C662 VTAIL.n204 VSUBS 0.010846f
C663 VTAIL.n205 VSUBS 0.463897f
C664 VTAIL.n206 VSUBS 0.020184f
C665 VTAIL.n207 VSUBS 0.010846f
C666 VTAIL.n208 VSUBS 0.011484f
C667 VTAIL.n209 VSUBS 0.025636f
C668 VTAIL.n210 VSUBS 0.025636f
C669 VTAIL.n211 VSUBS 0.011484f
C670 VTAIL.n212 VSUBS 0.010846f
C671 VTAIL.n213 VSUBS 0.020184f
C672 VTAIL.n214 VSUBS 0.020184f
C673 VTAIL.n215 VSUBS 0.010846f
C674 VTAIL.n216 VSUBS 0.011484f
C675 VTAIL.n217 VSUBS 0.025636f
C676 VTAIL.n218 VSUBS 0.062065f
C677 VTAIL.n219 VSUBS 0.011484f
C678 VTAIL.n220 VSUBS 0.010846f
C679 VTAIL.n221 VSUBS 0.04693f
C680 VTAIL.n222 VSUBS 0.031221f
C681 VTAIL.n223 VSUBS 0.754112f
C682 VTAIL.n224 VSUBS 0.022179f
C683 VTAIL.n225 VSUBS 0.020184f
C684 VTAIL.n226 VSUBS 0.010846f
C685 VTAIL.n227 VSUBS 0.025636f
C686 VTAIL.n228 VSUBS 0.011484f
C687 VTAIL.n229 VSUBS 0.020184f
C688 VTAIL.n230 VSUBS 0.010846f
C689 VTAIL.n231 VSUBS 0.025636f
C690 VTAIL.n232 VSUBS 0.011484f
C691 VTAIL.n233 VSUBS 0.089313f
C692 VTAIL.t2 VSUBS 0.055019f
C693 VTAIL.n234 VSUBS 0.019227f
C694 VTAIL.n235 VSUBS 0.0163f
C695 VTAIL.n236 VSUBS 0.010846f
C696 VTAIL.n237 VSUBS 0.463897f
C697 VTAIL.n238 VSUBS 0.020184f
C698 VTAIL.n239 VSUBS 0.010846f
C699 VTAIL.n240 VSUBS 0.011484f
C700 VTAIL.n241 VSUBS 0.025636f
C701 VTAIL.n242 VSUBS 0.025636f
C702 VTAIL.n243 VSUBS 0.011484f
C703 VTAIL.n244 VSUBS 0.010846f
C704 VTAIL.n245 VSUBS 0.020184f
C705 VTAIL.n246 VSUBS 0.020184f
C706 VTAIL.n247 VSUBS 0.010846f
C707 VTAIL.n248 VSUBS 0.011484f
C708 VTAIL.n249 VSUBS 0.025636f
C709 VTAIL.n250 VSUBS 0.062065f
C710 VTAIL.n251 VSUBS 0.011484f
C711 VTAIL.n252 VSUBS 0.010846f
C712 VTAIL.n253 VSUBS 0.04693f
C713 VTAIL.n254 VSUBS 0.031221f
C714 VTAIL.n255 VSUBS 0.718931f
C715 VP.n0 VSUBS 0.042092f
C716 VP.t3 VSUBS 0.601891f
C717 VP.t2 VSUBS 0.601953f
C718 VP.n1 VSUBS 1.13415f
C719 VP.n2 VSUBS 2.17093f
C720 VP.t1 VSUBS 0.579946f
C721 VP.n3 VSUBS 0.263403f
C722 VP.n4 VSUBS 0.009551f
C723 VP.t0 VSUBS 0.579946f
C724 VP.n5 VSUBS 0.263403f
C725 VP.n6 VSUBS 0.032619f
.ends

