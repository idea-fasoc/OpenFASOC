* NGSPICE file created from diff_pair_sample_1044.ext - technology: sky130A

.subckt diff_pair_sample_1044 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=1.24
X1 B.t8 B.t6 B.t7 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=1.24
X2 VDD1.t7 VP.t0 VTAIL.t6 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=1.24
X3 VTAIL.t9 VP.t1 VDD1.t6 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=1.24
X4 VTAIL.t10 VP.t2 VDD1.t5 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=1.24
X5 VTAIL.t0 VN.t0 VDD2.t7 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=1.24
X6 VDD1.t4 VP.t3 VTAIL.t11 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
X7 B.t5 B.t3 B.t4 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=1.24
X8 VTAIL.t12 VP.t4 VDD1.t3 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
X9 VDD2.t6 VN.t1 VTAIL.t1 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=1.24
X10 VTAIL.t5 VN.t2 VDD2.t5 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
X11 VDD2.t4 VN.t3 VTAIL.t4 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
X12 VTAIL.t3 VN.t4 VDD2.t3 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0.396 ps=2.73 w=2.4 l=1.24
X13 VDD2.t2 VN.t5 VTAIL.t2 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
X14 B.t2 B.t0 B.t1 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.936 pd=5.58 as=0 ps=0 w=2.4 l=1.24
X15 VDD2.t1 VN.t6 VTAIL.t14 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=1.24
X16 VDD1.t2 VP.t5 VTAIL.t7 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.936 ps=5.58 w=2.4 l=1.24
X17 VDD1.t1 VP.t6 VTAIL.t8 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
X18 VTAIL.t15 VN.t7 VDD2.t0 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
X19 VTAIL.t13 VP.t7 VDD1.t0 w_n2540_n1448# sky130_fd_pr__pfet_01v8 ad=0.396 pd=2.73 as=0.396 ps=2.73 w=2.4 l=1.24
R0 B.n305 B.n304 585
R1 B.n306 B.n39 585
R2 B.n308 B.n307 585
R3 B.n309 B.n38 585
R4 B.n311 B.n310 585
R5 B.n312 B.n37 585
R6 B.n314 B.n313 585
R7 B.n315 B.n36 585
R8 B.n317 B.n316 585
R9 B.n318 B.n35 585
R10 B.n320 B.n319 585
R11 B.n321 B.n34 585
R12 B.n323 B.n322 585
R13 B.n325 B.n31 585
R14 B.n327 B.n326 585
R15 B.n328 B.n30 585
R16 B.n330 B.n329 585
R17 B.n331 B.n29 585
R18 B.n333 B.n332 585
R19 B.n334 B.n28 585
R20 B.n336 B.n335 585
R21 B.n337 B.n27 585
R22 B.n339 B.n338 585
R23 B.n341 B.n340 585
R24 B.n342 B.n23 585
R25 B.n344 B.n343 585
R26 B.n345 B.n22 585
R27 B.n347 B.n346 585
R28 B.n348 B.n21 585
R29 B.n350 B.n349 585
R30 B.n351 B.n20 585
R31 B.n353 B.n352 585
R32 B.n354 B.n19 585
R33 B.n356 B.n355 585
R34 B.n357 B.n18 585
R35 B.n359 B.n358 585
R36 B.n303 B.n40 585
R37 B.n302 B.n301 585
R38 B.n300 B.n41 585
R39 B.n299 B.n298 585
R40 B.n297 B.n42 585
R41 B.n296 B.n295 585
R42 B.n294 B.n43 585
R43 B.n293 B.n292 585
R44 B.n291 B.n44 585
R45 B.n290 B.n289 585
R46 B.n288 B.n45 585
R47 B.n287 B.n286 585
R48 B.n285 B.n46 585
R49 B.n284 B.n283 585
R50 B.n282 B.n47 585
R51 B.n281 B.n280 585
R52 B.n279 B.n48 585
R53 B.n278 B.n277 585
R54 B.n276 B.n49 585
R55 B.n275 B.n274 585
R56 B.n273 B.n50 585
R57 B.n272 B.n271 585
R58 B.n270 B.n51 585
R59 B.n269 B.n268 585
R60 B.n267 B.n52 585
R61 B.n266 B.n265 585
R62 B.n264 B.n53 585
R63 B.n263 B.n262 585
R64 B.n261 B.n54 585
R65 B.n260 B.n259 585
R66 B.n258 B.n55 585
R67 B.n257 B.n256 585
R68 B.n255 B.n56 585
R69 B.n254 B.n253 585
R70 B.n252 B.n57 585
R71 B.n251 B.n250 585
R72 B.n249 B.n58 585
R73 B.n248 B.n247 585
R74 B.n246 B.n59 585
R75 B.n245 B.n244 585
R76 B.n243 B.n60 585
R77 B.n242 B.n241 585
R78 B.n240 B.n61 585
R79 B.n239 B.n238 585
R80 B.n237 B.n62 585
R81 B.n236 B.n235 585
R82 B.n234 B.n63 585
R83 B.n233 B.n232 585
R84 B.n231 B.n64 585
R85 B.n230 B.n229 585
R86 B.n228 B.n65 585
R87 B.n227 B.n226 585
R88 B.n225 B.n66 585
R89 B.n224 B.n223 585
R90 B.n222 B.n67 585
R91 B.n221 B.n220 585
R92 B.n219 B.n68 585
R93 B.n218 B.n217 585
R94 B.n216 B.n69 585
R95 B.n215 B.n214 585
R96 B.n213 B.n70 585
R97 B.n212 B.n211 585
R98 B.n210 B.n71 585
R99 B.n155 B.n154 585
R100 B.n156 B.n93 585
R101 B.n158 B.n157 585
R102 B.n159 B.n92 585
R103 B.n161 B.n160 585
R104 B.n162 B.n91 585
R105 B.n164 B.n163 585
R106 B.n165 B.n90 585
R107 B.n167 B.n166 585
R108 B.n168 B.n89 585
R109 B.n170 B.n169 585
R110 B.n171 B.n88 585
R111 B.n173 B.n172 585
R112 B.n175 B.n85 585
R113 B.n177 B.n176 585
R114 B.n178 B.n84 585
R115 B.n180 B.n179 585
R116 B.n181 B.n83 585
R117 B.n183 B.n182 585
R118 B.n184 B.n82 585
R119 B.n186 B.n185 585
R120 B.n187 B.n81 585
R121 B.n189 B.n188 585
R122 B.n191 B.n190 585
R123 B.n192 B.n77 585
R124 B.n194 B.n193 585
R125 B.n195 B.n76 585
R126 B.n197 B.n196 585
R127 B.n198 B.n75 585
R128 B.n200 B.n199 585
R129 B.n201 B.n74 585
R130 B.n203 B.n202 585
R131 B.n204 B.n73 585
R132 B.n206 B.n205 585
R133 B.n207 B.n72 585
R134 B.n209 B.n208 585
R135 B.n153 B.n94 585
R136 B.n152 B.n151 585
R137 B.n150 B.n95 585
R138 B.n149 B.n148 585
R139 B.n147 B.n96 585
R140 B.n146 B.n145 585
R141 B.n144 B.n97 585
R142 B.n143 B.n142 585
R143 B.n141 B.n98 585
R144 B.n140 B.n139 585
R145 B.n138 B.n99 585
R146 B.n137 B.n136 585
R147 B.n135 B.n100 585
R148 B.n134 B.n133 585
R149 B.n132 B.n101 585
R150 B.n131 B.n130 585
R151 B.n129 B.n102 585
R152 B.n128 B.n127 585
R153 B.n126 B.n103 585
R154 B.n125 B.n124 585
R155 B.n123 B.n104 585
R156 B.n122 B.n121 585
R157 B.n120 B.n105 585
R158 B.n119 B.n118 585
R159 B.n117 B.n106 585
R160 B.n116 B.n115 585
R161 B.n114 B.n107 585
R162 B.n113 B.n112 585
R163 B.n111 B.n108 585
R164 B.n110 B.n109 585
R165 B.n2 B.n0 585
R166 B.n405 B.n1 585
R167 B.n404 B.n403 585
R168 B.n402 B.n3 585
R169 B.n401 B.n400 585
R170 B.n399 B.n4 585
R171 B.n398 B.n397 585
R172 B.n396 B.n5 585
R173 B.n395 B.n394 585
R174 B.n393 B.n6 585
R175 B.n392 B.n391 585
R176 B.n390 B.n7 585
R177 B.n389 B.n388 585
R178 B.n387 B.n8 585
R179 B.n386 B.n385 585
R180 B.n384 B.n9 585
R181 B.n383 B.n382 585
R182 B.n381 B.n10 585
R183 B.n380 B.n379 585
R184 B.n378 B.n11 585
R185 B.n377 B.n376 585
R186 B.n375 B.n12 585
R187 B.n374 B.n373 585
R188 B.n372 B.n13 585
R189 B.n371 B.n370 585
R190 B.n369 B.n14 585
R191 B.n368 B.n367 585
R192 B.n366 B.n15 585
R193 B.n365 B.n364 585
R194 B.n363 B.n16 585
R195 B.n362 B.n361 585
R196 B.n360 B.n17 585
R197 B.n407 B.n406 585
R198 B.n154 B.n153 559.769
R199 B.n358 B.n17 559.769
R200 B.n208 B.n71 559.769
R201 B.n304 B.n303 559.769
R202 B.n78 B.t5 252.761
R203 B.n32 B.t7 252.761
R204 B.n86 B.t2 252.761
R205 B.n24 B.t10 252.761
R206 B.n78 B.t3 250.965
R207 B.n86 B.t0 250.965
R208 B.n24 B.t9 250.965
R209 B.n32 B.t6 250.965
R210 B.n79 B.t4 222.311
R211 B.n33 B.t8 222.311
R212 B.n87 B.t1 222.311
R213 B.n25 B.t11 222.311
R214 B.n153 B.n152 163.367
R215 B.n152 B.n95 163.367
R216 B.n148 B.n95 163.367
R217 B.n148 B.n147 163.367
R218 B.n147 B.n146 163.367
R219 B.n146 B.n97 163.367
R220 B.n142 B.n97 163.367
R221 B.n142 B.n141 163.367
R222 B.n141 B.n140 163.367
R223 B.n140 B.n99 163.367
R224 B.n136 B.n99 163.367
R225 B.n136 B.n135 163.367
R226 B.n135 B.n134 163.367
R227 B.n134 B.n101 163.367
R228 B.n130 B.n101 163.367
R229 B.n130 B.n129 163.367
R230 B.n129 B.n128 163.367
R231 B.n128 B.n103 163.367
R232 B.n124 B.n103 163.367
R233 B.n124 B.n123 163.367
R234 B.n123 B.n122 163.367
R235 B.n122 B.n105 163.367
R236 B.n118 B.n105 163.367
R237 B.n118 B.n117 163.367
R238 B.n117 B.n116 163.367
R239 B.n116 B.n107 163.367
R240 B.n112 B.n107 163.367
R241 B.n112 B.n111 163.367
R242 B.n111 B.n110 163.367
R243 B.n110 B.n2 163.367
R244 B.n406 B.n2 163.367
R245 B.n406 B.n405 163.367
R246 B.n405 B.n404 163.367
R247 B.n404 B.n3 163.367
R248 B.n400 B.n3 163.367
R249 B.n400 B.n399 163.367
R250 B.n399 B.n398 163.367
R251 B.n398 B.n5 163.367
R252 B.n394 B.n5 163.367
R253 B.n394 B.n393 163.367
R254 B.n393 B.n392 163.367
R255 B.n392 B.n7 163.367
R256 B.n388 B.n7 163.367
R257 B.n388 B.n387 163.367
R258 B.n387 B.n386 163.367
R259 B.n386 B.n9 163.367
R260 B.n382 B.n9 163.367
R261 B.n382 B.n381 163.367
R262 B.n381 B.n380 163.367
R263 B.n380 B.n11 163.367
R264 B.n376 B.n11 163.367
R265 B.n376 B.n375 163.367
R266 B.n375 B.n374 163.367
R267 B.n374 B.n13 163.367
R268 B.n370 B.n13 163.367
R269 B.n370 B.n369 163.367
R270 B.n369 B.n368 163.367
R271 B.n368 B.n15 163.367
R272 B.n364 B.n15 163.367
R273 B.n364 B.n363 163.367
R274 B.n363 B.n362 163.367
R275 B.n362 B.n17 163.367
R276 B.n154 B.n93 163.367
R277 B.n158 B.n93 163.367
R278 B.n159 B.n158 163.367
R279 B.n160 B.n159 163.367
R280 B.n160 B.n91 163.367
R281 B.n164 B.n91 163.367
R282 B.n165 B.n164 163.367
R283 B.n166 B.n165 163.367
R284 B.n166 B.n89 163.367
R285 B.n170 B.n89 163.367
R286 B.n171 B.n170 163.367
R287 B.n172 B.n171 163.367
R288 B.n172 B.n85 163.367
R289 B.n177 B.n85 163.367
R290 B.n178 B.n177 163.367
R291 B.n179 B.n178 163.367
R292 B.n179 B.n83 163.367
R293 B.n183 B.n83 163.367
R294 B.n184 B.n183 163.367
R295 B.n185 B.n184 163.367
R296 B.n185 B.n81 163.367
R297 B.n189 B.n81 163.367
R298 B.n190 B.n189 163.367
R299 B.n190 B.n77 163.367
R300 B.n194 B.n77 163.367
R301 B.n195 B.n194 163.367
R302 B.n196 B.n195 163.367
R303 B.n196 B.n75 163.367
R304 B.n200 B.n75 163.367
R305 B.n201 B.n200 163.367
R306 B.n202 B.n201 163.367
R307 B.n202 B.n73 163.367
R308 B.n206 B.n73 163.367
R309 B.n207 B.n206 163.367
R310 B.n208 B.n207 163.367
R311 B.n212 B.n71 163.367
R312 B.n213 B.n212 163.367
R313 B.n214 B.n213 163.367
R314 B.n214 B.n69 163.367
R315 B.n218 B.n69 163.367
R316 B.n219 B.n218 163.367
R317 B.n220 B.n219 163.367
R318 B.n220 B.n67 163.367
R319 B.n224 B.n67 163.367
R320 B.n225 B.n224 163.367
R321 B.n226 B.n225 163.367
R322 B.n226 B.n65 163.367
R323 B.n230 B.n65 163.367
R324 B.n231 B.n230 163.367
R325 B.n232 B.n231 163.367
R326 B.n232 B.n63 163.367
R327 B.n236 B.n63 163.367
R328 B.n237 B.n236 163.367
R329 B.n238 B.n237 163.367
R330 B.n238 B.n61 163.367
R331 B.n242 B.n61 163.367
R332 B.n243 B.n242 163.367
R333 B.n244 B.n243 163.367
R334 B.n244 B.n59 163.367
R335 B.n248 B.n59 163.367
R336 B.n249 B.n248 163.367
R337 B.n250 B.n249 163.367
R338 B.n250 B.n57 163.367
R339 B.n254 B.n57 163.367
R340 B.n255 B.n254 163.367
R341 B.n256 B.n255 163.367
R342 B.n256 B.n55 163.367
R343 B.n260 B.n55 163.367
R344 B.n261 B.n260 163.367
R345 B.n262 B.n261 163.367
R346 B.n262 B.n53 163.367
R347 B.n266 B.n53 163.367
R348 B.n267 B.n266 163.367
R349 B.n268 B.n267 163.367
R350 B.n268 B.n51 163.367
R351 B.n272 B.n51 163.367
R352 B.n273 B.n272 163.367
R353 B.n274 B.n273 163.367
R354 B.n274 B.n49 163.367
R355 B.n278 B.n49 163.367
R356 B.n279 B.n278 163.367
R357 B.n280 B.n279 163.367
R358 B.n280 B.n47 163.367
R359 B.n284 B.n47 163.367
R360 B.n285 B.n284 163.367
R361 B.n286 B.n285 163.367
R362 B.n286 B.n45 163.367
R363 B.n290 B.n45 163.367
R364 B.n291 B.n290 163.367
R365 B.n292 B.n291 163.367
R366 B.n292 B.n43 163.367
R367 B.n296 B.n43 163.367
R368 B.n297 B.n296 163.367
R369 B.n298 B.n297 163.367
R370 B.n298 B.n41 163.367
R371 B.n302 B.n41 163.367
R372 B.n303 B.n302 163.367
R373 B.n358 B.n357 163.367
R374 B.n357 B.n356 163.367
R375 B.n356 B.n19 163.367
R376 B.n352 B.n19 163.367
R377 B.n352 B.n351 163.367
R378 B.n351 B.n350 163.367
R379 B.n350 B.n21 163.367
R380 B.n346 B.n21 163.367
R381 B.n346 B.n345 163.367
R382 B.n345 B.n344 163.367
R383 B.n344 B.n23 163.367
R384 B.n340 B.n23 163.367
R385 B.n340 B.n339 163.367
R386 B.n339 B.n27 163.367
R387 B.n335 B.n27 163.367
R388 B.n335 B.n334 163.367
R389 B.n334 B.n333 163.367
R390 B.n333 B.n29 163.367
R391 B.n329 B.n29 163.367
R392 B.n329 B.n328 163.367
R393 B.n328 B.n327 163.367
R394 B.n327 B.n31 163.367
R395 B.n322 B.n31 163.367
R396 B.n322 B.n321 163.367
R397 B.n321 B.n320 163.367
R398 B.n320 B.n35 163.367
R399 B.n316 B.n35 163.367
R400 B.n316 B.n315 163.367
R401 B.n315 B.n314 163.367
R402 B.n314 B.n37 163.367
R403 B.n310 B.n37 163.367
R404 B.n310 B.n309 163.367
R405 B.n309 B.n308 163.367
R406 B.n308 B.n39 163.367
R407 B.n304 B.n39 163.367
R408 B.n80 B.n79 59.5399
R409 B.n174 B.n87 59.5399
R410 B.n26 B.n25 59.5399
R411 B.n324 B.n33 59.5399
R412 B.n360 B.n359 36.3712
R413 B.n305 B.n40 36.3712
R414 B.n210 B.n209 36.3712
R415 B.n155 B.n94 36.3712
R416 B.n79 B.n78 30.449
R417 B.n87 B.n86 30.449
R418 B.n25 B.n24 30.449
R419 B.n33 B.n32 30.449
R420 B B.n407 18.0485
R421 B.n359 B.n18 10.6151
R422 B.n355 B.n18 10.6151
R423 B.n355 B.n354 10.6151
R424 B.n354 B.n353 10.6151
R425 B.n353 B.n20 10.6151
R426 B.n349 B.n20 10.6151
R427 B.n349 B.n348 10.6151
R428 B.n348 B.n347 10.6151
R429 B.n347 B.n22 10.6151
R430 B.n343 B.n22 10.6151
R431 B.n343 B.n342 10.6151
R432 B.n342 B.n341 10.6151
R433 B.n338 B.n337 10.6151
R434 B.n337 B.n336 10.6151
R435 B.n336 B.n28 10.6151
R436 B.n332 B.n28 10.6151
R437 B.n332 B.n331 10.6151
R438 B.n331 B.n330 10.6151
R439 B.n330 B.n30 10.6151
R440 B.n326 B.n30 10.6151
R441 B.n326 B.n325 10.6151
R442 B.n323 B.n34 10.6151
R443 B.n319 B.n34 10.6151
R444 B.n319 B.n318 10.6151
R445 B.n318 B.n317 10.6151
R446 B.n317 B.n36 10.6151
R447 B.n313 B.n36 10.6151
R448 B.n313 B.n312 10.6151
R449 B.n312 B.n311 10.6151
R450 B.n311 B.n38 10.6151
R451 B.n307 B.n38 10.6151
R452 B.n307 B.n306 10.6151
R453 B.n306 B.n305 10.6151
R454 B.n211 B.n210 10.6151
R455 B.n211 B.n70 10.6151
R456 B.n215 B.n70 10.6151
R457 B.n216 B.n215 10.6151
R458 B.n217 B.n216 10.6151
R459 B.n217 B.n68 10.6151
R460 B.n221 B.n68 10.6151
R461 B.n222 B.n221 10.6151
R462 B.n223 B.n222 10.6151
R463 B.n223 B.n66 10.6151
R464 B.n227 B.n66 10.6151
R465 B.n228 B.n227 10.6151
R466 B.n229 B.n228 10.6151
R467 B.n229 B.n64 10.6151
R468 B.n233 B.n64 10.6151
R469 B.n234 B.n233 10.6151
R470 B.n235 B.n234 10.6151
R471 B.n235 B.n62 10.6151
R472 B.n239 B.n62 10.6151
R473 B.n240 B.n239 10.6151
R474 B.n241 B.n240 10.6151
R475 B.n241 B.n60 10.6151
R476 B.n245 B.n60 10.6151
R477 B.n246 B.n245 10.6151
R478 B.n247 B.n246 10.6151
R479 B.n247 B.n58 10.6151
R480 B.n251 B.n58 10.6151
R481 B.n252 B.n251 10.6151
R482 B.n253 B.n252 10.6151
R483 B.n253 B.n56 10.6151
R484 B.n257 B.n56 10.6151
R485 B.n258 B.n257 10.6151
R486 B.n259 B.n258 10.6151
R487 B.n259 B.n54 10.6151
R488 B.n263 B.n54 10.6151
R489 B.n264 B.n263 10.6151
R490 B.n265 B.n264 10.6151
R491 B.n265 B.n52 10.6151
R492 B.n269 B.n52 10.6151
R493 B.n270 B.n269 10.6151
R494 B.n271 B.n270 10.6151
R495 B.n271 B.n50 10.6151
R496 B.n275 B.n50 10.6151
R497 B.n276 B.n275 10.6151
R498 B.n277 B.n276 10.6151
R499 B.n277 B.n48 10.6151
R500 B.n281 B.n48 10.6151
R501 B.n282 B.n281 10.6151
R502 B.n283 B.n282 10.6151
R503 B.n283 B.n46 10.6151
R504 B.n287 B.n46 10.6151
R505 B.n288 B.n287 10.6151
R506 B.n289 B.n288 10.6151
R507 B.n289 B.n44 10.6151
R508 B.n293 B.n44 10.6151
R509 B.n294 B.n293 10.6151
R510 B.n295 B.n294 10.6151
R511 B.n295 B.n42 10.6151
R512 B.n299 B.n42 10.6151
R513 B.n300 B.n299 10.6151
R514 B.n301 B.n300 10.6151
R515 B.n301 B.n40 10.6151
R516 B.n156 B.n155 10.6151
R517 B.n157 B.n156 10.6151
R518 B.n157 B.n92 10.6151
R519 B.n161 B.n92 10.6151
R520 B.n162 B.n161 10.6151
R521 B.n163 B.n162 10.6151
R522 B.n163 B.n90 10.6151
R523 B.n167 B.n90 10.6151
R524 B.n168 B.n167 10.6151
R525 B.n169 B.n168 10.6151
R526 B.n169 B.n88 10.6151
R527 B.n173 B.n88 10.6151
R528 B.n176 B.n175 10.6151
R529 B.n176 B.n84 10.6151
R530 B.n180 B.n84 10.6151
R531 B.n181 B.n180 10.6151
R532 B.n182 B.n181 10.6151
R533 B.n182 B.n82 10.6151
R534 B.n186 B.n82 10.6151
R535 B.n187 B.n186 10.6151
R536 B.n188 B.n187 10.6151
R537 B.n192 B.n191 10.6151
R538 B.n193 B.n192 10.6151
R539 B.n193 B.n76 10.6151
R540 B.n197 B.n76 10.6151
R541 B.n198 B.n197 10.6151
R542 B.n199 B.n198 10.6151
R543 B.n199 B.n74 10.6151
R544 B.n203 B.n74 10.6151
R545 B.n204 B.n203 10.6151
R546 B.n205 B.n204 10.6151
R547 B.n205 B.n72 10.6151
R548 B.n209 B.n72 10.6151
R549 B.n151 B.n94 10.6151
R550 B.n151 B.n150 10.6151
R551 B.n150 B.n149 10.6151
R552 B.n149 B.n96 10.6151
R553 B.n145 B.n96 10.6151
R554 B.n145 B.n144 10.6151
R555 B.n144 B.n143 10.6151
R556 B.n143 B.n98 10.6151
R557 B.n139 B.n98 10.6151
R558 B.n139 B.n138 10.6151
R559 B.n138 B.n137 10.6151
R560 B.n137 B.n100 10.6151
R561 B.n133 B.n100 10.6151
R562 B.n133 B.n132 10.6151
R563 B.n132 B.n131 10.6151
R564 B.n131 B.n102 10.6151
R565 B.n127 B.n102 10.6151
R566 B.n127 B.n126 10.6151
R567 B.n126 B.n125 10.6151
R568 B.n125 B.n104 10.6151
R569 B.n121 B.n104 10.6151
R570 B.n121 B.n120 10.6151
R571 B.n120 B.n119 10.6151
R572 B.n119 B.n106 10.6151
R573 B.n115 B.n106 10.6151
R574 B.n115 B.n114 10.6151
R575 B.n114 B.n113 10.6151
R576 B.n113 B.n108 10.6151
R577 B.n109 B.n108 10.6151
R578 B.n109 B.n0 10.6151
R579 B.n403 B.n1 10.6151
R580 B.n403 B.n402 10.6151
R581 B.n402 B.n401 10.6151
R582 B.n401 B.n4 10.6151
R583 B.n397 B.n4 10.6151
R584 B.n397 B.n396 10.6151
R585 B.n396 B.n395 10.6151
R586 B.n395 B.n6 10.6151
R587 B.n391 B.n6 10.6151
R588 B.n391 B.n390 10.6151
R589 B.n390 B.n389 10.6151
R590 B.n389 B.n8 10.6151
R591 B.n385 B.n8 10.6151
R592 B.n385 B.n384 10.6151
R593 B.n384 B.n383 10.6151
R594 B.n383 B.n10 10.6151
R595 B.n379 B.n10 10.6151
R596 B.n379 B.n378 10.6151
R597 B.n378 B.n377 10.6151
R598 B.n377 B.n12 10.6151
R599 B.n373 B.n12 10.6151
R600 B.n373 B.n372 10.6151
R601 B.n372 B.n371 10.6151
R602 B.n371 B.n14 10.6151
R603 B.n367 B.n14 10.6151
R604 B.n367 B.n366 10.6151
R605 B.n366 B.n365 10.6151
R606 B.n365 B.n16 10.6151
R607 B.n361 B.n16 10.6151
R608 B.n361 B.n360 10.6151
R609 B.n341 B.n26 9.36635
R610 B.n324 B.n323 9.36635
R611 B.n174 B.n173 9.36635
R612 B.n191 B.n80 9.36635
R613 B.n407 B.n0 2.81026
R614 B.n407 B.n1 2.81026
R615 B.n338 B.n26 1.24928
R616 B.n325 B.n324 1.24928
R617 B.n175 B.n174 1.24928
R618 B.n188 B.n80 1.24928
R619 VP.n11 VP.n10 161.3
R620 VP.n12 VP.n7 161.3
R621 VP.n14 VP.n13 161.3
R622 VP.n16 VP.n15 161.3
R623 VP.n17 VP.n5 161.3
R624 VP.n32 VP.n0 161.3
R625 VP.n31 VP.n30 161.3
R626 VP.n29 VP.n28 161.3
R627 VP.n27 VP.n2 161.3
R628 VP.n26 VP.n25 161.3
R629 VP.n24 VP.n23 161.3
R630 VP.n22 VP.n4 161.3
R631 VP.n9 VP.t2 98.0805
R632 VP.n19 VP.n18 80.6037
R633 VP.n34 VP.n33 80.6037
R634 VP.n21 VP.n20 80.6037
R635 VP.n21 VP.t1 78.3255
R636 VP.n33 VP.t0 78.3255
R637 VP.n18 VP.t5 78.3255
R638 VP.n3 VP.t3 46.6457
R639 VP.n1 VP.t7 46.6457
R640 VP.n6 VP.t4 46.6457
R641 VP.n8 VP.t6 46.6457
R642 VP.n9 VP.n8 43.6464
R643 VP.n27 VP.n26 40.577
R644 VP.n28 VP.n27 40.577
R645 VP.n13 VP.n12 40.577
R646 VP.n12 VP.n11 40.577
R647 VP.n20 VP.n19 37.4256
R648 VP.n22 VP.n21 34.3247
R649 VP.n33 VP.n32 34.3247
R650 VP.n18 VP.n17 34.3247
R651 VP.n23 VP.n22 33.7956
R652 VP.n32 VP.n31 33.7956
R653 VP.n17 VP.n16 33.7956
R654 VP.n10 VP.n9 29.3018
R655 VP.n26 VP.n3 14.0178
R656 VP.n28 VP.n1 14.0178
R657 VP.n13 VP.n6 14.0178
R658 VP.n11 VP.n8 14.0178
R659 VP.n23 VP.n3 10.575
R660 VP.n31 VP.n1 10.575
R661 VP.n16 VP.n6 10.575
R662 VP.n19 VP.n5 0.285035
R663 VP.n20 VP.n4 0.285035
R664 VP.n34 VP.n0 0.285035
R665 VP.n10 VP.n7 0.189894
R666 VP.n14 VP.n7 0.189894
R667 VP.n15 VP.n14 0.189894
R668 VP.n15 VP.n5 0.189894
R669 VP.n24 VP.n4 0.189894
R670 VP.n25 VP.n24 0.189894
R671 VP.n25 VP.n2 0.189894
R672 VP.n29 VP.n2 0.189894
R673 VP.n30 VP.n29 0.189894
R674 VP.n30 VP.n0 0.189894
R675 VP VP.n34 0.146778
R676 VTAIL.n98 VTAIL.n92 756.745
R677 VTAIL.n8 VTAIL.n2 756.745
R678 VTAIL.n20 VTAIL.n14 756.745
R679 VTAIL.n34 VTAIL.n28 756.745
R680 VTAIL.n86 VTAIL.n80 756.745
R681 VTAIL.n72 VTAIL.n66 756.745
R682 VTAIL.n60 VTAIL.n54 756.745
R683 VTAIL.n46 VTAIL.n40 756.745
R684 VTAIL.n97 VTAIL.n96 585
R685 VTAIL.n99 VTAIL.n98 585
R686 VTAIL.n7 VTAIL.n6 585
R687 VTAIL.n9 VTAIL.n8 585
R688 VTAIL.n19 VTAIL.n18 585
R689 VTAIL.n21 VTAIL.n20 585
R690 VTAIL.n33 VTAIL.n32 585
R691 VTAIL.n35 VTAIL.n34 585
R692 VTAIL.n87 VTAIL.n86 585
R693 VTAIL.n85 VTAIL.n84 585
R694 VTAIL.n73 VTAIL.n72 585
R695 VTAIL.n71 VTAIL.n70 585
R696 VTAIL.n61 VTAIL.n60 585
R697 VTAIL.n59 VTAIL.n58 585
R698 VTAIL.n47 VTAIL.n46 585
R699 VTAIL.n45 VTAIL.n44 585
R700 VTAIL.n95 VTAIL.t14 355.474
R701 VTAIL.n5 VTAIL.t3 355.474
R702 VTAIL.n17 VTAIL.t6 355.474
R703 VTAIL.n31 VTAIL.t9 355.474
R704 VTAIL.n83 VTAIL.t7 355.474
R705 VTAIL.n69 VTAIL.t10 355.474
R706 VTAIL.n57 VTAIL.t1 355.474
R707 VTAIL.n43 VTAIL.t0 355.474
R708 VTAIL.n98 VTAIL.n97 171.744
R709 VTAIL.n8 VTAIL.n7 171.744
R710 VTAIL.n20 VTAIL.n19 171.744
R711 VTAIL.n34 VTAIL.n33 171.744
R712 VTAIL.n86 VTAIL.n85 171.744
R713 VTAIL.n72 VTAIL.n71 171.744
R714 VTAIL.n60 VTAIL.n59 171.744
R715 VTAIL.n46 VTAIL.n45 171.744
R716 VTAIL.n79 VTAIL.n78 135.042
R717 VTAIL.n53 VTAIL.n52 135.042
R718 VTAIL.n1 VTAIL.n0 135.042
R719 VTAIL.n27 VTAIL.n26 135.042
R720 VTAIL.n97 VTAIL.t14 85.8723
R721 VTAIL.n7 VTAIL.t3 85.8723
R722 VTAIL.n19 VTAIL.t6 85.8723
R723 VTAIL.n33 VTAIL.t9 85.8723
R724 VTAIL.n85 VTAIL.t7 85.8723
R725 VTAIL.n71 VTAIL.t10 85.8723
R726 VTAIL.n59 VTAIL.t1 85.8723
R727 VTAIL.n45 VTAIL.t0 85.8723
R728 VTAIL.n103 VTAIL.n102 32.1853
R729 VTAIL.n13 VTAIL.n12 32.1853
R730 VTAIL.n25 VTAIL.n24 32.1853
R731 VTAIL.n39 VTAIL.n38 32.1853
R732 VTAIL.n91 VTAIL.n90 32.1853
R733 VTAIL.n77 VTAIL.n76 32.1853
R734 VTAIL.n65 VTAIL.n64 32.1853
R735 VTAIL.n51 VTAIL.n50 32.1853
R736 VTAIL.n96 VTAIL.n95 15.8418
R737 VTAIL.n6 VTAIL.n5 15.8418
R738 VTAIL.n18 VTAIL.n17 15.8418
R739 VTAIL.n32 VTAIL.n31 15.8418
R740 VTAIL.n84 VTAIL.n83 15.8418
R741 VTAIL.n70 VTAIL.n69 15.8418
R742 VTAIL.n58 VTAIL.n57 15.8418
R743 VTAIL.n44 VTAIL.n43 15.8418
R744 VTAIL.n103 VTAIL.n91 15.7893
R745 VTAIL.n51 VTAIL.n39 15.7893
R746 VTAIL.n0 VTAIL.t4 13.5442
R747 VTAIL.n0 VTAIL.t5 13.5442
R748 VTAIL.n26 VTAIL.t11 13.5442
R749 VTAIL.n26 VTAIL.t13 13.5442
R750 VTAIL.n78 VTAIL.t8 13.5442
R751 VTAIL.n78 VTAIL.t12 13.5442
R752 VTAIL.n52 VTAIL.t2 13.5442
R753 VTAIL.n52 VTAIL.t15 13.5442
R754 VTAIL.n99 VTAIL.n94 12.8005
R755 VTAIL.n9 VTAIL.n4 12.8005
R756 VTAIL.n21 VTAIL.n16 12.8005
R757 VTAIL.n35 VTAIL.n30 12.8005
R758 VTAIL.n87 VTAIL.n82 12.8005
R759 VTAIL.n73 VTAIL.n68 12.8005
R760 VTAIL.n61 VTAIL.n56 12.8005
R761 VTAIL.n47 VTAIL.n42 12.8005
R762 VTAIL.n100 VTAIL.n92 12.0247
R763 VTAIL.n10 VTAIL.n2 12.0247
R764 VTAIL.n22 VTAIL.n14 12.0247
R765 VTAIL.n36 VTAIL.n28 12.0247
R766 VTAIL.n88 VTAIL.n80 12.0247
R767 VTAIL.n74 VTAIL.n66 12.0247
R768 VTAIL.n62 VTAIL.n54 12.0247
R769 VTAIL.n48 VTAIL.n40 12.0247
R770 VTAIL.n102 VTAIL.n101 9.45567
R771 VTAIL.n12 VTAIL.n11 9.45567
R772 VTAIL.n24 VTAIL.n23 9.45567
R773 VTAIL.n38 VTAIL.n37 9.45567
R774 VTAIL.n90 VTAIL.n89 9.45567
R775 VTAIL.n76 VTAIL.n75 9.45567
R776 VTAIL.n64 VTAIL.n63 9.45567
R777 VTAIL.n50 VTAIL.n49 9.45567
R778 VTAIL.n101 VTAIL.n100 9.3005
R779 VTAIL.n94 VTAIL.n93 9.3005
R780 VTAIL.n11 VTAIL.n10 9.3005
R781 VTAIL.n4 VTAIL.n3 9.3005
R782 VTAIL.n23 VTAIL.n22 9.3005
R783 VTAIL.n16 VTAIL.n15 9.3005
R784 VTAIL.n37 VTAIL.n36 9.3005
R785 VTAIL.n30 VTAIL.n29 9.3005
R786 VTAIL.n89 VTAIL.n88 9.3005
R787 VTAIL.n82 VTAIL.n81 9.3005
R788 VTAIL.n75 VTAIL.n74 9.3005
R789 VTAIL.n68 VTAIL.n67 9.3005
R790 VTAIL.n63 VTAIL.n62 9.3005
R791 VTAIL.n56 VTAIL.n55 9.3005
R792 VTAIL.n49 VTAIL.n48 9.3005
R793 VTAIL.n42 VTAIL.n41 9.3005
R794 VTAIL.n83 VTAIL.n81 4.29255
R795 VTAIL.n69 VTAIL.n67 4.29255
R796 VTAIL.n57 VTAIL.n55 4.29255
R797 VTAIL.n43 VTAIL.n41 4.29255
R798 VTAIL.n95 VTAIL.n93 4.29255
R799 VTAIL.n5 VTAIL.n3 4.29255
R800 VTAIL.n17 VTAIL.n15 4.29255
R801 VTAIL.n31 VTAIL.n29 4.29255
R802 VTAIL.n102 VTAIL.n92 1.93989
R803 VTAIL.n12 VTAIL.n2 1.93989
R804 VTAIL.n24 VTAIL.n14 1.93989
R805 VTAIL.n38 VTAIL.n28 1.93989
R806 VTAIL.n90 VTAIL.n80 1.93989
R807 VTAIL.n76 VTAIL.n66 1.93989
R808 VTAIL.n64 VTAIL.n54 1.93989
R809 VTAIL.n50 VTAIL.n40 1.93989
R810 VTAIL.n53 VTAIL.n51 1.35395
R811 VTAIL.n65 VTAIL.n53 1.35395
R812 VTAIL.n79 VTAIL.n77 1.35395
R813 VTAIL.n91 VTAIL.n79 1.35395
R814 VTAIL.n39 VTAIL.n27 1.35395
R815 VTAIL.n27 VTAIL.n25 1.35395
R816 VTAIL.n13 VTAIL.n1 1.35395
R817 VTAIL VTAIL.n103 1.29576
R818 VTAIL.n100 VTAIL.n99 1.16414
R819 VTAIL.n10 VTAIL.n9 1.16414
R820 VTAIL.n22 VTAIL.n21 1.16414
R821 VTAIL.n36 VTAIL.n35 1.16414
R822 VTAIL.n88 VTAIL.n87 1.16414
R823 VTAIL.n74 VTAIL.n73 1.16414
R824 VTAIL.n62 VTAIL.n61 1.16414
R825 VTAIL.n48 VTAIL.n47 1.16414
R826 VTAIL.n77 VTAIL.n65 0.470328
R827 VTAIL.n25 VTAIL.n13 0.470328
R828 VTAIL.n96 VTAIL.n94 0.388379
R829 VTAIL.n6 VTAIL.n4 0.388379
R830 VTAIL.n18 VTAIL.n16 0.388379
R831 VTAIL.n32 VTAIL.n30 0.388379
R832 VTAIL.n84 VTAIL.n82 0.388379
R833 VTAIL.n70 VTAIL.n68 0.388379
R834 VTAIL.n58 VTAIL.n56 0.388379
R835 VTAIL.n44 VTAIL.n42 0.388379
R836 VTAIL.n101 VTAIL.n93 0.155672
R837 VTAIL.n11 VTAIL.n3 0.155672
R838 VTAIL.n23 VTAIL.n15 0.155672
R839 VTAIL.n37 VTAIL.n29 0.155672
R840 VTAIL.n89 VTAIL.n81 0.155672
R841 VTAIL.n75 VTAIL.n67 0.155672
R842 VTAIL.n63 VTAIL.n55 0.155672
R843 VTAIL.n49 VTAIL.n41 0.155672
R844 VTAIL VTAIL.n1 0.0586897
R845 VDD1 VDD1.n0 152.456
R846 VDD1.n3 VDD1.n2 152.341
R847 VDD1.n3 VDD1.n1 152.341
R848 VDD1.n5 VDD1.n4 151.72
R849 VDD1.n5 VDD1.n3 32.4578
R850 VDD1.n4 VDD1.t3 13.5442
R851 VDD1.n4 VDD1.t2 13.5442
R852 VDD1.n0 VDD1.t5 13.5442
R853 VDD1.n0 VDD1.t1 13.5442
R854 VDD1.n2 VDD1.t0 13.5442
R855 VDD1.n2 VDD1.t7 13.5442
R856 VDD1.n1 VDD1.t6 13.5442
R857 VDD1.n1 VDD1.t4 13.5442
R858 VDD1 VDD1.n5 0.619035
R859 VN.n27 VN.n15 161.3
R860 VN.n26 VN.n25 161.3
R861 VN.n24 VN.n23 161.3
R862 VN.n22 VN.n17 161.3
R863 VN.n21 VN.n20 161.3
R864 VN.n12 VN.n0 161.3
R865 VN.n11 VN.n10 161.3
R866 VN.n9 VN.n8 161.3
R867 VN.n7 VN.n2 161.3
R868 VN.n6 VN.n5 161.3
R869 VN.n4 VN.t4 98.0805
R870 VN.n19 VN.t1 98.0805
R871 VN.n29 VN.n28 80.6037
R872 VN.n14 VN.n13 80.6037
R873 VN.n13 VN.t6 78.3255
R874 VN.n28 VN.t0 78.3255
R875 VN.n3 VN.t3 46.6457
R876 VN.n1 VN.t2 46.6457
R877 VN.n18 VN.t7 46.6457
R878 VN.n16 VN.t5 46.6457
R879 VN.n4 VN.n3 43.6464
R880 VN.n19 VN.n18 43.6464
R881 VN.n7 VN.n6 40.577
R882 VN.n8 VN.n7 40.577
R883 VN.n22 VN.n21 40.577
R884 VN.n23 VN.n22 40.577
R885 VN VN.n29 37.7112
R886 VN.n13 VN.n12 34.3247
R887 VN.n28 VN.n27 34.3247
R888 VN.n12 VN.n11 33.7956
R889 VN.n27 VN.n26 33.7956
R890 VN.n20 VN.n19 29.3018
R891 VN.n5 VN.n4 29.3018
R892 VN.n6 VN.n3 14.0178
R893 VN.n8 VN.n1 14.0178
R894 VN.n21 VN.n18 14.0178
R895 VN.n23 VN.n16 14.0178
R896 VN.n11 VN.n1 10.575
R897 VN.n26 VN.n16 10.575
R898 VN.n29 VN.n15 0.285035
R899 VN.n14 VN.n0 0.285035
R900 VN.n25 VN.n15 0.189894
R901 VN.n25 VN.n24 0.189894
R902 VN.n24 VN.n17 0.189894
R903 VN.n20 VN.n17 0.189894
R904 VN.n5 VN.n2 0.189894
R905 VN.n9 VN.n2 0.189894
R906 VN.n10 VN.n9 0.189894
R907 VN.n10 VN.n0 0.189894
R908 VN VN.n14 0.146778
R909 VDD2.n2 VDD2.n1 152.341
R910 VDD2.n2 VDD2.n0 152.341
R911 VDD2 VDD2.n5 152.339
R912 VDD2.n4 VDD2.n3 151.72
R913 VDD2.n4 VDD2.n2 31.8748
R914 VDD2.n5 VDD2.t0 13.5442
R915 VDD2.n5 VDD2.t6 13.5442
R916 VDD2.n3 VDD2.t7 13.5442
R917 VDD2.n3 VDD2.t2 13.5442
R918 VDD2.n1 VDD2.t5 13.5442
R919 VDD2.n1 VDD2.t1 13.5442
R920 VDD2.n0 VDD2.t3 13.5442
R921 VDD2.n0 VDD2.t4 13.5442
R922 VDD2 VDD2.n4 0.735414
C0 B VP 1.33239f
C1 w_n2540_n1448# VDD2 1.29121f
C2 VP VN 4.2236f
C3 VTAIL VDD2 3.94813f
C4 w_n2540_n1448# VTAIL 1.81052f
C5 VDD1 VDD2 1.09481f
C6 B VDD2 1.02886f
C7 w_n2540_n1448# VDD1 1.23432f
C8 VN VDD2 1.75328f
C9 VTAIL VDD1 3.90283f
C10 B w_n2540_n1448# 5.3494f
C11 w_n2540_n1448# VN 4.59093f
C12 B VTAIL 1.38547f
C13 VTAIL VN 2.23811f
C14 VP VDD2 0.381168f
C15 B VDD1 0.97529f
C16 VDD1 VN 0.154751f
C17 w_n2540_n1448# VP 4.91324f
C18 B VN 0.794205f
C19 VTAIL VP 2.25221f
C20 VP VDD1 1.97817f
C21 VDD2 VSUBS 0.827411f
C22 VDD1 VSUBS 1.218283f
C23 VTAIL VSUBS 0.416741f
C24 VN VSUBS 4.50796f
C25 VP VSUBS 1.709877f
C26 B VSUBS 2.536203f
C27 w_n2540_n1448# VSUBS 46.7868f
C28 VDD2.t3 VSUBS 0.032225f
C29 VDD2.t4 VSUBS 0.032225f
C30 VDD2.n0 VSUBS 0.15728f
C31 VDD2.t5 VSUBS 0.032225f
C32 VDD2.t1 VSUBS 0.032225f
C33 VDD2.n1 VSUBS 0.15728f
C34 VDD2.n2 VSUBS 1.4123f
C35 VDD2.t7 VSUBS 0.032225f
C36 VDD2.t2 VSUBS 0.032225f
C37 VDD2.n3 VSUBS 0.156018f
C38 VDD2.n4 VSUBS 1.22054f
C39 VDD2.t0 VSUBS 0.032225f
C40 VDD2.t6 VSUBS 0.032225f
C41 VDD2.n5 VSUBS 0.157271f
C42 VN.n0 VSUBS 0.070285f
C43 VN.t2 VSUBS 0.378282f
C44 VN.n1 VSUBS 0.194652f
C45 VN.n2 VSUBS 0.052672f
C46 VN.t3 VSUBS 0.378282f
C47 VN.n3 VSUBS 0.264378f
C48 VN.t4 VSUBS 0.539833f
C49 VN.n4 VSUBS 0.282052f
C50 VN.n5 VSUBS 0.275477f
C51 VN.n6 VSUBS 0.0834f
C52 VN.n7 VSUBS 0.042542f
C53 VN.n8 VSUBS 0.0834f
C54 VN.n9 VSUBS 0.052672f
C55 VN.n10 VSUBS 0.052672f
C56 VN.n11 VSUBS 0.078332f
C57 VN.n12 VSUBS 0.036793f
C58 VN.t6 VSUBS 0.477734f
C59 VN.n13 VSUBS 0.296255f
C60 VN.n14 VSUBS 0.04933f
C61 VN.n15 VSUBS 0.070285f
C62 VN.t5 VSUBS 0.378282f
C63 VN.n16 VSUBS 0.194652f
C64 VN.n17 VSUBS 0.052672f
C65 VN.t7 VSUBS 0.378282f
C66 VN.n18 VSUBS 0.264378f
C67 VN.t1 VSUBS 0.539833f
C68 VN.n19 VSUBS 0.282052f
C69 VN.n20 VSUBS 0.275477f
C70 VN.n21 VSUBS 0.0834f
C71 VN.n22 VSUBS 0.042542f
C72 VN.n23 VSUBS 0.0834f
C73 VN.n24 VSUBS 0.052672f
C74 VN.n25 VSUBS 0.052672f
C75 VN.n26 VSUBS 0.078332f
C76 VN.n27 VSUBS 0.036793f
C77 VN.t0 VSUBS 0.477734f
C78 VN.n28 VSUBS 0.296255f
C79 VN.n29 VSUBS 1.82808f
C80 VDD1.t5 VSUBS 0.031715f
C81 VDD1.t1 VSUBS 0.031715f
C82 VDD1.n0 VSUBS 0.155042f
C83 VDD1.t6 VSUBS 0.031715f
C84 VDD1.t4 VSUBS 0.031715f
C85 VDD1.n1 VSUBS 0.154789f
C86 VDD1.t0 VSUBS 0.031715f
C87 VDD1.t7 VSUBS 0.031715f
C88 VDD1.n2 VSUBS 0.154789f
C89 VDD1.n3 VSUBS 1.42549f
C90 VDD1.t3 VSUBS 0.031715f
C91 VDD1.t2 VSUBS 0.031715f
C92 VDD1.n4 VSUBS 0.153547f
C93 VDD1.n5 VSUBS 1.22114f
C94 VTAIL.t4 VSUBS 0.050536f
C95 VTAIL.t5 VSUBS 0.050536f
C96 VTAIL.n0 VSUBS 0.207746f
C97 VTAIL.n1 VSUBS 0.425895f
C98 VTAIL.n2 VSUBS 0.026908f
C99 VTAIL.n3 VSUBS 0.179936f
C100 VTAIL.n4 VSUBS 0.014318f
C101 VTAIL.t3 VSUBS 0.07349f
C102 VTAIL.n5 VSUBS 0.085804f
C103 VTAIL.n6 VSUBS 0.019955f
C104 VTAIL.n7 VSUBS 0.025383f
C105 VTAIL.n8 VSUBS 0.073857f
C106 VTAIL.n9 VSUBS 0.015161f
C107 VTAIL.n10 VSUBS 0.014318f
C108 VTAIL.n11 VSUBS 0.061591f
C109 VTAIL.n12 VSUBS 0.036784f
C110 VTAIL.n13 VSUBS 0.179303f
C111 VTAIL.n14 VSUBS 0.026908f
C112 VTAIL.n15 VSUBS 0.179936f
C113 VTAIL.n16 VSUBS 0.014318f
C114 VTAIL.t6 VSUBS 0.07349f
C115 VTAIL.n17 VSUBS 0.085804f
C116 VTAIL.n18 VSUBS 0.019955f
C117 VTAIL.n19 VSUBS 0.025383f
C118 VTAIL.n20 VSUBS 0.073857f
C119 VTAIL.n21 VSUBS 0.015161f
C120 VTAIL.n22 VSUBS 0.014318f
C121 VTAIL.n23 VSUBS 0.061591f
C122 VTAIL.n24 VSUBS 0.036784f
C123 VTAIL.n25 VSUBS 0.179303f
C124 VTAIL.t11 VSUBS 0.050536f
C125 VTAIL.t13 VSUBS 0.050536f
C126 VTAIL.n26 VSUBS 0.207746f
C127 VTAIL.n27 VSUBS 0.537105f
C128 VTAIL.n28 VSUBS 0.026908f
C129 VTAIL.n29 VSUBS 0.179936f
C130 VTAIL.n30 VSUBS 0.014318f
C131 VTAIL.t9 VSUBS 0.07349f
C132 VTAIL.n31 VSUBS 0.085804f
C133 VTAIL.n32 VSUBS 0.019955f
C134 VTAIL.n33 VSUBS 0.025383f
C135 VTAIL.n34 VSUBS 0.073857f
C136 VTAIL.n35 VSUBS 0.015161f
C137 VTAIL.n36 VSUBS 0.014318f
C138 VTAIL.n37 VSUBS 0.061591f
C139 VTAIL.n38 VSUBS 0.036784f
C140 VTAIL.n39 VSUBS 0.794765f
C141 VTAIL.n40 VSUBS 0.026908f
C142 VTAIL.n41 VSUBS 0.179936f
C143 VTAIL.n42 VSUBS 0.014318f
C144 VTAIL.t0 VSUBS 0.07349f
C145 VTAIL.n43 VSUBS 0.085804f
C146 VTAIL.n44 VSUBS 0.019955f
C147 VTAIL.n45 VSUBS 0.025383f
C148 VTAIL.n46 VSUBS 0.073857f
C149 VTAIL.n47 VSUBS 0.015161f
C150 VTAIL.n48 VSUBS 0.014318f
C151 VTAIL.n49 VSUBS 0.061591f
C152 VTAIL.n50 VSUBS 0.036784f
C153 VTAIL.n51 VSUBS 0.794765f
C154 VTAIL.t2 VSUBS 0.050536f
C155 VTAIL.t15 VSUBS 0.050536f
C156 VTAIL.n52 VSUBS 0.207747f
C157 VTAIL.n53 VSUBS 0.537104f
C158 VTAIL.n54 VSUBS 0.026908f
C159 VTAIL.n55 VSUBS 0.179936f
C160 VTAIL.n56 VSUBS 0.014318f
C161 VTAIL.t1 VSUBS 0.07349f
C162 VTAIL.n57 VSUBS 0.085804f
C163 VTAIL.n58 VSUBS 0.019955f
C164 VTAIL.n59 VSUBS 0.025383f
C165 VTAIL.n60 VSUBS 0.073857f
C166 VTAIL.n61 VSUBS 0.015161f
C167 VTAIL.n62 VSUBS 0.014318f
C168 VTAIL.n63 VSUBS 0.061591f
C169 VTAIL.n64 VSUBS 0.036784f
C170 VTAIL.n65 VSUBS 0.179303f
C171 VTAIL.n66 VSUBS 0.026908f
C172 VTAIL.n67 VSUBS 0.179936f
C173 VTAIL.n68 VSUBS 0.014318f
C174 VTAIL.t10 VSUBS 0.07349f
C175 VTAIL.n69 VSUBS 0.085804f
C176 VTAIL.n70 VSUBS 0.019955f
C177 VTAIL.n71 VSUBS 0.025383f
C178 VTAIL.n72 VSUBS 0.073857f
C179 VTAIL.n73 VSUBS 0.015161f
C180 VTAIL.n74 VSUBS 0.014318f
C181 VTAIL.n75 VSUBS 0.061591f
C182 VTAIL.n76 VSUBS 0.036784f
C183 VTAIL.n77 VSUBS 0.179303f
C184 VTAIL.t8 VSUBS 0.050536f
C185 VTAIL.t12 VSUBS 0.050536f
C186 VTAIL.n78 VSUBS 0.207747f
C187 VTAIL.n79 VSUBS 0.537104f
C188 VTAIL.n80 VSUBS 0.026908f
C189 VTAIL.n81 VSUBS 0.179936f
C190 VTAIL.n82 VSUBS 0.014318f
C191 VTAIL.t7 VSUBS 0.07349f
C192 VTAIL.n83 VSUBS 0.085804f
C193 VTAIL.n84 VSUBS 0.019955f
C194 VTAIL.n85 VSUBS 0.025383f
C195 VTAIL.n86 VSUBS 0.073857f
C196 VTAIL.n87 VSUBS 0.015161f
C197 VTAIL.n88 VSUBS 0.014318f
C198 VTAIL.n89 VSUBS 0.061591f
C199 VTAIL.n90 VSUBS 0.036784f
C200 VTAIL.n91 VSUBS 0.794765f
C201 VTAIL.n92 VSUBS 0.026908f
C202 VTAIL.n93 VSUBS 0.179936f
C203 VTAIL.n94 VSUBS 0.014318f
C204 VTAIL.t14 VSUBS 0.07349f
C205 VTAIL.n95 VSUBS 0.085804f
C206 VTAIL.n96 VSUBS 0.019955f
C207 VTAIL.n97 VSUBS 0.025383f
C208 VTAIL.n98 VSUBS 0.073857f
C209 VTAIL.n99 VSUBS 0.015161f
C210 VTAIL.n100 VSUBS 0.014318f
C211 VTAIL.n101 VSUBS 0.061591f
C212 VTAIL.n102 VSUBS 0.036784f
C213 VTAIL.n103 VSUBS 0.789769f
C214 VP.n0 VSUBS 0.073334f
C215 VP.t7 VSUBS 0.394695f
C216 VP.n1 VSUBS 0.203097f
C217 VP.n2 VSUBS 0.054958f
C218 VP.t3 VSUBS 0.394695f
C219 VP.n3 VSUBS 0.203097f
C220 VP.n4 VSUBS 0.073334f
C221 VP.n5 VSUBS 0.073334f
C222 VP.t5 VSUBS 0.498461f
C223 VP.t4 VSUBS 0.394695f
C224 VP.n6 VSUBS 0.203097f
C225 VP.n7 VSUBS 0.054958f
C226 VP.t6 VSUBS 0.394695f
C227 VP.n8 VSUBS 0.275849f
C228 VP.t2 VSUBS 0.563255f
C229 VP.n9 VSUBS 0.294289f
C230 VP.n10 VSUBS 0.28743f
C231 VP.n11 VSUBS 0.087018f
C232 VP.n12 VSUBS 0.044387f
C233 VP.n13 VSUBS 0.087018f
C234 VP.n14 VSUBS 0.054958f
C235 VP.n15 VSUBS 0.054958f
C236 VP.n16 VSUBS 0.081731f
C237 VP.n17 VSUBS 0.038389f
C238 VP.n18 VSUBS 0.309109f
C239 VP.n19 VSUBS 1.8759f
C240 VP.n20 VSUBS 1.92884f
C241 VP.t1 VSUBS 0.498461f
C242 VP.n21 VSUBS 0.309109f
C243 VP.n22 VSUBS 0.038389f
C244 VP.n23 VSUBS 0.081731f
C245 VP.n24 VSUBS 0.054958f
C246 VP.n25 VSUBS 0.054958f
C247 VP.n26 VSUBS 0.087018f
C248 VP.n27 VSUBS 0.044387f
C249 VP.n28 VSUBS 0.087018f
C250 VP.n29 VSUBS 0.054958f
C251 VP.n30 VSUBS 0.054958f
C252 VP.n31 VSUBS 0.081731f
C253 VP.n32 VSUBS 0.038389f
C254 VP.t0 VSUBS 0.498461f
C255 VP.n33 VSUBS 0.309109f
C256 VP.n34 VSUBS 0.05147f
C257 B.n0 VSUBS 0.005193f
C258 B.n1 VSUBS 0.005193f
C259 B.n2 VSUBS 0.008212f
C260 B.n3 VSUBS 0.008212f
C261 B.n4 VSUBS 0.008212f
C262 B.n5 VSUBS 0.008212f
C263 B.n6 VSUBS 0.008212f
C264 B.n7 VSUBS 0.008212f
C265 B.n8 VSUBS 0.008212f
C266 B.n9 VSUBS 0.008212f
C267 B.n10 VSUBS 0.008212f
C268 B.n11 VSUBS 0.008212f
C269 B.n12 VSUBS 0.008212f
C270 B.n13 VSUBS 0.008212f
C271 B.n14 VSUBS 0.008212f
C272 B.n15 VSUBS 0.008212f
C273 B.n16 VSUBS 0.008212f
C274 B.n17 VSUBS 0.020215f
C275 B.n18 VSUBS 0.008212f
C276 B.n19 VSUBS 0.008212f
C277 B.n20 VSUBS 0.008212f
C278 B.n21 VSUBS 0.008212f
C279 B.n22 VSUBS 0.008212f
C280 B.n23 VSUBS 0.008212f
C281 B.t11 VSUBS 0.043493f
C282 B.t10 VSUBS 0.052407f
C283 B.t9 VSUBS 0.167443f
C284 B.n24 VSUBS 0.094626f
C285 B.n25 VSUBS 0.08571f
C286 B.n26 VSUBS 0.019026f
C287 B.n27 VSUBS 0.008212f
C288 B.n28 VSUBS 0.008212f
C289 B.n29 VSUBS 0.008212f
C290 B.n30 VSUBS 0.008212f
C291 B.n31 VSUBS 0.008212f
C292 B.t8 VSUBS 0.043493f
C293 B.t7 VSUBS 0.052407f
C294 B.t6 VSUBS 0.167443f
C295 B.n32 VSUBS 0.094626f
C296 B.n33 VSUBS 0.08571f
C297 B.n34 VSUBS 0.008212f
C298 B.n35 VSUBS 0.008212f
C299 B.n36 VSUBS 0.008212f
C300 B.n37 VSUBS 0.008212f
C301 B.n38 VSUBS 0.008212f
C302 B.n39 VSUBS 0.008212f
C303 B.n40 VSUBS 0.021086f
C304 B.n41 VSUBS 0.008212f
C305 B.n42 VSUBS 0.008212f
C306 B.n43 VSUBS 0.008212f
C307 B.n44 VSUBS 0.008212f
C308 B.n45 VSUBS 0.008212f
C309 B.n46 VSUBS 0.008212f
C310 B.n47 VSUBS 0.008212f
C311 B.n48 VSUBS 0.008212f
C312 B.n49 VSUBS 0.008212f
C313 B.n50 VSUBS 0.008212f
C314 B.n51 VSUBS 0.008212f
C315 B.n52 VSUBS 0.008212f
C316 B.n53 VSUBS 0.008212f
C317 B.n54 VSUBS 0.008212f
C318 B.n55 VSUBS 0.008212f
C319 B.n56 VSUBS 0.008212f
C320 B.n57 VSUBS 0.008212f
C321 B.n58 VSUBS 0.008212f
C322 B.n59 VSUBS 0.008212f
C323 B.n60 VSUBS 0.008212f
C324 B.n61 VSUBS 0.008212f
C325 B.n62 VSUBS 0.008212f
C326 B.n63 VSUBS 0.008212f
C327 B.n64 VSUBS 0.008212f
C328 B.n65 VSUBS 0.008212f
C329 B.n66 VSUBS 0.008212f
C330 B.n67 VSUBS 0.008212f
C331 B.n68 VSUBS 0.008212f
C332 B.n69 VSUBS 0.008212f
C333 B.n70 VSUBS 0.008212f
C334 B.n71 VSUBS 0.020215f
C335 B.n72 VSUBS 0.008212f
C336 B.n73 VSUBS 0.008212f
C337 B.n74 VSUBS 0.008212f
C338 B.n75 VSUBS 0.008212f
C339 B.n76 VSUBS 0.008212f
C340 B.n77 VSUBS 0.008212f
C341 B.t4 VSUBS 0.043493f
C342 B.t5 VSUBS 0.052407f
C343 B.t3 VSUBS 0.167443f
C344 B.n78 VSUBS 0.094626f
C345 B.n79 VSUBS 0.08571f
C346 B.n80 VSUBS 0.019026f
C347 B.n81 VSUBS 0.008212f
C348 B.n82 VSUBS 0.008212f
C349 B.n83 VSUBS 0.008212f
C350 B.n84 VSUBS 0.008212f
C351 B.n85 VSUBS 0.008212f
C352 B.t1 VSUBS 0.043493f
C353 B.t2 VSUBS 0.052407f
C354 B.t0 VSUBS 0.167443f
C355 B.n86 VSUBS 0.094626f
C356 B.n87 VSUBS 0.08571f
C357 B.n88 VSUBS 0.008212f
C358 B.n89 VSUBS 0.008212f
C359 B.n90 VSUBS 0.008212f
C360 B.n91 VSUBS 0.008212f
C361 B.n92 VSUBS 0.008212f
C362 B.n93 VSUBS 0.008212f
C363 B.n94 VSUBS 0.020215f
C364 B.n95 VSUBS 0.008212f
C365 B.n96 VSUBS 0.008212f
C366 B.n97 VSUBS 0.008212f
C367 B.n98 VSUBS 0.008212f
C368 B.n99 VSUBS 0.008212f
C369 B.n100 VSUBS 0.008212f
C370 B.n101 VSUBS 0.008212f
C371 B.n102 VSUBS 0.008212f
C372 B.n103 VSUBS 0.008212f
C373 B.n104 VSUBS 0.008212f
C374 B.n105 VSUBS 0.008212f
C375 B.n106 VSUBS 0.008212f
C376 B.n107 VSUBS 0.008212f
C377 B.n108 VSUBS 0.008212f
C378 B.n109 VSUBS 0.008212f
C379 B.n110 VSUBS 0.008212f
C380 B.n111 VSUBS 0.008212f
C381 B.n112 VSUBS 0.008212f
C382 B.n113 VSUBS 0.008212f
C383 B.n114 VSUBS 0.008212f
C384 B.n115 VSUBS 0.008212f
C385 B.n116 VSUBS 0.008212f
C386 B.n117 VSUBS 0.008212f
C387 B.n118 VSUBS 0.008212f
C388 B.n119 VSUBS 0.008212f
C389 B.n120 VSUBS 0.008212f
C390 B.n121 VSUBS 0.008212f
C391 B.n122 VSUBS 0.008212f
C392 B.n123 VSUBS 0.008212f
C393 B.n124 VSUBS 0.008212f
C394 B.n125 VSUBS 0.008212f
C395 B.n126 VSUBS 0.008212f
C396 B.n127 VSUBS 0.008212f
C397 B.n128 VSUBS 0.008212f
C398 B.n129 VSUBS 0.008212f
C399 B.n130 VSUBS 0.008212f
C400 B.n131 VSUBS 0.008212f
C401 B.n132 VSUBS 0.008212f
C402 B.n133 VSUBS 0.008212f
C403 B.n134 VSUBS 0.008212f
C404 B.n135 VSUBS 0.008212f
C405 B.n136 VSUBS 0.008212f
C406 B.n137 VSUBS 0.008212f
C407 B.n138 VSUBS 0.008212f
C408 B.n139 VSUBS 0.008212f
C409 B.n140 VSUBS 0.008212f
C410 B.n141 VSUBS 0.008212f
C411 B.n142 VSUBS 0.008212f
C412 B.n143 VSUBS 0.008212f
C413 B.n144 VSUBS 0.008212f
C414 B.n145 VSUBS 0.008212f
C415 B.n146 VSUBS 0.008212f
C416 B.n147 VSUBS 0.008212f
C417 B.n148 VSUBS 0.008212f
C418 B.n149 VSUBS 0.008212f
C419 B.n150 VSUBS 0.008212f
C420 B.n151 VSUBS 0.008212f
C421 B.n152 VSUBS 0.008212f
C422 B.n153 VSUBS 0.020215f
C423 B.n154 VSUBS 0.021086f
C424 B.n155 VSUBS 0.021086f
C425 B.n156 VSUBS 0.008212f
C426 B.n157 VSUBS 0.008212f
C427 B.n158 VSUBS 0.008212f
C428 B.n159 VSUBS 0.008212f
C429 B.n160 VSUBS 0.008212f
C430 B.n161 VSUBS 0.008212f
C431 B.n162 VSUBS 0.008212f
C432 B.n163 VSUBS 0.008212f
C433 B.n164 VSUBS 0.008212f
C434 B.n165 VSUBS 0.008212f
C435 B.n166 VSUBS 0.008212f
C436 B.n167 VSUBS 0.008212f
C437 B.n168 VSUBS 0.008212f
C438 B.n169 VSUBS 0.008212f
C439 B.n170 VSUBS 0.008212f
C440 B.n171 VSUBS 0.008212f
C441 B.n172 VSUBS 0.008212f
C442 B.n173 VSUBS 0.007729f
C443 B.n174 VSUBS 0.019026f
C444 B.n175 VSUBS 0.004589f
C445 B.n176 VSUBS 0.008212f
C446 B.n177 VSUBS 0.008212f
C447 B.n178 VSUBS 0.008212f
C448 B.n179 VSUBS 0.008212f
C449 B.n180 VSUBS 0.008212f
C450 B.n181 VSUBS 0.008212f
C451 B.n182 VSUBS 0.008212f
C452 B.n183 VSUBS 0.008212f
C453 B.n184 VSUBS 0.008212f
C454 B.n185 VSUBS 0.008212f
C455 B.n186 VSUBS 0.008212f
C456 B.n187 VSUBS 0.008212f
C457 B.n188 VSUBS 0.004589f
C458 B.n189 VSUBS 0.008212f
C459 B.n190 VSUBS 0.008212f
C460 B.n191 VSUBS 0.007729f
C461 B.n192 VSUBS 0.008212f
C462 B.n193 VSUBS 0.008212f
C463 B.n194 VSUBS 0.008212f
C464 B.n195 VSUBS 0.008212f
C465 B.n196 VSUBS 0.008212f
C466 B.n197 VSUBS 0.008212f
C467 B.n198 VSUBS 0.008212f
C468 B.n199 VSUBS 0.008212f
C469 B.n200 VSUBS 0.008212f
C470 B.n201 VSUBS 0.008212f
C471 B.n202 VSUBS 0.008212f
C472 B.n203 VSUBS 0.008212f
C473 B.n204 VSUBS 0.008212f
C474 B.n205 VSUBS 0.008212f
C475 B.n206 VSUBS 0.008212f
C476 B.n207 VSUBS 0.008212f
C477 B.n208 VSUBS 0.021086f
C478 B.n209 VSUBS 0.021086f
C479 B.n210 VSUBS 0.020215f
C480 B.n211 VSUBS 0.008212f
C481 B.n212 VSUBS 0.008212f
C482 B.n213 VSUBS 0.008212f
C483 B.n214 VSUBS 0.008212f
C484 B.n215 VSUBS 0.008212f
C485 B.n216 VSUBS 0.008212f
C486 B.n217 VSUBS 0.008212f
C487 B.n218 VSUBS 0.008212f
C488 B.n219 VSUBS 0.008212f
C489 B.n220 VSUBS 0.008212f
C490 B.n221 VSUBS 0.008212f
C491 B.n222 VSUBS 0.008212f
C492 B.n223 VSUBS 0.008212f
C493 B.n224 VSUBS 0.008212f
C494 B.n225 VSUBS 0.008212f
C495 B.n226 VSUBS 0.008212f
C496 B.n227 VSUBS 0.008212f
C497 B.n228 VSUBS 0.008212f
C498 B.n229 VSUBS 0.008212f
C499 B.n230 VSUBS 0.008212f
C500 B.n231 VSUBS 0.008212f
C501 B.n232 VSUBS 0.008212f
C502 B.n233 VSUBS 0.008212f
C503 B.n234 VSUBS 0.008212f
C504 B.n235 VSUBS 0.008212f
C505 B.n236 VSUBS 0.008212f
C506 B.n237 VSUBS 0.008212f
C507 B.n238 VSUBS 0.008212f
C508 B.n239 VSUBS 0.008212f
C509 B.n240 VSUBS 0.008212f
C510 B.n241 VSUBS 0.008212f
C511 B.n242 VSUBS 0.008212f
C512 B.n243 VSUBS 0.008212f
C513 B.n244 VSUBS 0.008212f
C514 B.n245 VSUBS 0.008212f
C515 B.n246 VSUBS 0.008212f
C516 B.n247 VSUBS 0.008212f
C517 B.n248 VSUBS 0.008212f
C518 B.n249 VSUBS 0.008212f
C519 B.n250 VSUBS 0.008212f
C520 B.n251 VSUBS 0.008212f
C521 B.n252 VSUBS 0.008212f
C522 B.n253 VSUBS 0.008212f
C523 B.n254 VSUBS 0.008212f
C524 B.n255 VSUBS 0.008212f
C525 B.n256 VSUBS 0.008212f
C526 B.n257 VSUBS 0.008212f
C527 B.n258 VSUBS 0.008212f
C528 B.n259 VSUBS 0.008212f
C529 B.n260 VSUBS 0.008212f
C530 B.n261 VSUBS 0.008212f
C531 B.n262 VSUBS 0.008212f
C532 B.n263 VSUBS 0.008212f
C533 B.n264 VSUBS 0.008212f
C534 B.n265 VSUBS 0.008212f
C535 B.n266 VSUBS 0.008212f
C536 B.n267 VSUBS 0.008212f
C537 B.n268 VSUBS 0.008212f
C538 B.n269 VSUBS 0.008212f
C539 B.n270 VSUBS 0.008212f
C540 B.n271 VSUBS 0.008212f
C541 B.n272 VSUBS 0.008212f
C542 B.n273 VSUBS 0.008212f
C543 B.n274 VSUBS 0.008212f
C544 B.n275 VSUBS 0.008212f
C545 B.n276 VSUBS 0.008212f
C546 B.n277 VSUBS 0.008212f
C547 B.n278 VSUBS 0.008212f
C548 B.n279 VSUBS 0.008212f
C549 B.n280 VSUBS 0.008212f
C550 B.n281 VSUBS 0.008212f
C551 B.n282 VSUBS 0.008212f
C552 B.n283 VSUBS 0.008212f
C553 B.n284 VSUBS 0.008212f
C554 B.n285 VSUBS 0.008212f
C555 B.n286 VSUBS 0.008212f
C556 B.n287 VSUBS 0.008212f
C557 B.n288 VSUBS 0.008212f
C558 B.n289 VSUBS 0.008212f
C559 B.n290 VSUBS 0.008212f
C560 B.n291 VSUBS 0.008212f
C561 B.n292 VSUBS 0.008212f
C562 B.n293 VSUBS 0.008212f
C563 B.n294 VSUBS 0.008212f
C564 B.n295 VSUBS 0.008212f
C565 B.n296 VSUBS 0.008212f
C566 B.n297 VSUBS 0.008212f
C567 B.n298 VSUBS 0.008212f
C568 B.n299 VSUBS 0.008212f
C569 B.n300 VSUBS 0.008212f
C570 B.n301 VSUBS 0.008212f
C571 B.n302 VSUBS 0.008212f
C572 B.n303 VSUBS 0.020215f
C573 B.n304 VSUBS 0.021086f
C574 B.n305 VSUBS 0.020215f
C575 B.n306 VSUBS 0.008212f
C576 B.n307 VSUBS 0.008212f
C577 B.n308 VSUBS 0.008212f
C578 B.n309 VSUBS 0.008212f
C579 B.n310 VSUBS 0.008212f
C580 B.n311 VSUBS 0.008212f
C581 B.n312 VSUBS 0.008212f
C582 B.n313 VSUBS 0.008212f
C583 B.n314 VSUBS 0.008212f
C584 B.n315 VSUBS 0.008212f
C585 B.n316 VSUBS 0.008212f
C586 B.n317 VSUBS 0.008212f
C587 B.n318 VSUBS 0.008212f
C588 B.n319 VSUBS 0.008212f
C589 B.n320 VSUBS 0.008212f
C590 B.n321 VSUBS 0.008212f
C591 B.n322 VSUBS 0.008212f
C592 B.n323 VSUBS 0.007729f
C593 B.n324 VSUBS 0.019026f
C594 B.n325 VSUBS 0.004589f
C595 B.n326 VSUBS 0.008212f
C596 B.n327 VSUBS 0.008212f
C597 B.n328 VSUBS 0.008212f
C598 B.n329 VSUBS 0.008212f
C599 B.n330 VSUBS 0.008212f
C600 B.n331 VSUBS 0.008212f
C601 B.n332 VSUBS 0.008212f
C602 B.n333 VSUBS 0.008212f
C603 B.n334 VSUBS 0.008212f
C604 B.n335 VSUBS 0.008212f
C605 B.n336 VSUBS 0.008212f
C606 B.n337 VSUBS 0.008212f
C607 B.n338 VSUBS 0.004589f
C608 B.n339 VSUBS 0.008212f
C609 B.n340 VSUBS 0.008212f
C610 B.n341 VSUBS 0.007729f
C611 B.n342 VSUBS 0.008212f
C612 B.n343 VSUBS 0.008212f
C613 B.n344 VSUBS 0.008212f
C614 B.n345 VSUBS 0.008212f
C615 B.n346 VSUBS 0.008212f
C616 B.n347 VSUBS 0.008212f
C617 B.n348 VSUBS 0.008212f
C618 B.n349 VSUBS 0.008212f
C619 B.n350 VSUBS 0.008212f
C620 B.n351 VSUBS 0.008212f
C621 B.n352 VSUBS 0.008212f
C622 B.n353 VSUBS 0.008212f
C623 B.n354 VSUBS 0.008212f
C624 B.n355 VSUBS 0.008212f
C625 B.n356 VSUBS 0.008212f
C626 B.n357 VSUBS 0.008212f
C627 B.n358 VSUBS 0.021086f
C628 B.n359 VSUBS 0.021086f
C629 B.n360 VSUBS 0.020215f
C630 B.n361 VSUBS 0.008212f
C631 B.n362 VSUBS 0.008212f
C632 B.n363 VSUBS 0.008212f
C633 B.n364 VSUBS 0.008212f
C634 B.n365 VSUBS 0.008212f
C635 B.n366 VSUBS 0.008212f
C636 B.n367 VSUBS 0.008212f
C637 B.n368 VSUBS 0.008212f
C638 B.n369 VSUBS 0.008212f
C639 B.n370 VSUBS 0.008212f
C640 B.n371 VSUBS 0.008212f
C641 B.n372 VSUBS 0.008212f
C642 B.n373 VSUBS 0.008212f
C643 B.n374 VSUBS 0.008212f
C644 B.n375 VSUBS 0.008212f
C645 B.n376 VSUBS 0.008212f
C646 B.n377 VSUBS 0.008212f
C647 B.n378 VSUBS 0.008212f
C648 B.n379 VSUBS 0.008212f
C649 B.n380 VSUBS 0.008212f
C650 B.n381 VSUBS 0.008212f
C651 B.n382 VSUBS 0.008212f
C652 B.n383 VSUBS 0.008212f
C653 B.n384 VSUBS 0.008212f
C654 B.n385 VSUBS 0.008212f
C655 B.n386 VSUBS 0.008212f
C656 B.n387 VSUBS 0.008212f
C657 B.n388 VSUBS 0.008212f
C658 B.n389 VSUBS 0.008212f
C659 B.n390 VSUBS 0.008212f
C660 B.n391 VSUBS 0.008212f
C661 B.n392 VSUBS 0.008212f
C662 B.n393 VSUBS 0.008212f
C663 B.n394 VSUBS 0.008212f
C664 B.n395 VSUBS 0.008212f
C665 B.n396 VSUBS 0.008212f
C666 B.n397 VSUBS 0.008212f
C667 B.n398 VSUBS 0.008212f
C668 B.n399 VSUBS 0.008212f
C669 B.n400 VSUBS 0.008212f
C670 B.n401 VSUBS 0.008212f
C671 B.n402 VSUBS 0.008212f
C672 B.n403 VSUBS 0.008212f
C673 B.n404 VSUBS 0.008212f
C674 B.n405 VSUBS 0.008212f
C675 B.n406 VSUBS 0.008212f
C676 B.n407 VSUBS 0.018594f
.ends

