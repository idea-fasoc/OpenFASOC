* NGSPICE file created from diff_pair_sample_0568.ext - technology: sky130A

.subckt diff_pair_sample_0568 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t0 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=2.1945 pd=13.63 as=5.187 ps=27.38 w=13.3 l=1.64
X1 VDD1.t2 VP.t1 VTAIL.t1 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=2.1945 pd=13.63 as=5.187 ps=27.38 w=13.3 l=1.64
X2 B.t11 B.t9 B.t10 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=0 ps=0 w=13.3 l=1.64
X3 B.t8 B.t6 B.t7 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=0 ps=0 w=13.3 l=1.64
X4 VTAIL.t4 VN.t0 VDD2.t3 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=2.1945 ps=13.63 w=13.3 l=1.64
X5 VTAIL.t5 VN.t1 VDD2.t2 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=2.1945 ps=13.63 w=13.3 l=1.64
X6 B.t5 B.t3 B.t4 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=0 ps=0 w=13.3 l=1.64
X7 VTAIL.t3 VP.t2 VDD1.t1 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=2.1945 ps=13.63 w=13.3 l=1.64
X8 VDD2.t1 VN.t2 VTAIL.t7 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=2.1945 pd=13.63 as=5.187 ps=27.38 w=13.3 l=1.64
X9 VDD2.t0 VN.t3 VTAIL.t6 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=2.1945 pd=13.63 as=5.187 ps=27.38 w=13.3 l=1.64
X10 B.t2 B.t0 B.t1 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=0 ps=0 w=13.3 l=1.64
X11 VTAIL.t2 VP.t3 VDD1.t0 w_n2152_n3628# sky130_fd_pr__pfet_01v8 ad=5.187 pd=27.38 as=2.1945 ps=13.63 w=13.3 l=1.64
R0 VP.n2 VP.t2 233.706
R1 VP.n2 VP.t1 233.377
R2 VP.n4 VP.t3 195.446
R3 VP.n11 VP.t0 195.446
R4 VP.n4 VP.n3 174.202
R5 VP.n12 VP.n11 174.202
R6 VP.n10 VP.n0 161.3
R7 VP.n9 VP.n8 161.3
R8 VP.n7 VP.n1 161.3
R9 VP.n6 VP.n5 161.3
R10 VP.n3 VP.n2 56.9317
R11 VP.n9 VP.n1 56.4773
R12 VP.n5 VP.n1 24.3439
R13 VP.n10 VP.n9 24.3439
R14 VP.n5 VP.n4 11.4419
R15 VP.n11 VP.n10 11.4419
R16 VP.n6 VP.n3 0.189894
R17 VP.n7 VP.n6 0.189894
R18 VP.n8 VP.n7 0.189894
R19 VP.n8 VP.n0 0.189894
R20 VP.n12 VP.n0 0.189894
R21 VP VP.n12 0.0516364
R22 VTAIL.n529 VTAIL.n528 585
R23 VTAIL.n531 VTAIL.n530 585
R24 VTAIL.n524 VTAIL.n523 585
R25 VTAIL.n537 VTAIL.n536 585
R26 VTAIL.n539 VTAIL.n538 585
R27 VTAIL.n520 VTAIL.n519 585
R28 VTAIL.n545 VTAIL.n544 585
R29 VTAIL.n547 VTAIL.n546 585
R30 VTAIL.n516 VTAIL.n515 585
R31 VTAIL.n553 VTAIL.n552 585
R32 VTAIL.n555 VTAIL.n554 585
R33 VTAIL.n512 VTAIL.n511 585
R34 VTAIL.n561 VTAIL.n560 585
R35 VTAIL.n563 VTAIL.n562 585
R36 VTAIL.n508 VTAIL.n507 585
R37 VTAIL.n569 VTAIL.n568 585
R38 VTAIL.n571 VTAIL.n570 585
R39 VTAIL.n25 VTAIL.n24 585
R40 VTAIL.n27 VTAIL.n26 585
R41 VTAIL.n20 VTAIL.n19 585
R42 VTAIL.n33 VTAIL.n32 585
R43 VTAIL.n35 VTAIL.n34 585
R44 VTAIL.n16 VTAIL.n15 585
R45 VTAIL.n41 VTAIL.n40 585
R46 VTAIL.n43 VTAIL.n42 585
R47 VTAIL.n12 VTAIL.n11 585
R48 VTAIL.n49 VTAIL.n48 585
R49 VTAIL.n51 VTAIL.n50 585
R50 VTAIL.n8 VTAIL.n7 585
R51 VTAIL.n57 VTAIL.n56 585
R52 VTAIL.n59 VTAIL.n58 585
R53 VTAIL.n4 VTAIL.n3 585
R54 VTAIL.n65 VTAIL.n64 585
R55 VTAIL.n67 VTAIL.n66 585
R56 VTAIL.n97 VTAIL.n96 585
R57 VTAIL.n99 VTAIL.n98 585
R58 VTAIL.n92 VTAIL.n91 585
R59 VTAIL.n105 VTAIL.n104 585
R60 VTAIL.n107 VTAIL.n106 585
R61 VTAIL.n88 VTAIL.n87 585
R62 VTAIL.n113 VTAIL.n112 585
R63 VTAIL.n115 VTAIL.n114 585
R64 VTAIL.n84 VTAIL.n83 585
R65 VTAIL.n121 VTAIL.n120 585
R66 VTAIL.n123 VTAIL.n122 585
R67 VTAIL.n80 VTAIL.n79 585
R68 VTAIL.n129 VTAIL.n128 585
R69 VTAIL.n131 VTAIL.n130 585
R70 VTAIL.n76 VTAIL.n75 585
R71 VTAIL.n137 VTAIL.n136 585
R72 VTAIL.n139 VTAIL.n138 585
R73 VTAIL.n169 VTAIL.n168 585
R74 VTAIL.n171 VTAIL.n170 585
R75 VTAIL.n164 VTAIL.n163 585
R76 VTAIL.n177 VTAIL.n176 585
R77 VTAIL.n179 VTAIL.n178 585
R78 VTAIL.n160 VTAIL.n159 585
R79 VTAIL.n185 VTAIL.n184 585
R80 VTAIL.n187 VTAIL.n186 585
R81 VTAIL.n156 VTAIL.n155 585
R82 VTAIL.n193 VTAIL.n192 585
R83 VTAIL.n195 VTAIL.n194 585
R84 VTAIL.n152 VTAIL.n151 585
R85 VTAIL.n201 VTAIL.n200 585
R86 VTAIL.n203 VTAIL.n202 585
R87 VTAIL.n148 VTAIL.n147 585
R88 VTAIL.n209 VTAIL.n208 585
R89 VTAIL.n211 VTAIL.n210 585
R90 VTAIL.n499 VTAIL.n498 585
R91 VTAIL.n497 VTAIL.n496 585
R92 VTAIL.n436 VTAIL.n435 585
R93 VTAIL.n491 VTAIL.n490 585
R94 VTAIL.n489 VTAIL.n488 585
R95 VTAIL.n440 VTAIL.n439 585
R96 VTAIL.n483 VTAIL.n482 585
R97 VTAIL.n481 VTAIL.n480 585
R98 VTAIL.n444 VTAIL.n443 585
R99 VTAIL.n475 VTAIL.n474 585
R100 VTAIL.n473 VTAIL.n472 585
R101 VTAIL.n448 VTAIL.n447 585
R102 VTAIL.n467 VTAIL.n466 585
R103 VTAIL.n465 VTAIL.n464 585
R104 VTAIL.n452 VTAIL.n451 585
R105 VTAIL.n459 VTAIL.n458 585
R106 VTAIL.n457 VTAIL.n456 585
R107 VTAIL.n427 VTAIL.n426 585
R108 VTAIL.n425 VTAIL.n424 585
R109 VTAIL.n364 VTAIL.n363 585
R110 VTAIL.n419 VTAIL.n418 585
R111 VTAIL.n417 VTAIL.n416 585
R112 VTAIL.n368 VTAIL.n367 585
R113 VTAIL.n411 VTAIL.n410 585
R114 VTAIL.n409 VTAIL.n408 585
R115 VTAIL.n372 VTAIL.n371 585
R116 VTAIL.n403 VTAIL.n402 585
R117 VTAIL.n401 VTAIL.n400 585
R118 VTAIL.n376 VTAIL.n375 585
R119 VTAIL.n395 VTAIL.n394 585
R120 VTAIL.n393 VTAIL.n392 585
R121 VTAIL.n380 VTAIL.n379 585
R122 VTAIL.n387 VTAIL.n386 585
R123 VTAIL.n385 VTAIL.n384 585
R124 VTAIL.n355 VTAIL.n354 585
R125 VTAIL.n353 VTAIL.n352 585
R126 VTAIL.n292 VTAIL.n291 585
R127 VTAIL.n347 VTAIL.n346 585
R128 VTAIL.n345 VTAIL.n344 585
R129 VTAIL.n296 VTAIL.n295 585
R130 VTAIL.n339 VTAIL.n338 585
R131 VTAIL.n337 VTAIL.n336 585
R132 VTAIL.n300 VTAIL.n299 585
R133 VTAIL.n331 VTAIL.n330 585
R134 VTAIL.n329 VTAIL.n328 585
R135 VTAIL.n304 VTAIL.n303 585
R136 VTAIL.n323 VTAIL.n322 585
R137 VTAIL.n321 VTAIL.n320 585
R138 VTAIL.n308 VTAIL.n307 585
R139 VTAIL.n315 VTAIL.n314 585
R140 VTAIL.n313 VTAIL.n312 585
R141 VTAIL.n283 VTAIL.n282 585
R142 VTAIL.n281 VTAIL.n280 585
R143 VTAIL.n220 VTAIL.n219 585
R144 VTAIL.n275 VTAIL.n274 585
R145 VTAIL.n273 VTAIL.n272 585
R146 VTAIL.n224 VTAIL.n223 585
R147 VTAIL.n267 VTAIL.n266 585
R148 VTAIL.n265 VTAIL.n264 585
R149 VTAIL.n228 VTAIL.n227 585
R150 VTAIL.n259 VTAIL.n258 585
R151 VTAIL.n257 VTAIL.n256 585
R152 VTAIL.n232 VTAIL.n231 585
R153 VTAIL.n251 VTAIL.n250 585
R154 VTAIL.n249 VTAIL.n248 585
R155 VTAIL.n236 VTAIL.n235 585
R156 VTAIL.n243 VTAIL.n242 585
R157 VTAIL.n241 VTAIL.n240 585
R158 VTAIL.n570 VTAIL.n504 498.474
R159 VTAIL.n66 VTAIL.n0 498.474
R160 VTAIL.n138 VTAIL.n72 498.474
R161 VTAIL.n210 VTAIL.n144 498.474
R162 VTAIL.n498 VTAIL.n432 498.474
R163 VTAIL.n426 VTAIL.n360 498.474
R164 VTAIL.n354 VTAIL.n288 498.474
R165 VTAIL.n282 VTAIL.n216 498.474
R166 VTAIL.n527 VTAIL.t6 327.466
R167 VTAIL.n23 VTAIL.t4 327.466
R168 VTAIL.n95 VTAIL.t0 327.466
R169 VTAIL.n167 VTAIL.t2 327.466
R170 VTAIL.n455 VTAIL.t1 327.466
R171 VTAIL.n383 VTAIL.t3 327.466
R172 VTAIL.n311 VTAIL.t7 327.466
R173 VTAIL.n239 VTAIL.t5 327.466
R174 VTAIL.n530 VTAIL.n529 171.744
R175 VTAIL.n530 VTAIL.n523 171.744
R176 VTAIL.n537 VTAIL.n523 171.744
R177 VTAIL.n538 VTAIL.n537 171.744
R178 VTAIL.n538 VTAIL.n519 171.744
R179 VTAIL.n545 VTAIL.n519 171.744
R180 VTAIL.n546 VTAIL.n545 171.744
R181 VTAIL.n546 VTAIL.n515 171.744
R182 VTAIL.n553 VTAIL.n515 171.744
R183 VTAIL.n554 VTAIL.n553 171.744
R184 VTAIL.n554 VTAIL.n511 171.744
R185 VTAIL.n561 VTAIL.n511 171.744
R186 VTAIL.n562 VTAIL.n561 171.744
R187 VTAIL.n562 VTAIL.n507 171.744
R188 VTAIL.n569 VTAIL.n507 171.744
R189 VTAIL.n570 VTAIL.n569 171.744
R190 VTAIL.n26 VTAIL.n25 171.744
R191 VTAIL.n26 VTAIL.n19 171.744
R192 VTAIL.n33 VTAIL.n19 171.744
R193 VTAIL.n34 VTAIL.n33 171.744
R194 VTAIL.n34 VTAIL.n15 171.744
R195 VTAIL.n41 VTAIL.n15 171.744
R196 VTAIL.n42 VTAIL.n41 171.744
R197 VTAIL.n42 VTAIL.n11 171.744
R198 VTAIL.n49 VTAIL.n11 171.744
R199 VTAIL.n50 VTAIL.n49 171.744
R200 VTAIL.n50 VTAIL.n7 171.744
R201 VTAIL.n57 VTAIL.n7 171.744
R202 VTAIL.n58 VTAIL.n57 171.744
R203 VTAIL.n58 VTAIL.n3 171.744
R204 VTAIL.n65 VTAIL.n3 171.744
R205 VTAIL.n66 VTAIL.n65 171.744
R206 VTAIL.n98 VTAIL.n97 171.744
R207 VTAIL.n98 VTAIL.n91 171.744
R208 VTAIL.n105 VTAIL.n91 171.744
R209 VTAIL.n106 VTAIL.n105 171.744
R210 VTAIL.n106 VTAIL.n87 171.744
R211 VTAIL.n113 VTAIL.n87 171.744
R212 VTAIL.n114 VTAIL.n113 171.744
R213 VTAIL.n114 VTAIL.n83 171.744
R214 VTAIL.n121 VTAIL.n83 171.744
R215 VTAIL.n122 VTAIL.n121 171.744
R216 VTAIL.n122 VTAIL.n79 171.744
R217 VTAIL.n129 VTAIL.n79 171.744
R218 VTAIL.n130 VTAIL.n129 171.744
R219 VTAIL.n130 VTAIL.n75 171.744
R220 VTAIL.n137 VTAIL.n75 171.744
R221 VTAIL.n138 VTAIL.n137 171.744
R222 VTAIL.n170 VTAIL.n169 171.744
R223 VTAIL.n170 VTAIL.n163 171.744
R224 VTAIL.n177 VTAIL.n163 171.744
R225 VTAIL.n178 VTAIL.n177 171.744
R226 VTAIL.n178 VTAIL.n159 171.744
R227 VTAIL.n185 VTAIL.n159 171.744
R228 VTAIL.n186 VTAIL.n185 171.744
R229 VTAIL.n186 VTAIL.n155 171.744
R230 VTAIL.n193 VTAIL.n155 171.744
R231 VTAIL.n194 VTAIL.n193 171.744
R232 VTAIL.n194 VTAIL.n151 171.744
R233 VTAIL.n201 VTAIL.n151 171.744
R234 VTAIL.n202 VTAIL.n201 171.744
R235 VTAIL.n202 VTAIL.n147 171.744
R236 VTAIL.n209 VTAIL.n147 171.744
R237 VTAIL.n210 VTAIL.n209 171.744
R238 VTAIL.n498 VTAIL.n497 171.744
R239 VTAIL.n497 VTAIL.n435 171.744
R240 VTAIL.n490 VTAIL.n435 171.744
R241 VTAIL.n490 VTAIL.n489 171.744
R242 VTAIL.n489 VTAIL.n439 171.744
R243 VTAIL.n482 VTAIL.n439 171.744
R244 VTAIL.n482 VTAIL.n481 171.744
R245 VTAIL.n481 VTAIL.n443 171.744
R246 VTAIL.n474 VTAIL.n443 171.744
R247 VTAIL.n474 VTAIL.n473 171.744
R248 VTAIL.n473 VTAIL.n447 171.744
R249 VTAIL.n466 VTAIL.n447 171.744
R250 VTAIL.n466 VTAIL.n465 171.744
R251 VTAIL.n465 VTAIL.n451 171.744
R252 VTAIL.n458 VTAIL.n451 171.744
R253 VTAIL.n458 VTAIL.n457 171.744
R254 VTAIL.n426 VTAIL.n425 171.744
R255 VTAIL.n425 VTAIL.n363 171.744
R256 VTAIL.n418 VTAIL.n363 171.744
R257 VTAIL.n418 VTAIL.n417 171.744
R258 VTAIL.n417 VTAIL.n367 171.744
R259 VTAIL.n410 VTAIL.n367 171.744
R260 VTAIL.n410 VTAIL.n409 171.744
R261 VTAIL.n409 VTAIL.n371 171.744
R262 VTAIL.n402 VTAIL.n371 171.744
R263 VTAIL.n402 VTAIL.n401 171.744
R264 VTAIL.n401 VTAIL.n375 171.744
R265 VTAIL.n394 VTAIL.n375 171.744
R266 VTAIL.n394 VTAIL.n393 171.744
R267 VTAIL.n393 VTAIL.n379 171.744
R268 VTAIL.n386 VTAIL.n379 171.744
R269 VTAIL.n386 VTAIL.n385 171.744
R270 VTAIL.n354 VTAIL.n353 171.744
R271 VTAIL.n353 VTAIL.n291 171.744
R272 VTAIL.n346 VTAIL.n291 171.744
R273 VTAIL.n346 VTAIL.n345 171.744
R274 VTAIL.n345 VTAIL.n295 171.744
R275 VTAIL.n338 VTAIL.n295 171.744
R276 VTAIL.n338 VTAIL.n337 171.744
R277 VTAIL.n337 VTAIL.n299 171.744
R278 VTAIL.n330 VTAIL.n299 171.744
R279 VTAIL.n330 VTAIL.n329 171.744
R280 VTAIL.n329 VTAIL.n303 171.744
R281 VTAIL.n322 VTAIL.n303 171.744
R282 VTAIL.n322 VTAIL.n321 171.744
R283 VTAIL.n321 VTAIL.n307 171.744
R284 VTAIL.n314 VTAIL.n307 171.744
R285 VTAIL.n314 VTAIL.n313 171.744
R286 VTAIL.n282 VTAIL.n281 171.744
R287 VTAIL.n281 VTAIL.n219 171.744
R288 VTAIL.n274 VTAIL.n219 171.744
R289 VTAIL.n274 VTAIL.n273 171.744
R290 VTAIL.n273 VTAIL.n223 171.744
R291 VTAIL.n266 VTAIL.n223 171.744
R292 VTAIL.n266 VTAIL.n265 171.744
R293 VTAIL.n265 VTAIL.n227 171.744
R294 VTAIL.n258 VTAIL.n227 171.744
R295 VTAIL.n258 VTAIL.n257 171.744
R296 VTAIL.n257 VTAIL.n231 171.744
R297 VTAIL.n250 VTAIL.n231 171.744
R298 VTAIL.n250 VTAIL.n249 171.744
R299 VTAIL.n249 VTAIL.n235 171.744
R300 VTAIL.n242 VTAIL.n235 171.744
R301 VTAIL.n242 VTAIL.n241 171.744
R302 VTAIL.n529 VTAIL.t6 85.8723
R303 VTAIL.n25 VTAIL.t4 85.8723
R304 VTAIL.n97 VTAIL.t0 85.8723
R305 VTAIL.n169 VTAIL.t2 85.8723
R306 VTAIL.n457 VTAIL.t1 85.8723
R307 VTAIL.n385 VTAIL.t3 85.8723
R308 VTAIL.n313 VTAIL.t7 85.8723
R309 VTAIL.n241 VTAIL.t5 85.8723
R310 VTAIL.n575 VTAIL.n574 34.1247
R311 VTAIL.n71 VTAIL.n70 34.1247
R312 VTAIL.n143 VTAIL.n142 34.1247
R313 VTAIL.n215 VTAIL.n214 34.1247
R314 VTAIL.n503 VTAIL.n502 34.1247
R315 VTAIL.n431 VTAIL.n430 34.1247
R316 VTAIL.n359 VTAIL.n358 34.1247
R317 VTAIL.n287 VTAIL.n286 34.1247
R318 VTAIL.n575 VTAIL.n503 25.5307
R319 VTAIL.n287 VTAIL.n215 25.5307
R320 VTAIL.n528 VTAIL.n527 16.3895
R321 VTAIL.n24 VTAIL.n23 16.3895
R322 VTAIL.n96 VTAIL.n95 16.3895
R323 VTAIL.n168 VTAIL.n167 16.3895
R324 VTAIL.n456 VTAIL.n455 16.3895
R325 VTAIL.n384 VTAIL.n383 16.3895
R326 VTAIL.n312 VTAIL.n311 16.3895
R327 VTAIL.n240 VTAIL.n239 16.3895
R328 VTAIL.n531 VTAIL.n526 12.8005
R329 VTAIL.n572 VTAIL.n571 12.8005
R330 VTAIL.n27 VTAIL.n22 12.8005
R331 VTAIL.n68 VTAIL.n67 12.8005
R332 VTAIL.n99 VTAIL.n94 12.8005
R333 VTAIL.n140 VTAIL.n139 12.8005
R334 VTAIL.n171 VTAIL.n166 12.8005
R335 VTAIL.n212 VTAIL.n211 12.8005
R336 VTAIL.n500 VTAIL.n499 12.8005
R337 VTAIL.n459 VTAIL.n454 12.8005
R338 VTAIL.n428 VTAIL.n427 12.8005
R339 VTAIL.n387 VTAIL.n382 12.8005
R340 VTAIL.n356 VTAIL.n355 12.8005
R341 VTAIL.n315 VTAIL.n310 12.8005
R342 VTAIL.n284 VTAIL.n283 12.8005
R343 VTAIL.n243 VTAIL.n238 12.8005
R344 VTAIL.n532 VTAIL.n524 12.0247
R345 VTAIL.n568 VTAIL.n506 12.0247
R346 VTAIL.n28 VTAIL.n20 12.0247
R347 VTAIL.n64 VTAIL.n2 12.0247
R348 VTAIL.n100 VTAIL.n92 12.0247
R349 VTAIL.n136 VTAIL.n74 12.0247
R350 VTAIL.n172 VTAIL.n164 12.0247
R351 VTAIL.n208 VTAIL.n146 12.0247
R352 VTAIL.n496 VTAIL.n434 12.0247
R353 VTAIL.n460 VTAIL.n452 12.0247
R354 VTAIL.n424 VTAIL.n362 12.0247
R355 VTAIL.n388 VTAIL.n380 12.0247
R356 VTAIL.n352 VTAIL.n290 12.0247
R357 VTAIL.n316 VTAIL.n308 12.0247
R358 VTAIL.n280 VTAIL.n218 12.0247
R359 VTAIL.n244 VTAIL.n236 12.0247
R360 VTAIL.n536 VTAIL.n535 11.249
R361 VTAIL.n567 VTAIL.n508 11.249
R362 VTAIL.n32 VTAIL.n31 11.249
R363 VTAIL.n63 VTAIL.n4 11.249
R364 VTAIL.n104 VTAIL.n103 11.249
R365 VTAIL.n135 VTAIL.n76 11.249
R366 VTAIL.n176 VTAIL.n175 11.249
R367 VTAIL.n207 VTAIL.n148 11.249
R368 VTAIL.n495 VTAIL.n436 11.249
R369 VTAIL.n464 VTAIL.n463 11.249
R370 VTAIL.n423 VTAIL.n364 11.249
R371 VTAIL.n392 VTAIL.n391 11.249
R372 VTAIL.n351 VTAIL.n292 11.249
R373 VTAIL.n320 VTAIL.n319 11.249
R374 VTAIL.n279 VTAIL.n220 11.249
R375 VTAIL.n248 VTAIL.n247 11.249
R376 VTAIL.n539 VTAIL.n522 10.4732
R377 VTAIL.n564 VTAIL.n563 10.4732
R378 VTAIL.n35 VTAIL.n18 10.4732
R379 VTAIL.n60 VTAIL.n59 10.4732
R380 VTAIL.n107 VTAIL.n90 10.4732
R381 VTAIL.n132 VTAIL.n131 10.4732
R382 VTAIL.n179 VTAIL.n162 10.4732
R383 VTAIL.n204 VTAIL.n203 10.4732
R384 VTAIL.n492 VTAIL.n491 10.4732
R385 VTAIL.n467 VTAIL.n450 10.4732
R386 VTAIL.n420 VTAIL.n419 10.4732
R387 VTAIL.n395 VTAIL.n378 10.4732
R388 VTAIL.n348 VTAIL.n347 10.4732
R389 VTAIL.n323 VTAIL.n306 10.4732
R390 VTAIL.n276 VTAIL.n275 10.4732
R391 VTAIL.n251 VTAIL.n234 10.4732
R392 VTAIL.n540 VTAIL.n520 9.69747
R393 VTAIL.n560 VTAIL.n510 9.69747
R394 VTAIL.n36 VTAIL.n16 9.69747
R395 VTAIL.n56 VTAIL.n6 9.69747
R396 VTAIL.n108 VTAIL.n88 9.69747
R397 VTAIL.n128 VTAIL.n78 9.69747
R398 VTAIL.n180 VTAIL.n160 9.69747
R399 VTAIL.n200 VTAIL.n150 9.69747
R400 VTAIL.n488 VTAIL.n438 9.69747
R401 VTAIL.n468 VTAIL.n448 9.69747
R402 VTAIL.n416 VTAIL.n366 9.69747
R403 VTAIL.n396 VTAIL.n376 9.69747
R404 VTAIL.n344 VTAIL.n294 9.69747
R405 VTAIL.n324 VTAIL.n304 9.69747
R406 VTAIL.n272 VTAIL.n222 9.69747
R407 VTAIL.n252 VTAIL.n232 9.69747
R408 VTAIL.n574 VTAIL.n573 9.45567
R409 VTAIL.n70 VTAIL.n69 9.45567
R410 VTAIL.n142 VTAIL.n141 9.45567
R411 VTAIL.n214 VTAIL.n213 9.45567
R412 VTAIL.n502 VTAIL.n501 9.45567
R413 VTAIL.n430 VTAIL.n429 9.45567
R414 VTAIL.n358 VTAIL.n357 9.45567
R415 VTAIL.n286 VTAIL.n285 9.45567
R416 VTAIL.n549 VTAIL.n548 9.3005
R417 VTAIL.n518 VTAIL.n517 9.3005
R418 VTAIL.n543 VTAIL.n542 9.3005
R419 VTAIL.n541 VTAIL.n540 9.3005
R420 VTAIL.n522 VTAIL.n521 9.3005
R421 VTAIL.n535 VTAIL.n534 9.3005
R422 VTAIL.n533 VTAIL.n532 9.3005
R423 VTAIL.n526 VTAIL.n525 9.3005
R424 VTAIL.n551 VTAIL.n550 9.3005
R425 VTAIL.n514 VTAIL.n513 9.3005
R426 VTAIL.n557 VTAIL.n556 9.3005
R427 VTAIL.n559 VTAIL.n558 9.3005
R428 VTAIL.n510 VTAIL.n509 9.3005
R429 VTAIL.n565 VTAIL.n564 9.3005
R430 VTAIL.n567 VTAIL.n566 9.3005
R431 VTAIL.n506 VTAIL.n505 9.3005
R432 VTAIL.n573 VTAIL.n572 9.3005
R433 VTAIL.n45 VTAIL.n44 9.3005
R434 VTAIL.n14 VTAIL.n13 9.3005
R435 VTAIL.n39 VTAIL.n38 9.3005
R436 VTAIL.n37 VTAIL.n36 9.3005
R437 VTAIL.n18 VTAIL.n17 9.3005
R438 VTAIL.n31 VTAIL.n30 9.3005
R439 VTAIL.n29 VTAIL.n28 9.3005
R440 VTAIL.n22 VTAIL.n21 9.3005
R441 VTAIL.n47 VTAIL.n46 9.3005
R442 VTAIL.n10 VTAIL.n9 9.3005
R443 VTAIL.n53 VTAIL.n52 9.3005
R444 VTAIL.n55 VTAIL.n54 9.3005
R445 VTAIL.n6 VTAIL.n5 9.3005
R446 VTAIL.n61 VTAIL.n60 9.3005
R447 VTAIL.n63 VTAIL.n62 9.3005
R448 VTAIL.n2 VTAIL.n1 9.3005
R449 VTAIL.n69 VTAIL.n68 9.3005
R450 VTAIL.n117 VTAIL.n116 9.3005
R451 VTAIL.n86 VTAIL.n85 9.3005
R452 VTAIL.n111 VTAIL.n110 9.3005
R453 VTAIL.n109 VTAIL.n108 9.3005
R454 VTAIL.n90 VTAIL.n89 9.3005
R455 VTAIL.n103 VTAIL.n102 9.3005
R456 VTAIL.n101 VTAIL.n100 9.3005
R457 VTAIL.n94 VTAIL.n93 9.3005
R458 VTAIL.n119 VTAIL.n118 9.3005
R459 VTAIL.n82 VTAIL.n81 9.3005
R460 VTAIL.n125 VTAIL.n124 9.3005
R461 VTAIL.n127 VTAIL.n126 9.3005
R462 VTAIL.n78 VTAIL.n77 9.3005
R463 VTAIL.n133 VTAIL.n132 9.3005
R464 VTAIL.n135 VTAIL.n134 9.3005
R465 VTAIL.n74 VTAIL.n73 9.3005
R466 VTAIL.n141 VTAIL.n140 9.3005
R467 VTAIL.n189 VTAIL.n188 9.3005
R468 VTAIL.n158 VTAIL.n157 9.3005
R469 VTAIL.n183 VTAIL.n182 9.3005
R470 VTAIL.n181 VTAIL.n180 9.3005
R471 VTAIL.n162 VTAIL.n161 9.3005
R472 VTAIL.n175 VTAIL.n174 9.3005
R473 VTAIL.n173 VTAIL.n172 9.3005
R474 VTAIL.n166 VTAIL.n165 9.3005
R475 VTAIL.n191 VTAIL.n190 9.3005
R476 VTAIL.n154 VTAIL.n153 9.3005
R477 VTAIL.n197 VTAIL.n196 9.3005
R478 VTAIL.n199 VTAIL.n198 9.3005
R479 VTAIL.n150 VTAIL.n149 9.3005
R480 VTAIL.n205 VTAIL.n204 9.3005
R481 VTAIL.n207 VTAIL.n206 9.3005
R482 VTAIL.n146 VTAIL.n145 9.3005
R483 VTAIL.n213 VTAIL.n212 9.3005
R484 VTAIL.n442 VTAIL.n441 9.3005
R485 VTAIL.n485 VTAIL.n484 9.3005
R486 VTAIL.n487 VTAIL.n486 9.3005
R487 VTAIL.n438 VTAIL.n437 9.3005
R488 VTAIL.n493 VTAIL.n492 9.3005
R489 VTAIL.n495 VTAIL.n494 9.3005
R490 VTAIL.n434 VTAIL.n433 9.3005
R491 VTAIL.n501 VTAIL.n500 9.3005
R492 VTAIL.n479 VTAIL.n478 9.3005
R493 VTAIL.n477 VTAIL.n476 9.3005
R494 VTAIL.n446 VTAIL.n445 9.3005
R495 VTAIL.n471 VTAIL.n470 9.3005
R496 VTAIL.n469 VTAIL.n468 9.3005
R497 VTAIL.n450 VTAIL.n449 9.3005
R498 VTAIL.n463 VTAIL.n462 9.3005
R499 VTAIL.n461 VTAIL.n460 9.3005
R500 VTAIL.n454 VTAIL.n453 9.3005
R501 VTAIL.n370 VTAIL.n369 9.3005
R502 VTAIL.n413 VTAIL.n412 9.3005
R503 VTAIL.n415 VTAIL.n414 9.3005
R504 VTAIL.n366 VTAIL.n365 9.3005
R505 VTAIL.n421 VTAIL.n420 9.3005
R506 VTAIL.n423 VTAIL.n422 9.3005
R507 VTAIL.n362 VTAIL.n361 9.3005
R508 VTAIL.n429 VTAIL.n428 9.3005
R509 VTAIL.n407 VTAIL.n406 9.3005
R510 VTAIL.n405 VTAIL.n404 9.3005
R511 VTAIL.n374 VTAIL.n373 9.3005
R512 VTAIL.n399 VTAIL.n398 9.3005
R513 VTAIL.n397 VTAIL.n396 9.3005
R514 VTAIL.n378 VTAIL.n377 9.3005
R515 VTAIL.n391 VTAIL.n390 9.3005
R516 VTAIL.n389 VTAIL.n388 9.3005
R517 VTAIL.n382 VTAIL.n381 9.3005
R518 VTAIL.n298 VTAIL.n297 9.3005
R519 VTAIL.n341 VTAIL.n340 9.3005
R520 VTAIL.n343 VTAIL.n342 9.3005
R521 VTAIL.n294 VTAIL.n293 9.3005
R522 VTAIL.n349 VTAIL.n348 9.3005
R523 VTAIL.n351 VTAIL.n350 9.3005
R524 VTAIL.n290 VTAIL.n289 9.3005
R525 VTAIL.n357 VTAIL.n356 9.3005
R526 VTAIL.n335 VTAIL.n334 9.3005
R527 VTAIL.n333 VTAIL.n332 9.3005
R528 VTAIL.n302 VTAIL.n301 9.3005
R529 VTAIL.n327 VTAIL.n326 9.3005
R530 VTAIL.n325 VTAIL.n324 9.3005
R531 VTAIL.n306 VTAIL.n305 9.3005
R532 VTAIL.n319 VTAIL.n318 9.3005
R533 VTAIL.n317 VTAIL.n316 9.3005
R534 VTAIL.n310 VTAIL.n309 9.3005
R535 VTAIL.n226 VTAIL.n225 9.3005
R536 VTAIL.n269 VTAIL.n268 9.3005
R537 VTAIL.n271 VTAIL.n270 9.3005
R538 VTAIL.n222 VTAIL.n221 9.3005
R539 VTAIL.n277 VTAIL.n276 9.3005
R540 VTAIL.n279 VTAIL.n278 9.3005
R541 VTAIL.n218 VTAIL.n217 9.3005
R542 VTAIL.n285 VTAIL.n284 9.3005
R543 VTAIL.n263 VTAIL.n262 9.3005
R544 VTAIL.n261 VTAIL.n260 9.3005
R545 VTAIL.n230 VTAIL.n229 9.3005
R546 VTAIL.n255 VTAIL.n254 9.3005
R547 VTAIL.n253 VTAIL.n252 9.3005
R548 VTAIL.n234 VTAIL.n233 9.3005
R549 VTAIL.n247 VTAIL.n246 9.3005
R550 VTAIL.n245 VTAIL.n244 9.3005
R551 VTAIL.n238 VTAIL.n237 9.3005
R552 VTAIL.n544 VTAIL.n543 8.92171
R553 VTAIL.n559 VTAIL.n512 8.92171
R554 VTAIL.n40 VTAIL.n39 8.92171
R555 VTAIL.n55 VTAIL.n8 8.92171
R556 VTAIL.n112 VTAIL.n111 8.92171
R557 VTAIL.n127 VTAIL.n80 8.92171
R558 VTAIL.n184 VTAIL.n183 8.92171
R559 VTAIL.n199 VTAIL.n152 8.92171
R560 VTAIL.n487 VTAIL.n440 8.92171
R561 VTAIL.n472 VTAIL.n471 8.92171
R562 VTAIL.n415 VTAIL.n368 8.92171
R563 VTAIL.n400 VTAIL.n399 8.92171
R564 VTAIL.n343 VTAIL.n296 8.92171
R565 VTAIL.n328 VTAIL.n327 8.92171
R566 VTAIL.n271 VTAIL.n224 8.92171
R567 VTAIL.n256 VTAIL.n255 8.92171
R568 VTAIL.n547 VTAIL.n518 8.14595
R569 VTAIL.n556 VTAIL.n555 8.14595
R570 VTAIL.n43 VTAIL.n14 8.14595
R571 VTAIL.n52 VTAIL.n51 8.14595
R572 VTAIL.n115 VTAIL.n86 8.14595
R573 VTAIL.n124 VTAIL.n123 8.14595
R574 VTAIL.n187 VTAIL.n158 8.14595
R575 VTAIL.n196 VTAIL.n195 8.14595
R576 VTAIL.n484 VTAIL.n483 8.14595
R577 VTAIL.n475 VTAIL.n446 8.14595
R578 VTAIL.n412 VTAIL.n411 8.14595
R579 VTAIL.n403 VTAIL.n374 8.14595
R580 VTAIL.n340 VTAIL.n339 8.14595
R581 VTAIL.n331 VTAIL.n302 8.14595
R582 VTAIL.n268 VTAIL.n267 8.14595
R583 VTAIL.n259 VTAIL.n230 8.14595
R584 VTAIL.n574 VTAIL.n504 7.75445
R585 VTAIL.n70 VTAIL.n0 7.75445
R586 VTAIL.n142 VTAIL.n72 7.75445
R587 VTAIL.n214 VTAIL.n144 7.75445
R588 VTAIL.n502 VTAIL.n432 7.75445
R589 VTAIL.n430 VTAIL.n360 7.75445
R590 VTAIL.n358 VTAIL.n288 7.75445
R591 VTAIL.n286 VTAIL.n216 7.75445
R592 VTAIL.n548 VTAIL.n516 7.3702
R593 VTAIL.n552 VTAIL.n514 7.3702
R594 VTAIL.n44 VTAIL.n12 7.3702
R595 VTAIL.n48 VTAIL.n10 7.3702
R596 VTAIL.n116 VTAIL.n84 7.3702
R597 VTAIL.n120 VTAIL.n82 7.3702
R598 VTAIL.n188 VTAIL.n156 7.3702
R599 VTAIL.n192 VTAIL.n154 7.3702
R600 VTAIL.n480 VTAIL.n442 7.3702
R601 VTAIL.n476 VTAIL.n444 7.3702
R602 VTAIL.n408 VTAIL.n370 7.3702
R603 VTAIL.n404 VTAIL.n372 7.3702
R604 VTAIL.n336 VTAIL.n298 7.3702
R605 VTAIL.n332 VTAIL.n300 7.3702
R606 VTAIL.n264 VTAIL.n226 7.3702
R607 VTAIL.n260 VTAIL.n228 7.3702
R608 VTAIL.n551 VTAIL.n516 6.59444
R609 VTAIL.n552 VTAIL.n551 6.59444
R610 VTAIL.n47 VTAIL.n12 6.59444
R611 VTAIL.n48 VTAIL.n47 6.59444
R612 VTAIL.n119 VTAIL.n84 6.59444
R613 VTAIL.n120 VTAIL.n119 6.59444
R614 VTAIL.n191 VTAIL.n156 6.59444
R615 VTAIL.n192 VTAIL.n191 6.59444
R616 VTAIL.n480 VTAIL.n479 6.59444
R617 VTAIL.n479 VTAIL.n444 6.59444
R618 VTAIL.n408 VTAIL.n407 6.59444
R619 VTAIL.n407 VTAIL.n372 6.59444
R620 VTAIL.n336 VTAIL.n335 6.59444
R621 VTAIL.n335 VTAIL.n300 6.59444
R622 VTAIL.n264 VTAIL.n263 6.59444
R623 VTAIL.n263 VTAIL.n228 6.59444
R624 VTAIL.n572 VTAIL.n504 6.08283
R625 VTAIL.n68 VTAIL.n0 6.08283
R626 VTAIL.n140 VTAIL.n72 6.08283
R627 VTAIL.n212 VTAIL.n144 6.08283
R628 VTAIL.n500 VTAIL.n432 6.08283
R629 VTAIL.n428 VTAIL.n360 6.08283
R630 VTAIL.n356 VTAIL.n288 6.08283
R631 VTAIL.n284 VTAIL.n216 6.08283
R632 VTAIL.n548 VTAIL.n547 5.81868
R633 VTAIL.n555 VTAIL.n514 5.81868
R634 VTAIL.n44 VTAIL.n43 5.81868
R635 VTAIL.n51 VTAIL.n10 5.81868
R636 VTAIL.n116 VTAIL.n115 5.81868
R637 VTAIL.n123 VTAIL.n82 5.81868
R638 VTAIL.n188 VTAIL.n187 5.81868
R639 VTAIL.n195 VTAIL.n154 5.81868
R640 VTAIL.n483 VTAIL.n442 5.81868
R641 VTAIL.n476 VTAIL.n475 5.81868
R642 VTAIL.n411 VTAIL.n370 5.81868
R643 VTAIL.n404 VTAIL.n403 5.81868
R644 VTAIL.n339 VTAIL.n298 5.81868
R645 VTAIL.n332 VTAIL.n331 5.81868
R646 VTAIL.n267 VTAIL.n226 5.81868
R647 VTAIL.n260 VTAIL.n259 5.81868
R648 VTAIL.n544 VTAIL.n518 5.04292
R649 VTAIL.n556 VTAIL.n512 5.04292
R650 VTAIL.n40 VTAIL.n14 5.04292
R651 VTAIL.n52 VTAIL.n8 5.04292
R652 VTAIL.n112 VTAIL.n86 5.04292
R653 VTAIL.n124 VTAIL.n80 5.04292
R654 VTAIL.n184 VTAIL.n158 5.04292
R655 VTAIL.n196 VTAIL.n152 5.04292
R656 VTAIL.n484 VTAIL.n440 5.04292
R657 VTAIL.n472 VTAIL.n446 5.04292
R658 VTAIL.n412 VTAIL.n368 5.04292
R659 VTAIL.n400 VTAIL.n374 5.04292
R660 VTAIL.n340 VTAIL.n296 5.04292
R661 VTAIL.n328 VTAIL.n302 5.04292
R662 VTAIL.n268 VTAIL.n224 5.04292
R663 VTAIL.n256 VTAIL.n230 5.04292
R664 VTAIL.n543 VTAIL.n520 4.26717
R665 VTAIL.n560 VTAIL.n559 4.26717
R666 VTAIL.n39 VTAIL.n16 4.26717
R667 VTAIL.n56 VTAIL.n55 4.26717
R668 VTAIL.n111 VTAIL.n88 4.26717
R669 VTAIL.n128 VTAIL.n127 4.26717
R670 VTAIL.n183 VTAIL.n160 4.26717
R671 VTAIL.n200 VTAIL.n199 4.26717
R672 VTAIL.n488 VTAIL.n487 4.26717
R673 VTAIL.n471 VTAIL.n448 4.26717
R674 VTAIL.n416 VTAIL.n415 4.26717
R675 VTAIL.n399 VTAIL.n376 4.26717
R676 VTAIL.n344 VTAIL.n343 4.26717
R677 VTAIL.n327 VTAIL.n304 4.26717
R678 VTAIL.n272 VTAIL.n271 4.26717
R679 VTAIL.n255 VTAIL.n232 4.26717
R680 VTAIL.n527 VTAIL.n525 3.70982
R681 VTAIL.n23 VTAIL.n21 3.70982
R682 VTAIL.n95 VTAIL.n93 3.70982
R683 VTAIL.n167 VTAIL.n165 3.70982
R684 VTAIL.n455 VTAIL.n453 3.70982
R685 VTAIL.n383 VTAIL.n381 3.70982
R686 VTAIL.n311 VTAIL.n309 3.70982
R687 VTAIL.n239 VTAIL.n237 3.70982
R688 VTAIL.n540 VTAIL.n539 3.49141
R689 VTAIL.n563 VTAIL.n510 3.49141
R690 VTAIL.n36 VTAIL.n35 3.49141
R691 VTAIL.n59 VTAIL.n6 3.49141
R692 VTAIL.n108 VTAIL.n107 3.49141
R693 VTAIL.n131 VTAIL.n78 3.49141
R694 VTAIL.n180 VTAIL.n179 3.49141
R695 VTAIL.n203 VTAIL.n150 3.49141
R696 VTAIL.n491 VTAIL.n438 3.49141
R697 VTAIL.n468 VTAIL.n467 3.49141
R698 VTAIL.n419 VTAIL.n366 3.49141
R699 VTAIL.n396 VTAIL.n395 3.49141
R700 VTAIL.n347 VTAIL.n294 3.49141
R701 VTAIL.n324 VTAIL.n323 3.49141
R702 VTAIL.n275 VTAIL.n222 3.49141
R703 VTAIL.n252 VTAIL.n251 3.49141
R704 VTAIL.n536 VTAIL.n522 2.71565
R705 VTAIL.n564 VTAIL.n508 2.71565
R706 VTAIL.n32 VTAIL.n18 2.71565
R707 VTAIL.n60 VTAIL.n4 2.71565
R708 VTAIL.n104 VTAIL.n90 2.71565
R709 VTAIL.n132 VTAIL.n76 2.71565
R710 VTAIL.n176 VTAIL.n162 2.71565
R711 VTAIL.n204 VTAIL.n148 2.71565
R712 VTAIL.n492 VTAIL.n436 2.71565
R713 VTAIL.n464 VTAIL.n450 2.71565
R714 VTAIL.n420 VTAIL.n364 2.71565
R715 VTAIL.n392 VTAIL.n378 2.71565
R716 VTAIL.n348 VTAIL.n292 2.71565
R717 VTAIL.n320 VTAIL.n306 2.71565
R718 VTAIL.n276 VTAIL.n220 2.71565
R719 VTAIL.n248 VTAIL.n234 2.71565
R720 VTAIL.n535 VTAIL.n524 1.93989
R721 VTAIL.n568 VTAIL.n567 1.93989
R722 VTAIL.n31 VTAIL.n20 1.93989
R723 VTAIL.n64 VTAIL.n63 1.93989
R724 VTAIL.n103 VTAIL.n92 1.93989
R725 VTAIL.n136 VTAIL.n135 1.93989
R726 VTAIL.n175 VTAIL.n164 1.93989
R727 VTAIL.n208 VTAIL.n207 1.93989
R728 VTAIL.n496 VTAIL.n495 1.93989
R729 VTAIL.n463 VTAIL.n452 1.93989
R730 VTAIL.n424 VTAIL.n423 1.93989
R731 VTAIL.n391 VTAIL.n380 1.93989
R732 VTAIL.n352 VTAIL.n351 1.93989
R733 VTAIL.n319 VTAIL.n308 1.93989
R734 VTAIL.n280 VTAIL.n279 1.93989
R735 VTAIL.n247 VTAIL.n236 1.93989
R736 VTAIL.n359 VTAIL.n287 1.69878
R737 VTAIL.n503 VTAIL.n431 1.69878
R738 VTAIL.n215 VTAIL.n143 1.69878
R739 VTAIL.n532 VTAIL.n531 1.16414
R740 VTAIL.n571 VTAIL.n506 1.16414
R741 VTAIL.n28 VTAIL.n27 1.16414
R742 VTAIL.n67 VTAIL.n2 1.16414
R743 VTAIL.n100 VTAIL.n99 1.16414
R744 VTAIL.n139 VTAIL.n74 1.16414
R745 VTAIL.n172 VTAIL.n171 1.16414
R746 VTAIL.n211 VTAIL.n146 1.16414
R747 VTAIL.n499 VTAIL.n434 1.16414
R748 VTAIL.n460 VTAIL.n459 1.16414
R749 VTAIL.n427 VTAIL.n362 1.16414
R750 VTAIL.n388 VTAIL.n387 1.16414
R751 VTAIL.n355 VTAIL.n290 1.16414
R752 VTAIL.n316 VTAIL.n315 1.16414
R753 VTAIL.n283 VTAIL.n218 1.16414
R754 VTAIL.n244 VTAIL.n243 1.16414
R755 VTAIL VTAIL.n71 0.907828
R756 VTAIL VTAIL.n575 0.791448
R757 VTAIL.n431 VTAIL.n359 0.470328
R758 VTAIL.n143 VTAIL.n71 0.470328
R759 VTAIL.n528 VTAIL.n526 0.388379
R760 VTAIL.n24 VTAIL.n22 0.388379
R761 VTAIL.n96 VTAIL.n94 0.388379
R762 VTAIL.n168 VTAIL.n166 0.388379
R763 VTAIL.n456 VTAIL.n454 0.388379
R764 VTAIL.n384 VTAIL.n382 0.388379
R765 VTAIL.n312 VTAIL.n310 0.388379
R766 VTAIL.n240 VTAIL.n238 0.388379
R767 VTAIL.n533 VTAIL.n525 0.155672
R768 VTAIL.n534 VTAIL.n533 0.155672
R769 VTAIL.n534 VTAIL.n521 0.155672
R770 VTAIL.n541 VTAIL.n521 0.155672
R771 VTAIL.n542 VTAIL.n541 0.155672
R772 VTAIL.n542 VTAIL.n517 0.155672
R773 VTAIL.n549 VTAIL.n517 0.155672
R774 VTAIL.n550 VTAIL.n549 0.155672
R775 VTAIL.n550 VTAIL.n513 0.155672
R776 VTAIL.n557 VTAIL.n513 0.155672
R777 VTAIL.n558 VTAIL.n557 0.155672
R778 VTAIL.n558 VTAIL.n509 0.155672
R779 VTAIL.n565 VTAIL.n509 0.155672
R780 VTAIL.n566 VTAIL.n565 0.155672
R781 VTAIL.n566 VTAIL.n505 0.155672
R782 VTAIL.n573 VTAIL.n505 0.155672
R783 VTAIL.n29 VTAIL.n21 0.155672
R784 VTAIL.n30 VTAIL.n29 0.155672
R785 VTAIL.n30 VTAIL.n17 0.155672
R786 VTAIL.n37 VTAIL.n17 0.155672
R787 VTAIL.n38 VTAIL.n37 0.155672
R788 VTAIL.n38 VTAIL.n13 0.155672
R789 VTAIL.n45 VTAIL.n13 0.155672
R790 VTAIL.n46 VTAIL.n45 0.155672
R791 VTAIL.n46 VTAIL.n9 0.155672
R792 VTAIL.n53 VTAIL.n9 0.155672
R793 VTAIL.n54 VTAIL.n53 0.155672
R794 VTAIL.n54 VTAIL.n5 0.155672
R795 VTAIL.n61 VTAIL.n5 0.155672
R796 VTAIL.n62 VTAIL.n61 0.155672
R797 VTAIL.n62 VTAIL.n1 0.155672
R798 VTAIL.n69 VTAIL.n1 0.155672
R799 VTAIL.n101 VTAIL.n93 0.155672
R800 VTAIL.n102 VTAIL.n101 0.155672
R801 VTAIL.n102 VTAIL.n89 0.155672
R802 VTAIL.n109 VTAIL.n89 0.155672
R803 VTAIL.n110 VTAIL.n109 0.155672
R804 VTAIL.n110 VTAIL.n85 0.155672
R805 VTAIL.n117 VTAIL.n85 0.155672
R806 VTAIL.n118 VTAIL.n117 0.155672
R807 VTAIL.n118 VTAIL.n81 0.155672
R808 VTAIL.n125 VTAIL.n81 0.155672
R809 VTAIL.n126 VTAIL.n125 0.155672
R810 VTAIL.n126 VTAIL.n77 0.155672
R811 VTAIL.n133 VTAIL.n77 0.155672
R812 VTAIL.n134 VTAIL.n133 0.155672
R813 VTAIL.n134 VTAIL.n73 0.155672
R814 VTAIL.n141 VTAIL.n73 0.155672
R815 VTAIL.n173 VTAIL.n165 0.155672
R816 VTAIL.n174 VTAIL.n173 0.155672
R817 VTAIL.n174 VTAIL.n161 0.155672
R818 VTAIL.n181 VTAIL.n161 0.155672
R819 VTAIL.n182 VTAIL.n181 0.155672
R820 VTAIL.n182 VTAIL.n157 0.155672
R821 VTAIL.n189 VTAIL.n157 0.155672
R822 VTAIL.n190 VTAIL.n189 0.155672
R823 VTAIL.n190 VTAIL.n153 0.155672
R824 VTAIL.n197 VTAIL.n153 0.155672
R825 VTAIL.n198 VTAIL.n197 0.155672
R826 VTAIL.n198 VTAIL.n149 0.155672
R827 VTAIL.n205 VTAIL.n149 0.155672
R828 VTAIL.n206 VTAIL.n205 0.155672
R829 VTAIL.n206 VTAIL.n145 0.155672
R830 VTAIL.n213 VTAIL.n145 0.155672
R831 VTAIL.n501 VTAIL.n433 0.155672
R832 VTAIL.n494 VTAIL.n433 0.155672
R833 VTAIL.n494 VTAIL.n493 0.155672
R834 VTAIL.n493 VTAIL.n437 0.155672
R835 VTAIL.n486 VTAIL.n437 0.155672
R836 VTAIL.n486 VTAIL.n485 0.155672
R837 VTAIL.n485 VTAIL.n441 0.155672
R838 VTAIL.n478 VTAIL.n441 0.155672
R839 VTAIL.n478 VTAIL.n477 0.155672
R840 VTAIL.n477 VTAIL.n445 0.155672
R841 VTAIL.n470 VTAIL.n445 0.155672
R842 VTAIL.n470 VTAIL.n469 0.155672
R843 VTAIL.n469 VTAIL.n449 0.155672
R844 VTAIL.n462 VTAIL.n449 0.155672
R845 VTAIL.n462 VTAIL.n461 0.155672
R846 VTAIL.n461 VTAIL.n453 0.155672
R847 VTAIL.n429 VTAIL.n361 0.155672
R848 VTAIL.n422 VTAIL.n361 0.155672
R849 VTAIL.n422 VTAIL.n421 0.155672
R850 VTAIL.n421 VTAIL.n365 0.155672
R851 VTAIL.n414 VTAIL.n365 0.155672
R852 VTAIL.n414 VTAIL.n413 0.155672
R853 VTAIL.n413 VTAIL.n369 0.155672
R854 VTAIL.n406 VTAIL.n369 0.155672
R855 VTAIL.n406 VTAIL.n405 0.155672
R856 VTAIL.n405 VTAIL.n373 0.155672
R857 VTAIL.n398 VTAIL.n373 0.155672
R858 VTAIL.n398 VTAIL.n397 0.155672
R859 VTAIL.n397 VTAIL.n377 0.155672
R860 VTAIL.n390 VTAIL.n377 0.155672
R861 VTAIL.n390 VTAIL.n389 0.155672
R862 VTAIL.n389 VTAIL.n381 0.155672
R863 VTAIL.n357 VTAIL.n289 0.155672
R864 VTAIL.n350 VTAIL.n289 0.155672
R865 VTAIL.n350 VTAIL.n349 0.155672
R866 VTAIL.n349 VTAIL.n293 0.155672
R867 VTAIL.n342 VTAIL.n293 0.155672
R868 VTAIL.n342 VTAIL.n341 0.155672
R869 VTAIL.n341 VTAIL.n297 0.155672
R870 VTAIL.n334 VTAIL.n297 0.155672
R871 VTAIL.n334 VTAIL.n333 0.155672
R872 VTAIL.n333 VTAIL.n301 0.155672
R873 VTAIL.n326 VTAIL.n301 0.155672
R874 VTAIL.n326 VTAIL.n325 0.155672
R875 VTAIL.n325 VTAIL.n305 0.155672
R876 VTAIL.n318 VTAIL.n305 0.155672
R877 VTAIL.n318 VTAIL.n317 0.155672
R878 VTAIL.n317 VTAIL.n309 0.155672
R879 VTAIL.n285 VTAIL.n217 0.155672
R880 VTAIL.n278 VTAIL.n217 0.155672
R881 VTAIL.n278 VTAIL.n277 0.155672
R882 VTAIL.n277 VTAIL.n221 0.155672
R883 VTAIL.n270 VTAIL.n221 0.155672
R884 VTAIL.n270 VTAIL.n269 0.155672
R885 VTAIL.n269 VTAIL.n225 0.155672
R886 VTAIL.n262 VTAIL.n225 0.155672
R887 VTAIL.n262 VTAIL.n261 0.155672
R888 VTAIL.n261 VTAIL.n229 0.155672
R889 VTAIL.n254 VTAIL.n229 0.155672
R890 VTAIL.n254 VTAIL.n253 0.155672
R891 VTAIL.n253 VTAIL.n233 0.155672
R892 VTAIL.n246 VTAIL.n233 0.155672
R893 VTAIL.n246 VTAIL.n245 0.155672
R894 VTAIL.n245 VTAIL.n237 0.155672
R895 VDD1 VDD1.n1 114.706
R896 VDD1 VDD1.n0 73.964
R897 VDD1.n0 VDD1.t1 2.44448
R898 VDD1.n0 VDD1.t2 2.44448
R899 VDD1.n1 VDD1.t0 2.44448
R900 VDD1.n1 VDD1.t3 2.44448
R901 B.n348 B.n95 585
R902 B.n347 B.n346 585
R903 B.n345 B.n96 585
R904 B.n344 B.n343 585
R905 B.n342 B.n97 585
R906 B.n341 B.n340 585
R907 B.n339 B.n98 585
R908 B.n338 B.n337 585
R909 B.n336 B.n99 585
R910 B.n335 B.n334 585
R911 B.n333 B.n100 585
R912 B.n332 B.n331 585
R913 B.n330 B.n101 585
R914 B.n329 B.n328 585
R915 B.n327 B.n102 585
R916 B.n326 B.n325 585
R917 B.n324 B.n103 585
R918 B.n323 B.n322 585
R919 B.n321 B.n104 585
R920 B.n320 B.n319 585
R921 B.n318 B.n105 585
R922 B.n317 B.n316 585
R923 B.n315 B.n106 585
R924 B.n314 B.n313 585
R925 B.n312 B.n107 585
R926 B.n311 B.n310 585
R927 B.n309 B.n108 585
R928 B.n308 B.n307 585
R929 B.n306 B.n109 585
R930 B.n305 B.n304 585
R931 B.n303 B.n110 585
R932 B.n302 B.n301 585
R933 B.n300 B.n111 585
R934 B.n299 B.n298 585
R935 B.n297 B.n112 585
R936 B.n296 B.n295 585
R937 B.n294 B.n113 585
R938 B.n293 B.n292 585
R939 B.n291 B.n114 585
R940 B.n290 B.n289 585
R941 B.n288 B.n115 585
R942 B.n287 B.n286 585
R943 B.n285 B.n116 585
R944 B.n284 B.n283 585
R945 B.n282 B.n117 585
R946 B.n280 B.n279 585
R947 B.n278 B.n120 585
R948 B.n277 B.n276 585
R949 B.n275 B.n121 585
R950 B.n274 B.n273 585
R951 B.n272 B.n122 585
R952 B.n271 B.n270 585
R953 B.n269 B.n123 585
R954 B.n268 B.n267 585
R955 B.n266 B.n124 585
R956 B.n265 B.n264 585
R957 B.n260 B.n125 585
R958 B.n259 B.n258 585
R959 B.n257 B.n126 585
R960 B.n256 B.n255 585
R961 B.n254 B.n127 585
R962 B.n253 B.n252 585
R963 B.n251 B.n128 585
R964 B.n250 B.n249 585
R965 B.n248 B.n129 585
R966 B.n247 B.n246 585
R967 B.n245 B.n130 585
R968 B.n244 B.n243 585
R969 B.n242 B.n131 585
R970 B.n241 B.n240 585
R971 B.n239 B.n132 585
R972 B.n238 B.n237 585
R973 B.n236 B.n133 585
R974 B.n235 B.n234 585
R975 B.n233 B.n134 585
R976 B.n232 B.n231 585
R977 B.n230 B.n135 585
R978 B.n229 B.n228 585
R979 B.n227 B.n136 585
R980 B.n226 B.n225 585
R981 B.n224 B.n137 585
R982 B.n223 B.n222 585
R983 B.n221 B.n138 585
R984 B.n220 B.n219 585
R985 B.n218 B.n139 585
R986 B.n217 B.n216 585
R987 B.n215 B.n140 585
R988 B.n214 B.n213 585
R989 B.n212 B.n141 585
R990 B.n211 B.n210 585
R991 B.n209 B.n142 585
R992 B.n208 B.n207 585
R993 B.n206 B.n143 585
R994 B.n205 B.n204 585
R995 B.n203 B.n144 585
R996 B.n202 B.n201 585
R997 B.n200 B.n145 585
R998 B.n199 B.n198 585
R999 B.n197 B.n146 585
R1000 B.n196 B.n195 585
R1001 B.n350 B.n349 585
R1002 B.n351 B.n94 585
R1003 B.n353 B.n352 585
R1004 B.n354 B.n93 585
R1005 B.n356 B.n355 585
R1006 B.n357 B.n92 585
R1007 B.n359 B.n358 585
R1008 B.n360 B.n91 585
R1009 B.n362 B.n361 585
R1010 B.n363 B.n90 585
R1011 B.n365 B.n364 585
R1012 B.n366 B.n89 585
R1013 B.n368 B.n367 585
R1014 B.n369 B.n88 585
R1015 B.n371 B.n370 585
R1016 B.n372 B.n87 585
R1017 B.n374 B.n373 585
R1018 B.n375 B.n86 585
R1019 B.n377 B.n376 585
R1020 B.n378 B.n85 585
R1021 B.n380 B.n379 585
R1022 B.n381 B.n84 585
R1023 B.n383 B.n382 585
R1024 B.n384 B.n83 585
R1025 B.n386 B.n385 585
R1026 B.n387 B.n82 585
R1027 B.n389 B.n388 585
R1028 B.n390 B.n81 585
R1029 B.n392 B.n391 585
R1030 B.n393 B.n80 585
R1031 B.n395 B.n394 585
R1032 B.n396 B.n79 585
R1033 B.n398 B.n397 585
R1034 B.n399 B.n78 585
R1035 B.n401 B.n400 585
R1036 B.n402 B.n77 585
R1037 B.n404 B.n403 585
R1038 B.n405 B.n76 585
R1039 B.n407 B.n406 585
R1040 B.n408 B.n75 585
R1041 B.n410 B.n409 585
R1042 B.n411 B.n74 585
R1043 B.n413 B.n412 585
R1044 B.n414 B.n73 585
R1045 B.n416 B.n415 585
R1046 B.n417 B.n72 585
R1047 B.n419 B.n418 585
R1048 B.n420 B.n71 585
R1049 B.n422 B.n421 585
R1050 B.n423 B.n70 585
R1051 B.n425 B.n424 585
R1052 B.n426 B.n69 585
R1053 B.n578 B.n577 585
R1054 B.n576 B.n15 585
R1055 B.n575 B.n574 585
R1056 B.n573 B.n16 585
R1057 B.n572 B.n571 585
R1058 B.n570 B.n17 585
R1059 B.n569 B.n568 585
R1060 B.n567 B.n18 585
R1061 B.n566 B.n565 585
R1062 B.n564 B.n19 585
R1063 B.n563 B.n562 585
R1064 B.n561 B.n20 585
R1065 B.n560 B.n559 585
R1066 B.n558 B.n21 585
R1067 B.n557 B.n556 585
R1068 B.n555 B.n22 585
R1069 B.n554 B.n553 585
R1070 B.n552 B.n23 585
R1071 B.n551 B.n550 585
R1072 B.n549 B.n24 585
R1073 B.n548 B.n547 585
R1074 B.n546 B.n25 585
R1075 B.n545 B.n544 585
R1076 B.n543 B.n26 585
R1077 B.n542 B.n541 585
R1078 B.n540 B.n27 585
R1079 B.n539 B.n538 585
R1080 B.n537 B.n28 585
R1081 B.n536 B.n535 585
R1082 B.n534 B.n29 585
R1083 B.n533 B.n532 585
R1084 B.n531 B.n30 585
R1085 B.n530 B.n529 585
R1086 B.n528 B.n31 585
R1087 B.n527 B.n526 585
R1088 B.n525 B.n32 585
R1089 B.n524 B.n523 585
R1090 B.n522 B.n33 585
R1091 B.n521 B.n520 585
R1092 B.n519 B.n34 585
R1093 B.n518 B.n517 585
R1094 B.n516 B.n35 585
R1095 B.n515 B.n514 585
R1096 B.n513 B.n36 585
R1097 B.n512 B.n511 585
R1098 B.n509 B.n37 585
R1099 B.n508 B.n507 585
R1100 B.n506 B.n40 585
R1101 B.n505 B.n504 585
R1102 B.n503 B.n41 585
R1103 B.n502 B.n501 585
R1104 B.n500 B.n42 585
R1105 B.n499 B.n498 585
R1106 B.n497 B.n43 585
R1107 B.n496 B.n495 585
R1108 B.n494 B.n493 585
R1109 B.n492 B.n47 585
R1110 B.n491 B.n490 585
R1111 B.n489 B.n48 585
R1112 B.n488 B.n487 585
R1113 B.n486 B.n49 585
R1114 B.n485 B.n484 585
R1115 B.n483 B.n50 585
R1116 B.n482 B.n481 585
R1117 B.n480 B.n51 585
R1118 B.n479 B.n478 585
R1119 B.n477 B.n52 585
R1120 B.n476 B.n475 585
R1121 B.n474 B.n53 585
R1122 B.n473 B.n472 585
R1123 B.n471 B.n54 585
R1124 B.n470 B.n469 585
R1125 B.n468 B.n55 585
R1126 B.n467 B.n466 585
R1127 B.n465 B.n56 585
R1128 B.n464 B.n463 585
R1129 B.n462 B.n57 585
R1130 B.n461 B.n460 585
R1131 B.n459 B.n58 585
R1132 B.n458 B.n457 585
R1133 B.n456 B.n59 585
R1134 B.n455 B.n454 585
R1135 B.n453 B.n60 585
R1136 B.n452 B.n451 585
R1137 B.n450 B.n61 585
R1138 B.n449 B.n448 585
R1139 B.n447 B.n62 585
R1140 B.n446 B.n445 585
R1141 B.n444 B.n63 585
R1142 B.n443 B.n442 585
R1143 B.n441 B.n64 585
R1144 B.n440 B.n439 585
R1145 B.n438 B.n65 585
R1146 B.n437 B.n436 585
R1147 B.n435 B.n66 585
R1148 B.n434 B.n433 585
R1149 B.n432 B.n67 585
R1150 B.n431 B.n430 585
R1151 B.n429 B.n68 585
R1152 B.n428 B.n427 585
R1153 B.n579 B.n14 585
R1154 B.n581 B.n580 585
R1155 B.n582 B.n13 585
R1156 B.n584 B.n583 585
R1157 B.n585 B.n12 585
R1158 B.n587 B.n586 585
R1159 B.n588 B.n11 585
R1160 B.n590 B.n589 585
R1161 B.n591 B.n10 585
R1162 B.n593 B.n592 585
R1163 B.n594 B.n9 585
R1164 B.n596 B.n595 585
R1165 B.n597 B.n8 585
R1166 B.n599 B.n598 585
R1167 B.n600 B.n7 585
R1168 B.n602 B.n601 585
R1169 B.n603 B.n6 585
R1170 B.n605 B.n604 585
R1171 B.n606 B.n5 585
R1172 B.n608 B.n607 585
R1173 B.n609 B.n4 585
R1174 B.n611 B.n610 585
R1175 B.n612 B.n3 585
R1176 B.n614 B.n613 585
R1177 B.n615 B.n0 585
R1178 B.n2 B.n1 585
R1179 B.n160 B.n159 585
R1180 B.n161 B.n158 585
R1181 B.n163 B.n162 585
R1182 B.n164 B.n157 585
R1183 B.n166 B.n165 585
R1184 B.n167 B.n156 585
R1185 B.n169 B.n168 585
R1186 B.n170 B.n155 585
R1187 B.n172 B.n171 585
R1188 B.n173 B.n154 585
R1189 B.n175 B.n174 585
R1190 B.n176 B.n153 585
R1191 B.n178 B.n177 585
R1192 B.n179 B.n152 585
R1193 B.n181 B.n180 585
R1194 B.n182 B.n151 585
R1195 B.n184 B.n183 585
R1196 B.n185 B.n150 585
R1197 B.n187 B.n186 585
R1198 B.n188 B.n149 585
R1199 B.n190 B.n189 585
R1200 B.n191 B.n148 585
R1201 B.n193 B.n192 585
R1202 B.n194 B.n147 585
R1203 B.n196 B.n147 535.745
R1204 B.n350 B.n95 535.745
R1205 B.n428 B.n69 535.745
R1206 B.n579 B.n578 535.745
R1207 B.n118 B.t7 437.067
R1208 B.n44 B.t11 437.067
R1209 B.n261 B.t4 437.067
R1210 B.n38 B.t2 437.067
R1211 B.n261 B.t3 401.37
R1212 B.n118 B.t6 401.37
R1213 B.n44 B.t9 401.37
R1214 B.n38 B.t0 401.37
R1215 B.n119 B.t8 398.861
R1216 B.n45 B.t10 398.861
R1217 B.n262 B.t5 398.861
R1218 B.n39 B.t1 398.861
R1219 B.n617 B.n616 256.663
R1220 B.n616 B.n615 235.042
R1221 B.n616 B.n2 235.042
R1222 B.n197 B.n196 163.367
R1223 B.n198 B.n197 163.367
R1224 B.n198 B.n145 163.367
R1225 B.n202 B.n145 163.367
R1226 B.n203 B.n202 163.367
R1227 B.n204 B.n203 163.367
R1228 B.n204 B.n143 163.367
R1229 B.n208 B.n143 163.367
R1230 B.n209 B.n208 163.367
R1231 B.n210 B.n209 163.367
R1232 B.n210 B.n141 163.367
R1233 B.n214 B.n141 163.367
R1234 B.n215 B.n214 163.367
R1235 B.n216 B.n215 163.367
R1236 B.n216 B.n139 163.367
R1237 B.n220 B.n139 163.367
R1238 B.n221 B.n220 163.367
R1239 B.n222 B.n221 163.367
R1240 B.n222 B.n137 163.367
R1241 B.n226 B.n137 163.367
R1242 B.n227 B.n226 163.367
R1243 B.n228 B.n227 163.367
R1244 B.n228 B.n135 163.367
R1245 B.n232 B.n135 163.367
R1246 B.n233 B.n232 163.367
R1247 B.n234 B.n233 163.367
R1248 B.n234 B.n133 163.367
R1249 B.n238 B.n133 163.367
R1250 B.n239 B.n238 163.367
R1251 B.n240 B.n239 163.367
R1252 B.n240 B.n131 163.367
R1253 B.n244 B.n131 163.367
R1254 B.n245 B.n244 163.367
R1255 B.n246 B.n245 163.367
R1256 B.n246 B.n129 163.367
R1257 B.n250 B.n129 163.367
R1258 B.n251 B.n250 163.367
R1259 B.n252 B.n251 163.367
R1260 B.n252 B.n127 163.367
R1261 B.n256 B.n127 163.367
R1262 B.n257 B.n256 163.367
R1263 B.n258 B.n257 163.367
R1264 B.n258 B.n125 163.367
R1265 B.n265 B.n125 163.367
R1266 B.n266 B.n265 163.367
R1267 B.n267 B.n266 163.367
R1268 B.n267 B.n123 163.367
R1269 B.n271 B.n123 163.367
R1270 B.n272 B.n271 163.367
R1271 B.n273 B.n272 163.367
R1272 B.n273 B.n121 163.367
R1273 B.n277 B.n121 163.367
R1274 B.n278 B.n277 163.367
R1275 B.n279 B.n278 163.367
R1276 B.n279 B.n117 163.367
R1277 B.n284 B.n117 163.367
R1278 B.n285 B.n284 163.367
R1279 B.n286 B.n285 163.367
R1280 B.n286 B.n115 163.367
R1281 B.n290 B.n115 163.367
R1282 B.n291 B.n290 163.367
R1283 B.n292 B.n291 163.367
R1284 B.n292 B.n113 163.367
R1285 B.n296 B.n113 163.367
R1286 B.n297 B.n296 163.367
R1287 B.n298 B.n297 163.367
R1288 B.n298 B.n111 163.367
R1289 B.n302 B.n111 163.367
R1290 B.n303 B.n302 163.367
R1291 B.n304 B.n303 163.367
R1292 B.n304 B.n109 163.367
R1293 B.n308 B.n109 163.367
R1294 B.n309 B.n308 163.367
R1295 B.n310 B.n309 163.367
R1296 B.n310 B.n107 163.367
R1297 B.n314 B.n107 163.367
R1298 B.n315 B.n314 163.367
R1299 B.n316 B.n315 163.367
R1300 B.n316 B.n105 163.367
R1301 B.n320 B.n105 163.367
R1302 B.n321 B.n320 163.367
R1303 B.n322 B.n321 163.367
R1304 B.n322 B.n103 163.367
R1305 B.n326 B.n103 163.367
R1306 B.n327 B.n326 163.367
R1307 B.n328 B.n327 163.367
R1308 B.n328 B.n101 163.367
R1309 B.n332 B.n101 163.367
R1310 B.n333 B.n332 163.367
R1311 B.n334 B.n333 163.367
R1312 B.n334 B.n99 163.367
R1313 B.n338 B.n99 163.367
R1314 B.n339 B.n338 163.367
R1315 B.n340 B.n339 163.367
R1316 B.n340 B.n97 163.367
R1317 B.n344 B.n97 163.367
R1318 B.n345 B.n344 163.367
R1319 B.n346 B.n345 163.367
R1320 B.n346 B.n95 163.367
R1321 B.n424 B.n69 163.367
R1322 B.n424 B.n423 163.367
R1323 B.n423 B.n422 163.367
R1324 B.n422 B.n71 163.367
R1325 B.n418 B.n71 163.367
R1326 B.n418 B.n417 163.367
R1327 B.n417 B.n416 163.367
R1328 B.n416 B.n73 163.367
R1329 B.n412 B.n73 163.367
R1330 B.n412 B.n411 163.367
R1331 B.n411 B.n410 163.367
R1332 B.n410 B.n75 163.367
R1333 B.n406 B.n75 163.367
R1334 B.n406 B.n405 163.367
R1335 B.n405 B.n404 163.367
R1336 B.n404 B.n77 163.367
R1337 B.n400 B.n77 163.367
R1338 B.n400 B.n399 163.367
R1339 B.n399 B.n398 163.367
R1340 B.n398 B.n79 163.367
R1341 B.n394 B.n79 163.367
R1342 B.n394 B.n393 163.367
R1343 B.n393 B.n392 163.367
R1344 B.n392 B.n81 163.367
R1345 B.n388 B.n81 163.367
R1346 B.n388 B.n387 163.367
R1347 B.n387 B.n386 163.367
R1348 B.n386 B.n83 163.367
R1349 B.n382 B.n83 163.367
R1350 B.n382 B.n381 163.367
R1351 B.n381 B.n380 163.367
R1352 B.n380 B.n85 163.367
R1353 B.n376 B.n85 163.367
R1354 B.n376 B.n375 163.367
R1355 B.n375 B.n374 163.367
R1356 B.n374 B.n87 163.367
R1357 B.n370 B.n87 163.367
R1358 B.n370 B.n369 163.367
R1359 B.n369 B.n368 163.367
R1360 B.n368 B.n89 163.367
R1361 B.n364 B.n89 163.367
R1362 B.n364 B.n363 163.367
R1363 B.n363 B.n362 163.367
R1364 B.n362 B.n91 163.367
R1365 B.n358 B.n91 163.367
R1366 B.n358 B.n357 163.367
R1367 B.n357 B.n356 163.367
R1368 B.n356 B.n93 163.367
R1369 B.n352 B.n93 163.367
R1370 B.n352 B.n351 163.367
R1371 B.n351 B.n350 163.367
R1372 B.n578 B.n15 163.367
R1373 B.n574 B.n15 163.367
R1374 B.n574 B.n573 163.367
R1375 B.n573 B.n572 163.367
R1376 B.n572 B.n17 163.367
R1377 B.n568 B.n17 163.367
R1378 B.n568 B.n567 163.367
R1379 B.n567 B.n566 163.367
R1380 B.n566 B.n19 163.367
R1381 B.n562 B.n19 163.367
R1382 B.n562 B.n561 163.367
R1383 B.n561 B.n560 163.367
R1384 B.n560 B.n21 163.367
R1385 B.n556 B.n21 163.367
R1386 B.n556 B.n555 163.367
R1387 B.n555 B.n554 163.367
R1388 B.n554 B.n23 163.367
R1389 B.n550 B.n23 163.367
R1390 B.n550 B.n549 163.367
R1391 B.n549 B.n548 163.367
R1392 B.n548 B.n25 163.367
R1393 B.n544 B.n25 163.367
R1394 B.n544 B.n543 163.367
R1395 B.n543 B.n542 163.367
R1396 B.n542 B.n27 163.367
R1397 B.n538 B.n27 163.367
R1398 B.n538 B.n537 163.367
R1399 B.n537 B.n536 163.367
R1400 B.n536 B.n29 163.367
R1401 B.n532 B.n29 163.367
R1402 B.n532 B.n531 163.367
R1403 B.n531 B.n530 163.367
R1404 B.n530 B.n31 163.367
R1405 B.n526 B.n31 163.367
R1406 B.n526 B.n525 163.367
R1407 B.n525 B.n524 163.367
R1408 B.n524 B.n33 163.367
R1409 B.n520 B.n33 163.367
R1410 B.n520 B.n519 163.367
R1411 B.n519 B.n518 163.367
R1412 B.n518 B.n35 163.367
R1413 B.n514 B.n35 163.367
R1414 B.n514 B.n513 163.367
R1415 B.n513 B.n512 163.367
R1416 B.n512 B.n37 163.367
R1417 B.n507 B.n37 163.367
R1418 B.n507 B.n506 163.367
R1419 B.n506 B.n505 163.367
R1420 B.n505 B.n41 163.367
R1421 B.n501 B.n41 163.367
R1422 B.n501 B.n500 163.367
R1423 B.n500 B.n499 163.367
R1424 B.n499 B.n43 163.367
R1425 B.n495 B.n43 163.367
R1426 B.n495 B.n494 163.367
R1427 B.n494 B.n47 163.367
R1428 B.n490 B.n47 163.367
R1429 B.n490 B.n489 163.367
R1430 B.n489 B.n488 163.367
R1431 B.n488 B.n49 163.367
R1432 B.n484 B.n49 163.367
R1433 B.n484 B.n483 163.367
R1434 B.n483 B.n482 163.367
R1435 B.n482 B.n51 163.367
R1436 B.n478 B.n51 163.367
R1437 B.n478 B.n477 163.367
R1438 B.n477 B.n476 163.367
R1439 B.n476 B.n53 163.367
R1440 B.n472 B.n53 163.367
R1441 B.n472 B.n471 163.367
R1442 B.n471 B.n470 163.367
R1443 B.n470 B.n55 163.367
R1444 B.n466 B.n55 163.367
R1445 B.n466 B.n465 163.367
R1446 B.n465 B.n464 163.367
R1447 B.n464 B.n57 163.367
R1448 B.n460 B.n57 163.367
R1449 B.n460 B.n459 163.367
R1450 B.n459 B.n458 163.367
R1451 B.n458 B.n59 163.367
R1452 B.n454 B.n59 163.367
R1453 B.n454 B.n453 163.367
R1454 B.n453 B.n452 163.367
R1455 B.n452 B.n61 163.367
R1456 B.n448 B.n61 163.367
R1457 B.n448 B.n447 163.367
R1458 B.n447 B.n446 163.367
R1459 B.n446 B.n63 163.367
R1460 B.n442 B.n63 163.367
R1461 B.n442 B.n441 163.367
R1462 B.n441 B.n440 163.367
R1463 B.n440 B.n65 163.367
R1464 B.n436 B.n65 163.367
R1465 B.n436 B.n435 163.367
R1466 B.n435 B.n434 163.367
R1467 B.n434 B.n67 163.367
R1468 B.n430 B.n67 163.367
R1469 B.n430 B.n429 163.367
R1470 B.n429 B.n428 163.367
R1471 B.n580 B.n579 163.367
R1472 B.n580 B.n13 163.367
R1473 B.n584 B.n13 163.367
R1474 B.n585 B.n584 163.367
R1475 B.n586 B.n585 163.367
R1476 B.n586 B.n11 163.367
R1477 B.n590 B.n11 163.367
R1478 B.n591 B.n590 163.367
R1479 B.n592 B.n591 163.367
R1480 B.n592 B.n9 163.367
R1481 B.n596 B.n9 163.367
R1482 B.n597 B.n596 163.367
R1483 B.n598 B.n597 163.367
R1484 B.n598 B.n7 163.367
R1485 B.n602 B.n7 163.367
R1486 B.n603 B.n602 163.367
R1487 B.n604 B.n603 163.367
R1488 B.n604 B.n5 163.367
R1489 B.n608 B.n5 163.367
R1490 B.n609 B.n608 163.367
R1491 B.n610 B.n609 163.367
R1492 B.n610 B.n3 163.367
R1493 B.n614 B.n3 163.367
R1494 B.n615 B.n614 163.367
R1495 B.n160 B.n2 163.367
R1496 B.n161 B.n160 163.367
R1497 B.n162 B.n161 163.367
R1498 B.n162 B.n157 163.367
R1499 B.n166 B.n157 163.367
R1500 B.n167 B.n166 163.367
R1501 B.n168 B.n167 163.367
R1502 B.n168 B.n155 163.367
R1503 B.n172 B.n155 163.367
R1504 B.n173 B.n172 163.367
R1505 B.n174 B.n173 163.367
R1506 B.n174 B.n153 163.367
R1507 B.n178 B.n153 163.367
R1508 B.n179 B.n178 163.367
R1509 B.n180 B.n179 163.367
R1510 B.n180 B.n151 163.367
R1511 B.n184 B.n151 163.367
R1512 B.n185 B.n184 163.367
R1513 B.n186 B.n185 163.367
R1514 B.n186 B.n149 163.367
R1515 B.n190 B.n149 163.367
R1516 B.n191 B.n190 163.367
R1517 B.n192 B.n191 163.367
R1518 B.n192 B.n147 163.367
R1519 B.n263 B.n262 59.5399
R1520 B.n281 B.n119 59.5399
R1521 B.n46 B.n45 59.5399
R1522 B.n510 B.n39 59.5399
R1523 B.n262 B.n261 38.2066
R1524 B.n119 B.n118 38.2066
R1525 B.n45 B.n44 38.2066
R1526 B.n39 B.n38 38.2066
R1527 B.n577 B.n14 34.8103
R1528 B.n427 B.n426 34.8103
R1529 B.n349 B.n348 34.8103
R1530 B.n195 B.n194 34.8103
R1531 B B.n617 18.0485
R1532 B.n581 B.n14 10.6151
R1533 B.n582 B.n581 10.6151
R1534 B.n583 B.n582 10.6151
R1535 B.n583 B.n12 10.6151
R1536 B.n587 B.n12 10.6151
R1537 B.n588 B.n587 10.6151
R1538 B.n589 B.n588 10.6151
R1539 B.n589 B.n10 10.6151
R1540 B.n593 B.n10 10.6151
R1541 B.n594 B.n593 10.6151
R1542 B.n595 B.n594 10.6151
R1543 B.n595 B.n8 10.6151
R1544 B.n599 B.n8 10.6151
R1545 B.n600 B.n599 10.6151
R1546 B.n601 B.n600 10.6151
R1547 B.n601 B.n6 10.6151
R1548 B.n605 B.n6 10.6151
R1549 B.n606 B.n605 10.6151
R1550 B.n607 B.n606 10.6151
R1551 B.n607 B.n4 10.6151
R1552 B.n611 B.n4 10.6151
R1553 B.n612 B.n611 10.6151
R1554 B.n613 B.n612 10.6151
R1555 B.n613 B.n0 10.6151
R1556 B.n577 B.n576 10.6151
R1557 B.n576 B.n575 10.6151
R1558 B.n575 B.n16 10.6151
R1559 B.n571 B.n16 10.6151
R1560 B.n571 B.n570 10.6151
R1561 B.n570 B.n569 10.6151
R1562 B.n569 B.n18 10.6151
R1563 B.n565 B.n18 10.6151
R1564 B.n565 B.n564 10.6151
R1565 B.n564 B.n563 10.6151
R1566 B.n563 B.n20 10.6151
R1567 B.n559 B.n20 10.6151
R1568 B.n559 B.n558 10.6151
R1569 B.n558 B.n557 10.6151
R1570 B.n557 B.n22 10.6151
R1571 B.n553 B.n22 10.6151
R1572 B.n553 B.n552 10.6151
R1573 B.n552 B.n551 10.6151
R1574 B.n551 B.n24 10.6151
R1575 B.n547 B.n24 10.6151
R1576 B.n547 B.n546 10.6151
R1577 B.n546 B.n545 10.6151
R1578 B.n545 B.n26 10.6151
R1579 B.n541 B.n26 10.6151
R1580 B.n541 B.n540 10.6151
R1581 B.n540 B.n539 10.6151
R1582 B.n539 B.n28 10.6151
R1583 B.n535 B.n28 10.6151
R1584 B.n535 B.n534 10.6151
R1585 B.n534 B.n533 10.6151
R1586 B.n533 B.n30 10.6151
R1587 B.n529 B.n30 10.6151
R1588 B.n529 B.n528 10.6151
R1589 B.n528 B.n527 10.6151
R1590 B.n527 B.n32 10.6151
R1591 B.n523 B.n32 10.6151
R1592 B.n523 B.n522 10.6151
R1593 B.n522 B.n521 10.6151
R1594 B.n521 B.n34 10.6151
R1595 B.n517 B.n34 10.6151
R1596 B.n517 B.n516 10.6151
R1597 B.n516 B.n515 10.6151
R1598 B.n515 B.n36 10.6151
R1599 B.n511 B.n36 10.6151
R1600 B.n509 B.n508 10.6151
R1601 B.n508 B.n40 10.6151
R1602 B.n504 B.n40 10.6151
R1603 B.n504 B.n503 10.6151
R1604 B.n503 B.n502 10.6151
R1605 B.n502 B.n42 10.6151
R1606 B.n498 B.n42 10.6151
R1607 B.n498 B.n497 10.6151
R1608 B.n497 B.n496 10.6151
R1609 B.n493 B.n492 10.6151
R1610 B.n492 B.n491 10.6151
R1611 B.n491 B.n48 10.6151
R1612 B.n487 B.n48 10.6151
R1613 B.n487 B.n486 10.6151
R1614 B.n486 B.n485 10.6151
R1615 B.n485 B.n50 10.6151
R1616 B.n481 B.n50 10.6151
R1617 B.n481 B.n480 10.6151
R1618 B.n480 B.n479 10.6151
R1619 B.n479 B.n52 10.6151
R1620 B.n475 B.n52 10.6151
R1621 B.n475 B.n474 10.6151
R1622 B.n474 B.n473 10.6151
R1623 B.n473 B.n54 10.6151
R1624 B.n469 B.n54 10.6151
R1625 B.n469 B.n468 10.6151
R1626 B.n468 B.n467 10.6151
R1627 B.n467 B.n56 10.6151
R1628 B.n463 B.n56 10.6151
R1629 B.n463 B.n462 10.6151
R1630 B.n462 B.n461 10.6151
R1631 B.n461 B.n58 10.6151
R1632 B.n457 B.n58 10.6151
R1633 B.n457 B.n456 10.6151
R1634 B.n456 B.n455 10.6151
R1635 B.n455 B.n60 10.6151
R1636 B.n451 B.n60 10.6151
R1637 B.n451 B.n450 10.6151
R1638 B.n450 B.n449 10.6151
R1639 B.n449 B.n62 10.6151
R1640 B.n445 B.n62 10.6151
R1641 B.n445 B.n444 10.6151
R1642 B.n444 B.n443 10.6151
R1643 B.n443 B.n64 10.6151
R1644 B.n439 B.n64 10.6151
R1645 B.n439 B.n438 10.6151
R1646 B.n438 B.n437 10.6151
R1647 B.n437 B.n66 10.6151
R1648 B.n433 B.n66 10.6151
R1649 B.n433 B.n432 10.6151
R1650 B.n432 B.n431 10.6151
R1651 B.n431 B.n68 10.6151
R1652 B.n427 B.n68 10.6151
R1653 B.n426 B.n425 10.6151
R1654 B.n425 B.n70 10.6151
R1655 B.n421 B.n70 10.6151
R1656 B.n421 B.n420 10.6151
R1657 B.n420 B.n419 10.6151
R1658 B.n419 B.n72 10.6151
R1659 B.n415 B.n72 10.6151
R1660 B.n415 B.n414 10.6151
R1661 B.n414 B.n413 10.6151
R1662 B.n413 B.n74 10.6151
R1663 B.n409 B.n74 10.6151
R1664 B.n409 B.n408 10.6151
R1665 B.n408 B.n407 10.6151
R1666 B.n407 B.n76 10.6151
R1667 B.n403 B.n76 10.6151
R1668 B.n403 B.n402 10.6151
R1669 B.n402 B.n401 10.6151
R1670 B.n401 B.n78 10.6151
R1671 B.n397 B.n78 10.6151
R1672 B.n397 B.n396 10.6151
R1673 B.n396 B.n395 10.6151
R1674 B.n395 B.n80 10.6151
R1675 B.n391 B.n80 10.6151
R1676 B.n391 B.n390 10.6151
R1677 B.n390 B.n389 10.6151
R1678 B.n389 B.n82 10.6151
R1679 B.n385 B.n82 10.6151
R1680 B.n385 B.n384 10.6151
R1681 B.n384 B.n383 10.6151
R1682 B.n383 B.n84 10.6151
R1683 B.n379 B.n84 10.6151
R1684 B.n379 B.n378 10.6151
R1685 B.n378 B.n377 10.6151
R1686 B.n377 B.n86 10.6151
R1687 B.n373 B.n86 10.6151
R1688 B.n373 B.n372 10.6151
R1689 B.n372 B.n371 10.6151
R1690 B.n371 B.n88 10.6151
R1691 B.n367 B.n88 10.6151
R1692 B.n367 B.n366 10.6151
R1693 B.n366 B.n365 10.6151
R1694 B.n365 B.n90 10.6151
R1695 B.n361 B.n90 10.6151
R1696 B.n361 B.n360 10.6151
R1697 B.n360 B.n359 10.6151
R1698 B.n359 B.n92 10.6151
R1699 B.n355 B.n92 10.6151
R1700 B.n355 B.n354 10.6151
R1701 B.n354 B.n353 10.6151
R1702 B.n353 B.n94 10.6151
R1703 B.n349 B.n94 10.6151
R1704 B.n159 B.n1 10.6151
R1705 B.n159 B.n158 10.6151
R1706 B.n163 B.n158 10.6151
R1707 B.n164 B.n163 10.6151
R1708 B.n165 B.n164 10.6151
R1709 B.n165 B.n156 10.6151
R1710 B.n169 B.n156 10.6151
R1711 B.n170 B.n169 10.6151
R1712 B.n171 B.n170 10.6151
R1713 B.n171 B.n154 10.6151
R1714 B.n175 B.n154 10.6151
R1715 B.n176 B.n175 10.6151
R1716 B.n177 B.n176 10.6151
R1717 B.n177 B.n152 10.6151
R1718 B.n181 B.n152 10.6151
R1719 B.n182 B.n181 10.6151
R1720 B.n183 B.n182 10.6151
R1721 B.n183 B.n150 10.6151
R1722 B.n187 B.n150 10.6151
R1723 B.n188 B.n187 10.6151
R1724 B.n189 B.n188 10.6151
R1725 B.n189 B.n148 10.6151
R1726 B.n193 B.n148 10.6151
R1727 B.n194 B.n193 10.6151
R1728 B.n195 B.n146 10.6151
R1729 B.n199 B.n146 10.6151
R1730 B.n200 B.n199 10.6151
R1731 B.n201 B.n200 10.6151
R1732 B.n201 B.n144 10.6151
R1733 B.n205 B.n144 10.6151
R1734 B.n206 B.n205 10.6151
R1735 B.n207 B.n206 10.6151
R1736 B.n207 B.n142 10.6151
R1737 B.n211 B.n142 10.6151
R1738 B.n212 B.n211 10.6151
R1739 B.n213 B.n212 10.6151
R1740 B.n213 B.n140 10.6151
R1741 B.n217 B.n140 10.6151
R1742 B.n218 B.n217 10.6151
R1743 B.n219 B.n218 10.6151
R1744 B.n219 B.n138 10.6151
R1745 B.n223 B.n138 10.6151
R1746 B.n224 B.n223 10.6151
R1747 B.n225 B.n224 10.6151
R1748 B.n225 B.n136 10.6151
R1749 B.n229 B.n136 10.6151
R1750 B.n230 B.n229 10.6151
R1751 B.n231 B.n230 10.6151
R1752 B.n231 B.n134 10.6151
R1753 B.n235 B.n134 10.6151
R1754 B.n236 B.n235 10.6151
R1755 B.n237 B.n236 10.6151
R1756 B.n237 B.n132 10.6151
R1757 B.n241 B.n132 10.6151
R1758 B.n242 B.n241 10.6151
R1759 B.n243 B.n242 10.6151
R1760 B.n243 B.n130 10.6151
R1761 B.n247 B.n130 10.6151
R1762 B.n248 B.n247 10.6151
R1763 B.n249 B.n248 10.6151
R1764 B.n249 B.n128 10.6151
R1765 B.n253 B.n128 10.6151
R1766 B.n254 B.n253 10.6151
R1767 B.n255 B.n254 10.6151
R1768 B.n255 B.n126 10.6151
R1769 B.n259 B.n126 10.6151
R1770 B.n260 B.n259 10.6151
R1771 B.n264 B.n260 10.6151
R1772 B.n268 B.n124 10.6151
R1773 B.n269 B.n268 10.6151
R1774 B.n270 B.n269 10.6151
R1775 B.n270 B.n122 10.6151
R1776 B.n274 B.n122 10.6151
R1777 B.n275 B.n274 10.6151
R1778 B.n276 B.n275 10.6151
R1779 B.n276 B.n120 10.6151
R1780 B.n280 B.n120 10.6151
R1781 B.n283 B.n282 10.6151
R1782 B.n283 B.n116 10.6151
R1783 B.n287 B.n116 10.6151
R1784 B.n288 B.n287 10.6151
R1785 B.n289 B.n288 10.6151
R1786 B.n289 B.n114 10.6151
R1787 B.n293 B.n114 10.6151
R1788 B.n294 B.n293 10.6151
R1789 B.n295 B.n294 10.6151
R1790 B.n295 B.n112 10.6151
R1791 B.n299 B.n112 10.6151
R1792 B.n300 B.n299 10.6151
R1793 B.n301 B.n300 10.6151
R1794 B.n301 B.n110 10.6151
R1795 B.n305 B.n110 10.6151
R1796 B.n306 B.n305 10.6151
R1797 B.n307 B.n306 10.6151
R1798 B.n307 B.n108 10.6151
R1799 B.n311 B.n108 10.6151
R1800 B.n312 B.n311 10.6151
R1801 B.n313 B.n312 10.6151
R1802 B.n313 B.n106 10.6151
R1803 B.n317 B.n106 10.6151
R1804 B.n318 B.n317 10.6151
R1805 B.n319 B.n318 10.6151
R1806 B.n319 B.n104 10.6151
R1807 B.n323 B.n104 10.6151
R1808 B.n324 B.n323 10.6151
R1809 B.n325 B.n324 10.6151
R1810 B.n325 B.n102 10.6151
R1811 B.n329 B.n102 10.6151
R1812 B.n330 B.n329 10.6151
R1813 B.n331 B.n330 10.6151
R1814 B.n331 B.n100 10.6151
R1815 B.n335 B.n100 10.6151
R1816 B.n336 B.n335 10.6151
R1817 B.n337 B.n336 10.6151
R1818 B.n337 B.n98 10.6151
R1819 B.n341 B.n98 10.6151
R1820 B.n342 B.n341 10.6151
R1821 B.n343 B.n342 10.6151
R1822 B.n343 B.n96 10.6151
R1823 B.n347 B.n96 10.6151
R1824 B.n348 B.n347 10.6151
R1825 B.n511 B.n510 9.36635
R1826 B.n493 B.n46 9.36635
R1827 B.n264 B.n263 9.36635
R1828 B.n282 B.n281 9.36635
R1829 B.n617 B.n0 8.11757
R1830 B.n617 B.n1 8.11757
R1831 B.n510 B.n509 1.24928
R1832 B.n496 B.n46 1.24928
R1833 B.n263 B.n124 1.24928
R1834 B.n281 B.n280 1.24928
R1835 VN.n0 VN.t0 233.706
R1836 VN.n1 VN.t2 233.706
R1837 VN.n0 VN.t3 233.377
R1838 VN.n1 VN.t1 233.377
R1839 VN VN.n1 57.3123
R1840 VN VN.n0 12.5964
R1841 VDD2.n2 VDD2.n0 114.18
R1842 VDD2.n2 VDD2.n1 73.9058
R1843 VDD2.n1 VDD2.t2 2.44448
R1844 VDD2.n1 VDD2.t1 2.44448
R1845 VDD2.n0 VDD2.t3 2.44448
R1846 VDD2.n0 VDD2.t0 2.44448
R1847 VDD2 VDD2.n2 0.0586897
C0 VN B 0.938796f
C1 B w_n2152_n3628# 8.428901f
C2 B VDD2 1.16444f
C3 VN VDD1 0.147919f
C4 VDD1 w_n2152_n3628# 1.30128f
C5 VDD2 VDD1 0.794225f
C6 B VP 1.38938f
C7 VTAIL B 4.85412f
C8 VP VDD1 4.90343f
C9 VN w_n2152_n3628# 3.48461f
C10 VN VDD2 4.71884f
C11 VTAIL VDD1 5.84227f
C12 VDD2 w_n2152_n3628# 1.33592f
C13 VN VP 5.73954f
C14 VTAIL VN 4.44051f
C15 VP w_n2152_n3628# 3.75884f
C16 VP VDD2 0.333006f
C17 VTAIL w_n2152_n3628# 4.296f
C18 VTAIL VDD2 5.89004f
C19 B VDD1 1.12797f
C20 VTAIL VP 4.45462f
C21 VDD2 VSUBS 0.829914f
C22 VDD1 VSUBS 5.359685f
C23 VTAIL VSUBS 1.12936f
C24 VN VSUBS 5.23765f
C25 VP VSUBS 1.821087f
C26 B VSUBS 3.555265f
C27 w_n2152_n3628# VSUBS 95.9362f
C28 VDD2.t3 VSUBS 0.279884f
C29 VDD2.t0 VSUBS 0.279884f
C30 VDD2.n0 VSUBS 2.92884f
C31 VDD2.t2 VSUBS 0.279884f
C32 VDD2.t1 VSUBS 0.279884f
C33 VDD2.n1 VSUBS 2.23893f
C34 VDD2.n2 VSUBS 4.16123f
C35 VN.t0 VSUBS 2.60306f
C36 VN.t3 VSUBS 2.60158f
C37 VN.n0 VSUBS 1.82766f
C38 VN.t2 VSUBS 2.60306f
C39 VN.t1 VSUBS 2.60158f
C40 VN.n1 VSUBS 3.46718f
C41 B.n0 VSUBS 0.00634f
C42 B.n1 VSUBS 0.00634f
C43 B.n2 VSUBS 0.009377f
C44 B.n3 VSUBS 0.007186f
C45 B.n4 VSUBS 0.007186f
C46 B.n5 VSUBS 0.007186f
C47 B.n6 VSUBS 0.007186f
C48 B.n7 VSUBS 0.007186f
C49 B.n8 VSUBS 0.007186f
C50 B.n9 VSUBS 0.007186f
C51 B.n10 VSUBS 0.007186f
C52 B.n11 VSUBS 0.007186f
C53 B.n12 VSUBS 0.007186f
C54 B.n13 VSUBS 0.007186f
C55 B.n14 VSUBS 0.017318f
C56 B.n15 VSUBS 0.007186f
C57 B.n16 VSUBS 0.007186f
C58 B.n17 VSUBS 0.007186f
C59 B.n18 VSUBS 0.007186f
C60 B.n19 VSUBS 0.007186f
C61 B.n20 VSUBS 0.007186f
C62 B.n21 VSUBS 0.007186f
C63 B.n22 VSUBS 0.007186f
C64 B.n23 VSUBS 0.007186f
C65 B.n24 VSUBS 0.007186f
C66 B.n25 VSUBS 0.007186f
C67 B.n26 VSUBS 0.007186f
C68 B.n27 VSUBS 0.007186f
C69 B.n28 VSUBS 0.007186f
C70 B.n29 VSUBS 0.007186f
C71 B.n30 VSUBS 0.007186f
C72 B.n31 VSUBS 0.007186f
C73 B.n32 VSUBS 0.007186f
C74 B.n33 VSUBS 0.007186f
C75 B.n34 VSUBS 0.007186f
C76 B.n35 VSUBS 0.007186f
C77 B.n36 VSUBS 0.007186f
C78 B.n37 VSUBS 0.007186f
C79 B.t1 VSUBS 0.246489f
C80 B.t2 VSUBS 0.269441f
C81 B.t0 VSUBS 0.979132f
C82 B.n38 VSUBS 0.407198f
C83 B.n39 VSUBS 0.272813f
C84 B.n40 VSUBS 0.007186f
C85 B.n41 VSUBS 0.007186f
C86 B.n42 VSUBS 0.007186f
C87 B.n43 VSUBS 0.007186f
C88 B.t10 VSUBS 0.246493f
C89 B.t11 VSUBS 0.269444f
C90 B.t9 VSUBS 0.979132f
C91 B.n44 VSUBS 0.407195f
C92 B.n45 VSUBS 0.27281f
C93 B.n46 VSUBS 0.016649f
C94 B.n47 VSUBS 0.007186f
C95 B.n48 VSUBS 0.007186f
C96 B.n49 VSUBS 0.007186f
C97 B.n50 VSUBS 0.007186f
C98 B.n51 VSUBS 0.007186f
C99 B.n52 VSUBS 0.007186f
C100 B.n53 VSUBS 0.007186f
C101 B.n54 VSUBS 0.007186f
C102 B.n55 VSUBS 0.007186f
C103 B.n56 VSUBS 0.007186f
C104 B.n57 VSUBS 0.007186f
C105 B.n58 VSUBS 0.007186f
C106 B.n59 VSUBS 0.007186f
C107 B.n60 VSUBS 0.007186f
C108 B.n61 VSUBS 0.007186f
C109 B.n62 VSUBS 0.007186f
C110 B.n63 VSUBS 0.007186f
C111 B.n64 VSUBS 0.007186f
C112 B.n65 VSUBS 0.007186f
C113 B.n66 VSUBS 0.007186f
C114 B.n67 VSUBS 0.007186f
C115 B.n68 VSUBS 0.007186f
C116 B.n69 VSUBS 0.017318f
C117 B.n70 VSUBS 0.007186f
C118 B.n71 VSUBS 0.007186f
C119 B.n72 VSUBS 0.007186f
C120 B.n73 VSUBS 0.007186f
C121 B.n74 VSUBS 0.007186f
C122 B.n75 VSUBS 0.007186f
C123 B.n76 VSUBS 0.007186f
C124 B.n77 VSUBS 0.007186f
C125 B.n78 VSUBS 0.007186f
C126 B.n79 VSUBS 0.007186f
C127 B.n80 VSUBS 0.007186f
C128 B.n81 VSUBS 0.007186f
C129 B.n82 VSUBS 0.007186f
C130 B.n83 VSUBS 0.007186f
C131 B.n84 VSUBS 0.007186f
C132 B.n85 VSUBS 0.007186f
C133 B.n86 VSUBS 0.007186f
C134 B.n87 VSUBS 0.007186f
C135 B.n88 VSUBS 0.007186f
C136 B.n89 VSUBS 0.007186f
C137 B.n90 VSUBS 0.007186f
C138 B.n91 VSUBS 0.007186f
C139 B.n92 VSUBS 0.007186f
C140 B.n93 VSUBS 0.007186f
C141 B.n94 VSUBS 0.007186f
C142 B.n95 VSUBS 0.017765f
C143 B.n96 VSUBS 0.007186f
C144 B.n97 VSUBS 0.007186f
C145 B.n98 VSUBS 0.007186f
C146 B.n99 VSUBS 0.007186f
C147 B.n100 VSUBS 0.007186f
C148 B.n101 VSUBS 0.007186f
C149 B.n102 VSUBS 0.007186f
C150 B.n103 VSUBS 0.007186f
C151 B.n104 VSUBS 0.007186f
C152 B.n105 VSUBS 0.007186f
C153 B.n106 VSUBS 0.007186f
C154 B.n107 VSUBS 0.007186f
C155 B.n108 VSUBS 0.007186f
C156 B.n109 VSUBS 0.007186f
C157 B.n110 VSUBS 0.007186f
C158 B.n111 VSUBS 0.007186f
C159 B.n112 VSUBS 0.007186f
C160 B.n113 VSUBS 0.007186f
C161 B.n114 VSUBS 0.007186f
C162 B.n115 VSUBS 0.007186f
C163 B.n116 VSUBS 0.007186f
C164 B.n117 VSUBS 0.007186f
C165 B.t8 VSUBS 0.246493f
C166 B.t7 VSUBS 0.269444f
C167 B.t6 VSUBS 0.979132f
C168 B.n118 VSUBS 0.407195f
C169 B.n119 VSUBS 0.27281f
C170 B.n120 VSUBS 0.007186f
C171 B.n121 VSUBS 0.007186f
C172 B.n122 VSUBS 0.007186f
C173 B.n123 VSUBS 0.007186f
C174 B.n124 VSUBS 0.004016f
C175 B.n125 VSUBS 0.007186f
C176 B.n126 VSUBS 0.007186f
C177 B.n127 VSUBS 0.007186f
C178 B.n128 VSUBS 0.007186f
C179 B.n129 VSUBS 0.007186f
C180 B.n130 VSUBS 0.007186f
C181 B.n131 VSUBS 0.007186f
C182 B.n132 VSUBS 0.007186f
C183 B.n133 VSUBS 0.007186f
C184 B.n134 VSUBS 0.007186f
C185 B.n135 VSUBS 0.007186f
C186 B.n136 VSUBS 0.007186f
C187 B.n137 VSUBS 0.007186f
C188 B.n138 VSUBS 0.007186f
C189 B.n139 VSUBS 0.007186f
C190 B.n140 VSUBS 0.007186f
C191 B.n141 VSUBS 0.007186f
C192 B.n142 VSUBS 0.007186f
C193 B.n143 VSUBS 0.007186f
C194 B.n144 VSUBS 0.007186f
C195 B.n145 VSUBS 0.007186f
C196 B.n146 VSUBS 0.007186f
C197 B.n147 VSUBS 0.017318f
C198 B.n148 VSUBS 0.007186f
C199 B.n149 VSUBS 0.007186f
C200 B.n150 VSUBS 0.007186f
C201 B.n151 VSUBS 0.007186f
C202 B.n152 VSUBS 0.007186f
C203 B.n153 VSUBS 0.007186f
C204 B.n154 VSUBS 0.007186f
C205 B.n155 VSUBS 0.007186f
C206 B.n156 VSUBS 0.007186f
C207 B.n157 VSUBS 0.007186f
C208 B.n158 VSUBS 0.007186f
C209 B.n159 VSUBS 0.007186f
C210 B.n160 VSUBS 0.007186f
C211 B.n161 VSUBS 0.007186f
C212 B.n162 VSUBS 0.007186f
C213 B.n163 VSUBS 0.007186f
C214 B.n164 VSUBS 0.007186f
C215 B.n165 VSUBS 0.007186f
C216 B.n166 VSUBS 0.007186f
C217 B.n167 VSUBS 0.007186f
C218 B.n168 VSUBS 0.007186f
C219 B.n169 VSUBS 0.007186f
C220 B.n170 VSUBS 0.007186f
C221 B.n171 VSUBS 0.007186f
C222 B.n172 VSUBS 0.007186f
C223 B.n173 VSUBS 0.007186f
C224 B.n174 VSUBS 0.007186f
C225 B.n175 VSUBS 0.007186f
C226 B.n176 VSUBS 0.007186f
C227 B.n177 VSUBS 0.007186f
C228 B.n178 VSUBS 0.007186f
C229 B.n179 VSUBS 0.007186f
C230 B.n180 VSUBS 0.007186f
C231 B.n181 VSUBS 0.007186f
C232 B.n182 VSUBS 0.007186f
C233 B.n183 VSUBS 0.007186f
C234 B.n184 VSUBS 0.007186f
C235 B.n185 VSUBS 0.007186f
C236 B.n186 VSUBS 0.007186f
C237 B.n187 VSUBS 0.007186f
C238 B.n188 VSUBS 0.007186f
C239 B.n189 VSUBS 0.007186f
C240 B.n190 VSUBS 0.007186f
C241 B.n191 VSUBS 0.007186f
C242 B.n192 VSUBS 0.007186f
C243 B.n193 VSUBS 0.007186f
C244 B.n194 VSUBS 0.017318f
C245 B.n195 VSUBS 0.017765f
C246 B.n196 VSUBS 0.017765f
C247 B.n197 VSUBS 0.007186f
C248 B.n198 VSUBS 0.007186f
C249 B.n199 VSUBS 0.007186f
C250 B.n200 VSUBS 0.007186f
C251 B.n201 VSUBS 0.007186f
C252 B.n202 VSUBS 0.007186f
C253 B.n203 VSUBS 0.007186f
C254 B.n204 VSUBS 0.007186f
C255 B.n205 VSUBS 0.007186f
C256 B.n206 VSUBS 0.007186f
C257 B.n207 VSUBS 0.007186f
C258 B.n208 VSUBS 0.007186f
C259 B.n209 VSUBS 0.007186f
C260 B.n210 VSUBS 0.007186f
C261 B.n211 VSUBS 0.007186f
C262 B.n212 VSUBS 0.007186f
C263 B.n213 VSUBS 0.007186f
C264 B.n214 VSUBS 0.007186f
C265 B.n215 VSUBS 0.007186f
C266 B.n216 VSUBS 0.007186f
C267 B.n217 VSUBS 0.007186f
C268 B.n218 VSUBS 0.007186f
C269 B.n219 VSUBS 0.007186f
C270 B.n220 VSUBS 0.007186f
C271 B.n221 VSUBS 0.007186f
C272 B.n222 VSUBS 0.007186f
C273 B.n223 VSUBS 0.007186f
C274 B.n224 VSUBS 0.007186f
C275 B.n225 VSUBS 0.007186f
C276 B.n226 VSUBS 0.007186f
C277 B.n227 VSUBS 0.007186f
C278 B.n228 VSUBS 0.007186f
C279 B.n229 VSUBS 0.007186f
C280 B.n230 VSUBS 0.007186f
C281 B.n231 VSUBS 0.007186f
C282 B.n232 VSUBS 0.007186f
C283 B.n233 VSUBS 0.007186f
C284 B.n234 VSUBS 0.007186f
C285 B.n235 VSUBS 0.007186f
C286 B.n236 VSUBS 0.007186f
C287 B.n237 VSUBS 0.007186f
C288 B.n238 VSUBS 0.007186f
C289 B.n239 VSUBS 0.007186f
C290 B.n240 VSUBS 0.007186f
C291 B.n241 VSUBS 0.007186f
C292 B.n242 VSUBS 0.007186f
C293 B.n243 VSUBS 0.007186f
C294 B.n244 VSUBS 0.007186f
C295 B.n245 VSUBS 0.007186f
C296 B.n246 VSUBS 0.007186f
C297 B.n247 VSUBS 0.007186f
C298 B.n248 VSUBS 0.007186f
C299 B.n249 VSUBS 0.007186f
C300 B.n250 VSUBS 0.007186f
C301 B.n251 VSUBS 0.007186f
C302 B.n252 VSUBS 0.007186f
C303 B.n253 VSUBS 0.007186f
C304 B.n254 VSUBS 0.007186f
C305 B.n255 VSUBS 0.007186f
C306 B.n256 VSUBS 0.007186f
C307 B.n257 VSUBS 0.007186f
C308 B.n258 VSUBS 0.007186f
C309 B.n259 VSUBS 0.007186f
C310 B.n260 VSUBS 0.007186f
C311 B.t5 VSUBS 0.246489f
C312 B.t4 VSUBS 0.269441f
C313 B.t3 VSUBS 0.979132f
C314 B.n261 VSUBS 0.407198f
C315 B.n262 VSUBS 0.272813f
C316 B.n263 VSUBS 0.016649f
C317 B.n264 VSUBS 0.006763f
C318 B.n265 VSUBS 0.007186f
C319 B.n266 VSUBS 0.007186f
C320 B.n267 VSUBS 0.007186f
C321 B.n268 VSUBS 0.007186f
C322 B.n269 VSUBS 0.007186f
C323 B.n270 VSUBS 0.007186f
C324 B.n271 VSUBS 0.007186f
C325 B.n272 VSUBS 0.007186f
C326 B.n273 VSUBS 0.007186f
C327 B.n274 VSUBS 0.007186f
C328 B.n275 VSUBS 0.007186f
C329 B.n276 VSUBS 0.007186f
C330 B.n277 VSUBS 0.007186f
C331 B.n278 VSUBS 0.007186f
C332 B.n279 VSUBS 0.007186f
C333 B.n280 VSUBS 0.004016f
C334 B.n281 VSUBS 0.016649f
C335 B.n282 VSUBS 0.006763f
C336 B.n283 VSUBS 0.007186f
C337 B.n284 VSUBS 0.007186f
C338 B.n285 VSUBS 0.007186f
C339 B.n286 VSUBS 0.007186f
C340 B.n287 VSUBS 0.007186f
C341 B.n288 VSUBS 0.007186f
C342 B.n289 VSUBS 0.007186f
C343 B.n290 VSUBS 0.007186f
C344 B.n291 VSUBS 0.007186f
C345 B.n292 VSUBS 0.007186f
C346 B.n293 VSUBS 0.007186f
C347 B.n294 VSUBS 0.007186f
C348 B.n295 VSUBS 0.007186f
C349 B.n296 VSUBS 0.007186f
C350 B.n297 VSUBS 0.007186f
C351 B.n298 VSUBS 0.007186f
C352 B.n299 VSUBS 0.007186f
C353 B.n300 VSUBS 0.007186f
C354 B.n301 VSUBS 0.007186f
C355 B.n302 VSUBS 0.007186f
C356 B.n303 VSUBS 0.007186f
C357 B.n304 VSUBS 0.007186f
C358 B.n305 VSUBS 0.007186f
C359 B.n306 VSUBS 0.007186f
C360 B.n307 VSUBS 0.007186f
C361 B.n308 VSUBS 0.007186f
C362 B.n309 VSUBS 0.007186f
C363 B.n310 VSUBS 0.007186f
C364 B.n311 VSUBS 0.007186f
C365 B.n312 VSUBS 0.007186f
C366 B.n313 VSUBS 0.007186f
C367 B.n314 VSUBS 0.007186f
C368 B.n315 VSUBS 0.007186f
C369 B.n316 VSUBS 0.007186f
C370 B.n317 VSUBS 0.007186f
C371 B.n318 VSUBS 0.007186f
C372 B.n319 VSUBS 0.007186f
C373 B.n320 VSUBS 0.007186f
C374 B.n321 VSUBS 0.007186f
C375 B.n322 VSUBS 0.007186f
C376 B.n323 VSUBS 0.007186f
C377 B.n324 VSUBS 0.007186f
C378 B.n325 VSUBS 0.007186f
C379 B.n326 VSUBS 0.007186f
C380 B.n327 VSUBS 0.007186f
C381 B.n328 VSUBS 0.007186f
C382 B.n329 VSUBS 0.007186f
C383 B.n330 VSUBS 0.007186f
C384 B.n331 VSUBS 0.007186f
C385 B.n332 VSUBS 0.007186f
C386 B.n333 VSUBS 0.007186f
C387 B.n334 VSUBS 0.007186f
C388 B.n335 VSUBS 0.007186f
C389 B.n336 VSUBS 0.007186f
C390 B.n337 VSUBS 0.007186f
C391 B.n338 VSUBS 0.007186f
C392 B.n339 VSUBS 0.007186f
C393 B.n340 VSUBS 0.007186f
C394 B.n341 VSUBS 0.007186f
C395 B.n342 VSUBS 0.007186f
C396 B.n343 VSUBS 0.007186f
C397 B.n344 VSUBS 0.007186f
C398 B.n345 VSUBS 0.007186f
C399 B.n346 VSUBS 0.007186f
C400 B.n347 VSUBS 0.007186f
C401 B.n348 VSUBS 0.016968f
C402 B.n349 VSUBS 0.018115f
C403 B.n350 VSUBS 0.017318f
C404 B.n351 VSUBS 0.007186f
C405 B.n352 VSUBS 0.007186f
C406 B.n353 VSUBS 0.007186f
C407 B.n354 VSUBS 0.007186f
C408 B.n355 VSUBS 0.007186f
C409 B.n356 VSUBS 0.007186f
C410 B.n357 VSUBS 0.007186f
C411 B.n358 VSUBS 0.007186f
C412 B.n359 VSUBS 0.007186f
C413 B.n360 VSUBS 0.007186f
C414 B.n361 VSUBS 0.007186f
C415 B.n362 VSUBS 0.007186f
C416 B.n363 VSUBS 0.007186f
C417 B.n364 VSUBS 0.007186f
C418 B.n365 VSUBS 0.007186f
C419 B.n366 VSUBS 0.007186f
C420 B.n367 VSUBS 0.007186f
C421 B.n368 VSUBS 0.007186f
C422 B.n369 VSUBS 0.007186f
C423 B.n370 VSUBS 0.007186f
C424 B.n371 VSUBS 0.007186f
C425 B.n372 VSUBS 0.007186f
C426 B.n373 VSUBS 0.007186f
C427 B.n374 VSUBS 0.007186f
C428 B.n375 VSUBS 0.007186f
C429 B.n376 VSUBS 0.007186f
C430 B.n377 VSUBS 0.007186f
C431 B.n378 VSUBS 0.007186f
C432 B.n379 VSUBS 0.007186f
C433 B.n380 VSUBS 0.007186f
C434 B.n381 VSUBS 0.007186f
C435 B.n382 VSUBS 0.007186f
C436 B.n383 VSUBS 0.007186f
C437 B.n384 VSUBS 0.007186f
C438 B.n385 VSUBS 0.007186f
C439 B.n386 VSUBS 0.007186f
C440 B.n387 VSUBS 0.007186f
C441 B.n388 VSUBS 0.007186f
C442 B.n389 VSUBS 0.007186f
C443 B.n390 VSUBS 0.007186f
C444 B.n391 VSUBS 0.007186f
C445 B.n392 VSUBS 0.007186f
C446 B.n393 VSUBS 0.007186f
C447 B.n394 VSUBS 0.007186f
C448 B.n395 VSUBS 0.007186f
C449 B.n396 VSUBS 0.007186f
C450 B.n397 VSUBS 0.007186f
C451 B.n398 VSUBS 0.007186f
C452 B.n399 VSUBS 0.007186f
C453 B.n400 VSUBS 0.007186f
C454 B.n401 VSUBS 0.007186f
C455 B.n402 VSUBS 0.007186f
C456 B.n403 VSUBS 0.007186f
C457 B.n404 VSUBS 0.007186f
C458 B.n405 VSUBS 0.007186f
C459 B.n406 VSUBS 0.007186f
C460 B.n407 VSUBS 0.007186f
C461 B.n408 VSUBS 0.007186f
C462 B.n409 VSUBS 0.007186f
C463 B.n410 VSUBS 0.007186f
C464 B.n411 VSUBS 0.007186f
C465 B.n412 VSUBS 0.007186f
C466 B.n413 VSUBS 0.007186f
C467 B.n414 VSUBS 0.007186f
C468 B.n415 VSUBS 0.007186f
C469 B.n416 VSUBS 0.007186f
C470 B.n417 VSUBS 0.007186f
C471 B.n418 VSUBS 0.007186f
C472 B.n419 VSUBS 0.007186f
C473 B.n420 VSUBS 0.007186f
C474 B.n421 VSUBS 0.007186f
C475 B.n422 VSUBS 0.007186f
C476 B.n423 VSUBS 0.007186f
C477 B.n424 VSUBS 0.007186f
C478 B.n425 VSUBS 0.007186f
C479 B.n426 VSUBS 0.017318f
C480 B.n427 VSUBS 0.017765f
C481 B.n428 VSUBS 0.017765f
C482 B.n429 VSUBS 0.007186f
C483 B.n430 VSUBS 0.007186f
C484 B.n431 VSUBS 0.007186f
C485 B.n432 VSUBS 0.007186f
C486 B.n433 VSUBS 0.007186f
C487 B.n434 VSUBS 0.007186f
C488 B.n435 VSUBS 0.007186f
C489 B.n436 VSUBS 0.007186f
C490 B.n437 VSUBS 0.007186f
C491 B.n438 VSUBS 0.007186f
C492 B.n439 VSUBS 0.007186f
C493 B.n440 VSUBS 0.007186f
C494 B.n441 VSUBS 0.007186f
C495 B.n442 VSUBS 0.007186f
C496 B.n443 VSUBS 0.007186f
C497 B.n444 VSUBS 0.007186f
C498 B.n445 VSUBS 0.007186f
C499 B.n446 VSUBS 0.007186f
C500 B.n447 VSUBS 0.007186f
C501 B.n448 VSUBS 0.007186f
C502 B.n449 VSUBS 0.007186f
C503 B.n450 VSUBS 0.007186f
C504 B.n451 VSUBS 0.007186f
C505 B.n452 VSUBS 0.007186f
C506 B.n453 VSUBS 0.007186f
C507 B.n454 VSUBS 0.007186f
C508 B.n455 VSUBS 0.007186f
C509 B.n456 VSUBS 0.007186f
C510 B.n457 VSUBS 0.007186f
C511 B.n458 VSUBS 0.007186f
C512 B.n459 VSUBS 0.007186f
C513 B.n460 VSUBS 0.007186f
C514 B.n461 VSUBS 0.007186f
C515 B.n462 VSUBS 0.007186f
C516 B.n463 VSUBS 0.007186f
C517 B.n464 VSUBS 0.007186f
C518 B.n465 VSUBS 0.007186f
C519 B.n466 VSUBS 0.007186f
C520 B.n467 VSUBS 0.007186f
C521 B.n468 VSUBS 0.007186f
C522 B.n469 VSUBS 0.007186f
C523 B.n470 VSUBS 0.007186f
C524 B.n471 VSUBS 0.007186f
C525 B.n472 VSUBS 0.007186f
C526 B.n473 VSUBS 0.007186f
C527 B.n474 VSUBS 0.007186f
C528 B.n475 VSUBS 0.007186f
C529 B.n476 VSUBS 0.007186f
C530 B.n477 VSUBS 0.007186f
C531 B.n478 VSUBS 0.007186f
C532 B.n479 VSUBS 0.007186f
C533 B.n480 VSUBS 0.007186f
C534 B.n481 VSUBS 0.007186f
C535 B.n482 VSUBS 0.007186f
C536 B.n483 VSUBS 0.007186f
C537 B.n484 VSUBS 0.007186f
C538 B.n485 VSUBS 0.007186f
C539 B.n486 VSUBS 0.007186f
C540 B.n487 VSUBS 0.007186f
C541 B.n488 VSUBS 0.007186f
C542 B.n489 VSUBS 0.007186f
C543 B.n490 VSUBS 0.007186f
C544 B.n491 VSUBS 0.007186f
C545 B.n492 VSUBS 0.007186f
C546 B.n493 VSUBS 0.006763f
C547 B.n494 VSUBS 0.007186f
C548 B.n495 VSUBS 0.007186f
C549 B.n496 VSUBS 0.004016f
C550 B.n497 VSUBS 0.007186f
C551 B.n498 VSUBS 0.007186f
C552 B.n499 VSUBS 0.007186f
C553 B.n500 VSUBS 0.007186f
C554 B.n501 VSUBS 0.007186f
C555 B.n502 VSUBS 0.007186f
C556 B.n503 VSUBS 0.007186f
C557 B.n504 VSUBS 0.007186f
C558 B.n505 VSUBS 0.007186f
C559 B.n506 VSUBS 0.007186f
C560 B.n507 VSUBS 0.007186f
C561 B.n508 VSUBS 0.007186f
C562 B.n509 VSUBS 0.004016f
C563 B.n510 VSUBS 0.016649f
C564 B.n511 VSUBS 0.006763f
C565 B.n512 VSUBS 0.007186f
C566 B.n513 VSUBS 0.007186f
C567 B.n514 VSUBS 0.007186f
C568 B.n515 VSUBS 0.007186f
C569 B.n516 VSUBS 0.007186f
C570 B.n517 VSUBS 0.007186f
C571 B.n518 VSUBS 0.007186f
C572 B.n519 VSUBS 0.007186f
C573 B.n520 VSUBS 0.007186f
C574 B.n521 VSUBS 0.007186f
C575 B.n522 VSUBS 0.007186f
C576 B.n523 VSUBS 0.007186f
C577 B.n524 VSUBS 0.007186f
C578 B.n525 VSUBS 0.007186f
C579 B.n526 VSUBS 0.007186f
C580 B.n527 VSUBS 0.007186f
C581 B.n528 VSUBS 0.007186f
C582 B.n529 VSUBS 0.007186f
C583 B.n530 VSUBS 0.007186f
C584 B.n531 VSUBS 0.007186f
C585 B.n532 VSUBS 0.007186f
C586 B.n533 VSUBS 0.007186f
C587 B.n534 VSUBS 0.007186f
C588 B.n535 VSUBS 0.007186f
C589 B.n536 VSUBS 0.007186f
C590 B.n537 VSUBS 0.007186f
C591 B.n538 VSUBS 0.007186f
C592 B.n539 VSUBS 0.007186f
C593 B.n540 VSUBS 0.007186f
C594 B.n541 VSUBS 0.007186f
C595 B.n542 VSUBS 0.007186f
C596 B.n543 VSUBS 0.007186f
C597 B.n544 VSUBS 0.007186f
C598 B.n545 VSUBS 0.007186f
C599 B.n546 VSUBS 0.007186f
C600 B.n547 VSUBS 0.007186f
C601 B.n548 VSUBS 0.007186f
C602 B.n549 VSUBS 0.007186f
C603 B.n550 VSUBS 0.007186f
C604 B.n551 VSUBS 0.007186f
C605 B.n552 VSUBS 0.007186f
C606 B.n553 VSUBS 0.007186f
C607 B.n554 VSUBS 0.007186f
C608 B.n555 VSUBS 0.007186f
C609 B.n556 VSUBS 0.007186f
C610 B.n557 VSUBS 0.007186f
C611 B.n558 VSUBS 0.007186f
C612 B.n559 VSUBS 0.007186f
C613 B.n560 VSUBS 0.007186f
C614 B.n561 VSUBS 0.007186f
C615 B.n562 VSUBS 0.007186f
C616 B.n563 VSUBS 0.007186f
C617 B.n564 VSUBS 0.007186f
C618 B.n565 VSUBS 0.007186f
C619 B.n566 VSUBS 0.007186f
C620 B.n567 VSUBS 0.007186f
C621 B.n568 VSUBS 0.007186f
C622 B.n569 VSUBS 0.007186f
C623 B.n570 VSUBS 0.007186f
C624 B.n571 VSUBS 0.007186f
C625 B.n572 VSUBS 0.007186f
C626 B.n573 VSUBS 0.007186f
C627 B.n574 VSUBS 0.007186f
C628 B.n575 VSUBS 0.007186f
C629 B.n576 VSUBS 0.007186f
C630 B.n577 VSUBS 0.017765f
C631 B.n578 VSUBS 0.017765f
C632 B.n579 VSUBS 0.017318f
C633 B.n580 VSUBS 0.007186f
C634 B.n581 VSUBS 0.007186f
C635 B.n582 VSUBS 0.007186f
C636 B.n583 VSUBS 0.007186f
C637 B.n584 VSUBS 0.007186f
C638 B.n585 VSUBS 0.007186f
C639 B.n586 VSUBS 0.007186f
C640 B.n587 VSUBS 0.007186f
C641 B.n588 VSUBS 0.007186f
C642 B.n589 VSUBS 0.007186f
C643 B.n590 VSUBS 0.007186f
C644 B.n591 VSUBS 0.007186f
C645 B.n592 VSUBS 0.007186f
C646 B.n593 VSUBS 0.007186f
C647 B.n594 VSUBS 0.007186f
C648 B.n595 VSUBS 0.007186f
C649 B.n596 VSUBS 0.007186f
C650 B.n597 VSUBS 0.007186f
C651 B.n598 VSUBS 0.007186f
C652 B.n599 VSUBS 0.007186f
C653 B.n600 VSUBS 0.007186f
C654 B.n601 VSUBS 0.007186f
C655 B.n602 VSUBS 0.007186f
C656 B.n603 VSUBS 0.007186f
C657 B.n604 VSUBS 0.007186f
C658 B.n605 VSUBS 0.007186f
C659 B.n606 VSUBS 0.007186f
C660 B.n607 VSUBS 0.007186f
C661 B.n608 VSUBS 0.007186f
C662 B.n609 VSUBS 0.007186f
C663 B.n610 VSUBS 0.007186f
C664 B.n611 VSUBS 0.007186f
C665 B.n612 VSUBS 0.007186f
C666 B.n613 VSUBS 0.007186f
C667 B.n614 VSUBS 0.007186f
C668 B.n615 VSUBS 0.009377f
C669 B.n616 VSUBS 0.009989f
C670 B.n617 VSUBS 0.019864f
C671 VDD1.t1 VSUBS 0.279927f
C672 VDD1.t2 VSUBS 0.279927f
C673 VDD1.n0 VSUBS 2.23979f
C674 VDD1.t0 VSUBS 0.279927f
C675 VDD1.t3 VSUBS 0.279927f
C676 VDD1.n1 VSUBS 2.95406f
C677 VTAIL.n0 VSUBS 0.023845f
C678 VTAIL.n1 VSUBS 0.022702f
C679 VTAIL.n2 VSUBS 0.012199f
C680 VTAIL.n3 VSUBS 0.028834f
C681 VTAIL.n4 VSUBS 0.012917f
C682 VTAIL.n5 VSUBS 0.022702f
C683 VTAIL.n6 VSUBS 0.012199f
C684 VTAIL.n7 VSUBS 0.028834f
C685 VTAIL.n8 VSUBS 0.012917f
C686 VTAIL.n9 VSUBS 0.022702f
C687 VTAIL.n10 VSUBS 0.012199f
C688 VTAIL.n11 VSUBS 0.028834f
C689 VTAIL.n12 VSUBS 0.012917f
C690 VTAIL.n13 VSUBS 0.022702f
C691 VTAIL.n14 VSUBS 0.012199f
C692 VTAIL.n15 VSUBS 0.028834f
C693 VTAIL.n16 VSUBS 0.012917f
C694 VTAIL.n17 VSUBS 0.022702f
C695 VTAIL.n18 VSUBS 0.012199f
C696 VTAIL.n19 VSUBS 0.028834f
C697 VTAIL.n20 VSUBS 0.012917f
C698 VTAIL.n21 VSUBS 1.27436f
C699 VTAIL.n22 VSUBS 0.012199f
C700 VTAIL.t4 VSUBS 0.061633f
C701 VTAIL.n23 VSUBS 0.148646f
C702 VTAIL.n24 VSUBS 0.018343f
C703 VTAIL.n25 VSUBS 0.021625f
C704 VTAIL.n26 VSUBS 0.028834f
C705 VTAIL.n27 VSUBS 0.012917f
C706 VTAIL.n28 VSUBS 0.012199f
C707 VTAIL.n29 VSUBS 0.022702f
C708 VTAIL.n30 VSUBS 0.022702f
C709 VTAIL.n31 VSUBS 0.012199f
C710 VTAIL.n32 VSUBS 0.012917f
C711 VTAIL.n33 VSUBS 0.028834f
C712 VTAIL.n34 VSUBS 0.028834f
C713 VTAIL.n35 VSUBS 0.012917f
C714 VTAIL.n36 VSUBS 0.012199f
C715 VTAIL.n37 VSUBS 0.022702f
C716 VTAIL.n38 VSUBS 0.022702f
C717 VTAIL.n39 VSUBS 0.012199f
C718 VTAIL.n40 VSUBS 0.012917f
C719 VTAIL.n41 VSUBS 0.028834f
C720 VTAIL.n42 VSUBS 0.028834f
C721 VTAIL.n43 VSUBS 0.012917f
C722 VTAIL.n44 VSUBS 0.012199f
C723 VTAIL.n45 VSUBS 0.022702f
C724 VTAIL.n46 VSUBS 0.022702f
C725 VTAIL.n47 VSUBS 0.012199f
C726 VTAIL.n48 VSUBS 0.012917f
C727 VTAIL.n49 VSUBS 0.028834f
C728 VTAIL.n50 VSUBS 0.028834f
C729 VTAIL.n51 VSUBS 0.012917f
C730 VTAIL.n52 VSUBS 0.012199f
C731 VTAIL.n53 VSUBS 0.022702f
C732 VTAIL.n54 VSUBS 0.022702f
C733 VTAIL.n55 VSUBS 0.012199f
C734 VTAIL.n56 VSUBS 0.012917f
C735 VTAIL.n57 VSUBS 0.028834f
C736 VTAIL.n58 VSUBS 0.028834f
C737 VTAIL.n59 VSUBS 0.012917f
C738 VTAIL.n60 VSUBS 0.012199f
C739 VTAIL.n61 VSUBS 0.022702f
C740 VTAIL.n62 VSUBS 0.022702f
C741 VTAIL.n63 VSUBS 0.012199f
C742 VTAIL.n64 VSUBS 0.012917f
C743 VTAIL.n65 VSUBS 0.028834f
C744 VTAIL.n66 VSUBS 0.070508f
C745 VTAIL.n67 VSUBS 0.012917f
C746 VTAIL.n68 VSUBS 0.023956f
C747 VTAIL.n69 VSUBS 0.055576f
C748 VTAIL.n70 VSUBS 0.053411f
C749 VTAIL.n71 VSUBS 0.121881f
C750 VTAIL.n72 VSUBS 0.023845f
C751 VTAIL.n73 VSUBS 0.022702f
C752 VTAIL.n74 VSUBS 0.012199f
C753 VTAIL.n75 VSUBS 0.028834f
C754 VTAIL.n76 VSUBS 0.012917f
C755 VTAIL.n77 VSUBS 0.022702f
C756 VTAIL.n78 VSUBS 0.012199f
C757 VTAIL.n79 VSUBS 0.028834f
C758 VTAIL.n80 VSUBS 0.012917f
C759 VTAIL.n81 VSUBS 0.022702f
C760 VTAIL.n82 VSUBS 0.012199f
C761 VTAIL.n83 VSUBS 0.028834f
C762 VTAIL.n84 VSUBS 0.012917f
C763 VTAIL.n85 VSUBS 0.022702f
C764 VTAIL.n86 VSUBS 0.012199f
C765 VTAIL.n87 VSUBS 0.028834f
C766 VTAIL.n88 VSUBS 0.012917f
C767 VTAIL.n89 VSUBS 0.022702f
C768 VTAIL.n90 VSUBS 0.012199f
C769 VTAIL.n91 VSUBS 0.028834f
C770 VTAIL.n92 VSUBS 0.012917f
C771 VTAIL.n93 VSUBS 1.27436f
C772 VTAIL.n94 VSUBS 0.012199f
C773 VTAIL.t0 VSUBS 0.061633f
C774 VTAIL.n95 VSUBS 0.148646f
C775 VTAIL.n96 VSUBS 0.018343f
C776 VTAIL.n97 VSUBS 0.021625f
C777 VTAIL.n98 VSUBS 0.028834f
C778 VTAIL.n99 VSUBS 0.012917f
C779 VTAIL.n100 VSUBS 0.012199f
C780 VTAIL.n101 VSUBS 0.022702f
C781 VTAIL.n102 VSUBS 0.022702f
C782 VTAIL.n103 VSUBS 0.012199f
C783 VTAIL.n104 VSUBS 0.012917f
C784 VTAIL.n105 VSUBS 0.028834f
C785 VTAIL.n106 VSUBS 0.028834f
C786 VTAIL.n107 VSUBS 0.012917f
C787 VTAIL.n108 VSUBS 0.012199f
C788 VTAIL.n109 VSUBS 0.022702f
C789 VTAIL.n110 VSUBS 0.022702f
C790 VTAIL.n111 VSUBS 0.012199f
C791 VTAIL.n112 VSUBS 0.012917f
C792 VTAIL.n113 VSUBS 0.028834f
C793 VTAIL.n114 VSUBS 0.028834f
C794 VTAIL.n115 VSUBS 0.012917f
C795 VTAIL.n116 VSUBS 0.012199f
C796 VTAIL.n117 VSUBS 0.022702f
C797 VTAIL.n118 VSUBS 0.022702f
C798 VTAIL.n119 VSUBS 0.012199f
C799 VTAIL.n120 VSUBS 0.012917f
C800 VTAIL.n121 VSUBS 0.028834f
C801 VTAIL.n122 VSUBS 0.028834f
C802 VTAIL.n123 VSUBS 0.012917f
C803 VTAIL.n124 VSUBS 0.012199f
C804 VTAIL.n125 VSUBS 0.022702f
C805 VTAIL.n126 VSUBS 0.022702f
C806 VTAIL.n127 VSUBS 0.012199f
C807 VTAIL.n128 VSUBS 0.012917f
C808 VTAIL.n129 VSUBS 0.028834f
C809 VTAIL.n130 VSUBS 0.028834f
C810 VTAIL.n131 VSUBS 0.012917f
C811 VTAIL.n132 VSUBS 0.012199f
C812 VTAIL.n133 VSUBS 0.022702f
C813 VTAIL.n134 VSUBS 0.022702f
C814 VTAIL.n135 VSUBS 0.012199f
C815 VTAIL.n136 VSUBS 0.012917f
C816 VTAIL.n137 VSUBS 0.028834f
C817 VTAIL.n138 VSUBS 0.070508f
C818 VTAIL.n139 VSUBS 0.012917f
C819 VTAIL.n140 VSUBS 0.023956f
C820 VTAIL.n141 VSUBS 0.055576f
C821 VTAIL.n142 VSUBS 0.053411f
C822 VTAIL.n143 VSUBS 0.17974f
C823 VTAIL.n144 VSUBS 0.023845f
C824 VTAIL.n145 VSUBS 0.022702f
C825 VTAIL.n146 VSUBS 0.012199f
C826 VTAIL.n147 VSUBS 0.028834f
C827 VTAIL.n148 VSUBS 0.012917f
C828 VTAIL.n149 VSUBS 0.022702f
C829 VTAIL.n150 VSUBS 0.012199f
C830 VTAIL.n151 VSUBS 0.028834f
C831 VTAIL.n152 VSUBS 0.012917f
C832 VTAIL.n153 VSUBS 0.022702f
C833 VTAIL.n154 VSUBS 0.012199f
C834 VTAIL.n155 VSUBS 0.028834f
C835 VTAIL.n156 VSUBS 0.012917f
C836 VTAIL.n157 VSUBS 0.022702f
C837 VTAIL.n158 VSUBS 0.012199f
C838 VTAIL.n159 VSUBS 0.028834f
C839 VTAIL.n160 VSUBS 0.012917f
C840 VTAIL.n161 VSUBS 0.022702f
C841 VTAIL.n162 VSUBS 0.012199f
C842 VTAIL.n163 VSUBS 0.028834f
C843 VTAIL.n164 VSUBS 0.012917f
C844 VTAIL.n165 VSUBS 1.27436f
C845 VTAIL.n166 VSUBS 0.012199f
C846 VTAIL.t2 VSUBS 0.061633f
C847 VTAIL.n167 VSUBS 0.148646f
C848 VTAIL.n168 VSUBS 0.018343f
C849 VTAIL.n169 VSUBS 0.021625f
C850 VTAIL.n170 VSUBS 0.028834f
C851 VTAIL.n171 VSUBS 0.012917f
C852 VTAIL.n172 VSUBS 0.012199f
C853 VTAIL.n173 VSUBS 0.022702f
C854 VTAIL.n174 VSUBS 0.022702f
C855 VTAIL.n175 VSUBS 0.012199f
C856 VTAIL.n176 VSUBS 0.012917f
C857 VTAIL.n177 VSUBS 0.028834f
C858 VTAIL.n178 VSUBS 0.028834f
C859 VTAIL.n179 VSUBS 0.012917f
C860 VTAIL.n180 VSUBS 0.012199f
C861 VTAIL.n181 VSUBS 0.022702f
C862 VTAIL.n182 VSUBS 0.022702f
C863 VTAIL.n183 VSUBS 0.012199f
C864 VTAIL.n184 VSUBS 0.012917f
C865 VTAIL.n185 VSUBS 0.028834f
C866 VTAIL.n186 VSUBS 0.028834f
C867 VTAIL.n187 VSUBS 0.012917f
C868 VTAIL.n188 VSUBS 0.012199f
C869 VTAIL.n189 VSUBS 0.022702f
C870 VTAIL.n190 VSUBS 0.022702f
C871 VTAIL.n191 VSUBS 0.012199f
C872 VTAIL.n192 VSUBS 0.012917f
C873 VTAIL.n193 VSUBS 0.028834f
C874 VTAIL.n194 VSUBS 0.028834f
C875 VTAIL.n195 VSUBS 0.012917f
C876 VTAIL.n196 VSUBS 0.012199f
C877 VTAIL.n197 VSUBS 0.022702f
C878 VTAIL.n198 VSUBS 0.022702f
C879 VTAIL.n199 VSUBS 0.012199f
C880 VTAIL.n200 VSUBS 0.012917f
C881 VTAIL.n201 VSUBS 0.028834f
C882 VTAIL.n202 VSUBS 0.028834f
C883 VTAIL.n203 VSUBS 0.012917f
C884 VTAIL.n204 VSUBS 0.012199f
C885 VTAIL.n205 VSUBS 0.022702f
C886 VTAIL.n206 VSUBS 0.022702f
C887 VTAIL.n207 VSUBS 0.012199f
C888 VTAIL.n208 VSUBS 0.012917f
C889 VTAIL.n209 VSUBS 0.028834f
C890 VTAIL.n210 VSUBS 0.070508f
C891 VTAIL.n211 VSUBS 0.012917f
C892 VTAIL.n212 VSUBS 0.023956f
C893 VTAIL.n213 VSUBS 0.055576f
C894 VTAIL.n214 VSUBS 0.053411f
C895 VTAIL.n215 VSUBS 1.41669f
C896 VTAIL.n216 VSUBS 0.023845f
C897 VTAIL.n217 VSUBS 0.022702f
C898 VTAIL.n218 VSUBS 0.012199f
C899 VTAIL.n219 VSUBS 0.028834f
C900 VTAIL.n220 VSUBS 0.012917f
C901 VTAIL.n221 VSUBS 0.022702f
C902 VTAIL.n222 VSUBS 0.012199f
C903 VTAIL.n223 VSUBS 0.028834f
C904 VTAIL.n224 VSUBS 0.012917f
C905 VTAIL.n225 VSUBS 0.022702f
C906 VTAIL.n226 VSUBS 0.012199f
C907 VTAIL.n227 VSUBS 0.028834f
C908 VTAIL.n228 VSUBS 0.012917f
C909 VTAIL.n229 VSUBS 0.022702f
C910 VTAIL.n230 VSUBS 0.012199f
C911 VTAIL.n231 VSUBS 0.028834f
C912 VTAIL.n232 VSUBS 0.012917f
C913 VTAIL.n233 VSUBS 0.022702f
C914 VTAIL.n234 VSUBS 0.012199f
C915 VTAIL.n235 VSUBS 0.028834f
C916 VTAIL.n236 VSUBS 0.012917f
C917 VTAIL.n237 VSUBS 1.27436f
C918 VTAIL.n238 VSUBS 0.012199f
C919 VTAIL.t5 VSUBS 0.061633f
C920 VTAIL.n239 VSUBS 0.148646f
C921 VTAIL.n240 VSUBS 0.018343f
C922 VTAIL.n241 VSUBS 0.021625f
C923 VTAIL.n242 VSUBS 0.028834f
C924 VTAIL.n243 VSUBS 0.012917f
C925 VTAIL.n244 VSUBS 0.012199f
C926 VTAIL.n245 VSUBS 0.022702f
C927 VTAIL.n246 VSUBS 0.022702f
C928 VTAIL.n247 VSUBS 0.012199f
C929 VTAIL.n248 VSUBS 0.012917f
C930 VTAIL.n249 VSUBS 0.028834f
C931 VTAIL.n250 VSUBS 0.028834f
C932 VTAIL.n251 VSUBS 0.012917f
C933 VTAIL.n252 VSUBS 0.012199f
C934 VTAIL.n253 VSUBS 0.022702f
C935 VTAIL.n254 VSUBS 0.022702f
C936 VTAIL.n255 VSUBS 0.012199f
C937 VTAIL.n256 VSUBS 0.012917f
C938 VTAIL.n257 VSUBS 0.028834f
C939 VTAIL.n258 VSUBS 0.028834f
C940 VTAIL.n259 VSUBS 0.012917f
C941 VTAIL.n260 VSUBS 0.012199f
C942 VTAIL.n261 VSUBS 0.022702f
C943 VTAIL.n262 VSUBS 0.022702f
C944 VTAIL.n263 VSUBS 0.012199f
C945 VTAIL.n264 VSUBS 0.012917f
C946 VTAIL.n265 VSUBS 0.028834f
C947 VTAIL.n266 VSUBS 0.028834f
C948 VTAIL.n267 VSUBS 0.012917f
C949 VTAIL.n268 VSUBS 0.012199f
C950 VTAIL.n269 VSUBS 0.022702f
C951 VTAIL.n270 VSUBS 0.022702f
C952 VTAIL.n271 VSUBS 0.012199f
C953 VTAIL.n272 VSUBS 0.012917f
C954 VTAIL.n273 VSUBS 0.028834f
C955 VTAIL.n274 VSUBS 0.028834f
C956 VTAIL.n275 VSUBS 0.012917f
C957 VTAIL.n276 VSUBS 0.012199f
C958 VTAIL.n277 VSUBS 0.022702f
C959 VTAIL.n278 VSUBS 0.022702f
C960 VTAIL.n279 VSUBS 0.012199f
C961 VTAIL.n280 VSUBS 0.012917f
C962 VTAIL.n281 VSUBS 0.028834f
C963 VTAIL.n282 VSUBS 0.070508f
C964 VTAIL.n283 VSUBS 0.012917f
C965 VTAIL.n284 VSUBS 0.023956f
C966 VTAIL.n285 VSUBS 0.055576f
C967 VTAIL.n286 VSUBS 0.053411f
C968 VTAIL.n287 VSUBS 1.41669f
C969 VTAIL.n288 VSUBS 0.023845f
C970 VTAIL.n289 VSUBS 0.022702f
C971 VTAIL.n290 VSUBS 0.012199f
C972 VTAIL.n291 VSUBS 0.028834f
C973 VTAIL.n292 VSUBS 0.012917f
C974 VTAIL.n293 VSUBS 0.022702f
C975 VTAIL.n294 VSUBS 0.012199f
C976 VTAIL.n295 VSUBS 0.028834f
C977 VTAIL.n296 VSUBS 0.012917f
C978 VTAIL.n297 VSUBS 0.022702f
C979 VTAIL.n298 VSUBS 0.012199f
C980 VTAIL.n299 VSUBS 0.028834f
C981 VTAIL.n300 VSUBS 0.012917f
C982 VTAIL.n301 VSUBS 0.022702f
C983 VTAIL.n302 VSUBS 0.012199f
C984 VTAIL.n303 VSUBS 0.028834f
C985 VTAIL.n304 VSUBS 0.012917f
C986 VTAIL.n305 VSUBS 0.022702f
C987 VTAIL.n306 VSUBS 0.012199f
C988 VTAIL.n307 VSUBS 0.028834f
C989 VTAIL.n308 VSUBS 0.012917f
C990 VTAIL.n309 VSUBS 1.27436f
C991 VTAIL.n310 VSUBS 0.012199f
C992 VTAIL.t7 VSUBS 0.061633f
C993 VTAIL.n311 VSUBS 0.148646f
C994 VTAIL.n312 VSUBS 0.018343f
C995 VTAIL.n313 VSUBS 0.021625f
C996 VTAIL.n314 VSUBS 0.028834f
C997 VTAIL.n315 VSUBS 0.012917f
C998 VTAIL.n316 VSUBS 0.012199f
C999 VTAIL.n317 VSUBS 0.022702f
C1000 VTAIL.n318 VSUBS 0.022702f
C1001 VTAIL.n319 VSUBS 0.012199f
C1002 VTAIL.n320 VSUBS 0.012917f
C1003 VTAIL.n321 VSUBS 0.028834f
C1004 VTAIL.n322 VSUBS 0.028834f
C1005 VTAIL.n323 VSUBS 0.012917f
C1006 VTAIL.n324 VSUBS 0.012199f
C1007 VTAIL.n325 VSUBS 0.022702f
C1008 VTAIL.n326 VSUBS 0.022702f
C1009 VTAIL.n327 VSUBS 0.012199f
C1010 VTAIL.n328 VSUBS 0.012917f
C1011 VTAIL.n329 VSUBS 0.028834f
C1012 VTAIL.n330 VSUBS 0.028834f
C1013 VTAIL.n331 VSUBS 0.012917f
C1014 VTAIL.n332 VSUBS 0.012199f
C1015 VTAIL.n333 VSUBS 0.022702f
C1016 VTAIL.n334 VSUBS 0.022702f
C1017 VTAIL.n335 VSUBS 0.012199f
C1018 VTAIL.n336 VSUBS 0.012917f
C1019 VTAIL.n337 VSUBS 0.028834f
C1020 VTAIL.n338 VSUBS 0.028834f
C1021 VTAIL.n339 VSUBS 0.012917f
C1022 VTAIL.n340 VSUBS 0.012199f
C1023 VTAIL.n341 VSUBS 0.022702f
C1024 VTAIL.n342 VSUBS 0.022702f
C1025 VTAIL.n343 VSUBS 0.012199f
C1026 VTAIL.n344 VSUBS 0.012917f
C1027 VTAIL.n345 VSUBS 0.028834f
C1028 VTAIL.n346 VSUBS 0.028834f
C1029 VTAIL.n347 VSUBS 0.012917f
C1030 VTAIL.n348 VSUBS 0.012199f
C1031 VTAIL.n349 VSUBS 0.022702f
C1032 VTAIL.n350 VSUBS 0.022702f
C1033 VTAIL.n351 VSUBS 0.012199f
C1034 VTAIL.n352 VSUBS 0.012917f
C1035 VTAIL.n353 VSUBS 0.028834f
C1036 VTAIL.n354 VSUBS 0.070508f
C1037 VTAIL.n355 VSUBS 0.012917f
C1038 VTAIL.n356 VSUBS 0.023956f
C1039 VTAIL.n357 VSUBS 0.055576f
C1040 VTAIL.n358 VSUBS 0.053411f
C1041 VTAIL.n359 VSUBS 0.17974f
C1042 VTAIL.n360 VSUBS 0.023845f
C1043 VTAIL.n361 VSUBS 0.022702f
C1044 VTAIL.n362 VSUBS 0.012199f
C1045 VTAIL.n363 VSUBS 0.028834f
C1046 VTAIL.n364 VSUBS 0.012917f
C1047 VTAIL.n365 VSUBS 0.022702f
C1048 VTAIL.n366 VSUBS 0.012199f
C1049 VTAIL.n367 VSUBS 0.028834f
C1050 VTAIL.n368 VSUBS 0.012917f
C1051 VTAIL.n369 VSUBS 0.022702f
C1052 VTAIL.n370 VSUBS 0.012199f
C1053 VTAIL.n371 VSUBS 0.028834f
C1054 VTAIL.n372 VSUBS 0.012917f
C1055 VTAIL.n373 VSUBS 0.022702f
C1056 VTAIL.n374 VSUBS 0.012199f
C1057 VTAIL.n375 VSUBS 0.028834f
C1058 VTAIL.n376 VSUBS 0.012917f
C1059 VTAIL.n377 VSUBS 0.022702f
C1060 VTAIL.n378 VSUBS 0.012199f
C1061 VTAIL.n379 VSUBS 0.028834f
C1062 VTAIL.n380 VSUBS 0.012917f
C1063 VTAIL.n381 VSUBS 1.27436f
C1064 VTAIL.n382 VSUBS 0.012199f
C1065 VTAIL.t3 VSUBS 0.061633f
C1066 VTAIL.n383 VSUBS 0.148646f
C1067 VTAIL.n384 VSUBS 0.018343f
C1068 VTAIL.n385 VSUBS 0.021625f
C1069 VTAIL.n386 VSUBS 0.028834f
C1070 VTAIL.n387 VSUBS 0.012917f
C1071 VTAIL.n388 VSUBS 0.012199f
C1072 VTAIL.n389 VSUBS 0.022702f
C1073 VTAIL.n390 VSUBS 0.022702f
C1074 VTAIL.n391 VSUBS 0.012199f
C1075 VTAIL.n392 VSUBS 0.012917f
C1076 VTAIL.n393 VSUBS 0.028834f
C1077 VTAIL.n394 VSUBS 0.028834f
C1078 VTAIL.n395 VSUBS 0.012917f
C1079 VTAIL.n396 VSUBS 0.012199f
C1080 VTAIL.n397 VSUBS 0.022702f
C1081 VTAIL.n398 VSUBS 0.022702f
C1082 VTAIL.n399 VSUBS 0.012199f
C1083 VTAIL.n400 VSUBS 0.012917f
C1084 VTAIL.n401 VSUBS 0.028834f
C1085 VTAIL.n402 VSUBS 0.028834f
C1086 VTAIL.n403 VSUBS 0.012917f
C1087 VTAIL.n404 VSUBS 0.012199f
C1088 VTAIL.n405 VSUBS 0.022702f
C1089 VTAIL.n406 VSUBS 0.022702f
C1090 VTAIL.n407 VSUBS 0.012199f
C1091 VTAIL.n408 VSUBS 0.012917f
C1092 VTAIL.n409 VSUBS 0.028834f
C1093 VTAIL.n410 VSUBS 0.028834f
C1094 VTAIL.n411 VSUBS 0.012917f
C1095 VTAIL.n412 VSUBS 0.012199f
C1096 VTAIL.n413 VSUBS 0.022702f
C1097 VTAIL.n414 VSUBS 0.022702f
C1098 VTAIL.n415 VSUBS 0.012199f
C1099 VTAIL.n416 VSUBS 0.012917f
C1100 VTAIL.n417 VSUBS 0.028834f
C1101 VTAIL.n418 VSUBS 0.028834f
C1102 VTAIL.n419 VSUBS 0.012917f
C1103 VTAIL.n420 VSUBS 0.012199f
C1104 VTAIL.n421 VSUBS 0.022702f
C1105 VTAIL.n422 VSUBS 0.022702f
C1106 VTAIL.n423 VSUBS 0.012199f
C1107 VTAIL.n424 VSUBS 0.012917f
C1108 VTAIL.n425 VSUBS 0.028834f
C1109 VTAIL.n426 VSUBS 0.070508f
C1110 VTAIL.n427 VSUBS 0.012917f
C1111 VTAIL.n428 VSUBS 0.023956f
C1112 VTAIL.n429 VSUBS 0.055576f
C1113 VTAIL.n430 VSUBS 0.053411f
C1114 VTAIL.n431 VSUBS 0.17974f
C1115 VTAIL.n432 VSUBS 0.023845f
C1116 VTAIL.n433 VSUBS 0.022702f
C1117 VTAIL.n434 VSUBS 0.012199f
C1118 VTAIL.n435 VSUBS 0.028834f
C1119 VTAIL.n436 VSUBS 0.012917f
C1120 VTAIL.n437 VSUBS 0.022702f
C1121 VTAIL.n438 VSUBS 0.012199f
C1122 VTAIL.n439 VSUBS 0.028834f
C1123 VTAIL.n440 VSUBS 0.012917f
C1124 VTAIL.n441 VSUBS 0.022702f
C1125 VTAIL.n442 VSUBS 0.012199f
C1126 VTAIL.n443 VSUBS 0.028834f
C1127 VTAIL.n444 VSUBS 0.012917f
C1128 VTAIL.n445 VSUBS 0.022702f
C1129 VTAIL.n446 VSUBS 0.012199f
C1130 VTAIL.n447 VSUBS 0.028834f
C1131 VTAIL.n448 VSUBS 0.012917f
C1132 VTAIL.n449 VSUBS 0.022702f
C1133 VTAIL.n450 VSUBS 0.012199f
C1134 VTAIL.n451 VSUBS 0.028834f
C1135 VTAIL.n452 VSUBS 0.012917f
C1136 VTAIL.n453 VSUBS 1.27436f
C1137 VTAIL.n454 VSUBS 0.012199f
C1138 VTAIL.t1 VSUBS 0.061633f
C1139 VTAIL.n455 VSUBS 0.148646f
C1140 VTAIL.n456 VSUBS 0.018343f
C1141 VTAIL.n457 VSUBS 0.021625f
C1142 VTAIL.n458 VSUBS 0.028834f
C1143 VTAIL.n459 VSUBS 0.012917f
C1144 VTAIL.n460 VSUBS 0.012199f
C1145 VTAIL.n461 VSUBS 0.022702f
C1146 VTAIL.n462 VSUBS 0.022702f
C1147 VTAIL.n463 VSUBS 0.012199f
C1148 VTAIL.n464 VSUBS 0.012917f
C1149 VTAIL.n465 VSUBS 0.028834f
C1150 VTAIL.n466 VSUBS 0.028834f
C1151 VTAIL.n467 VSUBS 0.012917f
C1152 VTAIL.n468 VSUBS 0.012199f
C1153 VTAIL.n469 VSUBS 0.022702f
C1154 VTAIL.n470 VSUBS 0.022702f
C1155 VTAIL.n471 VSUBS 0.012199f
C1156 VTAIL.n472 VSUBS 0.012917f
C1157 VTAIL.n473 VSUBS 0.028834f
C1158 VTAIL.n474 VSUBS 0.028834f
C1159 VTAIL.n475 VSUBS 0.012917f
C1160 VTAIL.n476 VSUBS 0.012199f
C1161 VTAIL.n477 VSUBS 0.022702f
C1162 VTAIL.n478 VSUBS 0.022702f
C1163 VTAIL.n479 VSUBS 0.012199f
C1164 VTAIL.n480 VSUBS 0.012917f
C1165 VTAIL.n481 VSUBS 0.028834f
C1166 VTAIL.n482 VSUBS 0.028834f
C1167 VTAIL.n483 VSUBS 0.012917f
C1168 VTAIL.n484 VSUBS 0.012199f
C1169 VTAIL.n485 VSUBS 0.022702f
C1170 VTAIL.n486 VSUBS 0.022702f
C1171 VTAIL.n487 VSUBS 0.012199f
C1172 VTAIL.n488 VSUBS 0.012917f
C1173 VTAIL.n489 VSUBS 0.028834f
C1174 VTAIL.n490 VSUBS 0.028834f
C1175 VTAIL.n491 VSUBS 0.012917f
C1176 VTAIL.n492 VSUBS 0.012199f
C1177 VTAIL.n493 VSUBS 0.022702f
C1178 VTAIL.n494 VSUBS 0.022702f
C1179 VTAIL.n495 VSUBS 0.012199f
C1180 VTAIL.n496 VSUBS 0.012917f
C1181 VTAIL.n497 VSUBS 0.028834f
C1182 VTAIL.n498 VSUBS 0.070508f
C1183 VTAIL.n499 VSUBS 0.012917f
C1184 VTAIL.n500 VSUBS 0.023956f
C1185 VTAIL.n501 VSUBS 0.055576f
C1186 VTAIL.n502 VSUBS 0.053411f
C1187 VTAIL.n503 VSUBS 1.41669f
C1188 VTAIL.n504 VSUBS 0.023845f
C1189 VTAIL.n505 VSUBS 0.022702f
C1190 VTAIL.n506 VSUBS 0.012199f
C1191 VTAIL.n507 VSUBS 0.028834f
C1192 VTAIL.n508 VSUBS 0.012917f
C1193 VTAIL.n509 VSUBS 0.022702f
C1194 VTAIL.n510 VSUBS 0.012199f
C1195 VTAIL.n511 VSUBS 0.028834f
C1196 VTAIL.n512 VSUBS 0.012917f
C1197 VTAIL.n513 VSUBS 0.022702f
C1198 VTAIL.n514 VSUBS 0.012199f
C1199 VTAIL.n515 VSUBS 0.028834f
C1200 VTAIL.n516 VSUBS 0.012917f
C1201 VTAIL.n517 VSUBS 0.022702f
C1202 VTAIL.n518 VSUBS 0.012199f
C1203 VTAIL.n519 VSUBS 0.028834f
C1204 VTAIL.n520 VSUBS 0.012917f
C1205 VTAIL.n521 VSUBS 0.022702f
C1206 VTAIL.n522 VSUBS 0.012199f
C1207 VTAIL.n523 VSUBS 0.028834f
C1208 VTAIL.n524 VSUBS 0.012917f
C1209 VTAIL.n525 VSUBS 1.27436f
C1210 VTAIL.n526 VSUBS 0.012199f
C1211 VTAIL.t6 VSUBS 0.061633f
C1212 VTAIL.n527 VSUBS 0.148646f
C1213 VTAIL.n528 VSUBS 0.018343f
C1214 VTAIL.n529 VSUBS 0.021625f
C1215 VTAIL.n530 VSUBS 0.028834f
C1216 VTAIL.n531 VSUBS 0.012917f
C1217 VTAIL.n532 VSUBS 0.012199f
C1218 VTAIL.n533 VSUBS 0.022702f
C1219 VTAIL.n534 VSUBS 0.022702f
C1220 VTAIL.n535 VSUBS 0.012199f
C1221 VTAIL.n536 VSUBS 0.012917f
C1222 VTAIL.n537 VSUBS 0.028834f
C1223 VTAIL.n538 VSUBS 0.028834f
C1224 VTAIL.n539 VSUBS 0.012917f
C1225 VTAIL.n540 VSUBS 0.012199f
C1226 VTAIL.n541 VSUBS 0.022702f
C1227 VTAIL.n542 VSUBS 0.022702f
C1228 VTAIL.n543 VSUBS 0.012199f
C1229 VTAIL.n544 VSUBS 0.012917f
C1230 VTAIL.n545 VSUBS 0.028834f
C1231 VTAIL.n546 VSUBS 0.028834f
C1232 VTAIL.n547 VSUBS 0.012917f
C1233 VTAIL.n548 VSUBS 0.012199f
C1234 VTAIL.n549 VSUBS 0.022702f
C1235 VTAIL.n550 VSUBS 0.022702f
C1236 VTAIL.n551 VSUBS 0.012199f
C1237 VTAIL.n552 VSUBS 0.012917f
C1238 VTAIL.n553 VSUBS 0.028834f
C1239 VTAIL.n554 VSUBS 0.028834f
C1240 VTAIL.n555 VSUBS 0.012917f
C1241 VTAIL.n556 VSUBS 0.012199f
C1242 VTAIL.n557 VSUBS 0.022702f
C1243 VTAIL.n558 VSUBS 0.022702f
C1244 VTAIL.n559 VSUBS 0.012199f
C1245 VTAIL.n560 VSUBS 0.012917f
C1246 VTAIL.n561 VSUBS 0.028834f
C1247 VTAIL.n562 VSUBS 0.028834f
C1248 VTAIL.n563 VSUBS 0.012917f
C1249 VTAIL.n564 VSUBS 0.012199f
C1250 VTAIL.n565 VSUBS 0.022702f
C1251 VTAIL.n566 VSUBS 0.022702f
C1252 VTAIL.n567 VSUBS 0.012199f
C1253 VTAIL.n568 VSUBS 0.012917f
C1254 VTAIL.n569 VSUBS 0.028834f
C1255 VTAIL.n570 VSUBS 0.070508f
C1256 VTAIL.n571 VSUBS 0.012917f
C1257 VTAIL.n572 VSUBS 0.023956f
C1258 VTAIL.n573 VSUBS 0.055576f
C1259 VTAIL.n574 VSUBS 0.053411f
C1260 VTAIL.n575 VSUBS 1.35032f
C1261 VP.n0 VSUBS 0.042265f
C1262 VP.t0 VSUBS 2.5188f
C1263 VP.n1 VSUBS 0.061968f
C1264 VP.t2 VSUBS 2.69685f
C1265 VP.t1 VSUBS 2.69532f
C1266 VP.n2 VSUBS 3.56737f
C1267 VP.n3 VSUBS 2.42534f
C1268 VP.t3 VSUBS 2.5188f
C1269 VP.n4 VSUBS 1.00072f
C1270 VP.n5 VSUBS 0.05845f
C1271 VP.n6 VSUBS 0.042265f
C1272 VP.n7 VSUBS 0.042265f
C1273 VP.n8 VSUBS 0.042265f
C1274 VP.n9 VSUBS 0.061968f
C1275 VP.n10 VSUBS 0.05845f
C1276 VP.n11 VSUBS 1.00072f
C1277 VP.n12 VSUBS 0.040788f
.ends

