* NGSPICE file created from diff_pair_sample_1446.ext - technology: sky130A

.subckt diff_pair_sample_1446 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=4.3641 ps=23.16 w=11.19 l=0.65
X1 VDD2.t9 VN.t0 VTAIL.t8 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=4.3641 ps=23.16 w=11.19 l=0.65
X2 VDD1.t8 VP.t1 VTAIL.t14 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=4.3641 ps=23.16 w=11.19 l=0.65
X3 VTAIL.t3 VN.t1 VDD2.t8 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X4 VTAIL.t7 VN.t2 VDD2.t7 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X5 B.t11 B.t9 B.t10 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=0 ps=0 w=11.19 l=0.65
X6 VDD1.t7 VP.t2 VTAIL.t18 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=1.84635 ps=11.52 w=11.19 l=0.65
X7 VDD2.t6 VN.t3 VTAIL.t9 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=1.84635 ps=11.52 w=11.19 l=0.65
X8 B.t8 B.t6 B.t7 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=0 ps=0 w=11.19 l=0.65
X9 VTAIL.t17 VP.t3 VDD1.t6 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X10 VDD2.t5 VN.t4 VTAIL.t1 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=4.3641 ps=23.16 w=11.19 l=0.65
X11 VTAIL.t16 VP.t4 VDD1.t5 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X12 VDD1.t4 VP.t5 VTAIL.t10 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X13 VTAIL.t19 VP.t6 VDD1.t3 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X14 B.t5 B.t3 B.t4 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=0 ps=0 w=11.19 l=0.65
X15 VTAIL.t5 VN.t5 VDD2.t4 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X16 B.t2 B.t0 B.t1 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=0 ps=0 w=11.19 l=0.65
X17 VDD2.t3 VN.t6 VTAIL.t2 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=1.84635 ps=11.52 w=11.19 l=0.65
X18 VDD1.t2 VP.t7 VTAIL.t11 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X19 VDD1.t1 VP.t8 VTAIL.t12 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=4.3641 pd=23.16 as=1.84635 ps=11.52 w=11.19 l=0.65
X20 VDD2.t2 VN.t7 VTAIL.t4 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X21 VDD2.t1 VN.t8 VTAIL.t6 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X22 VTAIL.t0 VN.t9 VDD2.t0 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
X23 VTAIL.t13 VP.t9 VDD1.t0 w_n2146_n3206# sky130_fd_pr__pfet_01v8 ad=1.84635 pd=11.52 as=1.84635 ps=11.52 w=11.19 l=0.65
R0 VP.n4 VP.t2 502.519
R1 VP.n10 VP.t8 475.697
R2 VP.n1 VP.t6 475.697
R3 VP.n14 VP.t5 475.697
R4 VP.n15 VP.t4 475.697
R5 VP.n16 VP.t1 475.697
R6 VP.n8 VP.t0 475.697
R7 VP.n7 VP.t3 475.697
R8 VP.n6 VP.t7 475.697
R9 VP.n5 VP.t9 475.697
R10 VP.n17 VP.n16 161.3
R11 VP.n9 VP.n8 161.3
R12 VP.n11 VP.n10 161.3
R13 VP.n6 VP.n3 80.6037
R14 VP.n7 VP.n2 80.6037
R15 VP.n15 VP.n0 80.6037
R16 VP.n14 VP.n13 80.6037
R17 VP.n12 VP.n1 80.6037
R18 VP.n10 VP.n1 48.2005
R19 VP.n14 VP.n1 48.2005
R20 VP.n15 VP.n14 48.2005
R21 VP.n16 VP.n15 48.2005
R22 VP.n8 VP.n7 48.2005
R23 VP.n7 VP.n6 48.2005
R24 VP.n6 VP.n5 48.2005
R25 VP.n4 VP.n3 45.2318
R26 VP.n11 VP.n9 42.0005
R27 VP.n5 VP.n4 13.3799
R28 VP.n3 VP.n2 0.380177
R29 VP.n13 VP.n12 0.380177
R30 VP.n13 VP.n0 0.380177
R31 VP.n9 VP.n2 0.285035
R32 VP.n12 VP.n11 0.285035
R33 VP.n17 VP.n0 0.285035
R34 VP VP.n17 0.0516364
R35 VTAIL.n11 VTAIL.t1 64.4401
R36 VTAIL.n17 VTAIL.t8 64.44
R37 VTAIL.n2 VTAIL.t14 64.44
R38 VTAIL.n16 VTAIL.t15 64.44
R39 VTAIL.n15 VTAIL.n14 61.5354
R40 VTAIL.n13 VTAIL.n12 61.5354
R41 VTAIL.n10 VTAIL.n9 61.5354
R42 VTAIL.n8 VTAIL.n7 61.5354
R43 VTAIL.n19 VTAIL.n18 61.5351
R44 VTAIL.n1 VTAIL.n0 61.5351
R45 VTAIL.n4 VTAIL.n3 61.5351
R46 VTAIL.n6 VTAIL.n5 61.5351
R47 VTAIL.n8 VTAIL.n6 23.7031
R48 VTAIL.n17 VTAIL.n16 22.8583
R49 VTAIL.n18 VTAIL.t6 2.90533
R50 VTAIL.n18 VTAIL.t7 2.90533
R51 VTAIL.n0 VTAIL.t2 2.90533
R52 VTAIL.n0 VTAIL.t0 2.90533
R53 VTAIL.n3 VTAIL.t10 2.90533
R54 VTAIL.n3 VTAIL.t16 2.90533
R55 VTAIL.n5 VTAIL.t12 2.90533
R56 VTAIL.n5 VTAIL.t19 2.90533
R57 VTAIL.n14 VTAIL.t11 2.90533
R58 VTAIL.n14 VTAIL.t17 2.90533
R59 VTAIL.n12 VTAIL.t18 2.90533
R60 VTAIL.n12 VTAIL.t13 2.90533
R61 VTAIL.n9 VTAIL.t4 2.90533
R62 VTAIL.n9 VTAIL.t3 2.90533
R63 VTAIL.n7 VTAIL.t9 2.90533
R64 VTAIL.n7 VTAIL.t5 2.90533
R65 VTAIL.n13 VTAIL.n11 0.892741
R66 VTAIL.n2 VTAIL.n1 0.892741
R67 VTAIL.n10 VTAIL.n8 0.845328
R68 VTAIL.n11 VTAIL.n10 0.845328
R69 VTAIL.n15 VTAIL.n13 0.845328
R70 VTAIL.n16 VTAIL.n15 0.845328
R71 VTAIL.n6 VTAIL.n4 0.845328
R72 VTAIL.n4 VTAIL.n2 0.845328
R73 VTAIL.n19 VTAIL.n17 0.845328
R74 VTAIL VTAIL.n1 0.69231
R75 VTAIL VTAIL.n19 0.153517
R76 VDD1.n1 VDD1.t7 81.9637
R77 VDD1.n3 VDD1.t1 81.9636
R78 VDD1.n5 VDD1.n4 78.7922
R79 VDD1.n1 VDD1.n0 78.2141
R80 VDD1.n7 VDD1.n6 78.214
R81 VDD1.n3 VDD1.n2 78.2139
R82 VDD1.n7 VDD1.n5 38.3802
R83 VDD1.n6 VDD1.t6 2.90533
R84 VDD1.n6 VDD1.t9 2.90533
R85 VDD1.n0 VDD1.t0 2.90533
R86 VDD1.n0 VDD1.t2 2.90533
R87 VDD1.n4 VDD1.t5 2.90533
R88 VDD1.n4 VDD1.t8 2.90533
R89 VDD1.n2 VDD1.t3 2.90533
R90 VDD1.n2 VDD1.t4 2.90533
R91 VDD1 VDD1.n7 0.575931
R92 VDD1 VDD1.n1 0.269897
R93 VDD1.n5 VDD1.n3 0.156361
R94 VN.n2 VN.t6 502.519
R95 VN.n10 VN.t4 502.519
R96 VN.n1 VN.t9 475.697
R97 VN.n4 VN.t8 475.697
R98 VN.n5 VN.t2 475.697
R99 VN.n6 VN.t0 475.697
R100 VN.n9 VN.t1 475.697
R101 VN.n12 VN.t7 475.697
R102 VN.n13 VN.t5 475.697
R103 VN.n14 VN.t3 475.697
R104 VN.n7 VN.n6 161.3
R105 VN.n15 VN.n14 161.3
R106 VN.n13 VN.n8 80.6037
R107 VN.n12 VN.n11 80.6037
R108 VN.n5 VN.n0 80.6037
R109 VN.n4 VN.n3 80.6037
R110 VN.n4 VN.n1 48.2005
R111 VN.n5 VN.n4 48.2005
R112 VN.n6 VN.n5 48.2005
R113 VN.n12 VN.n9 48.2005
R114 VN.n13 VN.n12 48.2005
R115 VN.n14 VN.n13 48.2005
R116 VN.n11 VN.n10 45.2318
R117 VN.n3 VN.n2 45.2318
R118 VN VN.n15 42.3812
R119 VN.n10 VN.n9 13.3799
R120 VN.n2 VN.n1 13.3799
R121 VN.n11 VN.n8 0.380177
R122 VN.n3 VN.n0 0.380177
R123 VN.n15 VN.n8 0.285035
R124 VN.n7 VN.n0 0.285035
R125 VN VN.n7 0.0516364
R126 VDD2.n1 VDD2.t3 81.9636
R127 VDD2.n4 VDD2.t6 81.1189
R128 VDD2.n3 VDD2.n2 78.7922
R129 VDD2 VDD2.n7 78.7894
R130 VDD2.n6 VDD2.n5 78.2141
R131 VDD2.n1 VDD2.n0 78.2139
R132 VDD2.n4 VDD2.n3 37.3748
R133 VDD2.n7 VDD2.t8 2.90533
R134 VDD2.n7 VDD2.t5 2.90533
R135 VDD2.n5 VDD2.t4 2.90533
R136 VDD2.n5 VDD2.t2 2.90533
R137 VDD2.n2 VDD2.t7 2.90533
R138 VDD2.n2 VDD2.t9 2.90533
R139 VDD2.n0 VDD2.t0 2.90533
R140 VDD2.n0 VDD2.t1 2.90533
R141 VDD2.n6 VDD2.n4 0.845328
R142 VDD2 VDD2.n6 0.269897
R143 VDD2.n3 VDD2.n1 0.156361
R144 B.n114 B.t9 618.519
R145 B.n256 B.t6 618.519
R146 B.n42 B.t3 618.519
R147 B.n34 B.t0 618.519
R148 B.n318 B.n89 585
R149 B.n317 B.n316 585
R150 B.n315 B.n90 585
R151 B.n314 B.n313 585
R152 B.n312 B.n91 585
R153 B.n311 B.n310 585
R154 B.n309 B.n92 585
R155 B.n308 B.n307 585
R156 B.n306 B.n93 585
R157 B.n305 B.n304 585
R158 B.n303 B.n94 585
R159 B.n302 B.n301 585
R160 B.n300 B.n95 585
R161 B.n299 B.n298 585
R162 B.n297 B.n96 585
R163 B.n296 B.n295 585
R164 B.n294 B.n97 585
R165 B.n293 B.n292 585
R166 B.n291 B.n98 585
R167 B.n290 B.n289 585
R168 B.n288 B.n99 585
R169 B.n287 B.n286 585
R170 B.n285 B.n100 585
R171 B.n284 B.n283 585
R172 B.n282 B.n101 585
R173 B.n281 B.n280 585
R174 B.n279 B.n102 585
R175 B.n278 B.n277 585
R176 B.n276 B.n103 585
R177 B.n275 B.n274 585
R178 B.n273 B.n104 585
R179 B.n272 B.n271 585
R180 B.n270 B.n105 585
R181 B.n269 B.n268 585
R182 B.n267 B.n106 585
R183 B.n266 B.n265 585
R184 B.n264 B.n107 585
R185 B.n263 B.n262 585
R186 B.n261 B.n108 585
R187 B.n260 B.n259 585
R188 B.n255 B.n109 585
R189 B.n254 B.n253 585
R190 B.n252 B.n110 585
R191 B.n251 B.n250 585
R192 B.n249 B.n111 585
R193 B.n248 B.n247 585
R194 B.n246 B.n112 585
R195 B.n245 B.n244 585
R196 B.n243 B.n113 585
R197 B.n241 B.n240 585
R198 B.n239 B.n116 585
R199 B.n238 B.n237 585
R200 B.n236 B.n117 585
R201 B.n235 B.n234 585
R202 B.n233 B.n118 585
R203 B.n232 B.n231 585
R204 B.n230 B.n119 585
R205 B.n229 B.n228 585
R206 B.n227 B.n120 585
R207 B.n226 B.n225 585
R208 B.n224 B.n121 585
R209 B.n223 B.n222 585
R210 B.n221 B.n122 585
R211 B.n220 B.n219 585
R212 B.n218 B.n123 585
R213 B.n217 B.n216 585
R214 B.n215 B.n124 585
R215 B.n214 B.n213 585
R216 B.n212 B.n125 585
R217 B.n211 B.n210 585
R218 B.n209 B.n126 585
R219 B.n208 B.n207 585
R220 B.n206 B.n127 585
R221 B.n205 B.n204 585
R222 B.n203 B.n128 585
R223 B.n202 B.n201 585
R224 B.n200 B.n129 585
R225 B.n199 B.n198 585
R226 B.n197 B.n130 585
R227 B.n196 B.n195 585
R228 B.n194 B.n131 585
R229 B.n193 B.n192 585
R230 B.n191 B.n132 585
R231 B.n190 B.n189 585
R232 B.n188 B.n133 585
R233 B.n187 B.n186 585
R234 B.n185 B.n134 585
R235 B.n184 B.n183 585
R236 B.n320 B.n319 585
R237 B.n321 B.n88 585
R238 B.n323 B.n322 585
R239 B.n324 B.n87 585
R240 B.n326 B.n325 585
R241 B.n327 B.n86 585
R242 B.n329 B.n328 585
R243 B.n330 B.n85 585
R244 B.n332 B.n331 585
R245 B.n333 B.n84 585
R246 B.n335 B.n334 585
R247 B.n336 B.n83 585
R248 B.n338 B.n337 585
R249 B.n339 B.n82 585
R250 B.n341 B.n340 585
R251 B.n342 B.n81 585
R252 B.n344 B.n343 585
R253 B.n345 B.n80 585
R254 B.n347 B.n346 585
R255 B.n348 B.n79 585
R256 B.n350 B.n349 585
R257 B.n351 B.n78 585
R258 B.n353 B.n352 585
R259 B.n354 B.n77 585
R260 B.n356 B.n355 585
R261 B.n357 B.n76 585
R262 B.n359 B.n358 585
R263 B.n360 B.n75 585
R264 B.n362 B.n361 585
R265 B.n363 B.n74 585
R266 B.n365 B.n364 585
R267 B.n366 B.n73 585
R268 B.n368 B.n367 585
R269 B.n369 B.n72 585
R270 B.n371 B.n370 585
R271 B.n372 B.n71 585
R272 B.n374 B.n373 585
R273 B.n375 B.n70 585
R274 B.n377 B.n376 585
R275 B.n378 B.n69 585
R276 B.n380 B.n379 585
R277 B.n381 B.n68 585
R278 B.n383 B.n382 585
R279 B.n384 B.n67 585
R280 B.n386 B.n385 585
R281 B.n387 B.n66 585
R282 B.n389 B.n388 585
R283 B.n390 B.n65 585
R284 B.n392 B.n391 585
R285 B.n393 B.n64 585
R286 B.n395 B.n394 585
R287 B.n396 B.n63 585
R288 B.n530 B.n529 585
R289 B.n528 B.n15 585
R290 B.n527 B.n526 585
R291 B.n525 B.n16 585
R292 B.n524 B.n523 585
R293 B.n522 B.n17 585
R294 B.n521 B.n520 585
R295 B.n519 B.n18 585
R296 B.n518 B.n517 585
R297 B.n516 B.n19 585
R298 B.n515 B.n514 585
R299 B.n513 B.n20 585
R300 B.n512 B.n511 585
R301 B.n510 B.n21 585
R302 B.n509 B.n508 585
R303 B.n507 B.n22 585
R304 B.n506 B.n505 585
R305 B.n504 B.n23 585
R306 B.n503 B.n502 585
R307 B.n501 B.n24 585
R308 B.n500 B.n499 585
R309 B.n498 B.n25 585
R310 B.n497 B.n496 585
R311 B.n495 B.n26 585
R312 B.n494 B.n493 585
R313 B.n492 B.n27 585
R314 B.n491 B.n490 585
R315 B.n489 B.n28 585
R316 B.n488 B.n487 585
R317 B.n486 B.n29 585
R318 B.n485 B.n484 585
R319 B.n483 B.n30 585
R320 B.n482 B.n481 585
R321 B.n480 B.n31 585
R322 B.n479 B.n478 585
R323 B.n477 B.n32 585
R324 B.n476 B.n475 585
R325 B.n474 B.n33 585
R326 B.n473 B.n472 585
R327 B.n471 B.n470 585
R328 B.n469 B.n37 585
R329 B.n468 B.n467 585
R330 B.n466 B.n38 585
R331 B.n465 B.n464 585
R332 B.n463 B.n39 585
R333 B.n462 B.n461 585
R334 B.n460 B.n40 585
R335 B.n459 B.n458 585
R336 B.n457 B.n41 585
R337 B.n455 B.n454 585
R338 B.n453 B.n44 585
R339 B.n452 B.n451 585
R340 B.n450 B.n45 585
R341 B.n449 B.n448 585
R342 B.n447 B.n46 585
R343 B.n446 B.n445 585
R344 B.n444 B.n47 585
R345 B.n443 B.n442 585
R346 B.n441 B.n48 585
R347 B.n440 B.n439 585
R348 B.n438 B.n49 585
R349 B.n437 B.n436 585
R350 B.n435 B.n50 585
R351 B.n434 B.n433 585
R352 B.n432 B.n51 585
R353 B.n431 B.n430 585
R354 B.n429 B.n52 585
R355 B.n428 B.n427 585
R356 B.n426 B.n53 585
R357 B.n425 B.n424 585
R358 B.n423 B.n54 585
R359 B.n422 B.n421 585
R360 B.n420 B.n55 585
R361 B.n419 B.n418 585
R362 B.n417 B.n56 585
R363 B.n416 B.n415 585
R364 B.n414 B.n57 585
R365 B.n413 B.n412 585
R366 B.n411 B.n58 585
R367 B.n410 B.n409 585
R368 B.n408 B.n59 585
R369 B.n407 B.n406 585
R370 B.n405 B.n60 585
R371 B.n404 B.n403 585
R372 B.n402 B.n61 585
R373 B.n401 B.n400 585
R374 B.n399 B.n62 585
R375 B.n398 B.n397 585
R376 B.n531 B.n14 585
R377 B.n533 B.n532 585
R378 B.n534 B.n13 585
R379 B.n536 B.n535 585
R380 B.n537 B.n12 585
R381 B.n539 B.n538 585
R382 B.n540 B.n11 585
R383 B.n542 B.n541 585
R384 B.n543 B.n10 585
R385 B.n545 B.n544 585
R386 B.n546 B.n9 585
R387 B.n548 B.n547 585
R388 B.n549 B.n8 585
R389 B.n551 B.n550 585
R390 B.n552 B.n7 585
R391 B.n554 B.n553 585
R392 B.n555 B.n6 585
R393 B.n557 B.n556 585
R394 B.n558 B.n5 585
R395 B.n560 B.n559 585
R396 B.n561 B.n4 585
R397 B.n563 B.n562 585
R398 B.n564 B.n3 585
R399 B.n566 B.n565 585
R400 B.n567 B.n0 585
R401 B.n2 B.n1 585
R402 B.n148 B.n147 585
R403 B.n149 B.n146 585
R404 B.n151 B.n150 585
R405 B.n152 B.n145 585
R406 B.n154 B.n153 585
R407 B.n155 B.n144 585
R408 B.n157 B.n156 585
R409 B.n158 B.n143 585
R410 B.n160 B.n159 585
R411 B.n161 B.n142 585
R412 B.n163 B.n162 585
R413 B.n164 B.n141 585
R414 B.n166 B.n165 585
R415 B.n167 B.n140 585
R416 B.n169 B.n168 585
R417 B.n170 B.n139 585
R418 B.n172 B.n171 585
R419 B.n173 B.n138 585
R420 B.n175 B.n174 585
R421 B.n176 B.n137 585
R422 B.n178 B.n177 585
R423 B.n179 B.n136 585
R424 B.n181 B.n180 585
R425 B.n182 B.n135 585
R426 B.n184 B.n135 487.695
R427 B.n320 B.n89 487.695
R428 B.n398 B.n63 487.695
R429 B.n531 B.n530 487.695
R430 B.n569 B.n568 256.663
R431 B.n568 B.n567 235.042
R432 B.n568 B.n2 235.042
R433 B.n185 B.n184 163.367
R434 B.n186 B.n185 163.367
R435 B.n186 B.n133 163.367
R436 B.n190 B.n133 163.367
R437 B.n191 B.n190 163.367
R438 B.n192 B.n191 163.367
R439 B.n192 B.n131 163.367
R440 B.n196 B.n131 163.367
R441 B.n197 B.n196 163.367
R442 B.n198 B.n197 163.367
R443 B.n198 B.n129 163.367
R444 B.n202 B.n129 163.367
R445 B.n203 B.n202 163.367
R446 B.n204 B.n203 163.367
R447 B.n204 B.n127 163.367
R448 B.n208 B.n127 163.367
R449 B.n209 B.n208 163.367
R450 B.n210 B.n209 163.367
R451 B.n210 B.n125 163.367
R452 B.n214 B.n125 163.367
R453 B.n215 B.n214 163.367
R454 B.n216 B.n215 163.367
R455 B.n216 B.n123 163.367
R456 B.n220 B.n123 163.367
R457 B.n221 B.n220 163.367
R458 B.n222 B.n221 163.367
R459 B.n222 B.n121 163.367
R460 B.n226 B.n121 163.367
R461 B.n227 B.n226 163.367
R462 B.n228 B.n227 163.367
R463 B.n228 B.n119 163.367
R464 B.n232 B.n119 163.367
R465 B.n233 B.n232 163.367
R466 B.n234 B.n233 163.367
R467 B.n234 B.n117 163.367
R468 B.n238 B.n117 163.367
R469 B.n239 B.n238 163.367
R470 B.n240 B.n239 163.367
R471 B.n240 B.n113 163.367
R472 B.n245 B.n113 163.367
R473 B.n246 B.n245 163.367
R474 B.n247 B.n246 163.367
R475 B.n247 B.n111 163.367
R476 B.n251 B.n111 163.367
R477 B.n252 B.n251 163.367
R478 B.n253 B.n252 163.367
R479 B.n253 B.n109 163.367
R480 B.n260 B.n109 163.367
R481 B.n261 B.n260 163.367
R482 B.n262 B.n261 163.367
R483 B.n262 B.n107 163.367
R484 B.n266 B.n107 163.367
R485 B.n267 B.n266 163.367
R486 B.n268 B.n267 163.367
R487 B.n268 B.n105 163.367
R488 B.n272 B.n105 163.367
R489 B.n273 B.n272 163.367
R490 B.n274 B.n273 163.367
R491 B.n274 B.n103 163.367
R492 B.n278 B.n103 163.367
R493 B.n279 B.n278 163.367
R494 B.n280 B.n279 163.367
R495 B.n280 B.n101 163.367
R496 B.n284 B.n101 163.367
R497 B.n285 B.n284 163.367
R498 B.n286 B.n285 163.367
R499 B.n286 B.n99 163.367
R500 B.n290 B.n99 163.367
R501 B.n291 B.n290 163.367
R502 B.n292 B.n291 163.367
R503 B.n292 B.n97 163.367
R504 B.n296 B.n97 163.367
R505 B.n297 B.n296 163.367
R506 B.n298 B.n297 163.367
R507 B.n298 B.n95 163.367
R508 B.n302 B.n95 163.367
R509 B.n303 B.n302 163.367
R510 B.n304 B.n303 163.367
R511 B.n304 B.n93 163.367
R512 B.n308 B.n93 163.367
R513 B.n309 B.n308 163.367
R514 B.n310 B.n309 163.367
R515 B.n310 B.n91 163.367
R516 B.n314 B.n91 163.367
R517 B.n315 B.n314 163.367
R518 B.n316 B.n315 163.367
R519 B.n316 B.n89 163.367
R520 B.n394 B.n63 163.367
R521 B.n394 B.n393 163.367
R522 B.n393 B.n392 163.367
R523 B.n392 B.n65 163.367
R524 B.n388 B.n65 163.367
R525 B.n388 B.n387 163.367
R526 B.n387 B.n386 163.367
R527 B.n386 B.n67 163.367
R528 B.n382 B.n67 163.367
R529 B.n382 B.n381 163.367
R530 B.n381 B.n380 163.367
R531 B.n380 B.n69 163.367
R532 B.n376 B.n69 163.367
R533 B.n376 B.n375 163.367
R534 B.n375 B.n374 163.367
R535 B.n374 B.n71 163.367
R536 B.n370 B.n71 163.367
R537 B.n370 B.n369 163.367
R538 B.n369 B.n368 163.367
R539 B.n368 B.n73 163.367
R540 B.n364 B.n73 163.367
R541 B.n364 B.n363 163.367
R542 B.n363 B.n362 163.367
R543 B.n362 B.n75 163.367
R544 B.n358 B.n75 163.367
R545 B.n358 B.n357 163.367
R546 B.n357 B.n356 163.367
R547 B.n356 B.n77 163.367
R548 B.n352 B.n77 163.367
R549 B.n352 B.n351 163.367
R550 B.n351 B.n350 163.367
R551 B.n350 B.n79 163.367
R552 B.n346 B.n79 163.367
R553 B.n346 B.n345 163.367
R554 B.n345 B.n344 163.367
R555 B.n344 B.n81 163.367
R556 B.n340 B.n81 163.367
R557 B.n340 B.n339 163.367
R558 B.n339 B.n338 163.367
R559 B.n338 B.n83 163.367
R560 B.n334 B.n83 163.367
R561 B.n334 B.n333 163.367
R562 B.n333 B.n332 163.367
R563 B.n332 B.n85 163.367
R564 B.n328 B.n85 163.367
R565 B.n328 B.n327 163.367
R566 B.n327 B.n326 163.367
R567 B.n326 B.n87 163.367
R568 B.n322 B.n87 163.367
R569 B.n322 B.n321 163.367
R570 B.n321 B.n320 163.367
R571 B.n530 B.n15 163.367
R572 B.n526 B.n15 163.367
R573 B.n526 B.n525 163.367
R574 B.n525 B.n524 163.367
R575 B.n524 B.n17 163.367
R576 B.n520 B.n17 163.367
R577 B.n520 B.n519 163.367
R578 B.n519 B.n518 163.367
R579 B.n518 B.n19 163.367
R580 B.n514 B.n19 163.367
R581 B.n514 B.n513 163.367
R582 B.n513 B.n512 163.367
R583 B.n512 B.n21 163.367
R584 B.n508 B.n21 163.367
R585 B.n508 B.n507 163.367
R586 B.n507 B.n506 163.367
R587 B.n506 B.n23 163.367
R588 B.n502 B.n23 163.367
R589 B.n502 B.n501 163.367
R590 B.n501 B.n500 163.367
R591 B.n500 B.n25 163.367
R592 B.n496 B.n25 163.367
R593 B.n496 B.n495 163.367
R594 B.n495 B.n494 163.367
R595 B.n494 B.n27 163.367
R596 B.n490 B.n27 163.367
R597 B.n490 B.n489 163.367
R598 B.n489 B.n488 163.367
R599 B.n488 B.n29 163.367
R600 B.n484 B.n29 163.367
R601 B.n484 B.n483 163.367
R602 B.n483 B.n482 163.367
R603 B.n482 B.n31 163.367
R604 B.n478 B.n31 163.367
R605 B.n478 B.n477 163.367
R606 B.n477 B.n476 163.367
R607 B.n476 B.n33 163.367
R608 B.n472 B.n33 163.367
R609 B.n472 B.n471 163.367
R610 B.n471 B.n37 163.367
R611 B.n467 B.n37 163.367
R612 B.n467 B.n466 163.367
R613 B.n466 B.n465 163.367
R614 B.n465 B.n39 163.367
R615 B.n461 B.n39 163.367
R616 B.n461 B.n460 163.367
R617 B.n460 B.n459 163.367
R618 B.n459 B.n41 163.367
R619 B.n454 B.n41 163.367
R620 B.n454 B.n453 163.367
R621 B.n453 B.n452 163.367
R622 B.n452 B.n45 163.367
R623 B.n448 B.n45 163.367
R624 B.n448 B.n447 163.367
R625 B.n447 B.n446 163.367
R626 B.n446 B.n47 163.367
R627 B.n442 B.n47 163.367
R628 B.n442 B.n441 163.367
R629 B.n441 B.n440 163.367
R630 B.n440 B.n49 163.367
R631 B.n436 B.n49 163.367
R632 B.n436 B.n435 163.367
R633 B.n435 B.n434 163.367
R634 B.n434 B.n51 163.367
R635 B.n430 B.n51 163.367
R636 B.n430 B.n429 163.367
R637 B.n429 B.n428 163.367
R638 B.n428 B.n53 163.367
R639 B.n424 B.n53 163.367
R640 B.n424 B.n423 163.367
R641 B.n423 B.n422 163.367
R642 B.n422 B.n55 163.367
R643 B.n418 B.n55 163.367
R644 B.n418 B.n417 163.367
R645 B.n417 B.n416 163.367
R646 B.n416 B.n57 163.367
R647 B.n412 B.n57 163.367
R648 B.n412 B.n411 163.367
R649 B.n411 B.n410 163.367
R650 B.n410 B.n59 163.367
R651 B.n406 B.n59 163.367
R652 B.n406 B.n405 163.367
R653 B.n405 B.n404 163.367
R654 B.n404 B.n61 163.367
R655 B.n400 B.n61 163.367
R656 B.n400 B.n399 163.367
R657 B.n399 B.n398 163.367
R658 B.n532 B.n531 163.367
R659 B.n532 B.n13 163.367
R660 B.n536 B.n13 163.367
R661 B.n537 B.n536 163.367
R662 B.n538 B.n537 163.367
R663 B.n538 B.n11 163.367
R664 B.n542 B.n11 163.367
R665 B.n543 B.n542 163.367
R666 B.n544 B.n543 163.367
R667 B.n544 B.n9 163.367
R668 B.n548 B.n9 163.367
R669 B.n549 B.n548 163.367
R670 B.n550 B.n549 163.367
R671 B.n550 B.n7 163.367
R672 B.n554 B.n7 163.367
R673 B.n555 B.n554 163.367
R674 B.n556 B.n555 163.367
R675 B.n556 B.n5 163.367
R676 B.n560 B.n5 163.367
R677 B.n561 B.n560 163.367
R678 B.n562 B.n561 163.367
R679 B.n562 B.n3 163.367
R680 B.n566 B.n3 163.367
R681 B.n567 B.n566 163.367
R682 B.n148 B.n2 163.367
R683 B.n149 B.n148 163.367
R684 B.n150 B.n149 163.367
R685 B.n150 B.n145 163.367
R686 B.n154 B.n145 163.367
R687 B.n155 B.n154 163.367
R688 B.n156 B.n155 163.367
R689 B.n156 B.n143 163.367
R690 B.n160 B.n143 163.367
R691 B.n161 B.n160 163.367
R692 B.n162 B.n161 163.367
R693 B.n162 B.n141 163.367
R694 B.n166 B.n141 163.367
R695 B.n167 B.n166 163.367
R696 B.n168 B.n167 163.367
R697 B.n168 B.n139 163.367
R698 B.n172 B.n139 163.367
R699 B.n173 B.n172 163.367
R700 B.n174 B.n173 163.367
R701 B.n174 B.n137 163.367
R702 B.n178 B.n137 163.367
R703 B.n179 B.n178 163.367
R704 B.n180 B.n179 163.367
R705 B.n180 B.n135 163.367
R706 B.n256 B.t7 132.327
R707 B.n42 B.t5 132.327
R708 B.n114 B.t10 132.315
R709 B.n34 B.t2 132.315
R710 B.n257 B.t8 113.32
R711 B.n43 B.t4 113.32
R712 B.n115 B.t11 113.308
R713 B.n35 B.t1 113.308
R714 B.n242 B.n115 59.5399
R715 B.n258 B.n257 59.5399
R716 B.n456 B.n43 59.5399
R717 B.n36 B.n35 59.5399
R718 B.n529 B.n14 31.6883
R719 B.n397 B.n396 31.6883
R720 B.n319 B.n318 31.6883
R721 B.n183 B.n182 31.6883
R722 B.n115 B.n114 19.0066
R723 B.n257 B.n256 19.0066
R724 B.n43 B.n42 19.0066
R725 B.n35 B.n34 19.0066
R726 B B.n569 18.0485
R727 B.n533 B.n14 10.6151
R728 B.n534 B.n533 10.6151
R729 B.n535 B.n534 10.6151
R730 B.n535 B.n12 10.6151
R731 B.n539 B.n12 10.6151
R732 B.n540 B.n539 10.6151
R733 B.n541 B.n540 10.6151
R734 B.n541 B.n10 10.6151
R735 B.n545 B.n10 10.6151
R736 B.n546 B.n545 10.6151
R737 B.n547 B.n546 10.6151
R738 B.n547 B.n8 10.6151
R739 B.n551 B.n8 10.6151
R740 B.n552 B.n551 10.6151
R741 B.n553 B.n552 10.6151
R742 B.n553 B.n6 10.6151
R743 B.n557 B.n6 10.6151
R744 B.n558 B.n557 10.6151
R745 B.n559 B.n558 10.6151
R746 B.n559 B.n4 10.6151
R747 B.n563 B.n4 10.6151
R748 B.n564 B.n563 10.6151
R749 B.n565 B.n564 10.6151
R750 B.n565 B.n0 10.6151
R751 B.n529 B.n528 10.6151
R752 B.n528 B.n527 10.6151
R753 B.n527 B.n16 10.6151
R754 B.n523 B.n16 10.6151
R755 B.n523 B.n522 10.6151
R756 B.n522 B.n521 10.6151
R757 B.n521 B.n18 10.6151
R758 B.n517 B.n18 10.6151
R759 B.n517 B.n516 10.6151
R760 B.n516 B.n515 10.6151
R761 B.n515 B.n20 10.6151
R762 B.n511 B.n20 10.6151
R763 B.n511 B.n510 10.6151
R764 B.n510 B.n509 10.6151
R765 B.n509 B.n22 10.6151
R766 B.n505 B.n22 10.6151
R767 B.n505 B.n504 10.6151
R768 B.n504 B.n503 10.6151
R769 B.n503 B.n24 10.6151
R770 B.n499 B.n24 10.6151
R771 B.n499 B.n498 10.6151
R772 B.n498 B.n497 10.6151
R773 B.n497 B.n26 10.6151
R774 B.n493 B.n26 10.6151
R775 B.n493 B.n492 10.6151
R776 B.n492 B.n491 10.6151
R777 B.n491 B.n28 10.6151
R778 B.n487 B.n28 10.6151
R779 B.n487 B.n486 10.6151
R780 B.n486 B.n485 10.6151
R781 B.n485 B.n30 10.6151
R782 B.n481 B.n30 10.6151
R783 B.n481 B.n480 10.6151
R784 B.n480 B.n479 10.6151
R785 B.n479 B.n32 10.6151
R786 B.n475 B.n32 10.6151
R787 B.n475 B.n474 10.6151
R788 B.n474 B.n473 10.6151
R789 B.n470 B.n469 10.6151
R790 B.n469 B.n468 10.6151
R791 B.n468 B.n38 10.6151
R792 B.n464 B.n38 10.6151
R793 B.n464 B.n463 10.6151
R794 B.n463 B.n462 10.6151
R795 B.n462 B.n40 10.6151
R796 B.n458 B.n40 10.6151
R797 B.n458 B.n457 10.6151
R798 B.n455 B.n44 10.6151
R799 B.n451 B.n44 10.6151
R800 B.n451 B.n450 10.6151
R801 B.n450 B.n449 10.6151
R802 B.n449 B.n46 10.6151
R803 B.n445 B.n46 10.6151
R804 B.n445 B.n444 10.6151
R805 B.n444 B.n443 10.6151
R806 B.n443 B.n48 10.6151
R807 B.n439 B.n48 10.6151
R808 B.n439 B.n438 10.6151
R809 B.n438 B.n437 10.6151
R810 B.n437 B.n50 10.6151
R811 B.n433 B.n50 10.6151
R812 B.n433 B.n432 10.6151
R813 B.n432 B.n431 10.6151
R814 B.n431 B.n52 10.6151
R815 B.n427 B.n52 10.6151
R816 B.n427 B.n426 10.6151
R817 B.n426 B.n425 10.6151
R818 B.n425 B.n54 10.6151
R819 B.n421 B.n54 10.6151
R820 B.n421 B.n420 10.6151
R821 B.n420 B.n419 10.6151
R822 B.n419 B.n56 10.6151
R823 B.n415 B.n56 10.6151
R824 B.n415 B.n414 10.6151
R825 B.n414 B.n413 10.6151
R826 B.n413 B.n58 10.6151
R827 B.n409 B.n58 10.6151
R828 B.n409 B.n408 10.6151
R829 B.n408 B.n407 10.6151
R830 B.n407 B.n60 10.6151
R831 B.n403 B.n60 10.6151
R832 B.n403 B.n402 10.6151
R833 B.n402 B.n401 10.6151
R834 B.n401 B.n62 10.6151
R835 B.n397 B.n62 10.6151
R836 B.n396 B.n395 10.6151
R837 B.n395 B.n64 10.6151
R838 B.n391 B.n64 10.6151
R839 B.n391 B.n390 10.6151
R840 B.n390 B.n389 10.6151
R841 B.n389 B.n66 10.6151
R842 B.n385 B.n66 10.6151
R843 B.n385 B.n384 10.6151
R844 B.n384 B.n383 10.6151
R845 B.n383 B.n68 10.6151
R846 B.n379 B.n68 10.6151
R847 B.n379 B.n378 10.6151
R848 B.n378 B.n377 10.6151
R849 B.n377 B.n70 10.6151
R850 B.n373 B.n70 10.6151
R851 B.n373 B.n372 10.6151
R852 B.n372 B.n371 10.6151
R853 B.n371 B.n72 10.6151
R854 B.n367 B.n72 10.6151
R855 B.n367 B.n366 10.6151
R856 B.n366 B.n365 10.6151
R857 B.n365 B.n74 10.6151
R858 B.n361 B.n74 10.6151
R859 B.n361 B.n360 10.6151
R860 B.n360 B.n359 10.6151
R861 B.n359 B.n76 10.6151
R862 B.n355 B.n76 10.6151
R863 B.n355 B.n354 10.6151
R864 B.n354 B.n353 10.6151
R865 B.n353 B.n78 10.6151
R866 B.n349 B.n78 10.6151
R867 B.n349 B.n348 10.6151
R868 B.n348 B.n347 10.6151
R869 B.n347 B.n80 10.6151
R870 B.n343 B.n80 10.6151
R871 B.n343 B.n342 10.6151
R872 B.n342 B.n341 10.6151
R873 B.n341 B.n82 10.6151
R874 B.n337 B.n82 10.6151
R875 B.n337 B.n336 10.6151
R876 B.n336 B.n335 10.6151
R877 B.n335 B.n84 10.6151
R878 B.n331 B.n84 10.6151
R879 B.n331 B.n330 10.6151
R880 B.n330 B.n329 10.6151
R881 B.n329 B.n86 10.6151
R882 B.n325 B.n86 10.6151
R883 B.n325 B.n324 10.6151
R884 B.n324 B.n323 10.6151
R885 B.n323 B.n88 10.6151
R886 B.n319 B.n88 10.6151
R887 B.n147 B.n1 10.6151
R888 B.n147 B.n146 10.6151
R889 B.n151 B.n146 10.6151
R890 B.n152 B.n151 10.6151
R891 B.n153 B.n152 10.6151
R892 B.n153 B.n144 10.6151
R893 B.n157 B.n144 10.6151
R894 B.n158 B.n157 10.6151
R895 B.n159 B.n158 10.6151
R896 B.n159 B.n142 10.6151
R897 B.n163 B.n142 10.6151
R898 B.n164 B.n163 10.6151
R899 B.n165 B.n164 10.6151
R900 B.n165 B.n140 10.6151
R901 B.n169 B.n140 10.6151
R902 B.n170 B.n169 10.6151
R903 B.n171 B.n170 10.6151
R904 B.n171 B.n138 10.6151
R905 B.n175 B.n138 10.6151
R906 B.n176 B.n175 10.6151
R907 B.n177 B.n176 10.6151
R908 B.n177 B.n136 10.6151
R909 B.n181 B.n136 10.6151
R910 B.n182 B.n181 10.6151
R911 B.n183 B.n134 10.6151
R912 B.n187 B.n134 10.6151
R913 B.n188 B.n187 10.6151
R914 B.n189 B.n188 10.6151
R915 B.n189 B.n132 10.6151
R916 B.n193 B.n132 10.6151
R917 B.n194 B.n193 10.6151
R918 B.n195 B.n194 10.6151
R919 B.n195 B.n130 10.6151
R920 B.n199 B.n130 10.6151
R921 B.n200 B.n199 10.6151
R922 B.n201 B.n200 10.6151
R923 B.n201 B.n128 10.6151
R924 B.n205 B.n128 10.6151
R925 B.n206 B.n205 10.6151
R926 B.n207 B.n206 10.6151
R927 B.n207 B.n126 10.6151
R928 B.n211 B.n126 10.6151
R929 B.n212 B.n211 10.6151
R930 B.n213 B.n212 10.6151
R931 B.n213 B.n124 10.6151
R932 B.n217 B.n124 10.6151
R933 B.n218 B.n217 10.6151
R934 B.n219 B.n218 10.6151
R935 B.n219 B.n122 10.6151
R936 B.n223 B.n122 10.6151
R937 B.n224 B.n223 10.6151
R938 B.n225 B.n224 10.6151
R939 B.n225 B.n120 10.6151
R940 B.n229 B.n120 10.6151
R941 B.n230 B.n229 10.6151
R942 B.n231 B.n230 10.6151
R943 B.n231 B.n118 10.6151
R944 B.n235 B.n118 10.6151
R945 B.n236 B.n235 10.6151
R946 B.n237 B.n236 10.6151
R947 B.n237 B.n116 10.6151
R948 B.n241 B.n116 10.6151
R949 B.n244 B.n243 10.6151
R950 B.n244 B.n112 10.6151
R951 B.n248 B.n112 10.6151
R952 B.n249 B.n248 10.6151
R953 B.n250 B.n249 10.6151
R954 B.n250 B.n110 10.6151
R955 B.n254 B.n110 10.6151
R956 B.n255 B.n254 10.6151
R957 B.n259 B.n255 10.6151
R958 B.n263 B.n108 10.6151
R959 B.n264 B.n263 10.6151
R960 B.n265 B.n264 10.6151
R961 B.n265 B.n106 10.6151
R962 B.n269 B.n106 10.6151
R963 B.n270 B.n269 10.6151
R964 B.n271 B.n270 10.6151
R965 B.n271 B.n104 10.6151
R966 B.n275 B.n104 10.6151
R967 B.n276 B.n275 10.6151
R968 B.n277 B.n276 10.6151
R969 B.n277 B.n102 10.6151
R970 B.n281 B.n102 10.6151
R971 B.n282 B.n281 10.6151
R972 B.n283 B.n282 10.6151
R973 B.n283 B.n100 10.6151
R974 B.n287 B.n100 10.6151
R975 B.n288 B.n287 10.6151
R976 B.n289 B.n288 10.6151
R977 B.n289 B.n98 10.6151
R978 B.n293 B.n98 10.6151
R979 B.n294 B.n293 10.6151
R980 B.n295 B.n294 10.6151
R981 B.n295 B.n96 10.6151
R982 B.n299 B.n96 10.6151
R983 B.n300 B.n299 10.6151
R984 B.n301 B.n300 10.6151
R985 B.n301 B.n94 10.6151
R986 B.n305 B.n94 10.6151
R987 B.n306 B.n305 10.6151
R988 B.n307 B.n306 10.6151
R989 B.n307 B.n92 10.6151
R990 B.n311 B.n92 10.6151
R991 B.n312 B.n311 10.6151
R992 B.n313 B.n312 10.6151
R993 B.n313 B.n90 10.6151
R994 B.n317 B.n90 10.6151
R995 B.n318 B.n317 10.6151
R996 B.n473 B.n36 9.36635
R997 B.n456 B.n455 9.36635
R998 B.n242 B.n241 9.36635
R999 B.n258 B.n108 9.36635
R1000 B.n569 B.n0 8.11757
R1001 B.n569 B.n1 8.11757
R1002 B.n470 B.n36 1.24928
R1003 B.n457 B.n456 1.24928
R1004 B.n243 B.n242 1.24928
R1005 B.n259 B.n258 1.24928
C0 VDD1 VP 6.19799f
C1 VTAIL VN 5.85774f
C2 VN VDD1 0.14903f
C3 VTAIL VDD1 13.859099f
C4 VDD2 w_n2146_n3206# 2.00371f
C5 VDD2 B 1.6652f
C6 B w_n2146_n3206# 7.04358f
C7 VDD2 VP 0.335225f
C8 w_n2146_n3206# VP 4.24059f
C9 VDD2 VN 6.01627f
C10 VN w_n2146_n3206# 3.96721f
C11 B VP 1.22494f
C12 VDD2 VTAIL 13.893201f
C13 B VN 0.775995f
C14 VTAIL w_n2146_n3206# 2.89734f
C15 VDD2 VDD1 0.941936f
C16 VN VP 5.37016f
C17 w_n2146_n3206# VDD1 1.96168f
C18 VTAIL B 2.55494f
C19 VTAIL VP 5.87233f
C20 B VDD1 1.62283f
C21 VDD2 VSUBS 1.417414f
C22 VDD1 VSUBS 1.113311f
C23 VTAIL VSUBS 0.729465f
C24 VN VSUBS 4.83222f
C25 VP VSUBS 1.737032f
C26 B VSUBS 2.880052f
C27 w_n2146_n3206# VSUBS 84.8013f
C28 B.n0 VSUBS 0.006583f
C29 B.n1 VSUBS 0.006583f
C30 B.n2 VSUBS 0.009735f
C31 B.n3 VSUBS 0.00746f
C32 B.n4 VSUBS 0.00746f
C33 B.n5 VSUBS 0.00746f
C34 B.n6 VSUBS 0.00746f
C35 B.n7 VSUBS 0.00746f
C36 B.n8 VSUBS 0.00746f
C37 B.n9 VSUBS 0.00746f
C38 B.n10 VSUBS 0.00746f
C39 B.n11 VSUBS 0.00746f
C40 B.n12 VSUBS 0.00746f
C41 B.n13 VSUBS 0.00746f
C42 B.n14 VSUBS 0.016771f
C43 B.n15 VSUBS 0.00746f
C44 B.n16 VSUBS 0.00746f
C45 B.n17 VSUBS 0.00746f
C46 B.n18 VSUBS 0.00746f
C47 B.n19 VSUBS 0.00746f
C48 B.n20 VSUBS 0.00746f
C49 B.n21 VSUBS 0.00746f
C50 B.n22 VSUBS 0.00746f
C51 B.n23 VSUBS 0.00746f
C52 B.n24 VSUBS 0.00746f
C53 B.n25 VSUBS 0.00746f
C54 B.n26 VSUBS 0.00746f
C55 B.n27 VSUBS 0.00746f
C56 B.n28 VSUBS 0.00746f
C57 B.n29 VSUBS 0.00746f
C58 B.n30 VSUBS 0.00746f
C59 B.n31 VSUBS 0.00746f
C60 B.n32 VSUBS 0.00746f
C61 B.n33 VSUBS 0.00746f
C62 B.t1 VSUBS 0.385622f
C63 B.t2 VSUBS 0.39384f
C64 B.t0 VSUBS 0.319505f
C65 B.n34 VSUBS 0.133226f
C66 B.n35 VSUBS 0.067851f
C67 B.n36 VSUBS 0.017285f
C68 B.n37 VSUBS 0.00746f
C69 B.n38 VSUBS 0.00746f
C70 B.n39 VSUBS 0.00746f
C71 B.n40 VSUBS 0.00746f
C72 B.n41 VSUBS 0.00746f
C73 B.t4 VSUBS 0.385615f
C74 B.t5 VSUBS 0.393834f
C75 B.t3 VSUBS 0.319505f
C76 B.n42 VSUBS 0.133232f
C77 B.n43 VSUBS 0.067858f
C78 B.n44 VSUBS 0.00746f
C79 B.n45 VSUBS 0.00746f
C80 B.n46 VSUBS 0.00746f
C81 B.n47 VSUBS 0.00746f
C82 B.n48 VSUBS 0.00746f
C83 B.n49 VSUBS 0.00746f
C84 B.n50 VSUBS 0.00746f
C85 B.n51 VSUBS 0.00746f
C86 B.n52 VSUBS 0.00746f
C87 B.n53 VSUBS 0.00746f
C88 B.n54 VSUBS 0.00746f
C89 B.n55 VSUBS 0.00746f
C90 B.n56 VSUBS 0.00746f
C91 B.n57 VSUBS 0.00746f
C92 B.n58 VSUBS 0.00746f
C93 B.n59 VSUBS 0.00746f
C94 B.n60 VSUBS 0.00746f
C95 B.n61 VSUBS 0.00746f
C96 B.n62 VSUBS 0.00746f
C97 B.n63 VSUBS 0.016771f
C98 B.n64 VSUBS 0.00746f
C99 B.n65 VSUBS 0.00746f
C100 B.n66 VSUBS 0.00746f
C101 B.n67 VSUBS 0.00746f
C102 B.n68 VSUBS 0.00746f
C103 B.n69 VSUBS 0.00746f
C104 B.n70 VSUBS 0.00746f
C105 B.n71 VSUBS 0.00746f
C106 B.n72 VSUBS 0.00746f
C107 B.n73 VSUBS 0.00746f
C108 B.n74 VSUBS 0.00746f
C109 B.n75 VSUBS 0.00746f
C110 B.n76 VSUBS 0.00746f
C111 B.n77 VSUBS 0.00746f
C112 B.n78 VSUBS 0.00746f
C113 B.n79 VSUBS 0.00746f
C114 B.n80 VSUBS 0.00746f
C115 B.n81 VSUBS 0.00746f
C116 B.n82 VSUBS 0.00746f
C117 B.n83 VSUBS 0.00746f
C118 B.n84 VSUBS 0.00746f
C119 B.n85 VSUBS 0.00746f
C120 B.n86 VSUBS 0.00746f
C121 B.n87 VSUBS 0.00746f
C122 B.n88 VSUBS 0.00746f
C123 B.n89 VSUBS 0.017458f
C124 B.n90 VSUBS 0.00746f
C125 B.n91 VSUBS 0.00746f
C126 B.n92 VSUBS 0.00746f
C127 B.n93 VSUBS 0.00746f
C128 B.n94 VSUBS 0.00746f
C129 B.n95 VSUBS 0.00746f
C130 B.n96 VSUBS 0.00746f
C131 B.n97 VSUBS 0.00746f
C132 B.n98 VSUBS 0.00746f
C133 B.n99 VSUBS 0.00746f
C134 B.n100 VSUBS 0.00746f
C135 B.n101 VSUBS 0.00746f
C136 B.n102 VSUBS 0.00746f
C137 B.n103 VSUBS 0.00746f
C138 B.n104 VSUBS 0.00746f
C139 B.n105 VSUBS 0.00746f
C140 B.n106 VSUBS 0.00746f
C141 B.n107 VSUBS 0.00746f
C142 B.n108 VSUBS 0.007021f
C143 B.n109 VSUBS 0.00746f
C144 B.n110 VSUBS 0.00746f
C145 B.n111 VSUBS 0.00746f
C146 B.n112 VSUBS 0.00746f
C147 B.n113 VSUBS 0.00746f
C148 B.t11 VSUBS 0.385622f
C149 B.t10 VSUBS 0.39384f
C150 B.t9 VSUBS 0.319505f
C151 B.n114 VSUBS 0.133226f
C152 B.n115 VSUBS 0.067851f
C153 B.n116 VSUBS 0.00746f
C154 B.n117 VSUBS 0.00746f
C155 B.n118 VSUBS 0.00746f
C156 B.n119 VSUBS 0.00746f
C157 B.n120 VSUBS 0.00746f
C158 B.n121 VSUBS 0.00746f
C159 B.n122 VSUBS 0.00746f
C160 B.n123 VSUBS 0.00746f
C161 B.n124 VSUBS 0.00746f
C162 B.n125 VSUBS 0.00746f
C163 B.n126 VSUBS 0.00746f
C164 B.n127 VSUBS 0.00746f
C165 B.n128 VSUBS 0.00746f
C166 B.n129 VSUBS 0.00746f
C167 B.n130 VSUBS 0.00746f
C168 B.n131 VSUBS 0.00746f
C169 B.n132 VSUBS 0.00746f
C170 B.n133 VSUBS 0.00746f
C171 B.n134 VSUBS 0.00746f
C172 B.n135 VSUBS 0.016771f
C173 B.n136 VSUBS 0.00746f
C174 B.n137 VSUBS 0.00746f
C175 B.n138 VSUBS 0.00746f
C176 B.n139 VSUBS 0.00746f
C177 B.n140 VSUBS 0.00746f
C178 B.n141 VSUBS 0.00746f
C179 B.n142 VSUBS 0.00746f
C180 B.n143 VSUBS 0.00746f
C181 B.n144 VSUBS 0.00746f
C182 B.n145 VSUBS 0.00746f
C183 B.n146 VSUBS 0.00746f
C184 B.n147 VSUBS 0.00746f
C185 B.n148 VSUBS 0.00746f
C186 B.n149 VSUBS 0.00746f
C187 B.n150 VSUBS 0.00746f
C188 B.n151 VSUBS 0.00746f
C189 B.n152 VSUBS 0.00746f
C190 B.n153 VSUBS 0.00746f
C191 B.n154 VSUBS 0.00746f
C192 B.n155 VSUBS 0.00746f
C193 B.n156 VSUBS 0.00746f
C194 B.n157 VSUBS 0.00746f
C195 B.n158 VSUBS 0.00746f
C196 B.n159 VSUBS 0.00746f
C197 B.n160 VSUBS 0.00746f
C198 B.n161 VSUBS 0.00746f
C199 B.n162 VSUBS 0.00746f
C200 B.n163 VSUBS 0.00746f
C201 B.n164 VSUBS 0.00746f
C202 B.n165 VSUBS 0.00746f
C203 B.n166 VSUBS 0.00746f
C204 B.n167 VSUBS 0.00746f
C205 B.n168 VSUBS 0.00746f
C206 B.n169 VSUBS 0.00746f
C207 B.n170 VSUBS 0.00746f
C208 B.n171 VSUBS 0.00746f
C209 B.n172 VSUBS 0.00746f
C210 B.n173 VSUBS 0.00746f
C211 B.n174 VSUBS 0.00746f
C212 B.n175 VSUBS 0.00746f
C213 B.n176 VSUBS 0.00746f
C214 B.n177 VSUBS 0.00746f
C215 B.n178 VSUBS 0.00746f
C216 B.n179 VSUBS 0.00746f
C217 B.n180 VSUBS 0.00746f
C218 B.n181 VSUBS 0.00746f
C219 B.n182 VSUBS 0.016771f
C220 B.n183 VSUBS 0.017458f
C221 B.n184 VSUBS 0.017458f
C222 B.n185 VSUBS 0.00746f
C223 B.n186 VSUBS 0.00746f
C224 B.n187 VSUBS 0.00746f
C225 B.n188 VSUBS 0.00746f
C226 B.n189 VSUBS 0.00746f
C227 B.n190 VSUBS 0.00746f
C228 B.n191 VSUBS 0.00746f
C229 B.n192 VSUBS 0.00746f
C230 B.n193 VSUBS 0.00746f
C231 B.n194 VSUBS 0.00746f
C232 B.n195 VSUBS 0.00746f
C233 B.n196 VSUBS 0.00746f
C234 B.n197 VSUBS 0.00746f
C235 B.n198 VSUBS 0.00746f
C236 B.n199 VSUBS 0.00746f
C237 B.n200 VSUBS 0.00746f
C238 B.n201 VSUBS 0.00746f
C239 B.n202 VSUBS 0.00746f
C240 B.n203 VSUBS 0.00746f
C241 B.n204 VSUBS 0.00746f
C242 B.n205 VSUBS 0.00746f
C243 B.n206 VSUBS 0.00746f
C244 B.n207 VSUBS 0.00746f
C245 B.n208 VSUBS 0.00746f
C246 B.n209 VSUBS 0.00746f
C247 B.n210 VSUBS 0.00746f
C248 B.n211 VSUBS 0.00746f
C249 B.n212 VSUBS 0.00746f
C250 B.n213 VSUBS 0.00746f
C251 B.n214 VSUBS 0.00746f
C252 B.n215 VSUBS 0.00746f
C253 B.n216 VSUBS 0.00746f
C254 B.n217 VSUBS 0.00746f
C255 B.n218 VSUBS 0.00746f
C256 B.n219 VSUBS 0.00746f
C257 B.n220 VSUBS 0.00746f
C258 B.n221 VSUBS 0.00746f
C259 B.n222 VSUBS 0.00746f
C260 B.n223 VSUBS 0.00746f
C261 B.n224 VSUBS 0.00746f
C262 B.n225 VSUBS 0.00746f
C263 B.n226 VSUBS 0.00746f
C264 B.n227 VSUBS 0.00746f
C265 B.n228 VSUBS 0.00746f
C266 B.n229 VSUBS 0.00746f
C267 B.n230 VSUBS 0.00746f
C268 B.n231 VSUBS 0.00746f
C269 B.n232 VSUBS 0.00746f
C270 B.n233 VSUBS 0.00746f
C271 B.n234 VSUBS 0.00746f
C272 B.n235 VSUBS 0.00746f
C273 B.n236 VSUBS 0.00746f
C274 B.n237 VSUBS 0.00746f
C275 B.n238 VSUBS 0.00746f
C276 B.n239 VSUBS 0.00746f
C277 B.n240 VSUBS 0.00746f
C278 B.n241 VSUBS 0.007021f
C279 B.n242 VSUBS 0.017285f
C280 B.n243 VSUBS 0.004169f
C281 B.n244 VSUBS 0.00746f
C282 B.n245 VSUBS 0.00746f
C283 B.n246 VSUBS 0.00746f
C284 B.n247 VSUBS 0.00746f
C285 B.n248 VSUBS 0.00746f
C286 B.n249 VSUBS 0.00746f
C287 B.n250 VSUBS 0.00746f
C288 B.n251 VSUBS 0.00746f
C289 B.n252 VSUBS 0.00746f
C290 B.n253 VSUBS 0.00746f
C291 B.n254 VSUBS 0.00746f
C292 B.n255 VSUBS 0.00746f
C293 B.t8 VSUBS 0.385615f
C294 B.t7 VSUBS 0.393834f
C295 B.t6 VSUBS 0.319505f
C296 B.n256 VSUBS 0.133232f
C297 B.n257 VSUBS 0.067858f
C298 B.n258 VSUBS 0.017285f
C299 B.n259 VSUBS 0.004169f
C300 B.n260 VSUBS 0.00746f
C301 B.n261 VSUBS 0.00746f
C302 B.n262 VSUBS 0.00746f
C303 B.n263 VSUBS 0.00746f
C304 B.n264 VSUBS 0.00746f
C305 B.n265 VSUBS 0.00746f
C306 B.n266 VSUBS 0.00746f
C307 B.n267 VSUBS 0.00746f
C308 B.n268 VSUBS 0.00746f
C309 B.n269 VSUBS 0.00746f
C310 B.n270 VSUBS 0.00746f
C311 B.n271 VSUBS 0.00746f
C312 B.n272 VSUBS 0.00746f
C313 B.n273 VSUBS 0.00746f
C314 B.n274 VSUBS 0.00746f
C315 B.n275 VSUBS 0.00746f
C316 B.n276 VSUBS 0.00746f
C317 B.n277 VSUBS 0.00746f
C318 B.n278 VSUBS 0.00746f
C319 B.n279 VSUBS 0.00746f
C320 B.n280 VSUBS 0.00746f
C321 B.n281 VSUBS 0.00746f
C322 B.n282 VSUBS 0.00746f
C323 B.n283 VSUBS 0.00746f
C324 B.n284 VSUBS 0.00746f
C325 B.n285 VSUBS 0.00746f
C326 B.n286 VSUBS 0.00746f
C327 B.n287 VSUBS 0.00746f
C328 B.n288 VSUBS 0.00746f
C329 B.n289 VSUBS 0.00746f
C330 B.n290 VSUBS 0.00746f
C331 B.n291 VSUBS 0.00746f
C332 B.n292 VSUBS 0.00746f
C333 B.n293 VSUBS 0.00746f
C334 B.n294 VSUBS 0.00746f
C335 B.n295 VSUBS 0.00746f
C336 B.n296 VSUBS 0.00746f
C337 B.n297 VSUBS 0.00746f
C338 B.n298 VSUBS 0.00746f
C339 B.n299 VSUBS 0.00746f
C340 B.n300 VSUBS 0.00746f
C341 B.n301 VSUBS 0.00746f
C342 B.n302 VSUBS 0.00746f
C343 B.n303 VSUBS 0.00746f
C344 B.n304 VSUBS 0.00746f
C345 B.n305 VSUBS 0.00746f
C346 B.n306 VSUBS 0.00746f
C347 B.n307 VSUBS 0.00746f
C348 B.n308 VSUBS 0.00746f
C349 B.n309 VSUBS 0.00746f
C350 B.n310 VSUBS 0.00746f
C351 B.n311 VSUBS 0.00746f
C352 B.n312 VSUBS 0.00746f
C353 B.n313 VSUBS 0.00746f
C354 B.n314 VSUBS 0.00746f
C355 B.n315 VSUBS 0.00746f
C356 B.n316 VSUBS 0.00746f
C357 B.n317 VSUBS 0.00746f
C358 B.n318 VSUBS 0.01655f
C359 B.n319 VSUBS 0.01768f
C360 B.n320 VSUBS 0.016771f
C361 B.n321 VSUBS 0.00746f
C362 B.n322 VSUBS 0.00746f
C363 B.n323 VSUBS 0.00746f
C364 B.n324 VSUBS 0.00746f
C365 B.n325 VSUBS 0.00746f
C366 B.n326 VSUBS 0.00746f
C367 B.n327 VSUBS 0.00746f
C368 B.n328 VSUBS 0.00746f
C369 B.n329 VSUBS 0.00746f
C370 B.n330 VSUBS 0.00746f
C371 B.n331 VSUBS 0.00746f
C372 B.n332 VSUBS 0.00746f
C373 B.n333 VSUBS 0.00746f
C374 B.n334 VSUBS 0.00746f
C375 B.n335 VSUBS 0.00746f
C376 B.n336 VSUBS 0.00746f
C377 B.n337 VSUBS 0.00746f
C378 B.n338 VSUBS 0.00746f
C379 B.n339 VSUBS 0.00746f
C380 B.n340 VSUBS 0.00746f
C381 B.n341 VSUBS 0.00746f
C382 B.n342 VSUBS 0.00746f
C383 B.n343 VSUBS 0.00746f
C384 B.n344 VSUBS 0.00746f
C385 B.n345 VSUBS 0.00746f
C386 B.n346 VSUBS 0.00746f
C387 B.n347 VSUBS 0.00746f
C388 B.n348 VSUBS 0.00746f
C389 B.n349 VSUBS 0.00746f
C390 B.n350 VSUBS 0.00746f
C391 B.n351 VSUBS 0.00746f
C392 B.n352 VSUBS 0.00746f
C393 B.n353 VSUBS 0.00746f
C394 B.n354 VSUBS 0.00746f
C395 B.n355 VSUBS 0.00746f
C396 B.n356 VSUBS 0.00746f
C397 B.n357 VSUBS 0.00746f
C398 B.n358 VSUBS 0.00746f
C399 B.n359 VSUBS 0.00746f
C400 B.n360 VSUBS 0.00746f
C401 B.n361 VSUBS 0.00746f
C402 B.n362 VSUBS 0.00746f
C403 B.n363 VSUBS 0.00746f
C404 B.n364 VSUBS 0.00746f
C405 B.n365 VSUBS 0.00746f
C406 B.n366 VSUBS 0.00746f
C407 B.n367 VSUBS 0.00746f
C408 B.n368 VSUBS 0.00746f
C409 B.n369 VSUBS 0.00746f
C410 B.n370 VSUBS 0.00746f
C411 B.n371 VSUBS 0.00746f
C412 B.n372 VSUBS 0.00746f
C413 B.n373 VSUBS 0.00746f
C414 B.n374 VSUBS 0.00746f
C415 B.n375 VSUBS 0.00746f
C416 B.n376 VSUBS 0.00746f
C417 B.n377 VSUBS 0.00746f
C418 B.n378 VSUBS 0.00746f
C419 B.n379 VSUBS 0.00746f
C420 B.n380 VSUBS 0.00746f
C421 B.n381 VSUBS 0.00746f
C422 B.n382 VSUBS 0.00746f
C423 B.n383 VSUBS 0.00746f
C424 B.n384 VSUBS 0.00746f
C425 B.n385 VSUBS 0.00746f
C426 B.n386 VSUBS 0.00746f
C427 B.n387 VSUBS 0.00746f
C428 B.n388 VSUBS 0.00746f
C429 B.n389 VSUBS 0.00746f
C430 B.n390 VSUBS 0.00746f
C431 B.n391 VSUBS 0.00746f
C432 B.n392 VSUBS 0.00746f
C433 B.n393 VSUBS 0.00746f
C434 B.n394 VSUBS 0.00746f
C435 B.n395 VSUBS 0.00746f
C436 B.n396 VSUBS 0.016771f
C437 B.n397 VSUBS 0.017458f
C438 B.n398 VSUBS 0.017458f
C439 B.n399 VSUBS 0.00746f
C440 B.n400 VSUBS 0.00746f
C441 B.n401 VSUBS 0.00746f
C442 B.n402 VSUBS 0.00746f
C443 B.n403 VSUBS 0.00746f
C444 B.n404 VSUBS 0.00746f
C445 B.n405 VSUBS 0.00746f
C446 B.n406 VSUBS 0.00746f
C447 B.n407 VSUBS 0.00746f
C448 B.n408 VSUBS 0.00746f
C449 B.n409 VSUBS 0.00746f
C450 B.n410 VSUBS 0.00746f
C451 B.n411 VSUBS 0.00746f
C452 B.n412 VSUBS 0.00746f
C453 B.n413 VSUBS 0.00746f
C454 B.n414 VSUBS 0.00746f
C455 B.n415 VSUBS 0.00746f
C456 B.n416 VSUBS 0.00746f
C457 B.n417 VSUBS 0.00746f
C458 B.n418 VSUBS 0.00746f
C459 B.n419 VSUBS 0.00746f
C460 B.n420 VSUBS 0.00746f
C461 B.n421 VSUBS 0.00746f
C462 B.n422 VSUBS 0.00746f
C463 B.n423 VSUBS 0.00746f
C464 B.n424 VSUBS 0.00746f
C465 B.n425 VSUBS 0.00746f
C466 B.n426 VSUBS 0.00746f
C467 B.n427 VSUBS 0.00746f
C468 B.n428 VSUBS 0.00746f
C469 B.n429 VSUBS 0.00746f
C470 B.n430 VSUBS 0.00746f
C471 B.n431 VSUBS 0.00746f
C472 B.n432 VSUBS 0.00746f
C473 B.n433 VSUBS 0.00746f
C474 B.n434 VSUBS 0.00746f
C475 B.n435 VSUBS 0.00746f
C476 B.n436 VSUBS 0.00746f
C477 B.n437 VSUBS 0.00746f
C478 B.n438 VSUBS 0.00746f
C479 B.n439 VSUBS 0.00746f
C480 B.n440 VSUBS 0.00746f
C481 B.n441 VSUBS 0.00746f
C482 B.n442 VSUBS 0.00746f
C483 B.n443 VSUBS 0.00746f
C484 B.n444 VSUBS 0.00746f
C485 B.n445 VSUBS 0.00746f
C486 B.n446 VSUBS 0.00746f
C487 B.n447 VSUBS 0.00746f
C488 B.n448 VSUBS 0.00746f
C489 B.n449 VSUBS 0.00746f
C490 B.n450 VSUBS 0.00746f
C491 B.n451 VSUBS 0.00746f
C492 B.n452 VSUBS 0.00746f
C493 B.n453 VSUBS 0.00746f
C494 B.n454 VSUBS 0.00746f
C495 B.n455 VSUBS 0.007021f
C496 B.n456 VSUBS 0.017285f
C497 B.n457 VSUBS 0.004169f
C498 B.n458 VSUBS 0.00746f
C499 B.n459 VSUBS 0.00746f
C500 B.n460 VSUBS 0.00746f
C501 B.n461 VSUBS 0.00746f
C502 B.n462 VSUBS 0.00746f
C503 B.n463 VSUBS 0.00746f
C504 B.n464 VSUBS 0.00746f
C505 B.n465 VSUBS 0.00746f
C506 B.n466 VSUBS 0.00746f
C507 B.n467 VSUBS 0.00746f
C508 B.n468 VSUBS 0.00746f
C509 B.n469 VSUBS 0.00746f
C510 B.n470 VSUBS 0.004169f
C511 B.n471 VSUBS 0.00746f
C512 B.n472 VSUBS 0.00746f
C513 B.n473 VSUBS 0.007021f
C514 B.n474 VSUBS 0.00746f
C515 B.n475 VSUBS 0.00746f
C516 B.n476 VSUBS 0.00746f
C517 B.n477 VSUBS 0.00746f
C518 B.n478 VSUBS 0.00746f
C519 B.n479 VSUBS 0.00746f
C520 B.n480 VSUBS 0.00746f
C521 B.n481 VSUBS 0.00746f
C522 B.n482 VSUBS 0.00746f
C523 B.n483 VSUBS 0.00746f
C524 B.n484 VSUBS 0.00746f
C525 B.n485 VSUBS 0.00746f
C526 B.n486 VSUBS 0.00746f
C527 B.n487 VSUBS 0.00746f
C528 B.n488 VSUBS 0.00746f
C529 B.n489 VSUBS 0.00746f
C530 B.n490 VSUBS 0.00746f
C531 B.n491 VSUBS 0.00746f
C532 B.n492 VSUBS 0.00746f
C533 B.n493 VSUBS 0.00746f
C534 B.n494 VSUBS 0.00746f
C535 B.n495 VSUBS 0.00746f
C536 B.n496 VSUBS 0.00746f
C537 B.n497 VSUBS 0.00746f
C538 B.n498 VSUBS 0.00746f
C539 B.n499 VSUBS 0.00746f
C540 B.n500 VSUBS 0.00746f
C541 B.n501 VSUBS 0.00746f
C542 B.n502 VSUBS 0.00746f
C543 B.n503 VSUBS 0.00746f
C544 B.n504 VSUBS 0.00746f
C545 B.n505 VSUBS 0.00746f
C546 B.n506 VSUBS 0.00746f
C547 B.n507 VSUBS 0.00746f
C548 B.n508 VSUBS 0.00746f
C549 B.n509 VSUBS 0.00746f
C550 B.n510 VSUBS 0.00746f
C551 B.n511 VSUBS 0.00746f
C552 B.n512 VSUBS 0.00746f
C553 B.n513 VSUBS 0.00746f
C554 B.n514 VSUBS 0.00746f
C555 B.n515 VSUBS 0.00746f
C556 B.n516 VSUBS 0.00746f
C557 B.n517 VSUBS 0.00746f
C558 B.n518 VSUBS 0.00746f
C559 B.n519 VSUBS 0.00746f
C560 B.n520 VSUBS 0.00746f
C561 B.n521 VSUBS 0.00746f
C562 B.n522 VSUBS 0.00746f
C563 B.n523 VSUBS 0.00746f
C564 B.n524 VSUBS 0.00746f
C565 B.n525 VSUBS 0.00746f
C566 B.n526 VSUBS 0.00746f
C567 B.n527 VSUBS 0.00746f
C568 B.n528 VSUBS 0.00746f
C569 B.n529 VSUBS 0.017458f
C570 B.n530 VSUBS 0.017458f
C571 B.n531 VSUBS 0.016771f
C572 B.n532 VSUBS 0.00746f
C573 B.n533 VSUBS 0.00746f
C574 B.n534 VSUBS 0.00746f
C575 B.n535 VSUBS 0.00746f
C576 B.n536 VSUBS 0.00746f
C577 B.n537 VSUBS 0.00746f
C578 B.n538 VSUBS 0.00746f
C579 B.n539 VSUBS 0.00746f
C580 B.n540 VSUBS 0.00746f
C581 B.n541 VSUBS 0.00746f
C582 B.n542 VSUBS 0.00746f
C583 B.n543 VSUBS 0.00746f
C584 B.n544 VSUBS 0.00746f
C585 B.n545 VSUBS 0.00746f
C586 B.n546 VSUBS 0.00746f
C587 B.n547 VSUBS 0.00746f
C588 B.n548 VSUBS 0.00746f
C589 B.n549 VSUBS 0.00746f
C590 B.n550 VSUBS 0.00746f
C591 B.n551 VSUBS 0.00746f
C592 B.n552 VSUBS 0.00746f
C593 B.n553 VSUBS 0.00746f
C594 B.n554 VSUBS 0.00746f
C595 B.n555 VSUBS 0.00746f
C596 B.n556 VSUBS 0.00746f
C597 B.n557 VSUBS 0.00746f
C598 B.n558 VSUBS 0.00746f
C599 B.n559 VSUBS 0.00746f
C600 B.n560 VSUBS 0.00746f
C601 B.n561 VSUBS 0.00746f
C602 B.n562 VSUBS 0.00746f
C603 B.n563 VSUBS 0.00746f
C604 B.n564 VSUBS 0.00746f
C605 B.n565 VSUBS 0.00746f
C606 B.n566 VSUBS 0.00746f
C607 B.n567 VSUBS 0.009735f
C608 B.n568 VSUBS 0.010371f
C609 B.n569 VSUBS 0.020623f
C610 VDD2.t3 VSUBS 2.45088f
C611 VDD2.t0 VSUBS 0.241102f
C612 VDD2.t1 VSUBS 0.241102f
C613 VDD2.n0 VSUBS 1.86832f
C614 VDD2.n1 VSUBS 1.24252f
C615 VDD2.t7 VSUBS 0.241102f
C616 VDD2.t9 VSUBS 0.241102f
C617 VDD2.n2 VSUBS 1.87296f
C618 VDD2.n3 VSUBS 2.26232f
C619 VDD2.t6 VSUBS 2.44406f
C620 VDD2.n4 VSUBS 2.79525f
C621 VDD2.t4 VSUBS 0.241102f
C622 VDD2.t2 VSUBS 0.241102f
C623 VDD2.n5 VSUBS 1.86833f
C624 VDD2.n6 VSUBS 0.593062f
C625 VDD2.t8 VSUBS 0.241102f
C626 VDD2.t5 VSUBS 0.241102f
C627 VDD2.n7 VSUBS 1.87293f
C628 VN.n0 VSUBS 0.090324f
C629 VN.t9 VSUBS 1.12644f
C630 VN.n1 VSUBS 0.468801f
C631 VN.t6 VSUBS 1.15082f
C632 VN.n2 VSUBS 0.433807f
C633 VN.n3 VSUBS 0.288512f
C634 VN.t8 VSUBS 1.12644f
C635 VN.n4 VSUBS 0.468801f
C636 VN.t2 VSUBS 1.12644f
C637 VN.n5 VSUBS 0.468801f
C638 VN.t0 VSUBS 1.12644f
C639 VN.n6 VSUBS 0.456495f
C640 VN.n7 VSUBS 0.060157f
C641 VN.n8 VSUBS 0.090324f
C642 VN.t1 VSUBS 1.12644f
C643 VN.n9 VSUBS 0.468801f
C644 VN.t7 VSUBS 1.12644f
C645 VN.t4 VSUBS 1.15082f
C646 VN.n10 VSUBS 0.433807f
C647 VN.n11 VSUBS 0.288512f
C648 VN.n12 VSUBS 0.468801f
C649 VN.t5 VSUBS 1.12644f
C650 VN.n13 VSUBS 0.468801f
C651 VN.t3 VSUBS 1.12644f
C652 VN.n14 VSUBS 0.456495f
C653 VN.n15 VSUBS 2.29214f
C654 VDD1.t7 VSUBS 2.23915f
C655 VDD1.t0 VSUBS 0.220272f
C656 VDD1.t2 VSUBS 0.220272f
C657 VDD1.n0 VSUBS 1.70692f
C658 VDD1.n1 VSUBS 1.14057f
C659 VDD1.t1 VSUBS 2.23914f
C660 VDD1.t3 VSUBS 0.220272f
C661 VDD1.t4 VSUBS 0.220272f
C662 VDD1.n2 VSUBS 1.70691f
C663 VDD1.n3 VSUBS 1.13518f
C664 VDD1.t5 VSUBS 0.220272f
C665 VDD1.t8 VSUBS 0.220272f
C666 VDD1.n4 VSUBS 1.71115f
C667 VDD1.n5 VSUBS 2.14218f
C668 VDD1.t6 VSUBS 0.220272f
C669 VDD1.t9 VSUBS 0.220272f
C670 VDD1.n6 VSUBS 1.70691f
C671 VDD1.n7 VSUBS 2.54191f
C672 VTAIL.t2 VSUBS 0.263777f
C673 VTAIL.t0 VSUBS 0.263777f
C674 VTAIL.n0 VSUBS 1.89873f
C675 VTAIL.n1 VSUBS 0.798757f
C676 VTAIL.t14 VSUBS 2.51199f
C677 VTAIL.n2 VSUBS 0.9196f
C678 VTAIL.t10 VSUBS 0.263777f
C679 VTAIL.t16 VSUBS 0.263777f
C680 VTAIL.n3 VSUBS 1.89873f
C681 VTAIL.n4 VSUBS 0.808908f
C682 VTAIL.t12 VSUBS 0.263777f
C683 VTAIL.t19 VSUBS 0.263777f
C684 VTAIL.n5 VSUBS 1.89873f
C685 VTAIL.n6 VSUBS 2.22253f
C686 VTAIL.t9 VSUBS 0.263777f
C687 VTAIL.t5 VSUBS 0.263777f
C688 VTAIL.n7 VSUBS 1.89874f
C689 VTAIL.n8 VSUBS 2.22252f
C690 VTAIL.t4 VSUBS 0.263777f
C691 VTAIL.t3 VSUBS 0.263777f
C692 VTAIL.n9 VSUBS 1.89874f
C693 VTAIL.n10 VSUBS 0.8089f
C694 VTAIL.t1 VSUBS 2.51201f
C695 VTAIL.n11 VSUBS 0.919583f
C696 VTAIL.t18 VSUBS 0.263777f
C697 VTAIL.t13 VSUBS 0.263777f
C698 VTAIL.n12 VSUBS 1.89874f
C699 VTAIL.n13 VSUBS 0.813458f
C700 VTAIL.t11 VSUBS 0.263777f
C701 VTAIL.t17 VSUBS 0.263777f
C702 VTAIL.n14 VSUBS 1.89874f
C703 VTAIL.n15 VSUBS 0.8089f
C704 VTAIL.t15 VSUBS 2.51199f
C705 VTAIL.n16 VSUBS 2.24746f
C706 VTAIL.t8 VSUBS 2.51199f
C707 VTAIL.n17 VSUBS 2.24746f
C708 VTAIL.t6 VSUBS 0.263777f
C709 VTAIL.t7 VSUBS 0.263777f
C710 VTAIL.n18 VSUBS 1.89873f
C711 VTAIL.n19 VSUBS 0.742412f
C712 VP.n0 VSUBS 0.09235f
C713 VP.t6 VSUBS 1.15172f
C714 VP.n1 VSUBS 0.47932f
C715 VP.n2 VSUBS 0.09235f
C716 VP.t0 VSUBS 1.15172f
C717 VP.t3 VSUBS 1.15172f
C718 VP.t7 VSUBS 1.15172f
C719 VP.n3 VSUBS 0.294986f
C720 VP.t9 VSUBS 1.15172f
C721 VP.t2 VSUBS 1.17664f
C722 VP.n4 VSUBS 0.443541f
C723 VP.n5 VSUBS 0.47932f
C724 VP.n6 VSUBS 0.47932f
C725 VP.n7 VSUBS 0.47932f
C726 VP.n8 VSUBS 0.466738f
C727 VP.n9 VSUBS 2.30718f
C728 VP.t8 VSUBS 1.15172f
C729 VP.n10 VSUBS 0.466738f
C730 VP.n11 VSUBS 2.35463f
C731 VP.n12 VSUBS 0.09235f
C732 VP.n13 VSUBS 0.11089f
C733 VP.t5 VSUBS 1.15172f
C734 VP.n14 VSUBS 0.47932f
C735 VP.t4 VSUBS 1.15172f
C736 VP.n15 VSUBS 0.47932f
C737 VP.t1 VSUBS 1.15172f
C738 VP.n16 VSUBS 0.466738f
C739 VP.n17 VSUBS 0.061507f
.ends

