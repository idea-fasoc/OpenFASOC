* NGSPICE file created from diff_pair_sample_0628.ext - technology: sky130A

.subckt diff_pair_sample_0628 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t12 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X1 VDD1.t6 VP.t1 VTAIL.t9 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=3.9
X2 VDD2.t7 VN.t0 VTAIL.t2 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X3 VDD2.t6 VN.t1 VTAIL.t3 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=3.9
X4 VTAIL.t6 VN.t2 VDD2.t5 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X5 VTAIL.t8 VP.t2 VDD1.t5 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X6 VDD2.t4 VN.t3 VTAIL.t5 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X7 B.t11 B.t9 B.t10 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=3.9
X8 B.t8 B.t6 B.t7 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=3.9
X9 VDD2.t3 VN.t4 VTAIL.t1 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=3.9
X10 VTAIL.t4 VN.t5 VDD2.t2 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=3.9
X11 VTAIL.t10 VP.t3 VDD1.t4 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=3.9
X12 B.t5 B.t3 B.t4 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=3.9
X13 VDD1.t3 VP.t4 VTAIL.t11 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X14 B.t2 B.t0 B.t1 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0 ps=0 w=5.99 l=3.9
X15 VTAIL.t13 VP.t5 VDD1.t2 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X16 VDD1.t1 VP.t6 VTAIL.t15 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=2.3361 ps=12.76 w=5.99 l=3.9
X17 VTAIL.t7 VN.t6 VDD2.t1 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=0.98835 pd=6.32 as=0.98835 ps=6.32 w=5.99 l=3.9
X18 VTAIL.t0 VN.t7 VDD2.t0 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=3.9
X19 VTAIL.t14 VP.t7 VDD1.t0 w_n5200_n2166# sky130_fd_pr__pfet_01v8 ad=2.3361 pd=12.76 as=0.98835 ps=6.32 w=5.99 l=3.9
R0 VP.n26 VP.n25 161.3
R1 VP.n27 VP.n22 161.3
R2 VP.n29 VP.n28 161.3
R3 VP.n30 VP.n21 161.3
R4 VP.n32 VP.n31 161.3
R5 VP.n33 VP.n20 161.3
R6 VP.n35 VP.n34 161.3
R7 VP.n36 VP.n19 161.3
R8 VP.n39 VP.n38 161.3
R9 VP.n40 VP.n18 161.3
R10 VP.n42 VP.n41 161.3
R11 VP.n43 VP.n17 161.3
R12 VP.n45 VP.n44 161.3
R13 VP.n46 VP.n16 161.3
R14 VP.n48 VP.n47 161.3
R15 VP.n49 VP.n15 161.3
R16 VP.n51 VP.n50 161.3
R17 VP.n95 VP.n94 161.3
R18 VP.n93 VP.n1 161.3
R19 VP.n92 VP.n91 161.3
R20 VP.n90 VP.n2 161.3
R21 VP.n89 VP.n88 161.3
R22 VP.n87 VP.n3 161.3
R23 VP.n86 VP.n85 161.3
R24 VP.n84 VP.n4 161.3
R25 VP.n83 VP.n82 161.3
R26 VP.n80 VP.n5 161.3
R27 VP.n79 VP.n78 161.3
R28 VP.n77 VP.n6 161.3
R29 VP.n76 VP.n75 161.3
R30 VP.n74 VP.n7 161.3
R31 VP.n73 VP.n72 161.3
R32 VP.n71 VP.n8 161.3
R33 VP.n70 VP.n69 161.3
R34 VP.n67 VP.n9 161.3
R35 VP.n66 VP.n65 161.3
R36 VP.n64 VP.n10 161.3
R37 VP.n63 VP.n62 161.3
R38 VP.n61 VP.n11 161.3
R39 VP.n60 VP.n59 161.3
R40 VP.n58 VP.n12 161.3
R41 VP.n57 VP.n56 161.3
R42 VP.n55 VP.n13 161.3
R43 VP.n54 VP.n53 85.4187
R44 VP.n96 VP.n0 85.4187
R45 VP.n52 VP.n14 85.4187
R46 VP.n23 VP.t3 70.3024
R47 VP.n24 VP.n23 57.2231
R48 VP.n75 VP.n74 56.5193
R49 VP.n31 VP.n30 56.5193
R50 VP.n53 VP.n52 52.5296
R51 VP.n62 VP.n61 42.4359
R52 VP.n88 VP.n87 42.4359
R53 VP.n44 VP.n43 42.4359
R54 VP.n61 VP.n60 38.5509
R55 VP.n88 VP.n2 38.5509
R56 VP.n44 VP.n16 38.5509
R57 VP.n54 VP.t7 37.0156
R58 VP.n68 VP.t4 37.0156
R59 VP.n81 VP.t2 37.0156
R60 VP.n0 VP.t6 37.0156
R61 VP.n14 VP.t1 37.0156
R62 VP.n37 VP.t5 37.0156
R63 VP.n24 VP.t0 37.0156
R64 VP.n56 VP.n55 24.4675
R65 VP.n56 VP.n12 24.4675
R66 VP.n60 VP.n12 24.4675
R67 VP.n62 VP.n10 24.4675
R68 VP.n66 VP.n10 24.4675
R69 VP.n67 VP.n66 24.4675
R70 VP.n69 VP.n8 24.4675
R71 VP.n73 VP.n8 24.4675
R72 VP.n74 VP.n73 24.4675
R73 VP.n75 VP.n6 24.4675
R74 VP.n79 VP.n6 24.4675
R75 VP.n80 VP.n79 24.4675
R76 VP.n82 VP.n4 24.4675
R77 VP.n86 VP.n4 24.4675
R78 VP.n87 VP.n86 24.4675
R79 VP.n92 VP.n2 24.4675
R80 VP.n93 VP.n92 24.4675
R81 VP.n94 VP.n93 24.4675
R82 VP.n48 VP.n16 24.4675
R83 VP.n49 VP.n48 24.4675
R84 VP.n50 VP.n49 24.4675
R85 VP.n31 VP.n20 24.4675
R86 VP.n35 VP.n20 24.4675
R87 VP.n36 VP.n35 24.4675
R88 VP.n38 VP.n18 24.4675
R89 VP.n42 VP.n18 24.4675
R90 VP.n43 VP.n42 24.4675
R91 VP.n25 VP.n22 24.4675
R92 VP.n29 VP.n22 24.4675
R93 VP.n30 VP.n29 24.4675
R94 VP.n69 VP.n68 17.8614
R95 VP.n81 VP.n80 17.8614
R96 VP.n37 VP.n36 17.8614
R97 VP.n25 VP.n24 17.8614
R98 VP.n68 VP.n67 6.60659
R99 VP.n82 VP.n81 6.60659
R100 VP.n38 VP.n37 6.60659
R101 VP.n55 VP.n54 4.64923
R102 VP.n94 VP.n0 4.64923
R103 VP.n50 VP.n14 4.64923
R104 VP.n26 VP.n23 2.42477
R105 VP.n52 VP.n51 0.354971
R106 VP.n53 VP.n13 0.354971
R107 VP.n96 VP.n95 0.354971
R108 VP VP.n96 0.26696
R109 VP.n27 VP.n26 0.189894
R110 VP.n28 VP.n27 0.189894
R111 VP.n28 VP.n21 0.189894
R112 VP.n32 VP.n21 0.189894
R113 VP.n33 VP.n32 0.189894
R114 VP.n34 VP.n33 0.189894
R115 VP.n34 VP.n19 0.189894
R116 VP.n39 VP.n19 0.189894
R117 VP.n40 VP.n39 0.189894
R118 VP.n41 VP.n40 0.189894
R119 VP.n41 VP.n17 0.189894
R120 VP.n45 VP.n17 0.189894
R121 VP.n46 VP.n45 0.189894
R122 VP.n47 VP.n46 0.189894
R123 VP.n47 VP.n15 0.189894
R124 VP.n51 VP.n15 0.189894
R125 VP.n57 VP.n13 0.189894
R126 VP.n58 VP.n57 0.189894
R127 VP.n59 VP.n58 0.189894
R128 VP.n59 VP.n11 0.189894
R129 VP.n63 VP.n11 0.189894
R130 VP.n64 VP.n63 0.189894
R131 VP.n65 VP.n64 0.189894
R132 VP.n65 VP.n9 0.189894
R133 VP.n70 VP.n9 0.189894
R134 VP.n71 VP.n70 0.189894
R135 VP.n72 VP.n71 0.189894
R136 VP.n72 VP.n7 0.189894
R137 VP.n76 VP.n7 0.189894
R138 VP.n77 VP.n76 0.189894
R139 VP.n78 VP.n77 0.189894
R140 VP.n78 VP.n5 0.189894
R141 VP.n83 VP.n5 0.189894
R142 VP.n84 VP.n83 0.189894
R143 VP.n85 VP.n84 0.189894
R144 VP.n85 VP.n3 0.189894
R145 VP.n89 VP.n3 0.189894
R146 VP.n90 VP.n89 0.189894
R147 VP.n91 VP.n90 0.189894
R148 VP.n91 VP.n1 0.189894
R149 VP.n95 VP.n1 0.189894
R150 VTAIL.n258 VTAIL.n232 756.745
R151 VTAIL.n28 VTAIL.n2 756.745
R152 VTAIL.n60 VTAIL.n34 756.745
R153 VTAIL.n94 VTAIL.n68 756.745
R154 VTAIL.n226 VTAIL.n200 756.745
R155 VTAIL.n192 VTAIL.n166 756.745
R156 VTAIL.n160 VTAIL.n134 756.745
R157 VTAIL.n126 VTAIL.n100 756.745
R158 VTAIL.n243 VTAIL.n242 585
R159 VTAIL.n240 VTAIL.n239 585
R160 VTAIL.n249 VTAIL.n248 585
R161 VTAIL.n251 VTAIL.n250 585
R162 VTAIL.n236 VTAIL.n235 585
R163 VTAIL.n257 VTAIL.n256 585
R164 VTAIL.n259 VTAIL.n258 585
R165 VTAIL.n13 VTAIL.n12 585
R166 VTAIL.n10 VTAIL.n9 585
R167 VTAIL.n19 VTAIL.n18 585
R168 VTAIL.n21 VTAIL.n20 585
R169 VTAIL.n6 VTAIL.n5 585
R170 VTAIL.n27 VTAIL.n26 585
R171 VTAIL.n29 VTAIL.n28 585
R172 VTAIL.n45 VTAIL.n44 585
R173 VTAIL.n42 VTAIL.n41 585
R174 VTAIL.n51 VTAIL.n50 585
R175 VTAIL.n53 VTAIL.n52 585
R176 VTAIL.n38 VTAIL.n37 585
R177 VTAIL.n59 VTAIL.n58 585
R178 VTAIL.n61 VTAIL.n60 585
R179 VTAIL.n79 VTAIL.n78 585
R180 VTAIL.n76 VTAIL.n75 585
R181 VTAIL.n85 VTAIL.n84 585
R182 VTAIL.n87 VTAIL.n86 585
R183 VTAIL.n72 VTAIL.n71 585
R184 VTAIL.n93 VTAIL.n92 585
R185 VTAIL.n95 VTAIL.n94 585
R186 VTAIL.n227 VTAIL.n226 585
R187 VTAIL.n225 VTAIL.n224 585
R188 VTAIL.n204 VTAIL.n203 585
R189 VTAIL.n219 VTAIL.n218 585
R190 VTAIL.n217 VTAIL.n216 585
R191 VTAIL.n208 VTAIL.n207 585
R192 VTAIL.n211 VTAIL.n210 585
R193 VTAIL.n193 VTAIL.n192 585
R194 VTAIL.n191 VTAIL.n190 585
R195 VTAIL.n170 VTAIL.n169 585
R196 VTAIL.n185 VTAIL.n184 585
R197 VTAIL.n183 VTAIL.n182 585
R198 VTAIL.n174 VTAIL.n173 585
R199 VTAIL.n177 VTAIL.n176 585
R200 VTAIL.n161 VTAIL.n160 585
R201 VTAIL.n159 VTAIL.n158 585
R202 VTAIL.n138 VTAIL.n137 585
R203 VTAIL.n153 VTAIL.n152 585
R204 VTAIL.n151 VTAIL.n150 585
R205 VTAIL.n142 VTAIL.n141 585
R206 VTAIL.n145 VTAIL.n144 585
R207 VTAIL.n127 VTAIL.n126 585
R208 VTAIL.n125 VTAIL.n124 585
R209 VTAIL.n104 VTAIL.n103 585
R210 VTAIL.n119 VTAIL.n118 585
R211 VTAIL.n117 VTAIL.n116 585
R212 VTAIL.n108 VTAIL.n107 585
R213 VTAIL.n111 VTAIL.n110 585
R214 VTAIL.t3 VTAIL.n241 327.601
R215 VTAIL.t0 VTAIL.n11 327.601
R216 VTAIL.t15 VTAIL.n43 327.601
R217 VTAIL.t14 VTAIL.n77 327.601
R218 VTAIL.t9 VTAIL.n209 327.601
R219 VTAIL.t10 VTAIL.n175 327.601
R220 VTAIL.t1 VTAIL.n143 327.601
R221 VTAIL.t4 VTAIL.n109 327.601
R222 VTAIL.n242 VTAIL.n239 171.744
R223 VTAIL.n249 VTAIL.n239 171.744
R224 VTAIL.n250 VTAIL.n249 171.744
R225 VTAIL.n250 VTAIL.n235 171.744
R226 VTAIL.n257 VTAIL.n235 171.744
R227 VTAIL.n258 VTAIL.n257 171.744
R228 VTAIL.n12 VTAIL.n9 171.744
R229 VTAIL.n19 VTAIL.n9 171.744
R230 VTAIL.n20 VTAIL.n19 171.744
R231 VTAIL.n20 VTAIL.n5 171.744
R232 VTAIL.n27 VTAIL.n5 171.744
R233 VTAIL.n28 VTAIL.n27 171.744
R234 VTAIL.n44 VTAIL.n41 171.744
R235 VTAIL.n51 VTAIL.n41 171.744
R236 VTAIL.n52 VTAIL.n51 171.744
R237 VTAIL.n52 VTAIL.n37 171.744
R238 VTAIL.n59 VTAIL.n37 171.744
R239 VTAIL.n60 VTAIL.n59 171.744
R240 VTAIL.n78 VTAIL.n75 171.744
R241 VTAIL.n85 VTAIL.n75 171.744
R242 VTAIL.n86 VTAIL.n85 171.744
R243 VTAIL.n86 VTAIL.n71 171.744
R244 VTAIL.n93 VTAIL.n71 171.744
R245 VTAIL.n94 VTAIL.n93 171.744
R246 VTAIL.n226 VTAIL.n225 171.744
R247 VTAIL.n225 VTAIL.n203 171.744
R248 VTAIL.n218 VTAIL.n203 171.744
R249 VTAIL.n218 VTAIL.n217 171.744
R250 VTAIL.n217 VTAIL.n207 171.744
R251 VTAIL.n210 VTAIL.n207 171.744
R252 VTAIL.n192 VTAIL.n191 171.744
R253 VTAIL.n191 VTAIL.n169 171.744
R254 VTAIL.n184 VTAIL.n169 171.744
R255 VTAIL.n184 VTAIL.n183 171.744
R256 VTAIL.n183 VTAIL.n173 171.744
R257 VTAIL.n176 VTAIL.n173 171.744
R258 VTAIL.n160 VTAIL.n159 171.744
R259 VTAIL.n159 VTAIL.n137 171.744
R260 VTAIL.n152 VTAIL.n137 171.744
R261 VTAIL.n152 VTAIL.n151 171.744
R262 VTAIL.n151 VTAIL.n141 171.744
R263 VTAIL.n144 VTAIL.n141 171.744
R264 VTAIL.n126 VTAIL.n125 171.744
R265 VTAIL.n125 VTAIL.n103 171.744
R266 VTAIL.n118 VTAIL.n103 171.744
R267 VTAIL.n118 VTAIL.n117 171.744
R268 VTAIL.n117 VTAIL.n107 171.744
R269 VTAIL.n110 VTAIL.n107 171.744
R270 VTAIL.n242 VTAIL.t3 85.8723
R271 VTAIL.n12 VTAIL.t0 85.8723
R272 VTAIL.n44 VTAIL.t15 85.8723
R273 VTAIL.n78 VTAIL.t14 85.8723
R274 VTAIL.n210 VTAIL.t9 85.8723
R275 VTAIL.n176 VTAIL.t10 85.8723
R276 VTAIL.n144 VTAIL.t1 85.8723
R277 VTAIL.n110 VTAIL.t4 85.8723
R278 VTAIL.n199 VTAIL.n198 75.4215
R279 VTAIL.n133 VTAIL.n132 75.4215
R280 VTAIL.n1 VTAIL.n0 75.4214
R281 VTAIL.n67 VTAIL.n66 75.4214
R282 VTAIL.n263 VTAIL.n262 31.9914
R283 VTAIL.n33 VTAIL.n32 31.9914
R284 VTAIL.n65 VTAIL.n64 31.9914
R285 VTAIL.n99 VTAIL.n98 31.9914
R286 VTAIL.n231 VTAIL.n230 31.9914
R287 VTAIL.n197 VTAIL.n196 31.9914
R288 VTAIL.n165 VTAIL.n164 31.9914
R289 VTAIL.n131 VTAIL.n130 31.9914
R290 VTAIL.n263 VTAIL.n231 21.1772
R291 VTAIL.n131 VTAIL.n99 21.1772
R292 VTAIL.n243 VTAIL.n241 16.3865
R293 VTAIL.n13 VTAIL.n11 16.3865
R294 VTAIL.n45 VTAIL.n43 16.3865
R295 VTAIL.n79 VTAIL.n77 16.3865
R296 VTAIL.n211 VTAIL.n209 16.3865
R297 VTAIL.n177 VTAIL.n175 16.3865
R298 VTAIL.n145 VTAIL.n143 16.3865
R299 VTAIL.n111 VTAIL.n109 16.3865
R300 VTAIL.n244 VTAIL.n240 12.8005
R301 VTAIL.n14 VTAIL.n10 12.8005
R302 VTAIL.n46 VTAIL.n42 12.8005
R303 VTAIL.n80 VTAIL.n76 12.8005
R304 VTAIL.n212 VTAIL.n208 12.8005
R305 VTAIL.n178 VTAIL.n174 12.8005
R306 VTAIL.n146 VTAIL.n142 12.8005
R307 VTAIL.n112 VTAIL.n108 12.8005
R308 VTAIL.n248 VTAIL.n247 12.0247
R309 VTAIL.n18 VTAIL.n17 12.0247
R310 VTAIL.n50 VTAIL.n49 12.0247
R311 VTAIL.n84 VTAIL.n83 12.0247
R312 VTAIL.n216 VTAIL.n215 12.0247
R313 VTAIL.n182 VTAIL.n181 12.0247
R314 VTAIL.n150 VTAIL.n149 12.0247
R315 VTAIL.n116 VTAIL.n115 12.0247
R316 VTAIL.n251 VTAIL.n238 11.249
R317 VTAIL.n21 VTAIL.n8 11.249
R318 VTAIL.n53 VTAIL.n40 11.249
R319 VTAIL.n87 VTAIL.n74 11.249
R320 VTAIL.n219 VTAIL.n206 11.249
R321 VTAIL.n185 VTAIL.n172 11.249
R322 VTAIL.n153 VTAIL.n140 11.249
R323 VTAIL.n119 VTAIL.n106 11.249
R324 VTAIL.n252 VTAIL.n236 10.4732
R325 VTAIL.n22 VTAIL.n6 10.4732
R326 VTAIL.n54 VTAIL.n38 10.4732
R327 VTAIL.n88 VTAIL.n72 10.4732
R328 VTAIL.n220 VTAIL.n204 10.4732
R329 VTAIL.n186 VTAIL.n170 10.4732
R330 VTAIL.n154 VTAIL.n138 10.4732
R331 VTAIL.n120 VTAIL.n104 10.4732
R332 VTAIL.n256 VTAIL.n255 9.69747
R333 VTAIL.n26 VTAIL.n25 9.69747
R334 VTAIL.n58 VTAIL.n57 9.69747
R335 VTAIL.n92 VTAIL.n91 9.69747
R336 VTAIL.n224 VTAIL.n223 9.69747
R337 VTAIL.n190 VTAIL.n189 9.69747
R338 VTAIL.n158 VTAIL.n157 9.69747
R339 VTAIL.n124 VTAIL.n123 9.69747
R340 VTAIL.n262 VTAIL.n261 9.45567
R341 VTAIL.n32 VTAIL.n31 9.45567
R342 VTAIL.n64 VTAIL.n63 9.45567
R343 VTAIL.n98 VTAIL.n97 9.45567
R344 VTAIL.n230 VTAIL.n229 9.45567
R345 VTAIL.n196 VTAIL.n195 9.45567
R346 VTAIL.n164 VTAIL.n163 9.45567
R347 VTAIL.n130 VTAIL.n129 9.45567
R348 VTAIL.n261 VTAIL.n260 9.3005
R349 VTAIL.n234 VTAIL.n233 9.3005
R350 VTAIL.n255 VTAIL.n254 9.3005
R351 VTAIL.n253 VTAIL.n252 9.3005
R352 VTAIL.n238 VTAIL.n237 9.3005
R353 VTAIL.n247 VTAIL.n246 9.3005
R354 VTAIL.n245 VTAIL.n244 9.3005
R355 VTAIL.n31 VTAIL.n30 9.3005
R356 VTAIL.n4 VTAIL.n3 9.3005
R357 VTAIL.n25 VTAIL.n24 9.3005
R358 VTAIL.n23 VTAIL.n22 9.3005
R359 VTAIL.n8 VTAIL.n7 9.3005
R360 VTAIL.n17 VTAIL.n16 9.3005
R361 VTAIL.n15 VTAIL.n14 9.3005
R362 VTAIL.n63 VTAIL.n62 9.3005
R363 VTAIL.n36 VTAIL.n35 9.3005
R364 VTAIL.n57 VTAIL.n56 9.3005
R365 VTAIL.n55 VTAIL.n54 9.3005
R366 VTAIL.n40 VTAIL.n39 9.3005
R367 VTAIL.n49 VTAIL.n48 9.3005
R368 VTAIL.n47 VTAIL.n46 9.3005
R369 VTAIL.n97 VTAIL.n96 9.3005
R370 VTAIL.n70 VTAIL.n69 9.3005
R371 VTAIL.n91 VTAIL.n90 9.3005
R372 VTAIL.n89 VTAIL.n88 9.3005
R373 VTAIL.n74 VTAIL.n73 9.3005
R374 VTAIL.n83 VTAIL.n82 9.3005
R375 VTAIL.n81 VTAIL.n80 9.3005
R376 VTAIL.n229 VTAIL.n228 9.3005
R377 VTAIL.n202 VTAIL.n201 9.3005
R378 VTAIL.n223 VTAIL.n222 9.3005
R379 VTAIL.n221 VTAIL.n220 9.3005
R380 VTAIL.n206 VTAIL.n205 9.3005
R381 VTAIL.n215 VTAIL.n214 9.3005
R382 VTAIL.n213 VTAIL.n212 9.3005
R383 VTAIL.n195 VTAIL.n194 9.3005
R384 VTAIL.n168 VTAIL.n167 9.3005
R385 VTAIL.n189 VTAIL.n188 9.3005
R386 VTAIL.n187 VTAIL.n186 9.3005
R387 VTAIL.n172 VTAIL.n171 9.3005
R388 VTAIL.n181 VTAIL.n180 9.3005
R389 VTAIL.n179 VTAIL.n178 9.3005
R390 VTAIL.n163 VTAIL.n162 9.3005
R391 VTAIL.n136 VTAIL.n135 9.3005
R392 VTAIL.n157 VTAIL.n156 9.3005
R393 VTAIL.n155 VTAIL.n154 9.3005
R394 VTAIL.n140 VTAIL.n139 9.3005
R395 VTAIL.n149 VTAIL.n148 9.3005
R396 VTAIL.n147 VTAIL.n146 9.3005
R397 VTAIL.n129 VTAIL.n128 9.3005
R398 VTAIL.n102 VTAIL.n101 9.3005
R399 VTAIL.n123 VTAIL.n122 9.3005
R400 VTAIL.n121 VTAIL.n120 9.3005
R401 VTAIL.n106 VTAIL.n105 9.3005
R402 VTAIL.n115 VTAIL.n114 9.3005
R403 VTAIL.n113 VTAIL.n112 9.3005
R404 VTAIL.n259 VTAIL.n234 8.92171
R405 VTAIL.n29 VTAIL.n4 8.92171
R406 VTAIL.n61 VTAIL.n36 8.92171
R407 VTAIL.n95 VTAIL.n70 8.92171
R408 VTAIL.n227 VTAIL.n202 8.92171
R409 VTAIL.n193 VTAIL.n168 8.92171
R410 VTAIL.n161 VTAIL.n136 8.92171
R411 VTAIL.n127 VTAIL.n102 8.92171
R412 VTAIL.n260 VTAIL.n232 8.14595
R413 VTAIL.n30 VTAIL.n2 8.14595
R414 VTAIL.n62 VTAIL.n34 8.14595
R415 VTAIL.n96 VTAIL.n68 8.14595
R416 VTAIL.n228 VTAIL.n200 8.14595
R417 VTAIL.n194 VTAIL.n166 8.14595
R418 VTAIL.n162 VTAIL.n134 8.14595
R419 VTAIL.n128 VTAIL.n100 8.14595
R420 VTAIL.n262 VTAIL.n232 5.81868
R421 VTAIL.n32 VTAIL.n2 5.81868
R422 VTAIL.n64 VTAIL.n34 5.81868
R423 VTAIL.n98 VTAIL.n68 5.81868
R424 VTAIL.n230 VTAIL.n200 5.81868
R425 VTAIL.n196 VTAIL.n166 5.81868
R426 VTAIL.n164 VTAIL.n134 5.81868
R427 VTAIL.n130 VTAIL.n100 5.81868
R428 VTAIL.n0 VTAIL.t5 5.42704
R429 VTAIL.n0 VTAIL.t7 5.42704
R430 VTAIL.n66 VTAIL.t11 5.42704
R431 VTAIL.n66 VTAIL.t8 5.42704
R432 VTAIL.n198 VTAIL.t12 5.42704
R433 VTAIL.n198 VTAIL.t13 5.42704
R434 VTAIL.n132 VTAIL.t2 5.42704
R435 VTAIL.n132 VTAIL.t6 5.42704
R436 VTAIL.n260 VTAIL.n259 5.04292
R437 VTAIL.n30 VTAIL.n29 5.04292
R438 VTAIL.n62 VTAIL.n61 5.04292
R439 VTAIL.n96 VTAIL.n95 5.04292
R440 VTAIL.n228 VTAIL.n227 5.04292
R441 VTAIL.n194 VTAIL.n193 5.04292
R442 VTAIL.n162 VTAIL.n161 5.04292
R443 VTAIL.n128 VTAIL.n127 5.04292
R444 VTAIL.n256 VTAIL.n234 4.26717
R445 VTAIL.n26 VTAIL.n4 4.26717
R446 VTAIL.n58 VTAIL.n36 4.26717
R447 VTAIL.n92 VTAIL.n70 4.26717
R448 VTAIL.n224 VTAIL.n202 4.26717
R449 VTAIL.n190 VTAIL.n168 4.26717
R450 VTAIL.n158 VTAIL.n136 4.26717
R451 VTAIL.n124 VTAIL.n102 4.26717
R452 VTAIL.n213 VTAIL.n209 3.71286
R453 VTAIL.n179 VTAIL.n175 3.71286
R454 VTAIL.n147 VTAIL.n143 3.71286
R455 VTAIL.n113 VTAIL.n109 3.71286
R456 VTAIL.n245 VTAIL.n241 3.71286
R457 VTAIL.n15 VTAIL.n11 3.71286
R458 VTAIL.n47 VTAIL.n43 3.71286
R459 VTAIL.n81 VTAIL.n77 3.71286
R460 VTAIL.n133 VTAIL.n131 3.64705
R461 VTAIL.n165 VTAIL.n133 3.64705
R462 VTAIL.n199 VTAIL.n197 3.64705
R463 VTAIL.n231 VTAIL.n199 3.64705
R464 VTAIL.n99 VTAIL.n67 3.64705
R465 VTAIL.n67 VTAIL.n65 3.64705
R466 VTAIL.n33 VTAIL.n1 3.64705
R467 VTAIL VTAIL.n263 3.58886
R468 VTAIL.n255 VTAIL.n236 3.49141
R469 VTAIL.n25 VTAIL.n6 3.49141
R470 VTAIL.n57 VTAIL.n38 3.49141
R471 VTAIL.n91 VTAIL.n72 3.49141
R472 VTAIL.n223 VTAIL.n204 3.49141
R473 VTAIL.n189 VTAIL.n170 3.49141
R474 VTAIL.n157 VTAIL.n138 3.49141
R475 VTAIL.n123 VTAIL.n104 3.49141
R476 VTAIL.n252 VTAIL.n251 2.71565
R477 VTAIL.n22 VTAIL.n21 2.71565
R478 VTAIL.n54 VTAIL.n53 2.71565
R479 VTAIL.n88 VTAIL.n87 2.71565
R480 VTAIL.n220 VTAIL.n219 2.71565
R481 VTAIL.n186 VTAIL.n185 2.71565
R482 VTAIL.n154 VTAIL.n153 2.71565
R483 VTAIL.n120 VTAIL.n119 2.71565
R484 VTAIL.n248 VTAIL.n238 1.93989
R485 VTAIL.n18 VTAIL.n8 1.93989
R486 VTAIL.n50 VTAIL.n40 1.93989
R487 VTAIL.n84 VTAIL.n74 1.93989
R488 VTAIL.n216 VTAIL.n206 1.93989
R489 VTAIL.n182 VTAIL.n172 1.93989
R490 VTAIL.n150 VTAIL.n140 1.93989
R491 VTAIL.n116 VTAIL.n106 1.93989
R492 VTAIL.n247 VTAIL.n240 1.16414
R493 VTAIL.n17 VTAIL.n10 1.16414
R494 VTAIL.n49 VTAIL.n42 1.16414
R495 VTAIL.n83 VTAIL.n76 1.16414
R496 VTAIL.n215 VTAIL.n208 1.16414
R497 VTAIL.n181 VTAIL.n174 1.16414
R498 VTAIL.n149 VTAIL.n142 1.16414
R499 VTAIL.n115 VTAIL.n108 1.16414
R500 VTAIL.n197 VTAIL.n165 0.470328
R501 VTAIL.n65 VTAIL.n33 0.470328
R502 VTAIL.n244 VTAIL.n243 0.388379
R503 VTAIL.n14 VTAIL.n13 0.388379
R504 VTAIL.n46 VTAIL.n45 0.388379
R505 VTAIL.n80 VTAIL.n79 0.388379
R506 VTAIL.n212 VTAIL.n211 0.388379
R507 VTAIL.n178 VTAIL.n177 0.388379
R508 VTAIL.n146 VTAIL.n145 0.388379
R509 VTAIL.n112 VTAIL.n111 0.388379
R510 VTAIL.n246 VTAIL.n245 0.155672
R511 VTAIL.n246 VTAIL.n237 0.155672
R512 VTAIL.n253 VTAIL.n237 0.155672
R513 VTAIL.n254 VTAIL.n253 0.155672
R514 VTAIL.n254 VTAIL.n233 0.155672
R515 VTAIL.n261 VTAIL.n233 0.155672
R516 VTAIL.n16 VTAIL.n15 0.155672
R517 VTAIL.n16 VTAIL.n7 0.155672
R518 VTAIL.n23 VTAIL.n7 0.155672
R519 VTAIL.n24 VTAIL.n23 0.155672
R520 VTAIL.n24 VTAIL.n3 0.155672
R521 VTAIL.n31 VTAIL.n3 0.155672
R522 VTAIL.n48 VTAIL.n47 0.155672
R523 VTAIL.n48 VTAIL.n39 0.155672
R524 VTAIL.n55 VTAIL.n39 0.155672
R525 VTAIL.n56 VTAIL.n55 0.155672
R526 VTAIL.n56 VTAIL.n35 0.155672
R527 VTAIL.n63 VTAIL.n35 0.155672
R528 VTAIL.n82 VTAIL.n81 0.155672
R529 VTAIL.n82 VTAIL.n73 0.155672
R530 VTAIL.n89 VTAIL.n73 0.155672
R531 VTAIL.n90 VTAIL.n89 0.155672
R532 VTAIL.n90 VTAIL.n69 0.155672
R533 VTAIL.n97 VTAIL.n69 0.155672
R534 VTAIL.n229 VTAIL.n201 0.155672
R535 VTAIL.n222 VTAIL.n201 0.155672
R536 VTAIL.n222 VTAIL.n221 0.155672
R537 VTAIL.n221 VTAIL.n205 0.155672
R538 VTAIL.n214 VTAIL.n205 0.155672
R539 VTAIL.n214 VTAIL.n213 0.155672
R540 VTAIL.n195 VTAIL.n167 0.155672
R541 VTAIL.n188 VTAIL.n167 0.155672
R542 VTAIL.n188 VTAIL.n187 0.155672
R543 VTAIL.n187 VTAIL.n171 0.155672
R544 VTAIL.n180 VTAIL.n171 0.155672
R545 VTAIL.n180 VTAIL.n179 0.155672
R546 VTAIL.n163 VTAIL.n135 0.155672
R547 VTAIL.n156 VTAIL.n135 0.155672
R548 VTAIL.n156 VTAIL.n155 0.155672
R549 VTAIL.n155 VTAIL.n139 0.155672
R550 VTAIL.n148 VTAIL.n139 0.155672
R551 VTAIL.n148 VTAIL.n147 0.155672
R552 VTAIL.n129 VTAIL.n101 0.155672
R553 VTAIL.n122 VTAIL.n101 0.155672
R554 VTAIL.n122 VTAIL.n121 0.155672
R555 VTAIL.n121 VTAIL.n105 0.155672
R556 VTAIL.n114 VTAIL.n105 0.155672
R557 VTAIL.n114 VTAIL.n113 0.155672
R558 VTAIL VTAIL.n1 0.0586897
R559 VDD1 VDD1.n0 93.9818
R560 VDD1.n3 VDD1.n2 93.8681
R561 VDD1.n3 VDD1.n1 93.8681
R562 VDD1.n5 VDD1.n4 92.1001
R563 VDD1.n5 VDD1.n3 45.8716
R564 VDD1.n4 VDD1.t2 5.42704
R565 VDD1.n4 VDD1.t6 5.42704
R566 VDD1.n0 VDD1.t4 5.42704
R567 VDD1.n0 VDD1.t7 5.42704
R568 VDD1.n2 VDD1.t5 5.42704
R569 VDD1.n2 VDD1.t1 5.42704
R570 VDD1.n1 VDD1.t0 5.42704
R571 VDD1.n1 VDD1.t3 5.42704
R572 VDD1 VDD1.n5 1.76559
R573 VN.n76 VN.n75 161.3
R574 VN.n74 VN.n40 161.3
R575 VN.n73 VN.n72 161.3
R576 VN.n71 VN.n41 161.3
R577 VN.n70 VN.n69 161.3
R578 VN.n68 VN.n42 161.3
R579 VN.n67 VN.n66 161.3
R580 VN.n65 VN.n43 161.3
R581 VN.n64 VN.n63 161.3
R582 VN.n61 VN.n44 161.3
R583 VN.n60 VN.n59 161.3
R584 VN.n58 VN.n45 161.3
R585 VN.n57 VN.n56 161.3
R586 VN.n55 VN.n46 161.3
R587 VN.n54 VN.n53 161.3
R588 VN.n52 VN.n47 161.3
R589 VN.n51 VN.n50 161.3
R590 VN.n37 VN.n36 161.3
R591 VN.n35 VN.n1 161.3
R592 VN.n34 VN.n33 161.3
R593 VN.n32 VN.n2 161.3
R594 VN.n31 VN.n30 161.3
R595 VN.n29 VN.n3 161.3
R596 VN.n28 VN.n27 161.3
R597 VN.n26 VN.n4 161.3
R598 VN.n25 VN.n24 161.3
R599 VN.n22 VN.n5 161.3
R600 VN.n21 VN.n20 161.3
R601 VN.n19 VN.n6 161.3
R602 VN.n18 VN.n17 161.3
R603 VN.n16 VN.n7 161.3
R604 VN.n15 VN.n14 161.3
R605 VN.n13 VN.n8 161.3
R606 VN.n12 VN.n11 161.3
R607 VN.n38 VN.n0 85.4187
R608 VN.n77 VN.n39 85.4187
R609 VN.n9 VN.t7 70.3026
R610 VN.n48 VN.t4 70.3026
R611 VN.n10 VN.n9 57.223
R612 VN.n49 VN.n48 57.223
R613 VN.n17 VN.n16 56.5193
R614 VN.n56 VN.n55 56.5193
R615 VN VN.n77 52.695
R616 VN.n30 VN.n29 42.4359
R617 VN.n69 VN.n68 42.4359
R618 VN.n30 VN.n2 38.5509
R619 VN.n69 VN.n41 38.5509
R620 VN.n10 VN.t3 37.0156
R621 VN.n23 VN.t6 37.0156
R622 VN.n0 VN.t1 37.0156
R623 VN.n49 VN.t2 37.0156
R624 VN.n62 VN.t0 37.0156
R625 VN.n39 VN.t5 37.0156
R626 VN.n11 VN.n8 24.4675
R627 VN.n15 VN.n8 24.4675
R628 VN.n16 VN.n15 24.4675
R629 VN.n17 VN.n6 24.4675
R630 VN.n21 VN.n6 24.4675
R631 VN.n22 VN.n21 24.4675
R632 VN.n24 VN.n4 24.4675
R633 VN.n28 VN.n4 24.4675
R634 VN.n29 VN.n28 24.4675
R635 VN.n34 VN.n2 24.4675
R636 VN.n35 VN.n34 24.4675
R637 VN.n36 VN.n35 24.4675
R638 VN.n55 VN.n54 24.4675
R639 VN.n54 VN.n47 24.4675
R640 VN.n50 VN.n47 24.4675
R641 VN.n68 VN.n67 24.4675
R642 VN.n67 VN.n43 24.4675
R643 VN.n63 VN.n43 24.4675
R644 VN.n61 VN.n60 24.4675
R645 VN.n60 VN.n45 24.4675
R646 VN.n56 VN.n45 24.4675
R647 VN.n75 VN.n74 24.4675
R648 VN.n74 VN.n73 24.4675
R649 VN.n73 VN.n41 24.4675
R650 VN.n11 VN.n10 17.8614
R651 VN.n23 VN.n22 17.8614
R652 VN.n50 VN.n49 17.8614
R653 VN.n62 VN.n61 17.8614
R654 VN.n24 VN.n23 6.60659
R655 VN.n63 VN.n62 6.60659
R656 VN.n36 VN.n0 4.64923
R657 VN.n75 VN.n39 4.64923
R658 VN.n12 VN.n9 2.42478
R659 VN.n51 VN.n48 2.42478
R660 VN.n77 VN.n76 0.354971
R661 VN.n38 VN.n37 0.354971
R662 VN VN.n38 0.26696
R663 VN.n76 VN.n40 0.189894
R664 VN.n72 VN.n40 0.189894
R665 VN.n72 VN.n71 0.189894
R666 VN.n71 VN.n70 0.189894
R667 VN.n70 VN.n42 0.189894
R668 VN.n66 VN.n42 0.189894
R669 VN.n66 VN.n65 0.189894
R670 VN.n65 VN.n64 0.189894
R671 VN.n64 VN.n44 0.189894
R672 VN.n59 VN.n44 0.189894
R673 VN.n59 VN.n58 0.189894
R674 VN.n58 VN.n57 0.189894
R675 VN.n57 VN.n46 0.189894
R676 VN.n53 VN.n46 0.189894
R677 VN.n53 VN.n52 0.189894
R678 VN.n52 VN.n51 0.189894
R679 VN.n13 VN.n12 0.189894
R680 VN.n14 VN.n13 0.189894
R681 VN.n14 VN.n7 0.189894
R682 VN.n18 VN.n7 0.189894
R683 VN.n19 VN.n18 0.189894
R684 VN.n20 VN.n19 0.189894
R685 VN.n20 VN.n5 0.189894
R686 VN.n25 VN.n5 0.189894
R687 VN.n26 VN.n25 0.189894
R688 VN.n27 VN.n26 0.189894
R689 VN.n27 VN.n3 0.189894
R690 VN.n31 VN.n3 0.189894
R691 VN.n32 VN.n31 0.189894
R692 VN.n33 VN.n32 0.189894
R693 VN.n33 VN.n1 0.189894
R694 VN.n37 VN.n1 0.189894
R695 VDD2.n2 VDD2.n1 93.8681
R696 VDD2.n2 VDD2.n0 93.8681
R697 VDD2 VDD2.n5 93.8652
R698 VDD2.n4 VDD2.n3 92.1003
R699 VDD2.n4 VDD2.n2 45.2886
R700 VDD2.n5 VDD2.t5 5.42704
R701 VDD2.n5 VDD2.t3 5.42704
R702 VDD2.n3 VDD2.t2 5.42704
R703 VDD2.n3 VDD2.t7 5.42704
R704 VDD2.n1 VDD2.t1 5.42704
R705 VDD2.n1 VDD2.t6 5.42704
R706 VDD2.n0 VDD2.t0 5.42704
R707 VDD2.n0 VDD2.t4 5.42704
R708 VDD2 VDD2.n4 1.88197
R709 B.n398 B.n397 585
R710 B.n396 B.n141 585
R711 B.n395 B.n394 585
R712 B.n393 B.n142 585
R713 B.n392 B.n391 585
R714 B.n390 B.n143 585
R715 B.n389 B.n388 585
R716 B.n387 B.n144 585
R717 B.n386 B.n385 585
R718 B.n384 B.n145 585
R719 B.n383 B.n382 585
R720 B.n381 B.n146 585
R721 B.n380 B.n379 585
R722 B.n378 B.n147 585
R723 B.n377 B.n376 585
R724 B.n375 B.n148 585
R725 B.n374 B.n373 585
R726 B.n372 B.n149 585
R727 B.n371 B.n370 585
R728 B.n369 B.n150 585
R729 B.n368 B.n367 585
R730 B.n366 B.n151 585
R731 B.n365 B.n364 585
R732 B.n363 B.n152 585
R733 B.n362 B.n361 585
R734 B.n357 B.n153 585
R735 B.n356 B.n355 585
R736 B.n354 B.n154 585
R737 B.n353 B.n352 585
R738 B.n351 B.n155 585
R739 B.n350 B.n349 585
R740 B.n348 B.n156 585
R741 B.n347 B.n346 585
R742 B.n344 B.n157 585
R743 B.n343 B.n342 585
R744 B.n341 B.n160 585
R745 B.n340 B.n339 585
R746 B.n338 B.n161 585
R747 B.n337 B.n336 585
R748 B.n335 B.n162 585
R749 B.n334 B.n333 585
R750 B.n332 B.n163 585
R751 B.n331 B.n330 585
R752 B.n329 B.n164 585
R753 B.n328 B.n327 585
R754 B.n326 B.n165 585
R755 B.n325 B.n324 585
R756 B.n323 B.n166 585
R757 B.n322 B.n321 585
R758 B.n320 B.n167 585
R759 B.n319 B.n318 585
R760 B.n317 B.n168 585
R761 B.n316 B.n315 585
R762 B.n314 B.n169 585
R763 B.n313 B.n312 585
R764 B.n311 B.n170 585
R765 B.n310 B.n309 585
R766 B.n399 B.n140 585
R767 B.n401 B.n400 585
R768 B.n402 B.n139 585
R769 B.n404 B.n403 585
R770 B.n405 B.n138 585
R771 B.n407 B.n406 585
R772 B.n408 B.n137 585
R773 B.n410 B.n409 585
R774 B.n411 B.n136 585
R775 B.n413 B.n412 585
R776 B.n414 B.n135 585
R777 B.n416 B.n415 585
R778 B.n417 B.n134 585
R779 B.n419 B.n418 585
R780 B.n420 B.n133 585
R781 B.n422 B.n421 585
R782 B.n423 B.n132 585
R783 B.n425 B.n424 585
R784 B.n426 B.n131 585
R785 B.n428 B.n427 585
R786 B.n429 B.n130 585
R787 B.n431 B.n430 585
R788 B.n432 B.n129 585
R789 B.n434 B.n433 585
R790 B.n435 B.n128 585
R791 B.n437 B.n436 585
R792 B.n438 B.n127 585
R793 B.n440 B.n439 585
R794 B.n441 B.n126 585
R795 B.n443 B.n442 585
R796 B.n444 B.n125 585
R797 B.n446 B.n445 585
R798 B.n447 B.n124 585
R799 B.n449 B.n448 585
R800 B.n450 B.n123 585
R801 B.n452 B.n451 585
R802 B.n453 B.n122 585
R803 B.n455 B.n454 585
R804 B.n456 B.n121 585
R805 B.n458 B.n457 585
R806 B.n459 B.n120 585
R807 B.n461 B.n460 585
R808 B.n462 B.n119 585
R809 B.n464 B.n463 585
R810 B.n465 B.n118 585
R811 B.n467 B.n466 585
R812 B.n468 B.n117 585
R813 B.n470 B.n469 585
R814 B.n471 B.n116 585
R815 B.n473 B.n472 585
R816 B.n474 B.n115 585
R817 B.n476 B.n475 585
R818 B.n477 B.n114 585
R819 B.n479 B.n478 585
R820 B.n480 B.n113 585
R821 B.n482 B.n481 585
R822 B.n483 B.n112 585
R823 B.n485 B.n484 585
R824 B.n486 B.n111 585
R825 B.n488 B.n487 585
R826 B.n489 B.n110 585
R827 B.n491 B.n490 585
R828 B.n492 B.n109 585
R829 B.n494 B.n493 585
R830 B.n495 B.n108 585
R831 B.n497 B.n496 585
R832 B.n498 B.n107 585
R833 B.n500 B.n499 585
R834 B.n501 B.n106 585
R835 B.n503 B.n502 585
R836 B.n504 B.n105 585
R837 B.n506 B.n505 585
R838 B.n507 B.n104 585
R839 B.n509 B.n508 585
R840 B.n510 B.n103 585
R841 B.n512 B.n511 585
R842 B.n513 B.n102 585
R843 B.n515 B.n514 585
R844 B.n516 B.n101 585
R845 B.n518 B.n517 585
R846 B.n519 B.n100 585
R847 B.n521 B.n520 585
R848 B.n522 B.n99 585
R849 B.n524 B.n523 585
R850 B.n525 B.n98 585
R851 B.n527 B.n526 585
R852 B.n528 B.n97 585
R853 B.n530 B.n529 585
R854 B.n531 B.n96 585
R855 B.n533 B.n532 585
R856 B.n534 B.n95 585
R857 B.n536 B.n535 585
R858 B.n537 B.n94 585
R859 B.n539 B.n538 585
R860 B.n540 B.n93 585
R861 B.n542 B.n541 585
R862 B.n543 B.n92 585
R863 B.n545 B.n544 585
R864 B.n546 B.n91 585
R865 B.n548 B.n547 585
R866 B.n549 B.n90 585
R867 B.n551 B.n550 585
R868 B.n552 B.n89 585
R869 B.n554 B.n553 585
R870 B.n555 B.n88 585
R871 B.n557 B.n556 585
R872 B.n558 B.n87 585
R873 B.n560 B.n559 585
R874 B.n561 B.n86 585
R875 B.n563 B.n562 585
R876 B.n564 B.n85 585
R877 B.n566 B.n565 585
R878 B.n567 B.n84 585
R879 B.n569 B.n568 585
R880 B.n570 B.n83 585
R881 B.n572 B.n571 585
R882 B.n573 B.n82 585
R883 B.n575 B.n574 585
R884 B.n576 B.n81 585
R885 B.n578 B.n577 585
R886 B.n579 B.n80 585
R887 B.n581 B.n580 585
R888 B.n582 B.n79 585
R889 B.n584 B.n583 585
R890 B.n585 B.n78 585
R891 B.n587 B.n586 585
R892 B.n588 B.n77 585
R893 B.n590 B.n589 585
R894 B.n591 B.n76 585
R895 B.n593 B.n592 585
R896 B.n594 B.n75 585
R897 B.n596 B.n595 585
R898 B.n597 B.n74 585
R899 B.n599 B.n598 585
R900 B.n600 B.n73 585
R901 B.n602 B.n601 585
R902 B.n603 B.n72 585
R903 B.n605 B.n604 585
R904 B.n606 B.n71 585
R905 B.n608 B.n607 585
R906 B.n609 B.n70 585
R907 B.n611 B.n610 585
R908 B.n698 B.n37 585
R909 B.n697 B.n696 585
R910 B.n695 B.n38 585
R911 B.n694 B.n693 585
R912 B.n692 B.n39 585
R913 B.n691 B.n690 585
R914 B.n689 B.n40 585
R915 B.n688 B.n687 585
R916 B.n686 B.n41 585
R917 B.n685 B.n684 585
R918 B.n683 B.n42 585
R919 B.n682 B.n681 585
R920 B.n680 B.n43 585
R921 B.n679 B.n678 585
R922 B.n677 B.n44 585
R923 B.n676 B.n675 585
R924 B.n674 B.n45 585
R925 B.n673 B.n672 585
R926 B.n671 B.n46 585
R927 B.n670 B.n669 585
R928 B.n668 B.n47 585
R929 B.n667 B.n666 585
R930 B.n665 B.n48 585
R931 B.n664 B.n663 585
R932 B.n661 B.n49 585
R933 B.n660 B.n659 585
R934 B.n658 B.n52 585
R935 B.n657 B.n656 585
R936 B.n655 B.n53 585
R937 B.n654 B.n653 585
R938 B.n652 B.n54 585
R939 B.n651 B.n650 585
R940 B.n649 B.n55 585
R941 B.n647 B.n646 585
R942 B.n645 B.n58 585
R943 B.n644 B.n643 585
R944 B.n642 B.n59 585
R945 B.n641 B.n640 585
R946 B.n639 B.n60 585
R947 B.n638 B.n637 585
R948 B.n636 B.n61 585
R949 B.n635 B.n634 585
R950 B.n633 B.n62 585
R951 B.n632 B.n631 585
R952 B.n630 B.n63 585
R953 B.n629 B.n628 585
R954 B.n627 B.n64 585
R955 B.n626 B.n625 585
R956 B.n624 B.n65 585
R957 B.n623 B.n622 585
R958 B.n621 B.n66 585
R959 B.n620 B.n619 585
R960 B.n618 B.n67 585
R961 B.n617 B.n616 585
R962 B.n615 B.n68 585
R963 B.n614 B.n613 585
R964 B.n612 B.n69 585
R965 B.n700 B.n699 585
R966 B.n701 B.n36 585
R967 B.n703 B.n702 585
R968 B.n704 B.n35 585
R969 B.n706 B.n705 585
R970 B.n707 B.n34 585
R971 B.n709 B.n708 585
R972 B.n710 B.n33 585
R973 B.n712 B.n711 585
R974 B.n713 B.n32 585
R975 B.n715 B.n714 585
R976 B.n716 B.n31 585
R977 B.n718 B.n717 585
R978 B.n719 B.n30 585
R979 B.n721 B.n720 585
R980 B.n722 B.n29 585
R981 B.n724 B.n723 585
R982 B.n725 B.n28 585
R983 B.n727 B.n726 585
R984 B.n728 B.n27 585
R985 B.n730 B.n729 585
R986 B.n731 B.n26 585
R987 B.n733 B.n732 585
R988 B.n734 B.n25 585
R989 B.n736 B.n735 585
R990 B.n737 B.n24 585
R991 B.n739 B.n738 585
R992 B.n740 B.n23 585
R993 B.n742 B.n741 585
R994 B.n743 B.n22 585
R995 B.n745 B.n744 585
R996 B.n746 B.n21 585
R997 B.n748 B.n747 585
R998 B.n749 B.n20 585
R999 B.n751 B.n750 585
R1000 B.n752 B.n19 585
R1001 B.n754 B.n753 585
R1002 B.n755 B.n18 585
R1003 B.n757 B.n756 585
R1004 B.n758 B.n17 585
R1005 B.n760 B.n759 585
R1006 B.n761 B.n16 585
R1007 B.n763 B.n762 585
R1008 B.n764 B.n15 585
R1009 B.n766 B.n765 585
R1010 B.n767 B.n14 585
R1011 B.n769 B.n768 585
R1012 B.n770 B.n13 585
R1013 B.n772 B.n771 585
R1014 B.n773 B.n12 585
R1015 B.n775 B.n774 585
R1016 B.n776 B.n11 585
R1017 B.n778 B.n777 585
R1018 B.n779 B.n10 585
R1019 B.n781 B.n780 585
R1020 B.n782 B.n9 585
R1021 B.n784 B.n783 585
R1022 B.n785 B.n8 585
R1023 B.n787 B.n786 585
R1024 B.n788 B.n7 585
R1025 B.n790 B.n789 585
R1026 B.n791 B.n6 585
R1027 B.n793 B.n792 585
R1028 B.n794 B.n5 585
R1029 B.n796 B.n795 585
R1030 B.n797 B.n4 585
R1031 B.n799 B.n798 585
R1032 B.n800 B.n3 585
R1033 B.n802 B.n801 585
R1034 B.n803 B.n0 585
R1035 B.n2 B.n1 585
R1036 B.n206 B.n205 585
R1037 B.n208 B.n207 585
R1038 B.n209 B.n204 585
R1039 B.n211 B.n210 585
R1040 B.n212 B.n203 585
R1041 B.n214 B.n213 585
R1042 B.n215 B.n202 585
R1043 B.n217 B.n216 585
R1044 B.n218 B.n201 585
R1045 B.n220 B.n219 585
R1046 B.n221 B.n200 585
R1047 B.n223 B.n222 585
R1048 B.n224 B.n199 585
R1049 B.n226 B.n225 585
R1050 B.n227 B.n198 585
R1051 B.n229 B.n228 585
R1052 B.n230 B.n197 585
R1053 B.n232 B.n231 585
R1054 B.n233 B.n196 585
R1055 B.n235 B.n234 585
R1056 B.n236 B.n195 585
R1057 B.n238 B.n237 585
R1058 B.n239 B.n194 585
R1059 B.n241 B.n240 585
R1060 B.n242 B.n193 585
R1061 B.n244 B.n243 585
R1062 B.n245 B.n192 585
R1063 B.n247 B.n246 585
R1064 B.n248 B.n191 585
R1065 B.n250 B.n249 585
R1066 B.n251 B.n190 585
R1067 B.n253 B.n252 585
R1068 B.n254 B.n189 585
R1069 B.n256 B.n255 585
R1070 B.n257 B.n188 585
R1071 B.n259 B.n258 585
R1072 B.n260 B.n187 585
R1073 B.n262 B.n261 585
R1074 B.n263 B.n186 585
R1075 B.n265 B.n264 585
R1076 B.n266 B.n185 585
R1077 B.n268 B.n267 585
R1078 B.n269 B.n184 585
R1079 B.n271 B.n270 585
R1080 B.n272 B.n183 585
R1081 B.n274 B.n273 585
R1082 B.n275 B.n182 585
R1083 B.n277 B.n276 585
R1084 B.n278 B.n181 585
R1085 B.n280 B.n279 585
R1086 B.n281 B.n180 585
R1087 B.n283 B.n282 585
R1088 B.n284 B.n179 585
R1089 B.n286 B.n285 585
R1090 B.n287 B.n178 585
R1091 B.n289 B.n288 585
R1092 B.n290 B.n177 585
R1093 B.n292 B.n291 585
R1094 B.n293 B.n176 585
R1095 B.n295 B.n294 585
R1096 B.n296 B.n175 585
R1097 B.n298 B.n297 585
R1098 B.n299 B.n174 585
R1099 B.n301 B.n300 585
R1100 B.n302 B.n173 585
R1101 B.n304 B.n303 585
R1102 B.n305 B.n172 585
R1103 B.n307 B.n306 585
R1104 B.n308 B.n171 585
R1105 B.n310 B.n171 506.916
R1106 B.n399 B.n398 506.916
R1107 B.n610 B.n69 506.916
R1108 B.n700 B.n37 506.916
R1109 B.n358 B.t4 350.036
R1110 B.n56 B.t8 350.036
R1111 B.n158 B.t10 350.036
R1112 B.n50 B.t2 350.036
R1113 B.n359 B.t5 268
R1114 B.n57 B.t7 268
R1115 B.n159 B.t11 267.998
R1116 B.n51 B.t1 267.998
R1117 B.n805 B.n804 256.663
R1118 B.n158 B.t9 246.435
R1119 B.n358 B.t3 246.435
R1120 B.n56 B.t6 246.435
R1121 B.n50 B.t0 246.435
R1122 B.n804 B.n803 235.042
R1123 B.n804 B.n2 235.042
R1124 B.n311 B.n310 163.367
R1125 B.n312 B.n311 163.367
R1126 B.n312 B.n169 163.367
R1127 B.n316 B.n169 163.367
R1128 B.n317 B.n316 163.367
R1129 B.n318 B.n317 163.367
R1130 B.n318 B.n167 163.367
R1131 B.n322 B.n167 163.367
R1132 B.n323 B.n322 163.367
R1133 B.n324 B.n323 163.367
R1134 B.n324 B.n165 163.367
R1135 B.n328 B.n165 163.367
R1136 B.n329 B.n328 163.367
R1137 B.n330 B.n329 163.367
R1138 B.n330 B.n163 163.367
R1139 B.n334 B.n163 163.367
R1140 B.n335 B.n334 163.367
R1141 B.n336 B.n335 163.367
R1142 B.n336 B.n161 163.367
R1143 B.n340 B.n161 163.367
R1144 B.n341 B.n340 163.367
R1145 B.n342 B.n341 163.367
R1146 B.n342 B.n157 163.367
R1147 B.n347 B.n157 163.367
R1148 B.n348 B.n347 163.367
R1149 B.n349 B.n348 163.367
R1150 B.n349 B.n155 163.367
R1151 B.n353 B.n155 163.367
R1152 B.n354 B.n353 163.367
R1153 B.n355 B.n354 163.367
R1154 B.n355 B.n153 163.367
R1155 B.n362 B.n153 163.367
R1156 B.n363 B.n362 163.367
R1157 B.n364 B.n363 163.367
R1158 B.n364 B.n151 163.367
R1159 B.n368 B.n151 163.367
R1160 B.n369 B.n368 163.367
R1161 B.n370 B.n369 163.367
R1162 B.n370 B.n149 163.367
R1163 B.n374 B.n149 163.367
R1164 B.n375 B.n374 163.367
R1165 B.n376 B.n375 163.367
R1166 B.n376 B.n147 163.367
R1167 B.n380 B.n147 163.367
R1168 B.n381 B.n380 163.367
R1169 B.n382 B.n381 163.367
R1170 B.n382 B.n145 163.367
R1171 B.n386 B.n145 163.367
R1172 B.n387 B.n386 163.367
R1173 B.n388 B.n387 163.367
R1174 B.n388 B.n143 163.367
R1175 B.n392 B.n143 163.367
R1176 B.n393 B.n392 163.367
R1177 B.n394 B.n393 163.367
R1178 B.n394 B.n141 163.367
R1179 B.n398 B.n141 163.367
R1180 B.n610 B.n609 163.367
R1181 B.n609 B.n608 163.367
R1182 B.n608 B.n71 163.367
R1183 B.n604 B.n71 163.367
R1184 B.n604 B.n603 163.367
R1185 B.n603 B.n602 163.367
R1186 B.n602 B.n73 163.367
R1187 B.n598 B.n73 163.367
R1188 B.n598 B.n597 163.367
R1189 B.n597 B.n596 163.367
R1190 B.n596 B.n75 163.367
R1191 B.n592 B.n75 163.367
R1192 B.n592 B.n591 163.367
R1193 B.n591 B.n590 163.367
R1194 B.n590 B.n77 163.367
R1195 B.n586 B.n77 163.367
R1196 B.n586 B.n585 163.367
R1197 B.n585 B.n584 163.367
R1198 B.n584 B.n79 163.367
R1199 B.n580 B.n79 163.367
R1200 B.n580 B.n579 163.367
R1201 B.n579 B.n578 163.367
R1202 B.n578 B.n81 163.367
R1203 B.n574 B.n81 163.367
R1204 B.n574 B.n573 163.367
R1205 B.n573 B.n572 163.367
R1206 B.n572 B.n83 163.367
R1207 B.n568 B.n83 163.367
R1208 B.n568 B.n567 163.367
R1209 B.n567 B.n566 163.367
R1210 B.n566 B.n85 163.367
R1211 B.n562 B.n85 163.367
R1212 B.n562 B.n561 163.367
R1213 B.n561 B.n560 163.367
R1214 B.n560 B.n87 163.367
R1215 B.n556 B.n87 163.367
R1216 B.n556 B.n555 163.367
R1217 B.n555 B.n554 163.367
R1218 B.n554 B.n89 163.367
R1219 B.n550 B.n89 163.367
R1220 B.n550 B.n549 163.367
R1221 B.n549 B.n548 163.367
R1222 B.n548 B.n91 163.367
R1223 B.n544 B.n91 163.367
R1224 B.n544 B.n543 163.367
R1225 B.n543 B.n542 163.367
R1226 B.n542 B.n93 163.367
R1227 B.n538 B.n93 163.367
R1228 B.n538 B.n537 163.367
R1229 B.n537 B.n536 163.367
R1230 B.n536 B.n95 163.367
R1231 B.n532 B.n95 163.367
R1232 B.n532 B.n531 163.367
R1233 B.n531 B.n530 163.367
R1234 B.n530 B.n97 163.367
R1235 B.n526 B.n97 163.367
R1236 B.n526 B.n525 163.367
R1237 B.n525 B.n524 163.367
R1238 B.n524 B.n99 163.367
R1239 B.n520 B.n99 163.367
R1240 B.n520 B.n519 163.367
R1241 B.n519 B.n518 163.367
R1242 B.n518 B.n101 163.367
R1243 B.n514 B.n101 163.367
R1244 B.n514 B.n513 163.367
R1245 B.n513 B.n512 163.367
R1246 B.n512 B.n103 163.367
R1247 B.n508 B.n103 163.367
R1248 B.n508 B.n507 163.367
R1249 B.n507 B.n506 163.367
R1250 B.n506 B.n105 163.367
R1251 B.n502 B.n105 163.367
R1252 B.n502 B.n501 163.367
R1253 B.n501 B.n500 163.367
R1254 B.n500 B.n107 163.367
R1255 B.n496 B.n107 163.367
R1256 B.n496 B.n495 163.367
R1257 B.n495 B.n494 163.367
R1258 B.n494 B.n109 163.367
R1259 B.n490 B.n109 163.367
R1260 B.n490 B.n489 163.367
R1261 B.n489 B.n488 163.367
R1262 B.n488 B.n111 163.367
R1263 B.n484 B.n111 163.367
R1264 B.n484 B.n483 163.367
R1265 B.n483 B.n482 163.367
R1266 B.n482 B.n113 163.367
R1267 B.n478 B.n113 163.367
R1268 B.n478 B.n477 163.367
R1269 B.n477 B.n476 163.367
R1270 B.n476 B.n115 163.367
R1271 B.n472 B.n115 163.367
R1272 B.n472 B.n471 163.367
R1273 B.n471 B.n470 163.367
R1274 B.n470 B.n117 163.367
R1275 B.n466 B.n117 163.367
R1276 B.n466 B.n465 163.367
R1277 B.n465 B.n464 163.367
R1278 B.n464 B.n119 163.367
R1279 B.n460 B.n119 163.367
R1280 B.n460 B.n459 163.367
R1281 B.n459 B.n458 163.367
R1282 B.n458 B.n121 163.367
R1283 B.n454 B.n121 163.367
R1284 B.n454 B.n453 163.367
R1285 B.n453 B.n452 163.367
R1286 B.n452 B.n123 163.367
R1287 B.n448 B.n123 163.367
R1288 B.n448 B.n447 163.367
R1289 B.n447 B.n446 163.367
R1290 B.n446 B.n125 163.367
R1291 B.n442 B.n125 163.367
R1292 B.n442 B.n441 163.367
R1293 B.n441 B.n440 163.367
R1294 B.n440 B.n127 163.367
R1295 B.n436 B.n127 163.367
R1296 B.n436 B.n435 163.367
R1297 B.n435 B.n434 163.367
R1298 B.n434 B.n129 163.367
R1299 B.n430 B.n129 163.367
R1300 B.n430 B.n429 163.367
R1301 B.n429 B.n428 163.367
R1302 B.n428 B.n131 163.367
R1303 B.n424 B.n131 163.367
R1304 B.n424 B.n423 163.367
R1305 B.n423 B.n422 163.367
R1306 B.n422 B.n133 163.367
R1307 B.n418 B.n133 163.367
R1308 B.n418 B.n417 163.367
R1309 B.n417 B.n416 163.367
R1310 B.n416 B.n135 163.367
R1311 B.n412 B.n135 163.367
R1312 B.n412 B.n411 163.367
R1313 B.n411 B.n410 163.367
R1314 B.n410 B.n137 163.367
R1315 B.n406 B.n137 163.367
R1316 B.n406 B.n405 163.367
R1317 B.n405 B.n404 163.367
R1318 B.n404 B.n139 163.367
R1319 B.n400 B.n139 163.367
R1320 B.n400 B.n399 163.367
R1321 B.n696 B.n37 163.367
R1322 B.n696 B.n695 163.367
R1323 B.n695 B.n694 163.367
R1324 B.n694 B.n39 163.367
R1325 B.n690 B.n39 163.367
R1326 B.n690 B.n689 163.367
R1327 B.n689 B.n688 163.367
R1328 B.n688 B.n41 163.367
R1329 B.n684 B.n41 163.367
R1330 B.n684 B.n683 163.367
R1331 B.n683 B.n682 163.367
R1332 B.n682 B.n43 163.367
R1333 B.n678 B.n43 163.367
R1334 B.n678 B.n677 163.367
R1335 B.n677 B.n676 163.367
R1336 B.n676 B.n45 163.367
R1337 B.n672 B.n45 163.367
R1338 B.n672 B.n671 163.367
R1339 B.n671 B.n670 163.367
R1340 B.n670 B.n47 163.367
R1341 B.n666 B.n47 163.367
R1342 B.n666 B.n665 163.367
R1343 B.n665 B.n664 163.367
R1344 B.n664 B.n49 163.367
R1345 B.n659 B.n49 163.367
R1346 B.n659 B.n658 163.367
R1347 B.n658 B.n657 163.367
R1348 B.n657 B.n53 163.367
R1349 B.n653 B.n53 163.367
R1350 B.n653 B.n652 163.367
R1351 B.n652 B.n651 163.367
R1352 B.n651 B.n55 163.367
R1353 B.n646 B.n55 163.367
R1354 B.n646 B.n645 163.367
R1355 B.n645 B.n644 163.367
R1356 B.n644 B.n59 163.367
R1357 B.n640 B.n59 163.367
R1358 B.n640 B.n639 163.367
R1359 B.n639 B.n638 163.367
R1360 B.n638 B.n61 163.367
R1361 B.n634 B.n61 163.367
R1362 B.n634 B.n633 163.367
R1363 B.n633 B.n632 163.367
R1364 B.n632 B.n63 163.367
R1365 B.n628 B.n63 163.367
R1366 B.n628 B.n627 163.367
R1367 B.n627 B.n626 163.367
R1368 B.n626 B.n65 163.367
R1369 B.n622 B.n65 163.367
R1370 B.n622 B.n621 163.367
R1371 B.n621 B.n620 163.367
R1372 B.n620 B.n67 163.367
R1373 B.n616 B.n67 163.367
R1374 B.n616 B.n615 163.367
R1375 B.n615 B.n614 163.367
R1376 B.n614 B.n69 163.367
R1377 B.n701 B.n700 163.367
R1378 B.n702 B.n701 163.367
R1379 B.n702 B.n35 163.367
R1380 B.n706 B.n35 163.367
R1381 B.n707 B.n706 163.367
R1382 B.n708 B.n707 163.367
R1383 B.n708 B.n33 163.367
R1384 B.n712 B.n33 163.367
R1385 B.n713 B.n712 163.367
R1386 B.n714 B.n713 163.367
R1387 B.n714 B.n31 163.367
R1388 B.n718 B.n31 163.367
R1389 B.n719 B.n718 163.367
R1390 B.n720 B.n719 163.367
R1391 B.n720 B.n29 163.367
R1392 B.n724 B.n29 163.367
R1393 B.n725 B.n724 163.367
R1394 B.n726 B.n725 163.367
R1395 B.n726 B.n27 163.367
R1396 B.n730 B.n27 163.367
R1397 B.n731 B.n730 163.367
R1398 B.n732 B.n731 163.367
R1399 B.n732 B.n25 163.367
R1400 B.n736 B.n25 163.367
R1401 B.n737 B.n736 163.367
R1402 B.n738 B.n737 163.367
R1403 B.n738 B.n23 163.367
R1404 B.n742 B.n23 163.367
R1405 B.n743 B.n742 163.367
R1406 B.n744 B.n743 163.367
R1407 B.n744 B.n21 163.367
R1408 B.n748 B.n21 163.367
R1409 B.n749 B.n748 163.367
R1410 B.n750 B.n749 163.367
R1411 B.n750 B.n19 163.367
R1412 B.n754 B.n19 163.367
R1413 B.n755 B.n754 163.367
R1414 B.n756 B.n755 163.367
R1415 B.n756 B.n17 163.367
R1416 B.n760 B.n17 163.367
R1417 B.n761 B.n760 163.367
R1418 B.n762 B.n761 163.367
R1419 B.n762 B.n15 163.367
R1420 B.n766 B.n15 163.367
R1421 B.n767 B.n766 163.367
R1422 B.n768 B.n767 163.367
R1423 B.n768 B.n13 163.367
R1424 B.n772 B.n13 163.367
R1425 B.n773 B.n772 163.367
R1426 B.n774 B.n773 163.367
R1427 B.n774 B.n11 163.367
R1428 B.n778 B.n11 163.367
R1429 B.n779 B.n778 163.367
R1430 B.n780 B.n779 163.367
R1431 B.n780 B.n9 163.367
R1432 B.n784 B.n9 163.367
R1433 B.n785 B.n784 163.367
R1434 B.n786 B.n785 163.367
R1435 B.n786 B.n7 163.367
R1436 B.n790 B.n7 163.367
R1437 B.n791 B.n790 163.367
R1438 B.n792 B.n791 163.367
R1439 B.n792 B.n5 163.367
R1440 B.n796 B.n5 163.367
R1441 B.n797 B.n796 163.367
R1442 B.n798 B.n797 163.367
R1443 B.n798 B.n3 163.367
R1444 B.n802 B.n3 163.367
R1445 B.n803 B.n802 163.367
R1446 B.n205 B.n2 163.367
R1447 B.n208 B.n205 163.367
R1448 B.n209 B.n208 163.367
R1449 B.n210 B.n209 163.367
R1450 B.n210 B.n203 163.367
R1451 B.n214 B.n203 163.367
R1452 B.n215 B.n214 163.367
R1453 B.n216 B.n215 163.367
R1454 B.n216 B.n201 163.367
R1455 B.n220 B.n201 163.367
R1456 B.n221 B.n220 163.367
R1457 B.n222 B.n221 163.367
R1458 B.n222 B.n199 163.367
R1459 B.n226 B.n199 163.367
R1460 B.n227 B.n226 163.367
R1461 B.n228 B.n227 163.367
R1462 B.n228 B.n197 163.367
R1463 B.n232 B.n197 163.367
R1464 B.n233 B.n232 163.367
R1465 B.n234 B.n233 163.367
R1466 B.n234 B.n195 163.367
R1467 B.n238 B.n195 163.367
R1468 B.n239 B.n238 163.367
R1469 B.n240 B.n239 163.367
R1470 B.n240 B.n193 163.367
R1471 B.n244 B.n193 163.367
R1472 B.n245 B.n244 163.367
R1473 B.n246 B.n245 163.367
R1474 B.n246 B.n191 163.367
R1475 B.n250 B.n191 163.367
R1476 B.n251 B.n250 163.367
R1477 B.n252 B.n251 163.367
R1478 B.n252 B.n189 163.367
R1479 B.n256 B.n189 163.367
R1480 B.n257 B.n256 163.367
R1481 B.n258 B.n257 163.367
R1482 B.n258 B.n187 163.367
R1483 B.n262 B.n187 163.367
R1484 B.n263 B.n262 163.367
R1485 B.n264 B.n263 163.367
R1486 B.n264 B.n185 163.367
R1487 B.n268 B.n185 163.367
R1488 B.n269 B.n268 163.367
R1489 B.n270 B.n269 163.367
R1490 B.n270 B.n183 163.367
R1491 B.n274 B.n183 163.367
R1492 B.n275 B.n274 163.367
R1493 B.n276 B.n275 163.367
R1494 B.n276 B.n181 163.367
R1495 B.n280 B.n181 163.367
R1496 B.n281 B.n280 163.367
R1497 B.n282 B.n281 163.367
R1498 B.n282 B.n179 163.367
R1499 B.n286 B.n179 163.367
R1500 B.n287 B.n286 163.367
R1501 B.n288 B.n287 163.367
R1502 B.n288 B.n177 163.367
R1503 B.n292 B.n177 163.367
R1504 B.n293 B.n292 163.367
R1505 B.n294 B.n293 163.367
R1506 B.n294 B.n175 163.367
R1507 B.n298 B.n175 163.367
R1508 B.n299 B.n298 163.367
R1509 B.n300 B.n299 163.367
R1510 B.n300 B.n173 163.367
R1511 B.n304 B.n173 163.367
R1512 B.n305 B.n304 163.367
R1513 B.n306 B.n305 163.367
R1514 B.n306 B.n171 163.367
R1515 B.n159 B.n158 82.0369
R1516 B.n359 B.n358 82.0369
R1517 B.n57 B.n56 82.0369
R1518 B.n51 B.n50 82.0369
R1519 B.n345 B.n159 59.5399
R1520 B.n360 B.n359 59.5399
R1521 B.n648 B.n57 59.5399
R1522 B.n662 B.n51 59.5399
R1523 B.n699 B.n698 32.9371
R1524 B.n612 B.n611 32.9371
R1525 B.n397 B.n140 32.9371
R1526 B.n309 B.n308 32.9371
R1527 B B.n805 18.0485
R1528 B.n699 B.n36 10.6151
R1529 B.n703 B.n36 10.6151
R1530 B.n704 B.n703 10.6151
R1531 B.n705 B.n704 10.6151
R1532 B.n705 B.n34 10.6151
R1533 B.n709 B.n34 10.6151
R1534 B.n710 B.n709 10.6151
R1535 B.n711 B.n710 10.6151
R1536 B.n711 B.n32 10.6151
R1537 B.n715 B.n32 10.6151
R1538 B.n716 B.n715 10.6151
R1539 B.n717 B.n716 10.6151
R1540 B.n717 B.n30 10.6151
R1541 B.n721 B.n30 10.6151
R1542 B.n722 B.n721 10.6151
R1543 B.n723 B.n722 10.6151
R1544 B.n723 B.n28 10.6151
R1545 B.n727 B.n28 10.6151
R1546 B.n728 B.n727 10.6151
R1547 B.n729 B.n728 10.6151
R1548 B.n729 B.n26 10.6151
R1549 B.n733 B.n26 10.6151
R1550 B.n734 B.n733 10.6151
R1551 B.n735 B.n734 10.6151
R1552 B.n735 B.n24 10.6151
R1553 B.n739 B.n24 10.6151
R1554 B.n740 B.n739 10.6151
R1555 B.n741 B.n740 10.6151
R1556 B.n741 B.n22 10.6151
R1557 B.n745 B.n22 10.6151
R1558 B.n746 B.n745 10.6151
R1559 B.n747 B.n746 10.6151
R1560 B.n747 B.n20 10.6151
R1561 B.n751 B.n20 10.6151
R1562 B.n752 B.n751 10.6151
R1563 B.n753 B.n752 10.6151
R1564 B.n753 B.n18 10.6151
R1565 B.n757 B.n18 10.6151
R1566 B.n758 B.n757 10.6151
R1567 B.n759 B.n758 10.6151
R1568 B.n759 B.n16 10.6151
R1569 B.n763 B.n16 10.6151
R1570 B.n764 B.n763 10.6151
R1571 B.n765 B.n764 10.6151
R1572 B.n765 B.n14 10.6151
R1573 B.n769 B.n14 10.6151
R1574 B.n770 B.n769 10.6151
R1575 B.n771 B.n770 10.6151
R1576 B.n771 B.n12 10.6151
R1577 B.n775 B.n12 10.6151
R1578 B.n776 B.n775 10.6151
R1579 B.n777 B.n776 10.6151
R1580 B.n777 B.n10 10.6151
R1581 B.n781 B.n10 10.6151
R1582 B.n782 B.n781 10.6151
R1583 B.n783 B.n782 10.6151
R1584 B.n783 B.n8 10.6151
R1585 B.n787 B.n8 10.6151
R1586 B.n788 B.n787 10.6151
R1587 B.n789 B.n788 10.6151
R1588 B.n789 B.n6 10.6151
R1589 B.n793 B.n6 10.6151
R1590 B.n794 B.n793 10.6151
R1591 B.n795 B.n794 10.6151
R1592 B.n795 B.n4 10.6151
R1593 B.n799 B.n4 10.6151
R1594 B.n800 B.n799 10.6151
R1595 B.n801 B.n800 10.6151
R1596 B.n801 B.n0 10.6151
R1597 B.n698 B.n697 10.6151
R1598 B.n697 B.n38 10.6151
R1599 B.n693 B.n38 10.6151
R1600 B.n693 B.n692 10.6151
R1601 B.n692 B.n691 10.6151
R1602 B.n691 B.n40 10.6151
R1603 B.n687 B.n40 10.6151
R1604 B.n687 B.n686 10.6151
R1605 B.n686 B.n685 10.6151
R1606 B.n685 B.n42 10.6151
R1607 B.n681 B.n42 10.6151
R1608 B.n681 B.n680 10.6151
R1609 B.n680 B.n679 10.6151
R1610 B.n679 B.n44 10.6151
R1611 B.n675 B.n44 10.6151
R1612 B.n675 B.n674 10.6151
R1613 B.n674 B.n673 10.6151
R1614 B.n673 B.n46 10.6151
R1615 B.n669 B.n46 10.6151
R1616 B.n669 B.n668 10.6151
R1617 B.n668 B.n667 10.6151
R1618 B.n667 B.n48 10.6151
R1619 B.n663 B.n48 10.6151
R1620 B.n661 B.n660 10.6151
R1621 B.n660 B.n52 10.6151
R1622 B.n656 B.n52 10.6151
R1623 B.n656 B.n655 10.6151
R1624 B.n655 B.n654 10.6151
R1625 B.n654 B.n54 10.6151
R1626 B.n650 B.n54 10.6151
R1627 B.n650 B.n649 10.6151
R1628 B.n647 B.n58 10.6151
R1629 B.n643 B.n58 10.6151
R1630 B.n643 B.n642 10.6151
R1631 B.n642 B.n641 10.6151
R1632 B.n641 B.n60 10.6151
R1633 B.n637 B.n60 10.6151
R1634 B.n637 B.n636 10.6151
R1635 B.n636 B.n635 10.6151
R1636 B.n635 B.n62 10.6151
R1637 B.n631 B.n62 10.6151
R1638 B.n631 B.n630 10.6151
R1639 B.n630 B.n629 10.6151
R1640 B.n629 B.n64 10.6151
R1641 B.n625 B.n64 10.6151
R1642 B.n625 B.n624 10.6151
R1643 B.n624 B.n623 10.6151
R1644 B.n623 B.n66 10.6151
R1645 B.n619 B.n66 10.6151
R1646 B.n619 B.n618 10.6151
R1647 B.n618 B.n617 10.6151
R1648 B.n617 B.n68 10.6151
R1649 B.n613 B.n68 10.6151
R1650 B.n613 B.n612 10.6151
R1651 B.n611 B.n70 10.6151
R1652 B.n607 B.n70 10.6151
R1653 B.n607 B.n606 10.6151
R1654 B.n606 B.n605 10.6151
R1655 B.n605 B.n72 10.6151
R1656 B.n601 B.n72 10.6151
R1657 B.n601 B.n600 10.6151
R1658 B.n600 B.n599 10.6151
R1659 B.n599 B.n74 10.6151
R1660 B.n595 B.n74 10.6151
R1661 B.n595 B.n594 10.6151
R1662 B.n594 B.n593 10.6151
R1663 B.n593 B.n76 10.6151
R1664 B.n589 B.n76 10.6151
R1665 B.n589 B.n588 10.6151
R1666 B.n588 B.n587 10.6151
R1667 B.n587 B.n78 10.6151
R1668 B.n583 B.n78 10.6151
R1669 B.n583 B.n582 10.6151
R1670 B.n582 B.n581 10.6151
R1671 B.n581 B.n80 10.6151
R1672 B.n577 B.n80 10.6151
R1673 B.n577 B.n576 10.6151
R1674 B.n576 B.n575 10.6151
R1675 B.n575 B.n82 10.6151
R1676 B.n571 B.n82 10.6151
R1677 B.n571 B.n570 10.6151
R1678 B.n570 B.n569 10.6151
R1679 B.n569 B.n84 10.6151
R1680 B.n565 B.n84 10.6151
R1681 B.n565 B.n564 10.6151
R1682 B.n564 B.n563 10.6151
R1683 B.n563 B.n86 10.6151
R1684 B.n559 B.n86 10.6151
R1685 B.n559 B.n558 10.6151
R1686 B.n558 B.n557 10.6151
R1687 B.n557 B.n88 10.6151
R1688 B.n553 B.n88 10.6151
R1689 B.n553 B.n552 10.6151
R1690 B.n552 B.n551 10.6151
R1691 B.n551 B.n90 10.6151
R1692 B.n547 B.n90 10.6151
R1693 B.n547 B.n546 10.6151
R1694 B.n546 B.n545 10.6151
R1695 B.n545 B.n92 10.6151
R1696 B.n541 B.n92 10.6151
R1697 B.n541 B.n540 10.6151
R1698 B.n540 B.n539 10.6151
R1699 B.n539 B.n94 10.6151
R1700 B.n535 B.n94 10.6151
R1701 B.n535 B.n534 10.6151
R1702 B.n534 B.n533 10.6151
R1703 B.n533 B.n96 10.6151
R1704 B.n529 B.n96 10.6151
R1705 B.n529 B.n528 10.6151
R1706 B.n528 B.n527 10.6151
R1707 B.n527 B.n98 10.6151
R1708 B.n523 B.n98 10.6151
R1709 B.n523 B.n522 10.6151
R1710 B.n522 B.n521 10.6151
R1711 B.n521 B.n100 10.6151
R1712 B.n517 B.n100 10.6151
R1713 B.n517 B.n516 10.6151
R1714 B.n516 B.n515 10.6151
R1715 B.n515 B.n102 10.6151
R1716 B.n511 B.n102 10.6151
R1717 B.n511 B.n510 10.6151
R1718 B.n510 B.n509 10.6151
R1719 B.n509 B.n104 10.6151
R1720 B.n505 B.n104 10.6151
R1721 B.n505 B.n504 10.6151
R1722 B.n504 B.n503 10.6151
R1723 B.n503 B.n106 10.6151
R1724 B.n499 B.n106 10.6151
R1725 B.n499 B.n498 10.6151
R1726 B.n498 B.n497 10.6151
R1727 B.n497 B.n108 10.6151
R1728 B.n493 B.n108 10.6151
R1729 B.n493 B.n492 10.6151
R1730 B.n492 B.n491 10.6151
R1731 B.n491 B.n110 10.6151
R1732 B.n487 B.n110 10.6151
R1733 B.n487 B.n486 10.6151
R1734 B.n486 B.n485 10.6151
R1735 B.n485 B.n112 10.6151
R1736 B.n481 B.n112 10.6151
R1737 B.n481 B.n480 10.6151
R1738 B.n480 B.n479 10.6151
R1739 B.n479 B.n114 10.6151
R1740 B.n475 B.n114 10.6151
R1741 B.n475 B.n474 10.6151
R1742 B.n474 B.n473 10.6151
R1743 B.n473 B.n116 10.6151
R1744 B.n469 B.n116 10.6151
R1745 B.n469 B.n468 10.6151
R1746 B.n468 B.n467 10.6151
R1747 B.n467 B.n118 10.6151
R1748 B.n463 B.n118 10.6151
R1749 B.n463 B.n462 10.6151
R1750 B.n462 B.n461 10.6151
R1751 B.n461 B.n120 10.6151
R1752 B.n457 B.n120 10.6151
R1753 B.n457 B.n456 10.6151
R1754 B.n456 B.n455 10.6151
R1755 B.n455 B.n122 10.6151
R1756 B.n451 B.n122 10.6151
R1757 B.n451 B.n450 10.6151
R1758 B.n450 B.n449 10.6151
R1759 B.n449 B.n124 10.6151
R1760 B.n445 B.n124 10.6151
R1761 B.n445 B.n444 10.6151
R1762 B.n444 B.n443 10.6151
R1763 B.n443 B.n126 10.6151
R1764 B.n439 B.n126 10.6151
R1765 B.n439 B.n438 10.6151
R1766 B.n438 B.n437 10.6151
R1767 B.n437 B.n128 10.6151
R1768 B.n433 B.n128 10.6151
R1769 B.n433 B.n432 10.6151
R1770 B.n432 B.n431 10.6151
R1771 B.n431 B.n130 10.6151
R1772 B.n427 B.n130 10.6151
R1773 B.n427 B.n426 10.6151
R1774 B.n426 B.n425 10.6151
R1775 B.n425 B.n132 10.6151
R1776 B.n421 B.n132 10.6151
R1777 B.n421 B.n420 10.6151
R1778 B.n420 B.n419 10.6151
R1779 B.n419 B.n134 10.6151
R1780 B.n415 B.n134 10.6151
R1781 B.n415 B.n414 10.6151
R1782 B.n414 B.n413 10.6151
R1783 B.n413 B.n136 10.6151
R1784 B.n409 B.n136 10.6151
R1785 B.n409 B.n408 10.6151
R1786 B.n408 B.n407 10.6151
R1787 B.n407 B.n138 10.6151
R1788 B.n403 B.n138 10.6151
R1789 B.n403 B.n402 10.6151
R1790 B.n402 B.n401 10.6151
R1791 B.n401 B.n140 10.6151
R1792 B.n206 B.n1 10.6151
R1793 B.n207 B.n206 10.6151
R1794 B.n207 B.n204 10.6151
R1795 B.n211 B.n204 10.6151
R1796 B.n212 B.n211 10.6151
R1797 B.n213 B.n212 10.6151
R1798 B.n213 B.n202 10.6151
R1799 B.n217 B.n202 10.6151
R1800 B.n218 B.n217 10.6151
R1801 B.n219 B.n218 10.6151
R1802 B.n219 B.n200 10.6151
R1803 B.n223 B.n200 10.6151
R1804 B.n224 B.n223 10.6151
R1805 B.n225 B.n224 10.6151
R1806 B.n225 B.n198 10.6151
R1807 B.n229 B.n198 10.6151
R1808 B.n230 B.n229 10.6151
R1809 B.n231 B.n230 10.6151
R1810 B.n231 B.n196 10.6151
R1811 B.n235 B.n196 10.6151
R1812 B.n236 B.n235 10.6151
R1813 B.n237 B.n236 10.6151
R1814 B.n237 B.n194 10.6151
R1815 B.n241 B.n194 10.6151
R1816 B.n242 B.n241 10.6151
R1817 B.n243 B.n242 10.6151
R1818 B.n243 B.n192 10.6151
R1819 B.n247 B.n192 10.6151
R1820 B.n248 B.n247 10.6151
R1821 B.n249 B.n248 10.6151
R1822 B.n249 B.n190 10.6151
R1823 B.n253 B.n190 10.6151
R1824 B.n254 B.n253 10.6151
R1825 B.n255 B.n254 10.6151
R1826 B.n255 B.n188 10.6151
R1827 B.n259 B.n188 10.6151
R1828 B.n260 B.n259 10.6151
R1829 B.n261 B.n260 10.6151
R1830 B.n261 B.n186 10.6151
R1831 B.n265 B.n186 10.6151
R1832 B.n266 B.n265 10.6151
R1833 B.n267 B.n266 10.6151
R1834 B.n267 B.n184 10.6151
R1835 B.n271 B.n184 10.6151
R1836 B.n272 B.n271 10.6151
R1837 B.n273 B.n272 10.6151
R1838 B.n273 B.n182 10.6151
R1839 B.n277 B.n182 10.6151
R1840 B.n278 B.n277 10.6151
R1841 B.n279 B.n278 10.6151
R1842 B.n279 B.n180 10.6151
R1843 B.n283 B.n180 10.6151
R1844 B.n284 B.n283 10.6151
R1845 B.n285 B.n284 10.6151
R1846 B.n285 B.n178 10.6151
R1847 B.n289 B.n178 10.6151
R1848 B.n290 B.n289 10.6151
R1849 B.n291 B.n290 10.6151
R1850 B.n291 B.n176 10.6151
R1851 B.n295 B.n176 10.6151
R1852 B.n296 B.n295 10.6151
R1853 B.n297 B.n296 10.6151
R1854 B.n297 B.n174 10.6151
R1855 B.n301 B.n174 10.6151
R1856 B.n302 B.n301 10.6151
R1857 B.n303 B.n302 10.6151
R1858 B.n303 B.n172 10.6151
R1859 B.n307 B.n172 10.6151
R1860 B.n308 B.n307 10.6151
R1861 B.n309 B.n170 10.6151
R1862 B.n313 B.n170 10.6151
R1863 B.n314 B.n313 10.6151
R1864 B.n315 B.n314 10.6151
R1865 B.n315 B.n168 10.6151
R1866 B.n319 B.n168 10.6151
R1867 B.n320 B.n319 10.6151
R1868 B.n321 B.n320 10.6151
R1869 B.n321 B.n166 10.6151
R1870 B.n325 B.n166 10.6151
R1871 B.n326 B.n325 10.6151
R1872 B.n327 B.n326 10.6151
R1873 B.n327 B.n164 10.6151
R1874 B.n331 B.n164 10.6151
R1875 B.n332 B.n331 10.6151
R1876 B.n333 B.n332 10.6151
R1877 B.n333 B.n162 10.6151
R1878 B.n337 B.n162 10.6151
R1879 B.n338 B.n337 10.6151
R1880 B.n339 B.n338 10.6151
R1881 B.n339 B.n160 10.6151
R1882 B.n343 B.n160 10.6151
R1883 B.n344 B.n343 10.6151
R1884 B.n346 B.n156 10.6151
R1885 B.n350 B.n156 10.6151
R1886 B.n351 B.n350 10.6151
R1887 B.n352 B.n351 10.6151
R1888 B.n352 B.n154 10.6151
R1889 B.n356 B.n154 10.6151
R1890 B.n357 B.n356 10.6151
R1891 B.n361 B.n357 10.6151
R1892 B.n365 B.n152 10.6151
R1893 B.n366 B.n365 10.6151
R1894 B.n367 B.n366 10.6151
R1895 B.n367 B.n150 10.6151
R1896 B.n371 B.n150 10.6151
R1897 B.n372 B.n371 10.6151
R1898 B.n373 B.n372 10.6151
R1899 B.n373 B.n148 10.6151
R1900 B.n377 B.n148 10.6151
R1901 B.n378 B.n377 10.6151
R1902 B.n379 B.n378 10.6151
R1903 B.n379 B.n146 10.6151
R1904 B.n383 B.n146 10.6151
R1905 B.n384 B.n383 10.6151
R1906 B.n385 B.n384 10.6151
R1907 B.n385 B.n144 10.6151
R1908 B.n389 B.n144 10.6151
R1909 B.n390 B.n389 10.6151
R1910 B.n391 B.n390 10.6151
R1911 B.n391 B.n142 10.6151
R1912 B.n395 B.n142 10.6151
R1913 B.n396 B.n395 10.6151
R1914 B.n397 B.n396 10.6151
R1915 B.n805 B.n0 8.11757
R1916 B.n805 B.n1 8.11757
R1917 B.n662 B.n661 6.5566
R1918 B.n649 B.n648 6.5566
R1919 B.n346 B.n345 6.5566
R1920 B.n361 B.n360 6.5566
R1921 B.n663 B.n662 4.05904
R1922 B.n648 B.n647 4.05904
R1923 B.n345 B.n344 4.05904
R1924 B.n360 B.n152 4.05904
C0 w_n5200_n2166# VDD1 2.20384f
C1 B VDD2 2.02192f
C2 VTAIL VDD2 7.08445f
C3 B VP 2.59575f
C4 VN VDD2 4.88907f
C5 VTAIL VP 6.25941f
C6 VDD1 VDD2 2.44979f
C7 VN VP 8.137799f
C8 VDD1 VP 5.39094f
C9 w_n5200_n2166# VDD2 2.37308f
C10 B VTAIL 3.40398f
C11 w_n5200_n2166# VP 11.5181f
C12 B VN 1.45075f
C13 B VDD1 1.88499f
C14 VN VTAIL 6.2453f
C15 VTAIL VDD1 7.02132f
C16 VN VDD1 0.153699f
C17 B w_n5200_n2166# 10.4358f
C18 VDD2 VP 0.657625f
C19 w_n5200_n2166# VTAIL 3.02354f
C20 w_n5200_n2166# VN 10.8392f
C21 VDD2 VSUBS 2.536212f
C22 VDD1 VSUBS 3.23287f
C23 VTAIL VSUBS 0.829044f
C24 VN VSUBS 8.27296f
C25 VP VSUBS 4.439299f
C26 B VSUBS 5.946345f
C27 w_n5200_n2166# VSUBS 0.140587p
C28 B.n0 VSUBS 0.009013f
C29 B.n1 VSUBS 0.009013f
C30 B.n2 VSUBS 0.01333f
C31 B.n3 VSUBS 0.010215f
C32 B.n4 VSUBS 0.010215f
C33 B.n5 VSUBS 0.010215f
C34 B.n6 VSUBS 0.010215f
C35 B.n7 VSUBS 0.010215f
C36 B.n8 VSUBS 0.010215f
C37 B.n9 VSUBS 0.010215f
C38 B.n10 VSUBS 0.010215f
C39 B.n11 VSUBS 0.010215f
C40 B.n12 VSUBS 0.010215f
C41 B.n13 VSUBS 0.010215f
C42 B.n14 VSUBS 0.010215f
C43 B.n15 VSUBS 0.010215f
C44 B.n16 VSUBS 0.010215f
C45 B.n17 VSUBS 0.010215f
C46 B.n18 VSUBS 0.010215f
C47 B.n19 VSUBS 0.010215f
C48 B.n20 VSUBS 0.010215f
C49 B.n21 VSUBS 0.010215f
C50 B.n22 VSUBS 0.010215f
C51 B.n23 VSUBS 0.010215f
C52 B.n24 VSUBS 0.010215f
C53 B.n25 VSUBS 0.010215f
C54 B.n26 VSUBS 0.010215f
C55 B.n27 VSUBS 0.010215f
C56 B.n28 VSUBS 0.010215f
C57 B.n29 VSUBS 0.010215f
C58 B.n30 VSUBS 0.010215f
C59 B.n31 VSUBS 0.010215f
C60 B.n32 VSUBS 0.010215f
C61 B.n33 VSUBS 0.010215f
C62 B.n34 VSUBS 0.010215f
C63 B.n35 VSUBS 0.010215f
C64 B.n36 VSUBS 0.010215f
C65 B.n37 VSUBS 0.024196f
C66 B.n38 VSUBS 0.010215f
C67 B.n39 VSUBS 0.010215f
C68 B.n40 VSUBS 0.010215f
C69 B.n41 VSUBS 0.010215f
C70 B.n42 VSUBS 0.010215f
C71 B.n43 VSUBS 0.010215f
C72 B.n44 VSUBS 0.010215f
C73 B.n45 VSUBS 0.010215f
C74 B.n46 VSUBS 0.010215f
C75 B.n47 VSUBS 0.010215f
C76 B.n48 VSUBS 0.010215f
C77 B.n49 VSUBS 0.010215f
C78 B.t1 VSUBS 0.130317f
C79 B.t2 VSUBS 0.182187f
C80 B.t0 VSUBS 1.64056f
C81 B.n50 VSUBS 0.29986f
C82 B.n51 VSUBS 0.235892f
C83 B.n52 VSUBS 0.010215f
C84 B.n53 VSUBS 0.010215f
C85 B.n54 VSUBS 0.010215f
C86 B.n55 VSUBS 0.010215f
C87 B.t7 VSUBS 0.13032f
C88 B.t8 VSUBS 0.182189f
C89 B.t6 VSUBS 1.64056f
C90 B.n56 VSUBS 0.299858f
C91 B.n57 VSUBS 0.235889f
C92 B.n58 VSUBS 0.010215f
C93 B.n59 VSUBS 0.010215f
C94 B.n60 VSUBS 0.010215f
C95 B.n61 VSUBS 0.010215f
C96 B.n62 VSUBS 0.010215f
C97 B.n63 VSUBS 0.010215f
C98 B.n64 VSUBS 0.010215f
C99 B.n65 VSUBS 0.010215f
C100 B.n66 VSUBS 0.010215f
C101 B.n67 VSUBS 0.010215f
C102 B.n68 VSUBS 0.010215f
C103 B.n69 VSUBS 0.024196f
C104 B.n70 VSUBS 0.010215f
C105 B.n71 VSUBS 0.010215f
C106 B.n72 VSUBS 0.010215f
C107 B.n73 VSUBS 0.010215f
C108 B.n74 VSUBS 0.010215f
C109 B.n75 VSUBS 0.010215f
C110 B.n76 VSUBS 0.010215f
C111 B.n77 VSUBS 0.010215f
C112 B.n78 VSUBS 0.010215f
C113 B.n79 VSUBS 0.010215f
C114 B.n80 VSUBS 0.010215f
C115 B.n81 VSUBS 0.010215f
C116 B.n82 VSUBS 0.010215f
C117 B.n83 VSUBS 0.010215f
C118 B.n84 VSUBS 0.010215f
C119 B.n85 VSUBS 0.010215f
C120 B.n86 VSUBS 0.010215f
C121 B.n87 VSUBS 0.010215f
C122 B.n88 VSUBS 0.010215f
C123 B.n89 VSUBS 0.010215f
C124 B.n90 VSUBS 0.010215f
C125 B.n91 VSUBS 0.010215f
C126 B.n92 VSUBS 0.010215f
C127 B.n93 VSUBS 0.010215f
C128 B.n94 VSUBS 0.010215f
C129 B.n95 VSUBS 0.010215f
C130 B.n96 VSUBS 0.010215f
C131 B.n97 VSUBS 0.010215f
C132 B.n98 VSUBS 0.010215f
C133 B.n99 VSUBS 0.010215f
C134 B.n100 VSUBS 0.010215f
C135 B.n101 VSUBS 0.010215f
C136 B.n102 VSUBS 0.010215f
C137 B.n103 VSUBS 0.010215f
C138 B.n104 VSUBS 0.010215f
C139 B.n105 VSUBS 0.010215f
C140 B.n106 VSUBS 0.010215f
C141 B.n107 VSUBS 0.010215f
C142 B.n108 VSUBS 0.010215f
C143 B.n109 VSUBS 0.010215f
C144 B.n110 VSUBS 0.010215f
C145 B.n111 VSUBS 0.010215f
C146 B.n112 VSUBS 0.010215f
C147 B.n113 VSUBS 0.010215f
C148 B.n114 VSUBS 0.010215f
C149 B.n115 VSUBS 0.010215f
C150 B.n116 VSUBS 0.010215f
C151 B.n117 VSUBS 0.010215f
C152 B.n118 VSUBS 0.010215f
C153 B.n119 VSUBS 0.010215f
C154 B.n120 VSUBS 0.010215f
C155 B.n121 VSUBS 0.010215f
C156 B.n122 VSUBS 0.010215f
C157 B.n123 VSUBS 0.010215f
C158 B.n124 VSUBS 0.010215f
C159 B.n125 VSUBS 0.010215f
C160 B.n126 VSUBS 0.010215f
C161 B.n127 VSUBS 0.010215f
C162 B.n128 VSUBS 0.010215f
C163 B.n129 VSUBS 0.010215f
C164 B.n130 VSUBS 0.010215f
C165 B.n131 VSUBS 0.010215f
C166 B.n132 VSUBS 0.010215f
C167 B.n133 VSUBS 0.010215f
C168 B.n134 VSUBS 0.010215f
C169 B.n135 VSUBS 0.010215f
C170 B.n136 VSUBS 0.010215f
C171 B.n137 VSUBS 0.010215f
C172 B.n138 VSUBS 0.010215f
C173 B.n139 VSUBS 0.010215f
C174 B.n140 VSUBS 0.025071f
C175 B.n141 VSUBS 0.010215f
C176 B.n142 VSUBS 0.010215f
C177 B.n143 VSUBS 0.010215f
C178 B.n144 VSUBS 0.010215f
C179 B.n145 VSUBS 0.010215f
C180 B.n146 VSUBS 0.010215f
C181 B.n147 VSUBS 0.010215f
C182 B.n148 VSUBS 0.010215f
C183 B.n149 VSUBS 0.010215f
C184 B.n150 VSUBS 0.010215f
C185 B.n151 VSUBS 0.010215f
C186 B.n152 VSUBS 0.00706f
C187 B.n153 VSUBS 0.010215f
C188 B.n154 VSUBS 0.010215f
C189 B.n155 VSUBS 0.010215f
C190 B.n156 VSUBS 0.010215f
C191 B.n157 VSUBS 0.010215f
C192 B.t11 VSUBS 0.130317f
C193 B.t10 VSUBS 0.182187f
C194 B.t9 VSUBS 1.64056f
C195 B.n158 VSUBS 0.29986f
C196 B.n159 VSUBS 0.235892f
C197 B.n160 VSUBS 0.010215f
C198 B.n161 VSUBS 0.010215f
C199 B.n162 VSUBS 0.010215f
C200 B.n163 VSUBS 0.010215f
C201 B.n164 VSUBS 0.010215f
C202 B.n165 VSUBS 0.010215f
C203 B.n166 VSUBS 0.010215f
C204 B.n167 VSUBS 0.010215f
C205 B.n168 VSUBS 0.010215f
C206 B.n169 VSUBS 0.010215f
C207 B.n170 VSUBS 0.010215f
C208 B.n171 VSUBS 0.023875f
C209 B.n172 VSUBS 0.010215f
C210 B.n173 VSUBS 0.010215f
C211 B.n174 VSUBS 0.010215f
C212 B.n175 VSUBS 0.010215f
C213 B.n176 VSUBS 0.010215f
C214 B.n177 VSUBS 0.010215f
C215 B.n178 VSUBS 0.010215f
C216 B.n179 VSUBS 0.010215f
C217 B.n180 VSUBS 0.010215f
C218 B.n181 VSUBS 0.010215f
C219 B.n182 VSUBS 0.010215f
C220 B.n183 VSUBS 0.010215f
C221 B.n184 VSUBS 0.010215f
C222 B.n185 VSUBS 0.010215f
C223 B.n186 VSUBS 0.010215f
C224 B.n187 VSUBS 0.010215f
C225 B.n188 VSUBS 0.010215f
C226 B.n189 VSUBS 0.010215f
C227 B.n190 VSUBS 0.010215f
C228 B.n191 VSUBS 0.010215f
C229 B.n192 VSUBS 0.010215f
C230 B.n193 VSUBS 0.010215f
C231 B.n194 VSUBS 0.010215f
C232 B.n195 VSUBS 0.010215f
C233 B.n196 VSUBS 0.010215f
C234 B.n197 VSUBS 0.010215f
C235 B.n198 VSUBS 0.010215f
C236 B.n199 VSUBS 0.010215f
C237 B.n200 VSUBS 0.010215f
C238 B.n201 VSUBS 0.010215f
C239 B.n202 VSUBS 0.010215f
C240 B.n203 VSUBS 0.010215f
C241 B.n204 VSUBS 0.010215f
C242 B.n205 VSUBS 0.010215f
C243 B.n206 VSUBS 0.010215f
C244 B.n207 VSUBS 0.010215f
C245 B.n208 VSUBS 0.010215f
C246 B.n209 VSUBS 0.010215f
C247 B.n210 VSUBS 0.010215f
C248 B.n211 VSUBS 0.010215f
C249 B.n212 VSUBS 0.010215f
C250 B.n213 VSUBS 0.010215f
C251 B.n214 VSUBS 0.010215f
C252 B.n215 VSUBS 0.010215f
C253 B.n216 VSUBS 0.010215f
C254 B.n217 VSUBS 0.010215f
C255 B.n218 VSUBS 0.010215f
C256 B.n219 VSUBS 0.010215f
C257 B.n220 VSUBS 0.010215f
C258 B.n221 VSUBS 0.010215f
C259 B.n222 VSUBS 0.010215f
C260 B.n223 VSUBS 0.010215f
C261 B.n224 VSUBS 0.010215f
C262 B.n225 VSUBS 0.010215f
C263 B.n226 VSUBS 0.010215f
C264 B.n227 VSUBS 0.010215f
C265 B.n228 VSUBS 0.010215f
C266 B.n229 VSUBS 0.010215f
C267 B.n230 VSUBS 0.010215f
C268 B.n231 VSUBS 0.010215f
C269 B.n232 VSUBS 0.010215f
C270 B.n233 VSUBS 0.010215f
C271 B.n234 VSUBS 0.010215f
C272 B.n235 VSUBS 0.010215f
C273 B.n236 VSUBS 0.010215f
C274 B.n237 VSUBS 0.010215f
C275 B.n238 VSUBS 0.010215f
C276 B.n239 VSUBS 0.010215f
C277 B.n240 VSUBS 0.010215f
C278 B.n241 VSUBS 0.010215f
C279 B.n242 VSUBS 0.010215f
C280 B.n243 VSUBS 0.010215f
C281 B.n244 VSUBS 0.010215f
C282 B.n245 VSUBS 0.010215f
C283 B.n246 VSUBS 0.010215f
C284 B.n247 VSUBS 0.010215f
C285 B.n248 VSUBS 0.010215f
C286 B.n249 VSUBS 0.010215f
C287 B.n250 VSUBS 0.010215f
C288 B.n251 VSUBS 0.010215f
C289 B.n252 VSUBS 0.010215f
C290 B.n253 VSUBS 0.010215f
C291 B.n254 VSUBS 0.010215f
C292 B.n255 VSUBS 0.010215f
C293 B.n256 VSUBS 0.010215f
C294 B.n257 VSUBS 0.010215f
C295 B.n258 VSUBS 0.010215f
C296 B.n259 VSUBS 0.010215f
C297 B.n260 VSUBS 0.010215f
C298 B.n261 VSUBS 0.010215f
C299 B.n262 VSUBS 0.010215f
C300 B.n263 VSUBS 0.010215f
C301 B.n264 VSUBS 0.010215f
C302 B.n265 VSUBS 0.010215f
C303 B.n266 VSUBS 0.010215f
C304 B.n267 VSUBS 0.010215f
C305 B.n268 VSUBS 0.010215f
C306 B.n269 VSUBS 0.010215f
C307 B.n270 VSUBS 0.010215f
C308 B.n271 VSUBS 0.010215f
C309 B.n272 VSUBS 0.010215f
C310 B.n273 VSUBS 0.010215f
C311 B.n274 VSUBS 0.010215f
C312 B.n275 VSUBS 0.010215f
C313 B.n276 VSUBS 0.010215f
C314 B.n277 VSUBS 0.010215f
C315 B.n278 VSUBS 0.010215f
C316 B.n279 VSUBS 0.010215f
C317 B.n280 VSUBS 0.010215f
C318 B.n281 VSUBS 0.010215f
C319 B.n282 VSUBS 0.010215f
C320 B.n283 VSUBS 0.010215f
C321 B.n284 VSUBS 0.010215f
C322 B.n285 VSUBS 0.010215f
C323 B.n286 VSUBS 0.010215f
C324 B.n287 VSUBS 0.010215f
C325 B.n288 VSUBS 0.010215f
C326 B.n289 VSUBS 0.010215f
C327 B.n290 VSUBS 0.010215f
C328 B.n291 VSUBS 0.010215f
C329 B.n292 VSUBS 0.010215f
C330 B.n293 VSUBS 0.010215f
C331 B.n294 VSUBS 0.010215f
C332 B.n295 VSUBS 0.010215f
C333 B.n296 VSUBS 0.010215f
C334 B.n297 VSUBS 0.010215f
C335 B.n298 VSUBS 0.010215f
C336 B.n299 VSUBS 0.010215f
C337 B.n300 VSUBS 0.010215f
C338 B.n301 VSUBS 0.010215f
C339 B.n302 VSUBS 0.010215f
C340 B.n303 VSUBS 0.010215f
C341 B.n304 VSUBS 0.010215f
C342 B.n305 VSUBS 0.010215f
C343 B.n306 VSUBS 0.010215f
C344 B.n307 VSUBS 0.010215f
C345 B.n308 VSUBS 0.023875f
C346 B.n309 VSUBS 0.024196f
C347 B.n310 VSUBS 0.024196f
C348 B.n311 VSUBS 0.010215f
C349 B.n312 VSUBS 0.010215f
C350 B.n313 VSUBS 0.010215f
C351 B.n314 VSUBS 0.010215f
C352 B.n315 VSUBS 0.010215f
C353 B.n316 VSUBS 0.010215f
C354 B.n317 VSUBS 0.010215f
C355 B.n318 VSUBS 0.010215f
C356 B.n319 VSUBS 0.010215f
C357 B.n320 VSUBS 0.010215f
C358 B.n321 VSUBS 0.010215f
C359 B.n322 VSUBS 0.010215f
C360 B.n323 VSUBS 0.010215f
C361 B.n324 VSUBS 0.010215f
C362 B.n325 VSUBS 0.010215f
C363 B.n326 VSUBS 0.010215f
C364 B.n327 VSUBS 0.010215f
C365 B.n328 VSUBS 0.010215f
C366 B.n329 VSUBS 0.010215f
C367 B.n330 VSUBS 0.010215f
C368 B.n331 VSUBS 0.010215f
C369 B.n332 VSUBS 0.010215f
C370 B.n333 VSUBS 0.010215f
C371 B.n334 VSUBS 0.010215f
C372 B.n335 VSUBS 0.010215f
C373 B.n336 VSUBS 0.010215f
C374 B.n337 VSUBS 0.010215f
C375 B.n338 VSUBS 0.010215f
C376 B.n339 VSUBS 0.010215f
C377 B.n340 VSUBS 0.010215f
C378 B.n341 VSUBS 0.010215f
C379 B.n342 VSUBS 0.010215f
C380 B.n343 VSUBS 0.010215f
C381 B.n344 VSUBS 0.00706f
C382 B.n345 VSUBS 0.023667f
C383 B.n346 VSUBS 0.008262f
C384 B.n347 VSUBS 0.010215f
C385 B.n348 VSUBS 0.010215f
C386 B.n349 VSUBS 0.010215f
C387 B.n350 VSUBS 0.010215f
C388 B.n351 VSUBS 0.010215f
C389 B.n352 VSUBS 0.010215f
C390 B.n353 VSUBS 0.010215f
C391 B.n354 VSUBS 0.010215f
C392 B.n355 VSUBS 0.010215f
C393 B.n356 VSUBS 0.010215f
C394 B.n357 VSUBS 0.010215f
C395 B.t5 VSUBS 0.13032f
C396 B.t4 VSUBS 0.182189f
C397 B.t3 VSUBS 1.64056f
C398 B.n358 VSUBS 0.299858f
C399 B.n359 VSUBS 0.235889f
C400 B.n360 VSUBS 0.023667f
C401 B.n361 VSUBS 0.008262f
C402 B.n362 VSUBS 0.010215f
C403 B.n363 VSUBS 0.010215f
C404 B.n364 VSUBS 0.010215f
C405 B.n365 VSUBS 0.010215f
C406 B.n366 VSUBS 0.010215f
C407 B.n367 VSUBS 0.010215f
C408 B.n368 VSUBS 0.010215f
C409 B.n369 VSUBS 0.010215f
C410 B.n370 VSUBS 0.010215f
C411 B.n371 VSUBS 0.010215f
C412 B.n372 VSUBS 0.010215f
C413 B.n373 VSUBS 0.010215f
C414 B.n374 VSUBS 0.010215f
C415 B.n375 VSUBS 0.010215f
C416 B.n376 VSUBS 0.010215f
C417 B.n377 VSUBS 0.010215f
C418 B.n378 VSUBS 0.010215f
C419 B.n379 VSUBS 0.010215f
C420 B.n380 VSUBS 0.010215f
C421 B.n381 VSUBS 0.010215f
C422 B.n382 VSUBS 0.010215f
C423 B.n383 VSUBS 0.010215f
C424 B.n384 VSUBS 0.010215f
C425 B.n385 VSUBS 0.010215f
C426 B.n386 VSUBS 0.010215f
C427 B.n387 VSUBS 0.010215f
C428 B.n388 VSUBS 0.010215f
C429 B.n389 VSUBS 0.010215f
C430 B.n390 VSUBS 0.010215f
C431 B.n391 VSUBS 0.010215f
C432 B.n392 VSUBS 0.010215f
C433 B.n393 VSUBS 0.010215f
C434 B.n394 VSUBS 0.010215f
C435 B.n395 VSUBS 0.010215f
C436 B.n396 VSUBS 0.010215f
C437 B.n397 VSUBS 0.022999f
C438 B.n398 VSUBS 0.024196f
C439 B.n399 VSUBS 0.023875f
C440 B.n400 VSUBS 0.010215f
C441 B.n401 VSUBS 0.010215f
C442 B.n402 VSUBS 0.010215f
C443 B.n403 VSUBS 0.010215f
C444 B.n404 VSUBS 0.010215f
C445 B.n405 VSUBS 0.010215f
C446 B.n406 VSUBS 0.010215f
C447 B.n407 VSUBS 0.010215f
C448 B.n408 VSUBS 0.010215f
C449 B.n409 VSUBS 0.010215f
C450 B.n410 VSUBS 0.010215f
C451 B.n411 VSUBS 0.010215f
C452 B.n412 VSUBS 0.010215f
C453 B.n413 VSUBS 0.010215f
C454 B.n414 VSUBS 0.010215f
C455 B.n415 VSUBS 0.010215f
C456 B.n416 VSUBS 0.010215f
C457 B.n417 VSUBS 0.010215f
C458 B.n418 VSUBS 0.010215f
C459 B.n419 VSUBS 0.010215f
C460 B.n420 VSUBS 0.010215f
C461 B.n421 VSUBS 0.010215f
C462 B.n422 VSUBS 0.010215f
C463 B.n423 VSUBS 0.010215f
C464 B.n424 VSUBS 0.010215f
C465 B.n425 VSUBS 0.010215f
C466 B.n426 VSUBS 0.010215f
C467 B.n427 VSUBS 0.010215f
C468 B.n428 VSUBS 0.010215f
C469 B.n429 VSUBS 0.010215f
C470 B.n430 VSUBS 0.010215f
C471 B.n431 VSUBS 0.010215f
C472 B.n432 VSUBS 0.010215f
C473 B.n433 VSUBS 0.010215f
C474 B.n434 VSUBS 0.010215f
C475 B.n435 VSUBS 0.010215f
C476 B.n436 VSUBS 0.010215f
C477 B.n437 VSUBS 0.010215f
C478 B.n438 VSUBS 0.010215f
C479 B.n439 VSUBS 0.010215f
C480 B.n440 VSUBS 0.010215f
C481 B.n441 VSUBS 0.010215f
C482 B.n442 VSUBS 0.010215f
C483 B.n443 VSUBS 0.010215f
C484 B.n444 VSUBS 0.010215f
C485 B.n445 VSUBS 0.010215f
C486 B.n446 VSUBS 0.010215f
C487 B.n447 VSUBS 0.010215f
C488 B.n448 VSUBS 0.010215f
C489 B.n449 VSUBS 0.010215f
C490 B.n450 VSUBS 0.010215f
C491 B.n451 VSUBS 0.010215f
C492 B.n452 VSUBS 0.010215f
C493 B.n453 VSUBS 0.010215f
C494 B.n454 VSUBS 0.010215f
C495 B.n455 VSUBS 0.010215f
C496 B.n456 VSUBS 0.010215f
C497 B.n457 VSUBS 0.010215f
C498 B.n458 VSUBS 0.010215f
C499 B.n459 VSUBS 0.010215f
C500 B.n460 VSUBS 0.010215f
C501 B.n461 VSUBS 0.010215f
C502 B.n462 VSUBS 0.010215f
C503 B.n463 VSUBS 0.010215f
C504 B.n464 VSUBS 0.010215f
C505 B.n465 VSUBS 0.010215f
C506 B.n466 VSUBS 0.010215f
C507 B.n467 VSUBS 0.010215f
C508 B.n468 VSUBS 0.010215f
C509 B.n469 VSUBS 0.010215f
C510 B.n470 VSUBS 0.010215f
C511 B.n471 VSUBS 0.010215f
C512 B.n472 VSUBS 0.010215f
C513 B.n473 VSUBS 0.010215f
C514 B.n474 VSUBS 0.010215f
C515 B.n475 VSUBS 0.010215f
C516 B.n476 VSUBS 0.010215f
C517 B.n477 VSUBS 0.010215f
C518 B.n478 VSUBS 0.010215f
C519 B.n479 VSUBS 0.010215f
C520 B.n480 VSUBS 0.010215f
C521 B.n481 VSUBS 0.010215f
C522 B.n482 VSUBS 0.010215f
C523 B.n483 VSUBS 0.010215f
C524 B.n484 VSUBS 0.010215f
C525 B.n485 VSUBS 0.010215f
C526 B.n486 VSUBS 0.010215f
C527 B.n487 VSUBS 0.010215f
C528 B.n488 VSUBS 0.010215f
C529 B.n489 VSUBS 0.010215f
C530 B.n490 VSUBS 0.010215f
C531 B.n491 VSUBS 0.010215f
C532 B.n492 VSUBS 0.010215f
C533 B.n493 VSUBS 0.010215f
C534 B.n494 VSUBS 0.010215f
C535 B.n495 VSUBS 0.010215f
C536 B.n496 VSUBS 0.010215f
C537 B.n497 VSUBS 0.010215f
C538 B.n498 VSUBS 0.010215f
C539 B.n499 VSUBS 0.010215f
C540 B.n500 VSUBS 0.010215f
C541 B.n501 VSUBS 0.010215f
C542 B.n502 VSUBS 0.010215f
C543 B.n503 VSUBS 0.010215f
C544 B.n504 VSUBS 0.010215f
C545 B.n505 VSUBS 0.010215f
C546 B.n506 VSUBS 0.010215f
C547 B.n507 VSUBS 0.010215f
C548 B.n508 VSUBS 0.010215f
C549 B.n509 VSUBS 0.010215f
C550 B.n510 VSUBS 0.010215f
C551 B.n511 VSUBS 0.010215f
C552 B.n512 VSUBS 0.010215f
C553 B.n513 VSUBS 0.010215f
C554 B.n514 VSUBS 0.010215f
C555 B.n515 VSUBS 0.010215f
C556 B.n516 VSUBS 0.010215f
C557 B.n517 VSUBS 0.010215f
C558 B.n518 VSUBS 0.010215f
C559 B.n519 VSUBS 0.010215f
C560 B.n520 VSUBS 0.010215f
C561 B.n521 VSUBS 0.010215f
C562 B.n522 VSUBS 0.010215f
C563 B.n523 VSUBS 0.010215f
C564 B.n524 VSUBS 0.010215f
C565 B.n525 VSUBS 0.010215f
C566 B.n526 VSUBS 0.010215f
C567 B.n527 VSUBS 0.010215f
C568 B.n528 VSUBS 0.010215f
C569 B.n529 VSUBS 0.010215f
C570 B.n530 VSUBS 0.010215f
C571 B.n531 VSUBS 0.010215f
C572 B.n532 VSUBS 0.010215f
C573 B.n533 VSUBS 0.010215f
C574 B.n534 VSUBS 0.010215f
C575 B.n535 VSUBS 0.010215f
C576 B.n536 VSUBS 0.010215f
C577 B.n537 VSUBS 0.010215f
C578 B.n538 VSUBS 0.010215f
C579 B.n539 VSUBS 0.010215f
C580 B.n540 VSUBS 0.010215f
C581 B.n541 VSUBS 0.010215f
C582 B.n542 VSUBS 0.010215f
C583 B.n543 VSUBS 0.010215f
C584 B.n544 VSUBS 0.010215f
C585 B.n545 VSUBS 0.010215f
C586 B.n546 VSUBS 0.010215f
C587 B.n547 VSUBS 0.010215f
C588 B.n548 VSUBS 0.010215f
C589 B.n549 VSUBS 0.010215f
C590 B.n550 VSUBS 0.010215f
C591 B.n551 VSUBS 0.010215f
C592 B.n552 VSUBS 0.010215f
C593 B.n553 VSUBS 0.010215f
C594 B.n554 VSUBS 0.010215f
C595 B.n555 VSUBS 0.010215f
C596 B.n556 VSUBS 0.010215f
C597 B.n557 VSUBS 0.010215f
C598 B.n558 VSUBS 0.010215f
C599 B.n559 VSUBS 0.010215f
C600 B.n560 VSUBS 0.010215f
C601 B.n561 VSUBS 0.010215f
C602 B.n562 VSUBS 0.010215f
C603 B.n563 VSUBS 0.010215f
C604 B.n564 VSUBS 0.010215f
C605 B.n565 VSUBS 0.010215f
C606 B.n566 VSUBS 0.010215f
C607 B.n567 VSUBS 0.010215f
C608 B.n568 VSUBS 0.010215f
C609 B.n569 VSUBS 0.010215f
C610 B.n570 VSUBS 0.010215f
C611 B.n571 VSUBS 0.010215f
C612 B.n572 VSUBS 0.010215f
C613 B.n573 VSUBS 0.010215f
C614 B.n574 VSUBS 0.010215f
C615 B.n575 VSUBS 0.010215f
C616 B.n576 VSUBS 0.010215f
C617 B.n577 VSUBS 0.010215f
C618 B.n578 VSUBS 0.010215f
C619 B.n579 VSUBS 0.010215f
C620 B.n580 VSUBS 0.010215f
C621 B.n581 VSUBS 0.010215f
C622 B.n582 VSUBS 0.010215f
C623 B.n583 VSUBS 0.010215f
C624 B.n584 VSUBS 0.010215f
C625 B.n585 VSUBS 0.010215f
C626 B.n586 VSUBS 0.010215f
C627 B.n587 VSUBS 0.010215f
C628 B.n588 VSUBS 0.010215f
C629 B.n589 VSUBS 0.010215f
C630 B.n590 VSUBS 0.010215f
C631 B.n591 VSUBS 0.010215f
C632 B.n592 VSUBS 0.010215f
C633 B.n593 VSUBS 0.010215f
C634 B.n594 VSUBS 0.010215f
C635 B.n595 VSUBS 0.010215f
C636 B.n596 VSUBS 0.010215f
C637 B.n597 VSUBS 0.010215f
C638 B.n598 VSUBS 0.010215f
C639 B.n599 VSUBS 0.010215f
C640 B.n600 VSUBS 0.010215f
C641 B.n601 VSUBS 0.010215f
C642 B.n602 VSUBS 0.010215f
C643 B.n603 VSUBS 0.010215f
C644 B.n604 VSUBS 0.010215f
C645 B.n605 VSUBS 0.010215f
C646 B.n606 VSUBS 0.010215f
C647 B.n607 VSUBS 0.010215f
C648 B.n608 VSUBS 0.010215f
C649 B.n609 VSUBS 0.010215f
C650 B.n610 VSUBS 0.023875f
C651 B.n611 VSUBS 0.023875f
C652 B.n612 VSUBS 0.024196f
C653 B.n613 VSUBS 0.010215f
C654 B.n614 VSUBS 0.010215f
C655 B.n615 VSUBS 0.010215f
C656 B.n616 VSUBS 0.010215f
C657 B.n617 VSUBS 0.010215f
C658 B.n618 VSUBS 0.010215f
C659 B.n619 VSUBS 0.010215f
C660 B.n620 VSUBS 0.010215f
C661 B.n621 VSUBS 0.010215f
C662 B.n622 VSUBS 0.010215f
C663 B.n623 VSUBS 0.010215f
C664 B.n624 VSUBS 0.010215f
C665 B.n625 VSUBS 0.010215f
C666 B.n626 VSUBS 0.010215f
C667 B.n627 VSUBS 0.010215f
C668 B.n628 VSUBS 0.010215f
C669 B.n629 VSUBS 0.010215f
C670 B.n630 VSUBS 0.010215f
C671 B.n631 VSUBS 0.010215f
C672 B.n632 VSUBS 0.010215f
C673 B.n633 VSUBS 0.010215f
C674 B.n634 VSUBS 0.010215f
C675 B.n635 VSUBS 0.010215f
C676 B.n636 VSUBS 0.010215f
C677 B.n637 VSUBS 0.010215f
C678 B.n638 VSUBS 0.010215f
C679 B.n639 VSUBS 0.010215f
C680 B.n640 VSUBS 0.010215f
C681 B.n641 VSUBS 0.010215f
C682 B.n642 VSUBS 0.010215f
C683 B.n643 VSUBS 0.010215f
C684 B.n644 VSUBS 0.010215f
C685 B.n645 VSUBS 0.010215f
C686 B.n646 VSUBS 0.010215f
C687 B.n647 VSUBS 0.00706f
C688 B.n648 VSUBS 0.023667f
C689 B.n649 VSUBS 0.008262f
C690 B.n650 VSUBS 0.010215f
C691 B.n651 VSUBS 0.010215f
C692 B.n652 VSUBS 0.010215f
C693 B.n653 VSUBS 0.010215f
C694 B.n654 VSUBS 0.010215f
C695 B.n655 VSUBS 0.010215f
C696 B.n656 VSUBS 0.010215f
C697 B.n657 VSUBS 0.010215f
C698 B.n658 VSUBS 0.010215f
C699 B.n659 VSUBS 0.010215f
C700 B.n660 VSUBS 0.010215f
C701 B.n661 VSUBS 0.008262f
C702 B.n662 VSUBS 0.023667f
C703 B.n663 VSUBS 0.00706f
C704 B.n664 VSUBS 0.010215f
C705 B.n665 VSUBS 0.010215f
C706 B.n666 VSUBS 0.010215f
C707 B.n667 VSUBS 0.010215f
C708 B.n668 VSUBS 0.010215f
C709 B.n669 VSUBS 0.010215f
C710 B.n670 VSUBS 0.010215f
C711 B.n671 VSUBS 0.010215f
C712 B.n672 VSUBS 0.010215f
C713 B.n673 VSUBS 0.010215f
C714 B.n674 VSUBS 0.010215f
C715 B.n675 VSUBS 0.010215f
C716 B.n676 VSUBS 0.010215f
C717 B.n677 VSUBS 0.010215f
C718 B.n678 VSUBS 0.010215f
C719 B.n679 VSUBS 0.010215f
C720 B.n680 VSUBS 0.010215f
C721 B.n681 VSUBS 0.010215f
C722 B.n682 VSUBS 0.010215f
C723 B.n683 VSUBS 0.010215f
C724 B.n684 VSUBS 0.010215f
C725 B.n685 VSUBS 0.010215f
C726 B.n686 VSUBS 0.010215f
C727 B.n687 VSUBS 0.010215f
C728 B.n688 VSUBS 0.010215f
C729 B.n689 VSUBS 0.010215f
C730 B.n690 VSUBS 0.010215f
C731 B.n691 VSUBS 0.010215f
C732 B.n692 VSUBS 0.010215f
C733 B.n693 VSUBS 0.010215f
C734 B.n694 VSUBS 0.010215f
C735 B.n695 VSUBS 0.010215f
C736 B.n696 VSUBS 0.010215f
C737 B.n697 VSUBS 0.010215f
C738 B.n698 VSUBS 0.024196f
C739 B.n699 VSUBS 0.023875f
C740 B.n700 VSUBS 0.023875f
C741 B.n701 VSUBS 0.010215f
C742 B.n702 VSUBS 0.010215f
C743 B.n703 VSUBS 0.010215f
C744 B.n704 VSUBS 0.010215f
C745 B.n705 VSUBS 0.010215f
C746 B.n706 VSUBS 0.010215f
C747 B.n707 VSUBS 0.010215f
C748 B.n708 VSUBS 0.010215f
C749 B.n709 VSUBS 0.010215f
C750 B.n710 VSUBS 0.010215f
C751 B.n711 VSUBS 0.010215f
C752 B.n712 VSUBS 0.010215f
C753 B.n713 VSUBS 0.010215f
C754 B.n714 VSUBS 0.010215f
C755 B.n715 VSUBS 0.010215f
C756 B.n716 VSUBS 0.010215f
C757 B.n717 VSUBS 0.010215f
C758 B.n718 VSUBS 0.010215f
C759 B.n719 VSUBS 0.010215f
C760 B.n720 VSUBS 0.010215f
C761 B.n721 VSUBS 0.010215f
C762 B.n722 VSUBS 0.010215f
C763 B.n723 VSUBS 0.010215f
C764 B.n724 VSUBS 0.010215f
C765 B.n725 VSUBS 0.010215f
C766 B.n726 VSUBS 0.010215f
C767 B.n727 VSUBS 0.010215f
C768 B.n728 VSUBS 0.010215f
C769 B.n729 VSUBS 0.010215f
C770 B.n730 VSUBS 0.010215f
C771 B.n731 VSUBS 0.010215f
C772 B.n732 VSUBS 0.010215f
C773 B.n733 VSUBS 0.010215f
C774 B.n734 VSUBS 0.010215f
C775 B.n735 VSUBS 0.010215f
C776 B.n736 VSUBS 0.010215f
C777 B.n737 VSUBS 0.010215f
C778 B.n738 VSUBS 0.010215f
C779 B.n739 VSUBS 0.010215f
C780 B.n740 VSUBS 0.010215f
C781 B.n741 VSUBS 0.010215f
C782 B.n742 VSUBS 0.010215f
C783 B.n743 VSUBS 0.010215f
C784 B.n744 VSUBS 0.010215f
C785 B.n745 VSUBS 0.010215f
C786 B.n746 VSUBS 0.010215f
C787 B.n747 VSUBS 0.010215f
C788 B.n748 VSUBS 0.010215f
C789 B.n749 VSUBS 0.010215f
C790 B.n750 VSUBS 0.010215f
C791 B.n751 VSUBS 0.010215f
C792 B.n752 VSUBS 0.010215f
C793 B.n753 VSUBS 0.010215f
C794 B.n754 VSUBS 0.010215f
C795 B.n755 VSUBS 0.010215f
C796 B.n756 VSUBS 0.010215f
C797 B.n757 VSUBS 0.010215f
C798 B.n758 VSUBS 0.010215f
C799 B.n759 VSUBS 0.010215f
C800 B.n760 VSUBS 0.010215f
C801 B.n761 VSUBS 0.010215f
C802 B.n762 VSUBS 0.010215f
C803 B.n763 VSUBS 0.010215f
C804 B.n764 VSUBS 0.010215f
C805 B.n765 VSUBS 0.010215f
C806 B.n766 VSUBS 0.010215f
C807 B.n767 VSUBS 0.010215f
C808 B.n768 VSUBS 0.010215f
C809 B.n769 VSUBS 0.010215f
C810 B.n770 VSUBS 0.010215f
C811 B.n771 VSUBS 0.010215f
C812 B.n772 VSUBS 0.010215f
C813 B.n773 VSUBS 0.010215f
C814 B.n774 VSUBS 0.010215f
C815 B.n775 VSUBS 0.010215f
C816 B.n776 VSUBS 0.010215f
C817 B.n777 VSUBS 0.010215f
C818 B.n778 VSUBS 0.010215f
C819 B.n779 VSUBS 0.010215f
C820 B.n780 VSUBS 0.010215f
C821 B.n781 VSUBS 0.010215f
C822 B.n782 VSUBS 0.010215f
C823 B.n783 VSUBS 0.010215f
C824 B.n784 VSUBS 0.010215f
C825 B.n785 VSUBS 0.010215f
C826 B.n786 VSUBS 0.010215f
C827 B.n787 VSUBS 0.010215f
C828 B.n788 VSUBS 0.010215f
C829 B.n789 VSUBS 0.010215f
C830 B.n790 VSUBS 0.010215f
C831 B.n791 VSUBS 0.010215f
C832 B.n792 VSUBS 0.010215f
C833 B.n793 VSUBS 0.010215f
C834 B.n794 VSUBS 0.010215f
C835 B.n795 VSUBS 0.010215f
C836 B.n796 VSUBS 0.010215f
C837 B.n797 VSUBS 0.010215f
C838 B.n798 VSUBS 0.010215f
C839 B.n799 VSUBS 0.010215f
C840 B.n800 VSUBS 0.010215f
C841 B.n801 VSUBS 0.010215f
C842 B.n802 VSUBS 0.010215f
C843 B.n803 VSUBS 0.01333f
C844 B.n804 VSUBS 0.0142f
C845 B.n805 VSUBS 0.028238f
C846 VDD2.t0 VSUBS 0.178564f
C847 VDD2.t4 VSUBS 0.178564f
C848 VDD2.n0 VSUBS 1.20607f
C849 VDD2.t1 VSUBS 0.178564f
C850 VDD2.t6 VSUBS 0.178564f
C851 VDD2.n1 VSUBS 1.20607f
C852 VDD2.n2 VSUBS 6.12371f
C853 VDD2.t2 VSUBS 0.178564f
C854 VDD2.t7 VSUBS 0.178564f
C855 VDD2.n3 VSUBS 1.18184f
C856 VDD2.n4 VSUBS 4.7425f
C857 VDD2.t5 VSUBS 0.178564f
C858 VDD2.t3 VSUBS 0.178564f
C859 VDD2.n5 VSUBS 1.20602f
C860 VN.t1 VSUBS 1.91532f
C861 VN.n0 VSUBS 0.826766f
C862 VN.n1 VSUBS 0.03098f
C863 VN.n2 VSUBS 0.06211f
C864 VN.n3 VSUBS 0.03098f
C865 VN.n4 VSUBS 0.057738f
C866 VN.n5 VSUBS 0.03098f
C867 VN.t6 VSUBS 1.91532f
C868 VN.n6 VSUBS 0.057738f
C869 VN.n7 VSUBS 0.03098f
C870 VN.n8 VSUBS 0.057738f
C871 VN.t7 VSUBS 2.36791f
C872 VN.n9 VSUBS 0.798205f
C873 VN.t3 VSUBS 1.91532f
C874 VN.n10 VSUBS 0.823674f
C875 VN.n11 VSUBS 0.05004f
C876 VN.n12 VSUBS 0.400826f
C877 VN.n13 VSUBS 0.03098f
C878 VN.n14 VSUBS 0.03098f
C879 VN.n15 VSUBS 0.057738f
C880 VN.n16 VSUBS 0.045225f
C881 VN.n17 VSUBS 0.045225f
C882 VN.n18 VSUBS 0.03098f
C883 VN.n19 VSUBS 0.03098f
C884 VN.n20 VSUBS 0.03098f
C885 VN.n21 VSUBS 0.057738f
C886 VN.n22 VSUBS 0.05004f
C887 VN.n23 VSUBS 0.704566f
C888 VN.n24 VSUBS 0.036928f
C889 VN.n25 VSUBS 0.03098f
C890 VN.n26 VSUBS 0.03098f
C891 VN.n27 VSUBS 0.03098f
C892 VN.n28 VSUBS 0.057738f
C893 VN.n29 VSUBS 0.060874f
C894 VN.n30 VSUBS 0.025204f
C895 VN.n31 VSUBS 0.03098f
C896 VN.n32 VSUBS 0.03098f
C897 VN.n33 VSUBS 0.03098f
C898 VN.n34 VSUBS 0.057738f
C899 VN.n35 VSUBS 0.057738f
C900 VN.n36 VSUBS 0.034647f
C901 VN.n37 VSUBS 0.05f
C902 VN.n38 VSUBS 0.095161f
C903 VN.t5 VSUBS 1.91532f
C904 VN.n39 VSUBS 0.826766f
C905 VN.n40 VSUBS 0.03098f
C906 VN.n41 VSUBS 0.06211f
C907 VN.n42 VSUBS 0.03098f
C908 VN.n43 VSUBS 0.057738f
C909 VN.n44 VSUBS 0.03098f
C910 VN.t0 VSUBS 1.91532f
C911 VN.n45 VSUBS 0.057738f
C912 VN.n46 VSUBS 0.03098f
C913 VN.n47 VSUBS 0.057738f
C914 VN.t4 VSUBS 2.36791f
C915 VN.n48 VSUBS 0.798205f
C916 VN.t2 VSUBS 1.91532f
C917 VN.n49 VSUBS 0.823674f
C918 VN.n50 VSUBS 0.05004f
C919 VN.n51 VSUBS 0.400826f
C920 VN.n52 VSUBS 0.03098f
C921 VN.n53 VSUBS 0.03098f
C922 VN.n54 VSUBS 0.057738f
C923 VN.n55 VSUBS 0.045225f
C924 VN.n56 VSUBS 0.045225f
C925 VN.n57 VSUBS 0.03098f
C926 VN.n58 VSUBS 0.03098f
C927 VN.n59 VSUBS 0.03098f
C928 VN.n60 VSUBS 0.057738f
C929 VN.n61 VSUBS 0.05004f
C930 VN.n62 VSUBS 0.704566f
C931 VN.n63 VSUBS 0.036928f
C932 VN.n64 VSUBS 0.03098f
C933 VN.n65 VSUBS 0.03098f
C934 VN.n66 VSUBS 0.03098f
C935 VN.n67 VSUBS 0.057738f
C936 VN.n68 VSUBS 0.060874f
C937 VN.n69 VSUBS 0.025204f
C938 VN.n70 VSUBS 0.03098f
C939 VN.n71 VSUBS 0.03098f
C940 VN.n72 VSUBS 0.03098f
C941 VN.n73 VSUBS 0.057738f
C942 VN.n74 VSUBS 0.057738f
C943 VN.n75 VSUBS 0.034647f
C944 VN.n76 VSUBS 0.05f
C945 VN.n77 VSUBS 1.92527f
C946 VDD1.t4 VSUBS 0.160279f
C947 VDD1.t7 VSUBS 0.160279f
C948 VDD1.n0 VSUBS 1.08419f
C949 VDD1.t0 VSUBS 0.160279f
C950 VDD1.t3 VSUBS 0.160279f
C951 VDD1.n1 VSUBS 1.08257f
C952 VDD1.t5 VSUBS 0.160279f
C953 VDD1.t1 VSUBS 0.160279f
C954 VDD1.n2 VSUBS 1.08257f
C955 VDD1.n3 VSUBS 5.5665f
C956 VDD1.t2 VSUBS 0.160279f
C957 VDD1.t6 VSUBS 0.160279f
C958 VDD1.n4 VSUBS 1.06081f
C959 VDD1.n5 VSUBS 4.29942f
C960 VTAIL.t5 VSUBS 0.147671f
C961 VTAIL.t7 VSUBS 0.147671f
C962 VTAIL.n0 VSUBS 0.866529f
C963 VTAIL.n1 VSUBS 0.947974f
C964 VTAIL.n2 VSUBS 0.034016f
C965 VTAIL.n3 VSUBS 0.031197f
C966 VTAIL.n4 VSUBS 0.016764f
C967 VTAIL.n5 VSUBS 0.039624f
C968 VTAIL.n6 VSUBS 0.01775f
C969 VTAIL.n7 VSUBS 0.031197f
C970 VTAIL.n8 VSUBS 0.016764f
C971 VTAIL.n9 VSUBS 0.039624f
C972 VTAIL.n10 VSUBS 0.01775f
C973 VTAIL.n11 VSUBS 0.137829f
C974 VTAIL.t0 VSUBS 0.085005f
C975 VTAIL.n12 VSUBS 0.029718f
C976 VTAIL.n13 VSUBS 0.025194f
C977 VTAIL.n14 VSUBS 0.016764f
C978 VTAIL.n15 VSUBS 0.714257f
C979 VTAIL.n16 VSUBS 0.031197f
C980 VTAIL.n17 VSUBS 0.016764f
C981 VTAIL.n18 VSUBS 0.01775f
C982 VTAIL.n19 VSUBS 0.039624f
C983 VTAIL.n20 VSUBS 0.039624f
C984 VTAIL.n21 VSUBS 0.01775f
C985 VTAIL.n22 VSUBS 0.016764f
C986 VTAIL.n23 VSUBS 0.031197f
C987 VTAIL.n24 VSUBS 0.031197f
C988 VTAIL.n25 VSUBS 0.016764f
C989 VTAIL.n26 VSUBS 0.01775f
C990 VTAIL.n27 VSUBS 0.039624f
C991 VTAIL.n28 VSUBS 0.09503f
C992 VTAIL.n29 VSUBS 0.01775f
C993 VTAIL.n30 VSUBS 0.016764f
C994 VTAIL.n31 VSUBS 0.071684f
C995 VTAIL.n32 VSUBS 0.047737f
C996 VTAIL.n33 VSUBS 0.440199f
C997 VTAIL.n34 VSUBS 0.034016f
C998 VTAIL.n35 VSUBS 0.031197f
C999 VTAIL.n36 VSUBS 0.016764f
C1000 VTAIL.n37 VSUBS 0.039624f
C1001 VTAIL.n38 VSUBS 0.01775f
C1002 VTAIL.n39 VSUBS 0.031197f
C1003 VTAIL.n40 VSUBS 0.016764f
C1004 VTAIL.n41 VSUBS 0.039624f
C1005 VTAIL.n42 VSUBS 0.01775f
C1006 VTAIL.n43 VSUBS 0.137829f
C1007 VTAIL.t15 VSUBS 0.085005f
C1008 VTAIL.n44 VSUBS 0.029718f
C1009 VTAIL.n45 VSUBS 0.025194f
C1010 VTAIL.n46 VSUBS 0.016764f
C1011 VTAIL.n47 VSUBS 0.714257f
C1012 VTAIL.n48 VSUBS 0.031197f
C1013 VTAIL.n49 VSUBS 0.016764f
C1014 VTAIL.n50 VSUBS 0.01775f
C1015 VTAIL.n51 VSUBS 0.039624f
C1016 VTAIL.n52 VSUBS 0.039624f
C1017 VTAIL.n53 VSUBS 0.01775f
C1018 VTAIL.n54 VSUBS 0.016764f
C1019 VTAIL.n55 VSUBS 0.031197f
C1020 VTAIL.n56 VSUBS 0.031197f
C1021 VTAIL.n57 VSUBS 0.016764f
C1022 VTAIL.n58 VSUBS 0.01775f
C1023 VTAIL.n59 VSUBS 0.039624f
C1024 VTAIL.n60 VSUBS 0.09503f
C1025 VTAIL.n61 VSUBS 0.01775f
C1026 VTAIL.n62 VSUBS 0.016764f
C1027 VTAIL.n63 VSUBS 0.071684f
C1028 VTAIL.n64 VSUBS 0.047737f
C1029 VTAIL.n65 VSUBS 0.440199f
C1030 VTAIL.t11 VSUBS 0.147671f
C1031 VTAIL.t8 VSUBS 0.147671f
C1032 VTAIL.n66 VSUBS 0.866529f
C1033 VTAIL.n67 VSUBS 1.30869f
C1034 VTAIL.n68 VSUBS 0.034016f
C1035 VTAIL.n69 VSUBS 0.031197f
C1036 VTAIL.n70 VSUBS 0.016764f
C1037 VTAIL.n71 VSUBS 0.039624f
C1038 VTAIL.n72 VSUBS 0.01775f
C1039 VTAIL.n73 VSUBS 0.031197f
C1040 VTAIL.n74 VSUBS 0.016764f
C1041 VTAIL.n75 VSUBS 0.039624f
C1042 VTAIL.n76 VSUBS 0.01775f
C1043 VTAIL.n77 VSUBS 0.137829f
C1044 VTAIL.t14 VSUBS 0.085005f
C1045 VTAIL.n78 VSUBS 0.029718f
C1046 VTAIL.n79 VSUBS 0.025194f
C1047 VTAIL.n80 VSUBS 0.016764f
C1048 VTAIL.n81 VSUBS 0.714257f
C1049 VTAIL.n82 VSUBS 0.031197f
C1050 VTAIL.n83 VSUBS 0.016764f
C1051 VTAIL.n84 VSUBS 0.01775f
C1052 VTAIL.n85 VSUBS 0.039624f
C1053 VTAIL.n86 VSUBS 0.039624f
C1054 VTAIL.n87 VSUBS 0.01775f
C1055 VTAIL.n88 VSUBS 0.016764f
C1056 VTAIL.n89 VSUBS 0.031197f
C1057 VTAIL.n90 VSUBS 0.031197f
C1058 VTAIL.n91 VSUBS 0.016764f
C1059 VTAIL.n92 VSUBS 0.01775f
C1060 VTAIL.n93 VSUBS 0.039624f
C1061 VTAIL.n94 VSUBS 0.09503f
C1062 VTAIL.n95 VSUBS 0.01775f
C1063 VTAIL.n96 VSUBS 0.016764f
C1064 VTAIL.n97 VSUBS 0.071684f
C1065 VTAIL.n98 VSUBS 0.047737f
C1066 VTAIL.n99 VSUBS 1.7024f
C1067 VTAIL.n100 VSUBS 0.034016f
C1068 VTAIL.n101 VSUBS 0.031197f
C1069 VTAIL.n102 VSUBS 0.016764f
C1070 VTAIL.n103 VSUBS 0.039624f
C1071 VTAIL.n104 VSUBS 0.01775f
C1072 VTAIL.n105 VSUBS 0.031197f
C1073 VTAIL.n106 VSUBS 0.016764f
C1074 VTAIL.n107 VSUBS 0.039624f
C1075 VTAIL.n108 VSUBS 0.01775f
C1076 VTAIL.n109 VSUBS 0.137829f
C1077 VTAIL.t4 VSUBS 0.085005f
C1078 VTAIL.n110 VSUBS 0.029718f
C1079 VTAIL.n111 VSUBS 0.025194f
C1080 VTAIL.n112 VSUBS 0.016764f
C1081 VTAIL.n113 VSUBS 0.714256f
C1082 VTAIL.n114 VSUBS 0.031197f
C1083 VTAIL.n115 VSUBS 0.016764f
C1084 VTAIL.n116 VSUBS 0.01775f
C1085 VTAIL.n117 VSUBS 0.039624f
C1086 VTAIL.n118 VSUBS 0.039624f
C1087 VTAIL.n119 VSUBS 0.01775f
C1088 VTAIL.n120 VSUBS 0.016764f
C1089 VTAIL.n121 VSUBS 0.031197f
C1090 VTAIL.n122 VSUBS 0.031197f
C1091 VTAIL.n123 VSUBS 0.016764f
C1092 VTAIL.n124 VSUBS 0.01775f
C1093 VTAIL.n125 VSUBS 0.039624f
C1094 VTAIL.n126 VSUBS 0.09503f
C1095 VTAIL.n127 VSUBS 0.01775f
C1096 VTAIL.n128 VSUBS 0.016764f
C1097 VTAIL.n129 VSUBS 0.071684f
C1098 VTAIL.n130 VSUBS 0.047737f
C1099 VTAIL.n131 VSUBS 1.7024f
C1100 VTAIL.t2 VSUBS 0.147671f
C1101 VTAIL.t6 VSUBS 0.147671f
C1102 VTAIL.n132 VSUBS 0.866536f
C1103 VTAIL.n133 VSUBS 1.30868f
C1104 VTAIL.n134 VSUBS 0.034016f
C1105 VTAIL.n135 VSUBS 0.031197f
C1106 VTAIL.n136 VSUBS 0.016764f
C1107 VTAIL.n137 VSUBS 0.039624f
C1108 VTAIL.n138 VSUBS 0.01775f
C1109 VTAIL.n139 VSUBS 0.031197f
C1110 VTAIL.n140 VSUBS 0.016764f
C1111 VTAIL.n141 VSUBS 0.039624f
C1112 VTAIL.n142 VSUBS 0.01775f
C1113 VTAIL.n143 VSUBS 0.137829f
C1114 VTAIL.t1 VSUBS 0.085005f
C1115 VTAIL.n144 VSUBS 0.029718f
C1116 VTAIL.n145 VSUBS 0.025194f
C1117 VTAIL.n146 VSUBS 0.016764f
C1118 VTAIL.n147 VSUBS 0.714256f
C1119 VTAIL.n148 VSUBS 0.031197f
C1120 VTAIL.n149 VSUBS 0.016764f
C1121 VTAIL.n150 VSUBS 0.01775f
C1122 VTAIL.n151 VSUBS 0.039624f
C1123 VTAIL.n152 VSUBS 0.039624f
C1124 VTAIL.n153 VSUBS 0.01775f
C1125 VTAIL.n154 VSUBS 0.016764f
C1126 VTAIL.n155 VSUBS 0.031197f
C1127 VTAIL.n156 VSUBS 0.031197f
C1128 VTAIL.n157 VSUBS 0.016764f
C1129 VTAIL.n158 VSUBS 0.01775f
C1130 VTAIL.n159 VSUBS 0.039624f
C1131 VTAIL.n160 VSUBS 0.09503f
C1132 VTAIL.n161 VSUBS 0.01775f
C1133 VTAIL.n162 VSUBS 0.016764f
C1134 VTAIL.n163 VSUBS 0.071684f
C1135 VTAIL.n164 VSUBS 0.047737f
C1136 VTAIL.n165 VSUBS 0.440199f
C1137 VTAIL.n166 VSUBS 0.034016f
C1138 VTAIL.n167 VSUBS 0.031197f
C1139 VTAIL.n168 VSUBS 0.016764f
C1140 VTAIL.n169 VSUBS 0.039624f
C1141 VTAIL.n170 VSUBS 0.01775f
C1142 VTAIL.n171 VSUBS 0.031197f
C1143 VTAIL.n172 VSUBS 0.016764f
C1144 VTAIL.n173 VSUBS 0.039624f
C1145 VTAIL.n174 VSUBS 0.01775f
C1146 VTAIL.n175 VSUBS 0.137829f
C1147 VTAIL.t10 VSUBS 0.085005f
C1148 VTAIL.n176 VSUBS 0.029718f
C1149 VTAIL.n177 VSUBS 0.025194f
C1150 VTAIL.n178 VSUBS 0.016764f
C1151 VTAIL.n179 VSUBS 0.714256f
C1152 VTAIL.n180 VSUBS 0.031197f
C1153 VTAIL.n181 VSUBS 0.016764f
C1154 VTAIL.n182 VSUBS 0.01775f
C1155 VTAIL.n183 VSUBS 0.039624f
C1156 VTAIL.n184 VSUBS 0.039624f
C1157 VTAIL.n185 VSUBS 0.01775f
C1158 VTAIL.n186 VSUBS 0.016764f
C1159 VTAIL.n187 VSUBS 0.031197f
C1160 VTAIL.n188 VSUBS 0.031197f
C1161 VTAIL.n189 VSUBS 0.016764f
C1162 VTAIL.n190 VSUBS 0.01775f
C1163 VTAIL.n191 VSUBS 0.039624f
C1164 VTAIL.n192 VSUBS 0.09503f
C1165 VTAIL.n193 VSUBS 0.01775f
C1166 VTAIL.n194 VSUBS 0.016764f
C1167 VTAIL.n195 VSUBS 0.071684f
C1168 VTAIL.n196 VSUBS 0.047737f
C1169 VTAIL.n197 VSUBS 0.440199f
C1170 VTAIL.t12 VSUBS 0.147671f
C1171 VTAIL.t13 VSUBS 0.147671f
C1172 VTAIL.n198 VSUBS 0.866536f
C1173 VTAIL.n199 VSUBS 1.30868f
C1174 VTAIL.n200 VSUBS 0.034016f
C1175 VTAIL.n201 VSUBS 0.031197f
C1176 VTAIL.n202 VSUBS 0.016764f
C1177 VTAIL.n203 VSUBS 0.039624f
C1178 VTAIL.n204 VSUBS 0.01775f
C1179 VTAIL.n205 VSUBS 0.031197f
C1180 VTAIL.n206 VSUBS 0.016764f
C1181 VTAIL.n207 VSUBS 0.039624f
C1182 VTAIL.n208 VSUBS 0.01775f
C1183 VTAIL.n209 VSUBS 0.137829f
C1184 VTAIL.t9 VSUBS 0.085005f
C1185 VTAIL.n210 VSUBS 0.029718f
C1186 VTAIL.n211 VSUBS 0.025194f
C1187 VTAIL.n212 VSUBS 0.016764f
C1188 VTAIL.n213 VSUBS 0.714256f
C1189 VTAIL.n214 VSUBS 0.031197f
C1190 VTAIL.n215 VSUBS 0.016764f
C1191 VTAIL.n216 VSUBS 0.01775f
C1192 VTAIL.n217 VSUBS 0.039624f
C1193 VTAIL.n218 VSUBS 0.039624f
C1194 VTAIL.n219 VSUBS 0.01775f
C1195 VTAIL.n220 VSUBS 0.016764f
C1196 VTAIL.n221 VSUBS 0.031197f
C1197 VTAIL.n222 VSUBS 0.031197f
C1198 VTAIL.n223 VSUBS 0.016764f
C1199 VTAIL.n224 VSUBS 0.01775f
C1200 VTAIL.n225 VSUBS 0.039624f
C1201 VTAIL.n226 VSUBS 0.09503f
C1202 VTAIL.n227 VSUBS 0.01775f
C1203 VTAIL.n228 VSUBS 0.016764f
C1204 VTAIL.n229 VSUBS 0.071684f
C1205 VTAIL.n230 VSUBS 0.047737f
C1206 VTAIL.n231 VSUBS 1.7024f
C1207 VTAIL.n232 VSUBS 0.034016f
C1208 VTAIL.n233 VSUBS 0.031197f
C1209 VTAIL.n234 VSUBS 0.016764f
C1210 VTAIL.n235 VSUBS 0.039624f
C1211 VTAIL.n236 VSUBS 0.01775f
C1212 VTAIL.n237 VSUBS 0.031197f
C1213 VTAIL.n238 VSUBS 0.016764f
C1214 VTAIL.n239 VSUBS 0.039624f
C1215 VTAIL.n240 VSUBS 0.01775f
C1216 VTAIL.n241 VSUBS 0.137829f
C1217 VTAIL.t3 VSUBS 0.085005f
C1218 VTAIL.n242 VSUBS 0.029718f
C1219 VTAIL.n243 VSUBS 0.025194f
C1220 VTAIL.n244 VSUBS 0.016764f
C1221 VTAIL.n245 VSUBS 0.714257f
C1222 VTAIL.n246 VSUBS 0.031197f
C1223 VTAIL.n247 VSUBS 0.016764f
C1224 VTAIL.n248 VSUBS 0.01775f
C1225 VTAIL.n249 VSUBS 0.039624f
C1226 VTAIL.n250 VSUBS 0.039624f
C1227 VTAIL.n251 VSUBS 0.01775f
C1228 VTAIL.n252 VSUBS 0.016764f
C1229 VTAIL.n253 VSUBS 0.031197f
C1230 VTAIL.n254 VSUBS 0.031197f
C1231 VTAIL.n255 VSUBS 0.016764f
C1232 VTAIL.n256 VSUBS 0.01775f
C1233 VTAIL.n257 VSUBS 0.039624f
C1234 VTAIL.n258 VSUBS 0.09503f
C1235 VTAIL.n259 VSUBS 0.01775f
C1236 VTAIL.n260 VSUBS 0.016764f
C1237 VTAIL.n261 VSUBS 0.071684f
C1238 VTAIL.n262 VSUBS 0.047737f
C1239 VTAIL.n263 VSUBS 1.69655f
C1240 VP.t6 VSUBS 2.16746f
C1241 VP.n0 VSUBS 0.935604f
C1242 VP.n1 VSUBS 0.035058f
C1243 VP.n2 VSUBS 0.070286f
C1244 VP.n3 VSUBS 0.035058f
C1245 VP.n4 VSUBS 0.065339f
C1246 VP.n5 VSUBS 0.035058f
C1247 VP.t2 VSUBS 2.16746f
C1248 VP.n6 VSUBS 0.065339f
C1249 VP.n7 VSUBS 0.035058f
C1250 VP.n8 VSUBS 0.065339f
C1251 VP.n9 VSUBS 0.035058f
C1252 VP.t4 VSUBS 2.16746f
C1253 VP.n10 VSUBS 0.065339f
C1254 VP.n11 VSUBS 0.035058f
C1255 VP.n12 VSUBS 0.065339f
C1256 VP.n13 VSUBS 0.056583f
C1257 VP.t7 VSUBS 2.16746f
C1258 VP.t1 VSUBS 2.16746f
C1259 VP.n14 VSUBS 0.935604f
C1260 VP.n15 VSUBS 0.035058f
C1261 VP.n16 VSUBS 0.070286f
C1262 VP.n17 VSUBS 0.035058f
C1263 VP.n18 VSUBS 0.065339f
C1264 VP.n19 VSUBS 0.035058f
C1265 VP.t5 VSUBS 2.16746f
C1266 VP.n20 VSUBS 0.065339f
C1267 VP.n21 VSUBS 0.035058f
C1268 VP.n22 VSUBS 0.065339f
C1269 VP.t3 VSUBS 2.67962f
C1270 VP.n23 VSUBS 0.903284f
C1271 VP.t0 VSUBS 2.16746f
C1272 VP.n24 VSUBS 0.932104f
C1273 VP.n25 VSUBS 0.056628f
C1274 VP.n26 VSUBS 0.453592f
C1275 VP.n27 VSUBS 0.035058f
C1276 VP.n28 VSUBS 0.035058f
C1277 VP.n29 VSUBS 0.065339f
C1278 VP.n30 VSUBS 0.051178f
C1279 VP.n31 VSUBS 0.051178f
C1280 VP.n32 VSUBS 0.035058f
C1281 VP.n33 VSUBS 0.035058f
C1282 VP.n34 VSUBS 0.035058f
C1283 VP.n35 VSUBS 0.065339f
C1284 VP.n36 VSUBS 0.056628f
C1285 VP.n37 VSUBS 0.797317f
C1286 VP.n38 VSUBS 0.041789f
C1287 VP.n39 VSUBS 0.035058f
C1288 VP.n40 VSUBS 0.035058f
C1289 VP.n41 VSUBS 0.035058f
C1290 VP.n42 VSUBS 0.065339f
C1291 VP.n43 VSUBS 0.068888f
C1292 VP.n44 VSUBS 0.028522f
C1293 VP.n45 VSUBS 0.035058f
C1294 VP.n46 VSUBS 0.035058f
C1295 VP.n47 VSUBS 0.035058f
C1296 VP.n48 VSUBS 0.065339f
C1297 VP.n49 VSUBS 0.065339f
C1298 VP.n50 VSUBS 0.039208f
C1299 VP.n51 VSUBS 0.056583f
C1300 VP.n52 VSUBS 2.16462f
C1301 VP.n53 VSUBS 2.18861f
C1302 VP.n54 VSUBS 0.935604f
C1303 VP.n55 VSUBS 0.039208f
C1304 VP.n56 VSUBS 0.065339f
C1305 VP.n57 VSUBS 0.035058f
C1306 VP.n58 VSUBS 0.035058f
C1307 VP.n59 VSUBS 0.035058f
C1308 VP.n60 VSUBS 0.070286f
C1309 VP.n61 VSUBS 0.028522f
C1310 VP.n62 VSUBS 0.068888f
C1311 VP.n63 VSUBS 0.035058f
C1312 VP.n64 VSUBS 0.035058f
C1313 VP.n65 VSUBS 0.035058f
C1314 VP.n66 VSUBS 0.065339f
C1315 VP.n67 VSUBS 0.041789f
C1316 VP.n68 VSUBS 0.797317f
C1317 VP.n69 VSUBS 0.056628f
C1318 VP.n70 VSUBS 0.035058f
C1319 VP.n71 VSUBS 0.035058f
C1320 VP.n72 VSUBS 0.035058f
C1321 VP.n73 VSUBS 0.065339f
C1322 VP.n74 VSUBS 0.051178f
C1323 VP.n75 VSUBS 0.051178f
C1324 VP.n76 VSUBS 0.035058f
C1325 VP.n77 VSUBS 0.035058f
C1326 VP.n78 VSUBS 0.035058f
C1327 VP.n79 VSUBS 0.065339f
C1328 VP.n80 VSUBS 0.056628f
C1329 VP.n81 VSUBS 0.797317f
C1330 VP.n82 VSUBS 0.041789f
C1331 VP.n83 VSUBS 0.035058f
C1332 VP.n84 VSUBS 0.035058f
C1333 VP.n85 VSUBS 0.035058f
C1334 VP.n86 VSUBS 0.065339f
C1335 VP.n87 VSUBS 0.068888f
C1336 VP.n88 VSUBS 0.028522f
C1337 VP.n89 VSUBS 0.035058f
C1338 VP.n90 VSUBS 0.035058f
C1339 VP.n91 VSUBS 0.035058f
C1340 VP.n92 VSUBS 0.065339f
C1341 VP.n93 VSUBS 0.065339f
C1342 VP.n94 VSUBS 0.039208f
C1343 VP.n95 VSUBS 0.056583f
C1344 VP.n96 VSUBS 0.107688f
.ends

