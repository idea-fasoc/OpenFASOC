* NGSPICE file created from diff_pair_sample_1133.ext - technology: sky130A

.subckt diff_pair_sample_1133 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t9 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=0 ps=0 w=19.48 l=3.54
X1 VTAIL.t7 VN.t0 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=3.2142 ps=19.81 w=19.48 l=3.54
X2 B.t14 B.t12 B.t13 B.t5 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=0 ps=0 w=19.48 l=3.54
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=0 ps=0 w=19.48 l=3.54
X4 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=0 ps=0 w=19.48 l=3.54
X5 VDD2.t3 VN.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2142 pd=19.81 as=7.5972 ps=39.74 w=19.48 l=3.54
X6 VTAIL.t5 VN.t2 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=3.2142 ps=19.81 w=19.48 l=3.54
X7 VDD2.t2 VN.t3 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2142 pd=19.81 as=7.5972 ps=39.74 w=19.48 l=3.54
X8 VTAIL.t3 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=3.2142 ps=19.81 w=19.48 l=3.54
X9 VDD1.t2 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=3.2142 pd=19.81 as=7.5972 ps=39.74 w=19.48 l=3.54
X10 VTAIL.t0 VP.t2 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=7.5972 pd=39.74 as=3.2142 ps=19.81 w=19.48 l=3.54
X11 VDD1.t0 VP.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=3.2142 pd=19.81 as=7.5972 ps=39.74 w=19.48 l=3.54
R0 B.n761 B.n151 585
R1 B.n151 B.n78 585
R2 B.n763 B.n762 585
R3 B.n765 B.n150 585
R4 B.n768 B.n767 585
R5 B.n769 B.n149 585
R6 B.n771 B.n770 585
R7 B.n773 B.n148 585
R8 B.n776 B.n775 585
R9 B.n777 B.n147 585
R10 B.n779 B.n778 585
R11 B.n781 B.n146 585
R12 B.n784 B.n783 585
R13 B.n785 B.n145 585
R14 B.n787 B.n786 585
R15 B.n789 B.n144 585
R16 B.n792 B.n791 585
R17 B.n793 B.n143 585
R18 B.n795 B.n794 585
R19 B.n797 B.n142 585
R20 B.n800 B.n799 585
R21 B.n801 B.n141 585
R22 B.n803 B.n802 585
R23 B.n805 B.n140 585
R24 B.n808 B.n807 585
R25 B.n809 B.n139 585
R26 B.n811 B.n810 585
R27 B.n813 B.n138 585
R28 B.n816 B.n815 585
R29 B.n817 B.n137 585
R30 B.n819 B.n818 585
R31 B.n821 B.n136 585
R32 B.n824 B.n823 585
R33 B.n825 B.n135 585
R34 B.n827 B.n826 585
R35 B.n829 B.n134 585
R36 B.n832 B.n831 585
R37 B.n833 B.n133 585
R38 B.n835 B.n834 585
R39 B.n837 B.n132 585
R40 B.n840 B.n839 585
R41 B.n841 B.n131 585
R42 B.n843 B.n842 585
R43 B.n845 B.n130 585
R44 B.n848 B.n847 585
R45 B.n849 B.n129 585
R46 B.n851 B.n850 585
R47 B.n853 B.n128 585
R48 B.n856 B.n855 585
R49 B.n857 B.n127 585
R50 B.n859 B.n858 585
R51 B.n861 B.n126 585
R52 B.n864 B.n863 585
R53 B.n865 B.n125 585
R54 B.n867 B.n866 585
R55 B.n869 B.n124 585
R56 B.n872 B.n871 585
R57 B.n873 B.n123 585
R58 B.n875 B.n874 585
R59 B.n877 B.n122 585
R60 B.n880 B.n879 585
R61 B.n881 B.n121 585
R62 B.n883 B.n882 585
R63 B.n885 B.n120 585
R64 B.n888 B.n887 585
R65 B.n890 B.n117 585
R66 B.n892 B.n891 585
R67 B.n894 B.n116 585
R68 B.n897 B.n896 585
R69 B.n898 B.n115 585
R70 B.n900 B.n899 585
R71 B.n902 B.n114 585
R72 B.n905 B.n904 585
R73 B.n906 B.n111 585
R74 B.n909 B.n908 585
R75 B.n911 B.n110 585
R76 B.n914 B.n913 585
R77 B.n915 B.n109 585
R78 B.n917 B.n916 585
R79 B.n919 B.n108 585
R80 B.n922 B.n921 585
R81 B.n923 B.n107 585
R82 B.n925 B.n924 585
R83 B.n927 B.n106 585
R84 B.n930 B.n929 585
R85 B.n931 B.n105 585
R86 B.n933 B.n932 585
R87 B.n935 B.n104 585
R88 B.n938 B.n937 585
R89 B.n939 B.n103 585
R90 B.n941 B.n940 585
R91 B.n943 B.n102 585
R92 B.n946 B.n945 585
R93 B.n947 B.n101 585
R94 B.n949 B.n948 585
R95 B.n951 B.n100 585
R96 B.n954 B.n953 585
R97 B.n955 B.n99 585
R98 B.n957 B.n956 585
R99 B.n959 B.n98 585
R100 B.n962 B.n961 585
R101 B.n963 B.n97 585
R102 B.n965 B.n964 585
R103 B.n967 B.n96 585
R104 B.n970 B.n969 585
R105 B.n971 B.n95 585
R106 B.n973 B.n972 585
R107 B.n975 B.n94 585
R108 B.n978 B.n977 585
R109 B.n979 B.n93 585
R110 B.n981 B.n980 585
R111 B.n983 B.n92 585
R112 B.n986 B.n985 585
R113 B.n987 B.n91 585
R114 B.n989 B.n988 585
R115 B.n991 B.n90 585
R116 B.n994 B.n993 585
R117 B.n995 B.n89 585
R118 B.n997 B.n996 585
R119 B.n999 B.n88 585
R120 B.n1002 B.n1001 585
R121 B.n1003 B.n87 585
R122 B.n1005 B.n1004 585
R123 B.n1007 B.n86 585
R124 B.n1010 B.n1009 585
R125 B.n1011 B.n85 585
R126 B.n1013 B.n1012 585
R127 B.n1015 B.n84 585
R128 B.n1018 B.n1017 585
R129 B.n1019 B.n83 585
R130 B.n1021 B.n1020 585
R131 B.n1023 B.n82 585
R132 B.n1026 B.n1025 585
R133 B.n1027 B.n81 585
R134 B.n1029 B.n1028 585
R135 B.n1031 B.n80 585
R136 B.n1034 B.n1033 585
R137 B.n1035 B.n79 585
R138 B.n760 B.n77 585
R139 B.n1038 B.n77 585
R140 B.n759 B.n76 585
R141 B.n1039 B.n76 585
R142 B.n758 B.n75 585
R143 B.n1040 B.n75 585
R144 B.n757 B.n756 585
R145 B.n756 B.n71 585
R146 B.n755 B.n70 585
R147 B.n1046 B.n70 585
R148 B.n754 B.n69 585
R149 B.n1047 B.n69 585
R150 B.n753 B.n68 585
R151 B.n1048 B.n68 585
R152 B.n752 B.n751 585
R153 B.n751 B.n64 585
R154 B.n750 B.n63 585
R155 B.n1054 B.n63 585
R156 B.n749 B.n62 585
R157 B.n1055 B.n62 585
R158 B.n748 B.n61 585
R159 B.n1056 B.n61 585
R160 B.n747 B.n746 585
R161 B.n746 B.n57 585
R162 B.n745 B.n56 585
R163 B.n1062 B.n56 585
R164 B.n744 B.n55 585
R165 B.n1063 B.n55 585
R166 B.n743 B.n54 585
R167 B.n1064 B.n54 585
R168 B.n742 B.n741 585
R169 B.n741 B.n50 585
R170 B.n740 B.n49 585
R171 B.n1070 B.n49 585
R172 B.n739 B.n48 585
R173 B.n1071 B.n48 585
R174 B.n738 B.n47 585
R175 B.n1072 B.n47 585
R176 B.n737 B.n736 585
R177 B.n736 B.n43 585
R178 B.n735 B.n42 585
R179 B.n1078 B.n42 585
R180 B.n734 B.n41 585
R181 B.n1079 B.n41 585
R182 B.n733 B.n40 585
R183 B.n1080 B.n40 585
R184 B.n732 B.n731 585
R185 B.n731 B.n39 585
R186 B.n730 B.n35 585
R187 B.n1086 B.n35 585
R188 B.n729 B.n34 585
R189 B.n1087 B.n34 585
R190 B.n728 B.n33 585
R191 B.n1088 B.n33 585
R192 B.n727 B.n726 585
R193 B.n726 B.n29 585
R194 B.n725 B.n28 585
R195 B.n1094 B.n28 585
R196 B.n724 B.n27 585
R197 B.n1095 B.n27 585
R198 B.n723 B.n26 585
R199 B.n1096 B.n26 585
R200 B.n722 B.n721 585
R201 B.n721 B.n22 585
R202 B.n720 B.n21 585
R203 B.n1102 B.n21 585
R204 B.n719 B.n20 585
R205 B.n1103 B.n20 585
R206 B.n718 B.n19 585
R207 B.n1104 B.n19 585
R208 B.n717 B.n716 585
R209 B.n716 B.n15 585
R210 B.n715 B.n14 585
R211 B.n1110 B.n14 585
R212 B.n714 B.n13 585
R213 B.n1111 B.n13 585
R214 B.n713 B.n12 585
R215 B.n1112 B.n12 585
R216 B.n712 B.n711 585
R217 B.n711 B.n8 585
R218 B.n710 B.n7 585
R219 B.n1118 B.n7 585
R220 B.n709 B.n6 585
R221 B.n1119 B.n6 585
R222 B.n708 B.n5 585
R223 B.n1120 B.n5 585
R224 B.n707 B.n706 585
R225 B.n706 B.n4 585
R226 B.n705 B.n152 585
R227 B.n705 B.n704 585
R228 B.n695 B.n153 585
R229 B.n154 B.n153 585
R230 B.n697 B.n696 585
R231 B.n698 B.n697 585
R232 B.n694 B.n159 585
R233 B.n159 B.n158 585
R234 B.n693 B.n692 585
R235 B.n692 B.n691 585
R236 B.n161 B.n160 585
R237 B.n162 B.n161 585
R238 B.n684 B.n683 585
R239 B.n685 B.n684 585
R240 B.n682 B.n167 585
R241 B.n167 B.n166 585
R242 B.n681 B.n680 585
R243 B.n680 B.n679 585
R244 B.n169 B.n168 585
R245 B.n170 B.n169 585
R246 B.n672 B.n671 585
R247 B.n673 B.n672 585
R248 B.n670 B.n175 585
R249 B.n175 B.n174 585
R250 B.n669 B.n668 585
R251 B.n668 B.n667 585
R252 B.n177 B.n176 585
R253 B.n178 B.n177 585
R254 B.n660 B.n659 585
R255 B.n661 B.n660 585
R256 B.n658 B.n183 585
R257 B.n183 B.n182 585
R258 B.n657 B.n656 585
R259 B.n656 B.n655 585
R260 B.n185 B.n184 585
R261 B.n648 B.n185 585
R262 B.n647 B.n646 585
R263 B.n649 B.n647 585
R264 B.n645 B.n190 585
R265 B.n190 B.n189 585
R266 B.n644 B.n643 585
R267 B.n643 B.n642 585
R268 B.n192 B.n191 585
R269 B.n193 B.n192 585
R270 B.n635 B.n634 585
R271 B.n636 B.n635 585
R272 B.n633 B.n198 585
R273 B.n198 B.n197 585
R274 B.n632 B.n631 585
R275 B.n631 B.n630 585
R276 B.n200 B.n199 585
R277 B.n201 B.n200 585
R278 B.n623 B.n622 585
R279 B.n624 B.n623 585
R280 B.n621 B.n206 585
R281 B.n206 B.n205 585
R282 B.n620 B.n619 585
R283 B.n619 B.n618 585
R284 B.n208 B.n207 585
R285 B.n209 B.n208 585
R286 B.n611 B.n610 585
R287 B.n612 B.n611 585
R288 B.n609 B.n214 585
R289 B.n214 B.n213 585
R290 B.n608 B.n607 585
R291 B.n607 B.n606 585
R292 B.n216 B.n215 585
R293 B.n217 B.n216 585
R294 B.n599 B.n598 585
R295 B.n600 B.n599 585
R296 B.n597 B.n222 585
R297 B.n222 B.n221 585
R298 B.n596 B.n595 585
R299 B.n595 B.n594 585
R300 B.n224 B.n223 585
R301 B.n225 B.n224 585
R302 B.n587 B.n586 585
R303 B.n588 B.n587 585
R304 B.n585 B.n230 585
R305 B.n230 B.n229 585
R306 B.n584 B.n583 585
R307 B.n583 B.n582 585
R308 B.n579 B.n234 585
R309 B.n578 B.n577 585
R310 B.n575 B.n235 585
R311 B.n575 B.n233 585
R312 B.n574 B.n573 585
R313 B.n572 B.n571 585
R314 B.n570 B.n237 585
R315 B.n568 B.n567 585
R316 B.n566 B.n238 585
R317 B.n565 B.n564 585
R318 B.n562 B.n239 585
R319 B.n560 B.n559 585
R320 B.n558 B.n240 585
R321 B.n557 B.n556 585
R322 B.n554 B.n241 585
R323 B.n552 B.n551 585
R324 B.n550 B.n242 585
R325 B.n549 B.n548 585
R326 B.n546 B.n243 585
R327 B.n544 B.n543 585
R328 B.n542 B.n244 585
R329 B.n541 B.n540 585
R330 B.n538 B.n245 585
R331 B.n536 B.n535 585
R332 B.n534 B.n246 585
R333 B.n533 B.n532 585
R334 B.n530 B.n247 585
R335 B.n528 B.n527 585
R336 B.n526 B.n248 585
R337 B.n525 B.n524 585
R338 B.n522 B.n249 585
R339 B.n520 B.n519 585
R340 B.n518 B.n250 585
R341 B.n517 B.n516 585
R342 B.n514 B.n251 585
R343 B.n512 B.n511 585
R344 B.n510 B.n252 585
R345 B.n509 B.n508 585
R346 B.n506 B.n253 585
R347 B.n504 B.n503 585
R348 B.n502 B.n254 585
R349 B.n501 B.n500 585
R350 B.n498 B.n255 585
R351 B.n496 B.n495 585
R352 B.n494 B.n256 585
R353 B.n493 B.n492 585
R354 B.n490 B.n257 585
R355 B.n488 B.n487 585
R356 B.n486 B.n258 585
R357 B.n485 B.n484 585
R358 B.n482 B.n259 585
R359 B.n480 B.n479 585
R360 B.n478 B.n260 585
R361 B.n477 B.n476 585
R362 B.n474 B.n261 585
R363 B.n472 B.n471 585
R364 B.n470 B.n262 585
R365 B.n469 B.n468 585
R366 B.n466 B.n263 585
R367 B.n464 B.n463 585
R368 B.n462 B.n264 585
R369 B.n461 B.n460 585
R370 B.n458 B.n265 585
R371 B.n456 B.n455 585
R372 B.n454 B.n266 585
R373 B.n452 B.n451 585
R374 B.n449 B.n269 585
R375 B.n447 B.n446 585
R376 B.n445 B.n270 585
R377 B.n444 B.n443 585
R378 B.n441 B.n271 585
R379 B.n439 B.n438 585
R380 B.n437 B.n272 585
R381 B.n436 B.n435 585
R382 B.n433 B.n432 585
R383 B.n431 B.n430 585
R384 B.n429 B.n277 585
R385 B.n427 B.n426 585
R386 B.n425 B.n278 585
R387 B.n424 B.n423 585
R388 B.n421 B.n279 585
R389 B.n419 B.n418 585
R390 B.n417 B.n280 585
R391 B.n416 B.n415 585
R392 B.n413 B.n281 585
R393 B.n411 B.n410 585
R394 B.n409 B.n282 585
R395 B.n408 B.n407 585
R396 B.n405 B.n283 585
R397 B.n403 B.n402 585
R398 B.n401 B.n284 585
R399 B.n400 B.n399 585
R400 B.n397 B.n285 585
R401 B.n395 B.n394 585
R402 B.n393 B.n286 585
R403 B.n392 B.n391 585
R404 B.n389 B.n287 585
R405 B.n387 B.n386 585
R406 B.n385 B.n288 585
R407 B.n384 B.n383 585
R408 B.n381 B.n289 585
R409 B.n379 B.n378 585
R410 B.n377 B.n290 585
R411 B.n376 B.n375 585
R412 B.n373 B.n291 585
R413 B.n371 B.n370 585
R414 B.n369 B.n292 585
R415 B.n368 B.n367 585
R416 B.n365 B.n293 585
R417 B.n363 B.n362 585
R418 B.n361 B.n294 585
R419 B.n360 B.n359 585
R420 B.n357 B.n295 585
R421 B.n355 B.n354 585
R422 B.n353 B.n296 585
R423 B.n352 B.n351 585
R424 B.n349 B.n297 585
R425 B.n347 B.n346 585
R426 B.n345 B.n298 585
R427 B.n344 B.n343 585
R428 B.n341 B.n299 585
R429 B.n339 B.n338 585
R430 B.n337 B.n300 585
R431 B.n336 B.n335 585
R432 B.n333 B.n301 585
R433 B.n331 B.n330 585
R434 B.n329 B.n302 585
R435 B.n328 B.n327 585
R436 B.n325 B.n303 585
R437 B.n323 B.n322 585
R438 B.n321 B.n304 585
R439 B.n320 B.n319 585
R440 B.n317 B.n305 585
R441 B.n315 B.n314 585
R442 B.n313 B.n306 585
R443 B.n312 B.n311 585
R444 B.n309 B.n307 585
R445 B.n232 B.n231 585
R446 B.n581 B.n580 585
R447 B.n582 B.n581 585
R448 B.n228 B.n227 585
R449 B.n229 B.n228 585
R450 B.n590 B.n589 585
R451 B.n589 B.n588 585
R452 B.n591 B.n226 585
R453 B.n226 B.n225 585
R454 B.n593 B.n592 585
R455 B.n594 B.n593 585
R456 B.n220 B.n219 585
R457 B.n221 B.n220 585
R458 B.n602 B.n601 585
R459 B.n601 B.n600 585
R460 B.n603 B.n218 585
R461 B.n218 B.n217 585
R462 B.n605 B.n604 585
R463 B.n606 B.n605 585
R464 B.n212 B.n211 585
R465 B.n213 B.n212 585
R466 B.n614 B.n613 585
R467 B.n613 B.n612 585
R468 B.n615 B.n210 585
R469 B.n210 B.n209 585
R470 B.n617 B.n616 585
R471 B.n618 B.n617 585
R472 B.n204 B.n203 585
R473 B.n205 B.n204 585
R474 B.n626 B.n625 585
R475 B.n625 B.n624 585
R476 B.n627 B.n202 585
R477 B.n202 B.n201 585
R478 B.n629 B.n628 585
R479 B.n630 B.n629 585
R480 B.n196 B.n195 585
R481 B.n197 B.n196 585
R482 B.n638 B.n637 585
R483 B.n637 B.n636 585
R484 B.n639 B.n194 585
R485 B.n194 B.n193 585
R486 B.n641 B.n640 585
R487 B.n642 B.n641 585
R488 B.n188 B.n187 585
R489 B.n189 B.n188 585
R490 B.n651 B.n650 585
R491 B.n650 B.n649 585
R492 B.n652 B.n186 585
R493 B.n648 B.n186 585
R494 B.n654 B.n653 585
R495 B.n655 B.n654 585
R496 B.n181 B.n180 585
R497 B.n182 B.n181 585
R498 B.n663 B.n662 585
R499 B.n662 B.n661 585
R500 B.n664 B.n179 585
R501 B.n179 B.n178 585
R502 B.n666 B.n665 585
R503 B.n667 B.n666 585
R504 B.n173 B.n172 585
R505 B.n174 B.n173 585
R506 B.n675 B.n674 585
R507 B.n674 B.n673 585
R508 B.n676 B.n171 585
R509 B.n171 B.n170 585
R510 B.n678 B.n677 585
R511 B.n679 B.n678 585
R512 B.n165 B.n164 585
R513 B.n166 B.n165 585
R514 B.n687 B.n686 585
R515 B.n686 B.n685 585
R516 B.n688 B.n163 585
R517 B.n163 B.n162 585
R518 B.n690 B.n689 585
R519 B.n691 B.n690 585
R520 B.n157 B.n156 585
R521 B.n158 B.n157 585
R522 B.n700 B.n699 585
R523 B.n699 B.n698 585
R524 B.n701 B.n155 585
R525 B.n155 B.n154 585
R526 B.n703 B.n702 585
R527 B.n704 B.n703 585
R528 B.n2 B.n0 585
R529 B.n4 B.n2 585
R530 B.n3 B.n1 585
R531 B.n1119 B.n3 585
R532 B.n1117 B.n1116 585
R533 B.n1118 B.n1117 585
R534 B.n1115 B.n9 585
R535 B.n9 B.n8 585
R536 B.n1114 B.n1113 585
R537 B.n1113 B.n1112 585
R538 B.n11 B.n10 585
R539 B.n1111 B.n11 585
R540 B.n1109 B.n1108 585
R541 B.n1110 B.n1109 585
R542 B.n1107 B.n16 585
R543 B.n16 B.n15 585
R544 B.n1106 B.n1105 585
R545 B.n1105 B.n1104 585
R546 B.n18 B.n17 585
R547 B.n1103 B.n18 585
R548 B.n1101 B.n1100 585
R549 B.n1102 B.n1101 585
R550 B.n1099 B.n23 585
R551 B.n23 B.n22 585
R552 B.n1098 B.n1097 585
R553 B.n1097 B.n1096 585
R554 B.n25 B.n24 585
R555 B.n1095 B.n25 585
R556 B.n1093 B.n1092 585
R557 B.n1094 B.n1093 585
R558 B.n1091 B.n30 585
R559 B.n30 B.n29 585
R560 B.n1090 B.n1089 585
R561 B.n1089 B.n1088 585
R562 B.n32 B.n31 585
R563 B.n1087 B.n32 585
R564 B.n1085 B.n1084 585
R565 B.n1086 B.n1085 585
R566 B.n1083 B.n36 585
R567 B.n39 B.n36 585
R568 B.n1082 B.n1081 585
R569 B.n1081 B.n1080 585
R570 B.n38 B.n37 585
R571 B.n1079 B.n38 585
R572 B.n1077 B.n1076 585
R573 B.n1078 B.n1077 585
R574 B.n1075 B.n44 585
R575 B.n44 B.n43 585
R576 B.n1074 B.n1073 585
R577 B.n1073 B.n1072 585
R578 B.n46 B.n45 585
R579 B.n1071 B.n46 585
R580 B.n1069 B.n1068 585
R581 B.n1070 B.n1069 585
R582 B.n1067 B.n51 585
R583 B.n51 B.n50 585
R584 B.n1066 B.n1065 585
R585 B.n1065 B.n1064 585
R586 B.n53 B.n52 585
R587 B.n1063 B.n53 585
R588 B.n1061 B.n1060 585
R589 B.n1062 B.n1061 585
R590 B.n1059 B.n58 585
R591 B.n58 B.n57 585
R592 B.n1058 B.n1057 585
R593 B.n1057 B.n1056 585
R594 B.n60 B.n59 585
R595 B.n1055 B.n60 585
R596 B.n1053 B.n1052 585
R597 B.n1054 B.n1053 585
R598 B.n1051 B.n65 585
R599 B.n65 B.n64 585
R600 B.n1050 B.n1049 585
R601 B.n1049 B.n1048 585
R602 B.n67 B.n66 585
R603 B.n1047 B.n67 585
R604 B.n1045 B.n1044 585
R605 B.n1046 B.n1045 585
R606 B.n1043 B.n72 585
R607 B.n72 B.n71 585
R608 B.n1042 B.n1041 585
R609 B.n1041 B.n1040 585
R610 B.n74 B.n73 585
R611 B.n1039 B.n74 585
R612 B.n1037 B.n1036 585
R613 B.n1038 B.n1037 585
R614 B.n1122 B.n1121 585
R615 B.n1121 B.n1120 585
R616 B.n581 B.n234 526.135
R617 B.n1037 B.n79 526.135
R618 B.n583 B.n232 526.135
R619 B.n151 B.n77 526.135
R620 B.n273 B.t14 485.899
R621 B.n267 B.t7 485.899
R622 B.n112 B.t16 485.899
R623 B.n118 B.t10 485.899
R624 B.n274 B.t13 410.844
R625 B.n119 B.t11 410.844
R626 B.n268 B.t6 410.844
R627 B.n113 B.t17 410.844
R628 B.n273 B.t12 341.748
R629 B.n267 B.t4 341.748
R630 B.n112 B.t15 341.748
R631 B.n118 B.t8 341.748
R632 B.n764 B.n78 256.663
R633 B.n766 B.n78 256.663
R634 B.n772 B.n78 256.663
R635 B.n774 B.n78 256.663
R636 B.n780 B.n78 256.663
R637 B.n782 B.n78 256.663
R638 B.n788 B.n78 256.663
R639 B.n790 B.n78 256.663
R640 B.n796 B.n78 256.663
R641 B.n798 B.n78 256.663
R642 B.n804 B.n78 256.663
R643 B.n806 B.n78 256.663
R644 B.n812 B.n78 256.663
R645 B.n814 B.n78 256.663
R646 B.n820 B.n78 256.663
R647 B.n822 B.n78 256.663
R648 B.n828 B.n78 256.663
R649 B.n830 B.n78 256.663
R650 B.n836 B.n78 256.663
R651 B.n838 B.n78 256.663
R652 B.n844 B.n78 256.663
R653 B.n846 B.n78 256.663
R654 B.n852 B.n78 256.663
R655 B.n854 B.n78 256.663
R656 B.n860 B.n78 256.663
R657 B.n862 B.n78 256.663
R658 B.n868 B.n78 256.663
R659 B.n870 B.n78 256.663
R660 B.n876 B.n78 256.663
R661 B.n878 B.n78 256.663
R662 B.n884 B.n78 256.663
R663 B.n886 B.n78 256.663
R664 B.n893 B.n78 256.663
R665 B.n895 B.n78 256.663
R666 B.n901 B.n78 256.663
R667 B.n903 B.n78 256.663
R668 B.n910 B.n78 256.663
R669 B.n912 B.n78 256.663
R670 B.n918 B.n78 256.663
R671 B.n920 B.n78 256.663
R672 B.n926 B.n78 256.663
R673 B.n928 B.n78 256.663
R674 B.n934 B.n78 256.663
R675 B.n936 B.n78 256.663
R676 B.n942 B.n78 256.663
R677 B.n944 B.n78 256.663
R678 B.n950 B.n78 256.663
R679 B.n952 B.n78 256.663
R680 B.n958 B.n78 256.663
R681 B.n960 B.n78 256.663
R682 B.n966 B.n78 256.663
R683 B.n968 B.n78 256.663
R684 B.n974 B.n78 256.663
R685 B.n976 B.n78 256.663
R686 B.n982 B.n78 256.663
R687 B.n984 B.n78 256.663
R688 B.n990 B.n78 256.663
R689 B.n992 B.n78 256.663
R690 B.n998 B.n78 256.663
R691 B.n1000 B.n78 256.663
R692 B.n1006 B.n78 256.663
R693 B.n1008 B.n78 256.663
R694 B.n1014 B.n78 256.663
R695 B.n1016 B.n78 256.663
R696 B.n1022 B.n78 256.663
R697 B.n1024 B.n78 256.663
R698 B.n1030 B.n78 256.663
R699 B.n1032 B.n78 256.663
R700 B.n576 B.n233 256.663
R701 B.n236 B.n233 256.663
R702 B.n569 B.n233 256.663
R703 B.n563 B.n233 256.663
R704 B.n561 B.n233 256.663
R705 B.n555 B.n233 256.663
R706 B.n553 B.n233 256.663
R707 B.n547 B.n233 256.663
R708 B.n545 B.n233 256.663
R709 B.n539 B.n233 256.663
R710 B.n537 B.n233 256.663
R711 B.n531 B.n233 256.663
R712 B.n529 B.n233 256.663
R713 B.n523 B.n233 256.663
R714 B.n521 B.n233 256.663
R715 B.n515 B.n233 256.663
R716 B.n513 B.n233 256.663
R717 B.n507 B.n233 256.663
R718 B.n505 B.n233 256.663
R719 B.n499 B.n233 256.663
R720 B.n497 B.n233 256.663
R721 B.n491 B.n233 256.663
R722 B.n489 B.n233 256.663
R723 B.n483 B.n233 256.663
R724 B.n481 B.n233 256.663
R725 B.n475 B.n233 256.663
R726 B.n473 B.n233 256.663
R727 B.n467 B.n233 256.663
R728 B.n465 B.n233 256.663
R729 B.n459 B.n233 256.663
R730 B.n457 B.n233 256.663
R731 B.n450 B.n233 256.663
R732 B.n448 B.n233 256.663
R733 B.n442 B.n233 256.663
R734 B.n440 B.n233 256.663
R735 B.n434 B.n233 256.663
R736 B.n276 B.n233 256.663
R737 B.n428 B.n233 256.663
R738 B.n422 B.n233 256.663
R739 B.n420 B.n233 256.663
R740 B.n414 B.n233 256.663
R741 B.n412 B.n233 256.663
R742 B.n406 B.n233 256.663
R743 B.n404 B.n233 256.663
R744 B.n398 B.n233 256.663
R745 B.n396 B.n233 256.663
R746 B.n390 B.n233 256.663
R747 B.n388 B.n233 256.663
R748 B.n382 B.n233 256.663
R749 B.n380 B.n233 256.663
R750 B.n374 B.n233 256.663
R751 B.n372 B.n233 256.663
R752 B.n366 B.n233 256.663
R753 B.n364 B.n233 256.663
R754 B.n358 B.n233 256.663
R755 B.n356 B.n233 256.663
R756 B.n350 B.n233 256.663
R757 B.n348 B.n233 256.663
R758 B.n342 B.n233 256.663
R759 B.n340 B.n233 256.663
R760 B.n334 B.n233 256.663
R761 B.n332 B.n233 256.663
R762 B.n326 B.n233 256.663
R763 B.n324 B.n233 256.663
R764 B.n318 B.n233 256.663
R765 B.n316 B.n233 256.663
R766 B.n310 B.n233 256.663
R767 B.n308 B.n233 256.663
R768 B.n581 B.n228 163.367
R769 B.n589 B.n228 163.367
R770 B.n589 B.n226 163.367
R771 B.n593 B.n226 163.367
R772 B.n593 B.n220 163.367
R773 B.n601 B.n220 163.367
R774 B.n601 B.n218 163.367
R775 B.n605 B.n218 163.367
R776 B.n605 B.n212 163.367
R777 B.n613 B.n212 163.367
R778 B.n613 B.n210 163.367
R779 B.n617 B.n210 163.367
R780 B.n617 B.n204 163.367
R781 B.n625 B.n204 163.367
R782 B.n625 B.n202 163.367
R783 B.n629 B.n202 163.367
R784 B.n629 B.n196 163.367
R785 B.n637 B.n196 163.367
R786 B.n637 B.n194 163.367
R787 B.n641 B.n194 163.367
R788 B.n641 B.n188 163.367
R789 B.n650 B.n188 163.367
R790 B.n650 B.n186 163.367
R791 B.n654 B.n186 163.367
R792 B.n654 B.n181 163.367
R793 B.n662 B.n181 163.367
R794 B.n662 B.n179 163.367
R795 B.n666 B.n179 163.367
R796 B.n666 B.n173 163.367
R797 B.n674 B.n173 163.367
R798 B.n674 B.n171 163.367
R799 B.n678 B.n171 163.367
R800 B.n678 B.n165 163.367
R801 B.n686 B.n165 163.367
R802 B.n686 B.n163 163.367
R803 B.n690 B.n163 163.367
R804 B.n690 B.n157 163.367
R805 B.n699 B.n157 163.367
R806 B.n699 B.n155 163.367
R807 B.n703 B.n155 163.367
R808 B.n703 B.n2 163.367
R809 B.n1121 B.n2 163.367
R810 B.n1121 B.n3 163.367
R811 B.n1117 B.n3 163.367
R812 B.n1117 B.n9 163.367
R813 B.n1113 B.n9 163.367
R814 B.n1113 B.n11 163.367
R815 B.n1109 B.n11 163.367
R816 B.n1109 B.n16 163.367
R817 B.n1105 B.n16 163.367
R818 B.n1105 B.n18 163.367
R819 B.n1101 B.n18 163.367
R820 B.n1101 B.n23 163.367
R821 B.n1097 B.n23 163.367
R822 B.n1097 B.n25 163.367
R823 B.n1093 B.n25 163.367
R824 B.n1093 B.n30 163.367
R825 B.n1089 B.n30 163.367
R826 B.n1089 B.n32 163.367
R827 B.n1085 B.n32 163.367
R828 B.n1085 B.n36 163.367
R829 B.n1081 B.n36 163.367
R830 B.n1081 B.n38 163.367
R831 B.n1077 B.n38 163.367
R832 B.n1077 B.n44 163.367
R833 B.n1073 B.n44 163.367
R834 B.n1073 B.n46 163.367
R835 B.n1069 B.n46 163.367
R836 B.n1069 B.n51 163.367
R837 B.n1065 B.n51 163.367
R838 B.n1065 B.n53 163.367
R839 B.n1061 B.n53 163.367
R840 B.n1061 B.n58 163.367
R841 B.n1057 B.n58 163.367
R842 B.n1057 B.n60 163.367
R843 B.n1053 B.n60 163.367
R844 B.n1053 B.n65 163.367
R845 B.n1049 B.n65 163.367
R846 B.n1049 B.n67 163.367
R847 B.n1045 B.n67 163.367
R848 B.n1045 B.n72 163.367
R849 B.n1041 B.n72 163.367
R850 B.n1041 B.n74 163.367
R851 B.n1037 B.n74 163.367
R852 B.n577 B.n575 163.367
R853 B.n575 B.n574 163.367
R854 B.n571 B.n570 163.367
R855 B.n568 B.n238 163.367
R856 B.n564 B.n562 163.367
R857 B.n560 B.n240 163.367
R858 B.n556 B.n554 163.367
R859 B.n552 B.n242 163.367
R860 B.n548 B.n546 163.367
R861 B.n544 B.n244 163.367
R862 B.n540 B.n538 163.367
R863 B.n536 B.n246 163.367
R864 B.n532 B.n530 163.367
R865 B.n528 B.n248 163.367
R866 B.n524 B.n522 163.367
R867 B.n520 B.n250 163.367
R868 B.n516 B.n514 163.367
R869 B.n512 B.n252 163.367
R870 B.n508 B.n506 163.367
R871 B.n504 B.n254 163.367
R872 B.n500 B.n498 163.367
R873 B.n496 B.n256 163.367
R874 B.n492 B.n490 163.367
R875 B.n488 B.n258 163.367
R876 B.n484 B.n482 163.367
R877 B.n480 B.n260 163.367
R878 B.n476 B.n474 163.367
R879 B.n472 B.n262 163.367
R880 B.n468 B.n466 163.367
R881 B.n464 B.n264 163.367
R882 B.n460 B.n458 163.367
R883 B.n456 B.n266 163.367
R884 B.n451 B.n449 163.367
R885 B.n447 B.n270 163.367
R886 B.n443 B.n441 163.367
R887 B.n439 B.n272 163.367
R888 B.n435 B.n433 163.367
R889 B.n430 B.n429 163.367
R890 B.n427 B.n278 163.367
R891 B.n423 B.n421 163.367
R892 B.n419 B.n280 163.367
R893 B.n415 B.n413 163.367
R894 B.n411 B.n282 163.367
R895 B.n407 B.n405 163.367
R896 B.n403 B.n284 163.367
R897 B.n399 B.n397 163.367
R898 B.n395 B.n286 163.367
R899 B.n391 B.n389 163.367
R900 B.n387 B.n288 163.367
R901 B.n383 B.n381 163.367
R902 B.n379 B.n290 163.367
R903 B.n375 B.n373 163.367
R904 B.n371 B.n292 163.367
R905 B.n367 B.n365 163.367
R906 B.n363 B.n294 163.367
R907 B.n359 B.n357 163.367
R908 B.n355 B.n296 163.367
R909 B.n351 B.n349 163.367
R910 B.n347 B.n298 163.367
R911 B.n343 B.n341 163.367
R912 B.n339 B.n300 163.367
R913 B.n335 B.n333 163.367
R914 B.n331 B.n302 163.367
R915 B.n327 B.n325 163.367
R916 B.n323 B.n304 163.367
R917 B.n319 B.n317 163.367
R918 B.n315 B.n306 163.367
R919 B.n311 B.n309 163.367
R920 B.n583 B.n230 163.367
R921 B.n587 B.n230 163.367
R922 B.n587 B.n224 163.367
R923 B.n595 B.n224 163.367
R924 B.n595 B.n222 163.367
R925 B.n599 B.n222 163.367
R926 B.n599 B.n216 163.367
R927 B.n607 B.n216 163.367
R928 B.n607 B.n214 163.367
R929 B.n611 B.n214 163.367
R930 B.n611 B.n208 163.367
R931 B.n619 B.n208 163.367
R932 B.n619 B.n206 163.367
R933 B.n623 B.n206 163.367
R934 B.n623 B.n200 163.367
R935 B.n631 B.n200 163.367
R936 B.n631 B.n198 163.367
R937 B.n635 B.n198 163.367
R938 B.n635 B.n192 163.367
R939 B.n643 B.n192 163.367
R940 B.n643 B.n190 163.367
R941 B.n647 B.n190 163.367
R942 B.n647 B.n185 163.367
R943 B.n656 B.n185 163.367
R944 B.n656 B.n183 163.367
R945 B.n660 B.n183 163.367
R946 B.n660 B.n177 163.367
R947 B.n668 B.n177 163.367
R948 B.n668 B.n175 163.367
R949 B.n672 B.n175 163.367
R950 B.n672 B.n169 163.367
R951 B.n680 B.n169 163.367
R952 B.n680 B.n167 163.367
R953 B.n684 B.n167 163.367
R954 B.n684 B.n161 163.367
R955 B.n692 B.n161 163.367
R956 B.n692 B.n159 163.367
R957 B.n697 B.n159 163.367
R958 B.n697 B.n153 163.367
R959 B.n705 B.n153 163.367
R960 B.n706 B.n705 163.367
R961 B.n706 B.n5 163.367
R962 B.n6 B.n5 163.367
R963 B.n7 B.n6 163.367
R964 B.n711 B.n7 163.367
R965 B.n711 B.n12 163.367
R966 B.n13 B.n12 163.367
R967 B.n14 B.n13 163.367
R968 B.n716 B.n14 163.367
R969 B.n716 B.n19 163.367
R970 B.n20 B.n19 163.367
R971 B.n21 B.n20 163.367
R972 B.n721 B.n21 163.367
R973 B.n721 B.n26 163.367
R974 B.n27 B.n26 163.367
R975 B.n28 B.n27 163.367
R976 B.n726 B.n28 163.367
R977 B.n726 B.n33 163.367
R978 B.n34 B.n33 163.367
R979 B.n35 B.n34 163.367
R980 B.n731 B.n35 163.367
R981 B.n731 B.n40 163.367
R982 B.n41 B.n40 163.367
R983 B.n42 B.n41 163.367
R984 B.n736 B.n42 163.367
R985 B.n736 B.n47 163.367
R986 B.n48 B.n47 163.367
R987 B.n49 B.n48 163.367
R988 B.n741 B.n49 163.367
R989 B.n741 B.n54 163.367
R990 B.n55 B.n54 163.367
R991 B.n56 B.n55 163.367
R992 B.n746 B.n56 163.367
R993 B.n746 B.n61 163.367
R994 B.n62 B.n61 163.367
R995 B.n63 B.n62 163.367
R996 B.n751 B.n63 163.367
R997 B.n751 B.n68 163.367
R998 B.n69 B.n68 163.367
R999 B.n70 B.n69 163.367
R1000 B.n756 B.n70 163.367
R1001 B.n756 B.n75 163.367
R1002 B.n76 B.n75 163.367
R1003 B.n77 B.n76 163.367
R1004 B.n1033 B.n1031 163.367
R1005 B.n1029 B.n81 163.367
R1006 B.n1025 B.n1023 163.367
R1007 B.n1021 B.n83 163.367
R1008 B.n1017 B.n1015 163.367
R1009 B.n1013 B.n85 163.367
R1010 B.n1009 B.n1007 163.367
R1011 B.n1005 B.n87 163.367
R1012 B.n1001 B.n999 163.367
R1013 B.n997 B.n89 163.367
R1014 B.n993 B.n991 163.367
R1015 B.n989 B.n91 163.367
R1016 B.n985 B.n983 163.367
R1017 B.n981 B.n93 163.367
R1018 B.n977 B.n975 163.367
R1019 B.n973 B.n95 163.367
R1020 B.n969 B.n967 163.367
R1021 B.n965 B.n97 163.367
R1022 B.n961 B.n959 163.367
R1023 B.n957 B.n99 163.367
R1024 B.n953 B.n951 163.367
R1025 B.n949 B.n101 163.367
R1026 B.n945 B.n943 163.367
R1027 B.n941 B.n103 163.367
R1028 B.n937 B.n935 163.367
R1029 B.n933 B.n105 163.367
R1030 B.n929 B.n927 163.367
R1031 B.n925 B.n107 163.367
R1032 B.n921 B.n919 163.367
R1033 B.n917 B.n109 163.367
R1034 B.n913 B.n911 163.367
R1035 B.n909 B.n111 163.367
R1036 B.n904 B.n902 163.367
R1037 B.n900 B.n115 163.367
R1038 B.n896 B.n894 163.367
R1039 B.n892 B.n117 163.367
R1040 B.n887 B.n885 163.367
R1041 B.n883 B.n121 163.367
R1042 B.n879 B.n877 163.367
R1043 B.n875 B.n123 163.367
R1044 B.n871 B.n869 163.367
R1045 B.n867 B.n125 163.367
R1046 B.n863 B.n861 163.367
R1047 B.n859 B.n127 163.367
R1048 B.n855 B.n853 163.367
R1049 B.n851 B.n129 163.367
R1050 B.n847 B.n845 163.367
R1051 B.n843 B.n131 163.367
R1052 B.n839 B.n837 163.367
R1053 B.n835 B.n133 163.367
R1054 B.n831 B.n829 163.367
R1055 B.n827 B.n135 163.367
R1056 B.n823 B.n821 163.367
R1057 B.n819 B.n137 163.367
R1058 B.n815 B.n813 163.367
R1059 B.n811 B.n139 163.367
R1060 B.n807 B.n805 163.367
R1061 B.n803 B.n141 163.367
R1062 B.n799 B.n797 163.367
R1063 B.n795 B.n143 163.367
R1064 B.n791 B.n789 163.367
R1065 B.n787 B.n145 163.367
R1066 B.n783 B.n781 163.367
R1067 B.n779 B.n147 163.367
R1068 B.n775 B.n773 163.367
R1069 B.n771 B.n149 163.367
R1070 B.n767 B.n765 163.367
R1071 B.n763 B.n151 163.367
R1072 B.n274 B.n273 75.0551
R1073 B.n268 B.n267 75.0551
R1074 B.n113 B.n112 75.0551
R1075 B.n119 B.n118 75.0551
R1076 B.n576 B.n234 71.676
R1077 B.n574 B.n236 71.676
R1078 B.n570 B.n569 71.676
R1079 B.n563 B.n238 71.676
R1080 B.n562 B.n561 71.676
R1081 B.n555 B.n240 71.676
R1082 B.n554 B.n553 71.676
R1083 B.n547 B.n242 71.676
R1084 B.n546 B.n545 71.676
R1085 B.n539 B.n244 71.676
R1086 B.n538 B.n537 71.676
R1087 B.n531 B.n246 71.676
R1088 B.n530 B.n529 71.676
R1089 B.n523 B.n248 71.676
R1090 B.n522 B.n521 71.676
R1091 B.n515 B.n250 71.676
R1092 B.n514 B.n513 71.676
R1093 B.n507 B.n252 71.676
R1094 B.n506 B.n505 71.676
R1095 B.n499 B.n254 71.676
R1096 B.n498 B.n497 71.676
R1097 B.n491 B.n256 71.676
R1098 B.n490 B.n489 71.676
R1099 B.n483 B.n258 71.676
R1100 B.n482 B.n481 71.676
R1101 B.n475 B.n260 71.676
R1102 B.n474 B.n473 71.676
R1103 B.n467 B.n262 71.676
R1104 B.n466 B.n465 71.676
R1105 B.n459 B.n264 71.676
R1106 B.n458 B.n457 71.676
R1107 B.n450 B.n266 71.676
R1108 B.n449 B.n448 71.676
R1109 B.n442 B.n270 71.676
R1110 B.n441 B.n440 71.676
R1111 B.n434 B.n272 71.676
R1112 B.n433 B.n276 71.676
R1113 B.n429 B.n428 71.676
R1114 B.n422 B.n278 71.676
R1115 B.n421 B.n420 71.676
R1116 B.n414 B.n280 71.676
R1117 B.n413 B.n412 71.676
R1118 B.n406 B.n282 71.676
R1119 B.n405 B.n404 71.676
R1120 B.n398 B.n284 71.676
R1121 B.n397 B.n396 71.676
R1122 B.n390 B.n286 71.676
R1123 B.n389 B.n388 71.676
R1124 B.n382 B.n288 71.676
R1125 B.n381 B.n380 71.676
R1126 B.n374 B.n290 71.676
R1127 B.n373 B.n372 71.676
R1128 B.n366 B.n292 71.676
R1129 B.n365 B.n364 71.676
R1130 B.n358 B.n294 71.676
R1131 B.n357 B.n356 71.676
R1132 B.n350 B.n296 71.676
R1133 B.n349 B.n348 71.676
R1134 B.n342 B.n298 71.676
R1135 B.n341 B.n340 71.676
R1136 B.n334 B.n300 71.676
R1137 B.n333 B.n332 71.676
R1138 B.n326 B.n302 71.676
R1139 B.n325 B.n324 71.676
R1140 B.n318 B.n304 71.676
R1141 B.n317 B.n316 71.676
R1142 B.n310 B.n306 71.676
R1143 B.n309 B.n308 71.676
R1144 B.n1032 B.n79 71.676
R1145 B.n1031 B.n1030 71.676
R1146 B.n1024 B.n81 71.676
R1147 B.n1023 B.n1022 71.676
R1148 B.n1016 B.n83 71.676
R1149 B.n1015 B.n1014 71.676
R1150 B.n1008 B.n85 71.676
R1151 B.n1007 B.n1006 71.676
R1152 B.n1000 B.n87 71.676
R1153 B.n999 B.n998 71.676
R1154 B.n992 B.n89 71.676
R1155 B.n991 B.n990 71.676
R1156 B.n984 B.n91 71.676
R1157 B.n983 B.n982 71.676
R1158 B.n976 B.n93 71.676
R1159 B.n975 B.n974 71.676
R1160 B.n968 B.n95 71.676
R1161 B.n967 B.n966 71.676
R1162 B.n960 B.n97 71.676
R1163 B.n959 B.n958 71.676
R1164 B.n952 B.n99 71.676
R1165 B.n951 B.n950 71.676
R1166 B.n944 B.n101 71.676
R1167 B.n943 B.n942 71.676
R1168 B.n936 B.n103 71.676
R1169 B.n935 B.n934 71.676
R1170 B.n928 B.n105 71.676
R1171 B.n927 B.n926 71.676
R1172 B.n920 B.n107 71.676
R1173 B.n919 B.n918 71.676
R1174 B.n912 B.n109 71.676
R1175 B.n911 B.n910 71.676
R1176 B.n903 B.n111 71.676
R1177 B.n902 B.n901 71.676
R1178 B.n895 B.n115 71.676
R1179 B.n894 B.n893 71.676
R1180 B.n886 B.n117 71.676
R1181 B.n885 B.n884 71.676
R1182 B.n878 B.n121 71.676
R1183 B.n877 B.n876 71.676
R1184 B.n870 B.n123 71.676
R1185 B.n869 B.n868 71.676
R1186 B.n862 B.n125 71.676
R1187 B.n861 B.n860 71.676
R1188 B.n854 B.n127 71.676
R1189 B.n853 B.n852 71.676
R1190 B.n846 B.n129 71.676
R1191 B.n845 B.n844 71.676
R1192 B.n838 B.n131 71.676
R1193 B.n837 B.n836 71.676
R1194 B.n830 B.n133 71.676
R1195 B.n829 B.n828 71.676
R1196 B.n822 B.n135 71.676
R1197 B.n821 B.n820 71.676
R1198 B.n814 B.n137 71.676
R1199 B.n813 B.n812 71.676
R1200 B.n806 B.n139 71.676
R1201 B.n805 B.n804 71.676
R1202 B.n798 B.n141 71.676
R1203 B.n797 B.n796 71.676
R1204 B.n790 B.n143 71.676
R1205 B.n789 B.n788 71.676
R1206 B.n782 B.n145 71.676
R1207 B.n781 B.n780 71.676
R1208 B.n774 B.n147 71.676
R1209 B.n773 B.n772 71.676
R1210 B.n766 B.n149 71.676
R1211 B.n765 B.n764 71.676
R1212 B.n764 B.n763 71.676
R1213 B.n767 B.n766 71.676
R1214 B.n772 B.n771 71.676
R1215 B.n775 B.n774 71.676
R1216 B.n780 B.n779 71.676
R1217 B.n783 B.n782 71.676
R1218 B.n788 B.n787 71.676
R1219 B.n791 B.n790 71.676
R1220 B.n796 B.n795 71.676
R1221 B.n799 B.n798 71.676
R1222 B.n804 B.n803 71.676
R1223 B.n807 B.n806 71.676
R1224 B.n812 B.n811 71.676
R1225 B.n815 B.n814 71.676
R1226 B.n820 B.n819 71.676
R1227 B.n823 B.n822 71.676
R1228 B.n828 B.n827 71.676
R1229 B.n831 B.n830 71.676
R1230 B.n836 B.n835 71.676
R1231 B.n839 B.n838 71.676
R1232 B.n844 B.n843 71.676
R1233 B.n847 B.n846 71.676
R1234 B.n852 B.n851 71.676
R1235 B.n855 B.n854 71.676
R1236 B.n860 B.n859 71.676
R1237 B.n863 B.n862 71.676
R1238 B.n868 B.n867 71.676
R1239 B.n871 B.n870 71.676
R1240 B.n876 B.n875 71.676
R1241 B.n879 B.n878 71.676
R1242 B.n884 B.n883 71.676
R1243 B.n887 B.n886 71.676
R1244 B.n893 B.n892 71.676
R1245 B.n896 B.n895 71.676
R1246 B.n901 B.n900 71.676
R1247 B.n904 B.n903 71.676
R1248 B.n910 B.n909 71.676
R1249 B.n913 B.n912 71.676
R1250 B.n918 B.n917 71.676
R1251 B.n921 B.n920 71.676
R1252 B.n926 B.n925 71.676
R1253 B.n929 B.n928 71.676
R1254 B.n934 B.n933 71.676
R1255 B.n937 B.n936 71.676
R1256 B.n942 B.n941 71.676
R1257 B.n945 B.n944 71.676
R1258 B.n950 B.n949 71.676
R1259 B.n953 B.n952 71.676
R1260 B.n958 B.n957 71.676
R1261 B.n961 B.n960 71.676
R1262 B.n966 B.n965 71.676
R1263 B.n969 B.n968 71.676
R1264 B.n974 B.n973 71.676
R1265 B.n977 B.n976 71.676
R1266 B.n982 B.n981 71.676
R1267 B.n985 B.n984 71.676
R1268 B.n990 B.n989 71.676
R1269 B.n993 B.n992 71.676
R1270 B.n998 B.n997 71.676
R1271 B.n1001 B.n1000 71.676
R1272 B.n1006 B.n1005 71.676
R1273 B.n1009 B.n1008 71.676
R1274 B.n1014 B.n1013 71.676
R1275 B.n1017 B.n1016 71.676
R1276 B.n1022 B.n1021 71.676
R1277 B.n1025 B.n1024 71.676
R1278 B.n1030 B.n1029 71.676
R1279 B.n1033 B.n1032 71.676
R1280 B.n577 B.n576 71.676
R1281 B.n571 B.n236 71.676
R1282 B.n569 B.n568 71.676
R1283 B.n564 B.n563 71.676
R1284 B.n561 B.n560 71.676
R1285 B.n556 B.n555 71.676
R1286 B.n553 B.n552 71.676
R1287 B.n548 B.n547 71.676
R1288 B.n545 B.n544 71.676
R1289 B.n540 B.n539 71.676
R1290 B.n537 B.n536 71.676
R1291 B.n532 B.n531 71.676
R1292 B.n529 B.n528 71.676
R1293 B.n524 B.n523 71.676
R1294 B.n521 B.n520 71.676
R1295 B.n516 B.n515 71.676
R1296 B.n513 B.n512 71.676
R1297 B.n508 B.n507 71.676
R1298 B.n505 B.n504 71.676
R1299 B.n500 B.n499 71.676
R1300 B.n497 B.n496 71.676
R1301 B.n492 B.n491 71.676
R1302 B.n489 B.n488 71.676
R1303 B.n484 B.n483 71.676
R1304 B.n481 B.n480 71.676
R1305 B.n476 B.n475 71.676
R1306 B.n473 B.n472 71.676
R1307 B.n468 B.n467 71.676
R1308 B.n465 B.n464 71.676
R1309 B.n460 B.n459 71.676
R1310 B.n457 B.n456 71.676
R1311 B.n451 B.n450 71.676
R1312 B.n448 B.n447 71.676
R1313 B.n443 B.n442 71.676
R1314 B.n440 B.n439 71.676
R1315 B.n435 B.n434 71.676
R1316 B.n430 B.n276 71.676
R1317 B.n428 B.n427 71.676
R1318 B.n423 B.n422 71.676
R1319 B.n420 B.n419 71.676
R1320 B.n415 B.n414 71.676
R1321 B.n412 B.n411 71.676
R1322 B.n407 B.n406 71.676
R1323 B.n404 B.n403 71.676
R1324 B.n399 B.n398 71.676
R1325 B.n396 B.n395 71.676
R1326 B.n391 B.n390 71.676
R1327 B.n388 B.n387 71.676
R1328 B.n383 B.n382 71.676
R1329 B.n380 B.n379 71.676
R1330 B.n375 B.n374 71.676
R1331 B.n372 B.n371 71.676
R1332 B.n367 B.n366 71.676
R1333 B.n364 B.n363 71.676
R1334 B.n359 B.n358 71.676
R1335 B.n356 B.n355 71.676
R1336 B.n351 B.n350 71.676
R1337 B.n348 B.n347 71.676
R1338 B.n343 B.n342 71.676
R1339 B.n340 B.n339 71.676
R1340 B.n335 B.n334 71.676
R1341 B.n332 B.n331 71.676
R1342 B.n327 B.n326 71.676
R1343 B.n324 B.n323 71.676
R1344 B.n319 B.n318 71.676
R1345 B.n316 B.n315 71.676
R1346 B.n311 B.n310 71.676
R1347 B.n308 B.n232 71.676
R1348 B.n582 B.n233 62.6545
R1349 B.n1038 B.n78 62.6545
R1350 B.n275 B.n274 59.5399
R1351 B.n453 B.n268 59.5399
R1352 B.n907 B.n113 59.5399
R1353 B.n889 B.n119 59.5399
R1354 B.n1036 B.n1035 34.1859
R1355 B.n761 B.n760 34.1859
R1356 B.n584 B.n231 34.1859
R1357 B.n580 B.n579 34.1859
R1358 B.n582 B.n229 30.2166
R1359 B.n588 B.n229 30.2166
R1360 B.n588 B.n225 30.2166
R1361 B.n594 B.n225 30.2166
R1362 B.n594 B.n221 30.2166
R1363 B.n600 B.n221 30.2166
R1364 B.n600 B.n217 30.2166
R1365 B.n606 B.n217 30.2166
R1366 B.n612 B.n213 30.2166
R1367 B.n612 B.n209 30.2166
R1368 B.n618 B.n209 30.2166
R1369 B.n618 B.n205 30.2166
R1370 B.n624 B.n205 30.2166
R1371 B.n624 B.n201 30.2166
R1372 B.n630 B.n201 30.2166
R1373 B.n630 B.n197 30.2166
R1374 B.n636 B.n197 30.2166
R1375 B.n636 B.n193 30.2166
R1376 B.n642 B.n193 30.2166
R1377 B.n642 B.n189 30.2166
R1378 B.n649 B.n189 30.2166
R1379 B.n649 B.n648 30.2166
R1380 B.n655 B.n182 30.2166
R1381 B.n661 B.n182 30.2166
R1382 B.n661 B.n178 30.2166
R1383 B.n667 B.n178 30.2166
R1384 B.n667 B.n174 30.2166
R1385 B.n673 B.n174 30.2166
R1386 B.n673 B.n170 30.2166
R1387 B.n679 B.n170 30.2166
R1388 B.n679 B.n166 30.2166
R1389 B.n685 B.n166 30.2166
R1390 B.n691 B.n162 30.2166
R1391 B.n691 B.n158 30.2166
R1392 B.n698 B.n158 30.2166
R1393 B.n698 B.n154 30.2166
R1394 B.n704 B.n154 30.2166
R1395 B.n704 B.n4 30.2166
R1396 B.n1120 B.n4 30.2166
R1397 B.n1120 B.n1119 30.2166
R1398 B.n1119 B.n1118 30.2166
R1399 B.n1118 B.n8 30.2166
R1400 B.n1112 B.n8 30.2166
R1401 B.n1112 B.n1111 30.2166
R1402 B.n1111 B.n1110 30.2166
R1403 B.n1110 B.n15 30.2166
R1404 B.n1104 B.n1103 30.2166
R1405 B.n1103 B.n1102 30.2166
R1406 B.n1102 B.n22 30.2166
R1407 B.n1096 B.n22 30.2166
R1408 B.n1096 B.n1095 30.2166
R1409 B.n1095 B.n1094 30.2166
R1410 B.n1094 B.n29 30.2166
R1411 B.n1088 B.n29 30.2166
R1412 B.n1088 B.n1087 30.2166
R1413 B.n1087 B.n1086 30.2166
R1414 B.n1080 B.n39 30.2166
R1415 B.n1080 B.n1079 30.2166
R1416 B.n1079 B.n1078 30.2166
R1417 B.n1078 B.n43 30.2166
R1418 B.n1072 B.n43 30.2166
R1419 B.n1072 B.n1071 30.2166
R1420 B.n1071 B.n1070 30.2166
R1421 B.n1070 B.n50 30.2166
R1422 B.n1064 B.n50 30.2166
R1423 B.n1064 B.n1063 30.2166
R1424 B.n1063 B.n1062 30.2166
R1425 B.n1062 B.n57 30.2166
R1426 B.n1056 B.n57 30.2166
R1427 B.n1056 B.n1055 30.2166
R1428 B.n1054 B.n64 30.2166
R1429 B.n1048 B.n64 30.2166
R1430 B.n1048 B.n1047 30.2166
R1431 B.n1047 B.n1046 30.2166
R1432 B.n1046 B.n71 30.2166
R1433 B.n1040 B.n71 30.2166
R1434 B.n1040 B.n1039 30.2166
R1435 B.n1039 B.n1038 30.2166
R1436 B.n606 B.t5 22.2182
R1437 B.t9 B.n1054 22.2182
R1438 B.n685 B.t1 21.3295
R1439 B.n1104 B.t0 21.3295
R1440 B.n655 B.t3 20.4408
R1441 B.n1086 B.t2 20.4408
R1442 B B.n1122 18.0485
R1443 B.n1035 B.n1034 10.6151
R1444 B.n1034 B.n80 10.6151
R1445 B.n1028 B.n80 10.6151
R1446 B.n1028 B.n1027 10.6151
R1447 B.n1027 B.n1026 10.6151
R1448 B.n1026 B.n82 10.6151
R1449 B.n1020 B.n82 10.6151
R1450 B.n1020 B.n1019 10.6151
R1451 B.n1019 B.n1018 10.6151
R1452 B.n1018 B.n84 10.6151
R1453 B.n1012 B.n84 10.6151
R1454 B.n1012 B.n1011 10.6151
R1455 B.n1011 B.n1010 10.6151
R1456 B.n1010 B.n86 10.6151
R1457 B.n1004 B.n86 10.6151
R1458 B.n1004 B.n1003 10.6151
R1459 B.n1003 B.n1002 10.6151
R1460 B.n1002 B.n88 10.6151
R1461 B.n996 B.n88 10.6151
R1462 B.n996 B.n995 10.6151
R1463 B.n995 B.n994 10.6151
R1464 B.n994 B.n90 10.6151
R1465 B.n988 B.n90 10.6151
R1466 B.n988 B.n987 10.6151
R1467 B.n987 B.n986 10.6151
R1468 B.n986 B.n92 10.6151
R1469 B.n980 B.n92 10.6151
R1470 B.n980 B.n979 10.6151
R1471 B.n979 B.n978 10.6151
R1472 B.n978 B.n94 10.6151
R1473 B.n972 B.n94 10.6151
R1474 B.n972 B.n971 10.6151
R1475 B.n971 B.n970 10.6151
R1476 B.n970 B.n96 10.6151
R1477 B.n964 B.n96 10.6151
R1478 B.n964 B.n963 10.6151
R1479 B.n963 B.n962 10.6151
R1480 B.n962 B.n98 10.6151
R1481 B.n956 B.n98 10.6151
R1482 B.n956 B.n955 10.6151
R1483 B.n955 B.n954 10.6151
R1484 B.n954 B.n100 10.6151
R1485 B.n948 B.n100 10.6151
R1486 B.n948 B.n947 10.6151
R1487 B.n947 B.n946 10.6151
R1488 B.n946 B.n102 10.6151
R1489 B.n940 B.n102 10.6151
R1490 B.n940 B.n939 10.6151
R1491 B.n939 B.n938 10.6151
R1492 B.n938 B.n104 10.6151
R1493 B.n932 B.n104 10.6151
R1494 B.n932 B.n931 10.6151
R1495 B.n931 B.n930 10.6151
R1496 B.n930 B.n106 10.6151
R1497 B.n924 B.n106 10.6151
R1498 B.n924 B.n923 10.6151
R1499 B.n923 B.n922 10.6151
R1500 B.n922 B.n108 10.6151
R1501 B.n916 B.n108 10.6151
R1502 B.n916 B.n915 10.6151
R1503 B.n915 B.n914 10.6151
R1504 B.n914 B.n110 10.6151
R1505 B.n908 B.n110 10.6151
R1506 B.n906 B.n905 10.6151
R1507 B.n905 B.n114 10.6151
R1508 B.n899 B.n114 10.6151
R1509 B.n899 B.n898 10.6151
R1510 B.n898 B.n897 10.6151
R1511 B.n897 B.n116 10.6151
R1512 B.n891 B.n116 10.6151
R1513 B.n891 B.n890 10.6151
R1514 B.n888 B.n120 10.6151
R1515 B.n882 B.n120 10.6151
R1516 B.n882 B.n881 10.6151
R1517 B.n881 B.n880 10.6151
R1518 B.n880 B.n122 10.6151
R1519 B.n874 B.n122 10.6151
R1520 B.n874 B.n873 10.6151
R1521 B.n873 B.n872 10.6151
R1522 B.n872 B.n124 10.6151
R1523 B.n866 B.n124 10.6151
R1524 B.n866 B.n865 10.6151
R1525 B.n865 B.n864 10.6151
R1526 B.n864 B.n126 10.6151
R1527 B.n858 B.n126 10.6151
R1528 B.n858 B.n857 10.6151
R1529 B.n857 B.n856 10.6151
R1530 B.n856 B.n128 10.6151
R1531 B.n850 B.n128 10.6151
R1532 B.n850 B.n849 10.6151
R1533 B.n849 B.n848 10.6151
R1534 B.n848 B.n130 10.6151
R1535 B.n842 B.n130 10.6151
R1536 B.n842 B.n841 10.6151
R1537 B.n841 B.n840 10.6151
R1538 B.n840 B.n132 10.6151
R1539 B.n834 B.n132 10.6151
R1540 B.n834 B.n833 10.6151
R1541 B.n833 B.n832 10.6151
R1542 B.n832 B.n134 10.6151
R1543 B.n826 B.n134 10.6151
R1544 B.n826 B.n825 10.6151
R1545 B.n825 B.n824 10.6151
R1546 B.n824 B.n136 10.6151
R1547 B.n818 B.n136 10.6151
R1548 B.n818 B.n817 10.6151
R1549 B.n817 B.n816 10.6151
R1550 B.n816 B.n138 10.6151
R1551 B.n810 B.n138 10.6151
R1552 B.n810 B.n809 10.6151
R1553 B.n809 B.n808 10.6151
R1554 B.n808 B.n140 10.6151
R1555 B.n802 B.n140 10.6151
R1556 B.n802 B.n801 10.6151
R1557 B.n801 B.n800 10.6151
R1558 B.n800 B.n142 10.6151
R1559 B.n794 B.n142 10.6151
R1560 B.n794 B.n793 10.6151
R1561 B.n793 B.n792 10.6151
R1562 B.n792 B.n144 10.6151
R1563 B.n786 B.n144 10.6151
R1564 B.n786 B.n785 10.6151
R1565 B.n785 B.n784 10.6151
R1566 B.n784 B.n146 10.6151
R1567 B.n778 B.n146 10.6151
R1568 B.n778 B.n777 10.6151
R1569 B.n777 B.n776 10.6151
R1570 B.n776 B.n148 10.6151
R1571 B.n770 B.n148 10.6151
R1572 B.n770 B.n769 10.6151
R1573 B.n769 B.n768 10.6151
R1574 B.n768 B.n150 10.6151
R1575 B.n762 B.n150 10.6151
R1576 B.n762 B.n761 10.6151
R1577 B.n585 B.n584 10.6151
R1578 B.n586 B.n585 10.6151
R1579 B.n586 B.n223 10.6151
R1580 B.n596 B.n223 10.6151
R1581 B.n597 B.n596 10.6151
R1582 B.n598 B.n597 10.6151
R1583 B.n598 B.n215 10.6151
R1584 B.n608 B.n215 10.6151
R1585 B.n609 B.n608 10.6151
R1586 B.n610 B.n609 10.6151
R1587 B.n610 B.n207 10.6151
R1588 B.n620 B.n207 10.6151
R1589 B.n621 B.n620 10.6151
R1590 B.n622 B.n621 10.6151
R1591 B.n622 B.n199 10.6151
R1592 B.n632 B.n199 10.6151
R1593 B.n633 B.n632 10.6151
R1594 B.n634 B.n633 10.6151
R1595 B.n634 B.n191 10.6151
R1596 B.n644 B.n191 10.6151
R1597 B.n645 B.n644 10.6151
R1598 B.n646 B.n645 10.6151
R1599 B.n646 B.n184 10.6151
R1600 B.n657 B.n184 10.6151
R1601 B.n658 B.n657 10.6151
R1602 B.n659 B.n658 10.6151
R1603 B.n659 B.n176 10.6151
R1604 B.n669 B.n176 10.6151
R1605 B.n670 B.n669 10.6151
R1606 B.n671 B.n670 10.6151
R1607 B.n671 B.n168 10.6151
R1608 B.n681 B.n168 10.6151
R1609 B.n682 B.n681 10.6151
R1610 B.n683 B.n682 10.6151
R1611 B.n683 B.n160 10.6151
R1612 B.n693 B.n160 10.6151
R1613 B.n694 B.n693 10.6151
R1614 B.n696 B.n694 10.6151
R1615 B.n696 B.n695 10.6151
R1616 B.n695 B.n152 10.6151
R1617 B.n707 B.n152 10.6151
R1618 B.n708 B.n707 10.6151
R1619 B.n709 B.n708 10.6151
R1620 B.n710 B.n709 10.6151
R1621 B.n712 B.n710 10.6151
R1622 B.n713 B.n712 10.6151
R1623 B.n714 B.n713 10.6151
R1624 B.n715 B.n714 10.6151
R1625 B.n717 B.n715 10.6151
R1626 B.n718 B.n717 10.6151
R1627 B.n719 B.n718 10.6151
R1628 B.n720 B.n719 10.6151
R1629 B.n722 B.n720 10.6151
R1630 B.n723 B.n722 10.6151
R1631 B.n724 B.n723 10.6151
R1632 B.n725 B.n724 10.6151
R1633 B.n727 B.n725 10.6151
R1634 B.n728 B.n727 10.6151
R1635 B.n729 B.n728 10.6151
R1636 B.n730 B.n729 10.6151
R1637 B.n732 B.n730 10.6151
R1638 B.n733 B.n732 10.6151
R1639 B.n734 B.n733 10.6151
R1640 B.n735 B.n734 10.6151
R1641 B.n737 B.n735 10.6151
R1642 B.n738 B.n737 10.6151
R1643 B.n739 B.n738 10.6151
R1644 B.n740 B.n739 10.6151
R1645 B.n742 B.n740 10.6151
R1646 B.n743 B.n742 10.6151
R1647 B.n744 B.n743 10.6151
R1648 B.n745 B.n744 10.6151
R1649 B.n747 B.n745 10.6151
R1650 B.n748 B.n747 10.6151
R1651 B.n749 B.n748 10.6151
R1652 B.n750 B.n749 10.6151
R1653 B.n752 B.n750 10.6151
R1654 B.n753 B.n752 10.6151
R1655 B.n754 B.n753 10.6151
R1656 B.n755 B.n754 10.6151
R1657 B.n757 B.n755 10.6151
R1658 B.n758 B.n757 10.6151
R1659 B.n759 B.n758 10.6151
R1660 B.n760 B.n759 10.6151
R1661 B.n579 B.n578 10.6151
R1662 B.n578 B.n235 10.6151
R1663 B.n573 B.n235 10.6151
R1664 B.n573 B.n572 10.6151
R1665 B.n572 B.n237 10.6151
R1666 B.n567 B.n237 10.6151
R1667 B.n567 B.n566 10.6151
R1668 B.n566 B.n565 10.6151
R1669 B.n565 B.n239 10.6151
R1670 B.n559 B.n239 10.6151
R1671 B.n559 B.n558 10.6151
R1672 B.n558 B.n557 10.6151
R1673 B.n557 B.n241 10.6151
R1674 B.n551 B.n241 10.6151
R1675 B.n551 B.n550 10.6151
R1676 B.n550 B.n549 10.6151
R1677 B.n549 B.n243 10.6151
R1678 B.n543 B.n243 10.6151
R1679 B.n543 B.n542 10.6151
R1680 B.n542 B.n541 10.6151
R1681 B.n541 B.n245 10.6151
R1682 B.n535 B.n245 10.6151
R1683 B.n535 B.n534 10.6151
R1684 B.n534 B.n533 10.6151
R1685 B.n533 B.n247 10.6151
R1686 B.n527 B.n247 10.6151
R1687 B.n527 B.n526 10.6151
R1688 B.n526 B.n525 10.6151
R1689 B.n525 B.n249 10.6151
R1690 B.n519 B.n249 10.6151
R1691 B.n519 B.n518 10.6151
R1692 B.n518 B.n517 10.6151
R1693 B.n517 B.n251 10.6151
R1694 B.n511 B.n251 10.6151
R1695 B.n511 B.n510 10.6151
R1696 B.n510 B.n509 10.6151
R1697 B.n509 B.n253 10.6151
R1698 B.n503 B.n253 10.6151
R1699 B.n503 B.n502 10.6151
R1700 B.n502 B.n501 10.6151
R1701 B.n501 B.n255 10.6151
R1702 B.n495 B.n255 10.6151
R1703 B.n495 B.n494 10.6151
R1704 B.n494 B.n493 10.6151
R1705 B.n493 B.n257 10.6151
R1706 B.n487 B.n257 10.6151
R1707 B.n487 B.n486 10.6151
R1708 B.n486 B.n485 10.6151
R1709 B.n485 B.n259 10.6151
R1710 B.n479 B.n259 10.6151
R1711 B.n479 B.n478 10.6151
R1712 B.n478 B.n477 10.6151
R1713 B.n477 B.n261 10.6151
R1714 B.n471 B.n261 10.6151
R1715 B.n471 B.n470 10.6151
R1716 B.n470 B.n469 10.6151
R1717 B.n469 B.n263 10.6151
R1718 B.n463 B.n263 10.6151
R1719 B.n463 B.n462 10.6151
R1720 B.n462 B.n461 10.6151
R1721 B.n461 B.n265 10.6151
R1722 B.n455 B.n265 10.6151
R1723 B.n455 B.n454 10.6151
R1724 B.n452 B.n269 10.6151
R1725 B.n446 B.n269 10.6151
R1726 B.n446 B.n445 10.6151
R1727 B.n445 B.n444 10.6151
R1728 B.n444 B.n271 10.6151
R1729 B.n438 B.n271 10.6151
R1730 B.n438 B.n437 10.6151
R1731 B.n437 B.n436 10.6151
R1732 B.n432 B.n431 10.6151
R1733 B.n431 B.n277 10.6151
R1734 B.n426 B.n277 10.6151
R1735 B.n426 B.n425 10.6151
R1736 B.n425 B.n424 10.6151
R1737 B.n424 B.n279 10.6151
R1738 B.n418 B.n279 10.6151
R1739 B.n418 B.n417 10.6151
R1740 B.n417 B.n416 10.6151
R1741 B.n416 B.n281 10.6151
R1742 B.n410 B.n281 10.6151
R1743 B.n410 B.n409 10.6151
R1744 B.n409 B.n408 10.6151
R1745 B.n408 B.n283 10.6151
R1746 B.n402 B.n283 10.6151
R1747 B.n402 B.n401 10.6151
R1748 B.n401 B.n400 10.6151
R1749 B.n400 B.n285 10.6151
R1750 B.n394 B.n285 10.6151
R1751 B.n394 B.n393 10.6151
R1752 B.n393 B.n392 10.6151
R1753 B.n392 B.n287 10.6151
R1754 B.n386 B.n287 10.6151
R1755 B.n386 B.n385 10.6151
R1756 B.n385 B.n384 10.6151
R1757 B.n384 B.n289 10.6151
R1758 B.n378 B.n289 10.6151
R1759 B.n378 B.n377 10.6151
R1760 B.n377 B.n376 10.6151
R1761 B.n376 B.n291 10.6151
R1762 B.n370 B.n291 10.6151
R1763 B.n370 B.n369 10.6151
R1764 B.n369 B.n368 10.6151
R1765 B.n368 B.n293 10.6151
R1766 B.n362 B.n293 10.6151
R1767 B.n362 B.n361 10.6151
R1768 B.n361 B.n360 10.6151
R1769 B.n360 B.n295 10.6151
R1770 B.n354 B.n295 10.6151
R1771 B.n354 B.n353 10.6151
R1772 B.n353 B.n352 10.6151
R1773 B.n352 B.n297 10.6151
R1774 B.n346 B.n297 10.6151
R1775 B.n346 B.n345 10.6151
R1776 B.n345 B.n344 10.6151
R1777 B.n344 B.n299 10.6151
R1778 B.n338 B.n299 10.6151
R1779 B.n338 B.n337 10.6151
R1780 B.n337 B.n336 10.6151
R1781 B.n336 B.n301 10.6151
R1782 B.n330 B.n301 10.6151
R1783 B.n330 B.n329 10.6151
R1784 B.n329 B.n328 10.6151
R1785 B.n328 B.n303 10.6151
R1786 B.n322 B.n303 10.6151
R1787 B.n322 B.n321 10.6151
R1788 B.n321 B.n320 10.6151
R1789 B.n320 B.n305 10.6151
R1790 B.n314 B.n305 10.6151
R1791 B.n314 B.n313 10.6151
R1792 B.n313 B.n312 10.6151
R1793 B.n312 B.n307 10.6151
R1794 B.n307 B.n231 10.6151
R1795 B.n580 B.n227 10.6151
R1796 B.n590 B.n227 10.6151
R1797 B.n591 B.n590 10.6151
R1798 B.n592 B.n591 10.6151
R1799 B.n592 B.n219 10.6151
R1800 B.n602 B.n219 10.6151
R1801 B.n603 B.n602 10.6151
R1802 B.n604 B.n603 10.6151
R1803 B.n604 B.n211 10.6151
R1804 B.n614 B.n211 10.6151
R1805 B.n615 B.n614 10.6151
R1806 B.n616 B.n615 10.6151
R1807 B.n616 B.n203 10.6151
R1808 B.n626 B.n203 10.6151
R1809 B.n627 B.n626 10.6151
R1810 B.n628 B.n627 10.6151
R1811 B.n628 B.n195 10.6151
R1812 B.n638 B.n195 10.6151
R1813 B.n639 B.n638 10.6151
R1814 B.n640 B.n639 10.6151
R1815 B.n640 B.n187 10.6151
R1816 B.n651 B.n187 10.6151
R1817 B.n652 B.n651 10.6151
R1818 B.n653 B.n652 10.6151
R1819 B.n653 B.n180 10.6151
R1820 B.n663 B.n180 10.6151
R1821 B.n664 B.n663 10.6151
R1822 B.n665 B.n664 10.6151
R1823 B.n665 B.n172 10.6151
R1824 B.n675 B.n172 10.6151
R1825 B.n676 B.n675 10.6151
R1826 B.n677 B.n676 10.6151
R1827 B.n677 B.n164 10.6151
R1828 B.n687 B.n164 10.6151
R1829 B.n688 B.n687 10.6151
R1830 B.n689 B.n688 10.6151
R1831 B.n689 B.n156 10.6151
R1832 B.n700 B.n156 10.6151
R1833 B.n701 B.n700 10.6151
R1834 B.n702 B.n701 10.6151
R1835 B.n702 B.n0 10.6151
R1836 B.n1116 B.n1 10.6151
R1837 B.n1116 B.n1115 10.6151
R1838 B.n1115 B.n1114 10.6151
R1839 B.n1114 B.n10 10.6151
R1840 B.n1108 B.n10 10.6151
R1841 B.n1108 B.n1107 10.6151
R1842 B.n1107 B.n1106 10.6151
R1843 B.n1106 B.n17 10.6151
R1844 B.n1100 B.n17 10.6151
R1845 B.n1100 B.n1099 10.6151
R1846 B.n1099 B.n1098 10.6151
R1847 B.n1098 B.n24 10.6151
R1848 B.n1092 B.n24 10.6151
R1849 B.n1092 B.n1091 10.6151
R1850 B.n1091 B.n1090 10.6151
R1851 B.n1090 B.n31 10.6151
R1852 B.n1084 B.n31 10.6151
R1853 B.n1084 B.n1083 10.6151
R1854 B.n1083 B.n1082 10.6151
R1855 B.n1082 B.n37 10.6151
R1856 B.n1076 B.n37 10.6151
R1857 B.n1076 B.n1075 10.6151
R1858 B.n1075 B.n1074 10.6151
R1859 B.n1074 B.n45 10.6151
R1860 B.n1068 B.n45 10.6151
R1861 B.n1068 B.n1067 10.6151
R1862 B.n1067 B.n1066 10.6151
R1863 B.n1066 B.n52 10.6151
R1864 B.n1060 B.n52 10.6151
R1865 B.n1060 B.n1059 10.6151
R1866 B.n1059 B.n1058 10.6151
R1867 B.n1058 B.n59 10.6151
R1868 B.n1052 B.n59 10.6151
R1869 B.n1052 B.n1051 10.6151
R1870 B.n1051 B.n1050 10.6151
R1871 B.n1050 B.n66 10.6151
R1872 B.n1044 B.n66 10.6151
R1873 B.n1044 B.n1043 10.6151
R1874 B.n1043 B.n1042 10.6151
R1875 B.n1042 B.n73 10.6151
R1876 B.n1036 B.n73 10.6151
R1877 B.n648 B.t3 9.7763
R1878 B.n39 B.t2 9.7763
R1879 B.t1 B.n162 8.88759
R1880 B.t0 B.n15 8.88759
R1881 B.t5 B.n213 7.99888
R1882 B.n1055 B.t9 7.99888
R1883 B.n907 B.n906 6.5566
R1884 B.n890 B.n889 6.5566
R1885 B.n453 B.n452 6.5566
R1886 B.n436 B.n275 6.5566
R1887 B.n908 B.n907 4.05904
R1888 B.n889 B.n888 4.05904
R1889 B.n454 B.n453 4.05904
R1890 B.n432 B.n275 4.05904
R1891 B.n1122 B.n0 2.81026
R1892 B.n1122 B.n1 2.81026
R1893 VN.n1 VN.t1 167.321
R1894 VN.n0 VN.t0 167.321
R1895 VN.n0 VN.t3 166.089
R1896 VN.n1 VN.t2 166.089
R1897 VN VN.n1 57.2316
R1898 VN VN.n0 2.15206
R1899 VDD2.n2 VDD2.n0 113.822
R1900 VDD2.n2 VDD2.n1 63.3047
R1901 VDD2.n1 VDD2.t1 1.01693
R1902 VDD2.n1 VDD2.t3 1.01693
R1903 VDD2.n0 VDD2.t0 1.01693
R1904 VDD2.n0 VDD2.t2 1.01693
R1905 VDD2 VDD2.n2 0.0586897
R1906 VTAIL.n842 VTAIL.n742 214.453
R1907 VTAIL.n100 VTAIL.n0 214.453
R1908 VTAIL.n206 VTAIL.n106 214.453
R1909 VTAIL.n312 VTAIL.n212 214.453
R1910 VTAIL.n736 VTAIL.n636 214.453
R1911 VTAIL.n630 VTAIL.n530 214.453
R1912 VTAIL.n524 VTAIL.n424 214.453
R1913 VTAIL.n418 VTAIL.n318 214.453
R1914 VTAIL.n777 VTAIL.n776 185
R1915 VTAIL.n774 VTAIL.n773 185
R1916 VTAIL.n783 VTAIL.n782 185
R1917 VTAIL.n785 VTAIL.n784 185
R1918 VTAIL.n770 VTAIL.n769 185
R1919 VTAIL.n791 VTAIL.n790 185
R1920 VTAIL.n794 VTAIL.n793 185
R1921 VTAIL.n792 VTAIL.n766 185
R1922 VTAIL.n799 VTAIL.n765 185
R1923 VTAIL.n801 VTAIL.n800 185
R1924 VTAIL.n803 VTAIL.n802 185
R1925 VTAIL.n762 VTAIL.n761 185
R1926 VTAIL.n809 VTAIL.n808 185
R1927 VTAIL.n811 VTAIL.n810 185
R1928 VTAIL.n758 VTAIL.n757 185
R1929 VTAIL.n817 VTAIL.n816 185
R1930 VTAIL.n819 VTAIL.n818 185
R1931 VTAIL.n754 VTAIL.n753 185
R1932 VTAIL.n825 VTAIL.n824 185
R1933 VTAIL.n827 VTAIL.n826 185
R1934 VTAIL.n750 VTAIL.n749 185
R1935 VTAIL.n833 VTAIL.n832 185
R1936 VTAIL.n835 VTAIL.n834 185
R1937 VTAIL.n746 VTAIL.n745 185
R1938 VTAIL.n841 VTAIL.n840 185
R1939 VTAIL.n843 VTAIL.n842 185
R1940 VTAIL.n35 VTAIL.n34 185
R1941 VTAIL.n32 VTAIL.n31 185
R1942 VTAIL.n41 VTAIL.n40 185
R1943 VTAIL.n43 VTAIL.n42 185
R1944 VTAIL.n28 VTAIL.n27 185
R1945 VTAIL.n49 VTAIL.n48 185
R1946 VTAIL.n52 VTAIL.n51 185
R1947 VTAIL.n50 VTAIL.n24 185
R1948 VTAIL.n57 VTAIL.n23 185
R1949 VTAIL.n59 VTAIL.n58 185
R1950 VTAIL.n61 VTAIL.n60 185
R1951 VTAIL.n20 VTAIL.n19 185
R1952 VTAIL.n67 VTAIL.n66 185
R1953 VTAIL.n69 VTAIL.n68 185
R1954 VTAIL.n16 VTAIL.n15 185
R1955 VTAIL.n75 VTAIL.n74 185
R1956 VTAIL.n77 VTAIL.n76 185
R1957 VTAIL.n12 VTAIL.n11 185
R1958 VTAIL.n83 VTAIL.n82 185
R1959 VTAIL.n85 VTAIL.n84 185
R1960 VTAIL.n8 VTAIL.n7 185
R1961 VTAIL.n91 VTAIL.n90 185
R1962 VTAIL.n93 VTAIL.n92 185
R1963 VTAIL.n4 VTAIL.n3 185
R1964 VTAIL.n99 VTAIL.n98 185
R1965 VTAIL.n101 VTAIL.n100 185
R1966 VTAIL.n141 VTAIL.n140 185
R1967 VTAIL.n138 VTAIL.n137 185
R1968 VTAIL.n147 VTAIL.n146 185
R1969 VTAIL.n149 VTAIL.n148 185
R1970 VTAIL.n134 VTAIL.n133 185
R1971 VTAIL.n155 VTAIL.n154 185
R1972 VTAIL.n158 VTAIL.n157 185
R1973 VTAIL.n156 VTAIL.n130 185
R1974 VTAIL.n163 VTAIL.n129 185
R1975 VTAIL.n165 VTAIL.n164 185
R1976 VTAIL.n167 VTAIL.n166 185
R1977 VTAIL.n126 VTAIL.n125 185
R1978 VTAIL.n173 VTAIL.n172 185
R1979 VTAIL.n175 VTAIL.n174 185
R1980 VTAIL.n122 VTAIL.n121 185
R1981 VTAIL.n181 VTAIL.n180 185
R1982 VTAIL.n183 VTAIL.n182 185
R1983 VTAIL.n118 VTAIL.n117 185
R1984 VTAIL.n189 VTAIL.n188 185
R1985 VTAIL.n191 VTAIL.n190 185
R1986 VTAIL.n114 VTAIL.n113 185
R1987 VTAIL.n197 VTAIL.n196 185
R1988 VTAIL.n199 VTAIL.n198 185
R1989 VTAIL.n110 VTAIL.n109 185
R1990 VTAIL.n205 VTAIL.n204 185
R1991 VTAIL.n207 VTAIL.n206 185
R1992 VTAIL.n247 VTAIL.n246 185
R1993 VTAIL.n244 VTAIL.n243 185
R1994 VTAIL.n253 VTAIL.n252 185
R1995 VTAIL.n255 VTAIL.n254 185
R1996 VTAIL.n240 VTAIL.n239 185
R1997 VTAIL.n261 VTAIL.n260 185
R1998 VTAIL.n264 VTAIL.n263 185
R1999 VTAIL.n262 VTAIL.n236 185
R2000 VTAIL.n269 VTAIL.n235 185
R2001 VTAIL.n271 VTAIL.n270 185
R2002 VTAIL.n273 VTAIL.n272 185
R2003 VTAIL.n232 VTAIL.n231 185
R2004 VTAIL.n279 VTAIL.n278 185
R2005 VTAIL.n281 VTAIL.n280 185
R2006 VTAIL.n228 VTAIL.n227 185
R2007 VTAIL.n287 VTAIL.n286 185
R2008 VTAIL.n289 VTAIL.n288 185
R2009 VTAIL.n224 VTAIL.n223 185
R2010 VTAIL.n295 VTAIL.n294 185
R2011 VTAIL.n297 VTAIL.n296 185
R2012 VTAIL.n220 VTAIL.n219 185
R2013 VTAIL.n303 VTAIL.n302 185
R2014 VTAIL.n305 VTAIL.n304 185
R2015 VTAIL.n216 VTAIL.n215 185
R2016 VTAIL.n311 VTAIL.n310 185
R2017 VTAIL.n313 VTAIL.n312 185
R2018 VTAIL.n737 VTAIL.n736 185
R2019 VTAIL.n735 VTAIL.n734 185
R2020 VTAIL.n640 VTAIL.n639 185
R2021 VTAIL.n729 VTAIL.n728 185
R2022 VTAIL.n727 VTAIL.n726 185
R2023 VTAIL.n644 VTAIL.n643 185
R2024 VTAIL.n721 VTAIL.n720 185
R2025 VTAIL.n719 VTAIL.n718 185
R2026 VTAIL.n648 VTAIL.n647 185
R2027 VTAIL.n713 VTAIL.n712 185
R2028 VTAIL.n711 VTAIL.n710 185
R2029 VTAIL.n652 VTAIL.n651 185
R2030 VTAIL.n705 VTAIL.n704 185
R2031 VTAIL.n703 VTAIL.n702 185
R2032 VTAIL.n656 VTAIL.n655 185
R2033 VTAIL.n697 VTAIL.n696 185
R2034 VTAIL.n695 VTAIL.n694 185
R2035 VTAIL.n693 VTAIL.n659 185
R2036 VTAIL.n663 VTAIL.n660 185
R2037 VTAIL.n688 VTAIL.n687 185
R2038 VTAIL.n686 VTAIL.n685 185
R2039 VTAIL.n665 VTAIL.n664 185
R2040 VTAIL.n680 VTAIL.n679 185
R2041 VTAIL.n678 VTAIL.n677 185
R2042 VTAIL.n669 VTAIL.n668 185
R2043 VTAIL.n672 VTAIL.n671 185
R2044 VTAIL.n631 VTAIL.n630 185
R2045 VTAIL.n629 VTAIL.n628 185
R2046 VTAIL.n534 VTAIL.n533 185
R2047 VTAIL.n623 VTAIL.n622 185
R2048 VTAIL.n621 VTAIL.n620 185
R2049 VTAIL.n538 VTAIL.n537 185
R2050 VTAIL.n615 VTAIL.n614 185
R2051 VTAIL.n613 VTAIL.n612 185
R2052 VTAIL.n542 VTAIL.n541 185
R2053 VTAIL.n607 VTAIL.n606 185
R2054 VTAIL.n605 VTAIL.n604 185
R2055 VTAIL.n546 VTAIL.n545 185
R2056 VTAIL.n599 VTAIL.n598 185
R2057 VTAIL.n597 VTAIL.n596 185
R2058 VTAIL.n550 VTAIL.n549 185
R2059 VTAIL.n591 VTAIL.n590 185
R2060 VTAIL.n589 VTAIL.n588 185
R2061 VTAIL.n587 VTAIL.n553 185
R2062 VTAIL.n557 VTAIL.n554 185
R2063 VTAIL.n582 VTAIL.n581 185
R2064 VTAIL.n580 VTAIL.n579 185
R2065 VTAIL.n559 VTAIL.n558 185
R2066 VTAIL.n574 VTAIL.n573 185
R2067 VTAIL.n572 VTAIL.n571 185
R2068 VTAIL.n563 VTAIL.n562 185
R2069 VTAIL.n566 VTAIL.n565 185
R2070 VTAIL.n525 VTAIL.n524 185
R2071 VTAIL.n523 VTAIL.n522 185
R2072 VTAIL.n428 VTAIL.n427 185
R2073 VTAIL.n517 VTAIL.n516 185
R2074 VTAIL.n515 VTAIL.n514 185
R2075 VTAIL.n432 VTAIL.n431 185
R2076 VTAIL.n509 VTAIL.n508 185
R2077 VTAIL.n507 VTAIL.n506 185
R2078 VTAIL.n436 VTAIL.n435 185
R2079 VTAIL.n501 VTAIL.n500 185
R2080 VTAIL.n499 VTAIL.n498 185
R2081 VTAIL.n440 VTAIL.n439 185
R2082 VTAIL.n493 VTAIL.n492 185
R2083 VTAIL.n491 VTAIL.n490 185
R2084 VTAIL.n444 VTAIL.n443 185
R2085 VTAIL.n485 VTAIL.n484 185
R2086 VTAIL.n483 VTAIL.n482 185
R2087 VTAIL.n481 VTAIL.n447 185
R2088 VTAIL.n451 VTAIL.n448 185
R2089 VTAIL.n476 VTAIL.n475 185
R2090 VTAIL.n474 VTAIL.n473 185
R2091 VTAIL.n453 VTAIL.n452 185
R2092 VTAIL.n468 VTAIL.n467 185
R2093 VTAIL.n466 VTAIL.n465 185
R2094 VTAIL.n457 VTAIL.n456 185
R2095 VTAIL.n460 VTAIL.n459 185
R2096 VTAIL.n419 VTAIL.n418 185
R2097 VTAIL.n417 VTAIL.n416 185
R2098 VTAIL.n322 VTAIL.n321 185
R2099 VTAIL.n411 VTAIL.n410 185
R2100 VTAIL.n409 VTAIL.n408 185
R2101 VTAIL.n326 VTAIL.n325 185
R2102 VTAIL.n403 VTAIL.n402 185
R2103 VTAIL.n401 VTAIL.n400 185
R2104 VTAIL.n330 VTAIL.n329 185
R2105 VTAIL.n395 VTAIL.n394 185
R2106 VTAIL.n393 VTAIL.n392 185
R2107 VTAIL.n334 VTAIL.n333 185
R2108 VTAIL.n387 VTAIL.n386 185
R2109 VTAIL.n385 VTAIL.n384 185
R2110 VTAIL.n338 VTAIL.n337 185
R2111 VTAIL.n379 VTAIL.n378 185
R2112 VTAIL.n377 VTAIL.n376 185
R2113 VTAIL.n375 VTAIL.n341 185
R2114 VTAIL.n345 VTAIL.n342 185
R2115 VTAIL.n370 VTAIL.n369 185
R2116 VTAIL.n368 VTAIL.n367 185
R2117 VTAIL.n347 VTAIL.n346 185
R2118 VTAIL.n362 VTAIL.n361 185
R2119 VTAIL.n360 VTAIL.n359 185
R2120 VTAIL.n351 VTAIL.n350 185
R2121 VTAIL.n354 VTAIL.n353 185
R2122 VTAIL.t4 VTAIL.n775 149.524
R2123 VTAIL.t7 VTAIL.n33 149.524
R2124 VTAIL.t1 VTAIL.n139 149.524
R2125 VTAIL.t3 VTAIL.n245 149.524
R2126 VTAIL.t2 VTAIL.n670 149.524
R2127 VTAIL.t0 VTAIL.n564 149.524
R2128 VTAIL.t6 VTAIL.n458 149.524
R2129 VTAIL.t5 VTAIL.n352 149.524
R2130 VTAIL.n776 VTAIL.n773 104.615
R2131 VTAIL.n783 VTAIL.n773 104.615
R2132 VTAIL.n784 VTAIL.n783 104.615
R2133 VTAIL.n784 VTAIL.n769 104.615
R2134 VTAIL.n791 VTAIL.n769 104.615
R2135 VTAIL.n793 VTAIL.n791 104.615
R2136 VTAIL.n793 VTAIL.n792 104.615
R2137 VTAIL.n792 VTAIL.n765 104.615
R2138 VTAIL.n801 VTAIL.n765 104.615
R2139 VTAIL.n802 VTAIL.n801 104.615
R2140 VTAIL.n802 VTAIL.n761 104.615
R2141 VTAIL.n809 VTAIL.n761 104.615
R2142 VTAIL.n810 VTAIL.n809 104.615
R2143 VTAIL.n810 VTAIL.n757 104.615
R2144 VTAIL.n817 VTAIL.n757 104.615
R2145 VTAIL.n818 VTAIL.n817 104.615
R2146 VTAIL.n818 VTAIL.n753 104.615
R2147 VTAIL.n825 VTAIL.n753 104.615
R2148 VTAIL.n826 VTAIL.n825 104.615
R2149 VTAIL.n826 VTAIL.n749 104.615
R2150 VTAIL.n833 VTAIL.n749 104.615
R2151 VTAIL.n834 VTAIL.n833 104.615
R2152 VTAIL.n834 VTAIL.n745 104.615
R2153 VTAIL.n841 VTAIL.n745 104.615
R2154 VTAIL.n842 VTAIL.n841 104.615
R2155 VTAIL.n34 VTAIL.n31 104.615
R2156 VTAIL.n41 VTAIL.n31 104.615
R2157 VTAIL.n42 VTAIL.n41 104.615
R2158 VTAIL.n42 VTAIL.n27 104.615
R2159 VTAIL.n49 VTAIL.n27 104.615
R2160 VTAIL.n51 VTAIL.n49 104.615
R2161 VTAIL.n51 VTAIL.n50 104.615
R2162 VTAIL.n50 VTAIL.n23 104.615
R2163 VTAIL.n59 VTAIL.n23 104.615
R2164 VTAIL.n60 VTAIL.n59 104.615
R2165 VTAIL.n60 VTAIL.n19 104.615
R2166 VTAIL.n67 VTAIL.n19 104.615
R2167 VTAIL.n68 VTAIL.n67 104.615
R2168 VTAIL.n68 VTAIL.n15 104.615
R2169 VTAIL.n75 VTAIL.n15 104.615
R2170 VTAIL.n76 VTAIL.n75 104.615
R2171 VTAIL.n76 VTAIL.n11 104.615
R2172 VTAIL.n83 VTAIL.n11 104.615
R2173 VTAIL.n84 VTAIL.n83 104.615
R2174 VTAIL.n84 VTAIL.n7 104.615
R2175 VTAIL.n91 VTAIL.n7 104.615
R2176 VTAIL.n92 VTAIL.n91 104.615
R2177 VTAIL.n92 VTAIL.n3 104.615
R2178 VTAIL.n99 VTAIL.n3 104.615
R2179 VTAIL.n100 VTAIL.n99 104.615
R2180 VTAIL.n140 VTAIL.n137 104.615
R2181 VTAIL.n147 VTAIL.n137 104.615
R2182 VTAIL.n148 VTAIL.n147 104.615
R2183 VTAIL.n148 VTAIL.n133 104.615
R2184 VTAIL.n155 VTAIL.n133 104.615
R2185 VTAIL.n157 VTAIL.n155 104.615
R2186 VTAIL.n157 VTAIL.n156 104.615
R2187 VTAIL.n156 VTAIL.n129 104.615
R2188 VTAIL.n165 VTAIL.n129 104.615
R2189 VTAIL.n166 VTAIL.n165 104.615
R2190 VTAIL.n166 VTAIL.n125 104.615
R2191 VTAIL.n173 VTAIL.n125 104.615
R2192 VTAIL.n174 VTAIL.n173 104.615
R2193 VTAIL.n174 VTAIL.n121 104.615
R2194 VTAIL.n181 VTAIL.n121 104.615
R2195 VTAIL.n182 VTAIL.n181 104.615
R2196 VTAIL.n182 VTAIL.n117 104.615
R2197 VTAIL.n189 VTAIL.n117 104.615
R2198 VTAIL.n190 VTAIL.n189 104.615
R2199 VTAIL.n190 VTAIL.n113 104.615
R2200 VTAIL.n197 VTAIL.n113 104.615
R2201 VTAIL.n198 VTAIL.n197 104.615
R2202 VTAIL.n198 VTAIL.n109 104.615
R2203 VTAIL.n205 VTAIL.n109 104.615
R2204 VTAIL.n206 VTAIL.n205 104.615
R2205 VTAIL.n246 VTAIL.n243 104.615
R2206 VTAIL.n253 VTAIL.n243 104.615
R2207 VTAIL.n254 VTAIL.n253 104.615
R2208 VTAIL.n254 VTAIL.n239 104.615
R2209 VTAIL.n261 VTAIL.n239 104.615
R2210 VTAIL.n263 VTAIL.n261 104.615
R2211 VTAIL.n263 VTAIL.n262 104.615
R2212 VTAIL.n262 VTAIL.n235 104.615
R2213 VTAIL.n271 VTAIL.n235 104.615
R2214 VTAIL.n272 VTAIL.n271 104.615
R2215 VTAIL.n272 VTAIL.n231 104.615
R2216 VTAIL.n279 VTAIL.n231 104.615
R2217 VTAIL.n280 VTAIL.n279 104.615
R2218 VTAIL.n280 VTAIL.n227 104.615
R2219 VTAIL.n287 VTAIL.n227 104.615
R2220 VTAIL.n288 VTAIL.n287 104.615
R2221 VTAIL.n288 VTAIL.n223 104.615
R2222 VTAIL.n295 VTAIL.n223 104.615
R2223 VTAIL.n296 VTAIL.n295 104.615
R2224 VTAIL.n296 VTAIL.n219 104.615
R2225 VTAIL.n303 VTAIL.n219 104.615
R2226 VTAIL.n304 VTAIL.n303 104.615
R2227 VTAIL.n304 VTAIL.n215 104.615
R2228 VTAIL.n311 VTAIL.n215 104.615
R2229 VTAIL.n312 VTAIL.n311 104.615
R2230 VTAIL.n736 VTAIL.n735 104.615
R2231 VTAIL.n735 VTAIL.n639 104.615
R2232 VTAIL.n728 VTAIL.n639 104.615
R2233 VTAIL.n728 VTAIL.n727 104.615
R2234 VTAIL.n727 VTAIL.n643 104.615
R2235 VTAIL.n720 VTAIL.n643 104.615
R2236 VTAIL.n720 VTAIL.n719 104.615
R2237 VTAIL.n719 VTAIL.n647 104.615
R2238 VTAIL.n712 VTAIL.n647 104.615
R2239 VTAIL.n712 VTAIL.n711 104.615
R2240 VTAIL.n711 VTAIL.n651 104.615
R2241 VTAIL.n704 VTAIL.n651 104.615
R2242 VTAIL.n704 VTAIL.n703 104.615
R2243 VTAIL.n703 VTAIL.n655 104.615
R2244 VTAIL.n696 VTAIL.n655 104.615
R2245 VTAIL.n696 VTAIL.n695 104.615
R2246 VTAIL.n695 VTAIL.n659 104.615
R2247 VTAIL.n663 VTAIL.n659 104.615
R2248 VTAIL.n687 VTAIL.n663 104.615
R2249 VTAIL.n687 VTAIL.n686 104.615
R2250 VTAIL.n686 VTAIL.n664 104.615
R2251 VTAIL.n679 VTAIL.n664 104.615
R2252 VTAIL.n679 VTAIL.n678 104.615
R2253 VTAIL.n678 VTAIL.n668 104.615
R2254 VTAIL.n671 VTAIL.n668 104.615
R2255 VTAIL.n630 VTAIL.n629 104.615
R2256 VTAIL.n629 VTAIL.n533 104.615
R2257 VTAIL.n622 VTAIL.n533 104.615
R2258 VTAIL.n622 VTAIL.n621 104.615
R2259 VTAIL.n621 VTAIL.n537 104.615
R2260 VTAIL.n614 VTAIL.n537 104.615
R2261 VTAIL.n614 VTAIL.n613 104.615
R2262 VTAIL.n613 VTAIL.n541 104.615
R2263 VTAIL.n606 VTAIL.n541 104.615
R2264 VTAIL.n606 VTAIL.n605 104.615
R2265 VTAIL.n605 VTAIL.n545 104.615
R2266 VTAIL.n598 VTAIL.n545 104.615
R2267 VTAIL.n598 VTAIL.n597 104.615
R2268 VTAIL.n597 VTAIL.n549 104.615
R2269 VTAIL.n590 VTAIL.n549 104.615
R2270 VTAIL.n590 VTAIL.n589 104.615
R2271 VTAIL.n589 VTAIL.n553 104.615
R2272 VTAIL.n557 VTAIL.n553 104.615
R2273 VTAIL.n581 VTAIL.n557 104.615
R2274 VTAIL.n581 VTAIL.n580 104.615
R2275 VTAIL.n580 VTAIL.n558 104.615
R2276 VTAIL.n573 VTAIL.n558 104.615
R2277 VTAIL.n573 VTAIL.n572 104.615
R2278 VTAIL.n572 VTAIL.n562 104.615
R2279 VTAIL.n565 VTAIL.n562 104.615
R2280 VTAIL.n524 VTAIL.n523 104.615
R2281 VTAIL.n523 VTAIL.n427 104.615
R2282 VTAIL.n516 VTAIL.n427 104.615
R2283 VTAIL.n516 VTAIL.n515 104.615
R2284 VTAIL.n515 VTAIL.n431 104.615
R2285 VTAIL.n508 VTAIL.n431 104.615
R2286 VTAIL.n508 VTAIL.n507 104.615
R2287 VTAIL.n507 VTAIL.n435 104.615
R2288 VTAIL.n500 VTAIL.n435 104.615
R2289 VTAIL.n500 VTAIL.n499 104.615
R2290 VTAIL.n499 VTAIL.n439 104.615
R2291 VTAIL.n492 VTAIL.n439 104.615
R2292 VTAIL.n492 VTAIL.n491 104.615
R2293 VTAIL.n491 VTAIL.n443 104.615
R2294 VTAIL.n484 VTAIL.n443 104.615
R2295 VTAIL.n484 VTAIL.n483 104.615
R2296 VTAIL.n483 VTAIL.n447 104.615
R2297 VTAIL.n451 VTAIL.n447 104.615
R2298 VTAIL.n475 VTAIL.n451 104.615
R2299 VTAIL.n475 VTAIL.n474 104.615
R2300 VTAIL.n474 VTAIL.n452 104.615
R2301 VTAIL.n467 VTAIL.n452 104.615
R2302 VTAIL.n467 VTAIL.n466 104.615
R2303 VTAIL.n466 VTAIL.n456 104.615
R2304 VTAIL.n459 VTAIL.n456 104.615
R2305 VTAIL.n418 VTAIL.n417 104.615
R2306 VTAIL.n417 VTAIL.n321 104.615
R2307 VTAIL.n410 VTAIL.n321 104.615
R2308 VTAIL.n410 VTAIL.n409 104.615
R2309 VTAIL.n409 VTAIL.n325 104.615
R2310 VTAIL.n402 VTAIL.n325 104.615
R2311 VTAIL.n402 VTAIL.n401 104.615
R2312 VTAIL.n401 VTAIL.n329 104.615
R2313 VTAIL.n394 VTAIL.n329 104.615
R2314 VTAIL.n394 VTAIL.n393 104.615
R2315 VTAIL.n393 VTAIL.n333 104.615
R2316 VTAIL.n386 VTAIL.n333 104.615
R2317 VTAIL.n386 VTAIL.n385 104.615
R2318 VTAIL.n385 VTAIL.n337 104.615
R2319 VTAIL.n378 VTAIL.n337 104.615
R2320 VTAIL.n378 VTAIL.n377 104.615
R2321 VTAIL.n377 VTAIL.n341 104.615
R2322 VTAIL.n345 VTAIL.n341 104.615
R2323 VTAIL.n369 VTAIL.n345 104.615
R2324 VTAIL.n369 VTAIL.n368 104.615
R2325 VTAIL.n368 VTAIL.n346 104.615
R2326 VTAIL.n361 VTAIL.n346 104.615
R2327 VTAIL.n361 VTAIL.n360 104.615
R2328 VTAIL.n360 VTAIL.n350 104.615
R2329 VTAIL.n353 VTAIL.n350 104.615
R2330 VTAIL.n776 VTAIL.t4 52.3082
R2331 VTAIL.n34 VTAIL.t7 52.3082
R2332 VTAIL.n140 VTAIL.t1 52.3082
R2333 VTAIL.n246 VTAIL.t3 52.3082
R2334 VTAIL.n671 VTAIL.t2 52.3082
R2335 VTAIL.n565 VTAIL.t0 52.3082
R2336 VTAIL.n459 VTAIL.t6 52.3082
R2337 VTAIL.n353 VTAIL.t5 52.3082
R2338 VTAIL.n847 VTAIL.n846 35.2884
R2339 VTAIL.n105 VTAIL.n104 35.2884
R2340 VTAIL.n211 VTAIL.n210 35.2884
R2341 VTAIL.n317 VTAIL.n316 35.2884
R2342 VTAIL.n741 VTAIL.n740 35.2884
R2343 VTAIL.n635 VTAIL.n634 35.2884
R2344 VTAIL.n529 VTAIL.n528 35.2884
R2345 VTAIL.n423 VTAIL.n422 35.2884
R2346 VTAIL.n847 VTAIL.n741 32.4962
R2347 VTAIL.n423 VTAIL.n317 32.4962
R2348 VTAIL.n800 VTAIL.n799 13.1884
R2349 VTAIL.n58 VTAIL.n57 13.1884
R2350 VTAIL.n164 VTAIL.n163 13.1884
R2351 VTAIL.n270 VTAIL.n269 13.1884
R2352 VTAIL.n694 VTAIL.n693 13.1884
R2353 VTAIL.n588 VTAIL.n587 13.1884
R2354 VTAIL.n482 VTAIL.n481 13.1884
R2355 VTAIL.n376 VTAIL.n375 13.1884
R2356 VTAIL.n798 VTAIL.n766 12.8005
R2357 VTAIL.n803 VTAIL.n764 12.8005
R2358 VTAIL.n844 VTAIL.n843 12.8005
R2359 VTAIL.n56 VTAIL.n24 12.8005
R2360 VTAIL.n61 VTAIL.n22 12.8005
R2361 VTAIL.n102 VTAIL.n101 12.8005
R2362 VTAIL.n162 VTAIL.n130 12.8005
R2363 VTAIL.n167 VTAIL.n128 12.8005
R2364 VTAIL.n208 VTAIL.n207 12.8005
R2365 VTAIL.n268 VTAIL.n236 12.8005
R2366 VTAIL.n273 VTAIL.n234 12.8005
R2367 VTAIL.n314 VTAIL.n313 12.8005
R2368 VTAIL.n738 VTAIL.n737 12.8005
R2369 VTAIL.n697 VTAIL.n658 12.8005
R2370 VTAIL.n692 VTAIL.n660 12.8005
R2371 VTAIL.n632 VTAIL.n631 12.8005
R2372 VTAIL.n591 VTAIL.n552 12.8005
R2373 VTAIL.n586 VTAIL.n554 12.8005
R2374 VTAIL.n526 VTAIL.n525 12.8005
R2375 VTAIL.n485 VTAIL.n446 12.8005
R2376 VTAIL.n480 VTAIL.n448 12.8005
R2377 VTAIL.n420 VTAIL.n419 12.8005
R2378 VTAIL.n379 VTAIL.n340 12.8005
R2379 VTAIL.n374 VTAIL.n342 12.8005
R2380 VTAIL.n795 VTAIL.n794 12.0247
R2381 VTAIL.n804 VTAIL.n762 12.0247
R2382 VTAIL.n840 VTAIL.n744 12.0247
R2383 VTAIL.n53 VTAIL.n52 12.0247
R2384 VTAIL.n62 VTAIL.n20 12.0247
R2385 VTAIL.n98 VTAIL.n2 12.0247
R2386 VTAIL.n159 VTAIL.n158 12.0247
R2387 VTAIL.n168 VTAIL.n126 12.0247
R2388 VTAIL.n204 VTAIL.n108 12.0247
R2389 VTAIL.n265 VTAIL.n264 12.0247
R2390 VTAIL.n274 VTAIL.n232 12.0247
R2391 VTAIL.n310 VTAIL.n214 12.0247
R2392 VTAIL.n734 VTAIL.n638 12.0247
R2393 VTAIL.n698 VTAIL.n656 12.0247
R2394 VTAIL.n689 VTAIL.n688 12.0247
R2395 VTAIL.n628 VTAIL.n532 12.0247
R2396 VTAIL.n592 VTAIL.n550 12.0247
R2397 VTAIL.n583 VTAIL.n582 12.0247
R2398 VTAIL.n522 VTAIL.n426 12.0247
R2399 VTAIL.n486 VTAIL.n444 12.0247
R2400 VTAIL.n477 VTAIL.n476 12.0247
R2401 VTAIL.n416 VTAIL.n320 12.0247
R2402 VTAIL.n380 VTAIL.n338 12.0247
R2403 VTAIL.n371 VTAIL.n370 12.0247
R2404 VTAIL.n790 VTAIL.n768 11.249
R2405 VTAIL.n808 VTAIL.n807 11.249
R2406 VTAIL.n839 VTAIL.n746 11.249
R2407 VTAIL.n48 VTAIL.n26 11.249
R2408 VTAIL.n66 VTAIL.n65 11.249
R2409 VTAIL.n97 VTAIL.n4 11.249
R2410 VTAIL.n154 VTAIL.n132 11.249
R2411 VTAIL.n172 VTAIL.n171 11.249
R2412 VTAIL.n203 VTAIL.n110 11.249
R2413 VTAIL.n260 VTAIL.n238 11.249
R2414 VTAIL.n278 VTAIL.n277 11.249
R2415 VTAIL.n309 VTAIL.n216 11.249
R2416 VTAIL.n733 VTAIL.n640 11.249
R2417 VTAIL.n702 VTAIL.n701 11.249
R2418 VTAIL.n685 VTAIL.n662 11.249
R2419 VTAIL.n627 VTAIL.n534 11.249
R2420 VTAIL.n596 VTAIL.n595 11.249
R2421 VTAIL.n579 VTAIL.n556 11.249
R2422 VTAIL.n521 VTAIL.n428 11.249
R2423 VTAIL.n490 VTAIL.n489 11.249
R2424 VTAIL.n473 VTAIL.n450 11.249
R2425 VTAIL.n415 VTAIL.n322 11.249
R2426 VTAIL.n384 VTAIL.n383 11.249
R2427 VTAIL.n367 VTAIL.n344 11.249
R2428 VTAIL.n789 VTAIL.n770 10.4732
R2429 VTAIL.n811 VTAIL.n760 10.4732
R2430 VTAIL.n836 VTAIL.n835 10.4732
R2431 VTAIL.n47 VTAIL.n28 10.4732
R2432 VTAIL.n69 VTAIL.n18 10.4732
R2433 VTAIL.n94 VTAIL.n93 10.4732
R2434 VTAIL.n153 VTAIL.n134 10.4732
R2435 VTAIL.n175 VTAIL.n124 10.4732
R2436 VTAIL.n200 VTAIL.n199 10.4732
R2437 VTAIL.n259 VTAIL.n240 10.4732
R2438 VTAIL.n281 VTAIL.n230 10.4732
R2439 VTAIL.n306 VTAIL.n305 10.4732
R2440 VTAIL.n730 VTAIL.n729 10.4732
R2441 VTAIL.n705 VTAIL.n654 10.4732
R2442 VTAIL.n684 VTAIL.n665 10.4732
R2443 VTAIL.n624 VTAIL.n623 10.4732
R2444 VTAIL.n599 VTAIL.n548 10.4732
R2445 VTAIL.n578 VTAIL.n559 10.4732
R2446 VTAIL.n518 VTAIL.n517 10.4732
R2447 VTAIL.n493 VTAIL.n442 10.4732
R2448 VTAIL.n472 VTAIL.n453 10.4732
R2449 VTAIL.n412 VTAIL.n411 10.4732
R2450 VTAIL.n387 VTAIL.n336 10.4732
R2451 VTAIL.n366 VTAIL.n347 10.4732
R2452 VTAIL.n777 VTAIL.n775 10.2747
R2453 VTAIL.n35 VTAIL.n33 10.2747
R2454 VTAIL.n141 VTAIL.n139 10.2747
R2455 VTAIL.n247 VTAIL.n245 10.2747
R2456 VTAIL.n672 VTAIL.n670 10.2747
R2457 VTAIL.n566 VTAIL.n564 10.2747
R2458 VTAIL.n460 VTAIL.n458 10.2747
R2459 VTAIL.n354 VTAIL.n352 10.2747
R2460 VTAIL.n786 VTAIL.n785 9.69747
R2461 VTAIL.n812 VTAIL.n758 9.69747
R2462 VTAIL.n832 VTAIL.n748 9.69747
R2463 VTAIL.n44 VTAIL.n43 9.69747
R2464 VTAIL.n70 VTAIL.n16 9.69747
R2465 VTAIL.n90 VTAIL.n6 9.69747
R2466 VTAIL.n150 VTAIL.n149 9.69747
R2467 VTAIL.n176 VTAIL.n122 9.69747
R2468 VTAIL.n196 VTAIL.n112 9.69747
R2469 VTAIL.n256 VTAIL.n255 9.69747
R2470 VTAIL.n282 VTAIL.n228 9.69747
R2471 VTAIL.n302 VTAIL.n218 9.69747
R2472 VTAIL.n726 VTAIL.n642 9.69747
R2473 VTAIL.n706 VTAIL.n652 9.69747
R2474 VTAIL.n681 VTAIL.n680 9.69747
R2475 VTAIL.n620 VTAIL.n536 9.69747
R2476 VTAIL.n600 VTAIL.n546 9.69747
R2477 VTAIL.n575 VTAIL.n574 9.69747
R2478 VTAIL.n514 VTAIL.n430 9.69747
R2479 VTAIL.n494 VTAIL.n440 9.69747
R2480 VTAIL.n469 VTAIL.n468 9.69747
R2481 VTAIL.n408 VTAIL.n324 9.69747
R2482 VTAIL.n388 VTAIL.n334 9.69747
R2483 VTAIL.n363 VTAIL.n362 9.69747
R2484 VTAIL.n846 VTAIL.n845 9.45567
R2485 VTAIL.n104 VTAIL.n103 9.45567
R2486 VTAIL.n210 VTAIL.n209 9.45567
R2487 VTAIL.n316 VTAIL.n315 9.45567
R2488 VTAIL.n740 VTAIL.n739 9.45567
R2489 VTAIL.n634 VTAIL.n633 9.45567
R2490 VTAIL.n528 VTAIL.n527 9.45567
R2491 VTAIL.n422 VTAIL.n421 9.45567
R2492 VTAIL.n821 VTAIL.n820 9.3005
R2493 VTAIL.n756 VTAIL.n755 9.3005
R2494 VTAIL.n815 VTAIL.n814 9.3005
R2495 VTAIL.n813 VTAIL.n812 9.3005
R2496 VTAIL.n760 VTAIL.n759 9.3005
R2497 VTAIL.n807 VTAIL.n806 9.3005
R2498 VTAIL.n805 VTAIL.n804 9.3005
R2499 VTAIL.n764 VTAIL.n763 9.3005
R2500 VTAIL.n779 VTAIL.n778 9.3005
R2501 VTAIL.n781 VTAIL.n780 9.3005
R2502 VTAIL.n772 VTAIL.n771 9.3005
R2503 VTAIL.n787 VTAIL.n786 9.3005
R2504 VTAIL.n789 VTAIL.n788 9.3005
R2505 VTAIL.n768 VTAIL.n767 9.3005
R2506 VTAIL.n796 VTAIL.n795 9.3005
R2507 VTAIL.n798 VTAIL.n797 9.3005
R2508 VTAIL.n823 VTAIL.n822 9.3005
R2509 VTAIL.n752 VTAIL.n751 9.3005
R2510 VTAIL.n829 VTAIL.n828 9.3005
R2511 VTAIL.n831 VTAIL.n830 9.3005
R2512 VTAIL.n748 VTAIL.n747 9.3005
R2513 VTAIL.n837 VTAIL.n836 9.3005
R2514 VTAIL.n839 VTAIL.n838 9.3005
R2515 VTAIL.n744 VTAIL.n743 9.3005
R2516 VTAIL.n845 VTAIL.n844 9.3005
R2517 VTAIL.n79 VTAIL.n78 9.3005
R2518 VTAIL.n14 VTAIL.n13 9.3005
R2519 VTAIL.n73 VTAIL.n72 9.3005
R2520 VTAIL.n71 VTAIL.n70 9.3005
R2521 VTAIL.n18 VTAIL.n17 9.3005
R2522 VTAIL.n65 VTAIL.n64 9.3005
R2523 VTAIL.n63 VTAIL.n62 9.3005
R2524 VTAIL.n22 VTAIL.n21 9.3005
R2525 VTAIL.n37 VTAIL.n36 9.3005
R2526 VTAIL.n39 VTAIL.n38 9.3005
R2527 VTAIL.n30 VTAIL.n29 9.3005
R2528 VTAIL.n45 VTAIL.n44 9.3005
R2529 VTAIL.n47 VTAIL.n46 9.3005
R2530 VTAIL.n26 VTAIL.n25 9.3005
R2531 VTAIL.n54 VTAIL.n53 9.3005
R2532 VTAIL.n56 VTAIL.n55 9.3005
R2533 VTAIL.n81 VTAIL.n80 9.3005
R2534 VTAIL.n10 VTAIL.n9 9.3005
R2535 VTAIL.n87 VTAIL.n86 9.3005
R2536 VTAIL.n89 VTAIL.n88 9.3005
R2537 VTAIL.n6 VTAIL.n5 9.3005
R2538 VTAIL.n95 VTAIL.n94 9.3005
R2539 VTAIL.n97 VTAIL.n96 9.3005
R2540 VTAIL.n2 VTAIL.n1 9.3005
R2541 VTAIL.n103 VTAIL.n102 9.3005
R2542 VTAIL.n185 VTAIL.n184 9.3005
R2543 VTAIL.n120 VTAIL.n119 9.3005
R2544 VTAIL.n179 VTAIL.n178 9.3005
R2545 VTAIL.n177 VTAIL.n176 9.3005
R2546 VTAIL.n124 VTAIL.n123 9.3005
R2547 VTAIL.n171 VTAIL.n170 9.3005
R2548 VTAIL.n169 VTAIL.n168 9.3005
R2549 VTAIL.n128 VTAIL.n127 9.3005
R2550 VTAIL.n143 VTAIL.n142 9.3005
R2551 VTAIL.n145 VTAIL.n144 9.3005
R2552 VTAIL.n136 VTAIL.n135 9.3005
R2553 VTAIL.n151 VTAIL.n150 9.3005
R2554 VTAIL.n153 VTAIL.n152 9.3005
R2555 VTAIL.n132 VTAIL.n131 9.3005
R2556 VTAIL.n160 VTAIL.n159 9.3005
R2557 VTAIL.n162 VTAIL.n161 9.3005
R2558 VTAIL.n187 VTAIL.n186 9.3005
R2559 VTAIL.n116 VTAIL.n115 9.3005
R2560 VTAIL.n193 VTAIL.n192 9.3005
R2561 VTAIL.n195 VTAIL.n194 9.3005
R2562 VTAIL.n112 VTAIL.n111 9.3005
R2563 VTAIL.n201 VTAIL.n200 9.3005
R2564 VTAIL.n203 VTAIL.n202 9.3005
R2565 VTAIL.n108 VTAIL.n107 9.3005
R2566 VTAIL.n209 VTAIL.n208 9.3005
R2567 VTAIL.n291 VTAIL.n290 9.3005
R2568 VTAIL.n226 VTAIL.n225 9.3005
R2569 VTAIL.n285 VTAIL.n284 9.3005
R2570 VTAIL.n283 VTAIL.n282 9.3005
R2571 VTAIL.n230 VTAIL.n229 9.3005
R2572 VTAIL.n277 VTAIL.n276 9.3005
R2573 VTAIL.n275 VTAIL.n274 9.3005
R2574 VTAIL.n234 VTAIL.n233 9.3005
R2575 VTAIL.n249 VTAIL.n248 9.3005
R2576 VTAIL.n251 VTAIL.n250 9.3005
R2577 VTAIL.n242 VTAIL.n241 9.3005
R2578 VTAIL.n257 VTAIL.n256 9.3005
R2579 VTAIL.n259 VTAIL.n258 9.3005
R2580 VTAIL.n238 VTAIL.n237 9.3005
R2581 VTAIL.n266 VTAIL.n265 9.3005
R2582 VTAIL.n268 VTAIL.n267 9.3005
R2583 VTAIL.n293 VTAIL.n292 9.3005
R2584 VTAIL.n222 VTAIL.n221 9.3005
R2585 VTAIL.n299 VTAIL.n298 9.3005
R2586 VTAIL.n301 VTAIL.n300 9.3005
R2587 VTAIL.n218 VTAIL.n217 9.3005
R2588 VTAIL.n307 VTAIL.n306 9.3005
R2589 VTAIL.n309 VTAIL.n308 9.3005
R2590 VTAIL.n214 VTAIL.n213 9.3005
R2591 VTAIL.n315 VTAIL.n314 9.3005
R2592 VTAIL.n674 VTAIL.n673 9.3005
R2593 VTAIL.n676 VTAIL.n675 9.3005
R2594 VTAIL.n667 VTAIL.n666 9.3005
R2595 VTAIL.n682 VTAIL.n681 9.3005
R2596 VTAIL.n684 VTAIL.n683 9.3005
R2597 VTAIL.n662 VTAIL.n661 9.3005
R2598 VTAIL.n690 VTAIL.n689 9.3005
R2599 VTAIL.n692 VTAIL.n691 9.3005
R2600 VTAIL.n646 VTAIL.n645 9.3005
R2601 VTAIL.n723 VTAIL.n722 9.3005
R2602 VTAIL.n725 VTAIL.n724 9.3005
R2603 VTAIL.n642 VTAIL.n641 9.3005
R2604 VTAIL.n731 VTAIL.n730 9.3005
R2605 VTAIL.n733 VTAIL.n732 9.3005
R2606 VTAIL.n638 VTAIL.n637 9.3005
R2607 VTAIL.n739 VTAIL.n738 9.3005
R2608 VTAIL.n717 VTAIL.n716 9.3005
R2609 VTAIL.n715 VTAIL.n714 9.3005
R2610 VTAIL.n650 VTAIL.n649 9.3005
R2611 VTAIL.n709 VTAIL.n708 9.3005
R2612 VTAIL.n707 VTAIL.n706 9.3005
R2613 VTAIL.n654 VTAIL.n653 9.3005
R2614 VTAIL.n701 VTAIL.n700 9.3005
R2615 VTAIL.n699 VTAIL.n698 9.3005
R2616 VTAIL.n658 VTAIL.n657 9.3005
R2617 VTAIL.n568 VTAIL.n567 9.3005
R2618 VTAIL.n570 VTAIL.n569 9.3005
R2619 VTAIL.n561 VTAIL.n560 9.3005
R2620 VTAIL.n576 VTAIL.n575 9.3005
R2621 VTAIL.n578 VTAIL.n577 9.3005
R2622 VTAIL.n556 VTAIL.n555 9.3005
R2623 VTAIL.n584 VTAIL.n583 9.3005
R2624 VTAIL.n586 VTAIL.n585 9.3005
R2625 VTAIL.n540 VTAIL.n539 9.3005
R2626 VTAIL.n617 VTAIL.n616 9.3005
R2627 VTAIL.n619 VTAIL.n618 9.3005
R2628 VTAIL.n536 VTAIL.n535 9.3005
R2629 VTAIL.n625 VTAIL.n624 9.3005
R2630 VTAIL.n627 VTAIL.n626 9.3005
R2631 VTAIL.n532 VTAIL.n531 9.3005
R2632 VTAIL.n633 VTAIL.n632 9.3005
R2633 VTAIL.n611 VTAIL.n610 9.3005
R2634 VTAIL.n609 VTAIL.n608 9.3005
R2635 VTAIL.n544 VTAIL.n543 9.3005
R2636 VTAIL.n603 VTAIL.n602 9.3005
R2637 VTAIL.n601 VTAIL.n600 9.3005
R2638 VTAIL.n548 VTAIL.n547 9.3005
R2639 VTAIL.n595 VTAIL.n594 9.3005
R2640 VTAIL.n593 VTAIL.n592 9.3005
R2641 VTAIL.n552 VTAIL.n551 9.3005
R2642 VTAIL.n462 VTAIL.n461 9.3005
R2643 VTAIL.n464 VTAIL.n463 9.3005
R2644 VTAIL.n455 VTAIL.n454 9.3005
R2645 VTAIL.n470 VTAIL.n469 9.3005
R2646 VTAIL.n472 VTAIL.n471 9.3005
R2647 VTAIL.n450 VTAIL.n449 9.3005
R2648 VTAIL.n478 VTAIL.n477 9.3005
R2649 VTAIL.n480 VTAIL.n479 9.3005
R2650 VTAIL.n434 VTAIL.n433 9.3005
R2651 VTAIL.n511 VTAIL.n510 9.3005
R2652 VTAIL.n513 VTAIL.n512 9.3005
R2653 VTAIL.n430 VTAIL.n429 9.3005
R2654 VTAIL.n519 VTAIL.n518 9.3005
R2655 VTAIL.n521 VTAIL.n520 9.3005
R2656 VTAIL.n426 VTAIL.n425 9.3005
R2657 VTAIL.n527 VTAIL.n526 9.3005
R2658 VTAIL.n505 VTAIL.n504 9.3005
R2659 VTAIL.n503 VTAIL.n502 9.3005
R2660 VTAIL.n438 VTAIL.n437 9.3005
R2661 VTAIL.n497 VTAIL.n496 9.3005
R2662 VTAIL.n495 VTAIL.n494 9.3005
R2663 VTAIL.n442 VTAIL.n441 9.3005
R2664 VTAIL.n489 VTAIL.n488 9.3005
R2665 VTAIL.n487 VTAIL.n486 9.3005
R2666 VTAIL.n446 VTAIL.n445 9.3005
R2667 VTAIL.n356 VTAIL.n355 9.3005
R2668 VTAIL.n358 VTAIL.n357 9.3005
R2669 VTAIL.n349 VTAIL.n348 9.3005
R2670 VTAIL.n364 VTAIL.n363 9.3005
R2671 VTAIL.n366 VTAIL.n365 9.3005
R2672 VTAIL.n344 VTAIL.n343 9.3005
R2673 VTAIL.n372 VTAIL.n371 9.3005
R2674 VTAIL.n374 VTAIL.n373 9.3005
R2675 VTAIL.n328 VTAIL.n327 9.3005
R2676 VTAIL.n405 VTAIL.n404 9.3005
R2677 VTAIL.n407 VTAIL.n406 9.3005
R2678 VTAIL.n324 VTAIL.n323 9.3005
R2679 VTAIL.n413 VTAIL.n412 9.3005
R2680 VTAIL.n415 VTAIL.n414 9.3005
R2681 VTAIL.n320 VTAIL.n319 9.3005
R2682 VTAIL.n421 VTAIL.n420 9.3005
R2683 VTAIL.n399 VTAIL.n398 9.3005
R2684 VTAIL.n397 VTAIL.n396 9.3005
R2685 VTAIL.n332 VTAIL.n331 9.3005
R2686 VTAIL.n391 VTAIL.n390 9.3005
R2687 VTAIL.n389 VTAIL.n388 9.3005
R2688 VTAIL.n336 VTAIL.n335 9.3005
R2689 VTAIL.n383 VTAIL.n382 9.3005
R2690 VTAIL.n381 VTAIL.n380 9.3005
R2691 VTAIL.n340 VTAIL.n339 9.3005
R2692 VTAIL.n782 VTAIL.n772 8.92171
R2693 VTAIL.n816 VTAIL.n815 8.92171
R2694 VTAIL.n831 VTAIL.n750 8.92171
R2695 VTAIL.n40 VTAIL.n30 8.92171
R2696 VTAIL.n74 VTAIL.n73 8.92171
R2697 VTAIL.n89 VTAIL.n8 8.92171
R2698 VTAIL.n146 VTAIL.n136 8.92171
R2699 VTAIL.n180 VTAIL.n179 8.92171
R2700 VTAIL.n195 VTAIL.n114 8.92171
R2701 VTAIL.n252 VTAIL.n242 8.92171
R2702 VTAIL.n286 VTAIL.n285 8.92171
R2703 VTAIL.n301 VTAIL.n220 8.92171
R2704 VTAIL.n725 VTAIL.n644 8.92171
R2705 VTAIL.n710 VTAIL.n709 8.92171
R2706 VTAIL.n677 VTAIL.n667 8.92171
R2707 VTAIL.n619 VTAIL.n538 8.92171
R2708 VTAIL.n604 VTAIL.n603 8.92171
R2709 VTAIL.n571 VTAIL.n561 8.92171
R2710 VTAIL.n513 VTAIL.n432 8.92171
R2711 VTAIL.n498 VTAIL.n497 8.92171
R2712 VTAIL.n465 VTAIL.n455 8.92171
R2713 VTAIL.n407 VTAIL.n326 8.92171
R2714 VTAIL.n392 VTAIL.n391 8.92171
R2715 VTAIL.n359 VTAIL.n349 8.92171
R2716 VTAIL.n846 VTAIL.n742 8.2187
R2717 VTAIL.n104 VTAIL.n0 8.2187
R2718 VTAIL.n210 VTAIL.n106 8.2187
R2719 VTAIL.n316 VTAIL.n212 8.2187
R2720 VTAIL.n740 VTAIL.n636 8.2187
R2721 VTAIL.n634 VTAIL.n530 8.2187
R2722 VTAIL.n528 VTAIL.n424 8.2187
R2723 VTAIL.n422 VTAIL.n318 8.2187
R2724 VTAIL.n781 VTAIL.n774 8.14595
R2725 VTAIL.n819 VTAIL.n756 8.14595
R2726 VTAIL.n828 VTAIL.n827 8.14595
R2727 VTAIL.n39 VTAIL.n32 8.14595
R2728 VTAIL.n77 VTAIL.n14 8.14595
R2729 VTAIL.n86 VTAIL.n85 8.14595
R2730 VTAIL.n145 VTAIL.n138 8.14595
R2731 VTAIL.n183 VTAIL.n120 8.14595
R2732 VTAIL.n192 VTAIL.n191 8.14595
R2733 VTAIL.n251 VTAIL.n244 8.14595
R2734 VTAIL.n289 VTAIL.n226 8.14595
R2735 VTAIL.n298 VTAIL.n297 8.14595
R2736 VTAIL.n722 VTAIL.n721 8.14595
R2737 VTAIL.n713 VTAIL.n650 8.14595
R2738 VTAIL.n676 VTAIL.n669 8.14595
R2739 VTAIL.n616 VTAIL.n615 8.14595
R2740 VTAIL.n607 VTAIL.n544 8.14595
R2741 VTAIL.n570 VTAIL.n563 8.14595
R2742 VTAIL.n510 VTAIL.n509 8.14595
R2743 VTAIL.n501 VTAIL.n438 8.14595
R2744 VTAIL.n464 VTAIL.n457 8.14595
R2745 VTAIL.n404 VTAIL.n403 8.14595
R2746 VTAIL.n395 VTAIL.n332 8.14595
R2747 VTAIL.n358 VTAIL.n351 8.14595
R2748 VTAIL.n778 VTAIL.n777 7.3702
R2749 VTAIL.n820 VTAIL.n754 7.3702
R2750 VTAIL.n824 VTAIL.n752 7.3702
R2751 VTAIL.n36 VTAIL.n35 7.3702
R2752 VTAIL.n78 VTAIL.n12 7.3702
R2753 VTAIL.n82 VTAIL.n10 7.3702
R2754 VTAIL.n142 VTAIL.n141 7.3702
R2755 VTAIL.n184 VTAIL.n118 7.3702
R2756 VTAIL.n188 VTAIL.n116 7.3702
R2757 VTAIL.n248 VTAIL.n247 7.3702
R2758 VTAIL.n290 VTAIL.n224 7.3702
R2759 VTAIL.n294 VTAIL.n222 7.3702
R2760 VTAIL.n718 VTAIL.n646 7.3702
R2761 VTAIL.n714 VTAIL.n648 7.3702
R2762 VTAIL.n673 VTAIL.n672 7.3702
R2763 VTAIL.n612 VTAIL.n540 7.3702
R2764 VTAIL.n608 VTAIL.n542 7.3702
R2765 VTAIL.n567 VTAIL.n566 7.3702
R2766 VTAIL.n506 VTAIL.n434 7.3702
R2767 VTAIL.n502 VTAIL.n436 7.3702
R2768 VTAIL.n461 VTAIL.n460 7.3702
R2769 VTAIL.n400 VTAIL.n328 7.3702
R2770 VTAIL.n396 VTAIL.n330 7.3702
R2771 VTAIL.n355 VTAIL.n354 7.3702
R2772 VTAIL.n823 VTAIL.n754 6.59444
R2773 VTAIL.n824 VTAIL.n823 6.59444
R2774 VTAIL.n81 VTAIL.n12 6.59444
R2775 VTAIL.n82 VTAIL.n81 6.59444
R2776 VTAIL.n187 VTAIL.n118 6.59444
R2777 VTAIL.n188 VTAIL.n187 6.59444
R2778 VTAIL.n293 VTAIL.n224 6.59444
R2779 VTAIL.n294 VTAIL.n293 6.59444
R2780 VTAIL.n718 VTAIL.n717 6.59444
R2781 VTAIL.n717 VTAIL.n648 6.59444
R2782 VTAIL.n612 VTAIL.n611 6.59444
R2783 VTAIL.n611 VTAIL.n542 6.59444
R2784 VTAIL.n506 VTAIL.n505 6.59444
R2785 VTAIL.n505 VTAIL.n436 6.59444
R2786 VTAIL.n400 VTAIL.n399 6.59444
R2787 VTAIL.n399 VTAIL.n330 6.59444
R2788 VTAIL.n778 VTAIL.n774 5.81868
R2789 VTAIL.n820 VTAIL.n819 5.81868
R2790 VTAIL.n827 VTAIL.n752 5.81868
R2791 VTAIL.n36 VTAIL.n32 5.81868
R2792 VTAIL.n78 VTAIL.n77 5.81868
R2793 VTAIL.n85 VTAIL.n10 5.81868
R2794 VTAIL.n142 VTAIL.n138 5.81868
R2795 VTAIL.n184 VTAIL.n183 5.81868
R2796 VTAIL.n191 VTAIL.n116 5.81868
R2797 VTAIL.n248 VTAIL.n244 5.81868
R2798 VTAIL.n290 VTAIL.n289 5.81868
R2799 VTAIL.n297 VTAIL.n222 5.81868
R2800 VTAIL.n721 VTAIL.n646 5.81868
R2801 VTAIL.n714 VTAIL.n713 5.81868
R2802 VTAIL.n673 VTAIL.n669 5.81868
R2803 VTAIL.n615 VTAIL.n540 5.81868
R2804 VTAIL.n608 VTAIL.n607 5.81868
R2805 VTAIL.n567 VTAIL.n563 5.81868
R2806 VTAIL.n509 VTAIL.n434 5.81868
R2807 VTAIL.n502 VTAIL.n501 5.81868
R2808 VTAIL.n461 VTAIL.n457 5.81868
R2809 VTAIL.n403 VTAIL.n328 5.81868
R2810 VTAIL.n396 VTAIL.n395 5.81868
R2811 VTAIL.n355 VTAIL.n351 5.81868
R2812 VTAIL.n844 VTAIL.n742 5.3904
R2813 VTAIL.n102 VTAIL.n0 5.3904
R2814 VTAIL.n208 VTAIL.n106 5.3904
R2815 VTAIL.n314 VTAIL.n212 5.3904
R2816 VTAIL.n738 VTAIL.n636 5.3904
R2817 VTAIL.n632 VTAIL.n530 5.3904
R2818 VTAIL.n526 VTAIL.n424 5.3904
R2819 VTAIL.n420 VTAIL.n318 5.3904
R2820 VTAIL.n782 VTAIL.n781 5.04292
R2821 VTAIL.n816 VTAIL.n756 5.04292
R2822 VTAIL.n828 VTAIL.n750 5.04292
R2823 VTAIL.n40 VTAIL.n39 5.04292
R2824 VTAIL.n74 VTAIL.n14 5.04292
R2825 VTAIL.n86 VTAIL.n8 5.04292
R2826 VTAIL.n146 VTAIL.n145 5.04292
R2827 VTAIL.n180 VTAIL.n120 5.04292
R2828 VTAIL.n192 VTAIL.n114 5.04292
R2829 VTAIL.n252 VTAIL.n251 5.04292
R2830 VTAIL.n286 VTAIL.n226 5.04292
R2831 VTAIL.n298 VTAIL.n220 5.04292
R2832 VTAIL.n722 VTAIL.n644 5.04292
R2833 VTAIL.n710 VTAIL.n650 5.04292
R2834 VTAIL.n677 VTAIL.n676 5.04292
R2835 VTAIL.n616 VTAIL.n538 5.04292
R2836 VTAIL.n604 VTAIL.n544 5.04292
R2837 VTAIL.n571 VTAIL.n570 5.04292
R2838 VTAIL.n510 VTAIL.n432 5.04292
R2839 VTAIL.n498 VTAIL.n438 5.04292
R2840 VTAIL.n465 VTAIL.n464 5.04292
R2841 VTAIL.n404 VTAIL.n326 5.04292
R2842 VTAIL.n392 VTAIL.n332 5.04292
R2843 VTAIL.n359 VTAIL.n358 5.04292
R2844 VTAIL.n785 VTAIL.n772 4.26717
R2845 VTAIL.n815 VTAIL.n758 4.26717
R2846 VTAIL.n832 VTAIL.n831 4.26717
R2847 VTAIL.n43 VTAIL.n30 4.26717
R2848 VTAIL.n73 VTAIL.n16 4.26717
R2849 VTAIL.n90 VTAIL.n89 4.26717
R2850 VTAIL.n149 VTAIL.n136 4.26717
R2851 VTAIL.n179 VTAIL.n122 4.26717
R2852 VTAIL.n196 VTAIL.n195 4.26717
R2853 VTAIL.n255 VTAIL.n242 4.26717
R2854 VTAIL.n285 VTAIL.n228 4.26717
R2855 VTAIL.n302 VTAIL.n301 4.26717
R2856 VTAIL.n726 VTAIL.n725 4.26717
R2857 VTAIL.n709 VTAIL.n652 4.26717
R2858 VTAIL.n680 VTAIL.n667 4.26717
R2859 VTAIL.n620 VTAIL.n619 4.26717
R2860 VTAIL.n603 VTAIL.n546 4.26717
R2861 VTAIL.n574 VTAIL.n561 4.26717
R2862 VTAIL.n514 VTAIL.n513 4.26717
R2863 VTAIL.n497 VTAIL.n440 4.26717
R2864 VTAIL.n468 VTAIL.n455 4.26717
R2865 VTAIL.n408 VTAIL.n407 4.26717
R2866 VTAIL.n391 VTAIL.n334 4.26717
R2867 VTAIL.n362 VTAIL.n349 4.26717
R2868 VTAIL.n786 VTAIL.n770 3.49141
R2869 VTAIL.n812 VTAIL.n811 3.49141
R2870 VTAIL.n835 VTAIL.n748 3.49141
R2871 VTAIL.n44 VTAIL.n28 3.49141
R2872 VTAIL.n70 VTAIL.n69 3.49141
R2873 VTAIL.n93 VTAIL.n6 3.49141
R2874 VTAIL.n150 VTAIL.n134 3.49141
R2875 VTAIL.n176 VTAIL.n175 3.49141
R2876 VTAIL.n199 VTAIL.n112 3.49141
R2877 VTAIL.n256 VTAIL.n240 3.49141
R2878 VTAIL.n282 VTAIL.n281 3.49141
R2879 VTAIL.n305 VTAIL.n218 3.49141
R2880 VTAIL.n729 VTAIL.n642 3.49141
R2881 VTAIL.n706 VTAIL.n705 3.49141
R2882 VTAIL.n681 VTAIL.n665 3.49141
R2883 VTAIL.n623 VTAIL.n536 3.49141
R2884 VTAIL.n600 VTAIL.n599 3.49141
R2885 VTAIL.n575 VTAIL.n559 3.49141
R2886 VTAIL.n517 VTAIL.n430 3.49141
R2887 VTAIL.n494 VTAIL.n493 3.49141
R2888 VTAIL.n469 VTAIL.n453 3.49141
R2889 VTAIL.n411 VTAIL.n324 3.49141
R2890 VTAIL.n388 VTAIL.n387 3.49141
R2891 VTAIL.n363 VTAIL.n347 3.49141
R2892 VTAIL.n529 VTAIL.n423 3.33671
R2893 VTAIL.n741 VTAIL.n635 3.33671
R2894 VTAIL.n317 VTAIL.n211 3.33671
R2895 VTAIL.n779 VTAIL.n775 2.84303
R2896 VTAIL.n37 VTAIL.n33 2.84303
R2897 VTAIL.n143 VTAIL.n139 2.84303
R2898 VTAIL.n249 VTAIL.n245 2.84303
R2899 VTAIL.n674 VTAIL.n670 2.84303
R2900 VTAIL.n568 VTAIL.n564 2.84303
R2901 VTAIL.n462 VTAIL.n458 2.84303
R2902 VTAIL.n356 VTAIL.n352 2.84303
R2903 VTAIL.n790 VTAIL.n789 2.71565
R2904 VTAIL.n808 VTAIL.n760 2.71565
R2905 VTAIL.n836 VTAIL.n746 2.71565
R2906 VTAIL.n48 VTAIL.n47 2.71565
R2907 VTAIL.n66 VTAIL.n18 2.71565
R2908 VTAIL.n94 VTAIL.n4 2.71565
R2909 VTAIL.n154 VTAIL.n153 2.71565
R2910 VTAIL.n172 VTAIL.n124 2.71565
R2911 VTAIL.n200 VTAIL.n110 2.71565
R2912 VTAIL.n260 VTAIL.n259 2.71565
R2913 VTAIL.n278 VTAIL.n230 2.71565
R2914 VTAIL.n306 VTAIL.n216 2.71565
R2915 VTAIL.n730 VTAIL.n640 2.71565
R2916 VTAIL.n702 VTAIL.n654 2.71565
R2917 VTAIL.n685 VTAIL.n684 2.71565
R2918 VTAIL.n624 VTAIL.n534 2.71565
R2919 VTAIL.n596 VTAIL.n548 2.71565
R2920 VTAIL.n579 VTAIL.n578 2.71565
R2921 VTAIL.n518 VTAIL.n428 2.71565
R2922 VTAIL.n490 VTAIL.n442 2.71565
R2923 VTAIL.n473 VTAIL.n472 2.71565
R2924 VTAIL.n412 VTAIL.n322 2.71565
R2925 VTAIL.n384 VTAIL.n336 2.71565
R2926 VTAIL.n367 VTAIL.n366 2.71565
R2927 VTAIL.n794 VTAIL.n768 1.93989
R2928 VTAIL.n807 VTAIL.n762 1.93989
R2929 VTAIL.n840 VTAIL.n839 1.93989
R2930 VTAIL.n52 VTAIL.n26 1.93989
R2931 VTAIL.n65 VTAIL.n20 1.93989
R2932 VTAIL.n98 VTAIL.n97 1.93989
R2933 VTAIL.n158 VTAIL.n132 1.93989
R2934 VTAIL.n171 VTAIL.n126 1.93989
R2935 VTAIL.n204 VTAIL.n203 1.93989
R2936 VTAIL.n264 VTAIL.n238 1.93989
R2937 VTAIL.n277 VTAIL.n232 1.93989
R2938 VTAIL.n310 VTAIL.n309 1.93989
R2939 VTAIL.n734 VTAIL.n733 1.93989
R2940 VTAIL.n701 VTAIL.n656 1.93989
R2941 VTAIL.n688 VTAIL.n662 1.93989
R2942 VTAIL.n628 VTAIL.n627 1.93989
R2943 VTAIL.n595 VTAIL.n550 1.93989
R2944 VTAIL.n582 VTAIL.n556 1.93989
R2945 VTAIL.n522 VTAIL.n521 1.93989
R2946 VTAIL.n489 VTAIL.n444 1.93989
R2947 VTAIL.n476 VTAIL.n450 1.93989
R2948 VTAIL.n416 VTAIL.n415 1.93989
R2949 VTAIL.n383 VTAIL.n338 1.93989
R2950 VTAIL.n370 VTAIL.n344 1.93989
R2951 VTAIL VTAIL.n105 1.72679
R2952 VTAIL VTAIL.n847 1.61041
R2953 VTAIL.n795 VTAIL.n766 1.16414
R2954 VTAIL.n804 VTAIL.n803 1.16414
R2955 VTAIL.n843 VTAIL.n744 1.16414
R2956 VTAIL.n53 VTAIL.n24 1.16414
R2957 VTAIL.n62 VTAIL.n61 1.16414
R2958 VTAIL.n101 VTAIL.n2 1.16414
R2959 VTAIL.n159 VTAIL.n130 1.16414
R2960 VTAIL.n168 VTAIL.n167 1.16414
R2961 VTAIL.n207 VTAIL.n108 1.16414
R2962 VTAIL.n265 VTAIL.n236 1.16414
R2963 VTAIL.n274 VTAIL.n273 1.16414
R2964 VTAIL.n313 VTAIL.n214 1.16414
R2965 VTAIL.n737 VTAIL.n638 1.16414
R2966 VTAIL.n698 VTAIL.n697 1.16414
R2967 VTAIL.n689 VTAIL.n660 1.16414
R2968 VTAIL.n631 VTAIL.n532 1.16414
R2969 VTAIL.n592 VTAIL.n591 1.16414
R2970 VTAIL.n583 VTAIL.n554 1.16414
R2971 VTAIL.n525 VTAIL.n426 1.16414
R2972 VTAIL.n486 VTAIL.n485 1.16414
R2973 VTAIL.n477 VTAIL.n448 1.16414
R2974 VTAIL.n419 VTAIL.n320 1.16414
R2975 VTAIL.n380 VTAIL.n379 1.16414
R2976 VTAIL.n371 VTAIL.n342 1.16414
R2977 VTAIL.n635 VTAIL.n529 0.470328
R2978 VTAIL.n211 VTAIL.n105 0.470328
R2979 VTAIL.n799 VTAIL.n798 0.388379
R2980 VTAIL.n800 VTAIL.n764 0.388379
R2981 VTAIL.n57 VTAIL.n56 0.388379
R2982 VTAIL.n58 VTAIL.n22 0.388379
R2983 VTAIL.n163 VTAIL.n162 0.388379
R2984 VTAIL.n164 VTAIL.n128 0.388379
R2985 VTAIL.n269 VTAIL.n268 0.388379
R2986 VTAIL.n270 VTAIL.n234 0.388379
R2987 VTAIL.n694 VTAIL.n658 0.388379
R2988 VTAIL.n693 VTAIL.n692 0.388379
R2989 VTAIL.n588 VTAIL.n552 0.388379
R2990 VTAIL.n587 VTAIL.n586 0.388379
R2991 VTAIL.n482 VTAIL.n446 0.388379
R2992 VTAIL.n481 VTAIL.n480 0.388379
R2993 VTAIL.n376 VTAIL.n340 0.388379
R2994 VTAIL.n375 VTAIL.n374 0.388379
R2995 VTAIL.n780 VTAIL.n779 0.155672
R2996 VTAIL.n780 VTAIL.n771 0.155672
R2997 VTAIL.n787 VTAIL.n771 0.155672
R2998 VTAIL.n788 VTAIL.n787 0.155672
R2999 VTAIL.n788 VTAIL.n767 0.155672
R3000 VTAIL.n796 VTAIL.n767 0.155672
R3001 VTAIL.n797 VTAIL.n796 0.155672
R3002 VTAIL.n797 VTAIL.n763 0.155672
R3003 VTAIL.n805 VTAIL.n763 0.155672
R3004 VTAIL.n806 VTAIL.n805 0.155672
R3005 VTAIL.n806 VTAIL.n759 0.155672
R3006 VTAIL.n813 VTAIL.n759 0.155672
R3007 VTAIL.n814 VTAIL.n813 0.155672
R3008 VTAIL.n814 VTAIL.n755 0.155672
R3009 VTAIL.n821 VTAIL.n755 0.155672
R3010 VTAIL.n822 VTAIL.n821 0.155672
R3011 VTAIL.n822 VTAIL.n751 0.155672
R3012 VTAIL.n829 VTAIL.n751 0.155672
R3013 VTAIL.n830 VTAIL.n829 0.155672
R3014 VTAIL.n830 VTAIL.n747 0.155672
R3015 VTAIL.n837 VTAIL.n747 0.155672
R3016 VTAIL.n838 VTAIL.n837 0.155672
R3017 VTAIL.n838 VTAIL.n743 0.155672
R3018 VTAIL.n845 VTAIL.n743 0.155672
R3019 VTAIL.n38 VTAIL.n37 0.155672
R3020 VTAIL.n38 VTAIL.n29 0.155672
R3021 VTAIL.n45 VTAIL.n29 0.155672
R3022 VTAIL.n46 VTAIL.n45 0.155672
R3023 VTAIL.n46 VTAIL.n25 0.155672
R3024 VTAIL.n54 VTAIL.n25 0.155672
R3025 VTAIL.n55 VTAIL.n54 0.155672
R3026 VTAIL.n55 VTAIL.n21 0.155672
R3027 VTAIL.n63 VTAIL.n21 0.155672
R3028 VTAIL.n64 VTAIL.n63 0.155672
R3029 VTAIL.n64 VTAIL.n17 0.155672
R3030 VTAIL.n71 VTAIL.n17 0.155672
R3031 VTAIL.n72 VTAIL.n71 0.155672
R3032 VTAIL.n72 VTAIL.n13 0.155672
R3033 VTAIL.n79 VTAIL.n13 0.155672
R3034 VTAIL.n80 VTAIL.n79 0.155672
R3035 VTAIL.n80 VTAIL.n9 0.155672
R3036 VTAIL.n87 VTAIL.n9 0.155672
R3037 VTAIL.n88 VTAIL.n87 0.155672
R3038 VTAIL.n88 VTAIL.n5 0.155672
R3039 VTAIL.n95 VTAIL.n5 0.155672
R3040 VTAIL.n96 VTAIL.n95 0.155672
R3041 VTAIL.n96 VTAIL.n1 0.155672
R3042 VTAIL.n103 VTAIL.n1 0.155672
R3043 VTAIL.n144 VTAIL.n143 0.155672
R3044 VTAIL.n144 VTAIL.n135 0.155672
R3045 VTAIL.n151 VTAIL.n135 0.155672
R3046 VTAIL.n152 VTAIL.n151 0.155672
R3047 VTAIL.n152 VTAIL.n131 0.155672
R3048 VTAIL.n160 VTAIL.n131 0.155672
R3049 VTAIL.n161 VTAIL.n160 0.155672
R3050 VTAIL.n161 VTAIL.n127 0.155672
R3051 VTAIL.n169 VTAIL.n127 0.155672
R3052 VTAIL.n170 VTAIL.n169 0.155672
R3053 VTAIL.n170 VTAIL.n123 0.155672
R3054 VTAIL.n177 VTAIL.n123 0.155672
R3055 VTAIL.n178 VTAIL.n177 0.155672
R3056 VTAIL.n178 VTAIL.n119 0.155672
R3057 VTAIL.n185 VTAIL.n119 0.155672
R3058 VTAIL.n186 VTAIL.n185 0.155672
R3059 VTAIL.n186 VTAIL.n115 0.155672
R3060 VTAIL.n193 VTAIL.n115 0.155672
R3061 VTAIL.n194 VTAIL.n193 0.155672
R3062 VTAIL.n194 VTAIL.n111 0.155672
R3063 VTAIL.n201 VTAIL.n111 0.155672
R3064 VTAIL.n202 VTAIL.n201 0.155672
R3065 VTAIL.n202 VTAIL.n107 0.155672
R3066 VTAIL.n209 VTAIL.n107 0.155672
R3067 VTAIL.n250 VTAIL.n249 0.155672
R3068 VTAIL.n250 VTAIL.n241 0.155672
R3069 VTAIL.n257 VTAIL.n241 0.155672
R3070 VTAIL.n258 VTAIL.n257 0.155672
R3071 VTAIL.n258 VTAIL.n237 0.155672
R3072 VTAIL.n266 VTAIL.n237 0.155672
R3073 VTAIL.n267 VTAIL.n266 0.155672
R3074 VTAIL.n267 VTAIL.n233 0.155672
R3075 VTAIL.n275 VTAIL.n233 0.155672
R3076 VTAIL.n276 VTAIL.n275 0.155672
R3077 VTAIL.n276 VTAIL.n229 0.155672
R3078 VTAIL.n283 VTAIL.n229 0.155672
R3079 VTAIL.n284 VTAIL.n283 0.155672
R3080 VTAIL.n284 VTAIL.n225 0.155672
R3081 VTAIL.n291 VTAIL.n225 0.155672
R3082 VTAIL.n292 VTAIL.n291 0.155672
R3083 VTAIL.n292 VTAIL.n221 0.155672
R3084 VTAIL.n299 VTAIL.n221 0.155672
R3085 VTAIL.n300 VTAIL.n299 0.155672
R3086 VTAIL.n300 VTAIL.n217 0.155672
R3087 VTAIL.n307 VTAIL.n217 0.155672
R3088 VTAIL.n308 VTAIL.n307 0.155672
R3089 VTAIL.n308 VTAIL.n213 0.155672
R3090 VTAIL.n315 VTAIL.n213 0.155672
R3091 VTAIL.n739 VTAIL.n637 0.155672
R3092 VTAIL.n732 VTAIL.n637 0.155672
R3093 VTAIL.n732 VTAIL.n731 0.155672
R3094 VTAIL.n731 VTAIL.n641 0.155672
R3095 VTAIL.n724 VTAIL.n641 0.155672
R3096 VTAIL.n724 VTAIL.n723 0.155672
R3097 VTAIL.n723 VTAIL.n645 0.155672
R3098 VTAIL.n716 VTAIL.n645 0.155672
R3099 VTAIL.n716 VTAIL.n715 0.155672
R3100 VTAIL.n715 VTAIL.n649 0.155672
R3101 VTAIL.n708 VTAIL.n649 0.155672
R3102 VTAIL.n708 VTAIL.n707 0.155672
R3103 VTAIL.n707 VTAIL.n653 0.155672
R3104 VTAIL.n700 VTAIL.n653 0.155672
R3105 VTAIL.n700 VTAIL.n699 0.155672
R3106 VTAIL.n699 VTAIL.n657 0.155672
R3107 VTAIL.n691 VTAIL.n657 0.155672
R3108 VTAIL.n691 VTAIL.n690 0.155672
R3109 VTAIL.n690 VTAIL.n661 0.155672
R3110 VTAIL.n683 VTAIL.n661 0.155672
R3111 VTAIL.n683 VTAIL.n682 0.155672
R3112 VTAIL.n682 VTAIL.n666 0.155672
R3113 VTAIL.n675 VTAIL.n666 0.155672
R3114 VTAIL.n675 VTAIL.n674 0.155672
R3115 VTAIL.n633 VTAIL.n531 0.155672
R3116 VTAIL.n626 VTAIL.n531 0.155672
R3117 VTAIL.n626 VTAIL.n625 0.155672
R3118 VTAIL.n625 VTAIL.n535 0.155672
R3119 VTAIL.n618 VTAIL.n535 0.155672
R3120 VTAIL.n618 VTAIL.n617 0.155672
R3121 VTAIL.n617 VTAIL.n539 0.155672
R3122 VTAIL.n610 VTAIL.n539 0.155672
R3123 VTAIL.n610 VTAIL.n609 0.155672
R3124 VTAIL.n609 VTAIL.n543 0.155672
R3125 VTAIL.n602 VTAIL.n543 0.155672
R3126 VTAIL.n602 VTAIL.n601 0.155672
R3127 VTAIL.n601 VTAIL.n547 0.155672
R3128 VTAIL.n594 VTAIL.n547 0.155672
R3129 VTAIL.n594 VTAIL.n593 0.155672
R3130 VTAIL.n593 VTAIL.n551 0.155672
R3131 VTAIL.n585 VTAIL.n551 0.155672
R3132 VTAIL.n585 VTAIL.n584 0.155672
R3133 VTAIL.n584 VTAIL.n555 0.155672
R3134 VTAIL.n577 VTAIL.n555 0.155672
R3135 VTAIL.n577 VTAIL.n576 0.155672
R3136 VTAIL.n576 VTAIL.n560 0.155672
R3137 VTAIL.n569 VTAIL.n560 0.155672
R3138 VTAIL.n569 VTAIL.n568 0.155672
R3139 VTAIL.n527 VTAIL.n425 0.155672
R3140 VTAIL.n520 VTAIL.n425 0.155672
R3141 VTAIL.n520 VTAIL.n519 0.155672
R3142 VTAIL.n519 VTAIL.n429 0.155672
R3143 VTAIL.n512 VTAIL.n429 0.155672
R3144 VTAIL.n512 VTAIL.n511 0.155672
R3145 VTAIL.n511 VTAIL.n433 0.155672
R3146 VTAIL.n504 VTAIL.n433 0.155672
R3147 VTAIL.n504 VTAIL.n503 0.155672
R3148 VTAIL.n503 VTAIL.n437 0.155672
R3149 VTAIL.n496 VTAIL.n437 0.155672
R3150 VTAIL.n496 VTAIL.n495 0.155672
R3151 VTAIL.n495 VTAIL.n441 0.155672
R3152 VTAIL.n488 VTAIL.n441 0.155672
R3153 VTAIL.n488 VTAIL.n487 0.155672
R3154 VTAIL.n487 VTAIL.n445 0.155672
R3155 VTAIL.n479 VTAIL.n445 0.155672
R3156 VTAIL.n479 VTAIL.n478 0.155672
R3157 VTAIL.n478 VTAIL.n449 0.155672
R3158 VTAIL.n471 VTAIL.n449 0.155672
R3159 VTAIL.n471 VTAIL.n470 0.155672
R3160 VTAIL.n470 VTAIL.n454 0.155672
R3161 VTAIL.n463 VTAIL.n454 0.155672
R3162 VTAIL.n463 VTAIL.n462 0.155672
R3163 VTAIL.n421 VTAIL.n319 0.155672
R3164 VTAIL.n414 VTAIL.n319 0.155672
R3165 VTAIL.n414 VTAIL.n413 0.155672
R3166 VTAIL.n413 VTAIL.n323 0.155672
R3167 VTAIL.n406 VTAIL.n323 0.155672
R3168 VTAIL.n406 VTAIL.n405 0.155672
R3169 VTAIL.n405 VTAIL.n327 0.155672
R3170 VTAIL.n398 VTAIL.n327 0.155672
R3171 VTAIL.n398 VTAIL.n397 0.155672
R3172 VTAIL.n397 VTAIL.n331 0.155672
R3173 VTAIL.n390 VTAIL.n331 0.155672
R3174 VTAIL.n390 VTAIL.n389 0.155672
R3175 VTAIL.n389 VTAIL.n335 0.155672
R3176 VTAIL.n382 VTAIL.n335 0.155672
R3177 VTAIL.n382 VTAIL.n381 0.155672
R3178 VTAIL.n381 VTAIL.n339 0.155672
R3179 VTAIL.n373 VTAIL.n339 0.155672
R3180 VTAIL.n373 VTAIL.n372 0.155672
R3181 VTAIL.n372 VTAIL.n343 0.155672
R3182 VTAIL.n365 VTAIL.n343 0.155672
R3183 VTAIL.n365 VTAIL.n364 0.155672
R3184 VTAIL.n364 VTAIL.n348 0.155672
R3185 VTAIL.n357 VTAIL.n348 0.155672
R3186 VTAIL.n357 VTAIL.n356 0.155672
R3187 VP.n5 VP.t2 167.32
R3188 VP.n5 VP.t1 166.089
R3189 VP.n19 VP.n18 161.3
R3190 VP.n17 VP.n1 161.3
R3191 VP.n16 VP.n15 161.3
R3192 VP.n14 VP.n2 161.3
R3193 VP.n13 VP.n12 161.3
R3194 VP.n11 VP.n3 161.3
R3195 VP.n10 VP.n9 161.3
R3196 VP.n8 VP.n4 161.3
R3197 VP.n6 VP.t0 132.619
R3198 VP.n0 VP.t3 132.619
R3199 VP.n7 VP.n6 81.1466
R3200 VP.n20 VP.n0 81.1466
R3201 VP.n7 VP.n5 57.0663
R3202 VP.n12 VP.n2 56.5617
R3203 VP.n10 VP.n4 24.5923
R3204 VP.n11 VP.n10 24.5923
R3205 VP.n12 VP.n11 24.5923
R3206 VP.n16 VP.n2 24.5923
R3207 VP.n17 VP.n16 24.5923
R3208 VP.n18 VP.n17 24.5923
R3209 VP.n6 VP.n4 9.09948
R3210 VP.n18 VP.n0 9.09948
R3211 VP.n8 VP.n7 0.354861
R3212 VP.n20 VP.n19 0.354861
R3213 VP VP.n20 0.267071
R3214 VP.n9 VP.n8 0.189894
R3215 VP.n9 VP.n3 0.189894
R3216 VP.n13 VP.n3 0.189894
R3217 VP.n14 VP.n13 0.189894
R3218 VP.n15 VP.n14 0.189894
R3219 VP.n15 VP.n1 0.189894
R3220 VP.n19 VP.n1 0.189894
R3221 VDD1 VDD1.n1 114.347
R3222 VDD1 VDD1.n0 63.3629
R3223 VDD1.n0 VDD1.t1 1.01693
R3224 VDD1.n0 VDD1.t2 1.01693
R3225 VDD1.n1 VDD1.t3 1.01693
R3226 VDD1.n1 VDD1.t0 1.01693
C0 VN VP 8.24953f
C1 VN VTAIL 7.588799f
C2 VTAIL VP 7.60291f
C3 VN VDD1 0.150334f
C4 VP VDD1 8.191171f
C5 VTAIL VDD1 7.24719f
C6 VN VDD2 7.88787f
C7 VP VDD2 0.454604f
C8 VTAIL VDD2 7.307701f
C9 VDD1 VDD2 1.252f
C10 VDD2 B 4.885053f
C11 VDD1 B 10.092211f
C12 VTAIL B 15.139033f
C13 VN B 13.095931f
C14 VP B 11.438688f
C15 VDD1.t1 B 0.412331f
C16 VDD1.t2 B 0.412331f
C17 VDD1.n0 B 3.77727f
C18 VDD1.t3 B 0.412331f
C19 VDD1.t0 B 0.412331f
C20 VDD1.n1 B 4.79915f
C21 VP.t3 B 3.72993f
C22 VP.n0 B 1.35789f
C23 VP.n1 B 0.019637f
C24 VP.n2 B 0.028545f
C25 VP.n3 B 0.019637f
C26 VP.n4 B 0.025089f
C27 VP.t2 B 4.02778f
C28 VP.t1 B 4.01763f
C29 VP.n5 B 3.89818f
C30 VP.t0 B 3.72993f
C31 VP.n6 B 1.35789f
C32 VP.n7 B 1.35246f
C33 VP.n8 B 0.031688f
C34 VP.n9 B 0.019637f
C35 VP.n10 B 0.036414f
C36 VP.n11 B 0.036414f
C37 VP.n12 B 0.028545f
C38 VP.n13 B 0.019637f
C39 VP.n14 B 0.019637f
C40 VP.n15 B 0.019637f
C41 VP.n16 B 0.036414f
C42 VP.n17 B 0.036414f
C43 VP.n18 B 0.025089f
C44 VP.n19 B 0.031688f
C45 VP.n20 B 0.053706f
C46 VTAIL.n0 B 0.021207f
C47 VTAIL.n1 B 0.015445f
C48 VTAIL.n2 B 0.008299f
C49 VTAIL.n3 B 0.019617f
C50 VTAIL.n4 B 0.008788f
C51 VTAIL.n5 B 0.015445f
C52 VTAIL.n6 B 0.008299f
C53 VTAIL.n7 B 0.019617f
C54 VTAIL.n8 B 0.008788f
C55 VTAIL.n9 B 0.015445f
C56 VTAIL.n10 B 0.008299f
C57 VTAIL.n11 B 0.019617f
C58 VTAIL.n12 B 0.008788f
C59 VTAIL.n13 B 0.015445f
C60 VTAIL.n14 B 0.008299f
C61 VTAIL.n15 B 0.019617f
C62 VTAIL.n16 B 0.008788f
C63 VTAIL.n17 B 0.015445f
C64 VTAIL.n18 B 0.008299f
C65 VTAIL.n19 B 0.019617f
C66 VTAIL.n20 B 0.008788f
C67 VTAIL.n21 B 0.015445f
C68 VTAIL.n22 B 0.008299f
C69 VTAIL.n23 B 0.019617f
C70 VTAIL.n24 B 0.008788f
C71 VTAIL.n25 B 0.015445f
C72 VTAIL.n26 B 0.008299f
C73 VTAIL.n27 B 0.019617f
C74 VTAIL.n28 B 0.008788f
C75 VTAIL.n29 B 0.015445f
C76 VTAIL.n30 B 0.008299f
C77 VTAIL.n31 B 0.019617f
C78 VTAIL.n32 B 0.008788f
C79 VTAIL.n33 B 0.155709f
C80 VTAIL.t7 B 0.033754f
C81 VTAIL.n34 B 0.014713f
C82 VTAIL.n35 B 0.013868f
C83 VTAIL.n36 B 0.008299f
C84 VTAIL.n37 B 1.29302f
C85 VTAIL.n38 B 0.015445f
C86 VTAIL.n39 B 0.008299f
C87 VTAIL.n40 B 0.008788f
C88 VTAIL.n41 B 0.019617f
C89 VTAIL.n42 B 0.019617f
C90 VTAIL.n43 B 0.008788f
C91 VTAIL.n44 B 0.008299f
C92 VTAIL.n45 B 0.015445f
C93 VTAIL.n46 B 0.015445f
C94 VTAIL.n47 B 0.008299f
C95 VTAIL.n48 B 0.008788f
C96 VTAIL.n49 B 0.019617f
C97 VTAIL.n50 B 0.019617f
C98 VTAIL.n51 B 0.019617f
C99 VTAIL.n52 B 0.008788f
C100 VTAIL.n53 B 0.008299f
C101 VTAIL.n54 B 0.015445f
C102 VTAIL.n55 B 0.015445f
C103 VTAIL.n56 B 0.008299f
C104 VTAIL.n57 B 0.008544f
C105 VTAIL.n58 B 0.008544f
C106 VTAIL.n59 B 0.019617f
C107 VTAIL.n60 B 0.019617f
C108 VTAIL.n61 B 0.008788f
C109 VTAIL.n62 B 0.008299f
C110 VTAIL.n63 B 0.015445f
C111 VTAIL.n64 B 0.015445f
C112 VTAIL.n65 B 0.008299f
C113 VTAIL.n66 B 0.008788f
C114 VTAIL.n67 B 0.019617f
C115 VTAIL.n68 B 0.019617f
C116 VTAIL.n69 B 0.008788f
C117 VTAIL.n70 B 0.008299f
C118 VTAIL.n71 B 0.015445f
C119 VTAIL.n72 B 0.015445f
C120 VTAIL.n73 B 0.008299f
C121 VTAIL.n74 B 0.008788f
C122 VTAIL.n75 B 0.019617f
C123 VTAIL.n76 B 0.019617f
C124 VTAIL.n77 B 0.008788f
C125 VTAIL.n78 B 0.008299f
C126 VTAIL.n79 B 0.015445f
C127 VTAIL.n80 B 0.015445f
C128 VTAIL.n81 B 0.008299f
C129 VTAIL.n82 B 0.008788f
C130 VTAIL.n83 B 0.019617f
C131 VTAIL.n84 B 0.019617f
C132 VTAIL.n85 B 0.008788f
C133 VTAIL.n86 B 0.008299f
C134 VTAIL.n87 B 0.015445f
C135 VTAIL.n88 B 0.015445f
C136 VTAIL.n89 B 0.008299f
C137 VTAIL.n90 B 0.008788f
C138 VTAIL.n91 B 0.019617f
C139 VTAIL.n92 B 0.019617f
C140 VTAIL.n93 B 0.008788f
C141 VTAIL.n94 B 0.008299f
C142 VTAIL.n95 B 0.015445f
C143 VTAIL.n96 B 0.015445f
C144 VTAIL.n97 B 0.008299f
C145 VTAIL.n98 B 0.008788f
C146 VTAIL.n99 B 0.019617f
C147 VTAIL.n100 B 0.040235f
C148 VTAIL.n101 B 0.008788f
C149 VTAIL.n102 B 0.016228f
C150 VTAIL.n103 B 0.039076f
C151 VTAIL.n104 B 0.041657f
C152 VTAIL.n105 B 0.124395f
C153 VTAIL.n106 B 0.021207f
C154 VTAIL.n107 B 0.015445f
C155 VTAIL.n108 B 0.008299f
C156 VTAIL.n109 B 0.019617f
C157 VTAIL.n110 B 0.008788f
C158 VTAIL.n111 B 0.015445f
C159 VTAIL.n112 B 0.008299f
C160 VTAIL.n113 B 0.019617f
C161 VTAIL.n114 B 0.008788f
C162 VTAIL.n115 B 0.015445f
C163 VTAIL.n116 B 0.008299f
C164 VTAIL.n117 B 0.019617f
C165 VTAIL.n118 B 0.008788f
C166 VTAIL.n119 B 0.015445f
C167 VTAIL.n120 B 0.008299f
C168 VTAIL.n121 B 0.019617f
C169 VTAIL.n122 B 0.008788f
C170 VTAIL.n123 B 0.015445f
C171 VTAIL.n124 B 0.008299f
C172 VTAIL.n125 B 0.019617f
C173 VTAIL.n126 B 0.008788f
C174 VTAIL.n127 B 0.015445f
C175 VTAIL.n128 B 0.008299f
C176 VTAIL.n129 B 0.019617f
C177 VTAIL.n130 B 0.008788f
C178 VTAIL.n131 B 0.015445f
C179 VTAIL.n132 B 0.008299f
C180 VTAIL.n133 B 0.019617f
C181 VTAIL.n134 B 0.008788f
C182 VTAIL.n135 B 0.015445f
C183 VTAIL.n136 B 0.008299f
C184 VTAIL.n137 B 0.019617f
C185 VTAIL.n138 B 0.008788f
C186 VTAIL.n139 B 0.155709f
C187 VTAIL.t1 B 0.033754f
C188 VTAIL.n140 B 0.014713f
C189 VTAIL.n141 B 0.013868f
C190 VTAIL.n142 B 0.008299f
C191 VTAIL.n143 B 1.29302f
C192 VTAIL.n144 B 0.015445f
C193 VTAIL.n145 B 0.008299f
C194 VTAIL.n146 B 0.008788f
C195 VTAIL.n147 B 0.019617f
C196 VTAIL.n148 B 0.019617f
C197 VTAIL.n149 B 0.008788f
C198 VTAIL.n150 B 0.008299f
C199 VTAIL.n151 B 0.015445f
C200 VTAIL.n152 B 0.015445f
C201 VTAIL.n153 B 0.008299f
C202 VTAIL.n154 B 0.008788f
C203 VTAIL.n155 B 0.019617f
C204 VTAIL.n156 B 0.019617f
C205 VTAIL.n157 B 0.019617f
C206 VTAIL.n158 B 0.008788f
C207 VTAIL.n159 B 0.008299f
C208 VTAIL.n160 B 0.015445f
C209 VTAIL.n161 B 0.015445f
C210 VTAIL.n162 B 0.008299f
C211 VTAIL.n163 B 0.008544f
C212 VTAIL.n164 B 0.008544f
C213 VTAIL.n165 B 0.019617f
C214 VTAIL.n166 B 0.019617f
C215 VTAIL.n167 B 0.008788f
C216 VTAIL.n168 B 0.008299f
C217 VTAIL.n169 B 0.015445f
C218 VTAIL.n170 B 0.015445f
C219 VTAIL.n171 B 0.008299f
C220 VTAIL.n172 B 0.008788f
C221 VTAIL.n173 B 0.019617f
C222 VTAIL.n174 B 0.019617f
C223 VTAIL.n175 B 0.008788f
C224 VTAIL.n176 B 0.008299f
C225 VTAIL.n177 B 0.015445f
C226 VTAIL.n178 B 0.015445f
C227 VTAIL.n179 B 0.008299f
C228 VTAIL.n180 B 0.008788f
C229 VTAIL.n181 B 0.019617f
C230 VTAIL.n182 B 0.019617f
C231 VTAIL.n183 B 0.008788f
C232 VTAIL.n184 B 0.008299f
C233 VTAIL.n185 B 0.015445f
C234 VTAIL.n186 B 0.015445f
C235 VTAIL.n187 B 0.008299f
C236 VTAIL.n188 B 0.008788f
C237 VTAIL.n189 B 0.019617f
C238 VTAIL.n190 B 0.019617f
C239 VTAIL.n191 B 0.008788f
C240 VTAIL.n192 B 0.008299f
C241 VTAIL.n193 B 0.015445f
C242 VTAIL.n194 B 0.015445f
C243 VTAIL.n195 B 0.008299f
C244 VTAIL.n196 B 0.008788f
C245 VTAIL.n197 B 0.019617f
C246 VTAIL.n198 B 0.019617f
C247 VTAIL.n199 B 0.008788f
C248 VTAIL.n200 B 0.008299f
C249 VTAIL.n201 B 0.015445f
C250 VTAIL.n202 B 0.015445f
C251 VTAIL.n203 B 0.008299f
C252 VTAIL.n204 B 0.008788f
C253 VTAIL.n205 B 0.019617f
C254 VTAIL.n206 B 0.040235f
C255 VTAIL.n207 B 0.008788f
C256 VTAIL.n208 B 0.016228f
C257 VTAIL.n209 B 0.039076f
C258 VTAIL.n210 B 0.041657f
C259 VTAIL.n211 B 0.204515f
C260 VTAIL.n212 B 0.021207f
C261 VTAIL.n213 B 0.015445f
C262 VTAIL.n214 B 0.008299f
C263 VTAIL.n215 B 0.019617f
C264 VTAIL.n216 B 0.008788f
C265 VTAIL.n217 B 0.015445f
C266 VTAIL.n218 B 0.008299f
C267 VTAIL.n219 B 0.019617f
C268 VTAIL.n220 B 0.008788f
C269 VTAIL.n221 B 0.015445f
C270 VTAIL.n222 B 0.008299f
C271 VTAIL.n223 B 0.019617f
C272 VTAIL.n224 B 0.008788f
C273 VTAIL.n225 B 0.015445f
C274 VTAIL.n226 B 0.008299f
C275 VTAIL.n227 B 0.019617f
C276 VTAIL.n228 B 0.008788f
C277 VTAIL.n229 B 0.015445f
C278 VTAIL.n230 B 0.008299f
C279 VTAIL.n231 B 0.019617f
C280 VTAIL.n232 B 0.008788f
C281 VTAIL.n233 B 0.015445f
C282 VTAIL.n234 B 0.008299f
C283 VTAIL.n235 B 0.019617f
C284 VTAIL.n236 B 0.008788f
C285 VTAIL.n237 B 0.015445f
C286 VTAIL.n238 B 0.008299f
C287 VTAIL.n239 B 0.019617f
C288 VTAIL.n240 B 0.008788f
C289 VTAIL.n241 B 0.015445f
C290 VTAIL.n242 B 0.008299f
C291 VTAIL.n243 B 0.019617f
C292 VTAIL.n244 B 0.008788f
C293 VTAIL.n245 B 0.155709f
C294 VTAIL.t3 B 0.033754f
C295 VTAIL.n246 B 0.014713f
C296 VTAIL.n247 B 0.013868f
C297 VTAIL.n248 B 0.008299f
C298 VTAIL.n249 B 1.29302f
C299 VTAIL.n250 B 0.015445f
C300 VTAIL.n251 B 0.008299f
C301 VTAIL.n252 B 0.008788f
C302 VTAIL.n253 B 0.019617f
C303 VTAIL.n254 B 0.019617f
C304 VTAIL.n255 B 0.008788f
C305 VTAIL.n256 B 0.008299f
C306 VTAIL.n257 B 0.015445f
C307 VTAIL.n258 B 0.015445f
C308 VTAIL.n259 B 0.008299f
C309 VTAIL.n260 B 0.008788f
C310 VTAIL.n261 B 0.019617f
C311 VTAIL.n262 B 0.019617f
C312 VTAIL.n263 B 0.019617f
C313 VTAIL.n264 B 0.008788f
C314 VTAIL.n265 B 0.008299f
C315 VTAIL.n266 B 0.015445f
C316 VTAIL.n267 B 0.015445f
C317 VTAIL.n268 B 0.008299f
C318 VTAIL.n269 B 0.008544f
C319 VTAIL.n270 B 0.008544f
C320 VTAIL.n271 B 0.019617f
C321 VTAIL.n272 B 0.019617f
C322 VTAIL.n273 B 0.008788f
C323 VTAIL.n274 B 0.008299f
C324 VTAIL.n275 B 0.015445f
C325 VTAIL.n276 B 0.015445f
C326 VTAIL.n277 B 0.008299f
C327 VTAIL.n278 B 0.008788f
C328 VTAIL.n279 B 0.019617f
C329 VTAIL.n280 B 0.019617f
C330 VTAIL.n281 B 0.008788f
C331 VTAIL.n282 B 0.008299f
C332 VTAIL.n283 B 0.015445f
C333 VTAIL.n284 B 0.015445f
C334 VTAIL.n285 B 0.008299f
C335 VTAIL.n286 B 0.008788f
C336 VTAIL.n287 B 0.019617f
C337 VTAIL.n288 B 0.019617f
C338 VTAIL.n289 B 0.008788f
C339 VTAIL.n290 B 0.008299f
C340 VTAIL.n291 B 0.015445f
C341 VTAIL.n292 B 0.015445f
C342 VTAIL.n293 B 0.008299f
C343 VTAIL.n294 B 0.008788f
C344 VTAIL.n295 B 0.019617f
C345 VTAIL.n296 B 0.019617f
C346 VTAIL.n297 B 0.008788f
C347 VTAIL.n298 B 0.008299f
C348 VTAIL.n299 B 0.015445f
C349 VTAIL.n300 B 0.015445f
C350 VTAIL.n301 B 0.008299f
C351 VTAIL.n302 B 0.008788f
C352 VTAIL.n303 B 0.019617f
C353 VTAIL.n304 B 0.019617f
C354 VTAIL.n305 B 0.008788f
C355 VTAIL.n306 B 0.008299f
C356 VTAIL.n307 B 0.015445f
C357 VTAIL.n308 B 0.015445f
C358 VTAIL.n309 B 0.008299f
C359 VTAIL.n310 B 0.008788f
C360 VTAIL.n311 B 0.019617f
C361 VTAIL.n312 B 0.040235f
C362 VTAIL.n313 B 0.008788f
C363 VTAIL.n314 B 0.016228f
C364 VTAIL.n315 B 0.039076f
C365 VTAIL.n316 B 0.041657f
C366 VTAIL.n317 B 1.39271f
C367 VTAIL.n318 B 0.021207f
C368 VTAIL.n319 B 0.015445f
C369 VTAIL.n320 B 0.008299f
C370 VTAIL.n321 B 0.019617f
C371 VTAIL.n322 B 0.008788f
C372 VTAIL.n323 B 0.015445f
C373 VTAIL.n324 B 0.008299f
C374 VTAIL.n325 B 0.019617f
C375 VTAIL.n326 B 0.008788f
C376 VTAIL.n327 B 0.015445f
C377 VTAIL.n328 B 0.008299f
C378 VTAIL.n329 B 0.019617f
C379 VTAIL.n330 B 0.008788f
C380 VTAIL.n331 B 0.015445f
C381 VTAIL.n332 B 0.008299f
C382 VTAIL.n333 B 0.019617f
C383 VTAIL.n334 B 0.008788f
C384 VTAIL.n335 B 0.015445f
C385 VTAIL.n336 B 0.008299f
C386 VTAIL.n337 B 0.019617f
C387 VTAIL.n338 B 0.008788f
C388 VTAIL.n339 B 0.015445f
C389 VTAIL.n340 B 0.008299f
C390 VTAIL.n341 B 0.019617f
C391 VTAIL.n342 B 0.008788f
C392 VTAIL.n343 B 0.015445f
C393 VTAIL.n344 B 0.008299f
C394 VTAIL.n345 B 0.019617f
C395 VTAIL.n346 B 0.019617f
C396 VTAIL.n347 B 0.008788f
C397 VTAIL.n348 B 0.015445f
C398 VTAIL.n349 B 0.008299f
C399 VTAIL.n350 B 0.019617f
C400 VTAIL.n351 B 0.008788f
C401 VTAIL.n352 B 0.155709f
C402 VTAIL.t5 B 0.033754f
C403 VTAIL.n353 B 0.014713f
C404 VTAIL.n354 B 0.013868f
C405 VTAIL.n355 B 0.008299f
C406 VTAIL.n356 B 1.29302f
C407 VTAIL.n357 B 0.015445f
C408 VTAIL.n358 B 0.008299f
C409 VTAIL.n359 B 0.008788f
C410 VTAIL.n360 B 0.019617f
C411 VTAIL.n361 B 0.019617f
C412 VTAIL.n362 B 0.008788f
C413 VTAIL.n363 B 0.008299f
C414 VTAIL.n364 B 0.015445f
C415 VTAIL.n365 B 0.015445f
C416 VTAIL.n366 B 0.008299f
C417 VTAIL.n367 B 0.008788f
C418 VTAIL.n368 B 0.019617f
C419 VTAIL.n369 B 0.019617f
C420 VTAIL.n370 B 0.008788f
C421 VTAIL.n371 B 0.008299f
C422 VTAIL.n372 B 0.015445f
C423 VTAIL.n373 B 0.015445f
C424 VTAIL.n374 B 0.008299f
C425 VTAIL.n375 B 0.008544f
C426 VTAIL.n376 B 0.008544f
C427 VTAIL.n377 B 0.019617f
C428 VTAIL.n378 B 0.019617f
C429 VTAIL.n379 B 0.008788f
C430 VTAIL.n380 B 0.008299f
C431 VTAIL.n381 B 0.015445f
C432 VTAIL.n382 B 0.015445f
C433 VTAIL.n383 B 0.008299f
C434 VTAIL.n384 B 0.008788f
C435 VTAIL.n385 B 0.019617f
C436 VTAIL.n386 B 0.019617f
C437 VTAIL.n387 B 0.008788f
C438 VTAIL.n388 B 0.008299f
C439 VTAIL.n389 B 0.015445f
C440 VTAIL.n390 B 0.015445f
C441 VTAIL.n391 B 0.008299f
C442 VTAIL.n392 B 0.008788f
C443 VTAIL.n393 B 0.019617f
C444 VTAIL.n394 B 0.019617f
C445 VTAIL.n395 B 0.008788f
C446 VTAIL.n396 B 0.008299f
C447 VTAIL.n397 B 0.015445f
C448 VTAIL.n398 B 0.015445f
C449 VTAIL.n399 B 0.008299f
C450 VTAIL.n400 B 0.008788f
C451 VTAIL.n401 B 0.019617f
C452 VTAIL.n402 B 0.019617f
C453 VTAIL.n403 B 0.008788f
C454 VTAIL.n404 B 0.008299f
C455 VTAIL.n405 B 0.015445f
C456 VTAIL.n406 B 0.015445f
C457 VTAIL.n407 B 0.008299f
C458 VTAIL.n408 B 0.008788f
C459 VTAIL.n409 B 0.019617f
C460 VTAIL.n410 B 0.019617f
C461 VTAIL.n411 B 0.008788f
C462 VTAIL.n412 B 0.008299f
C463 VTAIL.n413 B 0.015445f
C464 VTAIL.n414 B 0.015445f
C465 VTAIL.n415 B 0.008299f
C466 VTAIL.n416 B 0.008788f
C467 VTAIL.n417 B 0.019617f
C468 VTAIL.n418 B 0.040235f
C469 VTAIL.n419 B 0.008788f
C470 VTAIL.n420 B 0.016228f
C471 VTAIL.n421 B 0.039076f
C472 VTAIL.n422 B 0.041657f
C473 VTAIL.n423 B 1.39271f
C474 VTAIL.n424 B 0.021207f
C475 VTAIL.n425 B 0.015445f
C476 VTAIL.n426 B 0.008299f
C477 VTAIL.n427 B 0.019617f
C478 VTAIL.n428 B 0.008788f
C479 VTAIL.n429 B 0.015445f
C480 VTAIL.n430 B 0.008299f
C481 VTAIL.n431 B 0.019617f
C482 VTAIL.n432 B 0.008788f
C483 VTAIL.n433 B 0.015445f
C484 VTAIL.n434 B 0.008299f
C485 VTAIL.n435 B 0.019617f
C486 VTAIL.n436 B 0.008788f
C487 VTAIL.n437 B 0.015445f
C488 VTAIL.n438 B 0.008299f
C489 VTAIL.n439 B 0.019617f
C490 VTAIL.n440 B 0.008788f
C491 VTAIL.n441 B 0.015445f
C492 VTAIL.n442 B 0.008299f
C493 VTAIL.n443 B 0.019617f
C494 VTAIL.n444 B 0.008788f
C495 VTAIL.n445 B 0.015445f
C496 VTAIL.n446 B 0.008299f
C497 VTAIL.n447 B 0.019617f
C498 VTAIL.n448 B 0.008788f
C499 VTAIL.n449 B 0.015445f
C500 VTAIL.n450 B 0.008299f
C501 VTAIL.n451 B 0.019617f
C502 VTAIL.n452 B 0.019617f
C503 VTAIL.n453 B 0.008788f
C504 VTAIL.n454 B 0.015445f
C505 VTAIL.n455 B 0.008299f
C506 VTAIL.n456 B 0.019617f
C507 VTAIL.n457 B 0.008788f
C508 VTAIL.n458 B 0.155709f
C509 VTAIL.t6 B 0.033754f
C510 VTAIL.n459 B 0.014713f
C511 VTAIL.n460 B 0.013868f
C512 VTAIL.n461 B 0.008299f
C513 VTAIL.n462 B 1.29302f
C514 VTAIL.n463 B 0.015445f
C515 VTAIL.n464 B 0.008299f
C516 VTAIL.n465 B 0.008788f
C517 VTAIL.n466 B 0.019617f
C518 VTAIL.n467 B 0.019617f
C519 VTAIL.n468 B 0.008788f
C520 VTAIL.n469 B 0.008299f
C521 VTAIL.n470 B 0.015445f
C522 VTAIL.n471 B 0.015445f
C523 VTAIL.n472 B 0.008299f
C524 VTAIL.n473 B 0.008788f
C525 VTAIL.n474 B 0.019617f
C526 VTAIL.n475 B 0.019617f
C527 VTAIL.n476 B 0.008788f
C528 VTAIL.n477 B 0.008299f
C529 VTAIL.n478 B 0.015445f
C530 VTAIL.n479 B 0.015445f
C531 VTAIL.n480 B 0.008299f
C532 VTAIL.n481 B 0.008544f
C533 VTAIL.n482 B 0.008544f
C534 VTAIL.n483 B 0.019617f
C535 VTAIL.n484 B 0.019617f
C536 VTAIL.n485 B 0.008788f
C537 VTAIL.n486 B 0.008299f
C538 VTAIL.n487 B 0.015445f
C539 VTAIL.n488 B 0.015445f
C540 VTAIL.n489 B 0.008299f
C541 VTAIL.n490 B 0.008788f
C542 VTAIL.n491 B 0.019617f
C543 VTAIL.n492 B 0.019617f
C544 VTAIL.n493 B 0.008788f
C545 VTAIL.n494 B 0.008299f
C546 VTAIL.n495 B 0.015445f
C547 VTAIL.n496 B 0.015445f
C548 VTAIL.n497 B 0.008299f
C549 VTAIL.n498 B 0.008788f
C550 VTAIL.n499 B 0.019617f
C551 VTAIL.n500 B 0.019617f
C552 VTAIL.n501 B 0.008788f
C553 VTAIL.n502 B 0.008299f
C554 VTAIL.n503 B 0.015445f
C555 VTAIL.n504 B 0.015445f
C556 VTAIL.n505 B 0.008299f
C557 VTAIL.n506 B 0.008788f
C558 VTAIL.n507 B 0.019617f
C559 VTAIL.n508 B 0.019617f
C560 VTAIL.n509 B 0.008788f
C561 VTAIL.n510 B 0.008299f
C562 VTAIL.n511 B 0.015445f
C563 VTAIL.n512 B 0.015445f
C564 VTAIL.n513 B 0.008299f
C565 VTAIL.n514 B 0.008788f
C566 VTAIL.n515 B 0.019617f
C567 VTAIL.n516 B 0.019617f
C568 VTAIL.n517 B 0.008788f
C569 VTAIL.n518 B 0.008299f
C570 VTAIL.n519 B 0.015445f
C571 VTAIL.n520 B 0.015445f
C572 VTAIL.n521 B 0.008299f
C573 VTAIL.n522 B 0.008788f
C574 VTAIL.n523 B 0.019617f
C575 VTAIL.n524 B 0.040235f
C576 VTAIL.n525 B 0.008788f
C577 VTAIL.n526 B 0.016228f
C578 VTAIL.n527 B 0.039076f
C579 VTAIL.n528 B 0.041657f
C580 VTAIL.n529 B 0.204515f
C581 VTAIL.n530 B 0.021207f
C582 VTAIL.n531 B 0.015445f
C583 VTAIL.n532 B 0.008299f
C584 VTAIL.n533 B 0.019617f
C585 VTAIL.n534 B 0.008788f
C586 VTAIL.n535 B 0.015445f
C587 VTAIL.n536 B 0.008299f
C588 VTAIL.n537 B 0.019617f
C589 VTAIL.n538 B 0.008788f
C590 VTAIL.n539 B 0.015445f
C591 VTAIL.n540 B 0.008299f
C592 VTAIL.n541 B 0.019617f
C593 VTAIL.n542 B 0.008788f
C594 VTAIL.n543 B 0.015445f
C595 VTAIL.n544 B 0.008299f
C596 VTAIL.n545 B 0.019617f
C597 VTAIL.n546 B 0.008788f
C598 VTAIL.n547 B 0.015445f
C599 VTAIL.n548 B 0.008299f
C600 VTAIL.n549 B 0.019617f
C601 VTAIL.n550 B 0.008788f
C602 VTAIL.n551 B 0.015445f
C603 VTAIL.n552 B 0.008299f
C604 VTAIL.n553 B 0.019617f
C605 VTAIL.n554 B 0.008788f
C606 VTAIL.n555 B 0.015445f
C607 VTAIL.n556 B 0.008299f
C608 VTAIL.n557 B 0.019617f
C609 VTAIL.n558 B 0.019617f
C610 VTAIL.n559 B 0.008788f
C611 VTAIL.n560 B 0.015445f
C612 VTAIL.n561 B 0.008299f
C613 VTAIL.n562 B 0.019617f
C614 VTAIL.n563 B 0.008788f
C615 VTAIL.n564 B 0.155709f
C616 VTAIL.t0 B 0.033754f
C617 VTAIL.n565 B 0.014713f
C618 VTAIL.n566 B 0.013868f
C619 VTAIL.n567 B 0.008299f
C620 VTAIL.n568 B 1.29302f
C621 VTAIL.n569 B 0.015445f
C622 VTAIL.n570 B 0.008299f
C623 VTAIL.n571 B 0.008788f
C624 VTAIL.n572 B 0.019617f
C625 VTAIL.n573 B 0.019617f
C626 VTAIL.n574 B 0.008788f
C627 VTAIL.n575 B 0.008299f
C628 VTAIL.n576 B 0.015445f
C629 VTAIL.n577 B 0.015445f
C630 VTAIL.n578 B 0.008299f
C631 VTAIL.n579 B 0.008788f
C632 VTAIL.n580 B 0.019617f
C633 VTAIL.n581 B 0.019617f
C634 VTAIL.n582 B 0.008788f
C635 VTAIL.n583 B 0.008299f
C636 VTAIL.n584 B 0.015445f
C637 VTAIL.n585 B 0.015445f
C638 VTAIL.n586 B 0.008299f
C639 VTAIL.n587 B 0.008544f
C640 VTAIL.n588 B 0.008544f
C641 VTAIL.n589 B 0.019617f
C642 VTAIL.n590 B 0.019617f
C643 VTAIL.n591 B 0.008788f
C644 VTAIL.n592 B 0.008299f
C645 VTAIL.n593 B 0.015445f
C646 VTAIL.n594 B 0.015445f
C647 VTAIL.n595 B 0.008299f
C648 VTAIL.n596 B 0.008788f
C649 VTAIL.n597 B 0.019617f
C650 VTAIL.n598 B 0.019617f
C651 VTAIL.n599 B 0.008788f
C652 VTAIL.n600 B 0.008299f
C653 VTAIL.n601 B 0.015445f
C654 VTAIL.n602 B 0.015445f
C655 VTAIL.n603 B 0.008299f
C656 VTAIL.n604 B 0.008788f
C657 VTAIL.n605 B 0.019617f
C658 VTAIL.n606 B 0.019617f
C659 VTAIL.n607 B 0.008788f
C660 VTAIL.n608 B 0.008299f
C661 VTAIL.n609 B 0.015445f
C662 VTAIL.n610 B 0.015445f
C663 VTAIL.n611 B 0.008299f
C664 VTAIL.n612 B 0.008788f
C665 VTAIL.n613 B 0.019617f
C666 VTAIL.n614 B 0.019617f
C667 VTAIL.n615 B 0.008788f
C668 VTAIL.n616 B 0.008299f
C669 VTAIL.n617 B 0.015445f
C670 VTAIL.n618 B 0.015445f
C671 VTAIL.n619 B 0.008299f
C672 VTAIL.n620 B 0.008788f
C673 VTAIL.n621 B 0.019617f
C674 VTAIL.n622 B 0.019617f
C675 VTAIL.n623 B 0.008788f
C676 VTAIL.n624 B 0.008299f
C677 VTAIL.n625 B 0.015445f
C678 VTAIL.n626 B 0.015445f
C679 VTAIL.n627 B 0.008299f
C680 VTAIL.n628 B 0.008788f
C681 VTAIL.n629 B 0.019617f
C682 VTAIL.n630 B 0.040235f
C683 VTAIL.n631 B 0.008788f
C684 VTAIL.n632 B 0.016228f
C685 VTAIL.n633 B 0.039076f
C686 VTAIL.n634 B 0.041657f
C687 VTAIL.n635 B 0.204515f
C688 VTAIL.n636 B 0.021207f
C689 VTAIL.n637 B 0.015445f
C690 VTAIL.n638 B 0.008299f
C691 VTAIL.n639 B 0.019617f
C692 VTAIL.n640 B 0.008788f
C693 VTAIL.n641 B 0.015445f
C694 VTAIL.n642 B 0.008299f
C695 VTAIL.n643 B 0.019617f
C696 VTAIL.n644 B 0.008788f
C697 VTAIL.n645 B 0.015445f
C698 VTAIL.n646 B 0.008299f
C699 VTAIL.n647 B 0.019617f
C700 VTAIL.n648 B 0.008788f
C701 VTAIL.n649 B 0.015445f
C702 VTAIL.n650 B 0.008299f
C703 VTAIL.n651 B 0.019617f
C704 VTAIL.n652 B 0.008788f
C705 VTAIL.n653 B 0.015445f
C706 VTAIL.n654 B 0.008299f
C707 VTAIL.n655 B 0.019617f
C708 VTAIL.n656 B 0.008788f
C709 VTAIL.n657 B 0.015445f
C710 VTAIL.n658 B 0.008299f
C711 VTAIL.n659 B 0.019617f
C712 VTAIL.n660 B 0.008788f
C713 VTAIL.n661 B 0.015445f
C714 VTAIL.n662 B 0.008299f
C715 VTAIL.n663 B 0.019617f
C716 VTAIL.n664 B 0.019617f
C717 VTAIL.n665 B 0.008788f
C718 VTAIL.n666 B 0.015445f
C719 VTAIL.n667 B 0.008299f
C720 VTAIL.n668 B 0.019617f
C721 VTAIL.n669 B 0.008788f
C722 VTAIL.n670 B 0.155709f
C723 VTAIL.t2 B 0.033754f
C724 VTAIL.n671 B 0.014713f
C725 VTAIL.n672 B 0.013868f
C726 VTAIL.n673 B 0.008299f
C727 VTAIL.n674 B 1.29302f
C728 VTAIL.n675 B 0.015445f
C729 VTAIL.n676 B 0.008299f
C730 VTAIL.n677 B 0.008788f
C731 VTAIL.n678 B 0.019617f
C732 VTAIL.n679 B 0.019617f
C733 VTAIL.n680 B 0.008788f
C734 VTAIL.n681 B 0.008299f
C735 VTAIL.n682 B 0.015445f
C736 VTAIL.n683 B 0.015445f
C737 VTAIL.n684 B 0.008299f
C738 VTAIL.n685 B 0.008788f
C739 VTAIL.n686 B 0.019617f
C740 VTAIL.n687 B 0.019617f
C741 VTAIL.n688 B 0.008788f
C742 VTAIL.n689 B 0.008299f
C743 VTAIL.n690 B 0.015445f
C744 VTAIL.n691 B 0.015445f
C745 VTAIL.n692 B 0.008299f
C746 VTAIL.n693 B 0.008544f
C747 VTAIL.n694 B 0.008544f
C748 VTAIL.n695 B 0.019617f
C749 VTAIL.n696 B 0.019617f
C750 VTAIL.n697 B 0.008788f
C751 VTAIL.n698 B 0.008299f
C752 VTAIL.n699 B 0.015445f
C753 VTAIL.n700 B 0.015445f
C754 VTAIL.n701 B 0.008299f
C755 VTAIL.n702 B 0.008788f
C756 VTAIL.n703 B 0.019617f
C757 VTAIL.n704 B 0.019617f
C758 VTAIL.n705 B 0.008788f
C759 VTAIL.n706 B 0.008299f
C760 VTAIL.n707 B 0.015445f
C761 VTAIL.n708 B 0.015445f
C762 VTAIL.n709 B 0.008299f
C763 VTAIL.n710 B 0.008788f
C764 VTAIL.n711 B 0.019617f
C765 VTAIL.n712 B 0.019617f
C766 VTAIL.n713 B 0.008788f
C767 VTAIL.n714 B 0.008299f
C768 VTAIL.n715 B 0.015445f
C769 VTAIL.n716 B 0.015445f
C770 VTAIL.n717 B 0.008299f
C771 VTAIL.n718 B 0.008788f
C772 VTAIL.n719 B 0.019617f
C773 VTAIL.n720 B 0.019617f
C774 VTAIL.n721 B 0.008788f
C775 VTAIL.n722 B 0.008299f
C776 VTAIL.n723 B 0.015445f
C777 VTAIL.n724 B 0.015445f
C778 VTAIL.n725 B 0.008299f
C779 VTAIL.n726 B 0.008788f
C780 VTAIL.n727 B 0.019617f
C781 VTAIL.n728 B 0.019617f
C782 VTAIL.n729 B 0.008788f
C783 VTAIL.n730 B 0.008299f
C784 VTAIL.n731 B 0.015445f
C785 VTAIL.n732 B 0.015445f
C786 VTAIL.n733 B 0.008299f
C787 VTAIL.n734 B 0.008788f
C788 VTAIL.n735 B 0.019617f
C789 VTAIL.n736 B 0.040235f
C790 VTAIL.n737 B 0.008788f
C791 VTAIL.n738 B 0.016228f
C792 VTAIL.n739 B 0.039076f
C793 VTAIL.n740 B 0.041657f
C794 VTAIL.n741 B 1.39271f
C795 VTAIL.n742 B 0.021207f
C796 VTAIL.n743 B 0.015445f
C797 VTAIL.n744 B 0.008299f
C798 VTAIL.n745 B 0.019617f
C799 VTAIL.n746 B 0.008788f
C800 VTAIL.n747 B 0.015445f
C801 VTAIL.n748 B 0.008299f
C802 VTAIL.n749 B 0.019617f
C803 VTAIL.n750 B 0.008788f
C804 VTAIL.n751 B 0.015445f
C805 VTAIL.n752 B 0.008299f
C806 VTAIL.n753 B 0.019617f
C807 VTAIL.n754 B 0.008788f
C808 VTAIL.n755 B 0.015445f
C809 VTAIL.n756 B 0.008299f
C810 VTAIL.n757 B 0.019617f
C811 VTAIL.n758 B 0.008788f
C812 VTAIL.n759 B 0.015445f
C813 VTAIL.n760 B 0.008299f
C814 VTAIL.n761 B 0.019617f
C815 VTAIL.n762 B 0.008788f
C816 VTAIL.n763 B 0.015445f
C817 VTAIL.n764 B 0.008299f
C818 VTAIL.n765 B 0.019617f
C819 VTAIL.n766 B 0.008788f
C820 VTAIL.n767 B 0.015445f
C821 VTAIL.n768 B 0.008299f
C822 VTAIL.n769 B 0.019617f
C823 VTAIL.n770 B 0.008788f
C824 VTAIL.n771 B 0.015445f
C825 VTAIL.n772 B 0.008299f
C826 VTAIL.n773 B 0.019617f
C827 VTAIL.n774 B 0.008788f
C828 VTAIL.n775 B 0.155709f
C829 VTAIL.t4 B 0.033754f
C830 VTAIL.n776 B 0.014713f
C831 VTAIL.n777 B 0.013868f
C832 VTAIL.n778 B 0.008299f
C833 VTAIL.n779 B 1.29302f
C834 VTAIL.n780 B 0.015445f
C835 VTAIL.n781 B 0.008299f
C836 VTAIL.n782 B 0.008788f
C837 VTAIL.n783 B 0.019617f
C838 VTAIL.n784 B 0.019617f
C839 VTAIL.n785 B 0.008788f
C840 VTAIL.n786 B 0.008299f
C841 VTAIL.n787 B 0.015445f
C842 VTAIL.n788 B 0.015445f
C843 VTAIL.n789 B 0.008299f
C844 VTAIL.n790 B 0.008788f
C845 VTAIL.n791 B 0.019617f
C846 VTAIL.n792 B 0.019617f
C847 VTAIL.n793 B 0.019617f
C848 VTAIL.n794 B 0.008788f
C849 VTAIL.n795 B 0.008299f
C850 VTAIL.n796 B 0.015445f
C851 VTAIL.n797 B 0.015445f
C852 VTAIL.n798 B 0.008299f
C853 VTAIL.n799 B 0.008544f
C854 VTAIL.n800 B 0.008544f
C855 VTAIL.n801 B 0.019617f
C856 VTAIL.n802 B 0.019617f
C857 VTAIL.n803 B 0.008788f
C858 VTAIL.n804 B 0.008299f
C859 VTAIL.n805 B 0.015445f
C860 VTAIL.n806 B 0.015445f
C861 VTAIL.n807 B 0.008299f
C862 VTAIL.n808 B 0.008788f
C863 VTAIL.n809 B 0.019617f
C864 VTAIL.n810 B 0.019617f
C865 VTAIL.n811 B 0.008788f
C866 VTAIL.n812 B 0.008299f
C867 VTAIL.n813 B 0.015445f
C868 VTAIL.n814 B 0.015445f
C869 VTAIL.n815 B 0.008299f
C870 VTAIL.n816 B 0.008788f
C871 VTAIL.n817 B 0.019617f
C872 VTAIL.n818 B 0.019617f
C873 VTAIL.n819 B 0.008788f
C874 VTAIL.n820 B 0.008299f
C875 VTAIL.n821 B 0.015445f
C876 VTAIL.n822 B 0.015445f
C877 VTAIL.n823 B 0.008299f
C878 VTAIL.n824 B 0.008788f
C879 VTAIL.n825 B 0.019617f
C880 VTAIL.n826 B 0.019617f
C881 VTAIL.n827 B 0.008788f
C882 VTAIL.n828 B 0.008299f
C883 VTAIL.n829 B 0.015445f
C884 VTAIL.n830 B 0.015445f
C885 VTAIL.n831 B 0.008299f
C886 VTAIL.n832 B 0.008788f
C887 VTAIL.n833 B 0.019617f
C888 VTAIL.n834 B 0.019617f
C889 VTAIL.n835 B 0.008788f
C890 VTAIL.n836 B 0.008299f
C891 VTAIL.n837 B 0.015445f
C892 VTAIL.n838 B 0.015445f
C893 VTAIL.n839 B 0.008299f
C894 VTAIL.n840 B 0.008788f
C895 VTAIL.n841 B 0.019617f
C896 VTAIL.n842 B 0.040235f
C897 VTAIL.n843 B 0.008788f
C898 VTAIL.n844 B 0.016228f
C899 VTAIL.n845 B 0.039076f
C900 VTAIL.n846 B 0.041657f
C901 VTAIL.n847 B 1.30679f
C902 VDD2.t0 B 0.409607f
C903 VDD2.t2 B 0.409607f
C904 VDD2.n0 B 4.73865f
C905 VDD2.t1 B 0.409607f
C906 VDD2.t3 B 0.409607f
C907 VDD2.n1 B 3.75185f
C908 VDD2.n2 B 4.7793f
C909 VN.t3 B 3.96285f
C910 VN.t0 B 3.97287f
C911 VN.n0 B 2.43545f
C912 VN.t1 B 3.97287f
C913 VN.t2 B 3.96285f
C914 VN.n1 B 3.85258f
.ends

