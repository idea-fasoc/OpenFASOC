* NGSPICE file created from diff_pair_sample_0073.ext - technology: sky130A

.subckt diff_pair_sample_0073 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t7 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=3.69
X1 VDD2.t3 VN.t0 VTAIL.t3 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=3.69
X2 VTAIL.t2 VN.t1 VDD2.t2 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=3.69
X3 B.t11 B.t9 B.t10 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=3.69
X4 VDD2.t1 VN.t2 VTAIL.t1 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=3.69
X5 B.t8 B.t6 B.t7 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=3.69
X6 B.t5 B.t3 B.t4 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=3.69
X7 VTAIL.t0 VN.t3 VDD2.t0 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=3.69
X8 VDD1.t2 VP.t1 VTAIL.t5 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=0.55275 pd=3.68 as=1.3065 ps=7.48 w=3.35 l=3.69
X9 VTAIL.t6 VP.t2 VDD1.t1 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=3.69
X10 VTAIL.t4 VP.t3 VDD1.t0 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0.55275 ps=3.68 w=3.35 l=3.69
X11 B.t2 B.t0 B.t1 w_n3382_n1638# sky130_fd_pr__pfet_01v8 ad=1.3065 pd=7.48 as=0 ps=0 w=3.35 l=3.69
R0 VP.n21 VP.n20 161.3
R1 VP.n19 VP.n1 161.3
R2 VP.n18 VP.n17 161.3
R3 VP.n16 VP.n2 161.3
R4 VP.n15 VP.n14 161.3
R5 VP.n13 VP.n3 161.3
R6 VP.n12 VP.n11 161.3
R7 VP.n10 VP.n4 161.3
R8 VP.n9 VP.n8 161.3
R9 VP.n7 VP.n6 89.5781
R10 VP.n22 VP.n0 89.5781
R11 VP.n5 VP.t3 55.084
R12 VP.n5 VP.t0 53.7611
R13 VP.n6 VP.n5 45.017
R14 VP.n14 VP.n13 40.4934
R15 VP.n14 VP.n2 40.4934
R16 VP.n8 VP.n4 24.4675
R17 VP.n12 VP.n4 24.4675
R18 VP.n13 VP.n12 24.4675
R19 VP.n18 VP.n2 24.4675
R20 VP.n19 VP.n18 24.4675
R21 VP.n20 VP.n19 24.4675
R22 VP.n7 VP.t2 21.8799
R23 VP.n0 VP.t1 21.8799
R24 VP.n8 VP.n7 0.48984
R25 VP.n20 VP.n0 0.48984
R26 VP.n9 VP.n6 0.354971
R27 VP.n22 VP.n21 0.354971
R28 VP VP.n22 0.26696
R29 VP.n10 VP.n9 0.189894
R30 VP.n11 VP.n10 0.189894
R31 VP.n11 VP.n3 0.189894
R32 VP.n15 VP.n3 0.189894
R33 VP.n16 VP.n15 0.189894
R34 VP.n17 VP.n16 0.189894
R35 VP.n17 VP.n1 0.189894
R36 VP.n21 VP.n1 0.189894
R37 VTAIL.n122 VTAIL.n112 756.745
R38 VTAIL.n10 VTAIL.n0 756.745
R39 VTAIL.n26 VTAIL.n16 756.745
R40 VTAIL.n42 VTAIL.n32 756.745
R41 VTAIL.n106 VTAIL.n96 756.745
R42 VTAIL.n90 VTAIL.n80 756.745
R43 VTAIL.n74 VTAIL.n64 756.745
R44 VTAIL.n58 VTAIL.n48 756.745
R45 VTAIL.n116 VTAIL.n115 585
R46 VTAIL.n121 VTAIL.n120 585
R47 VTAIL.n123 VTAIL.n122 585
R48 VTAIL.n4 VTAIL.n3 585
R49 VTAIL.n9 VTAIL.n8 585
R50 VTAIL.n11 VTAIL.n10 585
R51 VTAIL.n20 VTAIL.n19 585
R52 VTAIL.n25 VTAIL.n24 585
R53 VTAIL.n27 VTAIL.n26 585
R54 VTAIL.n36 VTAIL.n35 585
R55 VTAIL.n41 VTAIL.n40 585
R56 VTAIL.n43 VTAIL.n42 585
R57 VTAIL.n107 VTAIL.n106 585
R58 VTAIL.n105 VTAIL.n104 585
R59 VTAIL.n100 VTAIL.n99 585
R60 VTAIL.n91 VTAIL.n90 585
R61 VTAIL.n89 VTAIL.n88 585
R62 VTAIL.n84 VTAIL.n83 585
R63 VTAIL.n75 VTAIL.n74 585
R64 VTAIL.n73 VTAIL.n72 585
R65 VTAIL.n68 VTAIL.n67 585
R66 VTAIL.n59 VTAIL.n58 585
R67 VTAIL.n57 VTAIL.n56 585
R68 VTAIL.n52 VTAIL.n51 585
R69 VTAIL.n117 VTAIL.t3 336.901
R70 VTAIL.n5 VTAIL.t2 336.901
R71 VTAIL.n21 VTAIL.t5 336.901
R72 VTAIL.n37 VTAIL.t6 336.901
R73 VTAIL.n101 VTAIL.t7 336.901
R74 VTAIL.n85 VTAIL.t4 336.901
R75 VTAIL.n69 VTAIL.t1 336.901
R76 VTAIL.n53 VTAIL.t0 336.901
R77 VTAIL.n121 VTAIL.n115 171.744
R78 VTAIL.n122 VTAIL.n121 171.744
R79 VTAIL.n9 VTAIL.n3 171.744
R80 VTAIL.n10 VTAIL.n9 171.744
R81 VTAIL.n25 VTAIL.n19 171.744
R82 VTAIL.n26 VTAIL.n25 171.744
R83 VTAIL.n41 VTAIL.n35 171.744
R84 VTAIL.n42 VTAIL.n41 171.744
R85 VTAIL.n106 VTAIL.n105 171.744
R86 VTAIL.n105 VTAIL.n99 171.744
R87 VTAIL.n90 VTAIL.n89 171.744
R88 VTAIL.n89 VTAIL.n83 171.744
R89 VTAIL.n74 VTAIL.n73 171.744
R90 VTAIL.n73 VTAIL.n67 171.744
R91 VTAIL.n58 VTAIL.n57 171.744
R92 VTAIL.n57 VTAIL.n51 171.744
R93 VTAIL.t3 VTAIL.n115 85.8723
R94 VTAIL.t2 VTAIL.n3 85.8723
R95 VTAIL.t5 VTAIL.n19 85.8723
R96 VTAIL.t6 VTAIL.n35 85.8723
R97 VTAIL.t7 VTAIL.n99 85.8723
R98 VTAIL.t4 VTAIL.n83 85.8723
R99 VTAIL.t1 VTAIL.n67 85.8723
R100 VTAIL.t0 VTAIL.n51 85.8723
R101 VTAIL.n127 VTAIL.n126 36.646
R102 VTAIL.n15 VTAIL.n14 36.646
R103 VTAIL.n31 VTAIL.n30 36.646
R104 VTAIL.n47 VTAIL.n46 36.646
R105 VTAIL.n111 VTAIL.n110 36.646
R106 VTAIL.n95 VTAIL.n94 36.646
R107 VTAIL.n79 VTAIL.n78 36.646
R108 VTAIL.n63 VTAIL.n62 36.646
R109 VTAIL.n127 VTAIL.n111 18.7203
R110 VTAIL.n63 VTAIL.n47 18.7203
R111 VTAIL.n117 VTAIL.n116 16.193
R112 VTAIL.n5 VTAIL.n4 16.193
R113 VTAIL.n21 VTAIL.n20 16.193
R114 VTAIL.n37 VTAIL.n36 16.193
R115 VTAIL.n101 VTAIL.n100 16.193
R116 VTAIL.n85 VTAIL.n84 16.193
R117 VTAIL.n69 VTAIL.n68 16.193
R118 VTAIL.n53 VTAIL.n52 16.193
R119 VTAIL.n120 VTAIL.n119 12.8005
R120 VTAIL.n8 VTAIL.n7 12.8005
R121 VTAIL.n24 VTAIL.n23 12.8005
R122 VTAIL.n40 VTAIL.n39 12.8005
R123 VTAIL.n104 VTAIL.n103 12.8005
R124 VTAIL.n88 VTAIL.n87 12.8005
R125 VTAIL.n72 VTAIL.n71 12.8005
R126 VTAIL.n56 VTAIL.n55 12.8005
R127 VTAIL.n123 VTAIL.n114 12.0247
R128 VTAIL.n11 VTAIL.n2 12.0247
R129 VTAIL.n27 VTAIL.n18 12.0247
R130 VTAIL.n43 VTAIL.n34 12.0247
R131 VTAIL.n107 VTAIL.n98 12.0247
R132 VTAIL.n91 VTAIL.n82 12.0247
R133 VTAIL.n75 VTAIL.n66 12.0247
R134 VTAIL.n59 VTAIL.n50 12.0247
R135 VTAIL.n124 VTAIL.n112 11.249
R136 VTAIL.n12 VTAIL.n0 11.249
R137 VTAIL.n28 VTAIL.n16 11.249
R138 VTAIL.n44 VTAIL.n32 11.249
R139 VTAIL.n108 VTAIL.n96 11.249
R140 VTAIL.n92 VTAIL.n80 11.249
R141 VTAIL.n76 VTAIL.n64 11.249
R142 VTAIL.n60 VTAIL.n48 11.249
R143 VTAIL.n126 VTAIL.n125 9.45567
R144 VTAIL.n14 VTAIL.n13 9.45567
R145 VTAIL.n30 VTAIL.n29 9.45567
R146 VTAIL.n46 VTAIL.n45 9.45567
R147 VTAIL.n110 VTAIL.n109 9.45567
R148 VTAIL.n94 VTAIL.n93 9.45567
R149 VTAIL.n78 VTAIL.n77 9.45567
R150 VTAIL.n62 VTAIL.n61 9.45567
R151 VTAIL.n125 VTAIL.n124 9.3005
R152 VTAIL.n114 VTAIL.n113 9.3005
R153 VTAIL.n119 VTAIL.n118 9.3005
R154 VTAIL.n13 VTAIL.n12 9.3005
R155 VTAIL.n2 VTAIL.n1 9.3005
R156 VTAIL.n7 VTAIL.n6 9.3005
R157 VTAIL.n29 VTAIL.n28 9.3005
R158 VTAIL.n18 VTAIL.n17 9.3005
R159 VTAIL.n23 VTAIL.n22 9.3005
R160 VTAIL.n45 VTAIL.n44 9.3005
R161 VTAIL.n34 VTAIL.n33 9.3005
R162 VTAIL.n39 VTAIL.n38 9.3005
R163 VTAIL.n109 VTAIL.n108 9.3005
R164 VTAIL.n98 VTAIL.n97 9.3005
R165 VTAIL.n103 VTAIL.n102 9.3005
R166 VTAIL.n93 VTAIL.n92 9.3005
R167 VTAIL.n82 VTAIL.n81 9.3005
R168 VTAIL.n87 VTAIL.n86 9.3005
R169 VTAIL.n77 VTAIL.n76 9.3005
R170 VTAIL.n66 VTAIL.n65 9.3005
R171 VTAIL.n71 VTAIL.n70 9.3005
R172 VTAIL.n61 VTAIL.n60 9.3005
R173 VTAIL.n50 VTAIL.n49 9.3005
R174 VTAIL.n55 VTAIL.n54 9.3005
R175 VTAIL.n102 VTAIL.n101 3.91276
R176 VTAIL.n86 VTAIL.n85 3.91276
R177 VTAIL.n70 VTAIL.n69 3.91276
R178 VTAIL.n54 VTAIL.n53 3.91276
R179 VTAIL.n118 VTAIL.n117 3.91276
R180 VTAIL.n6 VTAIL.n5 3.91276
R181 VTAIL.n22 VTAIL.n21 3.91276
R182 VTAIL.n38 VTAIL.n37 3.91276
R183 VTAIL.n79 VTAIL.n63 3.46602
R184 VTAIL.n111 VTAIL.n95 3.46602
R185 VTAIL.n47 VTAIL.n31 3.46602
R186 VTAIL.n126 VTAIL.n112 2.71565
R187 VTAIL.n14 VTAIL.n0 2.71565
R188 VTAIL.n30 VTAIL.n16 2.71565
R189 VTAIL.n46 VTAIL.n32 2.71565
R190 VTAIL.n110 VTAIL.n96 2.71565
R191 VTAIL.n94 VTAIL.n80 2.71565
R192 VTAIL.n78 VTAIL.n64 2.71565
R193 VTAIL.n62 VTAIL.n48 2.71565
R194 VTAIL.n124 VTAIL.n123 1.93989
R195 VTAIL.n12 VTAIL.n11 1.93989
R196 VTAIL.n28 VTAIL.n27 1.93989
R197 VTAIL.n44 VTAIL.n43 1.93989
R198 VTAIL.n108 VTAIL.n107 1.93989
R199 VTAIL.n92 VTAIL.n91 1.93989
R200 VTAIL.n76 VTAIL.n75 1.93989
R201 VTAIL.n60 VTAIL.n59 1.93989
R202 VTAIL VTAIL.n15 1.79145
R203 VTAIL VTAIL.n127 1.67507
R204 VTAIL.n120 VTAIL.n114 1.16414
R205 VTAIL.n8 VTAIL.n2 1.16414
R206 VTAIL.n24 VTAIL.n18 1.16414
R207 VTAIL.n40 VTAIL.n34 1.16414
R208 VTAIL.n104 VTAIL.n98 1.16414
R209 VTAIL.n88 VTAIL.n82 1.16414
R210 VTAIL.n72 VTAIL.n66 1.16414
R211 VTAIL.n56 VTAIL.n50 1.16414
R212 VTAIL.n95 VTAIL.n79 0.470328
R213 VTAIL.n31 VTAIL.n15 0.470328
R214 VTAIL.n119 VTAIL.n116 0.388379
R215 VTAIL.n7 VTAIL.n4 0.388379
R216 VTAIL.n23 VTAIL.n20 0.388379
R217 VTAIL.n39 VTAIL.n36 0.388379
R218 VTAIL.n103 VTAIL.n100 0.388379
R219 VTAIL.n87 VTAIL.n84 0.388379
R220 VTAIL.n71 VTAIL.n68 0.388379
R221 VTAIL.n55 VTAIL.n52 0.388379
R222 VTAIL.n118 VTAIL.n113 0.155672
R223 VTAIL.n125 VTAIL.n113 0.155672
R224 VTAIL.n6 VTAIL.n1 0.155672
R225 VTAIL.n13 VTAIL.n1 0.155672
R226 VTAIL.n22 VTAIL.n17 0.155672
R227 VTAIL.n29 VTAIL.n17 0.155672
R228 VTAIL.n38 VTAIL.n33 0.155672
R229 VTAIL.n45 VTAIL.n33 0.155672
R230 VTAIL.n109 VTAIL.n97 0.155672
R231 VTAIL.n102 VTAIL.n97 0.155672
R232 VTAIL.n93 VTAIL.n81 0.155672
R233 VTAIL.n86 VTAIL.n81 0.155672
R234 VTAIL.n77 VTAIL.n65 0.155672
R235 VTAIL.n70 VTAIL.n65 0.155672
R236 VTAIL.n61 VTAIL.n49 0.155672
R237 VTAIL.n54 VTAIL.n49 0.155672
R238 VDD1 VDD1.n1 169.835
R239 VDD1 VDD1.n0 132.369
R240 VDD1.n0 VDD1.t0 9.70349
R241 VDD1.n0 VDD1.t3 9.70349
R242 VDD1.n1 VDD1.t1 9.70349
R243 VDD1.n1 VDD1.t2 9.70349
R244 VN.n0 VN.t1 55.0842
R245 VN.n1 VN.t2 55.0842
R246 VN.n0 VN.t0 53.7611
R247 VN.n1 VN.t3 53.7611
R248 VN VN.n1 45.1823
R249 VN VN.n0 1.94371
R250 VDD2.n2 VDD2.n0 169.31
R251 VDD2.n2 VDD2.n1 132.311
R252 VDD2.n1 VDD2.t0 9.70349
R253 VDD2.n1 VDD2.t1 9.70349
R254 VDD2.n0 VDD2.t2 9.70349
R255 VDD2.n0 VDD2.t3 9.70349
R256 VDD2 VDD2.n2 0.0586897
R257 B.n267 B.n266 585
R258 B.n265 B.n94 585
R259 B.n264 B.n263 585
R260 B.n262 B.n95 585
R261 B.n261 B.n260 585
R262 B.n259 B.n96 585
R263 B.n258 B.n257 585
R264 B.n256 B.n97 585
R265 B.n255 B.n254 585
R266 B.n253 B.n98 585
R267 B.n252 B.n251 585
R268 B.n250 B.n99 585
R269 B.n249 B.n248 585
R270 B.n247 B.n100 585
R271 B.n246 B.n245 585
R272 B.n244 B.n101 585
R273 B.n243 B.n242 585
R274 B.n238 B.n102 585
R275 B.n237 B.n236 585
R276 B.n235 B.n103 585
R277 B.n234 B.n233 585
R278 B.n232 B.n104 585
R279 B.n231 B.n230 585
R280 B.n229 B.n105 585
R281 B.n228 B.n227 585
R282 B.n226 B.n106 585
R283 B.n224 B.n223 585
R284 B.n222 B.n109 585
R285 B.n221 B.n220 585
R286 B.n219 B.n110 585
R287 B.n218 B.n217 585
R288 B.n216 B.n111 585
R289 B.n215 B.n214 585
R290 B.n213 B.n112 585
R291 B.n212 B.n211 585
R292 B.n210 B.n113 585
R293 B.n209 B.n208 585
R294 B.n207 B.n114 585
R295 B.n206 B.n205 585
R296 B.n204 B.n115 585
R297 B.n203 B.n202 585
R298 B.n201 B.n116 585
R299 B.n268 B.n93 585
R300 B.n270 B.n269 585
R301 B.n271 B.n92 585
R302 B.n273 B.n272 585
R303 B.n274 B.n91 585
R304 B.n276 B.n275 585
R305 B.n277 B.n90 585
R306 B.n279 B.n278 585
R307 B.n280 B.n89 585
R308 B.n282 B.n281 585
R309 B.n283 B.n88 585
R310 B.n285 B.n284 585
R311 B.n286 B.n87 585
R312 B.n288 B.n287 585
R313 B.n289 B.n86 585
R314 B.n291 B.n290 585
R315 B.n292 B.n85 585
R316 B.n294 B.n293 585
R317 B.n295 B.n84 585
R318 B.n297 B.n296 585
R319 B.n298 B.n83 585
R320 B.n300 B.n299 585
R321 B.n301 B.n82 585
R322 B.n303 B.n302 585
R323 B.n304 B.n81 585
R324 B.n306 B.n305 585
R325 B.n307 B.n80 585
R326 B.n309 B.n308 585
R327 B.n310 B.n79 585
R328 B.n312 B.n311 585
R329 B.n313 B.n78 585
R330 B.n315 B.n314 585
R331 B.n316 B.n77 585
R332 B.n318 B.n317 585
R333 B.n319 B.n76 585
R334 B.n321 B.n320 585
R335 B.n322 B.n75 585
R336 B.n324 B.n323 585
R337 B.n325 B.n74 585
R338 B.n327 B.n326 585
R339 B.n328 B.n73 585
R340 B.n330 B.n329 585
R341 B.n331 B.n72 585
R342 B.n333 B.n332 585
R343 B.n334 B.n71 585
R344 B.n336 B.n335 585
R345 B.n337 B.n70 585
R346 B.n339 B.n338 585
R347 B.n340 B.n69 585
R348 B.n342 B.n341 585
R349 B.n343 B.n68 585
R350 B.n345 B.n344 585
R351 B.n346 B.n67 585
R352 B.n348 B.n347 585
R353 B.n349 B.n66 585
R354 B.n351 B.n350 585
R355 B.n352 B.n65 585
R356 B.n354 B.n353 585
R357 B.n355 B.n64 585
R358 B.n357 B.n356 585
R359 B.n358 B.n63 585
R360 B.n360 B.n359 585
R361 B.n361 B.n62 585
R362 B.n363 B.n362 585
R363 B.n364 B.n61 585
R364 B.n366 B.n365 585
R365 B.n367 B.n60 585
R366 B.n369 B.n368 585
R367 B.n370 B.n59 585
R368 B.n372 B.n371 585
R369 B.n373 B.n58 585
R370 B.n375 B.n374 585
R371 B.n376 B.n57 585
R372 B.n378 B.n377 585
R373 B.n379 B.n56 585
R374 B.n381 B.n380 585
R375 B.n382 B.n55 585
R376 B.n384 B.n383 585
R377 B.n385 B.n54 585
R378 B.n387 B.n386 585
R379 B.n388 B.n53 585
R380 B.n390 B.n389 585
R381 B.n391 B.n52 585
R382 B.n393 B.n392 585
R383 B.n394 B.n51 585
R384 B.n396 B.n395 585
R385 B.n397 B.n50 585
R386 B.n399 B.n398 585
R387 B.n463 B.n462 585
R388 B.n461 B.n24 585
R389 B.n460 B.n459 585
R390 B.n458 B.n25 585
R391 B.n457 B.n456 585
R392 B.n455 B.n26 585
R393 B.n454 B.n453 585
R394 B.n452 B.n27 585
R395 B.n451 B.n450 585
R396 B.n449 B.n28 585
R397 B.n448 B.n447 585
R398 B.n446 B.n29 585
R399 B.n445 B.n444 585
R400 B.n443 B.n30 585
R401 B.n442 B.n441 585
R402 B.n440 B.n31 585
R403 B.n438 B.n437 585
R404 B.n436 B.n34 585
R405 B.n435 B.n434 585
R406 B.n433 B.n35 585
R407 B.n432 B.n431 585
R408 B.n430 B.n36 585
R409 B.n429 B.n428 585
R410 B.n427 B.n37 585
R411 B.n426 B.n425 585
R412 B.n424 B.n38 585
R413 B.n423 B.n422 585
R414 B.n421 B.n39 585
R415 B.n420 B.n419 585
R416 B.n418 B.n43 585
R417 B.n417 B.n416 585
R418 B.n415 B.n44 585
R419 B.n414 B.n413 585
R420 B.n412 B.n45 585
R421 B.n411 B.n410 585
R422 B.n409 B.n46 585
R423 B.n408 B.n407 585
R424 B.n406 B.n47 585
R425 B.n405 B.n404 585
R426 B.n403 B.n48 585
R427 B.n402 B.n401 585
R428 B.n400 B.n49 585
R429 B.n464 B.n23 585
R430 B.n466 B.n465 585
R431 B.n467 B.n22 585
R432 B.n469 B.n468 585
R433 B.n470 B.n21 585
R434 B.n472 B.n471 585
R435 B.n473 B.n20 585
R436 B.n475 B.n474 585
R437 B.n476 B.n19 585
R438 B.n478 B.n477 585
R439 B.n479 B.n18 585
R440 B.n481 B.n480 585
R441 B.n482 B.n17 585
R442 B.n484 B.n483 585
R443 B.n485 B.n16 585
R444 B.n487 B.n486 585
R445 B.n488 B.n15 585
R446 B.n490 B.n489 585
R447 B.n491 B.n14 585
R448 B.n493 B.n492 585
R449 B.n494 B.n13 585
R450 B.n496 B.n495 585
R451 B.n497 B.n12 585
R452 B.n499 B.n498 585
R453 B.n500 B.n11 585
R454 B.n502 B.n501 585
R455 B.n503 B.n10 585
R456 B.n505 B.n504 585
R457 B.n506 B.n9 585
R458 B.n508 B.n507 585
R459 B.n509 B.n8 585
R460 B.n511 B.n510 585
R461 B.n512 B.n7 585
R462 B.n514 B.n513 585
R463 B.n515 B.n6 585
R464 B.n517 B.n516 585
R465 B.n518 B.n5 585
R466 B.n520 B.n519 585
R467 B.n521 B.n4 585
R468 B.n523 B.n522 585
R469 B.n524 B.n3 585
R470 B.n526 B.n525 585
R471 B.n527 B.n0 585
R472 B.n2 B.n1 585
R473 B.n138 B.n137 585
R474 B.n140 B.n139 585
R475 B.n141 B.n136 585
R476 B.n143 B.n142 585
R477 B.n144 B.n135 585
R478 B.n146 B.n145 585
R479 B.n147 B.n134 585
R480 B.n149 B.n148 585
R481 B.n150 B.n133 585
R482 B.n152 B.n151 585
R483 B.n153 B.n132 585
R484 B.n155 B.n154 585
R485 B.n156 B.n131 585
R486 B.n158 B.n157 585
R487 B.n159 B.n130 585
R488 B.n161 B.n160 585
R489 B.n162 B.n129 585
R490 B.n164 B.n163 585
R491 B.n165 B.n128 585
R492 B.n167 B.n166 585
R493 B.n168 B.n127 585
R494 B.n170 B.n169 585
R495 B.n171 B.n126 585
R496 B.n173 B.n172 585
R497 B.n174 B.n125 585
R498 B.n176 B.n175 585
R499 B.n177 B.n124 585
R500 B.n179 B.n178 585
R501 B.n180 B.n123 585
R502 B.n182 B.n181 585
R503 B.n183 B.n122 585
R504 B.n185 B.n184 585
R505 B.n186 B.n121 585
R506 B.n188 B.n187 585
R507 B.n189 B.n120 585
R508 B.n191 B.n190 585
R509 B.n192 B.n119 585
R510 B.n194 B.n193 585
R511 B.n195 B.n118 585
R512 B.n197 B.n196 585
R513 B.n198 B.n117 585
R514 B.n200 B.n199 585
R515 B.n199 B.n116 506.916
R516 B.n268 B.n267 506.916
R517 B.n400 B.n399 506.916
R518 B.n462 B.n23 506.916
R519 B.n239 B.t10 306.433
R520 B.n40 B.t8 306.433
R521 B.n107 B.t1 306.433
R522 B.n32 B.t5 306.433
R523 B.n529 B.n528 256.663
R524 B.n528 B.n527 235.042
R525 B.n528 B.n2 235.042
R526 B.n107 B.t0 231.136
R527 B.n239 B.t9 231.136
R528 B.n40 B.t6 231.136
R529 B.n32 B.t3 231.136
R530 B.n240 B.t11 228.47
R531 B.n41 B.t7 228.47
R532 B.n108 B.t2 228.47
R533 B.n33 B.t4 228.47
R534 B.n203 B.n116 163.367
R535 B.n204 B.n203 163.367
R536 B.n205 B.n204 163.367
R537 B.n205 B.n114 163.367
R538 B.n209 B.n114 163.367
R539 B.n210 B.n209 163.367
R540 B.n211 B.n210 163.367
R541 B.n211 B.n112 163.367
R542 B.n215 B.n112 163.367
R543 B.n216 B.n215 163.367
R544 B.n217 B.n216 163.367
R545 B.n217 B.n110 163.367
R546 B.n221 B.n110 163.367
R547 B.n222 B.n221 163.367
R548 B.n223 B.n222 163.367
R549 B.n223 B.n106 163.367
R550 B.n228 B.n106 163.367
R551 B.n229 B.n228 163.367
R552 B.n230 B.n229 163.367
R553 B.n230 B.n104 163.367
R554 B.n234 B.n104 163.367
R555 B.n235 B.n234 163.367
R556 B.n236 B.n235 163.367
R557 B.n236 B.n102 163.367
R558 B.n243 B.n102 163.367
R559 B.n244 B.n243 163.367
R560 B.n245 B.n244 163.367
R561 B.n245 B.n100 163.367
R562 B.n249 B.n100 163.367
R563 B.n250 B.n249 163.367
R564 B.n251 B.n250 163.367
R565 B.n251 B.n98 163.367
R566 B.n255 B.n98 163.367
R567 B.n256 B.n255 163.367
R568 B.n257 B.n256 163.367
R569 B.n257 B.n96 163.367
R570 B.n261 B.n96 163.367
R571 B.n262 B.n261 163.367
R572 B.n263 B.n262 163.367
R573 B.n263 B.n94 163.367
R574 B.n267 B.n94 163.367
R575 B.n399 B.n50 163.367
R576 B.n395 B.n50 163.367
R577 B.n395 B.n394 163.367
R578 B.n394 B.n393 163.367
R579 B.n393 B.n52 163.367
R580 B.n389 B.n52 163.367
R581 B.n389 B.n388 163.367
R582 B.n388 B.n387 163.367
R583 B.n387 B.n54 163.367
R584 B.n383 B.n54 163.367
R585 B.n383 B.n382 163.367
R586 B.n382 B.n381 163.367
R587 B.n381 B.n56 163.367
R588 B.n377 B.n56 163.367
R589 B.n377 B.n376 163.367
R590 B.n376 B.n375 163.367
R591 B.n375 B.n58 163.367
R592 B.n371 B.n58 163.367
R593 B.n371 B.n370 163.367
R594 B.n370 B.n369 163.367
R595 B.n369 B.n60 163.367
R596 B.n365 B.n60 163.367
R597 B.n365 B.n364 163.367
R598 B.n364 B.n363 163.367
R599 B.n363 B.n62 163.367
R600 B.n359 B.n62 163.367
R601 B.n359 B.n358 163.367
R602 B.n358 B.n357 163.367
R603 B.n357 B.n64 163.367
R604 B.n353 B.n64 163.367
R605 B.n353 B.n352 163.367
R606 B.n352 B.n351 163.367
R607 B.n351 B.n66 163.367
R608 B.n347 B.n66 163.367
R609 B.n347 B.n346 163.367
R610 B.n346 B.n345 163.367
R611 B.n345 B.n68 163.367
R612 B.n341 B.n68 163.367
R613 B.n341 B.n340 163.367
R614 B.n340 B.n339 163.367
R615 B.n339 B.n70 163.367
R616 B.n335 B.n70 163.367
R617 B.n335 B.n334 163.367
R618 B.n334 B.n333 163.367
R619 B.n333 B.n72 163.367
R620 B.n329 B.n72 163.367
R621 B.n329 B.n328 163.367
R622 B.n328 B.n327 163.367
R623 B.n327 B.n74 163.367
R624 B.n323 B.n74 163.367
R625 B.n323 B.n322 163.367
R626 B.n322 B.n321 163.367
R627 B.n321 B.n76 163.367
R628 B.n317 B.n76 163.367
R629 B.n317 B.n316 163.367
R630 B.n316 B.n315 163.367
R631 B.n315 B.n78 163.367
R632 B.n311 B.n78 163.367
R633 B.n311 B.n310 163.367
R634 B.n310 B.n309 163.367
R635 B.n309 B.n80 163.367
R636 B.n305 B.n80 163.367
R637 B.n305 B.n304 163.367
R638 B.n304 B.n303 163.367
R639 B.n303 B.n82 163.367
R640 B.n299 B.n82 163.367
R641 B.n299 B.n298 163.367
R642 B.n298 B.n297 163.367
R643 B.n297 B.n84 163.367
R644 B.n293 B.n84 163.367
R645 B.n293 B.n292 163.367
R646 B.n292 B.n291 163.367
R647 B.n291 B.n86 163.367
R648 B.n287 B.n86 163.367
R649 B.n287 B.n286 163.367
R650 B.n286 B.n285 163.367
R651 B.n285 B.n88 163.367
R652 B.n281 B.n88 163.367
R653 B.n281 B.n280 163.367
R654 B.n280 B.n279 163.367
R655 B.n279 B.n90 163.367
R656 B.n275 B.n90 163.367
R657 B.n275 B.n274 163.367
R658 B.n274 B.n273 163.367
R659 B.n273 B.n92 163.367
R660 B.n269 B.n92 163.367
R661 B.n269 B.n268 163.367
R662 B.n462 B.n461 163.367
R663 B.n461 B.n460 163.367
R664 B.n460 B.n25 163.367
R665 B.n456 B.n25 163.367
R666 B.n456 B.n455 163.367
R667 B.n455 B.n454 163.367
R668 B.n454 B.n27 163.367
R669 B.n450 B.n27 163.367
R670 B.n450 B.n449 163.367
R671 B.n449 B.n448 163.367
R672 B.n448 B.n29 163.367
R673 B.n444 B.n29 163.367
R674 B.n444 B.n443 163.367
R675 B.n443 B.n442 163.367
R676 B.n442 B.n31 163.367
R677 B.n437 B.n31 163.367
R678 B.n437 B.n436 163.367
R679 B.n436 B.n435 163.367
R680 B.n435 B.n35 163.367
R681 B.n431 B.n35 163.367
R682 B.n431 B.n430 163.367
R683 B.n430 B.n429 163.367
R684 B.n429 B.n37 163.367
R685 B.n425 B.n37 163.367
R686 B.n425 B.n424 163.367
R687 B.n424 B.n423 163.367
R688 B.n423 B.n39 163.367
R689 B.n419 B.n39 163.367
R690 B.n419 B.n418 163.367
R691 B.n418 B.n417 163.367
R692 B.n417 B.n44 163.367
R693 B.n413 B.n44 163.367
R694 B.n413 B.n412 163.367
R695 B.n412 B.n411 163.367
R696 B.n411 B.n46 163.367
R697 B.n407 B.n46 163.367
R698 B.n407 B.n406 163.367
R699 B.n406 B.n405 163.367
R700 B.n405 B.n48 163.367
R701 B.n401 B.n48 163.367
R702 B.n401 B.n400 163.367
R703 B.n466 B.n23 163.367
R704 B.n467 B.n466 163.367
R705 B.n468 B.n467 163.367
R706 B.n468 B.n21 163.367
R707 B.n472 B.n21 163.367
R708 B.n473 B.n472 163.367
R709 B.n474 B.n473 163.367
R710 B.n474 B.n19 163.367
R711 B.n478 B.n19 163.367
R712 B.n479 B.n478 163.367
R713 B.n480 B.n479 163.367
R714 B.n480 B.n17 163.367
R715 B.n484 B.n17 163.367
R716 B.n485 B.n484 163.367
R717 B.n486 B.n485 163.367
R718 B.n486 B.n15 163.367
R719 B.n490 B.n15 163.367
R720 B.n491 B.n490 163.367
R721 B.n492 B.n491 163.367
R722 B.n492 B.n13 163.367
R723 B.n496 B.n13 163.367
R724 B.n497 B.n496 163.367
R725 B.n498 B.n497 163.367
R726 B.n498 B.n11 163.367
R727 B.n502 B.n11 163.367
R728 B.n503 B.n502 163.367
R729 B.n504 B.n503 163.367
R730 B.n504 B.n9 163.367
R731 B.n508 B.n9 163.367
R732 B.n509 B.n508 163.367
R733 B.n510 B.n509 163.367
R734 B.n510 B.n7 163.367
R735 B.n514 B.n7 163.367
R736 B.n515 B.n514 163.367
R737 B.n516 B.n515 163.367
R738 B.n516 B.n5 163.367
R739 B.n520 B.n5 163.367
R740 B.n521 B.n520 163.367
R741 B.n522 B.n521 163.367
R742 B.n522 B.n3 163.367
R743 B.n526 B.n3 163.367
R744 B.n527 B.n526 163.367
R745 B.n138 B.n2 163.367
R746 B.n139 B.n138 163.367
R747 B.n139 B.n136 163.367
R748 B.n143 B.n136 163.367
R749 B.n144 B.n143 163.367
R750 B.n145 B.n144 163.367
R751 B.n145 B.n134 163.367
R752 B.n149 B.n134 163.367
R753 B.n150 B.n149 163.367
R754 B.n151 B.n150 163.367
R755 B.n151 B.n132 163.367
R756 B.n155 B.n132 163.367
R757 B.n156 B.n155 163.367
R758 B.n157 B.n156 163.367
R759 B.n157 B.n130 163.367
R760 B.n161 B.n130 163.367
R761 B.n162 B.n161 163.367
R762 B.n163 B.n162 163.367
R763 B.n163 B.n128 163.367
R764 B.n167 B.n128 163.367
R765 B.n168 B.n167 163.367
R766 B.n169 B.n168 163.367
R767 B.n169 B.n126 163.367
R768 B.n173 B.n126 163.367
R769 B.n174 B.n173 163.367
R770 B.n175 B.n174 163.367
R771 B.n175 B.n124 163.367
R772 B.n179 B.n124 163.367
R773 B.n180 B.n179 163.367
R774 B.n181 B.n180 163.367
R775 B.n181 B.n122 163.367
R776 B.n185 B.n122 163.367
R777 B.n186 B.n185 163.367
R778 B.n187 B.n186 163.367
R779 B.n187 B.n120 163.367
R780 B.n191 B.n120 163.367
R781 B.n192 B.n191 163.367
R782 B.n193 B.n192 163.367
R783 B.n193 B.n118 163.367
R784 B.n197 B.n118 163.367
R785 B.n198 B.n197 163.367
R786 B.n199 B.n198 163.367
R787 B.n108 B.n107 77.9641
R788 B.n240 B.n239 77.9641
R789 B.n41 B.n40 77.9641
R790 B.n33 B.n32 77.9641
R791 B.n225 B.n108 59.5399
R792 B.n241 B.n240 59.5399
R793 B.n42 B.n41 59.5399
R794 B.n439 B.n33 59.5399
R795 B.n464 B.n463 32.9371
R796 B.n398 B.n49 32.9371
R797 B.n266 B.n93 32.9371
R798 B.n201 B.n200 32.9371
R799 B B.n529 18.0485
R800 B.n465 B.n464 10.6151
R801 B.n465 B.n22 10.6151
R802 B.n469 B.n22 10.6151
R803 B.n470 B.n469 10.6151
R804 B.n471 B.n470 10.6151
R805 B.n471 B.n20 10.6151
R806 B.n475 B.n20 10.6151
R807 B.n476 B.n475 10.6151
R808 B.n477 B.n476 10.6151
R809 B.n477 B.n18 10.6151
R810 B.n481 B.n18 10.6151
R811 B.n482 B.n481 10.6151
R812 B.n483 B.n482 10.6151
R813 B.n483 B.n16 10.6151
R814 B.n487 B.n16 10.6151
R815 B.n488 B.n487 10.6151
R816 B.n489 B.n488 10.6151
R817 B.n489 B.n14 10.6151
R818 B.n493 B.n14 10.6151
R819 B.n494 B.n493 10.6151
R820 B.n495 B.n494 10.6151
R821 B.n495 B.n12 10.6151
R822 B.n499 B.n12 10.6151
R823 B.n500 B.n499 10.6151
R824 B.n501 B.n500 10.6151
R825 B.n501 B.n10 10.6151
R826 B.n505 B.n10 10.6151
R827 B.n506 B.n505 10.6151
R828 B.n507 B.n506 10.6151
R829 B.n507 B.n8 10.6151
R830 B.n511 B.n8 10.6151
R831 B.n512 B.n511 10.6151
R832 B.n513 B.n512 10.6151
R833 B.n513 B.n6 10.6151
R834 B.n517 B.n6 10.6151
R835 B.n518 B.n517 10.6151
R836 B.n519 B.n518 10.6151
R837 B.n519 B.n4 10.6151
R838 B.n523 B.n4 10.6151
R839 B.n524 B.n523 10.6151
R840 B.n525 B.n524 10.6151
R841 B.n525 B.n0 10.6151
R842 B.n463 B.n24 10.6151
R843 B.n459 B.n24 10.6151
R844 B.n459 B.n458 10.6151
R845 B.n458 B.n457 10.6151
R846 B.n457 B.n26 10.6151
R847 B.n453 B.n26 10.6151
R848 B.n453 B.n452 10.6151
R849 B.n452 B.n451 10.6151
R850 B.n451 B.n28 10.6151
R851 B.n447 B.n28 10.6151
R852 B.n447 B.n446 10.6151
R853 B.n446 B.n445 10.6151
R854 B.n445 B.n30 10.6151
R855 B.n441 B.n30 10.6151
R856 B.n441 B.n440 10.6151
R857 B.n438 B.n34 10.6151
R858 B.n434 B.n34 10.6151
R859 B.n434 B.n433 10.6151
R860 B.n433 B.n432 10.6151
R861 B.n432 B.n36 10.6151
R862 B.n428 B.n36 10.6151
R863 B.n428 B.n427 10.6151
R864 B.n427 B.n426 10.6151
R865 B.n426 B.n38 10.6151
R866 B.n422 B.n421 10.6151
R867 B.n421 B.n420 10.6151
R868 B.n420 B.n43 10.6151
R869 B.n416 B.n43 10.6151
R870 B.n416 B.n415 10.6151
R871 B.n415 B.n414 10.6151
R872 B.n414 B.n45 10.6151
R873 B.n410 B.n45 10.6151
R874 B.n410 B.n409 10.6151
R875 B.n409 B.n408 10.6151
R876 B.n408 B.n47 10.6151
R877 B.n404 B.n47 10.6151
R878 B.n404 B.n403 10.6151
R879 B.n403 B.n402 10.6151
R880 B.n402 B.n49 10.6151
R881 B.n398 B.n397 10.6151
R882 B.n397 B.n396 10.6151
R883 B.n396 B.n51 10.6151
R884 B.n392 B.n51 10.6151
R885 B.n392 B.n391 10.6151
R886 B.n391 B.n390 10.6151
R887 B.n390 B.n53 10.6151
R888 B.n386 B.n53 10.6151
R889 B.n386 B.n385 10.6151
R890 B.n385 B.n384 10.6151
R891 B.n384 B.n55 10.6151
R892 B.n380 B.n55 10.6151
R893 B.n380 B.n379 10.6151
R894 B.n379 B.n378 10.6151
R895 B.n378 B.n57 10.6151
R896 B.n374 B.n57 10.6151
R897 B.n374 B.n373 10.6151
R898 B.n373 B.n372 10.6151
R899 B.n372 B.n59 10.6151
R900 B.n368 B.n59 10.6151
R901 B.n368 B.n367 10.6151
R902 B.n367 B.n366 10.6151
R903 B.n366 B.n61 10.6151
R904 B.n362 B.n61 10.6151
R905 B.n362 B.n361 10.6151
R906 B.n361 B.n360 10.6151
R907 B.n360 B.n63 10.6151
R908 B.n356 B.n63 10.6151
R909 B.n356 B.n355 10.6151
R910 B.n355 B.n354 10.6151
R911 B.n354 B.n65 10.6151
R912 B.n350 B.n65 10.6151
R913 B.n350 B.n349 10.6151
R914 B.n349 B.n348 10.6151
R915 B.n348 B.n67 10.6151
R916 B.n344 B.n67 10.6151
R917 B.n344 B.n343 10.6151
R918 B.n343 B.n342 10.6151
R919 B.n342 B.n69 10.6151
R920 B.n338 B.n69 10.6151
R921 B.n338 B.n337 10.6151
R922 B.n337 B.n336 10.6151
R923 B.n336 B.n71 10.6151
R924 B.n332 B.n71 10.6151
R925 B.n332 B.n331 10.6151
R926 B.n331 B.n330 10.6151
R927 B.n330 B.n73 10.6151
R928 B.n326 B.n73 10.6151
R929 B.n326 B.n325 10.6151
R930 B.n325 B.n324 10.6151
R931 B.n324 B.n75 10.6151
R932 B.n320 B.n75 10.6151
R933 B.n320 B.n319 10.6151
R934 B.n319 B.n318 10.6151
R935 B.n318 B.n77 10.6151
R936 B.n314 B.n77 10.6151
R937 B.n314 B.n313 10.6151
R938 B.n313 B.n312 10.6151
R939 B.n312 B.n79 10.6151
R940 B.n308 B.n79 10.6151
R941 B.n308 B.n307 10.6151
R942 B.n307 B.n306 10.6151
R943 B.n306 B.n81 10.6151
R944 B.n302 B.n81 10.6151
R945 B.n302 B.n301 10.6151
R946 B.n301 B.n300 10.6151
R947 B.n300 B.n83 10.6151
R948 B.n296 B.n83 10.6151
R949 B.n296 B.n295 10.6151
R950 B.n295 B.n294 10.6151
R951 B.n294 B.n85 10.6151
R952 B.n290 B.n85 10.6151
R953 B.n290 B.n289 10.6151
R954 B.n289 B.n288 10.6151
R955 B.n288 B.n87 10.6151
R956 B.n284 B.n87 10.6151
R957 B.n284 B.n283 10.6151
R958 B.n283 B.n282 10.6151
R959 B.n282 B.n89 10.6151
R960 B.n278 B.n89 10.6151
R961 B.n278 B.n277 10.6151
R962 B.n277 B.n276 10.6151
R963 B.n276 B.n91 10.6151
R964 B.n272 B.n91 10.6151
R965 B.n272 B.n271 10.6151
R966 B.n271 B.n270 10.6151
R967 B.n270 B.n93 10.6151
R968 B.n137 B.n1 10.6151
R969 B.n140 B.n137 10.6151
R970 B.n141 B.n140 10.6151
R971 B.n142 B.n141 10.6151
R972 B.n142 B.n135 10.6151
R973 B.n146 B.n135 10.6151
R974 B.n147 B.n146 10.6151
R975 B.n148 B.n147 10.6151
R976 B.n148 B.n133 10.6151
R977 B.n152 B.n133 10.6151
R978 B.n153 B.n152 10.6151
R979 B.n154 B.n153 10.6151
R980 B.n154 B.n131 10.6151
R981 B.n158 B.n131 10.6151
R982 B.n159 B.n158 10.6151
R983 B.n160 B.n159 10.6151
R984 B.n160 B.n129 10.6151
R985 B.n164 B.n129 10.6151
R986 B.n165 B.n164 10.6151
R987 B.n166 B.n165 10.6151
R988 B.n166 B.n127 10.6151
R989 B.n170 B.n127 10.6151
R990 B.n171 B.n170 10.6151
R991 B.n172 B.n171 10.6151
R992 B.n172 B.n125 10.6151
R993 B.n176 B.n125 10.6151
R994 B.n177 B.n176 10.6151
R995 B.n178 B.n177 10.6151
R996 B.n178 B.n123 10.6151
R997 B.n182 B.n123 10.6151
R998 B.n183 B.n182 10.6151
R999 B.n184 B.n183 10.6151
R1000 B.n184 B.n121 10.6151
R1001 B.n188 B.n121 10.6151
R1002 B.n189 B.n188 10.6151
R1003 B.n190 B.n189 10.6151
R1004 B.n190 B.n119 10.6151
R1005 B.n194 B.n119 10.6151
R1006 B.n195 B.n194 10.6151
R1007 B.n196 B.n195 10.6151
R1008 B.n196 B.n117 10.6151
R1009 B.n200 B.n117 10.6151
R1010 B.n202 B.n201 10.6151
R1011 B.n202 B.n115 10.6151
R1012 B.n206 B.n115 10.6151
R1013 B.n207 B.n206 10.6151
R1014 B.n208 B.n207 10.6151
R1015 B.n208 B.n113 10.6151
R1016 B.n212 B.n113 10.6151
R1017 B.n213 B.n212 10.6151
R1018 B.n214 B.n213 10.6151
R1019 B.n214 B.n111 10.6151
R1020 B.n218 B.n111 10.6151
R1021 B.n219 B.n218 10.6151
R1022 B.n220 B.n219 10.6151
R1023 B.n220 B.n109 10.6151
R1024 B.n224 B.n109 10.6151
R1025 B.n227 B.n226 10.6151
R1026 B.n227 B.n105 10.6151
R1027 B.n231 B.n105 10.6151
R1028 B.n232 B.n231 10.6151
R1029 B.n233 B.n232 10.6151
R1030 B.n233 B.n103 10.6151
R1031 B.n237 B.n103 10.6151
R1032 B.n238 B.n237 10.6151
R1033 B.n242 B.n238 10.6151
R1034 B.n246 B.n101 10.6151
R1035 B.n247 B.n246 10.6151
R1036 B.n248 B.n247 10.6151
R1037 B.n248 B.n99 10.6151
R1038 B.n252 B.n99 10.6151
R1039 B.n253 B.n252 10.6151
R1040 B.n254 B.n253 10.6151
R1041 B.n254 B.n97 10.6151
R1042 B.n258 B.n97 10.6151
R1043 B.n259 B.n258 10.6151
R1044 B.n260 B.n259 10.6151
R1045 B.n260 B.n95 10.6151
R1046 B.n264 B.n95 10.6151
R1047 B.n265 B.n264 10.6151
R1048 B.n266 B.n265 10.6151
R1049 B.n440 B.n439 9.36635
R1050 B.n422 B.n42 9.36635
R1051 B.n225 B.n224 9.36635
R1052 B.n241 B.n101 9.36635
R1053 B.n529 B.n0 8.11757
R1054 B.n529 B.n1 8.11757
R1055 B.n439 B.n438 1.24928
R1056 B.n42 B.n38 1.24928
R1057 B.n226 B.n225 1.24928
R1058 B.n242 B.n241 1.24928
C0 VTAIL VDD2 3.95162f
C1 w_n3382_n1638# B 8.195951f
C2 VP VDD2 0.468803f
C3 VDD1 VN 0.154499f
C4 VTAIL B 2.33216f
C5 VTAIL w_n3382_n1638# 2.10215f
C6 VP B 1.94233f
C7 VDD1 VDD2 1.28899f
C8 w_n3382_n1638# VP 6.21579f
C9 VN VDD2 1.64607f
C10 VTAIL VP 2.34532f
C11 VDD1 B 1.22152f
C12 w_n3382_n1638# VDD1 1.41994f
C13 B VN 1.21154f
C14 w_n3382_n1638# VN 5.78004f
C15 VTAIL VDD1 3.89011f
C16 VTAIL VN 2.33122f
C17 B VDD2 1.29197f
C18 w_n3382_n1638# VDD2 1.49965f
C19 VDD1 VP 1.95863f
C20 VP VN 5.38482f
C21 VDD2 VSUBS 0.837658f
C22 VDD1 VSUBS 3.96035f
C23 VTAIL VSUBS 0.717599f
C24 VN VSUBS 5.95325f
C25 VP VSUBS 2.32122f
C26 B VSUBS 4.229924f
C27 w_n3382_n1638# VSUBS 70.00739f
C28 B.n0 VSUBS 0.008433f
C29 B.n1 VSUBS 0.008433f
C30 B.n2 VSUBS 0.012472f
C31 B.n3 VSUBS 0.009558f
C32 B.n4 VSUBS 0.009558f
C33 B.n5 VSUBS 0.009558f
C34 B.n6 VSUBS 0.009558f
C35 B.n7 VSUBS 0.009558f
C36 B.n8 VSUBS 0.009558f
C37 B.n9 VSUBS 0.009558f
C38 B.n10 VSUBS 0.009558f
C39 B.n11 VSUBS 0.009558f
C40 B.n12 VSUBS 0.009558f
C41 B.n13 VSUBS 0.009558f
C42 B.n14 VSUBS 0.009558f
C43 B.n15 VSUBS 0.009558f
C44 B.n16 VSUBS 0.009558f
C45 B.n17 VSUBS 0.009558f
C46 B.n18 VSUBS 0.009558f
C47 B.n19 VSUBS 0.009558f
C48 B.n20 VSUBS 0.009558f
C49 B.n21 VSUBS 0.009558f
C50 B.n22 VSUBS 0.009558f
C51 B.n23 VSUBS 0.021847f
C52 B.n24 VSUBS 0.009558f
C53 B.n25 VSUBS 0.009558f
C54 B.n26 VSUBS 0.009558f
C55 B.n27 VSUBS 0.009558f
C56 B.n28 VSUBS 0.009558f
C57 B.n29 VSUBS 0.009558f
C58 B.n30 VSUBS 0.009558f
C59 B.n31 VSUBS 0.009558f
C60 B.t4 VSUBS 0.067822f
C61 B.t5 VSUBS 0.100816f
C62 B.t3 VSUBS 0.82529f
C63 B.n32 VSUBS 0.171884f
C64 B.n33 VSUBS 0.143313f
C65 B.n34 VSUBS 0.009558f
C66 B.n35 VSUBS 0.009558f
C67 B.n36 VSUBS 0.009558f
C68 B.n37 VSUBS 0.009558f
C69 B.n38 VSUBS 0.005341f
C70 B.n39 VSUBS 0.009558f
C71 B.t7 VSUBS 0.067823f
C72 B.t8 VSUBS 0.100817f
C73 B.t6 VSUBS 0.82529f
C74 B.n40 VSUBS 0.171883f
C75 B.n41 VSUBS 0.143312f
C76 B.n42 VSUBS 0.022144f
C77 B.n43 VSUBS 0.009558f
C78 B.n44 VSUBS 0.009558f
C79 B.n45 VSUBS 0.009558f
C80 B.n46 VSUBS 0.009558f
C81 B.n47 VSUBS 0.009558f
C82 B.n48 VSUBS 0.009558f
C83 B.n49 VSUBS 0.023131f
C84 B.n50 VSUBS 0.009558f
C85 B.n51 VSUBS 0.009558f
C86 B.n52 VSUBS 0.009558f
C87 B.n53 VSUBS 0.009558f
C88 B.n54 VSUBS 0.009558f
C89 B.n55 VSUBS 0.009558f
C90 B.n56 VSUBS 0.009558f
C91 B.n57 VSUBS 0.009558f
C92 B.n58 VSUBS 0.009558f
C93 B.n59 VSUBS 0.009558f
C94 B.n60 VSUBS 0.009558f
C95 B.n61 VSUBS 0.009558f
C96 B.n62 VSUBS 0.009558f
C97 B.n63 VSUBS 0.009558f
C98 B.n64 VSUBS 0.009558f
C99 B.n65 VSUBS 0.009558f
C100 B.n66 VSUBS 0.009558f
C101 B.n67 VSUBS 0.009558f
C102 B.n68 VSUBS 0.009558f
C103 B.n69 VSUBS 0.009558f
C104 B.n70 VSUBS 0.009558f
C105 B.n71 VSUBS 0.009558f
C106 B.n72 VSUBS 0.009558f
C107 B.n73 VSUBS 0.009558f
C108 B.n74 VSUBS 0.009558f
C109 B.n75 VSUBS 0.009558f
C110 B.n76 VSUBS 0.009558f
C111 B.n77 VSUBS 0.009558f
C112 B.n78 VSUBS 0.009558f
C113 B.n79 VSUBS 0.009558f
C114 B.n80 VSUBS 0.009558f
C115 B.n81 VSUBS 0.009558f
C116 B.n82 VSUBS 0.009558f
C117 B.n83 VSUBS 0.009558f
C118 B.n84 VSUBS 0.009558f
C119 B.n85 VSUBS 0.009558f
C120 B.n86 VSUBS 0.009558f
C121 B.n87 VSUBS 0.009558f
C122 B.n88 VSUBS 0.009558f
C123 B.n89 VSUBS 0.009558f
C124 B.n90 VSUBS 0.009558f
C125 B.n91 VSUBS 0.009558f
C126 B.n92 VSUBS 0.009558f
C127 B.n93 VSUBS 0.022967f
C128 B.n94 VSUBS 0.009558f
C129 B.n95 VSUBS 0.009558f
C130 B.n96 VSUBS 0.009558f
C131 B.n97 VSUBS 0.009558f
C132 B.n98 VSUBS 0.009558f
C133 B.n99 VSUBS 0.009558f
C134 B.n100 VSUBS 0.009558f
C135 B.n101 VSUBS 0.008995f
C136 B.n102 VSUBS 0.009558f
C137 B.n103 VSUBS 0.009558f
C138 B.n104 VSUBS 0.009558f
C139 B.n105 VSUBS 0.009558f
C140 B.n106 VSUBS 0.009558f
C141 B.t2 VSUBS 0.067822f
C142 B.t1 VSUBS 0.100816f
C143 B.t0 VSUBS 0.82529f
C144 B.n107 VSUBS 0.171884f
C145 B.n108 VSUBS 0.143313f
C146 B.n109 VSUBS 0.009558f
C147 B.n110 VSUBS 0.009558f
C148 B.n111 VSUBS 0.009558f
C149 B.n112 VSUBS 0.009558f
C150 B.n113 VSUBS 0.009558f
C151 B.n114 VSUBS 0.009558f
C152 B.n115 VSUBS 0.009558f
C153 B.n116 VSUBS 0.023131f
C154 B.n117 VSUBS 0.009558f
C155 B.n118 VSUBS 0.009558f
C156 B.n119 VSUBS 0.009558f
C157 B.n120 VSUBS 0.009558f
C158 B.n121 VSUBS 0.009558f
C159 B.n122 VSUBS 0.009558f
C160 B.n123 VSUBS 0.009558f
C161 B.n124 VSUBS 0.009558f
C162 B.n125 VSUBS 0.009558f
C163 B.n126 VSUBS 0.009558f
C164 B.n127 VSUBS 0.009558f
C165 B.n128 VSUBS 0.009558f
C166 B.n129 VSUBS 0.009558f
C167 B.n130 VSUBS 0.009558f
C168 B.n131 VSUBS 0.009558f
C169 B.n132 VSUBS 0.009558f
C170 B.n133 VSUBS 0.009558f
C171 B.n134 VSUBS 0.009558f
C172 B.n135 VSUBS 0.009558f
C173 B.n136 VSUBS 0.009558f
C174 B.n137 VSUBS 0.009558f
C175 B.n138 VSUBS 0.009558f
C176 B.n139 VSUBS 0.009558f
C177 B.n140 VSUBS 0.009558f
C178 B.n141 VSUBS 0.009558f
C179 B.n142 VSUBS 0.009558f
C180 B.n143 VSUBS 0.009558f
C181 B.n144 VSUBS 0.009558f
C182 B.n145 VSUBS 0.009558f
C183 B.n146 VSUBS 0.009558f
C184 B.n147 VSUBS 0.009558f
C185 B.n148 VSUBS 0.009558f
C186 B.n149 VSUBS 0.009558f
C187 B.n150 VSUBS 0.009558f
C188 B.n151 VSUBS 0.009558f
C189 B.n152 VSUBS 0.009558f
C190 B.n153 VSUBS 0.009558f
C191 B.n154 VSUBS 0.009558f
C192 B.n155 VSUBS 0.009558f
C193 B.n156 VSUBS 0.009558f
C194 B.n157 VSUBS 0.009558f
C195 B.n158 VSUBS 0.009558f
C196 B.n159 VSUBS 0.009558f
C197 B.n160 VSUBS 0.009558f
C198 B.n161 VSUBS 0.009558f
C199 B.n162 VSUBS 0.009558f
C200 B.n163 VSUBS 0.009558f
C201 B.n164 VSUBS 0.009558f
C202 B.n165 VSUBS 0.009558f
C203 B.n166 VSUBS 0.009558f
C204 B.n167 VSUBS 0.009558f
C205 B.n168 VSUBS 0.009558f
C206 B.n169 VSUBS 0.009558f
C207 B.n170 VSUBS 0.009558f
C208 B.n171 VSUBS 0.009558f
C209 B.n172 VSUBS 0.009558f
C210 B.n173 VSUBS 0.009558f
C211 B.n174 VSUBS 0.009558f
C212 B.n175 VSUBS 0.009558f
C213 B.n176 VSUBS 0.009558f
C214 B.n177 VSUBS 0.009558f
C215 B.n178 VSUBS 0.009558f
C216 B.n179 VSUBS 0.009558f
C217 B.n180 VSUBS 0.009558f
C218 B.n181 VSUBS 0.009558f
C219 B.n182 VSUBS 0.009558f
C220 B.n183 VSUBS 0.009558f
C221 B.n184 VSUBS 0.009558f
C222 B.n185 VSUBS 0.009558f
C223 B.n186 VSUBS 0.009558f
C224 B.n187 VSUBS 0.009558f
C225 B.n188 VSUBS 0.009558f
C226 B.n189 VSUBS 0.009558f
C227 B.n190 VSUBS 0.009558f
C228 B.n191 VSUBS 0.009558f
C229 B.n192 VSUBS 0.009558f
C230 B.n193 VSUBS 0.009558f
C231 B.n194 VSUBS 0.009558f
C232 B.n195 VSUBS 0.009558f
C233 B.n196 VSUBS 0.009558f
C234 B.n197 VSUBS 0.009558f
C235 B.n198 VSUBS 0.009558f
C236 B.n199 VSUBS 0.021847f
C237 B.n200 VSUBS 0.021847f
C238 B.n201 VSUBS 0.023131f
C239 B.n202 VSUBS 0.009558f
C240 B.n203 VSUBS 0.009558f
C241 B.n204 VSUBS 0.009558f
C242 B.n205 VSUBS 0.009558f
C243 B.n206 VSUBS 0.009558f
C244 B.n207 VSUBS 0.009558f
C245 B.n208 VSUBS 0.009558f
C246 B.n209 VSUBS 0.009558f
C247 B.n210 VSUBS 0.009558f
C248 B.n211 VSUBS 0.009558f
C249 B.n212 VSUBS 0.009558f
C250 B.n213 VSUBS 0.009558f
C251 B.n214 VSUBS 0.009558f
C252 B.n215 VSUBS 0.009558f
C253 B.n216 VSUBS 0.009558f
C254 B.n217 VSUBS 0.009558f
C255 B.n218 VSUBS 0.009558f
C256 B.n219 VSUBS 0.009558f
C257 B.n220 VSUBS 0.009558f
C258 B.n221 VSUBS 0.009558f
C259 B.n222 VSUBS 0.009558f
C260 B.n223 VSUBS 0.009558f
C261 B.n224 VSUBS 0.008995f
C262 B.n225 VSUBS 0.022144f
C263 B.n226 VSUBS 0.005341f
C264 B.n227 VSUBS 0.009558f
C265 B.n228 VSUBS 0.009558f
C266 B.n229 VSUBS 0.009558f
C267 B.n230 VSUBS 0.009558f
C268 B.n231 VSUBS 0.009558f
C269 B.n232 VSUBS 0.009558f
C270 B.n233 VSUBS 0.009558f
C271 B.n234 VSUBS 0.009558f
C272 B.n235 VSUBS 0.009558f
C273 B.n236 VSUBS 0.009558f
C274 B.n237 VSUBS 0.009558f
C275 B.n238 VSUBS 0.009558f
C276 B.t11 VSUBS 0.067823f
C277 B.t10 VSUBS 0.100817f
C278 B.t9 VSUBS 0.82529f
C279 B.n239 VSUBS 0.171883f
C280 B.n240 VSUBS 0.143312f
C281 B.n241 VSUBS 0.022144f
C282 B.n242 VSUBS 0.005341f
C283 B.n243 VSUBS 0.009558f
C284 B.n244 VSUBS 0.009558f
C285 B.n245 VSUBS 0.009558f
C286 B.n246 VSUBS 0.009558f
C287 B.n247 VSUBS 0.009558f
C288 B.n248 VSUBS 0.009558f
C289 B.n249 VSUBS 0.009558f
C290 B.n250 VSUBS 0.009558f
C291 B.n251 VSUBS 0.009558f
C292 B.n252 VSUBS 0.009558f
C293 B.n253 VSUBS 0.009558f
C294 B.n254 VSUBS 0.009558f
C295 B.n255 VSUBS 0.009558f
C296 B.n256 VSUBS 0.009558f
C297 B.n257 VSUBS 0.009558f
C298 B.n258 VSUBS 0.009558f
C299 B.n259 VSUBS 0.009558f
C300 B.n260 VSUBS 0.009558f
C301 B.n261 VSUBS 0.009558f
C302 B.n262 VSUBS 0.009558f
C303 B.n263 VSUBS 0.009558f
C304 B.n264 VSUBS 0.009558f
C305 B.n265 VSUBS 0.009558f
C306 B.n266 VSUBS 0.022011f
C307 B.n267 VSUBS 0.023131f
C308 B.n268 VSUBS 0.021847f
C309 B.n269 VSUBS 0.009558f
C310 B.n270 VSUBS 0.009558f
C311 B.n271 VSUBS 0.009558f
C312 B.n272 VSUBS 0.009558f
C313 B.n273 VSUBS 0.009558f
C314 B.n274 VSUBS 0.009558f
C315 B.n275 VSUBS 0.009558f
C316 B.n276 VSUBS 0.009558f
C317 B.n277 VSUBS 0.009558f
C318 B.n278 VSUBS 0.009558f
C319 B.n279 VSUBS 0.009558f
C320 B.n280 VSUBS 0.009558f
C321 B.n281 VSUBS 0.009558f
C322 B.n282 VSUBS 0.009558f
C323 B.n283 VSUBS 0.009558f
C324 B.n284 VSUBS 0.009558f
C325 B.n285 VSUBS 0.009558f
C326 B.n286 VSUBS 0.009558f
C327 B.n287 VSUBS 0.009558f
C328 B.n288 VSUBS 0.009558f
C329 B.n289 VSUBS 0.009558f
C330 B.n290 VSUBS 0.009558f
C331 B.n291 VSUBS 0.009558f
C332 B.n292 VSUBS 0.009558f
C333 B.n293 VSUBS 0.009558f
C334 B.n294 VSUBS 0.009558f
C335 B.n295 VSUBS 0.009558f
C336 B.n296 VSUBS 0.009558f
C337 B.n297 VSUBS 0.009558f
C338 B.n298 VSUBS 0.009558f
C339 B.n299 VSUBS 0.009558f
C340 B.n300 VSUBS 0.009558f
C341 B.n301 VSUBS 0.009558f
C342 B.n302 VSUBS 0.009558f
C343 B.n303 VSUBS 0.009558f
C344 B.n304 VSUBS 0.009558f
C345 B.n305 VSUBS 0.009558f
C346 B.n306 VSUBS 0.009558f
C347 B.n307 VSUBS 0.009558f
C348 B.n308 VSUBS 0.009558f
C349 B.n309 VSUBS 0.009558f
C350 B.n310 VSUBS 0.009558f
C351 B.n311 VSUBS 0.009558f
C352 B.n312 VSUBS 0.009558f
C353 B.n313 VSUBS 0.009558f
C354 B.n314 VSUBS 0.009558f
C355 B.n315 VSUBS 0.009558f
C356 B.n316 VSUBS 0.009558f
C357 B.n317 VSUBS 0.009558f
C358 B.n318 VSUBS 0.009558f
C359 B.n319 VSUBS 0.009558f
C360 B.n320 VSUBS 0.009558f
C361 B.n321 VSUBS 0.009558f
C362 B.n322 VSUBS 0.009558f
C363 B.n323 VSUBS 0.009558f
C364 B.n324 VSUBS 0.009558f
C365 B.n325 VSUBS 0.009558f
C366 B.n326 VSUBS 0.009558f
C367 B.n327 VSUBS 0.009558f
C368 B.n328 VSUBS 0.009558f
C369 B.n329 VSUBS 0.009558f
C370 B.n330 VSUBS 0.009558f
C371 B.n331 VSUBS 0.009558f
C372 B.n332 VSUBS 0.009558f
C373 B.n333 VSUBS 0.009558f
C374 B.n334 VSUBS 0.009558f
C375 B.n335 VSUBS 0.009558f
C376 B.n336 VSUBS 0.009558f
C377 B.n337 VSUBS 0.009558f
C378 B.n338 VSUBS 0.009558f
C379 B.n339 VSUBS 0.009558f
C380 B.n340 VSUBS 0.009558f
C381 B.n341 VSUBS 0.009558f
C382 B.n342 VSUBS 0.009558f
C383 B.n343 VSUBS 0.009558f
C384 B.n344 VSUBS 0.009558f
C385 B.n345 VSUBS 0.009558f
C386 B.n346 VSUBS 0.009558f
C387 B.n347 VSUBS 0.009558f
C388 B.n348 VSUBS 0.009558f
C389 B.n349 VSUBS 0.009558f
C390 B.n350 VSUBS 0.009558f
C391 B.n351 VSUBS 0.009558f
C392 B.n352 VSUBS 0.009558f
C393 B.n353 VSUBS 0.009558f
C394 B.n354 VSUBS 0.009558f
C395 B.n355 VSUBS 0.009558f
C396 B.n356 VSUBS 0.009558f
C397 B.n357 VSUBS 0.009558f
C398 B.n358 VSUBS 0.009558f
C399 B.n359 VSUBS 0.009558f
C400 B.n360 VSUBS 0.009558f
C401 B.n361 VSUBS 0.009558f
C402 B.n362 VSUBS 0.009558f
C403 B.n363 VSUBS 0.009558f
C404 B.n364 VSUBS 0.009558f
C405 B.n365 VSUBS 0.009558f
C406 B.n366 VSUBS 0.009558f
C407 B.n367 VSUBS 0.009558f
C408 B.n368 VSUBS 0.009558f
C409 B.n369 VSUBS 0.009558f
C410 B.n370 VSUBS 0.009558f
C411 B.n371 VSUBS 0.009558f
C412 B.n372 VSUBS 0.009558f
C413 B.n373 VSUBS 0.009558f
C414 B.n374 VSUBS 0.009558f
C415 B.n375 VSUBS 0.009558f
C416 B.n376 VSUBS 0.009558f
C417 B.n377 VSUBS 0.009558f
C418 B.n378 VSUBS 0.009558f
C419 B.n379 VSUBS 0.009558f
C420 B.n380 VSUBS 0.009558f
C421 B.n381 VSUBS 0.009558f
C422 B.n382 VSUBS 0.009558f
C423 B.n383 VSUBS 0.009558f
C424 B.n384 VSUBS 0.009558f
C425 B.n385 VSUBS 0.009558f
C426 B.n386 VSUBS 0.009558f
C427 B.n387 VSUBS 0.009558f
C428 B.n388 VSUBS 0.009558f
C429 B.n389 VSUBS 0.009558f
C430 B.n390 VSUBS 0.009558f
C431 B.n391 VSUBS 0.009558f
C432 B.n392 VSUBS 0.009558f
C433 B.n393 VSUBS 0.009558f
C434 B.n394 VSUBS 0.009558f
C435 B.n395 VSUBS 0.009558f
C436 B.n396 VSUBS 0.009558f
C437 B.n397 VSUBS 0.009558f
C438 B.n398 VSUBS 0.021847f
C439 B.n399 VSUBS 0.021847f
C440 B.n400 VSUBS 0.023131f
C441 B.n401 VSUBS 0.009558f
C442 B.n402 VSUBS 0.009558f
C443 B.n403 VSUBS 0.009558f
C444 B.n404 VSUBS 0.009558f
C445 B.n405 VSUBS 0.009558f
C446 B.n406 VSUBS 0.009558f
C447 B.n407 VSUBS 0.009558f
C448 B.n408 VSUBS 0.009558f
C449 B.n409 VSUBS 0.009558f
C450 B.n410 VSUBS 0.009558f
C451 B.n411 VSUBS 0.009558f
C452 B.n412 VSUBS 0.009558f
C453 B.n413 VSUBS 0.009558f
C454 B.n414 VSUBS 0.009558f
C455 B.n415 VSUBS 0.009558f
C456 B.n416 VSUBS 0.009558f
C457 B.n417 VSUBS 0.009558f
C458 B.n418 VSUBS 0.009558f
C459 B.n419 VSUBS 0.009558f
C460 B.n420 VSUBS 0.009558f
C461 B.n421 VSUBS 0.009558f
C462 B.n422 VSUBS 0.008995f
C463 B.n423 VSUBS 0.009558f
C464 B.n424 VSUBS 0.009558f
C465 B.n425 VSUBS 0.009558f
C466 B.n426 VSUBS 0.009558f
C467 B.n427 VSUBS 0.009558f
C468 B.n428 VSUBS 0.009558f
C469 B.n429 VSUBS 0.009558f
C470 B.n430 VSUBS 0.009558f
C471 B.n431 VSUBS 0.009558f
C472 B.n432 VSUBS 0.009558f
C473 B.n433 VSUBS 0.009558f
C474 B.n434 VSUBS 0.009558f
C475 B.n435 VSUBS 0.009558f
C476 B.n436 VSUBS 0.009558f
C477 B.n437 VSUBS 0.009558f
C478 B.n438 VSUBS 0.005341f
C479 B.n439 VSUBS 0.022144f
C480 B.n440 VSUBS 0.008995f
C481 B.n441 VSUBS 0.009558f
C482 B.n442 VSUBS 0.009558f
C483 B.n443 VSUBS 0.009558f
C484 B.n444 VSUBS 0.009558f
C485 B.n445 VSUBS 0.009558f
C486 B.n446 VSUBS 0.009558f
C487 B.n447 VSUBS 0.009558f
C488 B.n448 VSUBS 0.009558f
C489 B.n449 VSUBS 0.009558f
C490 B.n450 VSUBS 0.009558f
C491 B.n451 VSUBS 0.009558f
C492 B.n452 VSUBS 0.009558f
C493 B.n453 VSUBS 0.009558f
C494 B.n454 VSUBS 0.009558f
C495 B.n455 VSUBS 0.009558f
C496 B.n456 VSUBS 0.009558f
C497 B.n457 VSUBS 0.009558f
C498 B.n458 VSUBS 0.009558f
C499 B.n459 VSUBS 0.009558f
C500 B.n460 VSUBS 0.009558f
C501 B.n461 VSUBS 0.009558f
C502 B.n462 VSUBS 0.023131f
C503 B.n463 VSUBS 0.023131f
C504 B.n464 VSUBS 0.021847f
C505 B.n465 VSUBS 0.009558f
C506 B.n466 VSUBS 0.009558f
C507 B.n467 VSUBS 0.009558f
C508 B.n468 VSUBS 0.009558f
C509 B.n469 VSUBS 0.009558f
C510 B.n470 VSUBS 0.009558f
C511 B.n471 VSUBS 0.009558f
C512 B.n472 VSUBS 0.009558f
C513 B.n473 VSUBS 0.009558f
C514 B.n474 VSUBS 0.009558f
C515 B.n475 VSUBS 0.009558f
C516 B.n476 VSUBS 0.009558f
C517 B.n477 VSUBS 0.009558f
C518 B.n478 VSUBS 0.009558f
C519 B.n479 VSUBS 0.009558f
C520 B.n480 VSUBS 0.009558f
C521 B.n481 VSUBS 0.009558f
C522 B.n482 VSUBS 0.009558f
C523 B.n483 VSUBS 0.009558f
C524 B.n484 VSUBS 0.009558f
C525 B.n485 VSUBS 0.009558f
C526 B.n486 VSUBS 0.009558f
C527 B.n487 VSUBS 0.009558f
C528 B.n488 VSUBS 0.009558f
C529 B.n489 VSUBS 0.009558f
C530 B.n490 VSUBS 0.009558f
C531 B.n491 VSUBS 0.009558f
C532 B.n492 VSUBS 0.009558f
C533 B.n493 VSUBS 0.009558f
C534 B.n494 VSUBS 0.009558f
C535 B.n495 VSUBS 0.009558f
C536 B.n496 VSUBS 0.009558f
C537 B.n497 VSUBS 0.009558f
C538 B.n498 VSUBS 0.009558f
C539 B.n499 VSUBS 0.009558f
C540 B.n500 VSUBS 0.009558f
C541 B.n501 VSUBS 0.009558f
C542 B.n502 VSUBS 0.009558f
C543 B.n503 VSUBS 0.009558f
C544 B.n504 VSUBS 0.009558f
C545 B.n505 VSUBS 0.009558f
C546 B.n506 VSUBS 0.009558f
C547 B.n507 VSUBS 0.009558f
C548 B.n508 VSUBS 0.009558f
C549 B.n509 VSUBS 0.009558f
C550 B.n510 VSUBS 0.009558f
C551 B.n511 VSUBS 0.009558f
C552 B.n512 VSUBS 0.009558f
C553 B.n513 VSUBS 0.009558f
C554 B.n514 VSUBS 0.009558f
C555 B.n515 VSUBS 0.009558f
C556 B.n516 VSUBS 0.009558f
C557 B.n517 VSUBS 0.009558f
C558 B.n518 VSUBS 0.009558f
C559 B.n519 VSUBS 0.009558f
C560 B.n520 VSUBS 0.009558f
C561 B.n521 VSUBS 0.009558f
C562 B.n522 VSUBS 0.009558f
C563 B.n523 VSUBS 0.009558f
C564 B.n524 VSUBS 0.009558f
C565 B.n525 VSUBS 0.009558f
C566 B.n526 VSUBS 0.009558f
C567 B.n527 VSUBS 0.012472f
C568 B.n528 VSUBS 0.013286f
C569 B.n529 VSUBS 0.026421f
C570 VDD2.t2 VSUBS 0.055686f
C571 VDD2.t3 VSUBS 0.055686f
C572 VDD2.n0 VSUBS 0.528357f
C573 VDD2.t0 VSUBS 0.055686f
C574 VDD2.t1 VSUBS 0.055686f
C575 VDD2.n1 VSUBS 0.304304f
C576 VDD2.n2 VSUBS 2.70518f
C577 VN.t0 VSUBS 1.69676f
C578 VN.t1 VSUBS 1.7168f
C579 VN.n0 VSUBS 1.08157f
C580 VN.t3 VSUBS 1.69676f
C581 VN.t2 VSUBS 1.7168f
C582 VN.n1 VSUBS 3.2238f
C583 VDD1.t0 VSUBS 0.053259f
C584 VDD1.t3 VSUBS 0.053259f
C585 VDD1.n0 VSUBS 0.291265f
C586 VDD1.t1 VSUBS 0.053259f
C587 VDD1.t2 VSUBS 0.053259f
C588 VDD1.n1 VSUBS 0.516596f
C589 VTAIL.n0 VSUBS 0.037973f
C590 VTAIL.n1 VSUBS 0.033775f
C591 VTAIL.n2 VSUBS 0.018149f
C592 VTAIL.n3 VSUBS 0.032174f
C593 VTAIL.n4 VSUBS 0.026484f
C594 VTAIL.t2 VSUBS 0.097879f
C595 VTAIL.n5 VSUBS 0.126493f
C596 VTAIL.n6 VSUBS 0.359636f
C597 VTAIL.n7 VSUBS 0.018149f
C598 VTAIL.n8 VSUBS 0.019217f
C599 VTAIL.n9 VSUBS 0.042898f
C600 VTAIL.n10 VSUBS 0.106785f
C601 VTAIL.n11 VSUBS 0.019217f
C602 VTAIL.n12 VSUBS 0.018149f
C603 VTAIL.n13 VSUBS 0.088682f
C604 VTAIL.n14 VSUBS 0.05414f
C605 VTAIL.n15 VSUBS 0.280897f
C606 VTAIL.n16 VSUBS 0.037973f
C607 VTAIL.n17 VSUBS 0.033775f
C608 VTAIL.n18 VSUBS 0.018149f
C609 VTAIL.n19 VSUBS 0.032174f
C610 VTAIL.n20 VSUBS 0.026484f
C611 VTAIL.t5 VSUBS 0.097879f
C612 VTAIL.n21 VSUBS 0.126493f
C613 VTAIL.n22 VSUBS 0.359636f
C614 VTAIL.n23 VSUBS 0.018149f
C615 VTAIL.n24 VSUBS 0.019217f
C616 VTAIL.n25 VSUBS 0.042898f
C617 VTAIL.n26 VSUBS 0.106785f
C618 VTAIL.n27 VSUBS 0.019217f
C619 VTAIL.n28 VSUBS 0.018149f
C620 VTAIL.n29 VSUBS 0.088682f
C621 VTAIL.n30 VSUBS 0.05414f
C622 VTAIL.n31 VSUBS 0.463142f
C623 VTAIL.n32 VSUBS 0.037973f
C624 VTAIL.n33 VSUBS 0.033775f
C625 VTAIL.n34 VSUBS 0.018149f
C626 VTAIL.n35 VSUBS 0.032174f
C627 VTAIL.n36 VSUBS 0.026484f
C628 VTAIL.t6 VSUBS 0.097879f
C629 VTAIL.n37 VSUBS 0.126493f
C630 VTAIL.n38 VSUBS 0.359636f
C631 VTAIL.n39 VSUBS 0.018149f
C632 VTAIL.n40 VSUBS 0.019217f
C633 VTAIL.n41 VSUBS 0.042898f
C634 VTAIL.n42 VSUBS 0.106785f
C635 VTAIL.n43 VSUBS 0.019217f
C636 VTAIL.n44 VSUBS 0.018149f
C637 VTAIL.n45 VSUBS 0.088682f
C638 VTAIL.n46 VSUBS 0.05414f
C639 VTAIL.n47 VSUBS 1.56226f
C640 VTAIL.n48 VSUBS 0.037973f
C641 VTAIL.n49 VSUBS 0.033775f
C642 VTAIL.n50 VSUBS 0.018149f
C643 VTAIL.n51 VSUBS 0.032174f
C644 VTAIL.n52 VSUBS 0.026484f
C645 VTAIL.t0 VSUBS 0.097879f
C646 VTAIL.n53 VSUBS 0.126493f
C647 VTAIL.n54 VSUBS 0.359636f
C648 VTAIL.n55 VSUBS 0.018149f
C649 VTAIL.n56 VSUBS 0.019217f
C650 VTAIL.n57 VSUBS 0.042898f
C651 VTAIL.n58 VSUBS 0.106785f
C652 VTAIL.n59 VSUBS 0.019217f
C653 VTAIL.n60 VSUBS 0.018149f
C654 VTAIL.n61 VSUBS 0.088682f
C655 VTAIL.n62 VSUBS 0.05414f
C656 VTAIL.n63 VSUBS 1.56226f
C657 VTAIL.n64 VSUBS 0.037973f
C658 VTAIL.n65 VSUBS 0.033775f
C659 VTAIL.n66 VSUBS 0.018149f
C660 VTAIL.n67 VSUBS 0.032174f
C661 VTAIL.n68 VSUBS 0.026484f
C662 VTAIL.t1 VSUBS 0.097879f
C663 VTAIL.n69 VSUBS 0.126493f
C664 VTAIL.n70 VSUBS 0.359636f
C665 VTAIL.n71 VSUBS 0.018149f
C666 VTAIL.n72 VSUBS 0.019217f
C667 VTAIL.n73 VSUBS 0.042898f
C668 VTAIL.n74 VSUBS 0.106785f
C669 VTAIL.n75 VSUBS 0.019217f
C670 VTAIL.n76 VSUBS 0.018149f
C671 VTAIL.n77 VSUBS 0.088682f
C672 VTAIL.n78 VSUBS 0.05414f
C673 VTAIL.n79 VSUBS 0.463142f
C674 VTAIL.n80 VSUBS 0.037973f
C675 VTAIL.n81 VSUBS 0.033775f
C676 VTAIL.n82 VSUBS 0.018149f
C677 VTAIL.n83 VSUBS 0.032174f
C678 VTAIL.n84 VSUBS 0.026484f
C679 VTAIL.t4 VSUBS 0.097879f
C680 VTAIL.n85 VSUBS 0.126493f
C681 VTAIL.n86 VSUBS 0.359636f
C682 VTAIL.n87 VSUBS 0.018149f
C683 VTAIL.n88 VSUBS 0.019217f
C684 VTAIL.n89 VSUBS 0.042898f
C685 VTAIL.n90 VSUBS 0.106785f
C686 VTAIL.n91 VSUBS 0.019217f
C687 VTAIL.n92 VSUBS 0.018149f
C688 VTAIL.n93 VSUBS 0.088682f
C689 VTAIL.n94 VSUBS 0.05414f
C690 VTAIL.n95 VSUBS 0.463142f
C691 VTAIL.n96 VSUBS 0.037973f
C692 VTAIL.n97 VSUBS 0.033775f
C693 VTAIL.n98 VSUBS 0.018149f
C694 VTAIL.n99 VSUBS 0.032174f
C695 VTAIL.n100 VSUBS 0.026484f
C696 VTAIL.t7 VSUBS 0.097879f
C697 VTAIL.n101 VSUBS 0.126493f
C698 VTAIL.n102 VSUBS 0.359636f
C699 VTAIL.n103 VSUBS 0.018149f
C700 VTAIL.n104 VSUBS 0.019217f
C701 VTAIL.n105 VSUBS 0.042898f
C702 VTAIL.n106 VSUBS 0.106785f
C703 VTAIL.n107 VSUBS 0.019217f
C704 VTAIL.n108 VSUBS 0.018149f
C705 VTAIL.n109 VSUBS 0.088682f
C706 VTAIL.n110 VSUBS 0.05414f
C707 VTAIL.n111 VSUBS 1.56226f
C708 VTAIL.n112 VSUBS 0.037973f
C709 VTAIL.n113 VSUBS 0.033775f
C710 VTAIL.n114 VSUBS 0.018149f
C711 VTAIL.n115 VSUBS 0.032174f
C712 VTAIL.n116 VSUBS 0.026484f
C713 VTAIL.t3 VSUBS 0.097879f
C714 VTAIL.n117 VSUBS 0.126493f
C715 VTAIL.n118 VSUBS 0.359636f
C716 VTAIL.n119 VSUBS 0.018149f
C717 VTAIL.n120 VSUBS 0.019217f
C718 VTAIL.n121 VSUBS 0.042898f
C719 VTAIL.n122 VSUBS 0.106785f
C720 VTAIL.n123 VSUBS 0.019217f
C721 VTAIL.n124 VSUBS 0.018149f
C722 VTAIL.n125 VSUBS 0.088682f
C723 VTAIL.n126 VSUBS 0.05414f
C724 VTAIL.n127 VSUBS 1.36735f
C725 VP.t1 VSUBS 1.26995f
C726 VP.n0 VSUBS 0.651236f
C727 VP.n1 VSUBS 0.040709f
C728 VP.n2 VSUBS 0.080909f
C729 VP.n3 VSUBS 0.040709f
C730 VP.n4 VSUBS 0.075872f
C731 VP.t3 VSUBS 1.77494f
C732 VP.t0 VSUBS 1.75423f
C733 VP.n5 VSUBS 3.31576f
C734 VP.n6 VSUBS 2.01845f
C735 VP.t2 VSUBS 1.26995f
C736 VP.n7 VSUBS 0.651236f
C737 VP.n8 VSUBS 0.039163f
C738 VP.n9 VSUBS 0.065704f
C739 VP.n10 VSUBS 0.040709f
C740 VP.n11 VSUBS 0.040709f
C741 VP.n12 VSUBS 0.075872f
C742 VP.n13 VSUBS 0.080909f
C743 VP.n14 VSUBS 0.03291f
C744 VP.n15 VSUBS 0.040709f
C745 VP.n16 VSUBS 0.040709f
C746 VP.n17 VSUBS 0.040709f
C747 VP.n18 VSUBS 0.075872f
C748 VP.n19 VSUBS 0.075872f
C749 VP.n20 VSUBS 0.039163f
C750 VP.n21 VSUBS 0.065704f
C751 VP.n22 VSUBS 0.1252f
.ends

