* NGSPICE file created from diff_pair_sample_0048.ext - technology: sky130A

.subckt diff_pair_sample_0048 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=0 ps=0 w=14.4 l=2.72
X1 VTAIL.t7 VP.t0 VDD1.t1 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=2.376 ps=14.73 w=14.4 l=2.72
X2 VDD1.t0 VP.t1 VTAIL.t6 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=2.376 pd=14.73 as=5.616 ps=29.58 w=14.4 l=2.72
X3 VTAIL.t0 VN.t0 VDD2.t3 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=2.376 ps=14.73 w=14.4 l=2.72
X4 VDD2.t2 VN.t1 VTAIL.t1 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=2.376 pd=14.73 as=5.616 ps=29.58 w=14.4 l=2.72
X5 VTAIL.t2 VN.t2 VDD2.t1 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=2.376 ps=14.73 w=14.4 l=2.72
X6 VTAIL.t5 VP.t2 VDD1.t3 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=2.376 ps=14.73 w=14.4 l=2.72
X7 VDD2.t0 VN.t3 VTAIL.t3 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=2.376 pd=14.73 as=5.616 ps=29.58 w=14.4 l=2.72
X8 VDD1.t2 VP.t3 VTAIL.t4 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=2.376 pd=14.73 as=5.616 ps=29.58 w=14.4 l=2.72
X9 B.t8 B.t6 B.t7 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=0 ps=0 w=14.4 l=2.72
X10 B.t5 B.t3 B.t4 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=0 ps=0 w=14.4 l=2.72
X11 B.t2 B.t0 B.t1 w_n2800_n3848# sky130_fd_pr__pfet_01v8 ad=5.616 pd=29.58 as=0 ps=0 w=14.4 l=2.72
R0 B.n508 B.n77 585
R1 B.n510 B.n509 585
R2 B.n511 B.n76 585
R3 B.n513 B.n512 585
R4 B.n514 B.n75 585
R5 B.n516 B.n515 585
R6 B.n517 B.n74 585
R7 B.n519 B.n518 585
R8 B.n520 B.n73 585
R9 B.n522 B.n521 585
R10 B.n523 B.n72 585
R11 B.n525 B.n524 585
R12 B.n526 B.n71 585
R13 B.n528 B.n527 585
R14 B.n529 B.n70 585
R15 B.n531 B.n530 585
R16 B.n532 B.n69 585
R17 B.n534 B.n533 585
R18 B.n535 B.n68 585
R19 B.n537 B.n536 585
R20 B.n538 B.n67 585
R21 B.n540 B.n539 585
R22 B.n541 B.n66 585
R23 B.n543 B.n542 585
R24 B.n544 B.n65 585
R25 B.n546 B.n545 585
R26 B.n547 B.n64 585
R27 B.n549 B.n548 585
R28 B.n550 B.n63 585
R29 B.n552 B.n551 585
R30 B.n553 B.n62 585
R31 B.n555 B.n554 585
R32 B.n556 B.n61 585
R33 B.n558 B.n557 585
R34 B.n559 B.n60 585
R35 B.n561 B.n560 585
R36 B.n562 B.n59 585
R37 B.n564 B.n563 585
R38 B.n565 B.n58 585
R39 B.n567 B.n566 585
R40 B.n568 B.n57 585
R41 B.n570 B.n569 585
R42 B.n571 B.n56 585
R43 B.n573 B.n572 585
R44 B.n574 B.n55 585
R45 B.n576 B.n575 585
R46 B.n577 B.n54 585
R47 B.n579 B.n578 585
R48 B.n580 B.n51 585
R49 B.n583 B.n582 585
R50 B.n584 B.n50 585
R51 B.n586 B.n585 585
R52 B.n587 B.n49 585
R53 B.n589 B.n588 585
R54 B.n590 B.n48 585
R55 B.n592 B.n591 585
R56 B.n593 B.n47 585
R57 B.n595 B.n594 585
R58 B.n597 B.n596 585
R59 B.n598 B.n43 585
R60 B.n600 B.n599 585
R61 B.n601 B.n42 585
R62 B.n603 B.n602 585
R63 B.n604 B.n41 585
R64 B.n606 B.n605 585
R65 B.n607 B.n40 585
R66 B.n609 B.n608 585
R67 B.n610 B.n39 585
R68 B.n612 B.n611 585
R69 B.n613 B.n38 585
R70 B.n615 B.n614 585
R71 B.n616 B.n37 585
R72 B.n618 B.n617 585
R73 B.n619 B.n36 585
R74 B.n621 B.n620 585
R75 B.n622 B.n35 585
R76 B.n624 B.n623 585
R77 B.n625 B.n34 585
R78 B.n627 B.n626 585
R79 B.n628 B.n33 585
R80 B.n630 B.n629 585
R81 B.n631 B.n32 585
R82 B.n633 B.n632 585
R83 B.n634 B.n31 585
R84 B.n636 B.n635 585
R85 B.n637 B.n30 585
R86 B.n639 B.n638 585
R87 B.n640 B.n29 585
R88 B.n642 B.n641 585
R89 B.n643 B.n28 585
R90 B.n645 B.n644 585
R91 B.n646 B.n27 585
R92 B.n648 B.n647 585
R93 B.n649 B.n26 585
R94 B.n651 B.n650 585
R95 B.n652 B.n25 585
R96 B.n654 B.n653 585
R97 B.n655 B.n24 585
R98 B.n657 B.n656 585
R99 B.n658 B.n23 585
R100 B.n660 B.n659 585
R101 B.n661 B.n22 585
R102 B.n663 B.n662 585
R103 B.n664 B.n21 585
R104 B.n666 B.n665 585
R105 B.n667 B.n20 585
R106 B.n669 B.n668 585
R107 B.n507 B.n506 585
R108 B.n505 B.n78 585
R109 B.n504 B.n503 585
R110 B.n502 B.n79 585
R111 B.n501 B.n500 585
R112 B.n499 B.n80 585
R113 B.n498 B.n497 585
R114 B.n496 B.n81 585
R115 B.n495 B.n494 585
R116 B.n493 B.n82 585
R117 B.n492 B.n491 585
R118 B.n490 B.n83 585
R119 B.n489 B.n488 585
R120 B.n487 B.n84 585
R121 B.n486 B.n485 585
R122 B.n484 B.n85 585
R123 B.n483 B.n482 585
R124 B.n481 B.n86 585
R125 B.n480 B.n479 585
R126 B.n478 B.n87 585
R127 B.n477 B.n476 585
R128 B.n475 B.n88 585
R129 B.n474 B.n473 585
R130 B.n472 B.n89 585
R131 B.n471 B.n470 585
R132 B.n469 B.n90 585
R133 B.n468 B.n467 585
R134 B.n466 B.n91 585
R135 B.n465 B.n464 585
R136 B.n463 B.n92 585
R137 B.n462 B.n461 585
R138 B.n460 B.n93 585
R139 B.n459 B.n458 585
R140 B.n457 B.n94 585
R141 B.n456 B.n455 585
R142 B.n454 B.n95 585
R143 B.n453 B.n452 585
R144 B.n451 B.n96 585
R145 B.n450 B.n449 585
R146 B.n448 B.n97 585
R147 B.n447 B.n446 585
R148 B.n445 B.n98 585
R149 B.n444 B.n443 585
R150 B.n442 B.n99 585
R151 B.n441 B.n440 585
R152 B.n439 B.n100 585
R153 B.n438 B.n437 585
R154 B.n436 B.n101 585
R155 B.n435 B.n434 585
R156 B.n433 B.n102 585
R157 B.n432 B.n431 585
R158 B.n430 B.n103 585
R159 B.n429 B.n428 585
R160 B.n427 B.n104 585
R161 B.n426 B.n425 585
R162 B.n424 B.n105 585
R163 B.n423 B.n422 585
R164 B.n421 B.n106 585
R165 B.n420 B.n419 585
R166 B.n418 B.n107 585
R167 B.n417 B.n416 585
R168 B.n415 B.n108 585
R169 B.n414 B.n413 585
R170 B.n412 B.n109 585
R171 B.n411 B.n410 585
R172 B.n409 B.n110 585
R173 B.n408 B.n407 585
R174 B.n406 B.n111 585
R175 B.n405 B.n404 585
R176 B.n403 B.n112 585
R177 B.n402 B.n401 585
R178 B.n240 B.n239 585
R179 B.n241 B.n170 585
R180 B.n243 B.n242 585
R181 B.n244 B.n169 585
R182 B.n246 B.n245 585
R183 B.n247 B.n168 585
R184 B.n249 B.n248 585
R185 B.n250 B.n167 585
R186 B.n252 B.n251 585
R187 B.n253 B.n166 585
R188 B.n255 B.n254 585
R189 B.n256 B.n165 585
R190 B.n258 B.n257 585
R191 B.n259 B.n164 585
R192 B.n261 B.n260 585
R193 B.n262 B.n163 585
R194 B.n264 B.n263 585
R195 B.n265 B.n162 585
R196 B.n267 B.n266 585
R197 B.n268 B.n161 585
R198 B.n270 B.n269 585
R199 B.n271 B.n160 585
R200 B.n273 B.n272 585
R201 B.n274 B.n159 585
R202 B.n276 B.n275 585
R203 B.n277 B.n158 585
R204 B.n279 B.n278 585
R205 B.n280 B.n157 585
R206 B.n282 B.n281 585
R207 B.n283 B.n156 585
R208 B.n285 B.n284 585
R209 B.n286 B.n155 585
R210 B.n288 B.n287 585
R211 B.n289 B.n154 585
R212 B.n291 B.n290 585
R213 B.n292 B.n153 585
R214 B.n294 B.n293 585
R215 B.n295 B.n152 585
R216 B.n297 B.n296 585
R217 B.n298 B.n151 585
R218 B.n300 B.n299 585
R219 B.n301 B.n150 585
R220 B.n303 B.n302 585
R221 B.n304 B.n149 585
R222 B.n306 B.n305 585
R223 B.n307 B.n148 585
R224 B.n309 B.n308 585
R225 B.n310 B.n147 585
R226 B.n312 B.n311 585
R227 B.n314 B.n313 585
R228 B.n315 B.n143 585
R229 B.n317 B.n316 585
R230 B.n318 B.n142 585
R231 B.n320 B.n319 585
R232 B.n321 B.n141 585
R233 B.n323 B.n322 585
R234 B.n324 B.n140 585
R235 B.n326 B.n325 585
R236 B.n328 B.n137 585
R237 B.n330 B.n329 585
R238 B.n331 B.n136 585
R239 B.n333 B.n332 585
R240 B.n334 B.n135 585
R241 B.n336 B.n335 585
R242 B.n337 B.n134 585
R243 B.n339 B.n338 585
R244 B.n340 B.n133 585
R245 B.n342 B.n341 585
R246 B.n343 B.n132 585
R247 B.n345 B.n344 585
R248 B.n346 B.n131 585
R249 B.n348 B.n347 585
R250 B.n349 B.n130 585
R251 B.n351 B.n350 585
R252 B.n352 B.n129 585
R253 B.n354 B.n353 585
R254 B.n355 B.n128 585
R255 B.n357 B.n356 585
R256 B.n358 B.n127 585
R257 B.n360 B.n359 585
R258 B.n361 B.n126 585
R259 B.n363 B.n362 585
R260 B.n364 B.n125 585
R261 B.n366 B.n365 585
R262 B.n367 B.n124 585
R263 B.n369 B.n368 585
R264 B.n370 B.n123 585
R265 B.n372 B.n371 585
R266 B.n373 B.n122 585
R267 B.n375 B.n374 585
R268 B.n376 B.n121 585
R269 B.n378 B.n377 585
R270 B.n379 B.n120 585
R271 B.n381 B.n380 585
R272 B.n382 B.n119 585
R273 B.n384 B.n383 585
R274 B.n385 B.n118 585
R275 B.n387 B.n386 585
R276 B.n388 B.n117 585
R277 B.n390 B.n389 585
R278 B.n391 B.n116 585
R279 B.n393 B.n392 585
R280 B.n394 B.n115 585
R281 B.n396 B.n395 585
R282 B.n397 B.n114 585
R283 B.n399 B.n398 585
R284 B.n400 B.n113 585
R285 B.n238 B.n171 585
R286 B.n237 B.n236 585
R287 B.n235 B.n172 585
R288 B.n234 B.n233 585
R289 B.n232 B.n173 585
R290 B.n231 B.n230 585
R291 B.n229 B.n174 585
R292 B.n228 B.n227 585
R293 B.n226 B.n175 585
R294 B.n225 B.n224 585
R295 B.n223 B.n176 585
R296 B.n222 B.n221 585
R297 B.n220 B.n177 585
R298 B.n219 B.n218 585
R299 B.n217 B.n178 585
R300 B.n216 B.n215 585
R301 B.n214 B.n179 585
R302 B.n213 B.n212 585
R303 B.n211 B.n180 585
R304 B.n210 B.n209 585
R305 B.n208 B.n181 585
R306 B.n207 B.n206 585
R307 B.n205 B.n182 585
R308 B.n204 B.n203 585
R309 B.n202 B.n183 585
R310 B.n201 B.n200 585
R311 B.n199 B.n184 585
R312 B.n198 B.n197 585
R313 B.n196 B.n185 585
R314 B.n195 B.n194 585
R315 B.n193 B.n186 585
R316 B.n192 B.n191 585
R317 B.n190 B.n187 585
R318 B.n189 B.n188 585
R319 B.n2 B.n0 585
R320 B.n721 B.n1 585
R321 B.n720 B.n719 585
R322 B.n718 B.n3 585
R323 B.n717 B.n716 585
R324 B.n715 B.n4 585
R325 B.n714 B.n713 585
R326 B.n712 B.n5 585
R327 B.n711 B.n710 585
R328 B.n709 B.n6 585
R329 B.n708 B.n707 585
R330 B.n706 B.n7 585
R331 B.n705 B.n704 585
R332 B.n703 B.n8 585
R333 B.n702 B.n701 585
R334 B.n700 B.n9 585
R335 B.n699 B.n698 585
R336 B.n697 B.n10 585
R337 B.n696 B.n695 585
R338 B.n694 B.n11 585
R339 B.n693 B.n692 585
R340 B.n691 B.n12 585
R341 B.n690 B.n689 585
R342 B.n688 B.n13 585
R343 B.n687 B.n686 585
R344 B.n685 B.n14 585
R345 B.n684 B.n683 585
R346 B.n682 B.n15 585
R347 B.n681 B.n680 585
R348 B.n679 B.n16 585
R349 B.n678 B.n677 585
R350 B.n676 B.n17 585
R351 B.n675 B.n674 585
R352 B.n673 B.n18 585
R353 B.n672 B.n671 585
R354 B.n670 B.n19 585
R355 B.n723 B.n722 585
R356 B.n240 B.n171 497.305
R357 B.n668 B.n19 497.305
R358 B.n402 B.n113 497.305
R359 B.n506 B.n77 497.305
R360 B.n138 B.t0 335.81
R361 B.n144 B.t3 335.81
R362 B.n44 B.t6 335.81
R363 B.n52 B.t9 335.81
R364 B.n138 B.t2 168.13
R365 B.n52 B.t10 168.13
R366 B.n144 B.t5 168.112
R367 B.n44 B.t7 168.112
R368 B.n236 B.n171 163.367
R369 B.n236 B.n235 163.367
R370 B.n235 B.n234 163.367
R371 B.n234 B.n173 163.367
R372 B.n230 B.n173 163.367
R373 B.n230 B.n229 163.367
R374 B.n229 B.n228 163.367
R375 B.n228 B.n175 163.367
R376 B.n224 B.n175 163.367
R377 B.n224 B.n223 163.367
R378 B.n223 B.n222 163.367
R379 B.n222 B.n177 163.367
R380 B.n218 B.n177 163.367
R381 B.n218 B.n217 163.367
R382 B.n217 B.n216 163.367
R383 B.n216 B.n179 163.367
R384 B.n212 B.n179 163.367
R385 B.n212 B.n211 163.367
R386 B.n211 B.n210 163.367
R387 B.n210 B.n181 163.367
R388 B.n206 B.n181 163.367
R389 B.n206 B.n205 163.367
R390 B.n205 B.n204 163.367
R391 B.n204 B.n183 163.367
R392 B.n200 B.n183 163.367
R393 B.n200 B.n199 163.367
R394 B.n199 B.n198 163.367
R395 B.n198 B.n185 163.367
R396 B.n194 B.n185 163.367
R397 B.n194 B.n193 163.367
R398 B.n193 B.n192 163.367
R399 B.n192 B.n187 163.367
R400 B.n188 B.n187 163.367
R401 B.n188 B.n2 163.367
R402 B.n722 B.n2 163.367
R403 B.n722 B.n721 163.367
R404 B.n721 B.n720 163.367
R405 B.n720 B.n3 163.367
R406 B.n716 B.n3 163.367
R407 B.n716 B.n715 163.367
R408 B.n715 B.n714 163.367
R409 B.n714 B.n5 163.367
R410 B.n710 B.n5 163.367
R411 B.n710 B.n709 163.367
R412 B.n709 B.n708 163.367
R413 B.n708 B.n7 163.367
R414 B.n704 B.n7 163.367
R415 B.n704 B.n703 163.367
R416 B.n703 B.n702 163.367
R417 B.n702 B.n9 163.367
R418 B.n698 B.n9 163.367
R419 B.n698 B.n697 163.367
R420 B.n697 B.n696 163.367
R421 B.n696 B.n11 163.367
R422 B.n692 B.n11 163.367
R423 B.n692 B.n691 163.367
R424 B.n691 B.n690 163.367
R425 B.n690 B.n13 163.367
R426 B.n686 B.n13 163.367
R427 B.n686 B.n685 163.367
R428 B.n685 B.n684 163.367
R429 B.n684 B.n15 163.367
R430 B.n680 B.n15 163.367
R431 B.n680 B.n679 163.367
R432 B.n679 B.n678 163.367
R433 B.n678 B.n17 163.367
R434 B.n674 B.n17 163.367
R435 B.n674 B.n673 163.367
R436 B.n673 B.n672 163.367
R437 B.n672 B.n19 163.367
R438 B.n241 B.n240 163.367
R439 B.n242 B.n241 163.367
R440 B.n242 B.n169 163.367
R441 B.n246 B.n169 163.367
R442 B.n247 B.n246 163.367
R443 B.n248 B.n247 163.367
R444 B.n248 B.n167 163.367
R445 B.n252 B.n167 163.367
R446 B.n253 B.n252 163.367
R447 B.n254 B.n253 163.367
R448 B.n254 B.n165 163.367
R449 B.n258 B.n165 163.367
R450 B.n259 B.n258 163.367
R451 B.n260 B.n259 163.367
R452 B.n260 B.n163 163.367
R453 B.n264 B.n163 163.367
R454 B.n265 B.n264 163.367
R455 B.n266 B.n265 163.367
R456 B.n266 B.n161 163.367
R457 B.n270 B.n161 163.367
R458 B.n271 B.n270 163.367
R459 B.n272 B.n271 163.367
R460 B.n272 B.n159 163.367
R461 B.n276 B.n159 163.367
R462 B.n277 B.n276 163.367
R463 B.n278 B.n277 163.367
R464 B.n278 B.n157 163.367
R465 B.n282 B.n157 163.367
R466 B.n283 B.n282 163.367
R467 B.n284 B.n283 163.367
R468 B.n284 B.n155 163.367
R469 B.n288 B.n155 163.367
R470 B.n289 B.n288 163.367
R471 B.n290 B.n289 163.367
R472 B.n290 B.n153 163.367
R473 B.n294 B.n153 163.367
R474 B.n295 B.n294 163.367
R475 B.n296 B.n295 163.367
R476 B.n296 B.n151 163.367
R477 B.n300 B.n151 163.367
R478 B.n301 B.n300 163.367
R479 B.n302 B.n301 163.367
R480 B.n302 B.n149 163.367
R481 B.n306 B.n149 163.367
R482 B.n307 B.n306 163.367
R483 B.n308 B.n307 163.367
R484 B.n308 B.n147 163.367
R485 B.n312 B.n147 163.367
R486 B.n313 B.n312 163.367
R487 B.n313 B.n143 163.367
R488 B.n317 B.n143 163.367
R489 B.n318 B.n317 163.367
R490 B.n319 B.n318 163.367
R491 B.n319 B.n141 163.367
R492 B.n323 B.n141 163.367
R493 B.n324 B.n323 163.367
R494 B.n325 B.n324 163.367
R495 B.n325 B.n137 163.367
R496 B.n330 B.n137 163.367
R497 B.n331 B.n330 163.367
R498 B.n332 B.n331 163.367
R499 B.n332 B.n135 163.367
R500 B.n336 B.n135 163.367
R501 B.n337 B.n336 163.367
R502 B.n338 B.n337 163.367
R503 B.n338 B.n133 163.367
R504 B.n342 B.n133 163.367
R505 B.n343 B.n342 163.367
R506 B.n344 B.n343 163.367
R507 B.n344 B.n131 163.367
R508 B.n348 B.n131 163.367
R509 B.n349 B.n348 163.367
R510 B.n350 B.n349 163.367
R511 B.n350 B.n129 163.367
R512 B.n354 B.n129 163.367
R513 B.n355 B.n354 163.367
R514 B.n356 B.n355 163.367
R515 B.n356 B.n127 163.367
R516 B.n360 B.n127 163.367
R517 B.n361 B.n360 163.367
R518 B.n362 B.n361 163.367
R519 B.n362 B.n125 163.367
R520 B.n366 B.n125 163.367
R521 B.n367 B.n366 163.367
R522 B.n368 B.n367 163.367
R523 B.n368 B.n123 163.367
R524 B.n372 B.n123 163.367
R525 B.n373 B.n372 163.367
R526 B.n374 B.n373 163.367
R527 B.n374 B.n121 163.367
R528 B.n378 B.n121 163.367
R529 B.n379 B.n378 163.367
R530 B.n380 B.n379 163.367
R531 B.n380 B.n119 163.367
R532 B.n384 B.n119 163.367
R533 B.n385 B.n384 163.367
R534 B.n386 B.n385 163.367
R535 B.n386 B.n117 163.367
R536 B.n390 B.n117 163.367
R537 B.n391 B.n390 163.367
R538 B.n392 B.n391 163.367
R539 B.n392 B.n115 163.367
R540 B.n396 B.n115 163.367
R541 B.n397 B.n396 163.367
R542 B.n398 B.n397 163.367
R543 B.n398 B.n113 163.367
R544 B.n403 B.n402 163.367
R545 B.n404 B.n403 163.367
R546 B.n404 B.n111 163.367
R547 B.n408 B.n111 163.367
R548 B.n409 B.n408 163.367
R549 B.n410 B.n409 163.367
R550 B.n410 B.n109 163.367
R551 B.n414 B.n109 163.367
R552 B.n415 B.n414 163.367
R553 B.n416 B.n415 163.367
R554 B.n416 B.n107 163.367
R555 B.n420 B.n107 163.367
R556 B.n421 B.n420 163.367
R557 B.n422 B.n421 163.367
R558 B.n422 B.n105 163.367
R559 B.n426 B.n105 163.367
R560 B.n427 B.n426 163.367
R561 B.n428 B.n427 163.367
R562 B.n428 B.n103 163.367
R563 B.n432 B.n103 163.367
R564 B.n433 B.n432 163.367
R565 B.n434 B.n433 163.367
R566 B.n434 B.n101 163.367
R567 B.n438 B.n101 163.367
R568 B.n439 B.n438 163.367
R569 B.n440 B.n439 163.367
R570 B.n440 B.n99 163.367
R571 B.n444 B.n99 163.367
R572 B.n445 B.n444 163.367
R573 B.n446 B.n445 163.367
R574 B.n446 B.n97 163.367
R575 B.n450 B.n97 163.367
R576 B.n451 B.n450 163.367
R577 B.n452 B.n451 163.367
R578 B.n452 B.n95 163.367
R579 B.n456 B.n95 163.367
R580 B.n457 B.n456 163.367
R581 B.n458 B.n457 163.367
R582 B.n458 B.n93 163.367
R583 B.n462 B.n93 163.367
R584 B.n463 B.n462 163.367
R585 B.n464 B.n463 163.367
R586 B.n464 B.n91 163.367
R587 B.n468 B.n91 163.367
R588 B.n469 B.n468 163.367
R589 B.n470 B.n469 163.367
R590 B.n470 B.n89 163.367
R591 B.n474 B.n89 163.367
R592 B.n475 B.n474 163.367
R593 B.n476 B.n475 163.367
R594 B.n476 B.n87 163.367
R595 B.n480 B.n87 163.367
R596 B.n481 B.n480 163.367
R597 B.n482 B.n481 163.367
R598 B.n482 B.n85 163.367
R599 B.n486 B.n85 163.367
R600 B.n487 B.n486 163.367
R601 B.n488 B.n487 163.367
R602 B.n488 B.n83 163.367
R603 B.n492 B.n83 163.367
R604 B.n493 B.n492 163.367
R605 B.n494 B.n493 163.367
R606 B.n494 B.n81 163.367
R607 B.n498 B.n81 163.367
R608 B.n499 B.n498 163.367
R609 B.n500 B.n499 163.367
R610 B.n500 B.n79 163.367
R611 B.n504 B.n79 163.367
R612 B.n505 B.n504 163.367
R613 B.n506 B.n505 163.367
R614 B.n668 B.n667 163.367
R615 B.n667 B.n666 163.367
R616 B.n666 B.n21 163.367
R617 B.n662 B.n21 163.367
R618 B.n662 B.n661 163.367
R619 B.n661 B.n660 163.367
R620 B.n660 B.n23 163.367
R621 B.n656 B.n23 163.367
R622 B.n656 B.n655 163.367
R623 B.n655 B.n654 163.367
R624 B.n654 B.n25 163.367
R625 B.n650 B.n25 163.367
R626 B.n650 B.n649 163.367
R627 B.n649 B.n648 163.367
R628 B.n648 B.n27 163.367
R629 B.n644 B.n27 163.367
R630 B.n644 B.n643 163.367
R631 B.n643 B.n642 163.367
R632 B.n642 B.n29 163.367
R633 B.n638 B.n29 163.367
R634 B.n638 B.n637 163.367
R635 B.n637 B.n636 163.367
R636 B.n636 B.n31 163.367
R637 B.n632 B.n31 163.367
R638 B.n632 B.n631 163.367
R639 B.n631 B.n630 163.367
R640 B.n630 B.n33 163.367
R641 B.n626 B.n33 163.367
R642 B.n626 B.n625 163.367
R643 B.n625 B.n624 163.367
R644 B.n624 B.n35 163.367
R645 B.n620 B.n35 163.367
R646 B.n620 B.n619 163.367
R647 B.n619 B.n618 163.367
R648 B.n618 B.n37 163.367
R649 B.n614 B.n37 163.367
R650 B.n614 B.n613 163.367
R651 B.n613 B.n612 163.367
R652 B.n612 B.n39 163.367
R653 B.n608 B.n39 163.367
R654 B.n608 B.n607 163.367
R655 B.n607 B.n606 163.367
R656 B.n606 B.n41 163.367
R657 B.n602 B.n41 163.367
R658 B.n602 B.n601 163.367
R659 B.n601 B.n600 163.367
R660 B.n600 B.n43 163.367
R661 B.n596 B.n43 163.367
R662 B.n596 B.n595 163.367
R663 B.n595 B.n47 163.367
R664 B.n591 B.n47 163.367
R665 B.n591 B.n590 163.367
R666 B.n590 B.n589 163.367
R667 B.n589 B.n49 163.367
R668 B.n585 B.n49 163.367
R669 B.n585 B.n584 163.367
R670 B.n584 B.n583 163.367
R671 B.n583 B.n51 163.367
R672 B.n578 B.n51 163.367
R673 B.n578 B.n577 163.367
R674 B.n577 B.n576 163.367
R675 B.n576 B.n55 163.367
R676 B.n572 B.n55 163.367
R677 B.n572 B.n571 163.367
R678 B.n571 B.n570 163.367
R679 B.n570 B.n57 163.367
R680 B.n566 B.n57 163.367
R681 B.n566 B.n565 163.367
R682 B.n565 B.n564 163.367
R683 B.n564 B.n59 163.367
R684 B.n560 B.n59 163.367
R685 B.n560 B.n559 163.367
R686 B.n559 B.n558 163.367
R687 B.n558 B.n61 163.367
R688 B.n554 B.n61 163.367
R689 B.n554 B.n553 163.367
R690 B.n553 B.n552 163.367
R691 B.n552 B.n63 163.367
R692 B.n548 B.n63 163.367
R693 B.n548 B.n547 163.367
R694 B.n547 B.n546 163.367
R695 B.n546 B.n65 163.367
R696 B.n542 B.n65 163.367
R697 B.n542 B.n541 163.367
R698 B.n541 B.n540 163.367
R699 B.n540 B.n67 163.367
R700 B.n536 B.n67 163.367
R701 B.n536 B.n535 163.367
R702 B.n535 B.n534 163.367
R703 B.n534 B.n69 163.367
R704 B.n530 B.n69 163.367
R705 B.n530 B.n529 163.367
R706 B.n529 B.n528 163.367
R707 B.n528 B.n71 163.367
R708 B.n524 B.n71 163.367
R709 B.n524 B.n523 163.367
R710 B.n523 B.n522 163.367
R711 B.n522 B.n73 163.367
R712 B.n518 B.n73 163.367
R713 B.n518 B.n517 163.367
R714 B.n517 B.n516 163.367
R715 B.n516 B.n75 163.367
R716 B.n512 B.n75 163.367
R717 B.n512 B.n511 163.367
R718 B.n511 B.n510 163.367
R719 B.n510 B.n77 163.367
R720 B.n139 B.t1 108.978
R721 B.n53 B.t11 108.978
R722 B.n145 B.t4 108.96
R723 B.n45 B.t8 108.96
R724 B.n327 B.n139 59.5399
R725 B.n146 B.n145 59.5399
R726 B.n46 B.n45 59.5399
R727 B.n581 B.n53 59.5399
R728 B.n139 B.n138 59.152
R729 B.n145 B.n144 59.152
R730 B.n45 B.n44 59.152
R731 B.n53 B.n52 59.152
R732 B.n670 B.n669 32.3127
R733 B.n508 B.n507 32.3127
R734 B.n401 B.n400 32.3127
R735 B.n239 B.n238 32.3127
R736 B B.n723 18.0485
R737 B.n669 B.n20 10.6151
R738 B.n665 B.n20 10.6151
R739 B.n665 B.n664 10.6151
R740 B.n664 B.n663 10.6151
R741 B.n663 B.n22 10.6151
R742 B.n659 B.n22 10.6151
R743 B.n659 B.n658 10.6151
R744 B.n658 B.n657 10.6151
R745 B.n657 B.n24 10.6151
R746 B.n653 B.n24 10.6151
R747 B.n653 B.n652 10.6151
R748 B.n652 B.n651 10.6151
R749 B.n651 B.n26 10.6151
R750 B.n647 B.n26 10.6151
R751 B.n647 B.n646 10.6151
R752 B.n646 B.n645 10.6151
R753 B.n645 B.n28 10.6151
R754 B.n641 B.n28 10.6151
R755 B.n641 B.n640 10.6151
R756 B.n640 B.n639 10.6151
R757 B.n639 B.n30 10.6151
R758 B.n635 B.n30 10.6151
R759 B.n635 B.n634 10.6151
R760 B.n634 B.n633 10.6151
R761 B.n633 B.n32 10.6151
R762 B.n629 B.n32 10.6151
R763 B.n629 B.n628 10.6151
R764 B.n628 B.n627 10.6151
R765 B.n627 B.n34 10.6151
R766 B.n623 B.n34 10.6151
R767 B.n623 B.n622 10.6151
R768 B.n622 B.n621 10.6151
R769 B.n621 B.n36 10.6151
R770 B.n617 B.n36 10.6151
R771 B.n617 B.n616 10.6151
R772 B.n616 B.n615 10.6151
R773 B.n615 B.n38 10.6151
R774 B.n611 B.n38 10.6151
R775 B.n611 B.n610 10.6151
R776 B.n610 B.n609 10.6151
R777 B.n609 B.n40 10.6151
R778 B.n605 B.n40 10.6151
R779 B.n605 B.n604 10.6151
R780 B.n604 B.n603 10.6151
R781 B.n603 B.n42 10.6151
R782 B.n599 B.n42 10.6151
R783 B.n599 B.n598 10.6151
R784 B.n598 B.n597 10.6151
R785 B.n594 B.n593 10.6151
R786 B.n593 B.n592 10.6151
R787 B.n592 B.n48 10.6151
R788 B.n588 B.n48 10.6151
R789 B.n588 B.n587 10.6151
R790 B.n587 B.n586 10.6151
R791 B.n586 B.n50 10.6151
R792 B.n582 B.n50 10.6151
R793 B.n580 B.n579 10.6151
R794 B.n579 B.n54 10.6151
R795 B.n575 B.n54 10.6151
R796 B.n575 B.n574 10.6151
R797 B.n574 B.n573 10.6151
R798 B.n573 B.n56 10.6151
R799 B.n569 B.n56 10.6151
R800 B.n569 B.n568 10.6151
R801 B.n568 B.n567 10.6151
R802 B.n567 B.n58 10.6151
R803 B.n563 B.n58 10.6151
R804 B.n563 B.n562 10.6151
R805 B.n562 B.n561 10.6151
R806 B.n561 B.n60 10.6151
R807 B.n557 B.n60 10.6151
R808 B.n557 B.n556 10.6151
R809 B.n556 B.n555 10.6151
R810 B.n555 B.n62 10.6151
R811 B.n551 B.n62 10.6151
R812 B.n551 B.n550 10.6151
R813 B.n550 B.n549 10.6151
R814 B.n549 B.n64 10.6151
R815 B.n545 B.n64 10.6151
R816 B.n545 B.n544 10.6151
R817 B.n544 B.n543 10.6151
R818 B.n543 B.n66 10.6151
R819 B.n539 B.n66 10.6151
R820 B.n539 B.n538 10.6151
R821 B.n538 B.n537 10.6151
R822 B.n537 B.n68 10.6151
R823 B.n533 B.n68 10.6151
R824 B.n533 B.n532 10.6151
R825 B.n532 B.n531 10.6151
R826 B.n531 B.n70 10.6151
R827 B.n527 B.n70 10.6151
R828 B.n527 B.n526 10.6151
R829 B.n526 B.n525 10.6151
R830 B.n525 B.n72 10.6151
R831 B.n521 B.n72 10.6151
R832 B.n521 B.n520 10.6151
R833 B.n520 B.n519 10.6151
R834 B.n519 B.n74 10.6151
R835 B.n515 B.n74 10.6151
R836 B.n515 B.n514 10.6151
R837 B.n514 B.n513 10.6151
R838 B.n513 B.n76 10.6151
R839 B.n509 B.n76 10.6151
R840 B.n509 B.n508 10.6151
R841 B.n401 B.n112 10.6151
R842 B.n405 B.n112 10.6151
R843 B.n406 B.n405 10.6151
R844 B.n407 B.n406 10.6151
R845 B.n407 B.n110 10.6151
R846 B.n411 B.n110 10.6151
R847 B.n412 B.n411 10.6151
R848 B.n413 B.n412 10.6151
R849 B.n413 B.n108 10.6151
R850 B.n417 B.n108 10.6151
R851 B.n418 B.n417 10.6151
R852 B.n419 B.n418 10.6151
R853 B.n419 B.n106 10.6151
R854 B.n423 B.n106 10.6151
R855 B.n424 B.n423 10.6151
R856 B.n425 B.n424 10.6151
R857 B.n425 B.n104 10.6151
R858 B.n429 B.n104 10.6151
R859 B.n430 B.n429 10.6151
R860 B.n431 B.n430 10.6151
R861 B.n431 B.n102 10.6151
R862 B.n435 B.n102 10.6151
R863 B.n436 B.n435 10.6151
R864 B.n437 B.n436 10.6151
R865 B.n437 B.n100 10.6151
R866 B.n441 B.n100 10.6151
R867 B.n442 B.n441 10.6151
R868 B.n443 B.n442 10.6151
R869 B.n443 B.n98 10.6151
R870 B.n447 B.n98 10.6151
R871 B.n448 B.n447 10.6151
R872 B.n449 B.n448 10.6151
R873 B.n449 B.n96 10.6151
R874 B.n453 B.n96 10.6151
R875 B.n454 B.n453 10.6151
R876 B.n455 B.n454 10.6151
R877 B.n455 B.n94 10.6151
R878 B.n459 B.n94 10.6151
R879 B.n460 B.n459 10.6151
R880 B.n461 B.n460 10.6151
R881 B.n461 B.n92 10.6151
R882 B.n465 B.n92 10.6151
R883 B.n466 B.n465 10.6151
R884 B.n467 B.n466 10.6151
R885 B.n467 B.n90 10.6151
R886 B.n471 B.n90 10.6151
R887 B.n472 B.n471 10.6151
R888 B.n473 B.n472 10.6151
R889 B.n473 B.n88 10.6151
R890 B.n477 B.n88 10.6151
R891 B.n478 B.n477 10.6151
R892 B.n479 B.n478 10.6151
R893 B.n479 B.n86 10.6151
R894 B.n483 B.n86 10.6151
R895 B.n484 B.n483 10.6151
R896 B.n485 B.n484 10.6151
R897 B.n485 B.n84 10.6151
R898 B.n489 B.n84 10.6151
R899 B.n490 B.n489 10.6151
R900 B.n491 B.n490 10.6151
R901 B.n491 B.n82 10.6151
R902 B.n495 B.n82 10.6151
R903 B.n496 B.n495 10.6151
R904 B.n497 B.n496 10.6151
R905 B.n497 B.n80 10.6151
R906 B.n501 B.n80 10.6151
R907 B.n502 B.n501 10.6151
R908 B.n503 B.n502 10.6151
R909 B.n503 B.n78 10.6151
R910 B.n507 B.n78 10.6151
R911 B.n239 B.n170 10.6151
R912 B.n243 B.n170 10.6151
R913 B.n244 B.n243 10.6151
R914 B.n245 B.n244 10.6151
R915 B.n245 B.n168 10.6151
R916 B.n249 B.n168 10.6151
R917 B.n250 B.n249 10.6151
R918 B.n251 B.n250 10.6151
R919 B.n251 B.n166 10.6151
R920 B.n255 B.n166 10.6151
R921 B.n256 B.n255 10.6151
R922 B.n257 B.n256 10.6151
R923 B.n257 B.n164 10.6151
R924 B.n261 B.n164 10.6151
R925 B.n262 B.n261 10.6151
R926 B.n263 B.n262 10.6151
R927 B.n263 B.n162 10.6151
R928 B.n267 B.n162 10.6151
R929 B.n268 B.n267 10.6151
R930 B.n269 B.n268 10.6151
R931 B.n269 B.n160 10.6151
R932 B.n273 B.n160 10.6151
R933 B.n274 B.n273 10.6151
R934 B.n275 B.n274 10.6151
R935 B.n275 B.n158 10.6151
R936 B.n279 B.n158 10.6151
R937 B.n280 B.n279 10.6151
R938 B.n281 B.n280 10.6151
R939 B.n281 B.n156 10.6151
R940 B.n285 B.n156 10.6151
R941 B.n286 B.n285 10.6151
R942 B.n287 B.n286 10.6151
R943 B.n287 B.n154 10.6151
R944 B.n291 B.n154 10.6151
R945 B.n292 B.n291 10.6151
R946 B.n293 B.n292 10.6151
R947 B.n293 B.n152 10.6151
R948 B.n297 B.n152 10.6151
R949 B.n298 B.n297 10.6151
R950 B.n299 B.n298 10.6151
R951 B.n299 B.n150 10.6151
R952 B.n303 B.n150 10.6151
R953 B.n304 B.n303 10.6151
R954 B.n305 B.n304 10.6151
R955 B.n305 B.n148 10.6151
R956 B.n309 B.n148 10.6151
R957 B.n310 B.n309 10.6151
R958 B.n311 B.n310 10.6151
R959 B.n315 B.n314 10.6151
R960 B.n316 B.n315 10.6151
R961 B.n316 B.n142 10.6151
R962 B.n320 B.n142 10.6151
R963 B.n321 B.n320 10.6151
R964 B.n322 B.n321 10.6151
R965 B.n322 B.n140 10.6151
R966 B.n326 B.n140 10.6151
R967 B.n329 B.n328 10.6151
R968 B.n329 B.n136 10.6151
R969 B.n333 B.n136 10.6151
R970 B.n334 B.n333 10.6151
R971 B.n335 B.n334 10.6151
R972 B.n335 B.n134 10.6151
R973 B.n339 B.n134 10.6151
R974 B.n340 B.n339 10.6151
R975 B.n341 B.n340 10.6151
R976 B.n341 B.n132 10.6151
R977 B.n345 B.n132 10.6151
R978 B.n346 B.n345 10.6151
R979 B.n347 B.n346 10.6151
R980 B.n347 B.n130 10.6151
R981 B.n351 B.n130 10.6151
R982 B.n352 B.n351 10.6151
R983 B.n353 B.n352 10.6151
R984 B.n353 B.n128 10.6151
R985 B.n357 B.n128 10.6151
R986 B.n358 B.n357 10.6151
R987 B.n359 B.n358 10.6151
R988 B.n359 B.n126 10.6151
R989 B.n363 B.n126 10.6151
R990 B.n364 B.n363 10.6151
R991 B.n365 B.n364 10.6151
R992 B.n365 B.n124 10.6151
R993 B.n369 B.n124 10.6151
R994 B.n370 B.n369 10.6151
R995 B.n371 B.n370 10.6151
R996 B.n371 B.n122 10.6151
R997 B.n375 B.n122 10.6151
R998 B.n376 B.n375 10.6151
R999 B.n377 B.n376 10.6151
R1000 B.n377 B.n120 10.6151
R1001 B.n381 B.n120 10.6151
R1002 B.n382 B.n381 10.6151
R1003 B.n383 B.n382 10.6151
R1004 B.n383 B.n118 10.6151
R1005 B.n387 B.n118 10.6151
R1006 B.n388 B.n387 10.6151
R1007 B.n389 B.n388 10.6151
R1008 B.n389 B.n116 10.6151
R1009 B.n393 B.n116 10.6151
R1010 B.n394 B.n393 10.6151
R1011 B.n395 B.n394 10.6151
R1012 B.n395 B.n114 10.6151
R1013 B.n399 B.n114 10.6151
R1014 B.n400 B.n399 10.6151
R1015 B.n238 B.n237 10.6151
R1016 B.n237 B.n172 10.6151
R1017 B.n233 B.n172 10.6151
R1018 B.n233 B.n232 10.6151
R1019 B.n232 B.n231 10.6151
R1020 B.n231 B.n174 10.6151
R1021 B.n227 B.n174 10.6151
R1022 B.n227 B.n226 10.6151
R1023 B.n226 B.n225 10.6151
R1024 B.n225 B.n176 10.6151
R1025 B.n221 B.n176 10.6151
R1026 B.n221 B.n220 10.6151
R1027 B.n220 B.n219 10.6151
R1028 B.n219 B.n178 10.6151
R1029 B.n215 B.n178 10.6151
R1030 B.n215 B.n214 10.6151
R1031 B.n214 B.n213 10.6151
R1032 B.n213 B.n180 10.6151
R1033 B.n209 B.n180 10.6151
R1034 B.n209 B.n208 10.6151
R1035 B.n208 B.n207 10.6151
R1036 B.n207 B.n182 10.6151
R1037 B.n203 B.n182 10.6151
R1038 B.n203 B.n202 10.6151
R1039 B.n202 B.n201 10.6151
R1040 B.n201 B.n184 10.6151
R1041 B.n197 B.n184 10.6151
R1042 B.n197 B.n196 10.6151
R1043 B.n196 B.n195 10.6151
R1044 B.n195 B.n186 10.6151
R1045 B.n191 B.n186 10.6151
R1046 B.n191 B.n190 10.6151
R1047 B.n190 B.n189 10.6151
R1048 B.n189 B.n0 10.6151
R1049 B.n719 B.n1 10.6151
R1050 B.n719 B.n718 10.6151
R1051 B.n718 B.n717 10.6151
R1052 B.n717 B.n4 10.6151
R1053 B.n713 B.n4 10.6151
R1054 B.n713 B.n712 10.6151
R1055 B.n712 B.n711 10.6151
R1056 B.n711 B.n6 10.6151
R1057 B.n707 B.n6 10.6151
R1058 B.n707 B.n706 10.6151
R1059 B.n706 B.n705 10.6151
R1060 B.n705 B.n8 10.6151
R1061 B.n701 B.n8 10.6151
R1062 B.n701 B.n700 10.6151
R1063 B.n700 B.n699 10.6151
R1064 B.n699 B.n10 10.6151
R1065 B.n695 B.n10 10.6151
R1066 B.n695 B.n694 10.6151
R1067 B.n694 B.n693 10.6151
R1068 B.n693 B.n12 10.6151
R1069 B.n689 B.n12 10.6151
R1070 B.n689 B.n688 10.6151
R1071 B.n688 B.n687 10.6151
R1072 B.n687 B.n14 10.6151
R1073 B.n683 B.n14 10.6151
R1074 B.n683 B.n682 10.6151
R1075 B.n682 B.n681 10.6151
R1076 B.n681 B.n16 10.6151
R1077 B.n677 B.n16 10.6151
R1078 B.n677 B.n676 10.6151
R1079 B.n676 B.n675 10.6151
R1080 B.n675 B.n18 10.6151
R1081 B.n671 B.n18 10.6151
R1082 B.n671 B.n670 10.6151
R1083 B.n594 B.n46 6.5566
R1084 B.n582 B.n581 6.5566
R1085 B.n314 B.n146 6.5566
R1086 B.n327 B.n326 6.5566
R1087 B.n597 B.n46 4.05904
R1088 B.n581 B.n580 4.05904
R1089 B.n311 B.n146 4.05904
R1090 B.n328 B.n327 4.05904
R1091 B.n723 B.n0 2.81026
R1092 B.n723 B.n1 2.81026
R1093 VP.n4 VP.t2 161.726
R1094 VP.n16 VP.n0 161.3
R1095 VP.n15 VP.n14 161.3
R1096 VP.n13 VP.n1 161.3
R1097 VP.n12 VP.n11 161.3
R1098 VP.n10 VP.n2 161.3
R1099 VP.n9 VP.n8 161.3
R1100 VP.n7 VP.n3 161.3
R1101 VP.n4 VP.t1 160.853
R1102 VP.n5 VP.t0 127.588
R1103 VP.n17 VP.t3 127.588
R1104 VP.n6 VP.n5 109.389
R1105 VP.n18 VP.n17 109.389
R1106 VP.n6 VP.n4 52.0497
R1107 VP.n11 VP.n10 40.4106
R1108 VP.n11 VP.n1 40.4106
R1109 VP.n9 VP.n3 24.3439
R1110 VP.n10 VP.n9 24.3439
R1111 VP.n15 VP.n1 24.3439
R1112 VP.n16 VP.n15 24.3439
R1113 VP.n5 VP.n3 1.21767
R1114 VP.n17 VP.n16 1.21767
R1115 VP.n7 VP.n6 0.278398
R1116 VP.n18 VP.n0 0.278398
R1117 VP.n8 VP.n7 0.189894
R1118 VP.n8 VP.n2 0.189894
R1119 VP.n12 VP.n2 0.189894
R1120 VP.n13 VP.n12 0.189894
R1121 VP.n14 VP.n13 0.189894
R1122 VP.n14 VP.n0 0.189894
R1123 VP VP.n18 0.153422
R1124 VDD1 VDD1.n1 117.91
R1125 VDD1 VDD1.n0 73.4279
R1126 VDD1.n0 VDD1.t3 2.25779
R1127 VDD1.n0 VDD1.t0 2.25779
R1128 VDD1.n1 VDD1.t1 2.25779
R1129 VDD1.n1 VDD1.t2 2.25779
R1130 VTAIL.n5 VTAIL.t5 58.9483
R1131 VTAIL.n4 VTAIL.t1 58.9483
R1132 VTAIL.n3 VTAIL.t0 58.9483
R1133 VTAIL.n7 VTAIL.t3 58.9482
R1134 VTAIL.n0 VTAIL.t2 58.9482
R1135 VTAIL.n1 VTAIL.t4 58.9482
R1136 VTAIL.n2 VTAIL.t7 58.9482
R1137 VTAIL.n6 VTAIL.t6 58.9482
R1138 VTAIL.n7 VTAIL.n6 27.41
R1139 VTAIL.n3 VTAIL.n2 27.41
R1140 VTAIL.n4 VTAIL.n3 2.62981
R1141 VTAIL.n6 VTAIL.n5 2.62981
R1142 VTAIL.n2 VTAIL.n1 2.62981
R1143 VTAIL VTAIL.n0 1.37334
R1144 VTAIL VTAIL.n7 1.25697
R1145 VTAIL.n5 VTAIL.n4 0.470328
R1146 VTAIL.n1 VTAIL.n0 0.470328
R1147 VN.n0 VN.t2 161.726
R1148 VN.n1 VN.t1 161.726
R1149 VN.n0 VN.t3 160.853
R1150 VN.n1 VN.t0 160.853
R1151 VN VN.n1 52.3286
R1152 VN VN.n0 3.63537
R1153 VDD2.n2 VDD2.n0 117.386
R1154 VDD2.n2 VDD2.n1 73.3697
R1155 VDD2.n1 VDD2.t3 2.25779
R1156 VDD2.n1 VDD2.t2 2.25779
R1157 VDD2.n0 VDD2.t1 2.25779
R1158 VDD2.n0 VDD2.t0 2.25779
R1159 VDD2 VDD2.n2 0.0586897
C0 VDD2 VDD1 1.04914f
C1 w_n2800_n3848# VDD2 1.59687f
C2 VP VDD2 0.401443f
C3 B VTAIL 5.79306f
C4 VTAIL VDD1 5.98952f
C5 VTAIL w_n2800_n3848# 4.51503f
C6 B VDD1 1.34681f
C7 VN VDD2 5.68683f
C8 VTAIL VP 5.51438f
C9 B w_n2800_n3848# 10.0666f
C10 B VP 1.75413f
C11 w_n2800_n3848# VDD1 1.53809f
C12 VP VDD1 5.9389f
C13 VTAIL VN 5.50027f
C14 VP w_n2800_n3848# 5.18351f
C15 B VN 1.15574f
C16 VTAIL VDD2 6.044529f
C17 B VDD2 1.40094f
C18 VN VDD1 0.14861f
C19 VN w_n2800_n3848# 4.82325f
C20 VP VN 6.7287f
C21 VDD2 VSUBS 1.028135f
C22 VDD1 VSUBS 6.09226f
C23 VTAIL VSUBS 1.340264f
C24 VN VSUBS 5.58196f
C25 VP VSUBS 2.425517f
C26 B VSUBS 4.583f
C27 w_n2800_n3848# VSUBS 0.132216p
C28 VDD2.t1 VSUBS 0.303154f
C29 VDD2.t0 VSUBS 0.303154f
C30 VDD2.n0 VSUBS 3.24503f
C31 VDD2.t3 VSUBS 0.303154f
C32 VDD2.t2 VSUBS 0.303154f
C33 VDD2.n1 VSUBS 2.45462f
C34 VDD2.n2 VSUBS 4.55629f
C35 VN.t2 VSUBS 3.56307f
C36 VN.t3 VSUBS 3.55589f
C37 VN.n0 VSUBS 2.28552f
C38 VN.t1 VSUBS 3.56307f
C39 VN.t0 VSUBS 3.55589f
C40 VN.n1 VSUBS 4.08543f
C41 VTAIL.t2 VSUBS 2.61742f
C42 VTAIL.n0 VSUBS 0.754745f
C43 VTAIL.t4 VSUBS 2.61742f
C44 VTAIL.n1 VSUBS 0.847979f
C45 VTAIL.t7 VSUBS 2.61742f
C46 VTAIL.n2 VSUBS 2.24218f
C47 VTAIL.t0 VSUBS 2.61744f
C48 VTAIL.n3 VSUBS 2.24216f
C49 VTAIL.t1 VSUBS 2.61744f
C50 VTAIL.n4 VSUBS 0.847959f
C51 VTAIL.t5 VSUBS 2.61744f
C52 VTAIL.n5 VSUBS 0.847959f
C53 VTAIL.t6 VSUBS 2.61742f
C54 VTAIL.n6 VSUBS 2.24218f
C55 VTAIL.t3 VSUBS 2.61742f
C56 VTAIL.n7 VSUBS 2.14032f
C57 VDD1.t3 VSUBS 0.305764f
C58 VDD1.t0 VSUBS 0.305764f
C59 VDD1.n0 VSUBS 2.47635f
C60 VDD1.t1 VSUBS 0.305764f
C61 VDD1.t2 VSUBS 0.305764f
C62 VDD1.n1 VSUBS 3.29897f
C63 VP.n0 VSUBS 0.041442f
C64 VP.t3 VSUBS 3.37026f
C65 VP.n1 VSUBS 0.062803f
C66 VP.n2 VSUBS 0.031431f
C67 VP.n3 VSUBS 0.031259f
C68 VP.t1 VSUBS 3.6568f
C69 VP.t2 VSUBS 3.66418f
C70 VP.n4 VSUBS 4.18482f
C71 VP.t0 VSUBS 3.37026f
C72 VP.n5 VSUBS 1.27548f
C73 VP.n6 VSUBS 1.83766f
C74 VP.n7 VSUBS 0.041442f
C75 VP.n8 VSUBS 0.031431f
C76 VP.n9 VSUBS 0.058874f
C77 VP.n10 VSUBS 0.062803f
C78 VP.n11 VSUBS 0.025435f
C79 VP.n12 VSUBS 0.031431f
C80 VP.n13 VSUBS 0.031431f
C81 VP.n14 VSUBS 0.031431f
C82 VP.n15 VSUBS 0.058874f
C83 VP.n16 VSUBS 0.031259f
C84 VP.n17 VSUBS 1.27548f
C85 VP.n18 VSUBS 0.058674f
C86 B.n0 VSUBS 0.004011f
C87 B.n1 VSUBS 0.004011f
C88 B.n2 VSUBS 0.006343f
C89 B.n3 VSUBS 0.006343f
C90 B.n4 VSUBS 0.006343f
C91 B.n5 VSUBS 0.006343f
C92 B.n6 VSUBS 0.006343f
C93 B.n7 VSUBS 0.006343f
C94 B.n8 VSUBS 0.006343f
C95 B.n9 VSUBS 0.006343f
C96 B.n10 VSUBS 0.006343f
C97 B.n11 VSUBS 0.006343f
C98 B.n12 VSUBS 0.006343f
C99 B.n13 VSUBS 0.006343f
C100 B.n14 VSUBS 0.006343f
C101 B.n15 VSUBS 0.006343f
C102 B.n16 VSUBS 0.006343f
C103 B.n17 VSUBS 0.006343f
C104 B.n18 VSUBS 0.006343f
C105 B.n19 VSUBS 0.014341f
C106 B.n20 VSUBS 0.006343f
C107 B.n21 VSUBS 0.006343f
C108 B.n22 VSUBS 0.006343f
C109 B.n23 VSUBS 0.006343f
C110 B.n24 VSUBS 0.006343f
C111 B.n25 VSUBS 0.006343f
C112 B.n26 VSUBS 0.006343f
C113 B.n27 VSUBS 0.006343f
C114 B.n28 VSUBS 0.006343f
C115 B.n29 VSUBS 0.006343f
C116 B.n30 VSUBS 0.006343f
C117 B.n31 VSUBS 0.006343f
C118 B.n32 VSUBS 0.006343f
C119 B.n33 VSUBS 0.006343f
C120 B.n34 VSUBS 0.006343f
C121 B.n35 VSUBS 0.006343f
C122 B.n36 VSUBS 0.006343f
C123 B.n37 VSUBS 0.006343f
C124 B.n38 VSUBS 0.006343f
C125 B.n39 VSUBS 0.006343f
C126 B.n40 VSUBS 0.006343f
C127 B.n41 VSUBS 0.006343f
C128 B.n42 VSUBS 0.006343f
C129 B.n43 VSUBS 0.006343f
C130 B.t8 VSUBS 0.432844f
C131 B.t7 VSUBS 0.452759f
C132 B.t6 VSUBS 1.60306f
C133 B.n44 VSUBS 0.243696f
C134 B.n45 VSUBS 0.065647f
C135 B.n46 VSUBS 0.014696f
C136 B.n47 VSUBS 0.006343f
C137 B.n48 VSUBS 0.006343f
C138 B.n49 VSUBS 0.006343f
C139 B.n50 VSUBS 0.006343f
C140 B.n51 VSUBS 0.006343f
C141 B.t11 VSUBS 0.432832f
C142 B.t10 VSUBS 0.45275f
C143 B.t9 VSUBS 1.60306f
C144 B.n52 VSUBS 0.243705f
C145 B.n53 VSUBS 0.065658f
C146 B.n54 VSUBS 0.006343f
C147 B.n55 VSUBS 0.006343f
C148 B.n56 VSUBS 0.006343f
C149 B.n57 VSUBS 0.006343f
C150 B.n58 VSUBS 0.006343f
C151 B.n59 VSUBS 0.006343f
C152 B.n60 VSUBS 0.006343f
C153 B.n61 VSUBS 0.006343f
C154 B.n62 VSUBS 0.006343f
C155 B.n63 VSUBS 0.006343f
C156 B.n64 VSUBS 0.006343f
C157 B.n65 VSUBS 0.006343f
C158 B.n66 VSUBS 0.006343f
C159 B.n67 VSUBS 0.006343f
C160 B.n68 VSUBS 0.006343f
C161 B.n69 VSUBS 0.006343f
C162 B.n70 VSUBS 0.006343f
C163 B.n71 VSUBS 0.006343f
C164 B.n72 VSUBS 0.006343f
C165 B.n73 VSUBS 0.006343f
C166 B.n74 VSUBS 0.006343f
C167 B.n75 VSUBS 0.006343f
C168 B.n76 VSUBS 0.006343f
C169 B.n77 VSUBS 0.015135f
C170 B.n78 VSUBS 0.006343f
C171 B.n79 VSUBS 0.006343f
C172 B.n80 VSUBS 0.006343f
C173 B.n81 VSUBS 0.006343f
C174 B.n82 VSUBS 0.006343f
C175 B.n83 VSUBS 0.006343f
C176 B.n84 VSUBS 0.006343f
C177 B.n85 VSUBS 0.006343f
C178 B.n86 VSUBS 0.006343f
C179 B.n87 VSUBS 0.006343f
C180 B.n88 VSUBS 0.006343f
C181 B.n89 VSUBS 0.006343f
C182 B.n90 VSUBS 0.006343f
C183 B.n91 VSUBS 0.006343f
C184 B.n92 VSUBS 0.006343f
C185 B.n93 VSUBS 0.006343f
C186 B.n94 VSUBS 0.006343f
C187 B.n95 VSUBS 0.006343f
C188 B.n96 VSUBS 0.006343f
C189 B.n97 VSUBS 0.006343f
C190 B.n98 VSUBS 0.006343f
C191 B.n99 VSUBS 0.006343f
C192 B.n100 VSUBS 0.006343f
C193 B.n101 VSUBS 0.006343f
C194 B.n102 VSUBS 0.006343f
C195 B.n103 VSUBS 0.006343f
C196 B.n104 VSUBS 0.006343f
C197 B.n105 VSUBS 0.006343f
C198 B.n106 VSUBS 0.006343f
C199 B.n107 VSUBS 0.006343f
C200 B.n108 VSUBS 0.006343f
C201 B.n109 VSUBS 0.006343f
C202 B.n110 VSUBS 0.006343f
C203 B.n111 VSUBS 0.006343f
C204 B.n112 VSUBS 0.006343f
C205 B.n113 VSUBS 0.015135f
C206 B.n114 VSUBS 0.006343f
C207 B.n115 VSUBS 0.006343f
C208 B.n116 VSUBS 0.006343f
C209 B.n117 VSUBS 0.006343f
C210 B.n118 VSUBS 0.006343f
C211 B.n119 VSUBS 0.006343f
C212 B.n120 VSUBS 0.006343f
C213 B.n121 VSUBS 0.006343f
C214 B.n122 VSUBS 0.006343f
C215 B.n123 VSUBS 0.006343f
C216 B.n124 VSUBS 0.006343f
C217 B.n125 VSUBS 0.006343f
C218 B.n126 VSUBS 0.006343f
C219 B.n127 VSUBS 0.006343f
C220 B.n128 VSUBS 0.006343f
C221 B.n129 VSUBS 0.006343f
C222 B.n130 VSUBS 0.006343f
C223 B.n131 VSUBS 0.006343f
C224 B.n132 VSUBS 0.006343f
C225 B.n133 VSUBS 0.006343f
C226 B.n134 VSUBS 0.006343f
C227 B.n135 VSUBS 0.006343f
C228 B.n136 VSUBS 0.006343f
C229 B.n137 VSUBS 0.006343f
C230 B.t1 VSUBS 0.432832f
C231 B.t2 VSUBS 0.45275f
C232 B.t0 VSUBS 1.60306f
C233 B.n138 VSUBS 0.243705f
C234 B.n139 VSUBS 0.065658f
C235 B.n140 VSUBS 0.006343f
C236 B.n141 VSUBS 0.006343f
C237 B.n142 VSUBS 0.006343f
C238 B.n143 VSUBS 0.006343f
C239 B.t4 VSUBS 0.432844f
C240 B.t5 VSUBS 0.452759f
C241 B.t3 VSUBS 1.60306f
C242 B.n144 VSUBS 0.243696f
C243 B.n145 VSUBS 0.065647f
C244 B.n146 VSUBS 0.014696f
C245 B.n147 VSUBS 0.006343f
C246 B.n148 VSUBS 0.006343f
C247 B.n149 VSUBS 0.006343f
C248 B.n150 VSUBS 0.006343f
C249 B.n151 VSUBS 0.006343f
C250 B.n152 VSUBS 0.006343f
C251 B.n153 VSUBS 0.006343f
C252 B.n154 VSUBS 0.006343f
C253 B.n155 VSUBS 0.006343f
C254 B.n156 VSUBS 0.006343f
C255 B.n157 VSUBS 0.006343f
C256 B.n158 VSUBS 0.006343f
C257 B.n159 VSUBS 0.006343f
C258 B.n160 VSUBS 0.006343f
C259 B.n161 VSUBS 0.006343f
C260 B.n162 VSUBS 0.006343f
C261 B.n163 VSUBS 0.006343f
C262 B.n164 VSUBS 0.006343f
C263 B.n165 VSUBS 0.006343f
C264 B.n166 VSUBS 0.006343f
C265 B.n167 VSUBS 0.006343f
C266 B.n168 VSUBS 0.006343f
C267 B.n169 VSUBS 0.006343f
C268 B.n170 VSUBS 0.006343f
C269 B.n171 VSUBS 0.014341f
C270 B.n172 VSUBS 0.006343f
C271 B.n173 VSUBS 0.006343f
C272 B.n174 VSUBS 0.006343f
C273 B.n175 VSUBS 0.006343f
C274 B.n176 VSUBS 0.006343f
C275 B.n177 VSUBS 0.006343f
C276 B.n178 VSUBS 0.006343f
C277 B.n179 VSUBS 0.006343f
C278 B.n180 VSUBS 0.006343f
C279 B.n181 VSUBS 0.006343f
C280 B.n182 VSUBS 0.006343f
C281 B.n183 VSUBS 0.006343f
C282 B.n184 VSUBS 0.006343f
C283 B.n185 VSUBS 0.006343f
C284 B.n186 VSUBS 0.006343f
C285 B.n187 VSUBS 0.006343f
C286 B.n188 VSUBS 0.006343f
C287 B.n189 VSUBS 0.006343f
C288 B.n190 VSUBS 0.006343f
C289 B.n191 VSUBS 0.006343f
C290 B.n192 VSUBS 0.006343f
C291 B.n193 VSUBS 0.006343f
C292 B.n194 VSUBS 0.006343f
C293 B.n195 VSUBS 0.006343f
C294 B.n196 VSUBS 0.006343f
C295 B.n197 VSUBS 0.006343f
C296 B.n198 VSUBS 0.006343f
C297 B.n199 VSUBS 0.006343f
C298 B.n200 VSUBS 0.006343f
C299 B.n201 VSUBS 0.006343f
C300 B.n202 VSUBS 0.006343f
C301 B.n203 VSUBS 0.006343f
C302 B.n204 VSUBS 0.006343f
C303 B.n205 VSUBS 0.006343f
C304 B.n206 VSUBS 0.006343f
C305 B.n207 VSUBS 0.006343f
C306 B.n208 VSUBS 0.006343f
C307 B.n209 VSUBS 0.006343f
C308 B.n210 VSUBS 0.006343f
C309 B.n211 VSUBS 0.006343f
C310 B.n212 VSUBS 0.006343f
C311 B.n213 VSUBS 0.006343f
C312 B.n214 VSUBS 0.006343f
C313 B.n215 VSUBS 0.006343f
C314 B.n216 VSUBS 0.006343f
C315 B.n217 VSUBS 0.006343f
C316 B.n218 VSUBS 0.006343f
C317 B.n219 VSUBS 0.006343f
C318 B.n220 VSUBS 0.006343f
C319 B.n221 VSUBS 0.006343f
C320 B.n222 VSUBS 0.006343f
C321 B.n223 VSUBS 0.006343f
C322 B.n224 VSUBS 0.006343f
C323 B.n225 VSUBS 0.006343f
C324 B.n226 VSUBS 0.006343f
C325 B.n227 VSUBS 0.006343f
C326 B.n228 VSUBS 0.006343f
C327 B.n229 VSUBS 0.006343f
C328 B.n230 VSUBS 0.006343f
C329 B.n231 VSUBS 0.006343f
C330 B.n232 VSUBS 0.006343f
C331 B.n233 VSUBS 0.006343f
C332 B.n234 VSUBS 0.006343f
C333 B.n235 VSUBS 0.006343f
C334 B.n236 VSUBS 0.006343f
C335 B.n237 VSUBS 0.006343f
C336 B.n238 VSUBS 0.014341f
C337 B.n239 VSUBS 0.015135f
C338 B.n240 VSUBS 0.015135f
C339 B.n241 VSUBS 0.006343f
C340 B.n242 VSUBS 0.006343f
C341 B.n243 VSUBS 0.006343f
C342 B.n244 VSUBS 0.006343f
C343 B.n245 VSUBS 0.006343f
C344 B.n246 VSUBS 0.006343f
C345 B.n247 VSUBS 0.006343f
C346 B.n248 VSUBS 0.006343f
C347 B.n249 VSUBS 0.006343f
C348 B.n250 VSUBS 0.006343f
C349 B.n251 VSUBS 0.006343f
C350 B.n252 VSUBS 0.006343f
C351 B.n253 VSUBS 0.006343f
C352 B.n254 VSUBS 0.006343f
C353 B.n255 VSUBS 0.006343f
C354 B.n256 VSUBS 0.006343f
C355 B.n257 VSUBS 0.006343f
C356 B.n258 VSUBS 0.006343f
C357 B.n259 VSUBS 0.006343f
C358 B.n260 VSUBS 0.006343f
C359 B.n261 VSUBS 0.006343f
C360 B.n262 VSUBS 0.006343f
C361 B.n263 VSUBS 0.006343f
C362 B.n264 VSUBS 0.006343f
C363 B.n265 VSUBS 0.006343f
C364 B.n266 VSUBS 0.006343f
C365 B.n267 VSUBS 0.006343f
C366 B.n268 VSUBS 0.006343f
C367 B.n269 VSUBS 0.006343f
C368 B.n270 VSUBS 0.006343f
C369 B.n271 VSUBS 0.006343f
C370 B.n272 VSUBS 0.006343f
C371 B.n273 VSUBS 0.006343f
C372 B.n274 VSUBS 0.006343f
C373 B.n275 VSUBS 0.006343f
C374 B.n276 VSUBS 0.006343f
C375 B.n277 VSUBS 0.006343f
C376 B.n278 VSUBS 0.006343f
C377 B.n279 VSUBS 0.006343f
C378 B.n280 VSUBS 0.006343f
C379 B.n281 VSUBS 0.006343f
C380 B.n282 VSUBS 0.006343f
C381 B.n283 VSUBS 0.006343f
C382 B.n284 VSUBS 0.006343f
C383 B.n285 VSUBS 0.006343f
C384 B.n286 VSUBS 0.006343f
C385 B.n287 VSUBS 0.006343f
C386 B.n288 VSUBS 0.006343f
C387 B.n289 VSUBS 0.006343f
C388 B.n290 VSUBS 0.006343f
C389 B.n291 VSUBS 0.006343f
C390 B.n292 VSUBS 0.006343f
C391 B.n293 VSUBS 0.006343f
C392 B.n294 VSUBS 0.006343f
C393 B.n295 VSUBS 0.006343f
C394 B.n296 VSUBS 0.006343f
C395 B.n297 VSUBS 0.006343f
C396 B.n298 VSUBS 0.006343f
C397 B.n299 VSUBS 0.006343f
C398 B.n300 VSUBS 0.006343f
C399 B.n301 VSUBS 0.006343f
C400 B.n302 VSUBS 0.006343f
C401 B.n303 VSUBS 0.006343f
C402 B.n304 VSUBS 0.006343f
C403 B.n305 VSUBS 0.006343f
C404 B.n306 VSUBS 0.006343f
C405 B.n307 VSUBS 0.006343f
C406 B.n308 VSUBS 0.006343f
C407 B.n309 VSUBS 0.006343f
C408 B.n310 VSUBS 0.006343f
C409 B.n311 VSUBS 0.004384f
C410 B.n312 VSUBS 0.006343f
C411 B.n313 VSUBS 0.006343f
C412 B.n314 VSUBS 0.00513f
C413 B.n315 VSUBS 0.006343f
C414 B.n316 VSUBS 0.006343f
C415 B.n317 VSUBS 0.006343f
C416 B.n318 VSUBS 0.006343f
C417 B.n319 VSUBS 0.006343f
C418 B.n320 VSUBS 0.006343f
C419 B.n321 VSUBS 0.006343f
C420 B.n322 VSUBS 0.006343f
C421 B.n323 VSUBS 0.006343f
C422 B.n324 VSUBS 0.006343f
C423 B.n325 VSUBS 0.006343f
C424 B.n326 VSUBS 0.00513f
C425 B.n327 VSUBS 0.014696f
C426 B.n328 VSUBS 0.004384f
C427 B.n329 VSUBS 0.006343f
C428 B.n330 VSUBS 0.006343f
C429 B.n331 VSUBS 0.006343f
C430 B.n332 VSUBS 0.006343f
C431 B.n333 VSUBS 0.006343f
C432 B.n334 VSUBS 0.006343f
C433 B.n335 VSUBS 0.006343f
C434 B.n336 VSUBS 0.006343f
C435 B.n337 VSUBS 0.006343f
C436 B.n338 VSUBS 0.006343f
C437 B.n339 VSUBS 0.006343f
C438 B.n340 VSUBS 0.006343f
C439 B.n341 VSUBS 0.006343f
C440 B.n342 VSUBS 0.006343f
C441 B.n343 VSUBS 0.006343f
C442 B.n344 VSUBS 0.006343f
C443 B.n345 VSUBS 0.006343f
C444 B.n346 VSUBS 0.006343f
C445 B.n347 VSUBS 0.006343f
C446 B.n348 VSUBS 0.006343f
C447 B.n349 VSUBS 0.006343f
C448 B.n350 VSUBS 0.006343f
C449 B.n351 VSUBS 0.006343f
C450 B.n352 VSUBS 0.006343f
C451 B.n353 VSUBS 0.006343f
C452 B.n354 VSUBS 0.006343f
C453 B.n355 VSUBS 0.006343f
C454 B.n356 VSUBS 0.006343f
C455 B.n357 VSUBS 0.006343f
C456 B.n358 VSUBS 0.006343f
C457 B.n359 VSUBS 0.006343f
C458 B.n360 VSUBS 0.006343f
C459 B.n361 VSUBS 0.006343f
C460 B.n362 VSUBS 0.006343f
C461 B.n363 VSUBS 0.006343f
C462 B.n364 VSUBS 0.006343f
C463 B.n365 VSUBS 0.006343f
C464 B.n366 VSUBS 0.006343f
C465 B.n367 VSUBS 0.006343f
C466 B.n368 VSUBS 0.006343f
C467 B.n369 VSUBS 0.006343f
C468 B.n370 VSUBS 0.006343f
C469 B.n371 VSUBS 0.006343f
C470 B.n372 VSUBS 0.006343f
C471 B.n373 VSUBS 0.006343f
C472 B.n374 VSUBS 0.006343f
C473 B.n375 VSUBS 0.006343f
C474 B.n376 VSUBS 0.006343f
C475 B.n377 VSUBS 0.006343f
C476 B.n378 VSUBS 0.006343f
C477 B.n379 VSUBS 0.006343f
C478 B.n380 VSUBS 0.006343f
C479 B.n381 VSUBS 0.006343f
C480 B.n382 VSUBS 0.006343f
C481 B.n383 VSUBS 0.006343f
C482 B.n384 VSUBS 0.006343f
C483 B.n385 VSUBS 0.006343f
C484 B.n386 VSUBS 0.006343f
C485 B.n387 VSUBS 0.006343f
C486 B.n388 VSUBS 0.006343f
C487 B.n389 VSUBS 0.006343f
C488 B.n390 VSUBS 0.006343f
C489 B.n391 VSUBS 0.006343f
C490 B.n392 VSUBS 0.006343f
C491 B.n393 VSUBS 0.006343f
C492 B.n394 VSUBS 0.006343f
C493 B.n395 VSUBS 0.006343f
C494 B.n396 VSUBS 0.006343f
C495 B.n397 VSUBS 0.006343f
C496 B.n398 VSUBS 0.006343f
C497 B.n399 VSUBS 0.006343f
C498 B.n400 VSUBS 0.015135f
C499 B.n401 VSUBS 0.014341f
C500 B.n402 VSUBS 0.014341f
C501 B.n403 VSUBS 0.006343f
C502 B.n404 VSUBS 0.006343f
C503 B.n405 VSUBS 0.006343f
C504 B.n406 VSUBS 0.006343f
C505 B.n407 VSUBS 0.006343f
C506 B.n408 VSUBS 0.006343f
C507 B.n409 VSUBS 0.006343f
C508 B.n410 VSUBS 0.006343f
C509 B.n411 VSUBS 0.006343f
C510 B.n412 VSUBS 0.006343f
C511 B.n413 VSUBS 0.006343f
C512 B.n414 VSUBS 0.006343f
C513 B.n415 VSUBS 0.006343f
C514 B.n416 VSUBS 0.006343f
C515 B.n417 VSUBS 0.006343f
C516 B.n418 VSUBS 0.006343f
C517 B.n419 VSUBS 0.006343f
C518 B.n420 VSUBS 0.006343f
C519 B.n421 VSUBS 0.006343f
C520 B.n422 VSUBS 0.006343f
C521 B.n423 VSUBS 0.006343f
C522 B.n424 VSUBS 0.006343f
C523 B.n425 VSUBS 0.006343f
C524 B.n426 VSUBS 0.006343f
C525 B.n427 VSUBS 0.006343f
C526 B.n428 VSUBS 0.006343f
C527 B.n429 VSUBS 0.006343f
C528 B.n430 VSUBS 0.006343f
C529 B.n431 VSUBS 0.006343f
C530 B.n432 VSUBS 0.006343f
C531 B.n433 VSUBS 0.006343f
C532 B.n434 VSUBS 0.006343f
C533 B.n435 VSUBS 0.006343f
C534 B.n436 VSUBS 0.006343f
C535 B.n437 VSUBS 0.006343f
C536 B.n438 VSUBS 0.006343f
C537 B.n439 VSUBS 0.006343f
C538 B.n440 VSUBS 0.006343f
C539 B.n441 VSUBS 0.006343f
C540 B.n442 VSUBS 0.006343f
C541 B.n443 VSUBS 0.006343f
C542 B.n444 VSUBS 0.006343f
C543 B.n445 VSUBS 0.006343f
C544 B.n446 VSUBS 0.006343f
C545 B.n447 VSUBS 0.006343f
C546 B.n448 VSUBS 0.006343f
C547 B.n449 VSUBS 0.006343f
C548 B.n450 VSUBS 0.006343f
C549 B.n451 VSUBS 0.006343f
C550 B.n452 VSUBS 0.006343f
C551 B.n453 VSUBS 0.006343f
C552 B.n454 VSUBS 0.006343f
C553 B.n455 VSUBS 0.006343f
C554 B.n456 VSUBS 0.006343f
C555 B.n457 VSUBS 0.006343f
C556 B.n458 VSUBS 0.006343f
C557 B.n459 VSUBS 0.006343f
C558 B.n460 VSUBS 0.006343f
C559 B.n461 VSUBS 0.006343f
C560 B.n462 VSUBS 0.006343f
C561 B.n463 VSUBS 0.006343f
C562 B.n464 VSUBS 0.006343f
C563 B.n465 VSUBS 0.006343f
C564 B.n466 VSUBS 0.006343f
C565 B.n467 VSUBS 0.006343f
C566 B.n468 VSUBS 0.006343f
C567 B.n469 VSUBS 0.006343f
C568 B.n470 VSUBS 0.006343f
C569 B.n471 VSUBS 0.006343f
C570 B.n472 VSUBS 0.006343f
C571 B.n473 VSUBS 0.006343f
C572 B.n474 VSUBS 0.006343f
C573 B.n475 VSUBS 0.006343f
C574 B.n476 VSUBS 0.006343f
C575 B.n477 VSUBS 0.006343f
C576 B.n478 VSUBS 0.006343f
C577 B.n479 VSUBS 0.006343f
C578 B.n480 VSUBS 0.006343f
C579 B.n481 VSUBS 0.006343f
C580 B.n482 VSUBS 0.006343f
C581 B.n483 VSUBS 0.006343f
C582 B.n484 VSUBS 0.006343f
C583 B.n485 VSUBS 0.006343f
C584 B.n486 VSUBS 0.006343f
C585 B.n487 VSUBS 0.006343f
C586 B.n488 VSUBS 0.006343f
C587 B.n489 VSUBS 0.006343f
C588 B.n490 VSUBS 0.006343f
C589 B.n491 VSUBS 0.006343f
C590 B.n492 VSUBS 0.006343f
C591 B.n493 VSUBS 0.006343f
C592 B.n494 VSUBS 0.006343f
C593 B.n495 VSUBS 0.006343f
C594 B.n496 VSUBS 0.006343f
C595 B.n497 VSUBS 0.006343f
C596 B.n498 VSUBS 0.006343f
C597 B.n499 VSUBS 0.006343f
C598 B.n500 VSUBS 0.006343f
C599 B.n501 VSUBS 0.006343f
C600 B.n502 VSUBS 0.006343f
C601 B.n503 VSUBS 0.006343f
C602 B.n504 VSUBS 0.006343f
C603 B.n505 VSUBS 0.006343f
C604 B.n506 VSUBS 0.014341f
C605 B.n507 VSUBS 0.015098f
C606 B.n508 VSUBS 0.014378f
C607 B.n509 VSUBS 0.006343f
C608 B.n510 VSUBS 0.006343f
C609 B.n511 VSUBS 0.006343f
C610 B.n512 VSUBS 0.006343f
C611 B.n513 VSUBS 0.006343f
C612 B.n514 VSUBS 0.006343f
C613 B.n515 VSUBS 0.006343f
C614 B.n516 VSUBS 0.006343f
C615 B.n517 VSUBS 0.006343f
C616 B.n518 VSUBS 0.006343f
C617 B.n519 VSUBS 0.006343f
C618 B.n520 VSUBS 0.006343f
C619 B.n521 VSUBS 0.006343f
C620 B.n522 VSUBS 0.006343f
C621 B.n523 VSUBS 0.006343f
C622 B.n524 VSUBS 0.006343f
C623 B.n525 VSUBS 0.006343f
C624 B.n526 VSUBS 0.006343f
C625 B.n527 VSUBS 0.006343f
C626 B.n528 VSUBS 0.006343f
C627 B.n529 VSUBS 0.006343f
C628 B.n530 VSUBS 0.006343f
C629 B.n531 VSUBS 0.006343f
C630 B.n532 VSUBS 0.006343f
C631 B.n533 VSUBS 0.006343f
C632 B.n534 VSUBS 0.006343f
C633 B.n535 VSUBS 0.006343f
C634 B.n536 VSUBS 0.006343f
C635 B.n537 VSUBS 0.006343f
C636 B.n538 VSUBS 0.006343f
C637 B.n539 VSUBS 0.006343f
C638 B.n540 VSUBS 0.006343f
C639 B.n541 VSUBS 0.006343f
C640 B.n542 VSUBS 0.006343f
C641 B.n543 VSUBS 0.006343f
C642 B.n544 VSUBS 0.006343f
C643 B.n545 VSUBS 0.006343f
C644 B.n546 VSUBS 0.006343f
C645 B.n547 VSUBS 0.006343f
C646 B.n548 VSUBS 0.006343f
C647 B.n549 VSUBS 0.006343f
C648 B.n550 VSUBS 0.006343f
C649 B.n551 VSUBS 0.006343f
C650 B.n552 VSUBS 0.006343f
C651 B.n553 VSUBS 0.006343f
C652 B.n554 VSUBS 0.006343f
C653 B.n555 VSUBS 0.006343f
C654 B.n556 VSUBS 0.006343f
C655 B.n557 VSUBS 0.006343f
C656 B.n558 VSUBS 0.006343f
C657 B.n559 VSUBS 0.006343f
C658 B.n560 VSUBS 0.006343f
C659 B.n561 VSUBS 0.006343f
C660 B.n562 VSUBS 0.006343f
C661 B.n563 VSUBS 0.006343f
C662 B.n564 VSUBS 0.006343f
C663 B.n565 VSUBS 0.006343f
C664 B.n566 VSUBS 0.006343f
C665 B.n567 VSUBS 0.006343f
C666 B.n568 VSUBS 0.006343f
C667 B.n569 VSUBS 0.006343f
C668 B.n570 VSUBS 0.006343f
C669 B.n571 VSUBS 0.006343f
C670 B.n572 VSUBS 0.006343f
C671 B.n573 VSUBS 0.006343f
C672 B.n574 VSUBS 0.006343f
C673 B.n575 VSUBS 0.006343f
C674 B.n576 VSUBS 0.006343f
C675 B.n577 VSUBS 0.006343f
C676 B.n578 VSUBS 0.006343f
C677 B.n579 VSUBS 0.006343f
C678 B.n580 VSUBS 0.004384f
C679 B.n581 VSUBS 0.014696f
C680 B.n582 VSUBS 0.00513f
C681 B.n583 VSUBS 0.006343f
C682 B.n584 VSUBS 0.006343f
C683 B.n585 VSUBS 0.006343f
C684 B.n586 VSUBS 0.006343f
C685 B.n587 VSUBS 0.006343f
C686 B.n588 VSUBS 0.006343f
C687 B.n589 VSUBS 0.006343f
C688 B.n590 VSUBS 0.006343f
C689 B.n591 VSUBS 0.006343f
C690 B.n592 VSUBS 0.006343f
C691 B.n593 VSUBS 0.006343f
C692 B.n594 VSUBS 0.00513f
C693 B.n595 VSUBS 0.006343f
C694 B.n596 VSUBS 0.006343f
C695 B.n597 VSUBS 0.004384f
C696 B.n598 VSUBS 0.006343f
C697 B.n599 VSUBS 0.006343f
C698 B.n600 VSUBS 0.006343f
C699 B.n601 VSUBS 0.006343f
C700 B.n602 VSUBS 0.006343f
C701 B.n603 VSUBS 0.006343f
C702 B.n604 VSUBS 0.006343f
C703 B.n605 VSUBS 0.006343f
C704 B.n606 VSUBS 0.006343f
C705 B.n607 VSUBS 0.006343f
C706 B.n608 VSUBS 0.006343f
C707 B.n609 VSUBS 0.006343f
C708 B.n610 VSUBS 0.006343f
C709 B.n611 VSUBS 0.006343f
C710 B.n612 VSUBS 0.006343f
C711 B.n613 VSUBS 0.006343f
C712 B.n614 VSUBS 0.006343f
C713 B.n615 VSUBS 0.006343f
C714 B.n616 VSUBS 0.006343f
C715 B.n617 VSUBS 0.006343f
C716 B.n618 VSUBS 0.006343f
C717 B.n619 VSUBS 0.006343f
C718 B.n620 VSUBS 0.006343f
C719 B.n621 VSUBS 0.006343f
C720 B.n622 VSUBS 0.006343f
C721 B.n623 VSUBS 0.006343f
C722 B.n624 VSUBS 0.006343f
C723 B.n625 VSUBS 0.006343f
C724 B.n626 VSUBS 0.006343f
C725 B.n627 VSUBS 0.006343f
C726 B.n628 VSUBS 0.006343f
C727 B.n629 VSUBS 0.006343f
C728 B.n630 VSUBS 0.006343f
C729 B.n631 VSUBS 0.006343f
C730 B.n632 VSUBS 0.006343f
C731 B.n633 VSUBS 0.006343f
C732 B.n634 VSUBS 0.006343f
C733 B.n635 VSUBS 0.006343f
C734 B.n636 VSUBS 0.006343f
C735 B.n637 VSUBS 0.006343f
C736 B.n638 VSUBS 0.006343f
C737 B.n639 VSUBS 0.006343f
C738 B.n640 VSUBS 0.006343f
C739 B.n641 VSUBS 0.006343f
C740 B.n642 VSUBS 0.006343f
C741 B.n643 VSUBS 0.006343f
C742 B.n644 VSUBS 0.006343f
C743 B.n645 VSUBS 0.006343f
C744 B.n646 VSUBS 0.006343f
C745 B.n647 VSUBS 0.006343f
C746 B.n648 VSUBS 0.006343f
C747 B.n649 VSUBS 0.006343f
C748 B.n650 VSUBS 0.006343f
C749 B.n651 VSUBS 0.006343f
C750 B.n652 VSUBS 0.006343f
C751 B.n653 VSUBS 0.006343f
C752 B.n654 VSUBS 0.006343f
C753 B.n655 VSUBS 0.006343f
C754 B.n656 VSUBS 0.006343f
C755 B.n657 VSUBS 0.006343f
C756 B.n658 VSUBS 0.006343f
C757 B.n659 VSUBS 0.006343f
C758 B.n660 VSUBS 0.006343f
C759 B.n661 VSUBS 0.006343f
C760 B.n662 VSUBS 0.006343f
C761 B.n663 VSUBS 0.006343f
C762 B.n664 VSUBS 0.006343f
C763 B.n665 VSUBS 0.006343f
C764 B.n666 VSUBS 0.006343f
C765 B.n667 VSUBS 0.006343f
C766 B.n668 VSUBS 0.015135f
C767 B.n669 VSUBS 0.015135f
C768 B.n670 VSUBS 0.014341f
C769 B.n671 VSUBS 0.006343f
C770 B.n672 VSUBS 0.006343f
C771 B.n673 VSUBS 0.006343f
C772 B.n674 VSUBS 0.006343f
C773 B.n675 VSUBS 0.006343f
C774 B.n676 VSUBS 0.006343f
C775 B.n677 VSUBS 0.006343f
C776 B.n678 VSUBS 0.006343f
C777 B.n679 VSUBS 0.006343f
C778 B.n680 VSUBS 0.006343f
C779 B.n681 VSUBS 0.006343f
C780 B.n682 VSUBS 0.006343f
C781 B.n683 VSUBS 0.006343f
C782 B.n684 VSUBS 0.006343f
C783 B.n685 VSUBS 0.006343f
C784 B.n686 VSUBS 0.006343f
C785 B.n687 VSUBS 0.006343f
C786 B.n688 VSUBS 0.006343f
C787 B.n689 VSUBS 0.006343f
C788 B.n690 VSUBS 0.006343f
C789 B.n691 VSUBS 0.006343f
C790 B.n692 VSUBS 0.006343f
C791 B.n693 VSUBS 0.006343f
C792 B.n694 VSUBS 0.006343f
C793 B.n695 VSUBS 0.006343f
C794 B.n696 VSUBS 0.006343f
C795 B.n697 VSUBS 0.006343f
C796 B.n698 VSUBS 0.006343f
C797 B.n699 VSUBS 0.006343f
C798 B.n700 VSUBS 0.006343f
C799 B.n701 VSUBS 0.006343f
C800 B.n702 VSUBS 0.006343f
C801 B.n703 VSUBS 0.006343f
C802 B.n704 VSUBS 0.006343f
C803 B.n705 VSUBS 0.006343f
C804 B.n706 VSUBS 0.006343f
C805 B.n707 VSUBS 0.006343f
C806 B.n708 VSUBS 0.006343f
C807 B.n709 VSUBS 0.006343f
C808 B.n710 VSUBS 0.006343f
C809 B.n711 VSUBS 0.006343f
C810 B.n712 VSUBS 0.006343f
C811 B.n713 VSUBS 0.006343f
C812 B.n714 VSUBS 0.006343f
C813 B.n715 VSUBS 0.006343f
C814 B.n716 VSUBS 0.006343f
C815 B.n717 VSUBS 0.006343f
C816 B.n718 VSUBS 0.006343f
C817 B.n719 VSUBS 0.006343f
C818 B.n720 VSUBS 0.006343f
C819 B.n721 VSUBS 0.006343f
C820 B.n722 VSUBS 0.006343f
C821 B.n723 VSUBS 0.014363f
.ends

