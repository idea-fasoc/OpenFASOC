* NGSPICE file created from tg_sample_0002.ext - technology: sky130A

.subckt tg_sample_0002 VIN VGN VGP VSS VCC VOUT
X0 VOUT.t9 VGP.t0 VIN.t9 VCC.t4 sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=3.276 ps=17.58 w=8.4 l=3.34
X1 VOUT.t8 VGP.t1 VIN.t5 VCC.t3 sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=1.386 ps=8.73 w=8.4 l=3.34
X2 VIN.t1 VGN.t0 VOUT.t1 VSS.t4 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=3.47
X3 VCC.t12 VCC.t9 VCC.t11 VCC.t10 sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=0 ps=0 w=8.4 l=3.34
X4 VOUT.t7 VGP.t2 VIN.t6 VCC.t2 sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=1.386 ps=8.73 w=8.4 l=3.34
X5 VCC.t8 VCC.t5 VCC.t7 VCC.t6 sky130_fd_pr__pfet_01v8 ad=3.276 pd=17.58 as=0 ps=0 w=8.4 l=3.34
X6 VSS.t12 VSS.t9 VSS.t11 VSS.t10 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0 ps=0 w=0.98 l=3.47
X7 VIN.t3 VGN.t1 VOUT.t3 VSS.t3 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=3.47
X8 VOUT.t0 VGN.t2 VIN.t0 VSS.t2 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.3822 ps=2.74 w=0.98 l=3.47
X9 VOUT.t2 VGN.t3 VIN.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.1617 pd=1.31 as=0.1617 ps=1.31 w=0.98 l=3.47
X10 VIN.t7 VGP.t3 VOUT.t6 VCC.t1 sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=1.386 ps=8.73 w=8.4 l=3.34
X11 VIN.t8 VGP.t4 VOUT.t5 VCC.t0 sky130_fd_pr__pfet_01v8 ad=1.386 pd=8.73 as=1.386 ps=8.73 w=8.4 l=3.34
X12 VSS.t8 VSS.t5 VSS.t7 VSS.t6 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0 ps=0 w=0.98 l=3.47
X13 VOUT.t4 VGN.t4 VIN.t4 VSS.t0 sky130_fd_pr__nfet_01v8 ad=0.3822 pd=2.74 as=0.1617 ps=1.31 w=0.98 l=3.47
R0 VGP.n47 VGP.n46 161.3
R1 VGP.n45 VGP.n1 161.3
R2 VGP.n44 VGP.n43 161.3
R3 VGP.n42 VGP.n2 161.3
R4 VGP.n41 VGP.n40 161.3
R5 VGP.n39 VGP.n3 161.3
R6 VGP.n38 VGP.n37 161.3
R7 VGP.n36 VGP.n35 161.3
R8 VGP.n34 VGP.n5 161.3
R9 VGP.n33 VGP.n32 161.3
R10 VGP.n31 VGP.n6 161.3
R11 VGP.n30 VGP.n29 161.3
R12 VGP.n28 VGP.n7 161.3
R13 VGP.n27 VGP.n26 161.3
R14 VGP.n25 VGP.n8 161.3
R15 VGP.n24 VGP.n23 161.3
R16 VGP.n22 VGP.n9 161.3
R17 VGP.n21 VGP.n20 161.3
R18 VGP.n19 VGP.n10 161.3
R19 VGP.n18 VGP.n17 161.3
R20 VGP.n16 VGP.n11 161.3
R21 VGP.n15 VGP.n14 161.3
R22 VGP.n13 VGP.t0 93.6256
R23 VGP.n48 VGP.n0 73.3375
R24 VGP.n13 VGP.n12 65.9526
R25 VGP.n8 VGP.t2 60.6113
R26 VGP.n12 VGP.t3 60.6113
R27 VGP.n4 VGP.t4 60.6113
R28 VGP.n0 VGP.t1 60.6113
R29 VGP.n21 VGP.n10 56.4773
R30 VGP.n29 VGP.n6 56.4773
R31 VGP.n44 VGP.n2 40.8975
R32 VGP.n40 VGP.n2 39.9237
R33 VGP.n17 VGP.n10 24.3439
R34 VGP.n17 VGP.n16 24.3439
R35 VGP.n16 VGP.n15 24.3439
R36 VGP.n29 VGP.n28 24.3439
R37 VGP.n28 VGP.n27 24.3439
R38 VGP.n27 VGP.n8 24.3439
R39 VGP.n23 VGP.n8 24.3439
R40 VGP.n23 VGP.n22 24.3439
R41 VGP.n22 VGP.n21 24.3439
R42 VGP.n40 VGP.n39 24.3439
R43 VGP.n39 VGP.n38 24.3439
R44 VGP.n35 VGP.n34 24.3439
R45 VGP.n34 VGP.n33 24.3439
R46 VGP.n33 VGP.n6 24.3439
R47 VGP.n46 VGP.n45 24.3439
R48 VGP.n45 VGP.n44 24.3439
R49 VGP.n46 VGP.n0 16.554
R50 VGP.n38 VGP.n4 16.0672
R51 VGP.n15 VGP.n12 8.27727
R52 VGP.n35 VGP.n4 8.27727
R53 VGP.n14 VGP.n13 4.08017
R54 VGP VGP.n48 0.35776
R55 VGP.n48 VGP.n47 0.355081
R56 VGP.n47 VGP.n1 0.189894
R57 VGP.n43 VGP.n1 0.189894
R58 VGP.n43 VGP.n42 0.189894
R59 VGP.n42 VGP.n41 0.189894
R60 VGP.n41 VGP.n3 0.189894
R61 VGP.n37 VGP.n3 0.189894
R62 VGP.n37 VGP.n36 0.189894
R63 VGP.n36 VGP.n5 0.189894
R64 VGP.n32 VGP.n5 0.189894
R65 VGP.n32 VGP.n31 0.189894
R66 VGP.n31 VGP.n30 0.189894
R67 VGP.n30 VGP.n7 0.189894
R68 VGP.n26 VGP.n7 0.189894
R69 VGP.n26 VGP.n25 0.189894
R70 VGP.n25 VGP.n24 0.189894
R71 VGP.n24 VGP.n9 0.189894
R72 VGP.n20 VGP.n9 0.189894
R73 VGP.n20 VGP.n19 0.189894
R74 VGP.n19 VGP.n18 0.189894
R75 VGP.n18 VGP.n11 0.189894
R76 VGP.n14 VGP.n11 0.189894
R77 VIN.n5 VIN.t0 246.547
R78 VIN.n5 VIN.n4 223.066
R79 VIN.n7 VIN.n6 223.066
R80 VIN.n1 VIN.t9 69.7266
R81 VIN.n1 VIN.n0 62.6931
R82 VIN.n3 VIN.n2 62.6931
R83 VIN.n4 VIN.t2 20.2046
R84 VIN.n4 VIN.t1 20.2046
R85 VIN.n6 VIN.t4 20.2046
R86 VIN.n6 VIN.t3 20.2046
R87 VIN VIN.n3 13.0889
R88 VIN.n0 VIN.t6 3.87014
R89 VIN.n0 VIN.t7 3.87014
R90 VIN.n2 VIN.t5 3.87014
R91 VIN.n2 VIN.t8 3.87014
R92 VIN.n7 VIN.n5 3.27636
R93 VIN.n3 VIN.n1 3.16429
R94 VIN VIN.n7 1.64274
R95 VOUT.n5 VOUT.t4 263.224
R96 VOUT.n7 VOUT.n6 239.745
R97 VOUT.n5 VOUT.n4 239.745
R98 VOUT.n1 VOUT.t8 86.4052
R99 VOUT.n1 VOUT.n0 79.3719
R100 VOUT.n3 VOUT.n2 79.3719
R101 VOUT.n6 VOUT.t1 20.2046
R102 VOUT.n6 VOUT.t0 20.2046
R103 VOUT.n4 VOUT.t3 20.2046
R104 VOUT.n4 VOUT.t2 20.2046
R105 VOUT VOUT.n7 12.5371
R106 VOUT.n2 VOUT.t6 3.87014
R107 VOUT.n2 VOUT.t9 3.87014
R108 VOUT.n0 VOUT.t5 3.87014
R109 VOUT.n0 VOUT.t7 3.87014
R110 VOUT.n7 VOUT.n5 3.27636
R111 VOUT.n3 VOUT.n1 3.16429
R112 VOUT VOUT.n3 1.70309
R113 VCC.n515 VCC.n39 389.269
R114 VCC.n513 VCC.n43 389.269
R115 VCC.n252 VCC.n172 389.269
R116 VCC.n254 VCC.n170 389.269
R117 VCC.n448 VCC.t9 269.555
R118 VCC.n187 VCC.t5 269.555
R119 VCC.n513 VCC.n512 185
R120 VCC.n514 VCC.n513 185
R121 VCC.n44 VCC.n42 185
R122 VCC.n42 VCC.n40 185
R123 VCC.n431 VCC.n430 185
R124 VCC.n430 VCC.n429 185
R125 VCC.n47 VCC.n46 185
R126 VCC.n428 VCC.n47 185
R127 VCC.n426 VCC.n425 185
R128 VCC.n427 VCC.n426 185
R129 VCC.n51 VCC.n50 185
R130 VCC.n50 VCC.n49 185
R131 VCC.n421 VCC.n420 185
R132 VCC.n420 VCC.n419 185
R133 VCC.n54 VCC.n53 185
R134 VCC.n418 VCC.n54 185
R135 VCC.n416 VCC.n415 185
R136 VCC.n417 VCC.n416 185
R137 VCC.n58 VCC.n57 185
R138 VCC.n57 VCC.n56 185
R139 VCC.n411 VCC.n410 185
R140 VCC.n410 VCC.n409 185
R141 VCC.n61 VCC.n60 185
R142 VCC.n408 VCC.n61 185
R143 VCC.n406 VCC.n405 185
R144 VCC.n407 VCC.n406 185
R145 VCC.n65 VCC.n64 185
R146 VCC.n64 VCC.n63 185
R147 VCC.n401 VCC.n400 185
R148 VCC.n400 VCC.n399 185
R149 VCC.n68 VCC.n67 185
R150 VCC.n398 VCC.n68 185
R151 VCC.n396 VCC.n395 185
R152 VCC.n397 VCC.n396 185
R153 VCC.n72 VCC.n71 185
R154 VCC.n71 VCC.n70 185
R155 VCC.n391 VCC.n390 185
R156 VCC.n390 VCC.n389 185
R157 VCC.n75 VCC.n74 185
R158 VCC.n388 VCC.n75 185
R159 VCC.n386 VCC.n385 185
R160 VCC.n387 VCC.n386 185
R161 VCC.n77 VCC.n76 185
R162 VCC.n378 VCC.n76 185
R163 VCC.n381 VCC.n380 185
R164 VCC.n380 VCC.n379 185
R165 VCC.n80 VCC.n79 185
R166 VCC.n376 VCC.n80 185
R167 VCC.n374 VCC.n373 185
R168 VCC.n375 VCC.n374 185
R169 VCC.n84 VCC.n83 185
R170 VCC.n83 VCC.n82 185
R171 VCC.n369 VCC.n368 185
R172 VCC.n368 VCC.n367 185
R173 VCC.n87 VCC.n86 185
R174 VCC.n366 VCC.n87 185
R175 VCC.n365 VCC.n364 185
R176 VCC.t2 VCC.n365 185
R177 VCC.n90 VCC.n89 185
R178 VCC.n89 VCC.n88 185
R179 VCC.n360 VCC.n359 185
R180 VCC.n359 VCC.n358 185
R181 VCC.n93 VCC.n92 185
R182 VCC.n94 VCC.n93 185
R183 VCC.n349 VCC.n348 185
R184 VCC.n350 VCC.n349 185
R185 VCC.n103 VCC.n102 185
R186 VCC.n102 VCC.n101 185
R187 VCC.n344 VCC.n343 185
R188 VCC.n343 VCC.n342 185
R189 VCC.n106 VCC.n105 185
R190 VCC.n107 VCC.n106 185
R191 VCC.n333 VCC.n332 185
R192 VCC.n334 VCC.n333 185
R193 VCC.n115 VCC.n114 185
R194 VCC.n114 VCC.n113 185
R195 VCC.n328 VCC.n327 185
R196 VCC.n327 VCC.n326 185
R197 VCC.n118 VCC.n117 185
R198 VCC.n119 VCC.n118 185
R199 VCC.n317 VCC.n316 185
R200 VCC.n318 VCC.n317 185
R201 VCC.n127 VCC.n126 185
R202 VCC.n126 VCC.n125 185
R203 VCC.n312 VCC.n311 185
R204 VCC.n311 VCC.n310 185
R205 VCC.n130 VCC.n129 185
R206 VCC.n301 VCC.n130 185
R207 VCC.n300 VCC.n299 185
R208 VCC.n302 VCC.n300 185
R209 VCC.n138 VCC.n137 185
R210 VCC.n137 VCC.n136 185
R211 VCC.n295 VCC.n294 185
R212 VCC.n294 VCC.n293 185
R213 VCC.n141 VCC.n140 185
R214 VCC.n142 VCC.n141 185
R215 VCC.n284 VCC.n283 185
R216 VCC.n285 VCC.n284 185
R217 VCC.n150 VCC.n149 185
R218 VCC.n149 VCC.n148 185
R219 VCC.n279 VCC.n278 185
R220 VCC.n278 VCC.n277 185
R221 VCC.n153 VCC.n152 185
R222 VCC.n154 VCC.n153 185
R223 VCC.n268 VCC.n267 185
R224 VCC.n269 VCC.n268 185
R225 VCC.n161 VCC.n160 185
R226 VCC.n166 VCC.n160 185
R227 VCC.n263 VCC.n262 185
R228 VCC.n262 VCC.n261 185
R229 VCC.n164 VCC.n163 185
R230 VCC.n165 VCC.n164 185
R231 VCC.n252 VCC.n251 185
R232 VCC.n253 VCC.n252 185
R233 VCC.n255 VCC.n254 185
R234 VCC.n254 VCC.n253 185
R235 VCC.n168 VCC.n167 185
R236 VCC.n167 VCC.n165 185
R237 VCC.n260 VCC.n259 185
R238 VCC.n261 VCC.n260 185
R239 VCC.n159 VCC.n158 185
R240 VCC.n166 VCC.n159 185
R241 VCC.n271 VCC.n270 185
R242 VCC.n270 VCC.n269 185
R243 VCC.n156 VCC.n155 185
R244 VCC.n155 VCC.n154 185
R245 VCC.n276 VCC.n275 185
R246 VCC.n277 VCC.n276 185
R247 VCC.n147 VCC.n146 185
R248 VCC.n148 VCC.n147 185
R249 VCC.n287 VCC.n286 185
R250 VCC.n286 VCC.n285 185
R251 VCC.n144 VCC.n143 185
R252 VCC.n143 VCC.n142 185
R253 VCC.n292 VCC.n291 185
R254 VCC.n293 VCC.n292 185
R255 VCC.n135 VCC.n134 185
R256 VCC.n136 VCC.n135 185
R257 VCC.n304 VCC.n303 185
R258 VCC.n303 VCC.n302 185
R259 VCC.n132 VCC.n131 185
R260 VCC.n301 VCC.n131 185
R261 VCC.n309 VCC.n308 185
R262 VCC.n310 VCC.n309 185
R263 VCC.n124 VCC.n123 185
R264 VCC.n125 VCC.n124 185
R265 VCC.n320 VCC.n319 185
R266 VCC.n319 VCC.n318 185
R267 VCC.n121 VCC.n120 185
R268 VCC.n120 VCC.n119 185
R269 VCC.n325 VCC.n324 185
R270 VCC.n326 VCC.n325 185
R271 VCC.n112 VCC.n111 185
R272 VCC.n113 VCC.n112 185
R273 VCC.n336 VCC.n335 185
R274 VCC.n335 VCC.n334 185
R275 VCC.n109 VCC.n108 185
R276 VCC.n108 VCC.n107 185
R277 VCC.n341 VCC.n340 185
R278 VCC.n342 VCC.n341 185
R279 VCC.n100 VCC.n99 185
R280 VCC.n101 VCC.n100 185
R281 VCC.n352 VCC.n351 185
R282 VCC.n351 VCC.n350 185
R283 VCC.n97 VCC.n95 185
R284 VCC.n95 VCC.n94 185
R285 VCC.n357 VCC.n356 185
R286 VCC.n358 VCC.n357 185
R287 VCC.n96 VCC.n2 185
R288 VCC.n96 VCC.n88 185
R289 VCC.n558 VCC.n3 185
R290 VCC.t2 VCC.n3 185
R291 VCC.n557 VCC.n4 185
R292 VCC.n366 VCC.n4 185
R293 VCC.n556 VCC.n5 185
R294 VCC.n367 VCC.n5 185
R295 VCC.n81 VCC.n6 185
R296 VCC.n82 VCC.n81 185
R297 VCC.n552 VCC.n8 185
R298 VCC.n375 VCC.n8 185
R299 VCC.n551 VCC.n9 185
R300 VCC.n376 VCC.n9 185
R301 VCC.n550 VCC.n10 185
R302 VCC.n379 VCC.n10 185
R303 VCC.n377 VCC.n11 185
R304 VCC.n378 VCC.n377 185
R305 VCC.n546 VCC.n13 185
R306 VCC.n387 VCC.n13 185
R307 VCC.n545 VCC.n14 185
R308 VCC.n388 VCC.n14 185
R309 VCC.n544 VCC.n15 185
R310 VCC.n389 VCC.n15 185
R311 VCC.n69 VCC.n16 185
R312 VCC.n70 VCC.n69 185
R313 VCC.n540 VCC.n18 185
R314 VCC.n397 VCC.n18 185
R315 VCC.n539 VCC.n19 185
R316 VCC.n398 VCC.n19 185
R317 VCC.n538 VCC.n20 185
R318 VCC.n399 VCC.n20 185
R319 VCC.n62 VCC.n21 185
R320 VCC.n63 VCC.n62 185
R321 VCC.n534 VCC.n23 185
R322 VCC.n407 VCC.n23 185
R323 VCC.n533 VCC.n24 185
R324 VCC.n408 VCC.n24 185
R325 VCC.n532 VCC.n25 185
R326 VCC.n409 VCC.n25 185
R327 VCC.n55 VCC.n26 185
R328 VCC.n56 VCC.n55 185
R329 VCC.n528 VCC.n28 185
R330 VCC.n417 VCC.n28 185
R331 VCC.n527 VCC.n29 185
R332 VCC.n418 VCC.n29 185
R333 VCC.n526 VCC.n30 185
R334 VCC.n419 VCC.n30 185
R335 VCC.n48 VCC.n31 185
R336 VCC.n49 VCC.n48 185
R337 VCC.n522 VCC.n33 185
R338 VCC.n427 VCC.n33 185
R339 VCC.n521 VCC.n34 185
R340 VCC.n428 VCC.n34 185
R341 VCC.n520 VCC.n35 185
R342 VCC.n429 VCC.n35 185
R343 VCC.n38 VCC.n36 185
R344 VCC.n40 VCC.n38 185
R345 VCC.n516 VCC.n515 185
R346 VCC.n515 VCC.n514 185
R347 VCC.n510 VCC.n43 185
R348 VCC.n509 VCC.n508 185
R349 VCC.n506 VCC.n434 185
R350 VCC.n504 VCC.n503 185
R351 VCC.n502 VCC.n435 185
R352 VCC.n501 VCC.n500 185
R353 VCC.n498 VCC.n436 185
R354 VCC.n496 VCC.n495 185
R355 VCC.n494 VCC.n437 185
R356 VCC.n493 VCC.n492 185
R357 VCC.n490 VCC.n438 185
R358 VCC.n488 VCC.n487 185
R359 VCC.n486 VCC.n439 185
R360 VCC.n485 VCC.n484 185
R361 VCC.n482 VCC.n440 185
R362 VCC.n480 VCC.n479 185
R363 VCC.n478 VCC.n441 185
R364 VCC.n477 VCC.n476 185
R365 VCC.n474 VCC.n442 185
R366 VCC.n472 VCC.n471 185
R367 VCC.n470 VCC.n443 185
R368 VCC.n469 VCC.n468 185
R369 VCC.n466 VCC.n444 185
R370 VCC.n464 VCC.n463 185
R371 VCC.n462 VCC.n445 185
R372 VCC.n461 VCC.n460 185
R373 VCC.n458 VCC.n446 185
R374 VCC.n456 VCC.n455 185
R375 VCC.n454 VCC.n447 185
R376 VCC.n452 VCC.n451 185
R377 VCC.n39 VCC.n37 185
R378 VCC.n41 VCC.n39 185
R379 VCC.n170 VCC.n169 185
R380 VCC.n191 VCC.n190 185
R381 VCC.n193 VCC.n186 185
R382 VCC.n186 VCC.n171 185
R383 VCC.n195 VCC.n194 185
R384 VCC.n197 VCC.n185 185
R385 VCC.n200 VCC.n199 185
R386 VCC.n201 VCC.n184 185
R387 VCC.n203 VCC.n202 185
R388 VCC.n205 VCC.n183 185
R389 VCC.n208 VCC.n207 185
R390 VCC.n209 VCC.n182 185
R391 VCC.n211 VCC.n210 185
R392 VCC.n213 VCC.n181 185
R393 VCC.n216 VCC.n215 185
R394 VCC.n217 VCC.n180 185
R395 VCC.n219 VCC.n218 185
R396 VCC.n221 VCC.n179 185
R397 VCC.n224 VCC.n223 185
R398 VCC.n225 VCC.n178 185
R399 VCC.n227 VCC.n226 185
R400 VCC.n229 VCC.n177 185
R401 VCC.n232 VCC.n231 185
R402 VCC.n233 VCC.n176 185
R403 VCC.n235 VCC.n234 185
R404 VCC.n237 VCC.n175 185
R405 VCC.n240 VCC.n239 185
R406 VCC.n241 VCC.n174 185
R407 VCC.n243 VCC.n242 185
R408 VCC.n245 VCC.n173 185
R409 VCC.n248 VCC.n247 185
R410 VCC.n249 VCC.n172 185
R411 VCC.n448 VCC.t11 184.262
R412 VCC.n187 VCC.t8 184.262
R413 VCC.n252 VCC.n164 146.341
R414 VCC.n262 VCC.n164 146.341
R415 VCC.n262 VCC.n160 146.341
R416 VCC.n268 VCC.n160 146.341
R417 VCC.n268 VCC.n153 146.341
R418 VCC.n278 VCC.n153 146.341
R419 VCC.n278 VCC.n149 146.341
R420 VCC.n284 VCC.n149 146.341
R421 VCC.n284 VCC.n141 146.341
R422 VCC.n294 VCC.n141 146.341
R423 VCC.n294 VCC.n137 146.341
R424 VCC.n300 VCC.n137 146.341
R425 VCC.n300 VCC.n130 146.341
R426 VCC.n311 VCC.n130 146.341
R427 VCC.n311 VCC.n126 146.341
R428 VCC.n317 VCC.n126 146.341
R429 VCC.n317 VCC.n118 146.341
R430 VCC.n327 VCC.n118 146.341
R431 VCC.n327 VCC.n114 146.341
R432 VCC.n333 VCC.n114 146.341
R433 VCC.n333 VCC.n106 146.341
R434 VCC.n343 VCC.n106 146.341
R435 VCC.n343 VCC.n102 146.341
R436 VCC.n349 VCC.n102 146.341
R437 VCC.n349 VCC.n93 146.341
R438 VCC.n359 VCC.n93 146.341
R439 VCC.n359 VCC.n89 146.341
R440 VCC.n365 VCC.n89 146.341
R441 VCC.n365 VCC.n87 146.341
R442 VCC.n368 VCC.n87 146.341
R443 VCC.n368 VCC.n83 146.341
R444 VCC.n374 VCC.n83 146.341
R445 VCC.n374 VCC.n80 146.341
R446 VCC.n380 VCC.n80 146.341
R447 VCC.n380 VCC.n76 146.341
R448 VCC.n386 VCC.n76 146.341
R449 VCC.n386 VCC.n75 146.341
R450 VCC.n390 VCC.n75 146.341
R451 VCC.n390 VCC.n71 146.341
R452 VCC.n396 VCC.n71 146.341
R453 VCC.n396 VCC.n68 146.341
R454 VCC.n400 VCC.n68 146.341
R455 VCC.n400 VCC.n64 146.341
R456 VCC.n406 VCC.n64 146.341
R457 VCC.n406 VCC.n61 146.341
R458 VCC.n410 VCC.n61 146.341
R459 VCC.n410 VCC.n57 146.341
R460 VCC.n416 VCC.n57 146.341
R461 VCC.n416 VCC.n54 146.341
R462 VCC.n420 VCC.n54 146.341
R463 VCC.n420 VCC.n50 146.341
R464 VCC.n426 VCC.n50 146.341
R465 VCC.n426 VCC.n47 146.341
R466 VCC.n430 VCC.n47 146.341
R467 VCC.n430 VCC.n42 146.341
R468 VCC.n513 VCC.n42 146.341
R469 VCC.n254 VCC.n167 146.341
R470 VCC.n260 VCC.n167 146.341
R471 VCC.n260 VCC.n159 146.341
R472 VCC.n270 VCC.n159 146.341
R473 VCC.n270 VCC.n155 146.341
R474 VCC.n276 VCC.n155 146.341
R475 VCC.n276 VCC.n147 146.341
R476 VCC.n286 VCC.n147 146.341
R477 VCC.n286 VCC.n143 146.341
R478 VCC.n292 VCC.n143 146.341
R479 VCC.n292 VCC.n135 146.341
R480 VCC.n303 VCC.n135 146.341
R481 VCC.n303 VCC.n131 146.341
R482 VCC.n309 VCC.n131 146.341
R483 VCC.n309 VCC.n124 146.341
R484 VCC.n319 VCC.n124 146.341
R485 VCC.n319 VCC.n120 146.341
R486 VCC.n325 VCC.n120 146.341
R487 VCC.n325 VCC.n112 146.341
R488 VCC.n335 VCC.n112 146.341
R489 VCC.n335 VCC.n108 146.341
R490 VCC.n341 VCC.n108 146.341
R491 VCC.n341 VCC.n100 146.341
R492 VCC.n351 VCC.n100 146.341
R493 VCC.n351 VCC.n95 146.341
R494 VCC.n357 VCC.n95 146.341
R495 VCC.n357 VCC.n96 146.341
R496 VCC.n96 VCC.n3 146.341
R497 VCC.n4 VCC.n3 146.341
R498 VCC.n5 VCC.n4 146.341
R499 VCC.n81 VCC.n5 146.341
R500 VCC.n81 VCC.n8 146.341
R501 VCC.n9 VCC.n8 146.341
R502 VCC.n10 VCC.n9 146.341
R503 VCC.n377 VCC.n10 146.341
R504 VCC.n377 VCC.n13 146.341
R505 VCC.n14 VCC.n13 146.341
R506 VCC.n15 VCC.n14 146.341
R507 VCC.n69 VCC.n15 146.341
R508 VCC.n69 VCC.n18 146.341
R509 VCC.n19 VCC.n18 146.341
R510 VCC.n20 VCC.n19 146.341
R511 VCC.n62 VCC.n20 146.341
R512 VCC.n62 VCC.n23 146.341
R513 VCC.n24 VCC.n23 146.341
R514 VCC.n25 VCC.n24 146.341
R515 VCC.n55 VCC.n25 146.341
R516 VCC.n55 VCC.n28 146.341
R517 VCC.n29 VCC.n28 146.341
R518 VCC.n30 VCC.n29 146.341
R519 VCC.n48 VCC.n30 146.341
R520 VCC.n48 VCC.n33 146.341
R521 VCC.n34 VCC.n33 146.341
R522 VCC.n35 VCC.n34 146.341
R523 VCC.n38 VCC.n35 146.341
R524 VCC.n515 VCC.n38 146.341
R525 VCC.n449 VCC.t12 113.085
R526 VCC.n188 VCC.t7 113.085
R527 VCC.n451 VCC.n39 99.5127
R528 VCC.n456 VCC.n447 99.5127
R529 VCC.n460 VCC.n458 99.5127
R530 VCC.n464 VCC.n445 99.5127
R531 VCC.n468 VCC.n466 99.5127
R532 VCC.n472 VCC.n443 99.5127
R533 VCC.n476 VCC.n474 99.5127
R534 VCC.n480 VCC.n441 99.5127
R535 VCC.n484 VCC.n482 99.5127
R536 VCC.n488 VCC.n439 99.5127
R537 VCC.n492 VCC.n490 99.5127
R538 VCC.n496 VCC.n437 99.5127
R539 VCC.n500 VCC.n498 99.5127
R540 VCC.n504 VCC.n435 99.5127
R541 VCC.n508 VCC.n506 99.5127
R542 VCC.n190 VCC.n186 99.5127
R543 VCC.n195 VCC.n186 99.5127
R544 VCC.n199 VCC.n197 99.5127
R545 VCC.n203 VCC.n184 99.5127
R546 VCC.n207 VCC.n205 99.5127
R547 VCC.n211 VCC.n182 99.5127
R548 VCC.n215 VCC.n213 99.5127
R549 VCC.n219 VCC.n180 99.5127
R550 VCC.n223 VCC.n221 99.5127
R551 VCC.n227 VCC.n178 99.5127
R552 VCC.n231 VCC.n229 99.5127
R553 VCC.n235 VCC.n176 99.5127
R554 VCC.n239 VCC.n237 99.5127
R555 VCC.n243 VCC.n174 99.5127
R556 VCC.n247 VCC.n245 99.5127
R557 VCC.n507 VCC.n41 72.8958
R558 VCC.n505 VCC.n41 72.8958
R559 VCC.n499 VCC.n41 72.8958
R560 VCC.n497 VCC.n41 72.8958
R561 VCC.n491 VCC.n41 72.8958
R562 VCC.n489 VCC.n41 72.8958
R563 VCC.n483 VCC.n41 72.8958
R564 VCC.n481 VCC.n41 72.8958
R565 VCC.n475 VCC.n41 72.8958
R566 VCC.n473 VCC.n41 72.8958
R567 VCC.n467 VCC.n41 72.8958
R568 VCC.n465 VCC.n41 72.8958
R569 VCC.n459 VCC.n41 72.8958
R570 VCC.n457 VCC.n41 72.8958
R571 VCC.n450 VCC.n41 72.8958
R572 VCC.n189 VCC.n171 72.8958
R573 VCC.n196 VCC.n171 72.8958
R574 VCC.n198 VCC.n171 72.8958
R575 VCC.n204 VCC.n171 72.8958
R576 VCC.n206 VCC.n171 72.8958
R577 VCC.n212 VCC.n171 72.8958
R578 VCC.n214 VCC.n171 72.8958
R579 VCC.n220 VCC.n171 72.8958
R580 VCC.n222 VCC.n171 72.8958
R581 VCC.n228 VCC.n171 72.8958
R582 VCC.n230 VCC.n171 72.8958
R583 VCC.n236 VCC.n171 72.8958
R584 VCC.n238 VCC.n171 72.8958
R585 VCC.n244 VCC.n171 72.8958
R586 VCC.n246 VCC.n171 72.8958
R587 VCC.n449 VCC.n448 71.1763
R588 VCC.n188 VCC.n187 71.1763
R589 VCC.n253 VCC.n171 67.9661
R590 VCC.n514 VCC.n41 67.9661
R591 VCC.n450 VCC.n447 39.2114
R592 VCC.n458 VCC.n457 39.2114
R593 VCC.n459 VCC.n445 39.2114
R594 VCC.n466 VCC.n465 39.2114
R595 VCC.n467 VCC.n443 39.2114
R596 VCC.n474 VCC.n473 39.2114
R597 VCC.n475 VCC.n441 39.2114
R598 VCC.n482 VCC.n481 39.2114
R599 VCC.n483 VCC.n439 39.2114
R600 VCC.n490 VCC.n489 39.2114
R601 VCC.n491 VCC.n437 39.2114
R602 VCC.n498 VCC.n497 39.2114
R603 VCC.n499 VCC.n435 39.2114
R604 VCC.n506 VCC.n505 39.2114
R605 VCC.n507 VCC.n43 39.2114
R606 VCC.n189 VCC.n170 39.2114
R607 VCC.n196 VCC.n195 39.2114
R608 VCC.n199 VCC.n198 39.2114
R609 VCC.n204 VCC.n203 39.2114
R610 VCC.n207 VCC.n206 39.2114
R611 VCC.n212 VCC.n211 39.2114
R612 VCC.n215 VCC.n214 39.2114
R613 VCC.n220 VCC.n219 39.2114
R614 VCC.n223 VCC.n222 39.2114
R615 VCC.n228 VCC.n227 39.2114
R616 VCC.n231 VCC.n230 39.2114
R617 VCC.n236 VCC.n235 39.2114
R618 VCC.n239 VCC.n238 39.2114
R619 VCC.n244 VCC.n243 39.2114
R620 VCC.n247 VCC.n246 39.2114
R621 VCC.n508 VCC.n507 39.2114
R622 VCC.n505 VCC.n504 39.2114
R623 VCC.n500 VCC.n499 39.2114
R624 VCC.n497 VCC.n496 39.2114
R625 VCC.n492 VCC.n491 39.2114
R626 VCC.n489 VCC.n488 39.2114
R627 VCC.n484 VCC.n483 39.2114
R628 VCC.n481 VCC.n480 39.2114
R629 VCC.n476 VCC.n475 39.2114
R630 VCC.n473 VCC.n472 39.2114
R631 VCC.n468 VCC.n467 39.2114
R632 VCC.n465 VCC.n464 39.2114
R633 VCC.n460 VCC.n459 39.2114
R634 VCC.n457 VCC.n456 39.2114
R635 VCC.n451 VCC.n450 39.2114
R636 VCC.n190 VCC.n189 39.2114
R637 VCC.n197 VCC.n196 39.2114
R638 VCC.n198 VCC.n184 39.2114
R639 VCC.n205 VCC.n204 39.2114
R640 VCC.n206 VCC.n182 39.2114
R641 VCC.n213 VCC.n212 39.2114
R642 VCC.n214 VCC.n180 39.2114
R643 VCC.n221 VCC.n220 39.2114
R644 VCC.n222 VCC.n178 39.2114
R645 VCC.n229 VCC.n228 39.2114
R646 VCC.n230 VCC.n176 39.2114
R647 VCC.n237 VCC.n236 39.2114
R648 VCC.n238 VCC.n174 39.2114
R649 VCC.n245 VCC.n244 39.2114
R650 VCC.n246 VCC.n172 39.2114
R651 VCC.n253 VCC.n165 37.9701
R652 VCC.n261 VCC.n165 37.9701
R653 VCC.n261 VCC.n166 37.9701
R654 VCC.n269 VCC.n154 37.9701
R655 VCC.n277 VCC.n154 37.9701
R656 VCC.n277 VCC.n148 37.9701
R657 VCC.n285 VCC.n148 37.9701
R658 VCC.n285 VCC.n142 37.9701
R659 VCC.n293 VCC.n142 37.9701
R660 VCC.n293 VCC.n136 37.9701
R661 VCC.n302 VCC.n136 37.9701
R662 VCC.n302 VCC.n301 37.9701
R663 VCC.n310 VCC.n125 37.9701
R664 VCC.n318 VCC.n125 37.9701
R665 VCC.n318 VCC.n119 37.9701
R666 VCC.n326 VCC.n119 37.9701
R667 VCC.n326 VCC.n113 37.9701
R668 VCC.n334 VCC.n113 37.9701
R669 VCC.n342 VCC.n107 37.9701
R670 VCC.n342 VCC.n101 37.9701
R671 VCC.n350 VCC.n101 37.9701
R672 VCC.n350 VCC.n94 37.9701
R673 VCC.n358 VCC.n94 37.9701
R674 VCC.n358 VCC.n88 37.9701
R675 VCC.t2 VCC.n88 37.9701
R676 VCC.n366 VCC.t2 37.9701
R677 VCC.n367 VCC.n366 37.9701
R678 VCC.n367 VCC.n82 37.9701
R679 VCC.n375 VCC.n82 37.9701
R680 VCC.n376 VCC.n375 37.9701
R681 VCC.n379 VCC.n376 37.9701
R682 VCC.n379 VCC.n378 37.9701
R683 VCC.n388 VCC.n387 37.9701
R684 VCC.n389 VCC.n388 37.9701
R685 VCC.n389 VCC.n70 37.9701
R686 VCC.n397 VCC.n70 37.9701
R687 VCC.n398 VCC.n397 37.9701
R688 VCC.n399 VCC.n398 37.9701
R689 VCC.n407 VCC.n63 37.9701
R690 VCC.n408 VCC.n407 37.9701
R691 VCC.n409 VCC.n408 37.9701
R692 VCC.n409 VCC.n56 37.9701
R693 VCC.n417 VCC.n56 37.9701
R694 VCC.n418 VCC.n417 37.9701
R695 VCC.n419 VCC.n418 37.9701
R696 VCC.n419 VCC.n49 37.9701
R697 VCC.n427 VCC.n49 37.9701
R698 VCC.n429 VCC.n428 37.9701
R699 VCC.n429 VCC.n40 37.9701
R700 VCC.n514 VCC.n40 37.9701
R701 VCC.n166 VCC.t6 30.3762
R702 VCC.n428 VCC.t10 30.3762
R703 VCC.n517 VCC.n37 29.5539
R704 VCC.n511 VCC.n510 29.5539
R705 VCC.n256 VCC.n169 29.5539
R706 VCC.n250 VCC.n249 29.5539
R707 VCC.n453 VCC.n449 29.2853
R708 VCC.n192 VCC.n188 29.2853
R709 VCC.n310 VCC.t3 25.8198
R710 VCC.n399 VCC.t4 25.8198
R711 VCC.n334 VCC.t0 25.0605
R712 VCC.n387 VCC.t1 25.0605
R713 VCC.n251 VCC.n163 19.3944
R714 VCC.n263 VCC.n163 19.3944
R715 VCC.n263 VCC.n161 19.3944
R716 VCC.n267 VCC.n161 19.3944
R717 VCC.n267 VCC.n152 19.3944
R718 VCC.n279 VCC.n152 19.3944
R719 VCC.n279 VCC.n150 19.3944
R720 VCC.n283 VCC.n150 19.3944
R721 VCC.n283 VCC.n140 19.3944
R722 VCC.n295 VCC.n140 19.3944
R723 VCC.n295 VCC.n138 19.3944
R724 VCC.n299 VCC.n138 19.3944
R725 VCC.n299 VCC.n129 19.3944
R726 VCC.n312 VCC.n129 19.3944
R727 VCC.n312 VCC.n127 19.3944
R728 VCC.n316 VCC.n127 19.3944
R729 VCC.n316 VCC.n117 19.3944
R730 VCC.n328 VCC.n117 19.3944
R731 VCC.n328 VCC.n115 19.3944
R732 VCC.n332 VCC.n115 19.3944
R733 VCC.n332 VCC.n105 19.3944
R734 VCC.n344 VCC.n105 19.3944
R735 VCC.n344 VCC.n103 19.3944
R736 VCC.n348 VCC.n103 19.3944
R737 VCC.n348 VCC.n92 19.3944
R738 VCC.n360 VCC.n92 19.3944
R739 VCC.n360 VCC.n90 19.3944
R740 VCC.n364 VCC.n90 19.3944
R741 VCC.n364 VCC.n86 19.3944
R742 VCC.n369 VCC.n86 19.3944
R743 VCC.n369 VCC.n84 19.3944
R744 VCC.n373 VCC.n84 19.3944
R745 VCC.n373 VCC.n79 19.3944
R746 VCC.n381 VCC.n79 19.3944
R747 VCC.n381 VCC.n77 19.3944
R748 VCC.n385 VCC.n77 19.3944
R749 VCC.n385 VCC.n74 19.3944
R750 VCC.n391 VCC.n74 19.3944
R751 VCC.n391 VCC.n72 19.3944
R752 VCC.n395 VCC.n72 19.3944
R753 VCC.n395 VCC.n67 19.3944
R754 VCC.n401 VCC.n67 19.3944
R755 VCC.n401 VCC.n65 19.3944
R756 VCC.n405 VCC.n65 19.3944
R757 VCC.n405 VCC.n60 19.3944
R758 VCC.n411 VCC.n60 19.3944
R759 VCC.n411 VCC.n58 19.3944
R760 VCC.n415 VCC.n58 19.3944
R761 VCC.n415 VCC.n53 19.3944
R762 VCC.n421 VCC.n53 19.3944
R763 VCC.n421 VCC.n51 19.3944
R764 VCC.n425 VCC.n51 19.3944
R765 VCC.n425 VCC.n46 19.3944
R766 VCC.n431 VCC.n46 19.3944
R767 VCC.n431 VCC.n44 19.3944
R768 VCC.n512 VCC.n44 19.3944
R769 VCC.n255 VCC.n168 19.3944
R770 VCC.n259 VCC.n168 19.3944
R771 VCC.n259 VCC.n158 19.3944
R772 VCC.n271 VCC.n158 19.3944
R773 VCC.n271 VCC.n156 19.3944
R774 VCC.n275 VCC.n156 19.3944
R775 VCC.n275 VCC.n146 19.3944
R776 VCC.n287 VCC.n146 19.3944
R777 VCC.n287 VCC.n144 19.3944
R778 VCC.n291 VCC.n144 19.3944
R779 VCC.n291 VCC.n134 19.3944
R780 VCC.n304 VCC.n134 19.3944
R781 VCC.n304 VCC.n132 19.3944
R782 VCC.n308 VCC.n132 19.3944
R783 VCC.n308 VCC.n123 19.3944
R784 VCC.n320 VCC.n123 19.3944
R785 VCC.n320 VCC.n121 19.3944
R786 VCC.n324 VCC.n121 19.3944
R787 VCC.n324 VCC.n111 19.3944
R788 VCC.n336 VCC.n111 19.3944
R789 VCC.n336 VCC.n109 19.3944
R790 VCC.n340 VCC.n109 19.3944
R791 VCC.n340 VCC.n99 19.3944
R792 VCC.n352 VCC.n99 19.3944
R793 VCC.n352 VCC.n97 19.3944
R794 VCC.n356 VCC.n97 19.3944
R795 VCC.n356 VCC.n2 19.3944
R796 VCC.n558 VCC.n2 19.3944
R797 VCC.n558 VCC.n557 19.3944
R798 VCC.n557 VCC.n556 19.3944
R799 VCC.n556 VCC.n6 19.3944
R800 VCC.n552 VCC.n6 19.3944
R801 VCC.n552 VCC.n551 19.3944
R802 VCC.n551 VCC.n550 19.3944
R803 VCC.n550 VCC.n11 19.3944
R804 VCC.n546 VCC.n11 19.3944
R805 VCC.n546 VCC.n545 19.3944
R806 VCC.n545 VCC.n544 19.3944
R807 VCC.n544 VCC.n16 19.3944
R808 VCC.n540 VCC.n16 19.3944
R809 VCC.n540 VCC.n539 19.3944
R810 VCC.n539 VCC.n538 19.3944
R811 VCC.n538 VCC.n21 19.3944
R812 VCC.n534 VCC.n21 19.3944
R813 VCC.n534 VCC.n533 19.3944
R814 VCC.n533 VCC.n532 19.3944
R815 VCC.n532 VCC.n26 19.3944
R816 VCC.n528 VCC.n26 19.3944
R817 VCC.n528 VCC.n527 19.3944
R818 VCC.n527 VCC.n526 19.3944
R819 VCC.n526 VCC.n31 19.3944
R820 VCC.n522 VCC.n31 19.3944
R821 VCC.n522 VCC.n521 19.3944
R822 VCC.n521 VCC.n520 19.3944
R823 VCC.n520 VCC.n36 19.3944
R824 VCC.n516 VCC.n36 19.3944
R825 VCC.t0 VCC.n107 12.9102
R826 VCC.n378 VCC.t1 12.9102
R827 VCC.n301 VCC.t3 12.1508
R828 VCC.t4 VCC.n63 12.1508
R829 VCC.n452 VCC.n37 10.6151
R830 VCC.n455 VCC.n454 10.6151
R831 VCC.n455 VCC.n446 10.6151
R832 VCC.n461 VCC.n446 10.6151
R833 VCC.n462 VCC.n461 10.6151
R834 VCC.n463 VCC.n462 10.6151
R835 VCC.n463 VCC.n444 10.6151
R836 VCC.n469 VCC.n444 10.6151
R837 VCC.n470 VCC.n469 10.6151
R838 VCC.n471 VCC.n470 10.6151
R839 VCC.n471 VCC.n442 10.6151
R840 VCC.n477 VCC.n442 10.6151
R841 VCC.n478 VCC.n477 10.6151
R842 VCC.n479 VCC.n478 10.6151
R843 VCC.n479 VCC.n440 10.6151
R844 VCC.n485 VCC.n440 10.6151
R845 VCC.n486 VCC.n485 10.6151
R846 VCC.n487 VCC.n486 10.6151
R847 VCC.n487 VCC.n438 10.6151
R848 VCC.n493 VCC.n438 10.6151
R849 VCC.n494 VCC.n493 10.6151
R850 VCC.n495 VCC.n494 10.6151
R851 VCC.n495 VCC.n436 10.6151
R852 VCC.n501 VCC.n436 10.6151
R853 VCC.n502 VCC.n501 10.6151
R854 VCC.n503 VCC.n502 10.6151
R855 VCC.n503 VCC.n434 10.6151
R856 VCC.n509 VCC.n434 10.6151
R857 VCC.n510 VCC.n509 10.6151
R858 VCC.n191 VCC.n169 10.6151
R859 VCC.n194 VCC.n193 10.6151
R860 VCC.n194 VCC.n185 10.6151
R861 VCC.n200 VCC.n185 10.6151
R862 VCC.n201 VCC.n200 10.6151
R863 VCC.n202 VCC.n201 10.6151
R864 VCC.n202 VCC.n183 10.6151
R865 VCC.n208 VCC.n183 10.6151
R866 VCC.n209 VCC.n208 10.6151
R867 VCC.n210 VCC.n209 10.6151
R868 VCC.n210 VCC.n181 10.6151
R869 VCC.n216 VCC.n181 10.6151
R870 VCC.n217 VCC.n216 10.6151
R871 VCC.n218 VCC.n217 10.6151
R872 VCC.n218 VCC.n179 10.6151
R873 VCC.n224 VCC.n179 10.6151
R874 VCC.n225 VCC.n224 10.6151
R875 VCC.n226 VCC.n225 10.6151
R876 VCC.n226 VCC.n177 10.6151
R877 VCC.n232 VCC.n177 10.6151
R878 VCC.n233 VCC.n232 10.6151
R879 VCC.n234 VCC.n233 10.6151
R880 VCC.n234 VCC.n175 10.6151
R881 VCC.n240 VCC.n175 10.6151
R882 VCC.n241 VCC.n240 10.6151
R883 VCC.n242 VCC.n241 10.6151
R884 VCC.n242 VCC.n173 10.6151
R885 VCC.n248 VCC.n173 10.6151
R886 VCC.n249 VCC.n248 10.6151
R887 VCC.n557 VCC.n0 9.3005
R888 VCC.n556 VCC.n555 9.3005
R889 VCC.n554 VCC.n6 9.3005
R890 VCC.n553 VCC.n552 9.3005
R891 VCC.n551 VCC.n7 9.3005
R892 VCC.n550 VCC.n549 9.3005
R893 VCC.n548 VCC.n11 9.3005
R894 VCC.n547 VCC.n546 9.3005
R895 VCC.n545 VCC.n12 9.3005
R896 VCC.n544 VCC.n543 9.3005
R897 VCC.n542 VCC.n16 9.3005
R898 VCC.n541 VCC.n540 9.3005
R899 VCC.n539 VCC.n17 9.3005
R900 VCC.n538 VCC.n537 9.3005
R901 VCC.n536 VCC.n21 9.3005
R902 VCC.n535 VCC.n534 9.3005
R903 VCC.n533 VCC.n22 9.3005
R904 VCC.n532 VCC.n531 9.3005
R905 VCC.n530 VCC.n26 9.3005
R906 VCC.n529 VCC.n528 9.3005
R907 VCC.n527 VCC.n27 9.3005
R908 VCC.n526 VCC.n525 9.3005
R909 VCC.n524 VCC.n31 9.3005
R910 VCC.n523 VCC.n522 9.3005
R911 VCC.n521 VCC.n32 9.3005
R912 VCC.n520 VCC.n519 9.3005
R913 VCC.n518 VCC.n36 9.3005
R914 VCC.n517 VCC.n516 9.3005
R915 VCC.n163 VCC.n162 9.3005
R916 VCC.n264 VCC.n263 9.3005
R917 VCC.n265 VCC.n161 9.3005
R918 VCC.n267 VCC.n266 9.3005
R919 VCC.n152 VCC.n151 9.3005
R920 VCC.n280 VCC.n279 9.3005
R921 VCC.n281 VCC.n150 9.3005
R922 VCC.n283 VCC.n282 9.3005
R923 VCC.n140 VCC.n139 9.3005
R924 VCC.n296 VCC.n295 9.3005
R925 VCC.n297 VCC.n138 9.3005
R926 VCC.n299 VCC.n298 9.3005
R927 VCC.n129 VCC.n128 9.3005
R928 VCC.n313 VCC.n312 9.3005
R929 VCC.n314 VCC.n127 9.3005
R930 VCC.n316 VCC.n315 9.3005
R931 VCC.n117 VCC.n116 9.3005
R932 VCC.n329 VCC.n328 9.3005
R933 VCC.n330 VCC.n115 9.3005
R934 VCC.n332 VCC.n331 9.3005
R935 VCC.n105 VCC.n104 9.3005
R936 VCC.n345 VCC.n344 9.3005
R937 VCC.n346 VCC.n103 9.3005
R938 VCC.n348 VCC.n347 9.3005
R939 VCC.n92 VCC.n91 9.3005
R940 VCC.n361 VCC.n360 9.3005
R941 VCC.n362 VCC.n90 9.3005
R942 VCC.n364 VCC.n363 9.3005
R943 VCC.n86 VCC.n85 9.3005
R944 VCC.n370 VCC.n369 9.3005
R945 VCC.n371 VCC.n84 9.3005
R946 VCC.n373 VCC.n372 9.3005
R947 VCC.n79 VCC.n78 9.3005
R948 VCC.n382 VCC.n381 9.3005
R949 VCC.n383 VCC.n77 9.3005
R950 VCC.n385 VCC.n384 9.3005
R951 VCC.n74 VCC.n73 9.3005
R952 VCC.n392 VCC.n391 9.3005
R953 VCC.n393 VCC.n72 9.3005
R954 VCC.n395 VCC.n394 9.3005
R955 VCC.n67 VCC.n66 9.3005
R956 VCC.n402 VCC.n401 9.3005
R957 VCC.n403 VCC.n65 9.3005
R958 VCC.n405 VCC.n404 9.3005
R959 VCC.n60 VCC.n59 9.3005
R960 VCC.n412 VCC.n411 9.3005
R961 VCC.n413 VCC.n58 9.3005
R962 VCC.n415 VCC.n414 9.3005
R963 VCC.n53 VCC.n52 9.3005
R964 VCC.n422 VCC.n421 9.3005
R965 VCC.n423 VCC.n51 9.3005
R966 VCC.n425 VCC.n424 9.3005
R967 VCC.n46 VCC.n45 9.3005
R968 VCC.n432 VCC.n431 9.3005
R969 VCC.n433 VCC.n44 9.3005
R970 VCC.n512 VCC.n511 9.3005
R971 VCC.n251 VCC.n250 9.3005
R972 VCC.n256 VCC.n255 9.3005
R973 VCC.n257 VCC.n168 9.3005
R974 VCC.n259 VCC.n258 9.3005
R975 VCC.n158 VCC.n157 9.3005
R976 VCC.n272 VCC.n271 9.3005
R977 VCC.n273 VCC.n156 9.3005
R978 VCC.n275 VCC.n274 9.3005
R979 VCC.n146 VCC.n145 9.3005
R980 VCC.n288 VCC.n287 9.3005
R981 VCC.n289 VCC.n144 9.3005
R982 VCC.n291 VCC.n290 9.3005
R983 VCC.n134 VCC.n133 9.3005
R984 VCC.n305 VCC.n304 9.3005
R985 VCC.n306 VCC.n132 9.3005
R986 VCC.n308 VCC.n307 9.3005
R987 VCC.n123 VCC.n122 9.3005
R988 VCC.n321 VCC.n320 9.3005
R989 VCC.n322 VCC.n121 9.3005
R990 VCC.n324 VCC.n323 9.3005
R991 VCC.n111 VCC.n110 9.3005
R992 VCC.n337 VCC.n336 9.3005
R993 VCC.n338 VCC.n109 9.3005
R994 VCC.n340 VCC.n339 9.3005
R995 VCC.n99 VCC.n98 9.3005
R996 VCC.n353 VCC.n352 9.3005
R997 VCC.n354 VCC.n97 9.3005
R998 VCC.n356 VCC.n355 9.3005
R999 VCC.n2 VCC.n1 9.3005
R1000 VCC.n559 VCC.n558 9.3005
R1001 VCC.n269 VCC.t6 7.59442
R1002 VCC.t10 VCC.n427 7.59442
R1003 VCC.n453 VCC.n452 6.7127
R1004 VCC.n192 VCC.n191 6.7127
R1005 VCC.n454 VCC.n453 3.90294
R1006 VCC.n193 VCC.n192 3.90294
R1007 VCC.n555 VCC.n0 0.152939
R1008 VCC.n555 VCC.n554 0.152939
R1009 VCC.n554 VCC.n553 0.152939
R1010 VCC.n553 VCC.n7 0.152939
R1011 VCC.n549 VCC.n7 0.152939
R1012 VCC.n549 VCC.n548 0.152939
R1013 VCC.n548 VCC.n547 0.152939
R1014 VCC.n547 VCC.n12 0.152939
R1015 VCC.n543 VCC.n12 0.152939
R1016 VCC.n543 VCC.n542 0.152939
R1017 VCC.n542 VCC.n541 0.152939
R1018 VCC.n541 VCC.n17 0.152939
R1019 VCC.n537 VCC.n17 0.152939
R1020 VCC.n537 VCC.n536 0.152939
R1021 VCC.n536 VCC.n535 0.152939
R1022 VCC.n535 VCC.n22 0.152939
R1023 VCC.n531 VCC.n22 0.152939
R1024 VCC.n531 VCC.n530 0.152939
R1025 VCC.n530 VCC.n529 0.152939
R1026 VCC.n529 VCC.n27 0.152939
R1027 VCC.n525 VCC.n27 0.152939
R1028 VCC.n525 VCC.n524 0.152939
R1029 VCC.n524 VCC.n523 0.152939
R1030 VCC.n523 VCC.n32 0.152939
R1031 VCC.n519 VCC.n32 0.152939
R1032 VCC.n519 VCC.n518 0.152939
R1033 VCC.n518 VCC.n517 0.152939
R1034 VCC.n250 VCC.n162 0.152939
R1035 VCC.n264 VCC.n162 0.152939
R1036 VCC.n265 VCC.n264 0.152939
R1037 VCC.n266 VCC.n265 0.152939
R1038 VCC.n266 VCC.n151 0.152939
R1039 VCC.n280 VCC.n151 0.152939
R1040 VCC.n281 VCC.n280 0.152939
R1041 VCC.n282 VCC.n281 0.152939
R1042 VCC.n282 VCC.n139 0.152939
R1043 VCC.n296 VCC.n139 0.152939
R1044 VCC.n297 VCC.n296 0.152939
R1045 VCC.n298 VCC.n297 0.152939
R1046 VCC.n298 VCC.n128 0.152939
R1047 VCC.n313 VCC.n128 0.152939
R1048 VCC.n314 VCC.n313 0.152939
R1049 VCC.n315 VCC.n314 0.152939
R1050 VCC.n315 VCC.n116 0.152939
R1051 VCC.n329 VCC.n116 0.152939
R1052 VCC.n330 VCC.n329 0.152939
R1053 VCC.n331 VCC.n330 0.152939
R1054 VCC.n331 VCC.n104 0.152939
R1055 VCC.n345 VCC.n104 0.152939
R1056 VCC.n346 VCC.n345 0.152939
R1057 VCC.n347 VCC.n346 0.152939
R1058 VCC.n347 VCC.n91 0.152939
R1059 VCC.n361 VCC.n91 0.152939
R1060 VCC.n362 VCC.n361 0.152939
R1061 VCC.n363 VCC.n362 0.152939
R1062 VCC.n363 VCC.n85 0.152939
R1063 VCC.n370 VCC.n85 0.152939
R1064 VCC.n371 VCC.n370 0.152939
R1065 VCC.n372 VCC.n371 0.152939
R1066 VCC.n372 VCC.n78 0.152939
R1067 VCC.n382 VCC.n78 0.152939
R1068 VCC.n383 VCC.n382 0.152939
R1069 VCC.n384 VCC.n383 0.152939
R1070 VCC.n384 VCC.n73 0.152939
R1071 VCC.n392 VCC.n73 0.152939
R1072 VCC.n393 VCC.n392 0.152939
R1073 VCC.n394 VCC.n393 0.152939
R1074 VCC.n394 VCC.n66 0.152939
R1075 VCC.n402 VCC.n66 0.152939
R1076 VCC.n403 VCC.n402 0.152939
R1077 VCC.n404 VCC.n403 0.152939
R1078 VCC.n404 VCC.n59 0.152939
R1079 VCC.n412 VCC.n59 0.152939
R1080 VCC.n413 VCC.n412 0.152939
R1081 VCC.n414 VCC.n413 0.152939
R1082 VCC.n414 VCC.n52 0.152939
R1083 VCC.n422 VCC.n52 0.152939
R1084 VCC.n423 VCC.n422 0.152939
R1085 VCC.n424 VCC.n423 0.152939
R1086 VCC.n424 VCC.n45 0.152939
R1087 VCC.n432 VCC.n45 0.152939
R1088 VCC.n433 VCC.n432 0.152939
R1089 VCC.n511 VCC.n433 0.152939
R1090 VCC.n257 VCC.n256 0.152939
R1091 VCC.n258 VCC.n257 0.152939
R1092 VCC.n258 VCC.n157 0.152939
R1093 VCC.n272 VCC.n157 0.152939
R1094 VCC.n273 VCC.n272 0.152939
R1095 VCC.n274 VCC.n273 0.152939
R1096 VCC.n274 VCC.n145 0.152939
R1097 VCC.n288 VCC.n145 0.152939
R1098 VCC.n289 VCC.n288 0.152939
R1099 VCC.n290 VCC.n289 0.152939
R1100 VCC.n290 VCC.n133 0.152939
R1101 VCC.n305 VCC.n133 0.152939
R1102 VCC.n306 VCC.n305 0.152939
R1103 VCC.n307 VCC.n306 0.152939
R1104 VCC.n307 VCC.n122 0.152939
R1105 VCC.n321 VCC.n122 0.152939
R1106 VCC.n322 VCC.n321 0.152939
R1107 VCC.n323 VCC.n322 0.152939
R1108 VCC.n323 VCC.n110 0.152939
R1109 VCC.n337 VCC.n110 0.152939
R1110 VCC.n338 VCC.n337 0.152939
R1111 VCC.n339 VCC.n338 0.152939
R1112 VCC.n339 VCC.n98 0.152939
R1113 VCC.n353 VCC.n98 0.152939
R1114 VCC.n354 VCC.n353 0.152939
R1115 VCC.n355 VCC.n354 0.152939
R1116 VCC.n355 VCC.n1 0.152939
R1117 VCC.n559 VCC.n1 0.13922
R1118 VCC VCC.n0 0.0767195
R1119 VCC VCC.n559 0.063
R1120 VGN.n49 VGN.n48 161.3
R1121 VGN.n47 VGN.n1 161.3
R1122 VGN.n46 VGN.n45 161.3
R1123 VGN.n44 VGN.n2 161.3
R1124 VGN.n43 VGN.n42 161.3
R1125 VGN.n41 VGN.n3 161.3
R1126 VGN.n40 VGN.n39 161.3
R1127 VGN.n38 VGN.n4 161.3
R1128 VGN.n37 VGN.n36 161.3
R1129 VGN.n35 VGN.n5 161.3
R1130 VGN.n34 VGN.n33 161.3
R1131 VGN.n32 VGN.n7 161.3
R1132 VGN.n31 VGN.n30 161.3
R1133 VGN.n29 VGN.n8 161.3
R1134 VGN.n28 VGN.n27 161.3
R1135 VGN.n26 VGN.n9 161.3
R1136 VGN.n25 VGN.n24 161.3
R1137 VGN.n23 VGN.n10 161.3
R1138 VGN.n22 VGN.n21 161.3
R1139 VGN.n20 VGN.n11 161.3
R1140 VGN.n19 VGN.n18 161.3
R1141 VGN.n17 VGN.n12 161.3
R1142 VGN.n16 VGN.n15 161.3
R1143 VGN.n50 VGN.n0 85.0223
R1144 VGN.n14 VGN.n13 59.6012
R1145 VGN.n42 VGN.n2 56.4773
R1146 VGN.n22 VGN.n11 50.148
R1147 VGN.n30 VGN.n7 50.148
R1148 VGN.n14 VGN.t2 39.14
R1149 VGN.n18 VGN.n11 30.6732
R1150 VGN.n34 VGN.n7 30.6732
R1151 VGN.n18 VGN.n17 24.3439
R1152 VGN.n17 VGN.n16 24.3439
R1153 VGN.n30 VGN.n29 24.3439
R1154 VGN.n29 VGN.n28 24.3439
R1155 VGN.n28 VGN.n9 24.3439
R1156 VGN.n24 VGN.n9 24.3439
R1157 VGN.n24 VGN.n23 24.3439
R1158 VGN.n23 VGN.n22 24.3439
R1159 VGN.n42 VGN.n41 24.3439
R1160 VGN.n41 VGN.n40 24.3439
R1161 VGN.n40 VGN.n4 24.3439
R1162 VGN.n36 VGN.n35 24.3439
R1163 VGN.n35 VGN.n34 24.3439
R1164 VGN.n48 VGN.n47 24.3439
R1165 VGN.n47 VGN.n46 24.3439
R1166 VGN.n46 VGN.n2 24.3439
R1167 VGN.n16 VGN.n13 14.6066
R1168 VGN.n36 VGN.n6 14.6066
R1169 VGN.n6 VGN.n4 9.73787
R1170 VGN.n9 VGN.t3 6.80684
R1171 VGN.n13 VGN.t0 6.80684
R1172 VGN.n6 VGN.t1 6.80684
R1173 VGN.n0 VGN.t4 6.80684
R1174 VGN.n48 VGN.n0 4.86919
R1175 VGN.n15 VGN.n14 3.33651
R1176 VGN.n50 VGN.n49 0.355081
R1177 VGN VGN.n50 0.291472
R1178 VGN.n49 VGN.n1 0.189894
R1179 VGN.n45 VGN.n1 0.189894
R1180 VGN.n45 VGN.n44 0.189894
R1181 VGN.n44 VGN.n43 0.189894
R1182 VGN.n43 VGN.n3 0.189894
R1183 VGN.n39 VGN.n3 0.189894
R1184 VGN.n39 VGN.n38 0.189894
R1185 VGN.n38 VGN.n37 0.189894
R1186 VGN.n37 VGN.n5 0.189894
R1187 VGN.n33 VGN.n5 0.189894
R1188 VGN.n33 VGN.n32 0.189894
R1189 VGN.n32 VGN.n31 0.189894
R1190 VGN.n31 VGN.n8 0.189894
R1191 VGN.n27 VGN.n8 0.189894
R1192 VGN.n27 VGN.n26 0.189894
R1193 VGN.n26 VGN.n25 0.189894
R1194 VGN.n25 VGN.n10 0.189894
R1195 VGN.n21 VGN.n10 0.189894
R1196 VGN.n21 VGN.n20 0.189894
R1197 VGN.n20 VGN.n19 0.189894
R1198 VGN.n19 VGN.n12 0.189894
R1199 VGN.n15 VGN.n12 0.189894
R1200 VSS.n195 VSS.n168 774.148
R1201 VSS.n422 VSS.n41 774.148
R1202 VSS.n197 VSS.n169 675.086
R1203 VSS.n176 VSS.n167 675.086
R1204 VSS.n421 VSS.n43 675.086
R1205 VSS.n423 VSS.n39 675.086
R1206 VSS.n170 VSS.n169 585
R1207 VSS.n169 VSS.n168 585
R1208 VSS.n202 VSS.n201 585
R1209 VSS.n203 VSS.n202 585
R1210 VSS.n161 VSS.n160 585
R1211 VSS.n162 VSS.n161 585
R1212 VSS.n214 VSS.n213 585
R1213 VSS.n213 VSS.n212 585
R1214 VSS.n158 VSS.n157 585
R1215 VSS.n211 VSS.n157 585
R1216 VSS.n219 VSS.n218 585
R1217 VSS.n220 VSS.n219 585
R1218 VSS.n150 VSS.n149 585
R1219 VSS.n151 VSS.n150 585
R1220 VSS.n230 VSS.n229 585
R1221 VSS.n229 VSS.n228 585
R1222 VSS.n147 VSS.n146 585
R1223 VSS.n146 VSS.n145 585
R1224 VSS.n235 VSS.n234 585
R1225 VSS.n236 VSS.n235 585
R1226 VSS.n138 VSS.n137 585
R1227 VSS.n139 VSS.n138 585
R1228 VSS.n246 VSS.n245 585
R1229 VSS.n245 VSS.n244 585
R1230 VSS.n135 VSS.n134 585
R1231 VSS.n134 VSS.n133 585
R1232 VSS.n251 VSS.n250 585
R1233 VSS.n252 VSS.n251 585
R1234 VSS.n126 VSS.n125 585
R1235 VSS.n127 VSS.n126 585
R1236 VSS.n262 VSS.n261 585
R1237 VSS.n261 VSS.n260 585
R1238 VSS.n123 VSS.n122 585
R1239 VSS.n122 VSS.n121 585
R1240 VSS.n267 VSS.n266 585
R1241 VSS.n268 VSS.n267 585
R1242 VSS.n114 VSS.n113 585
R1243 VSS.n115 VSS.n114 585
R1244 VSS.n278 VSS.n277 585
R1245 VSS.n277 VSS.n276 585
R1246 VSS.n111 VSS.n110 585
R1247 VSS.n110 VSS.n109 585
R1248 VSS.n283 VSS.n282 585
R1249 VSS.n284 VSS.n283 585
R1250 VSS.n102 VSS.n101 585
R1251 VSS.n103 VSS.n102 585
R1252 VSS.n294 VSS.n293 585
R1253 VSS.n293 VSS.n292 585
R1254 VSS.n98 VSS.n96 585
R1255 VSS.n96 VSS.n94 585
R1256 VSS.n300 VSS.n299 585
R1257 VSS.n301 VSS.n300 585
R1258 VSS.n99 VSS.n97 585
R1259 VSS.n97 VSS.n95 585
R1260 VSS.n87 VSS.n86 585
R1261 VSS.n88 VSS.n87 585
R1262 VSS.n312 VSS.n311 585
R1263 VSS.n311 VSS.n310 585
R1264 VSS.n84 VSS.n83 585
R1265 VSS.n83 VSS.t1 585
R1266 VSS.n317 VSS.n316 585
R1267 VSS.n318 VSS.n317 585
R1268 VSS.n82 VSS.n81 585
R1269 VSS.n319 VSS.n82 585
R1270 VSS.n323 VSS.n322 585
R1271 VSS.n322 VSS.n321 585
R1272 VSS.n79 VSS.n78 585
R1273 VSS.n78 VSS.n77 585
R1274 VSS.n328 VSS.n327 585
R1275 VSS.n329 VSS.n328 585
R1276 VSS.n76 VSS.n75 585
R1277 VSS.n330 VSS.n76 585
R1278 VSS.n334 VSS.n333 585
R1279 VSS.n333 VSS.n332 585
R1280 VSS.n73 VSS.n72 585
R1281 VSS.n72 VSS.n71 585
R1282 VSS.n339 VSS.n338 585
R1283 VSS.n340 VSS.n339 585
R1284 VSS.n70 VSS.n69 585
R1285 VSS.n341 VSS.n70 585
R1286 VSS.n345 VSS.n344 585
R1287 VSS.n344 VSS.n343 585
R1288 VSS.n67 VSS.n66 585
R1289 VSS.n66 VSS.n65 585
R1290 VSS.n350 VSS.n349 585
R1291 VSS.n351 VSS.n350 585
R1292 VSS.n64 VSS.n63 585
R1293 VSS.n352 VSS.n64 585
R1294 VSS.n356 VSS.n355 585
R1295 VSS.n355 VSS.n354 585
R1296 VSS.n61 VSS.n60 585
R1297 VSS.n60 VSS.n59 585
R1298 VSS.n361 VSS.n360 585
R1299 VSS.n362 VSS.n361 585
R1300 VSS.n58 VSS.n57 585
R1301 VSS.n363 VSS.n58 585
R1302 VSS.n367 VSS.n366 585
R1303 VSS.n366 VSS.n365 585
R1304 VSS.n55 VSS.n54 585
R1305 VSS.n54 VSS.n53 585
R1306 VSS.n372 VSS.n371 585
R1307 VSS.n373 VSS.n372 585
R1308 VSS.n52 VSS.n51 585
R1309 VSS.n374 VSS.n52 585
R1310 VSS.n379 VSS.n378 585
R1311 VSS.n378 VSS.n377 585
R1312 VSS.n49 VSS.n48 585
R1313 VSS.n376 VSS.n48 585
R1314 VSS.n384 VSS.n383 585
R1315 VSS.n385 VSS.n384 585
R1316 VSS.n47 VSS.n46 585
R1317 VSS.n386 VSS.n47 585
R1318 VSS.n390 VSS.n389 585
R1319 VSS.n389 VSS.n388 585
R1320 VSS.n44 VSS.n42 585
R1321 VSS.n42 VSS.n40 585
R1322 VSS.n421 VSS.n420 585
R1323 VSS.n422 VSS.n421 585
R1324 VSS.n424 VSS.n423 585
R1325 VSS.n423 VSS.n422 585
R1326 VSS.n425 VSS.n38 585
R1327 VSS.n40 VSS.n38 585
R1328 VSS.n387 VSS.n36 585
R1329 VSS.n388 VSS.n387 585
R1330 VSS.n429 VSS.n35 585
R1331 VSS.n386 VSS.n35 585
R1332 VSS.n430 VSS.n34 585
R1333 VSS.n385 VSS.n34 585
R1334 VSS.n431 VSS.n33 585
R1335 VSS.n376 VSS.n33 585
R1336 VSS.n375 VSS.n31 585
R1337 VSS.n377 VSS.n375 585
R1338 VSS.n435 VSS.n30 585
R1339 VSS.n374 VSS.n30 585
R1340 VSS.n436 VSS.n29 585
R1341 VSS.n373 VSS.n29 585
R1342 VSS.n437 VSS.n28 585
R1343 VSS.n53 VSS.n28 585
R1344 VSS.n364 VSS.n26 585
R1345 VSS.n365 VSS.n364 585
R1346 VSS.n441 VSS.n25 585
R1347 VSS.n363 VSS.n25 585
R1348 VSS.n442 VSS.n24 585
R1349 VSS.n362 VSS.n24 585
R1350 VSS.n443 VSS.n23 585
R1351 VSS.n59 VSS.n23 585
R1352 VSS.n353 VSS.n21 585
R1353 VSS.n354 VSS.n353 585
R1354 VSS.n447 VSS.n20 585
R1355 VSS.n352 VSS.n20 585
R1356 VSS.n448 VSS.n19 585
R1357 VSS.n351 VSS.n19 585
R1358 VSS.n449 VSS.n18 585
R1359 VSS.n65 VSS.n18 585
R1360 VSS.n342 VSS.n16 585
R1361 VSS.n343 VSS.n342 585
R1362 VSS.n453 VSS.n15 585
R1363 VSS.n341 VSS.n15 585
R1364 VSS.n454 VSS.n14 585
R1365 VSS.n340 VSS.n14 585
R1366 VSS.n455 VSS.n13 585
R1367 VSS.n71 VSS.n13 585
R1368 VSS.n331 VSS.n11 585
R1369 VSS.n332 VSS.n331 585
R1370 VSS.n459 VSS.n10 585
R1371 VSS.n330 VSS.n10 585
R1372 VSS.n460 VSS.n9 585
R1373 VSS.n329 VSS.n9 585
R1374 VSS.n461 VSS.n8 585
R1375 VSS.n77 VSS.n8 585
R1376 VSS.n320 VSS.n6 585
R1377 VSS.n321 VSS.n320 585
R1378 VSS.n465 VSS.n5 585
R1379 VSS.n319 VSS.n5 585
R1380 VSS.n466 VSS.n4 585
R1381 VSS.n318 VSS.n4 585
R1382 VSS.n467 VSS.n3 585
R1383 VSS.t1 VSS.n3 585
R1384 VSS.n309 VSS.n2 585
R1385 VSS.n310 VSS.n309 585
R1386 VSS.n308 VSS.n307 585
R1387 VSS.n308 VSS.n88 585
R1388 VSS.n90 VSS.n89 585
R1389 VSS.n95 VSS.n89 585
R1390 VSS.n303 VSS.n302 585
R1391 VSS.n302 VSS.n301 585
R1392 VSS.n93 VSS.n92 585
R1393 VSS.n94 VSS.n93 585
R1394 VSS.n291 VSS.n290 585
R1395 VSS.n292 VSS.n291 585
R1396 VSS.n105 VSS.n104 585
R1397 VSS.n104 VSS.n103 585
R1398 VSS.n286 VSS.n285 585
R1399 VSS.n285 VSS.n284 585
R1400 VSS.n108 VSS.n107 585
R1401 VSS.n109 VSS.n108 585
R1402 VSS.n275 VSS.n274 585
R1403 VSS.n276 VSS.n275 585
R1404 VSS.n117 VSS.n116 585
R1405 VSS.n116 VSS.n115 585
R1406 VSS.n270 VSS.n269 585
R1407 VSS.n269 VSS.n268 585
R1408 VSS.n120 VSS.n119 585
R1409 VSS.n121 VSS.n120 585
R1410 VSS.n259 VSS.n258 585
R1411 VSS.n260 VSS.n259 585
R1412 VSS.n129 VSS.n128 585
R1413 VSS.n128 VSS.n127 585
R1414 VSS.n254 VSS.n253 585
R1415 VSS.n253 VSS.n252 585
R1416 VSS.n132 VSS.n131 585
R1417 VSS.n133 VSS.n132 585
R1418 VSS.n243 VSS.n242 585
R1419 VSS.n244 VSS.n243 585
R1420 VSS.n141 VSS.n140 585
R1421 VSS.n140 VSS.n139 585
R1422 VSS.n238 VSS.n237 585
R1423 VSS.n237 VSS.n236 585
R1424 VSS.n144 VSS.n143 585
R1425 VSS.n145 VSS.n144 585
R1426 VSS.n227 VSS.n226 585
R1427 VSS.n228 VSS.n227 585
R1428 VSS.n153 VSS.n152 585
R1429 VSS.n152 VSS.n151 585
R1430 VSS.n222 VSS.n221 585
R1431 VSS.n221 VSS.n220 585
R1432 VSS.n156 VSS.n155 585
R1433 VSS.n211 VSS.n156 585
R1434 VSS.n210 VSS.n209 585
R1435 VSS.n212 VSS.n210 585
R1436 VSS.n164 VSS.n163 585
R1437 VSS.n163 VSS.n162 585
R1438 VSS.n205 VSS.n204 585
R1439 VSS.n204 VSS.n203 585
R1440 VSS.n167 VSS.n166 585
R1441 VSS.n168 VSS.n167 585
R1442 VSS.n403 VSS.n39 585
R1443 VSS.n404 VSS.n399 585
R1444 VSS.n406 VSS.n405 585
R1445 VSS.n408 VSS.n396 585
R1446 VSS.n410 VSS.n409 585
R1447 VSS.n411 VSS.n395 585
R1448 VSS.n413 VSS.n412 585
R1449 VSS.n415 VSS.n393 585
R1450 VSS.n417 VSS.n416 585
R1451 VSS.n418 VSS.n43 585
R1452 VSS.n198 VSS.n197 585
R1453 VSS.n172 VSS.n171 585
R1454 VSS.n194 VSS.n193 585
R1455 VSS.n195 VSS.n194 585
R1456 VSS.n192 VSS.n177 585
R1457 VSS.n191 VSS.n190 585
R1458 VSS.n189 VSS.n188 585
R1459 VSS.n187 VSS.n186 585
R1460 VSS.n185 VSS.n184 585
R1461 VSS.n183 VSS.n182 585
R1462 VSS.n181 VSS.n176 585
R1463 VSS.n195 VSS.n176 585
R1464 VSS.n203 VSS.n168 394.974
R1465 VSS.n203 VSS.n162 394.974
R1466 VSS.n212 VSS.n162 394.974
R1467 VSS.n212 VSS.n211 394.974
R1468 VSS.n220 VSS.n151 394.974
R1469 VSS.n228 VSS.n151 394.974
R1470 VSS.n228 VSS.n145 394.974
R1471 VSS.n236 VSS.n145 394.974
R1472 VSS.n236 VSS.n139 394.974
R1473 VSS.n244 VSS.n139 394.974
R1474 VSS.n244 VSS.n133 394.974
R1475 VSS.n252 VSS.n133 394.974
R1476 VSS.n260 VSS.n127 394.974
R1477 VSS.n260 VSS.n121 394.974
R1478 VSS.n268 VSS.n121 394.974
R1479 VSS.n268 VSS.n115 394.974
R1480 VSS.n276 VSS.n115 394.974
R1481 VSS.n276 VSS.n109 394.974
R1482 VSS.n284 VSS.n109 394.974
R1483 VSS.n292 VSS.n103 394.974
R1484 VSS.n292 VSS.n94 394.974
R1485 VSS.n301 VSS.n94 394.974
R1486 VSS.n301 VSS.n95 394.974
R1487 VSS.n95 VSS.n88 394.974
R1488 VSS.n310 VSS.n88 394.974
R1489 VSS.n310 VSS.t1 394.974
R1490 VSS.n318 VSS.t1 394.974
R1491 VSS.n319 VSS.n318 394.974
R1492 VSS.n321 VSS.n319 394.974
R1493 VSS.n321 VSS.n77 394.974
R1494 VSS.n329 VSS.n77 394.974
R1495 VSS.n330 VSS.n329 394.974
R1496 VSS.n332 VSS.n330 394.974
R1497 VSS.n340 VSS.n71 394.974
R1498 VSS.n341 VSS.n340 394.974
R1499 VSS.n343 VSS.n341 394.974
R1500 VSS.n343 VSS.n65 394.974
R1501 VSS.n351 VSS.n65 394.974
R1502 VSS.n352 VSS.n351 394.974
R1503 VSS.n354 VSS.n352 394.974
R1504 VSS.n362 VSS.n59 394.974
R1505 VSS.n363 VSS.n362 394.974
R1506 VSS.n365 VSS.n363 394.974
R1507 VSS.n365 VSS.n53 394.974
R1508 VSS.n373 VSS.n53 394.974
R1509 VSS.n374 VSS.n373 394.974
R1510 VSS.n377 VSS.n374 394.974
R1511 VSS.n377 VSS.n376 394.974
R1512 VSS.n386 VSS.n385 394.974
R1513 VSS.n388 VSS.n386 394.974
R1514 VSS.n388 VSS.n40 394.974
R1515 VSS.n422 VSS.n40 394.974
R1516 VSS.n220 VSS.t6 387.075
R1517 VSS.n376 VSS.t10 387.075
R1518 VSS.n252 VSS.t0 315.978
R1519 VSS.t2 VSS.n59 315.978
R1520 VSS.n400 VSS.t11 307.604
R1521 VSS.n178 VSS.t8 307.604
R1522 VSS.n398 VSS.n41 256.663
R1523 VSS.n407 VSS.n41 256.663
R1524 VSS.n397 VSS.n41 256.663
R1525 VSS.n414 VSS.n41 256.663
R1526 VSS.n394 VSS.n41 256.663
R1527 VSS.n196 VSS.n195 256.663
R1528 VSS.n195 VSS.n173 256.663
R1529 VSS.n195 VSS.n174 256.663
R1530 VSS.n195 VSS.n175 256.663
R1531 VSS.n202 VSS.n169 240.244
R1532 VSS.n202 VSS.n161 240.244
R1533 VSS.n213 VSS.n161 240.244
R1534 VSS.n213 VSS.n157 240.244
R1535 VSS.n219 VSS.n157 240.244
R1536 VSS.n219 VSS.n150 240.244
R1537 VSS.n229 VSS.n150 240.244
R1538 VSS.n229 VSS.n146 240.244
R1539 VSS.n235 VSS.n146 240.244
R1540 VSS.n235 VSS.n138 240.244
R1541 VSS.n245 VSS.n138 240.244
R1542 VSS.n245 VSS.n134 240.244
R1543 VSS.n251 VSS.n134 240.244
R1544 VSS.n251 VSS.n126 240.244
R1545 VSS.n261 VSS.n126 240.244
R1546 VSS.n261 VSS.n122 240.244
R1547 VSS.n267 VSS.n122 240.244
R1548 VSS.n267 VSS.n114 240.244
R1549 VSS.n277 VSS.n114 240.244
R1550 VSS.n277 VSS.n110 240.244
R1551 VSS.n283 VSS.n110 240.244
R1552 VSS.n283 VSS.n102 240.244
R1553 VSS.n293 VSS.n102 240.244
R1554 VSS.n293 VSS.n96 240.244
R1555 VSS.n300 VSS.n96 240.244
R1556 VSS.n300 VSS.n97 240.244
R1557 VSS.n97 VSS.n87 240.244
R1558 VSS.n311 VSS.n87 240.244
R1559 VSS.n311 VSS.n83 240.244
R1560 VSS.n317 VSS.n83 240.244
R1561 VSS.n317 VSS.n82 240.244
R1562 VSS.n322 VSS.n82 240.244
R1563 VSS.n322 VSS.n78 240.244
R1564 VSS.n328 VSS.n78 240.244
R1565 VSS.n328 VSS.n76 240.244
R1566 VSS.n333 VSS.n76 240.244
R1567 VSS.n333 VSS.n72 240.244
R1568 VSS.n339 VSS.n72 240.244
R1569 VSS.n339 VSS.n70 240.244
R1570 VSS.n344 VSS.n70 240.244
R1571 VSS.n344 VSS.n66 240.244
R1572 VSS.n350 VSS.n66 240.244
R1573 VSS.n350 VSS.n64 240.244
R1574 VSS.n355 VSS.n64 240.244
R1575 VSS.n355 VSS.n60 240.244
R1576 VSS.n361 VSS.n60 240.244
R1577 VSS.n361 VSS.n58 240.244
R1578 VSS.n366 VSS.n58 240.244
R1579 VSS.n366 VSS.n54 240.244
R1580 VSS.n372 VSS.n54 240.244
R1581 VSS.n372 VSS.n52 240.244
R1582 VSS.n378 VSS.n52 240.244
R1583 VSS.n378 VSS.n48 240.244
R1584 VSS.n384 VSS.n48 240.244
R1585 VSS.n384 VSS.n47 240.244
R1586 VSS.n389 VSS.n47 240.244
R1587 VSS.n389 VSS.n42 240.244
R1588 VSS.n421 VSS.n42 240.244
R1589 VSS.n204 VSS.n167 240.244
R1590 VSS.n204 VSS.n163 240.244
R1591 VSS.n210 VSS.n163 240.244
R1592 VSS.n210 VSS.n156 240.244
R1593 VSS.n221 VSS.n156 240.244
R1594 VSS.n221 VSS.n152 240.244
R1595 VSS.n227 VSS.n152 240.244
R1596 VSS.n227 VSS.n144 240.244
R1597 VSS.n237 VSS.n144 240.244
R1598 VSS.n237 VSS.n140 240.244
R1599 VSS.n243 VSS.n140 240.244
R1600 VSS.n243 VSS.n132 240.244
R1601 VSS.n253 VSS.n132 240.244
R1602 VSS.n253 VSS.n128 240.244
R1603 VSS.n259 VSS.n128 240.244
R1604 VSS.n259 VSS.n120 240.244
R1605 VSS.n269 VSS.n120 240.244
R1606 VSS.n269 VSS.n116 240.244
R1607 VSS.n275 VSS.n116 240.244
R1608 VSS.n275 VSS.n108 240.244
R1609 VSS.n285 VSS.n108 240.244
R1610 VSS.n285 VSS.n104 240.244
R1611 VSS.n291 VSS.n104 240.244
R1612 VSS.n291 VSS.n93 240.244
R1613 VSS.n302 VSS.n93 240.244
R1614 VSS.n302 VSS.n89 240.244
R1615 VSS.n308 VSS.n89 240.244
R1616 VSS.n309 VSS.n308 240.244
R1617 VSS.n309 VSS.n3 240.244
R1618 VSS.n4 VSS.n3 240.244
R1619 VSS.n5 VSS.n4 240.244
R1620 VSS.n320 VSS.n5 240.244
R1621 VSS.n320 VSS.n8 240.244
R1622 VSS.n9 VSS.n8 240.244
R1623 VSS.n10 VSS.n9 240.244
R1624 VSS.n331 VSS.n10 240.244
R1625 VSS.n331 VSS.n13 240.244
R1626 VSS.n14 VSS.n13 240.244
R1627 VSS.n15 VSS.n14 240.244
R1628 VSS.n342 VSS.n15 240.244
R1629 VSS.n342 VSS.n18 240.244
R1630 VSS.n19 VSS.n18 240.244
R1631 VSS.n20 VSS.n19 240.244
R1632 VSS.n353 VSS.n20 240.244
R1633 VSS.n353 VSS.n23 240.244
R1634 VSS.n24 VSS.n23 240.244
R1635 VSS.n25 VSS.n24 240.244
R1636 VSS.n364 VSS.n25 240.244
R1637 VSS.n364 VSS.n28 240.244
R1638 VSS.n29 VSS.n28 240.244
R1639 VSS.n30 VSS.n29 240.244
R1640 VSS.n375 VSS.n30 240.244
R1641 VSS.n375 VSS.n33 240.244
R1642 VSS.n34 VSS.n33 240.244
R1643 VSS.n35 VSS.n34 240.244
R1644 VSS.n387 VSS.n35 240.244
R1645 VSS.n387 VSS.n38 240.244
R1646 VSS.n423 VSS.n38 240.244
R1647 VSS.t3 VSS.n103 236.984
R1648 VSS.n332 VSS.t4 236.984
R1649 VSS.n401 VSS.t12 233.907
R1650 VSS.n179 VSS.t7 233.907
R1651 VSS.n400 VSS.t9 209.774
R1652 VSS.n178 VSS.t5 209.774
R1653 VSS.n194 VSS.n172 163.367
R1654 VSS.n194 VSS.n177 163.367
R1655 VSS.n190 VSS.n189 163.367
R1656 VSS.n186 VSS.n185 163.367
R1657 VSS.n182 VSS.n176 163.367
R1658 VSS.n416 VSS.n415 163.367
R1659 VSS.n413 VSS.n395 163.367
R1660 VSS.n409 VSS.n408 163.367
R1661 VSS.n406 VSS.n399 163.367
R1662 VSS.n284 VSS.t3 157.989
R1663 VSS.t4 VSS.n71 157.989
R1664 VSS.t0 VSS.n127 78.9951
R1665 VSS.n354 VSS.t2 78.9951
R1666 VSS.n401 VSS.n400 73.6975
R1667 VSS.n179 VSS.n178 73.6975
R1668 VSS.n197 VSS.n196 71.676
R1669 VSS.n177 VSS.n173 71.676
R1670 VSS.n189 VSS.n174 71.676
R1671 VSS.n185 VSS.n175 71.676
R1672 VSS.n416 VSS.n394 71.676
R1673 VSS.n414 VSS.n413 71.676
R1674 VSS.n409 VSS.n397 71.676
R1675 VSS.n407 VSS.n406 71.676
R1676 VSS.n398 VSS.n39 71.676
R1677 VSS.n399 VSS.n398 71.676
R1678 VSS.n408 VSS.n407 71.676
R1679 VSS.n397 VSS.n395 71.676
R1680 VSS.n415 VSS.n414 71.676
R1681 VSS.n394 VSS.n43 71.676
R1682 VSS.n196 VSS.n172 71.676
R1683 VSS.n190 VSS.n173 71.676
R1684 VSS.n186 VSS.n174 71.676
R1685 VSS.n182 VSS.n175 71.676
R1686 VSS.n402 VSS.n401 34.3278
R1687 VSS.n180 VSS.n179 34.3278
R1688 VSS.n419 VSS.n418 29.2676
R1689 VSS.n403 VSS.n37 29.2676
R1690 VSS.n199 VSS.n198 29.2676
R1691 VSS.n181 VSS.n165 29.2676
R1692 VSS.n201 VSS.n170 19.3944
R1693 VSS.n201 VSS.n160 19.3944
R1694 VSS.n214 VSS.n160 19.3944
R1695 VSS.n214 VSS.n158 19.3944
R1696 VSS.n218 VSS.n158 19.3944
R1697 VSS.n218 VSS.n149 19.3944
R1698 VSS.n230 VSS.n149 19.3944
R1699 VSS.n230 VSS.n147 19.3944
R1700 VSS.n234 VSS.n147 19.3944
R1701 VSS.n234 VSS.n137 19.3944
R1702 VSS.n246 VSS.n137 19.3944
R1703 VSS.n246 VSS.n135 19.3944
R1704 VSS.n250 VSS.n135 19.3944
R1705 VSS.n250 VSS.n125 19.3944
R1706 VSS.n262 VSS.n125 19.3944
R1707 VSS.n262 VSS.n123 19.3944
R1708 VSS.n266 VSS.n123 19.3944
R1709 VSS.n266 VSS.n113 19.3944
R1710 VSS.n278 VSS.n113 19.3944
R1711 VSS.n278 VSS.n111 19.3944
R1712 VSS.n282 VSS.n111 19.3944
R1713 VSS.n282 VSS.n101 19.3944
R1714 VSS.n294 VSS.n101 19.3944
R1715 VSS.n294 VSS.n98 19.3944
R1716 VSS.n299 VSS.n98 19.3944
R1717 VSS.n299 VSS.n99 19.3944
R1718 VSS.n99 VSS.n86 19.3944
R1719 VSS.n312 VSS.n86 19.3944
R1720 VSS.n312 VSS.n84 19.3944
R1721 VSS.n316 VSS.n84 19.3944
R1722 VSS.n316 VSS.n81 19.3944
R1723 VSS.n323 VSS.n81 19.3944
R1724 VSS.n323 VSS.n79 19.3944
R1725 VSS.n327 VSS.n79 19.3944
R1726 VSS.n327 VSS.n75 19.3944
R1727 VSS.n334 VSS.n75 19.3944
R1728 VSS.n334 VSS.n73 19.3944
R1729 VSS.n338 VSS.n73 19.3944
R1730 VSS.n338 VSS.n69 19.3944
R1731 VSS.n345 VSS.n69 19.3944
R1732 VSS.n345 VSS.n67 19.3944
R1733 VSS.n349 VSS.n67 19.3944
R1734 VSS.n349 VSS.n63 19.3944
R1735 VSS.n356 VSS.n63 19.3944
R1736 VSS.n356 VSS.n61 19.3944
R1737 VSS.n360 VSS.n61 19.3944
R1738 VSS.n360 VSS.n57 19.3944
R1739 VSS.n367 VSS.n57 19.3944
R1740 VSS.n367 VSS.n55 19.3944
R1741 VSS.n371 VSS.n55 19.3944
R1742 VSS.n371 VSS.n51 19.3944
R1743 VSS.n379 VSS.n51 19.3944
R1744 VSS.n379 VSS.n49 19.3944
R1745 VSS.n383 VSS.n49 19.3944
R1746 VSS.n383 VSS.n46 19.3944
R1747 VSS.n390 VSS.n46 19.3944
R1748 VSS.n390 VSS.n44 19.3944
R1749 VSS.n420 VSS.n44 19.3944
R1750 VSS.n205 VSS.n166 19.3944
R1751 VSS.n205 VSS.n164 19.3944
R1752 VSS.n209 VSS.n164 19.3944
R1753 VSS.n209 VSS.n155 19.3944
R1754 VSS.n222 VSS.n155 19.3944
R1755 VSS.n222 VSS.n153 19.3944
R1756 VSS.n226 VSS.n153 19.3944
R1757 VSS.n226 VSS.n143 19.3944
R1758 VSS.n238 VSS.n143 19.3944
R1759 VSS.n238 VSS.n141 19.3944
R1760 VSS.n242 VSS.n141 19.3944
R1761 VSS.n242 VSS.n131 19.3944
R1762 VSS.n254 VSS.n131 19.3944
R1763 VSS.n254 VSS.n129 19.3944
R1764 VSS.n258 VSS.n129 19.3944
R1765 VSS.n258 VSS.n119 19.3944
R1766 VSS.n270 VSS.n119 19.3944
R1767 VSS.n270 VSS.n117 19.3944
R1768 VSS.n274 VSS.n117 19.3944
R1769 VSS.n274 VSS.n107 19.3944
R1770 VSS.n286 VSS.n107 19.3944
R1771 VSS.n286 VSS.n105 19.3944
R1772 VSS.n290 VSS.n105 19.3944
R1773 VSS.n290 VSS.n92 19.3944
R1774 VSS.n303 VSS.n92 19.3944
R1775 VSS.n303 VSS.n90 19.3944
R1776 VSS.n307 VSS.n90 19.3944
R1777 VSS.n307 VSS.n2 19.3944
R1778 VSS.n467 VSS.n2 19.3944
R1779 VSS.n467 VSS.n466 19.3944
R1780 VSS.n466 VSS.n465 19.3944
R1781 VSS.n465 VSS.n6 19.3944
R1782 VSS.n461 VSS.n6 19.3944
R1783 VSS.n461 VSS.n460 19.3944
R1784 VSS.n460 VSS.n459 19.3944
R1785 VSS.n459 VSS.n11 19.3944
R1786 VSS.n455 VSS.n11 19.3944
R1787 VSS.n455 VSS.n454 19.3944
R1788 VSS.n454 VSS.n453 19.3944
R1789 VSS.n453 VSS.n16 19.3944
R1790 VSS.n449 VSS.n16 19.3944
R1791 VSS.n449 VSS.n448 19.3944
R1792 VSS.n448 VSS.n447 19.3944
R1793 VSS.n447 VSS.n21 19.3944
R1794 VSS.n443 VSS.n21 19.3944
R1795 VSS.n443 VSS.n442 19.3944
R1796 VSS.n442 VSS.n441 19.3944
R1797 VSS.n441 VSS.n26 19.3944
R1798 VSS.n437 VSS.n26 19.3944
R1799 VSS.n437 VSS.n436 19.3944
R1800 VSS.n436 VSS.n435 19.3944
R1801 VSS.n435 VSS.n31 19.3944
R1802 VSS.n431 VSS.n31 19.3944
R1803 VSS.n431 VSS.n430 19.3944
R1804 VSS.n430 VSS.n429 19.3944
R1805 VSS.n429 VSS.n36 19.3944
R1806 VSS.n425 VSS.n36 19.3944
R1807 VSS.n425 VSS.n424 19.3944
R1808 VSS.n418 VSS.n417 10.6151
R1809 VSS.n417 VSS.n393 10.6151
R1810 VSS.n412 VSS.n393 10.6151
R1811 VSS.n412 VSS.n411 10.6151
R1812 VSS.n411 VSS.n410 10.6151
R1813 VSS.n410 VSS.n396 10.6151
R1814 VSS.n405 VSS.n404 10.6151
R1815 VSS.n404 VSS.n403 10.6151
R1816 VSS.n198 VSS.n171 10.6151
R1817 VSS.n193 VSS.n171 10.6151
R1818 VSS.n193 VSS.n192 10.6151
R1819 VSS.n192 VSS.n191 10.6151
R1820 VSS.n191 VSS.n188 10.6151
R1821 VSS.n188 VSS.n187 10.6151
R1822 VSS.n184 VSS.n183 10.6151
R1823 VSS.n183 VSS.n181 10.6151
R1824 VSS.n402 VSS.n396 10.1468
R1825 VSS.n187 VSS.n180 10.1468
R1826 VSS.n466 VSS.n0 9.3005
R1827 VSS.n465 VSS.n464 9.3005
R1828 VSS.n463 VSS.n6 9.3005
R1829 VSS.n462 VSS.n461 9.3005
R1830 VSS.n460 VSS.n7 9.3005
R1831 VSS.n459 VSS.n458 9.3005
R1832 VSS.n457 VSS.n11 9.3005
R1833 VSS.n456 VSS.n455 9.3005
R1834 VSS.n454 VSS.n12 9.3005
R1835 VSS.n453 VSS.n452 9.3005
R1836 VSS.n451 VSS.n16 9.3005
R1837 VSS.n450 VSS.n449 9.3005
R1838 VSS.n448 VSS.n17 9.3005
R1839 VSS.n447 VSS.n446 9.3005
R1840 VSS.n445 VSS.n21 9.3005
R1841 VSS.n444 VSS.n443 9.3005
R1842 VSS.n442 VSS.n22 9.3005
R1843 VSS.n441 VSS.n440 9.3005
R1844 VSS.n439 VSS.n26 9.3005
R1845 VSS.n438 VSS.n437 9.3005
R1846 VSS.n436 VSS.n27 9.3005
R1847 VSS.n435 VSS.n434 9.3005
R1848 VSS.n433 VSS.n31 9.3005
R1849 VSS.n432 VSS.n431 9.3005
R1850 VSS.n430 VSS.n32 9.3005
R1851 VSS.n429 VSS.n428 9.3005
R1852 VSS.n427 VSS.n36 9.3005
R1853 VSS.n426 VSS.n425 9.3005
R1854 VSS.n424 VSS.n37 9.3005
R1855 VSS.n199 VSS.n170 9.3005
R1856 VSS.n201 VSS.n200 9.3005
R1857 VSS.n160 VSS.n159 9.3005
R1858 VSS.n215 VSS.n214 9.3005
R1859 VSS.n216 VSS.n158 9.3005
R1860 VSS.n218 VSS.n217 9.3005
R1861 VSS.n149 VSS.n148 9.3005
R1862 VSS.n231 VSS.n230 9.3005
R1863 VSS.n232 VSS.n147 9.3005
R1864 VSS.n234 VSS.n233 9.3005
R1865 VSS.n137 VSS.n136 9.3005
R1866 VSS.n247 VSS.n246 9.3005
R1867 VSS.n248 VSS.n135 9.3005
R1868 VSS.n250 VSS.n249 9.3005
R1869 VSS.n125 VSS.n124 9.3005
R1870 VSS.n263 VSS.n262 9.3005
R1871 VSS.n264 VSS.n123 9.3005
R1872 VSS.n266 VSS.n265 9.3005
R1873 VSS.n113 VSS.n112 9.3005
R1874 VSS.n279 VSS.n278 9.3005
R1875 VSS.n280 VSS.n111 9.3005
R1876 VSS.n282 VSS.n281 9.3005
R1877 VSS.n101 VSS.n100 9.3005
R1878 VSS.n295 VSS.n294 9.3005
R1879 VSS.n296 VSS.n98 9.3005
R1880 VSS.n299 VSS.n298 9.3005
R1881 VSS.n297 VSS.n99 9.3005
R1882 VSS.n86 VSS.n85 9.3005
R1883 VSS.n313 VSS.n312 9.3005
R1884 VSS.n314 VSS.n84 9.3005
R1885 VSS.n316 VSS.n315 9.3005
R1886 VSS.n81 VSS.n80 9.3005
R1887 VSS.n324 VSS.n323 9.3005
R1888 VSS.n325 VSS.n79 9.3005
R1889 VSS.n327 VSS.n326 9.3005
R1890 VSS.n75 VSS.n74 9.3005
R1891 VSS.n335 VSS.n334 9.3005
R1892 VSS.n336 VSS.n73 9.3005
R1893 VSS.n338 VSS.n337 9.3005
R1894 VSS.n69 VSS.n68 9.3005
R1895 VSS.n346 VSS.n345 9.3005
R1896 VSS.n347 VSS.n67 9.3005
R1897 VSS.n349 VSS.n348 9.3005
R1898 VSS.n63 VSS.n62 9.3005
R1899 VSS.n357 VSS.n356 9.3005
R1900 VSS.n358 VSS.n61 9.3005
R1901 VSS.n360 VSS.n359 9.3005
R1902 VSS.n57 VSS.n56 9.3005
R1903 VSS.n368 VSS.n367 9.3005
R1904 VSS.n369 VSS.n55 9.3005
R1905 VSS.n371 VSS.n370 9.3005
R1906 VSS.n51 VSS.n50 9.3005
R1907 VSS.n380 VSS.n379 9.3005
R1908 VSS.n381 VSS.n49 9.3005
R1909 VSS.n383 VSS.n382 9.3005
R1910 VSS.n46 VSS.n45 9.3005
R1911 VSS.n391 VSS.n390 9.3005
R1912 VSS.n392 VSS.n44 9.3005
R1913 VSS.n420 VSS.n419 9.3005
R1914 VSS.n206 VSS.n205 9.3005
R1915 VSS.n207 VSS.n164 9.3005
R1916 VSS.n209 VSS.n208 9.3005
R1917 VSS.n155 VSS.n154 9.3005
R1918 VSS.n223 VSS.n222 9.3005
R1919 VSS.n224 VSS.n153 9.3005
R1920 VSS.n226 VSS.n225 9.3005
R1921 VSS.n143 VSS.n142 9.3005
R1922 VSS.n239 VSS.n238 9.3005
R1923 VSS.n240 VSS.n141 9.3005
R1924 VSS.n242 VSS.n241 9.3005
R1925 VSS.n131 VSS.n130 9.3005
R1926 VSS.n255 VSS.n254 9.3005
R1927 VSS.n256 VSS.n129 9.3005
R1928 VSS.n258 VSS.n257 9.3005
R1929 VSS.n119 VSS.n118 9.3005
R1930 VSS.n271 VSS.n270 9.3005
R1931 VSS.n272 VSS.n117 9.3005
R1932 VSS.n274 VSS.n273 9.3005
R1933 VSS.n107 VSS.n106 9.3005
R1934 VSS.n287 VSS.n286 9.3005
R1935 VSS.n288 VSS.n105 9.3005
R1936 VSS.n290 VSS.n289 9.3005
R1937 VSS.n92 VSS.n91 9.3005
R1938 VSS.n304 VSS.n303 9.3005
R1939 VSS.n305 VSS.n90 9.3005
R1940 VSS.n307 VSS.n306 9.3005
R1941 VSS.n2 VSS.n1 9.3005
R1942 VSS.n166 VSS.n165 9.3005
R1943 VSS.n468 VSS.n467 9.3005
R1944 VSS.n211 VSS.t6 7.89996
R1945 VSS.n385 VSS.t10 7.89996
R1946 VSS.n405 VSS.n402 0.468793
R1947 VSS.n184 VSS.n180 0.468793
R1948 VSS.n464 VSS.n0 0.152939
R1949 VSS.n464 VSS.n463 0.152939
R1950 VSS.n463 VSS.n462 0.152939
R1951 VSS.n462 VSS.n7 0.152939
R1952 VSS.n458 VSS.n7 0.152939
R1953 VSS.n458 VSS.n457 0.152939
R1954 VSS.n457 VSS.n456 0.152939
R1955 VSS.n456 VSS.n12 0.152939
R1956 VSS.n452 VSS.n12 0.152939
R1957 VSS.n452 VSS.n451 0.152939
R1958 VSS.n451 VSS.n450 0.152939
R1959 VSS.n450 VSS.n17 0.152939
R1960 VSS.n446 VSS.n17 0.152939
R1961 VSS.n446 VSS.n445 0.152939
R1962 VSS.n445 VSS.n444 0.152939
R1963 VSS.n444 VSS.n22 0.152939
R1964 VSS.n440 VSS.n22 0.152939
R1965 VSS.n440 VSS.n439 0.152939
R1966 VSS.n439 VSS.n438 0.152939
R1967 VSS.n438 VSS.n27 0.152939
R1968 VSS.n434 VSS.n27 0.152939
R1969 VSS.n434 VSS.n433 0.152939
R1970 VSS.n433 VSS.n432 0.152939
R1971 VSS.n432 VSS.n32 0.152939
R1972 VSS.n428 VSS.n32 0.152939
R1973 VSS.n428 VSS.n427 0.152939
R1974 VSS.n427 VSS.n426 0.152939
R1975 VSS.n426 VSS.n37 0.152939
R1976 VSS.n200 VSS.n199 0.152939
R1977 VSS.n200 VSS.n159 0.152939
R1978 VSS.n215 VSS.n159 0.152939
R1979 VSS.n216 VSS.n215 0.152939
R1980 VSS.n217 VSS.n216 0.152939
R1981 VSS.n217 VSS.n148 0.152939
R1982 VSS.n231 VSS.n148 0.152939
R1983 VSS.n232 VSS.n231 0.152939
R1984 VSS.n233 VSS.n232 0.152939
R1985 VSS.n233 VSS.n136 0.152939
R1986 VSS.n247 VSS.n136 0.152939
R1987 VSS.n248 VSS.n247 0.152939
R1988 VSS.n249 VSS.n248 0.152939
R1989 VSS.n249 VSS.n124 0.152939
R1990 VSS.n263 VSS.n124 0.152939
R1991 VSS.n264 VSS.n263 0.152939
R1992 VSS.n265 VSS.n264 0.152939
R1993 VSS.n265 VSS.n112 0.152939
R1994 VSS.n279 VSS.n112 0.152939
R1995 VSS.n280 VSS.n279 0.152939
R1996 VSS.n281 VSS.n280 0.152939
R1997 VSS.n281 VSS.n100 0.152939
R1998 VSS.n295 VSS.n100 0.152939
R1999 VSS.n296 VSS.n295 0.152939
R2000 VSS.n298 VSS.n296 0.152939
R2001 VSS.n298 VSS.n297 0.152939
R2002 VSS.n297 VSS.n85 0.152939
R2003 VSS.n313 VSS.n85 0.152939
R2004 VSS.n314 VSS.n313 0.152939
R2005 VSS.n315 VSS.n314 0.152939
R2006 VSS.n315 VSS.n80 0.152939
R2007 VSS.n324 VSS.n80 0.152939
R2008 VSS.n325 VSS.n324 0.152939
R2009 VSS.n326 VSS.n325 0.152939
R2010 VSS.n326 VSS.n74 0.152939
R2011 VSS.n335 VSS.n74 0.152939
R2012 VSS.n336 VSS.n335 0.152939
R2013 VSS.n337 VSS.n336 0.152939
R2014 VSS.n337 VSS.n68 0.152939
R2015 VSS.n346 VSS.n68 0.152939
R2016 VSS.n347 VSS.n346 0.152939
R2017 VSS.n348 VSS.n347 0.152939
R2018 VSS.n348 VSS.n62 0.152939
R2019 VSS.n357 VSS.n62 0.152939
R2020 VSS.n358 VSS.n357 0.152939
R2021 VSS.n359 VSS.n358 0.152939
R2022 VSS.n359 VSS.n56 0.152939
R2023 VSS.n368 VSS.n56 0.152939
R2024 VSS.n369 VSS.n368 0.152939
R2025 VSS.n370 VSS.n369 0.152939
R2026 VSS.n370 VSS.n50 0.152939
R2027 VSS.n380 VSS.n50 0.152939
R2028 VSS.n381 VSS.n380 0.152939
R2029 VSS.n382 VSS.n381 0.152939
R2030 VSS.n382 VSS.n45 0.152939
R2031 VSS.n391 VSS.n45 0.152939
R2032 VSS.n392 VSS.n391 0.152939
R2033 VSS.n419 VSS.n392 0.152939
R2034 VSS.n206 VSS.n165 0.152939
R2035 VSS.n207 VSS.n206 0.152939
R2036 VSS.n208 VSS.n207 0.152939
R2037 VSS.n208 VSS.n154 0.152939
R2038 VSS.n223 VSS.n154 0.152939
R2039 VSS.n224 VSS.n223 0.152939
R2040 VSS.n225 VSS.n224 0.152939
R2041 VSS.n225 VSS.n142 0.152939
R2042 VSS.n239 VSS.n142 0.152939
R2043 VSS.n240 VSS.n239 0.152939
R2044 VSS.n241 VSS.n240 0.152939
R2045 VSS.n241 VSS.n130 0.152939
R2046 VSS.n255 VSS.n130 0.152939
R2047 VSS.n256 VSS.n255 0.152939
R2048 VSS.n257 VSS.n256 0.152939
R2049 VSS.n257 VSS.n118 0.152939
R2050 VSS.n271 VSS.n118 0.152939
R2051 VSS.n272 VSS.n271 0.152939
R2052 VSS.n273 VSS.n272 0.152939
R2053 VSS.n273 VSS.n106 0.152939
R2054 VSS.n287 VSS.n106 0.152939
R2055 VSS.n288 VSS.n287 0.152939
R2056 VSS.n289 VSS.n288 0.152939
R2057 VSS.n289 VSS.n91 0.152939
R2058 VSS.n304 VSS.n91 0.152939
R2059 VSS.n305 VSS.n304 0.152939
R2060 VSS.n306 VSS.n305 0.152939
R2061 VSS.n306 VSS.n1 0.152939
R2062 VSS.n468 VSS.n1 0.13922
R2063 VSS VSS.n0 0.0767195
R2064 VSS VSS.n468 0.063
C0 VGP VIN 4.4489f
C1 VGP VOUT 3.67101f
C2 VOUT VIN 5.67954f
C3 VGP VGN 0.066133f
C4 VGN VIN 1.56112f
C5 VGN VOUT 0.587269f
C6 VCC VGP 6.66074f
C7 VCC VIN 1.24824f
C8 VCC VOUT 2.82904f
C9 VCC VGN 0.06632f
C10 VGN VSS 8.85494f
C11 VOUT VSS 2.775231f
C12 VIN VSS 1.440425f
C13 VGP VSS 2.395531f
C14 VCC VSS 50.339638f
C15 VCC.n0 VSS 0.002624f
C16 VCC.n1 VSS 0.003499f
C17 VCC.n2 VSS 0.002817f
C18 VCC.n3 VSS 0.003499f
C19 VCC.n4 VSS 0.003499f
C20 VCC.n5 VSS 0.003499f
C21 VCC.n6 VSS 0.002817f
C22 VCC.n7 VSS 0.003499f
C23 VCC.n8 VSS 0.003499f
C24 VCC.n9 VSS 0.003499f
C25 VCC.n10 VSS 0.003499f
C26 VCC.n11 VSS 0.002817f
C27 VCC.n12 VSS 0.003499f
C28 VCC.n13 VSS 0.003499f
C29 VCC.n14 VSS 0.003499f
C30 VCC.n15 VSS 0.003499f
C31 VCC.n16 VSS 0.002817f
C32 VCC.n17 VSS 0.003499f
C33 VCC.n18 VSS 0.003499f
C34 VCC.n19 VSS 0.003499f
C35 VCC.n20 VSS 0.003499f
C36 VCC.n21 VSS 0.002817f
C37 VCC.n22 VSS 0.003499f
C38 VCC.n23 VSS 0.003499f
C39 VCC.n24 VSS 0.003499f
C40 VCC.n25 VSS 0.003499f
C41 VCC.n26 VSS 0.002817f
C42 VCC.n27 VSS 0.003499f
C43 VCC.n28 VSS 0.003499f
C44 VCC.n29 VSS 0.003499f
C45 VCC.n30 VSS 0.003499f
C46 VCC.n31 VSS 0.002817f
C47 VCC.n32 VSS 0.003499f
C48 VCC.n33 VSS 0.003499f
C49 VCC.n34 VSS 0.003499f
C50 VCC.n35 VSS 0.003499f
C51 VCC.n36 VSS 0.002817f
C52 VCC.n37 VSS 0.004662f
C53 VCC.n38 VSS 0.003499f
C54 VCC.n39 VSS 0.006809f
C55 VCC.n40 VSS 0.106772f
C56 VCC.n41 VSS 0.205536f
C57 VCC.n42 VSS 0.003499f
C58 VCC.n43 VSS 0.006809f
C59 VCC.n44 VSS 0.002817f
C60 VCC.n45 VSS 0.003499f
C61 VCC.n46 VSS 0.002817f
C62 VCC.n47 VSS 0.003499f
C63 VCC.n48 VSS 0.003499f
C64 VCC.n49 VSS 0.106772f
C65 VCC.n50 VSS 0.003499f
C66 VCC.n51 VSS 0.002817f
C67 VCC.n52 VSS 0.003499f
C68 VCC.n53 VSS 0.002817f
C69 VCC.n54 VSS 0.003499f
C70 VCC.n55 VSS 0.003499f
C71 VCC.n56 VSS 0.106772f
C72 VCC.n57 VSS 0.003499f
C73 VCC.n58 VSS 0.002817f
C74 VCC.n59 VSS 0.003499f
C75 VCC.n60 VSS 0.002817f
C76 VCC.n61 VSS 0.003499f
C77 VCC.n62 VSS 0.003499f
C78 VCC.n63 VSS 0.070469f
C79 VCC.n64 VSS 0.003499f
C80 VCC.n65 VSS 0.002817f
C81 VCC.n66 VSS 0.003499f
C82 VCC.n67 VSS 0.002817f
C83 VCC.n68 VSS 0.003499f
C84 VCC.n69 VSS 0.003499f
C85 VCC.n70 VSS 0.106772f
C86 VCC.n71 VSS 0.003499f
C87 VCC.n72 VSS 0.002817f
C88 VCC.n73 VSS 0.003499f
C89 VCC.n74 VSS 0.002817f
C90 VCC.n75 VSS 0.003499f
C91 VCC.t1 VSS 0.053386f
C92 VCC.n76 VSS 0.003499f
C93 VCC.n77 VSS 0.002817f
C94 VCC.n78 VSS 0.003499f
C95 VCC.n79 VSS 0.002817f
C96 VCC.n80 VSS 0.003499f
C97 VCC.n81 VSS 0.003499f
C98 VCC.n82 VSS 0.106772f
C99 VCC.n83 VSS 0.003499f
C100 VCC.n84 VSS 0.002817f
C101 VCC.n85 VSS 0.003499f
C102 VCC.n86 VSS 0.002817f
C103 VCC.n87 VSS 0.003499f
C104 VCC.n88 VSS 0.106772f
C105 VCC.n89 VSS 0.003499f
C106 VCC.n90 VSS 0.002817f
C107 VCC.n91 VSS 0.003499f
C108 VCC.n92 VSS 0.002817f
C109 VCC.n93 VSS 0.003499f
C110 VCC.n94 VSS 0.106772f
C111 VCC.n95 VSS 0.003499f
C112 VCC.n96 VSS 0.003499f
C113 VCC.n97 VSS 0.002817f
C114 VCC.n98 VSS 0.003499f
C115 VCC.n99 VSS 0.002817f
C116 VCC.n100 VSS 0.003499f
C117 VCC.n101 VSS 0.106772f
C118 VCC.n102 VSS 0.003499f
C119 VCC.n103 VSS 0.002817f
C120 VCC.n104 VSS 0.003499f
C121 VCC.n105 VSS 0.002817f
C122 VCC.n106 VSS 0.003499f
C123 VCC.n107 VSS 0.071537f
C124 VCC.n108 VSS 0.003499f
C125 VCC.n109 VSS 0.002817f
C126 VCC.n110 VSS 0.003499f
C127 VCC.n111 VSS 0.002817f
C128 VCC.n112 VSS 0.003499f
C129 VCC.n113 VSS 0.106772f
C130 VCC.n114 VSS 0.003499f
C131 VCC.n115 VSS 0.002817f
C132 VCC.n116 VSS 0.003499f
C133 VCC.n117 VSS 0.002817f
C134 VCC.n118 VSS 0.003499f
C135 VCC.n119 VSS 0.106772f
C136 VCC.n120 VSS 0.003499f
C137 VCC.n121 VSS 0.002817f
C138 VCC.n122 VSS 0.003499f
C139 VCC.n123 VSS 0.002817f
C140 VCC.n124 VSS 0.003499f
C141 VCC.n125 VSS 0.106772f
C142 VCC.n126 VSS 0.003499f
C143 VCC.n127 VSS 0.002817f
C144 VCC.n128 VSS 0.003499f
C145 VCC.n129 VSS 0.002817f
C146 VCC.n130 VSS 0.003499f
C147 VCC.t3 VSS 0.053386f
C148 VCC.n131 VSS 0.003499f
C149 VCC.n132 VSS 0.002817f
C150 VCC.n133 VSS 0.003499f
C151 VCC.n134 VSS 0.002817f
C152 VCC.n135 VSS 0.003499f
C153 VCC.n136 VSS 0.106772f
C154 VCC.n137 VSS 0.003499f
C155 VCC.n138 VSS 0.002817f
C156 VCC.n139 VSS 0.003499f
C157 VCC.n140 VSS 0.002817f
C158 VCC.n141 VSS 0.003499f
C159 VCC.n142 VSS 0.106772f
C160 VCC.n143 VSS 0.003499f
C161 VCC.n144 VSS 0.002817f
C162 VCC.n145 VSS 0.003499f
C163 VCC.n146 VSS 0.002817f
C164 VCC.n147 VSS 0.003499f
C165 VCC.n148 VSS 0.106772f
C166 VCC.n149 VSS 0.003499f
C167 VCC.n150 VSS 0.002817f
C168 VCC.n151 VSS 0.003499f
C169 VCC.n152 VSS 0.002817f
C170 VCC.n153 VSS 0.003499f
C171 VCC.n154 VSS 0.106772f
C172 VCC.n155 VSS 0.003499f
C173 VCC.n156 VSS 0.002817f
C174 VCC.n157 VSS 0.003499f
C175 VCC.n158 VSS 0.002817f
C176 VCC.n159 VSS 0.003499f
C177 VCC.t6 VSS 0.053386f
C178 VCC.n160 VSS 0.003499f
C179 VCC.n161 VSS 0.002817f
C180 VCC.n162 VSS 0.003499f
C181 VCC.n163 VSS 0.002817f
C182 VCC.n164 VSS 0.003499f
C183 VCC.n165 VSS 0.106772f
C184 VCC.n166 VSS 0.096095f
C185 VCC.n167 VSS 0.003499f
C186 VCC.n168 VSS 0.002817f
C187 VCC.n169 VSS 0.004662f
C188 VCC.n170 VSS 0.006809f
C189 VCC.n171 VSS 0.205536f
C190 VCC.n172 VSS 0.006809f
C191 VCC.n173 VSS 0.00238f
C192 VCC.n174 VSS 0.00238f
C193 VCC.n175 VSS 0.00238f
C194 VCC.n176 VSS 0.00238f
C195 VCC.n177 VSS 0.00238f
C196 VCC.n178 VSS 0.00238f
C197 VCC.n179 VSS 0.00238f
C198 VCC.n180 VSS 0.00238f
C199 VCC.n181 VSS 0.00238f
C200 VCC.n182 VSS 0.00238f
C201 VCC.n183 VSS 0.00238f
C202 VCC.n184 VSS 0.00238f
C203 VCC.n185 VSS 0.00238f
C204 VCC.n186 VSS 0.00238f
C205 VCC.t7 VSS 0.088796f
C206 VCC.t8 VSS 0.097274f
C207 VCC.t5 VSS 0.44962f
C208 VCC.n187 VSS 0.054957f
C209 VCC.n188 VSS 0.023145f
C210 VCC.n190 VSS 0.00238f
C211 VCC.n191 VSS 0.001942f
C212 VCC.n192 VSS 0.003316f
C213 VCC.n193 VSS 0.001627f
C214 VCC.n194 VSS 0.00238f
C215 VCC.n195 VSS 0.00238f
C216 VCC.n197 VSS 0.00238f
C217 VCC.n199 VSS 0.00238f
C218 VCC.n200 VSS 0.00238f
C219 VCC.n201 VSS 0.00238f
C220 VCC.n202 VSS 0.00238f
C221 VCC.n203 VSS 0.00238f
C222 VCC.n205 VSS 0.00238f
C223 VCC.n207 VSS 0.00238f
C224 VCC.n208 VSS 0.00238f
C225 VCC.n209 VSS 0.00238f
C226 VCC.n210 VSS 0.00238f
C227 VCC.n211 VSS 0.00238f
C228 VCC.n213 VSS 0.00238f
C229 VCC.n215 VSS 0.00238f
C230 VCC.n216 VSS 0.00238f
C231 VCC.n217 VSS 0.00238f
C232 VCC.n218 VSS 0.00238f
C233 VCC.n219 VSS 0.00238f
C234 VCC.n221 VSS 0.00238f
C235 VCC.n223 VSS 0.00238f
C236 VCC.n224 VSS 0.00238f
C237 VCC.n225 VSS 0.00238f
C238 VCC.n226 VSS 0.00238f
C239 VCC.n227 VSS 0.00238f
C240 VCC.n229 VSS 0.00238f
C241 VCC.n231 VSS 0.00238f
C242 VCC.n232 VSS 0.00238f
C243 VCC.n233 VSS 0.00238f
C244 VCC.n234 VSS 0.00238f
C245 VCC.n235 VSS 0.00238f
C246 VCC.n237 VSS 0.00238f
C247 VCC.n239 VSS 0.00238f
C248 VCC.n240 VSS 0.00238f
C249 VCC.n241 VSS 0.00238f
C250 VCC.n242 VSS 0.00238f
C251 VCC.n243 VSS 0.00238f
C252 VCC.n245 VSS 0.00238f
C253 VCC.n247 VSS 0.00238f
C254 VCC.n248 VSS 0.00238f
C255 VCC.n249 VSS 0.004662f
C256 VCC.n250 VSS 0.01189f
C257 VCC.n251 VSS 0.002338f
C258 VCC.n252 VSS 0.006873f
C259 VCC.n253 VSS 0.148947f
C260 VCC.n254 VSS 0.006873f
C261 VCC.n255 VSS 0.002338f
C262 VCC.n256 VSS 0.01189f
C263 VCC.n257 VSS 0.003499f
C264 VCC.n258 VSS 0.003499f
C265 VCC.n259 VSS 0.002817f
C266 VCC.n260 VSS 0.003499f
C267 VCC.n261 VSS 0.106772f
C268 VCC.n262 VSS 0.003499f
C269 VCC.n263 VSS 0.002817f
C270 VCC.n264 VSS 0.003499f
C271 VCC.n265 VSS 0.003499f
C272 VCC.n266 VSS 0.003499f
C273 VCC.n267 VSS 0.002817f
C274 VCC.n268 VSS 0.003499f
C275 VCC.n269 VSS 0.064063f
C276 VCC.n270 VSS 0.003499f
C277 VCC.n271 VSS 0.002817f
C278 VCC.n272 VSS 0.003499f
C279 VCC.n273 VSS 0.003499f
C280 VCC.n274 VSS 0.003499f
C281 VCC.n275 VSS 0.002817f
C282 VCC.n276 VSS 0.003499f
C283 VCC.n277 VSS 0.106772f
C284 VCC.n278 VSS 0.003499f
C285 VCC.n279 VSS 0.002817f
C286 VCC.n280 VSS 0.003499f
C287 VCC.n281 VSS 0.003499f
C288 VCC.n282 VSS 0.003499f
C289 VCC.n283 VSS 0.002817f
C290 VCC.n284 VSS 0.003499f
C291 VCC.n285 VSS 0.106772f
C292 VCC.n286 VSS 0.003499f
C293 VCC.n287 VSS 0.002817f
C294 VCC.n288 VSS 0.003499f
C295 VCC.n289 VSS 0.003499f
C296 VCC.n290 VSS 0.003499f
C297 VCC.n291 VSS 0.002817f
C298 VCC.n292 VSS 0.003499f
C299 VCC.n293 VSS 0.106772f
C300 VCC.n294 VSS 0.003499f
C301 VCC.n295 VSS 0.002817f
C302 VCC.n296 VSS 0.003499f
C303 VCC.n297 VSS 0.003499f
C304 VCC.n298 VSS 0.003499f
C305 VCC.n299 VSS 0.002817f
C306 VCC.n300 VSS 0.003499f
C307 VCC.n301 VSS 0.070469f
C308 VCC.n302 VSS 0.106772f
C309 VCC.n303 VSS 0.003499f
C310 VCC.n304 VSS 0.002817f
C311 VCC.n305 VSS 0.003499f
C312 VCC.n306 VSS 0.003499f
C313 VCC.n307 VSS 0.003499f
C314 VCC.n308 VSS 0.002817f
C315 VCC.n309 VSS 0.003499f
C316 VCC.n310 VSS 0.089688f
C317 VCC.n311 VSS 0.003499f
C318 VCC.n312 VSS 0.002817f
C319 VCC.n313 VSS 0.003499f
C320 VCC.n314 VSS 0.003499f
C321 VCC.n315 VSS 0.003499f
C322 VCC.n316 VSS 0.002817f
C323 VCC.n317 VSS 0.003499f
C324 VCC.n318 VSS 0.106772f
C325 VCC.n319 VSS 0.003499f
C326 VCC.n320 VSS 0.002817f
C327 VCC.n321 VSS 0.003499f
C328 VCC.n322 VSS 0.003499f
C329 VCC.n323 VSS 0.003499f
C330 VCC.n324 VSS 0.002817f
C331 VCC.n325 VSS 0.003499f
C332 VCC.n326 VSS 0.106772f
C333 VCC.n327 VSS 0.003499f
C334 VCC.n328 VSS 0.002817f
C335 VCC.n329 VSS 0.003499f
C336 VCC.n330 VSS 0.003499f
C337 VCC.n331 VSS 0.003499f
C338 VCC.n332 VSS 0.002817f
C339 VCC.n333 VSS 0.003499f
C340 VCC.t0 VSS 0.053386f
C341 VCC.n334 VSS 0.088621f
C342 VCC.n335 VSS 0.003499f
C343 VCC.n336 VSS 0.002817f
C344 VCC.n337 VSS 0.003499f
C345 VCC.n338 VSS 0.003499f
C346 VCC.n339 VSS 0.003499f
C347 VCC.n340 VSS 0.002817f
C348 VCC.n341 VSS 0.003499f
C349 VCC.n342 VSS 0.106772f
C350 VCC.n343 VSS 0.003499f
C351 VCC.n344 VSS 0.002817f
C352 VCC.n345 VSS 0.003499f
C353 VCC.n346 VSS 0.003499f
C354 VCC.n347 VSS 0.003499f
C355 VCC.n348 VSS 0.002817f
C356 VCC.n349 VSS 0.003499f
C357 VCC.n350 VSS 0.106772f
C358 VCC.n351 VSS 0.003499f
C359 VCC.n352 VSS 0.002817f
C360 VCC.n353 VSS 0.003499f
C361 VCC.n354 VSS 0.003499f
C362 VCC.n355 VSS 0.003499f
C363 VCC.n356 VSS 0.002817f
C364 VCC.n357 VSS 0.003499f
C365 VCC.n358 VSS 0.106772f
C366 VCC.n359 VSS 0.003499f
C367 VCC.n360 VSS 0.002817f
C368 VCC.n361 VSS 0.003499f
C369 VCC.n362 VSS 0.003499f
C370 VCC.n363 VSS 0.003499f
C371 VCC.n364 VSS 0.002817f
C372 VCC.n365 VSS 0.003499f
C373 VCC.t2 VSS 0.106772f
C374 VCC.n366 VSS 0.106772f
C375 VCC.n367 VSS 0.106772f
C376 VCC.n368 VSS 0.003499f
C377 VCC.n369 VSS 0.002817f
C378 VCC.n370 VSS 0.003499f
C379 VCC.n371 VSS 0.003499f
C380 VCC.n372 VSS 0.003499f
C381 VCC.n373 VSS 0.002817f
C382 VCC.n374 VSS 0.003499f
C383 VCC.n375 VSS 0.106772f
C384 VCC.n376 VSS 0.106772f
C385 VCC.n377 VSS 0.003499f
C386 VCC.n378 VSS 0.071537f
C387 VCC.n379 VSS 0.106772f
C388 VCC.n380 VSS 0.003499f
C389 VCC.n381 VSS 0.002817f
C390 VCC.n382 VSS 0.003499f
C391 VCC.n383 VSS 0.003499f
C392 VCC.n384 VSS 0.003499f
C393 VCC.n385 VSS 0.002817f
C394 VCC.n386 VSS 0.003499f
C395 VCC.n387 VSS 0.088621f
C396 VCC.n388 VSS 0.106772f
C397 VCC.n389 VSS 0.106772f
C398 VCC.n390 VSS 0.003499f
C399 VCC.n391 VSS 0.002817f
C400 VCC.n392 VSS 0.003499f
C401 VCC.n393 VSS 0.003499f
C402 VCC.n394 VSS 0.003499f
C403 VCC.n395 VSS 0.002817f
C404 VCC.n396 VSS 0.003499f
C405 VCC.n397 VSS 0.106772f
C406 VCC.n398 VSS 0.106772f
C407 VCC.t4 VSS 0.053386f
C408 VCC.n399 VSS 0.089688f
C409 VCC.n400 VSS 0.003499f
C410 VCC.n401 VSS 0.002817f
C411 VCC.n402 VSS 0.003499f
C412 VCC.n403 VSS 0.003499f
C413 VCC.n404 VSS 0.003499f
C414 VCC.n405 VSS 0.002817f
C415 VCC.n406 VSS 0.003499f
C416 VCC.n407 VSS 0.106772f
C417 VCC.n408 VSS 0.106772f
C418 VCC.n409 VSS 0.106772f
C419 VCC.n410 VSS 0.003499f
C420 VCC.n411 VSS 0.002817f
C421 VCC.n412 VSS 0.003499f
C422 VCC.n413 VSS 0.003499f
C423 VCC.n414 VSS 0.003499f
C424 VCC.n415 VSS 0.002817f
C425 VCC.n416 VSS 0.003499f
C426 VCC.n417 VSS 0.106772f
C427 VCC.n418 VSS 0.106772f
C428 VCC.n419 VSS 0.106772f
C429 VCC.n420 VSS 0.003499f
C430 VCC.n421 VSS 0.002817f
C431 VCC.n422 VSS 0.003499f
C432 VCC.n423 VSS 0.003499f
C433 VCC.n424 VSS 0.003499f
C434 VCC.n425 VSS 0.002817f
C435 VCC.n426 VSS 0.003499f
C436 VCC.n427 VSS 0.064063f
C437 VCC.t10 VSS 0.053386f
C438 VCC.n428 VSS 0.096095f
C439 VCC.n429 VSS 0.106772f
C440 VCC.n430 VSS 0.003499f
C441 VCC.n431 VSS 0.002817f
C442 VCC.n432 VSS 0.003499f
C443 VCC.n433 VSS 0.003499f
C444 VCC.n434 VSS 0.00238f
C445 VCC.n435 VSS 0.00238f
C446 VCC.n436 VSS 0.00238f
C447 VCC.n437 VSS 0.00238f
C448 VCC.n438 VSS 0.00238f
C449 VCC.n439 VSS 0.00238f
C450 VCC.n440 VSS 0.00238f
C451 VCC.n441 VSS 0.00238f
C452 VCC.n442 VSS 0.00238f
C453 VCC.n443 VSS 0.00238f
C454 VCC.n444 VSS 0.00238f
C455 VCC.n445 VSS 0.00238f
C456 VCC.n446 VSS 0.00238f
C457 VCC.n447 VSS 0.00238f
C458 VCC.t12 VSS 0.088796f
C459 VCC.t11 VSS 0.097274f
C460 VCC.t9 VSS 0.44962f
C461 VCC.n448 VSS 0.054957f
C462 VCC.n449 VSS 0.023145f
C463 VCC.n451 VSS 0.00238f
C464 VCC.n452 VSS 0.001942f
C465 VCC.n453 VSS 0.003316f
C466 VCC.n454 VSS 0.001627f
C467 VCC.n455 VSS 0.00238f
C468 VCC.n456 VSS 0.00238f
C469 VCC.n458 VSS 0.00238f
C470 VCC.n460 VSS 0.00238f
C471 VCC.n461 VSS 0.00238f
C472 VCC.n462 VSS 0.00238f
C473 VCC.n463 VSS 0.00238f
C474 VCC.n464 VSS 0.00238f
C475 VCC.n466 VSS 0.00238f
C476 VCC.n468 VSS 0.00238f
C477 VCC.n469 VSS 0.00238f
C478 VCC.n470 VSS 0.00238f
C479 VCC.n471 VSS 0.00238f
C480 VCC.n472 VSS 0.00238f
C481 VCC.n474 VSS 0.00238f
C482 VCC.n476 VSS 0.00238f
C483 VCC.n477 VSS 0.00238f
C484 VCC.n478 VSS 0.00238f
C485 VCC.n479 VSS 0.00238f
C486 VCC.n480 VSS 0.00238f
C487 VCC.n482 VSS 0.00238f
C488 VCC.n484 VSS 0.00238f
C489 VCC.n485 VSS 0.00238f
C490 VCC.n486 VSS 0.00238f
C491 VCC.n487 VSS 0.00238f
C492 VCC.n488 VSS 0.00238f
C493 VCC.n490 VSS 0.00238f
C494 VCC.n492 VSS 0.00238f
C495 VCC.n493 VSS 0.00238f
C496 VCC.n494 VSS 0.00238f
C497 VCC.n495 VSS 0.00238f
C498 VCC.n496 VSS 0.00238f
C499 VCC.n498 VSS 0.00238f
C500 VCC.n500 VSS 0.00238f
C501 VCC.n501 VSS 0.00238f
C502 VCC.n502 VSS 0.00238f
C503 VCC.n503 VSS 0.00238f
C504 VCC.n504 VSS 0.00238f
C505 VCC.n506 VSS 0.00238f
C506 VCC.n508 VSS 0.00238f
C507 VCC.n509 VSS 0.00238f
C508 VCC.n510 VSS 0.004662f
C509 VCC.n511 VSS 0.01189f
C510 VCC.n512 VSS 0.002338f
C511 VCC.n513 VSS 0.006873f
C512 VCC.n514 VSS 0.148947f
C513 VCC.n515 VSS 0.006873f
C514 VCC.n516 VSS 0.002338f
C515 VCC.n517 VSS 0.01189f
C516 VCC.n518 VSS 0.003499f
C517 VCC.n519 VSS 0.003499f
C518 VCC.n520 VSS 0.002817f
C519 VCC.n521 VSS 0.002817f
C520 VCC.n522 VSS 0.002817f
C521 VCC.n523 VSS 0.003499f
C522 VCC.n524 VSS 0.003499f
C523 VCC.n525 VSS 0.003499f
C524 VCC.n526 VSS 0.002817f
C525 VCC.n527 VSS 0.002817f
C526 VCC.n528 VSS 0.002817f
C527 VCC.n529 VSS 0.003499f
C528 VCC.n530 VSS 0.003499f
C529 VCC.n531 VSS 0.003499f
C530 VCC.n532 VSS 0.002817f
C531 VCC.n533 VSS 0.002817f
C532 VCC.n534 VSS 0.002817f
C533 VCC.n535 VSS 0.003499f
C534 VCC.n536 VSS 0.003499f
C535 VCC.n537 VSS 0.003499f
C536 VCC.n538 VSS 0.002817f
C537 VCC.n539 VSS 0.002817f
C538 VCC.n540 VSS 0.002817f
C539 VCC.n541 VSS 0.003499f
C540 VCC.n542 VSS 0.003499f
C541 VCC.n543 VSS 0.003499f
C542 VCC.n544 VSS 0.002817f
C543 VCC.n545 VSS 0.002817f
C544 VCC.n546 VSS 0.002817f
C545 VCC.n547 VSS 0.003499f
C546 VCC.n548 VSS 0.003499f
C547 VCC.n549 VSS 0.003499f
C548 VCC.n550 VSS 0.002817f
C549 VCC.n551 VSS 0.002817f
C550 VCC.n552 VSS 0.002817f
C551 VCC.n553 VSS 0.003499f
C552 VCC.n554 VSS 0.003499f
C553 VCC.n555 VSS 0.003499f
C554 VCC.n556 VSS 0.002817f
C555 VCC.n557 VSS 0.002817f
C556 VCC.n558 VSS 0.002817f
C557 VCC.n559 VSS 0.003201f
C558 VOUT.t8 VSS 1.95755f
C559 VOUT.t5 VSS 0.202576f
C560 VOUT.t7 VSS 0.202576f
C561 VOUT.n0 VSS 1.45381f
C562 VOUT.n1 VSS 2.09716f
C563 VOUT.t6 VSS 0.202576f
C564 VOUT.t9 VSS 0.202576f
C565 VOUT.n2 VSS 1.45381f
C566 VOUT.n3 VSS 1.02993f
C567 VOUT.t4 VSS 0.15286f
C568 VOUT.t3 VSS 0.023634f
C569 VOUT.t2 VSS 0.023634f
C570 VOUT.n4 VSS 0.091799f
C571 VOUT.n5 VSS 1.40356f
C572 VOUT.t1 VSS 0.023634f
C573 VOUT.t0 VSS 0.023634f
C574 VOUT.n6 VSS 0.091799f
C575 VOUT.n7 VSS 1.06764f
C576 VIN.t9 VSS 1.52032f
C577 VIN.t6 VSS 0.169826f
C578 VIN.t7 VSS 0.169826f
C579 VIN.n0 VSS 1.0971f
C580 VIN.n1 VSS 1.93099f
C581 VIN.t5 VSS 0.169826f
C582 VIN.t8 VSS 0.169826f
C583 VIN.n2 VSS 1.0971f
C584 VIN.n3 VSS 1.30564f
C585 VIN.t0 VSS 0.115871f
C586 VIN.t2 VSS 0.019813f
C587 VIN.t1 VSS 0.019813f
C588 VIN.n4 VSS 0.064112f
C589 VIN.n5 VSS 1.13222f
C590 VIN.t4 VSS 0.019813f
C591 VIN.t3 VSS 0.019813f
C592 VIN.n6 VSS 0.064112f
C593 VIN.n7 VSS 0.560176f
C594 VGP.t1 VSS 1.83623f
C595 VGP.n0 VSS 0.760412f
C596 VGP.n1 VSS 0.024319f
C597 VGP.n2 VSS 0.019687f
C598 VGP.n3 VSS 0.024319f
C599 VGP.t4 VSS 1.83623f
C600 VGP.n4 VSS 0.65986f
C601 VGP.n5 VSS 0.024319f
C602 VGP.n6 VSS 0.029855f
C603 VGP.n7 VSS 0.024319f
C604 VGP.t2 VSS 1.83623f
C605 VGP.n8 VSS 0.682921f
C606 VGP.n9 VSS 0.024319f
C607 VGP.n10 VSS 0.029855f
C608 VGP.n11 VSS 0.024319f
C609 VGP.t3 VSS 1.83623f
C610 VGP.n12 VSS 0.738766f
C611 VGP.t0 VSS 2.13178f
C612 VGP.n13 VSS 0.703486f
C613 VGP.n14 VSS 0.286207f
C614 VGP.n15 VSS 0.030708f
C615 VGP.n16 VSS 0.045552f
C616 VGP.n17 VSS 0.045552f
C617 VGP.n18 VSS 0.024319f
C618 VGP.n19 VSS 0.024319f
C619 VGP.n20 VSS 0.024319f
C620 VGP.n21 VSS 0.041457f
C621 VGP.n22 VSS 0.045552f
C622 VGP.n23 VSS 0.045552f
C623 VGP.n24 VSS 0.024319f
C624 VGP.n25 VSS 0.024319f
C625 VGP.n26 VSS 0.024319f
C626 VGP.n27 VSS 0.045552f
C627 VGP.n28 VSS 0.045552f
C628 VGP.n29 VSS 0.041457f
C629 VGP.n30 VSS 0.024319f
C630 VGP.n31 VSS 0.024319f
C631 VGP.n32 VSS 0.024319f
C632 VGP.n33 VSS 0.045552f
C633 VGP.n34 VSS 0.045552f
C634 VGP.n35 VSS 0.030708f
C635 VGP.n36 VSS 0.024319f
C636 VGP.n37 VSS 0.024319f
C637 VGP.n38 VSS 0.037905f
C638 VGP.n39 VSS 0.045552f
C639 VGP.n40 VSS 0.048711f
C640 VGP.n41 VSS 0.024319f
C641 VGP.n42 VSS 0.024319f
C642 VGP.n43 VSS 0.024319f
C643 VGP.n44 VSS 0.048465f
C644 VGP.n45 VSS 0.045552f
C645 VGP.n46 VSS 0.038355f
C646 VGP.n47 VSS 0.039257f
C647 VGP.n48 VSS 0.068747f
.ends

