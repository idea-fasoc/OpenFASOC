* NGSPICE file created from diff_pair_sample_0537.ext - technology: sky130A

.subckt diff_pair_sample_0537 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=0 ps=0 w=10.28 l=1.83
X1 VTAIL.t11 VN.t0 VDD2.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=1.6962 ps=10.61 w=10.28 l=1.83
X2 VDD1.t5 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=4.0092 ps=21.34 w=10.28 l=1.83
X3 VTAIL.t10 VN.t1 VDD2.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=1.6962 ps=10.61 w=10.28 l=1.83
X4 VDD2.t3 VN.t2 VTAIL.t9 B.t0 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=4.0092 ps=21.34 w=10.28 l=1.83
X5 VDD1.t4 VP.t1 VTAIL.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=1.6962 ps=10.61 w=10.28 l=1.83
X6 VDD1.t3 VP.t2 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=1.6962 ps=10.61 w=10.28 l=1.83
X7 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=0 ps=0 w=10.28 l=1.83
X8 VDD2.t4 VN.t3 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=4.0092 ps=21.34 w=10.28 l=1.83
X9 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=0 ps=0 w=10.28 l=1.83
X10 VDD1.t2 VP.t3 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=4.0092 ps=21.34 w=10.28 l=1.83
X11 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=0 ps=0 w=10.28 l=1.83
X12 VDD2.t0 VN.t4 VTAIL.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=1.6962 ps=10.61 w=10.28 l=1.83
X13 VDD2.t5 VN.t5 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=4.0092 pd=21.34 as=1.6962 ps=10.61 w=10.28 l=1.83
X14 VTAIL.t3 VP.t4 VDD1.t1 B.t5 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=1.6962 ps=10.61 w=10.28 l=1.83
X15 VTAIL.t1 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.6962 pd=10.61 as=1.6962 ps=10.61 w=10.28 l=1.83
R0 B.n696 B.n695 585
R1 B.n697 B.n696 585
R2 B.n274 B.n105 585
R3 B.n273 B.n272 585
R4 B.n271 B.n270 585
R5 B.n269 B.n268 585
R6 B.n267 B.n266 585
R7 B.n265 B.n264 585
R8 B.n263 B.n262 585
R9 B.n261 B.n260 585
R10 B.n259 B.n258 585
R11 B.n257 B.n256 585
R12 B.n255 B.n254 585
R13 B.n253 B.n252 585
R14 B.n251 B.n250 585
R15 B.n249 B.n248 585
R16 B.n247 B.n246 585
R17 B.n245 B.n244 585
R18 B.n243 B.n242 585
R19 B.n241 B.n240 585
R20 B.n239 B.n238 585
R21 B.n237 B.n236 585
R22 B.n235 B.n234 585
R23 B.n233 B.n232 585
R24 B.n231 B.n230 585
R25 B.n229 B.n228 585
R26 B.n227 B.n226 585
R27 B.n225 B.n224 585
R28 B.n223 B.n222 585
R29 B.n221 B.n220 585
R30 B.n219 B.n218 585
R31 B.n217 B.n216 585
R32 B.n215 B.n214 585
R33 B.n213 B.n212 585
R34 B.n211 B.n210 585
R35 B.n209 B.n208 585
R36 B.n207 B.n206 585
R37 B.n205 B.n204 585
R38 B.n203 B.n202 585
R39 B.n201 B.n200 585
R40 B.n199 B.n198 585
R41 B.n197 B.n196 585
R42 B.n195 B.n194 585
R43 B.n193 B.n192 585
R44 B.n191 B.n190 585
R45 B.n189 B.n188 585
R46 B.n187 B.n186 585
R47 B.n184 B.n183 585
R48 B.n182 B.n181 585
R49 B.n180 B.n179 585
R50 B.n178 B.n177 585
R51 B.n176 B.n175 585
R52 B.n174 B.n173 585
R53 B.n172 B.n171 585
R54 B.n170 B.n169 585
R55 B.n168 B.n167 585
R56 B.n166 B.n165 585
R57 B.n164 B.n163 585
R58 B.n162 B.n161 585
R59 B.n160 B.n159 585
R60 B.n158 B.n157 585
R61 B.n156 B.n155 585
R62 B.n154 B.n153 585
R63 B.n152 B.n151 585
R64 B.n150 B.n149 585
R65 B.n148 B.n147 585
R66 B.n146 B.n145 585
R67 B.n144 B.n143 585
R68 B.n142 B.n141 585
R69 B.n140 B.n139 585
R70 B.n138 B.n137 585
R71 B.n136 B.n135 585
R72 B.n134 B.n133 585
R73 B.n132 B.n131 585
R74 B.n130 B.n129 585
R75 B.n128 B.n127 585
R76 B.n126 B.n125 585
R77 B.n124 B.n123 585
R78 B.n122 B.n121 585
R79 B.n120 B.n119 585
R80 B.n118 B.n117 585
R81 B.n116 B.n115 585
R82 B.n114 B.n113 585
R83 B.n112 B.n111 585
R84 B.n694 B.n63 585
R85 B.n698 B.n63 585
R86 B.n693 B.n62 585
R87 B.n699 B.n62 585
R88 B.n692 B.n691 585
R89 B.n691 B.n58 585
R90 B.n690 B.n57 585
R91 B.n705 B.n57 585
R92 B.n689 B.n56 585
R93 B.n706 B.n56 585
R94 B.n688 B.n55 585
R95 B.n707 B.n55 585
R96 B.n687 B.n686 585
R97 B.n686 B.n54 585
R98 B.n685 B.n50 585
R99 B.n713 B.n50 585
R100 B.n684 B.n49 585
R101 B.n714 B.n49 585
R102 B.n683 B.n48 585
R103 B.n715 B.n48 585
R104 B.n682 B.n681 585
R105 B.n681 B.n44 585
R106 B.n680 B.n43 585
R107 B.n721 B.n43 585
R108 B.n679 B.n42 585
R109 B.n722 B.n42 585
R110 B.n678 B.n41 585
R111 B.n723 B.n41 585
R112 B.n677 B.n676 585
R113 B.n676 B.n37 585
R114 B.n675 B.n36 585
R115 B.n729 B.n36 585
R116 B.n674 B.n35 585
R117 B.n730 B.n35 585
R118 B.n673 B.n34 585
R119 B.n731 B.n34 585
R120 B.n672 B.n671 585
R121 B.n671 B.n30 585
R122 B.n670 B.n29 585
R123 B.n737 B.n29 585
R124 B.n669 B.n28 585
R125 B.n738 B.n28 585
R126 B.n668 B.n27 585
R127 B.n739 B.n27 585
R128 B.n667 B.n666 585
R129 B.n666 B.n26 585
R130 B.n665 B.n22 585
R131 B.n745 B.n22 585
R132 B.n664 B.n21 585
R133 B.n746 B.n21 585
R134 B.n663 B.n20 585
R135 B.n747 B.n20 585
R136 B.n662 B.n661 585
R137 B.n661 B.n16 585
R138 B.n660 B.n15 585
R139 B.n753 B.n15 585
R140 B.n659 B.n14 585
R141 B.n754 B.n14 585
R142 B.n658 B.n13 585
R143 B.n755 B.n13 585
R144 B.n657 B.n656 585
R145 B.n656 B.n12 585
R146 B.n655 B.n654 585
R147 B.n655 B.n8 585
R148 B.n653 B.n7 585
R149 B.n762 B.n7 585
R150 B.n652 B.n6 585
R151 B.n763 B.n6 585
R152 B.n651 B.n5 585
R153 B.n764 B.n5 585
R154 B.n650 B.n649 585
R155 B.n649 B.n4 585
R156 B.n648 B.n275 585
R157 B.n648 B.n647 585
R158 B.n638 B.n276 585
R159 B.n277 B.n276 585
R160 B.n640 B.n639 585
R161 B.n641 B.n640 585
R162 B.n637 B.n281 585
R163 B.n285 B.n281 585
R164 B.n636 B.n635 585
R165 B.n635 B.n634 585
R166 B.n283 B.n282 585
R167 B.n284 B.n283 585
R168 B.n627 B.n626 585
R169 B.n628 B.n627 585
R170 B.n625 B.n290 585
R171 B.n290 B.n289 585
R172 B.n624 B.n623 585
R173 B.n623 B.n622 585
R174 B.n292 B.n291 585
R175 B.n615 B.n292 585
R176 B.n614 B.n613 585
R177 B.n616 B.n614 585
R178 B.n612 B.n297 585
R179 B.n297 B.n296 585
R180 B.n611 B.n610 585
R181 B.n610 B.n609 585
R182 B.n299 B.n298 585
R183 B.n300 B.n299 585
R184 B.n602 B.n601 585
R185 B.n603 B.n602 585
R186 B.n600 B.n304 585
R187 B.n308 B.n304 585
R188 B.n599 B.n598 585
R189 B.n598 B.n597 585
R190 B.n306 B.n305 585
R191 B.n307 B.n306 585
R192 B.n590 B.n589 585
R193 B.n591 B.n590 585
R194 B.n588 B.n313 585
R195 B.n313 B.n312 585
R196 B.n587 B.n586 585
R197 B.n586 B.n585 585
R198 B.n315 B.n314 585
R199 B.n316 B.n315 585
R200 B.n578 B.n577 585
R201 B.n579 B.n578 585
R202 B.n576 B.n321 585
R203 B.n321 B.n320 585
R204 B.n575 B.n574 585
R205 B.n574 B.n573 585
R206 B.n323 B.n322 585
R207 B.n566 B.n323 585
R208 B.n565 B.n564 585
R209 B.n567 B.n565 585
R210 B.n563 B.n328 585
R211 B.n328 B.n327 585
R212 B.n562 B.n561 585
R213 B.n561 B.n560 585
R214 B.n330 B.n329 585
R215 B.n331 B.n330 585
R216 B.n553 B.n552 585
R217 B.n554 B.n553 585
R218 B.n551 B.n336 585
R219 B.n336 B.n335 585
R220 B.n545 B.n544 585
R221 B.n543 B.n379 585
R222 B.n542 B.n378 585
R223 B.n547 B.n378 585
R224 B.n541 B.n540 585
R225 B.n539 B.n538 585
R226 B.n537 B.n536 585
R227 B.n535 B.n534 585
R228 B.n533 B.n532 585
R229 B.n531 B.n530 585
R230 B.n529 B.n528 585
R231 B.n527 B.n526 585
R232 B.n525 B.n524 585
R233 B.n523 B.n522 585
R234 B.n521 B.n520 585
R235 B.n519 B.n518 585
R236 B.n517 B.n516 585
R237 B.n515 B.n514 585
R238 B.n513 B.n512 585
R239 B.n511 B.n510 585
R240 B.n509 B.n508 585
R241 B.n507 B.n506 585
R242 B.n505 B.n504 585
R243 B.n503 B.n502 585
R244 B.n501 B.n500 585
R245 B.n499 B.n498 585
R246 B.n497 B.n496 585
R247 B.n495 B.n494 585
R248 B.n493 B.n492 585
R249 B.n491 B.n490 585
R250 B.n489 B.n488 585
R251 B.n487 B.n486 585
R252 B.n485 B.n484 585
R253 B.n483 B.n482 585
R254 B.n481 B.n480 585
R255 B.n479 B.n478 585
R256 B.n477 B.n476 585
R257 B.n475 B.n474 585
R258 B.n473 B.n472 585
R259 B.n471 B.n470 585
R260 B.n469 B.n468 585
R261 B.n467 B.n466 585
R262 B.n465 B.n464 585
R263 B.n463 B.n462 585
R264 B.n461 B.n460 585
R265 B.n459 B.n458 585
R266 B.n457 B.n456 585
R267 B.n454 B.n453 585
R268 B.n452 B.n451 585
R269 B.n450 B.n449 585
R270 B.n448 B.n447 585
R271 B.n446 B.n445 585
R272 B.n444 B.n443 585
R273 B.n442 B.n441 585
R274 B.n440 B.n439 585
R275 B.n438 B.n437 585
R276 B.n436 B.n435 585
R277 B.n434 B.n433 585
R278 B.n432 B.n431 585
R279 B.n430 B.n429 585
R280 B.n428 B.n427 585
R281 B.n426 B.n425 585
R282 B.n424 B.n423 585
R283 B.n422 B.n421 585
R284 B.n420 B.n419 585
R285 B.n418 B.n417 585
R286 B.n416 B.n415 585
R287 B.n414 B.n413 585
R288 B.n412 B.n411 585
R289 B.n410 B.n409 585
R290 B.n408 B.n407 585
R291 B.n406 B.n405 585
R292 B.n404 B.n403 585
R293 B.n402 B.n401 585
R294 B.n400 B.n399 585
R295 B.n398 B.n397 585
R296 B.n396 B.n395 585
R297 B.n394 B.n393 585
R298 B.n392 B.n391 585
R299 B.n390 B.n389 585
R300 B.n388 B.n387 585
R301 B.n386 B.n385 585
R302 B.n338 B.n337 585
R303 B.n550 B.n549 585
R304 B.n334 B.n333 585
R305 B.n335 B.n334 585
R306 B.n556 B.n555 585
R307 B.n555 B.n554 585
R308 B.n557 B.n332 585
R309 B.n332 B.n331 585
R310 B.n559 B.n558 585
R311 B.n560 B.n559 585
R312 B.n326 B.n325 585
R313 B.n327 B.n326 585
R314 B.n569 B.n568 585
R315 B.n568 B.n567 585
R316 B.n570 B.n324 585
R317 B.n566 B.n324 585
R318 B.n572 B.n571 585
R319 B.n573 B.n572 585
R320 B.n319 B.n318 585
R321 B.n320 B.n319 585
R322 B.n581 B.n580 585
R323 B.n580 B.n579 585
R324 B.n582 B.n317 585
R325 B.n317 B.n316 585
R326 B.n584 B.n583 585
R327 B.n585 B.n584 585
R328 B.n311 B.n310 585
R329 B.n312 B.n311 585
R330 B.n593 B.n592 585
R331 B.n592 B.n591 585
R332 B.n594 B.n309 585
R333 B.n309 B.n307 585
R334 B.n596 B.n595 585
R335 B.n597 B.n596 585
R336 B.n303 B.n302 585
R337 B.n308 B.n303 585
R338 B.n605 B.n604 585
R339 B.n604 B.n603 585
R340 B.n606 B.n301 585
R341 B.n301 B.n300 585
R342 B.n608 B.n607 585
R343 B.n609 B.n608 585
R344 B.n295 B.n294 585
R345 B.n296 B.n295 585
R346 B.n618 B.n617 585
R347 B.n617 B.n616 585
R348 B.n619 B.n293 585
R349 B.n615 B.n293 585
R350 B.n621 B.n620 585
R351 B.n622 B.n621 585
R352 B.n288 B.n287 585
R353 B.n289 B.n288 585
R354 B.n630 B.n629 585
R355 B.n629 B.n628 585
R356 B.n631 B.n286 585
R357 B.n286 B.n284 585
R358 B.n633 B.n632 585
R359 B.n634 B.n633 585
R360 B.n280 B.n279 585
R361 B.n285 B.n280 585
R362 B.n643 B.n642 585
R363 B.n642 B.n641 585
R364 B.n644 B.n278 585
R365 B.n278 B.n277 585
R366 B.n646 B.n645 585
R367 B.n647 B.n646 585
R368 B.n3 B.n0 585
R369 B.n4 B.n3 585
R370 B.n761 B.n1 585
R371 B.n762 B.n761 585
R372 B.n760 B.n759 585
R373 B.n760 B.n8 585
R374 B.n758 B.n9 585
R375 B.n12 B.n9 585
R376 B.n757 B.n756 585
R377 B.n756 B.n755 585
R378 B.n11 B.n10 585
R379 B.n754 B.n11 585
R380 B.n752 B.n751 585
R381 B.n753 B.n752 585
R382 B.n750 B.n17 585
R383 B.n17 B.n16 585
R384 B.n749 B.n748 585
R385 B.n748 B.n747 585
R386 B.n19 B.n18 585
R387 B.n746 B.n19 585
R388 B.n744 B.n743 585
R389 B.n745 B.n744 585
R390 B.n742 B.n23 585
R391 B.n26 B.n23 585
R392 B.n741 B.n740 585
R393 B.n740 B.n739 585
R394 B.n25 B.n24 585
R395 B.n738 B.n25 585
R396 B.n736 B.n735 585
R397 B.n737 B.n736 585
R398 B.n734 B.n31 585
R399 B.n31 B.n30 585
R400 B.n733 B.n732 585
R401 B.n732 B.n731 585
R402 B.n33 B.n32 585
R403 B.n730 B.n33 585
R404 B.n728 B.n727 585
R405 B.n729 B.n728 585
R406 B.n726 B.n38 585
R407 B.n38 B.n37 585
R408 B.n725 B.n724 585
R409 B.n724 B.n723 585
R410 B.n40 B.n39 585
R411 B.n722 B.n40 585
R412 B.n720 B.n719 585
R413 B.n721 B.n720 585
R414 B.n718 B.n45 585
R415 B.n45 B.n44 585
R416 B.n717 B.n716 585
R417 B.n716 B.n715 585
R418 B.n47 B.n46 585
R419 B.n714 B.n47 585
R420 B.n712 B.n711 585
R421 B.n713 B.n712 585
R422 B.n710 B.n51 585
R423 B.n54 B.n51 585
R424 B.n709 B.n708 585
R425 B.n708 B.n707 585
R426 B.n53 B.n52 585
R427 B.n706 B.n53 585
R428 B.n704 B.n703 585
R429 B.n705 B.n704 585
R430 B.n702 B.n59 585
R431 B.n59 B.n58 585
R432 B.n701 B.n700 585
R433 B.n700 B.n699 585
R434 B.n61 B.n60 585
R435 B.n698 B.n61 585
R436 B.n765 B.n764 585
R437 B.n763 B.n2 585
R438 B.n111 B.n61 478.086
R439 B.n696 B.n63 478.086
R440 B.n549 B.n336 478.086
R441 B.n545 B.n334 478.086
R442 B.n109 B.t17 341.87
R443 B.n106 B.t13 341.87
R444 B.n383 B.t6 341.87
R445 B.n380 B.t10 341.87
R446 B.n697 B.n104 256.663
R447 B.n697 B.n103 256.663
R448 B.n697 B.n102 256.663
R449 B.n697 B.n101 256.663
R450 B.n697 B.n100 256.663
R451 B.n697 B.n99 256.663
R452 B.n697 B.n98 256.663
R453 B.n697 B.n97 256.663
R454 B.n697 B.n96 256.663
R455 B.n697 B.n95 256.663
R456 B.n697 B.n94 256.663
R457 B.n697 B.n93 256.663
R458 B.n697 B.n92 256.663
R459 B.n697 B.n91 256.663
R460 B.n697 B.n90 256.663
R461 B.n697 B.n89 256.663
R462 B.n697 B.n88 256.663
R463 B.n697 B.n87 256.663
R464 B.n697 B.n86 256.663
R465 B.n697 B.n85 256.663
R466 B.n697 B.n84 256.663
R467 B.n697 B.n83 256.663
R468 B.n697 B.n82 256.663
R469 B.n697 B.n81 256.663
R470 B.n697 B.n80 256.663
R471 B.n697 B.n79 256.663
R472 B.n697 B.n78 256.663
R473 B.n697 B.n77 256.663
R474 B.n697 B.n76 256.663
R475 B.n697 B.n75 256.663
R476 B.n697 B.n74 256.663
R477 B.n697 B.n73 256.663
R478 B.n697 B.n72 256.663
R479 B.n697 B.n71 256.663
R480 B.n697 B.n70 256.663
R481 B.n697 B.n69 256.663
R482 B.n697 B.n68 256.663
R483 B.n697 B.n67 256.663
R484 B.n697 B.n66 256.663
R485 B.n697 B.n65 256.663
R486 B.n697 B.n64 256.663
R487 B.n547 B.n546 256.663
R488 B.n547 B.n339 256.663
R489 B.n547 B.n340 256.663
R490 B.n547 B.n341 256.663
R491 B.n547 B.n342 256.663
R492 B.n547 B.n343 256.663
R493 B.n547 B.n344 256.663
R494 B.n547 B.n345 256.663
R495 B.n547 B.n346 256.663
R496 B.n547 B.n347 256.663
R497 B.n547 B.n348 256.663
R498 B.n547 B.n349 256.663
R499 B.n547 B.n350 256.663
R500 B.n547 B.n351 256.663
R501 B.n547 B.n352 256.663
R502 B.n547 B.n353 256.663
R503 B.n547 B.n354 256.663
R504 B.n547 B.n355 256.663
R505 B.n547 B.n356 256.663
R506 B.n547 B.n357 256.663
R507 B.n547 B.n358 256.663
R508 B.n547 B.n359 256.663
R509 B.n547 B.n360 256.663
R510 B.n547 B.n361 256.663
R511 B.n547 B.n362 256.663
R512 B.n547 B.n363 256.663
R513 B.n547 B.n364 256.663
R514 B.n547 B.n365 256.663
R515 B.n547 B.n366 256.663
R516 B.n547 B.n367 256.663
R517 B.n547 B.n368 256.663
R518 B.n547 B.n369 256.663
R519 B.n547 B.n370 256.663
R520 B.n547 B.n371 256.663
R521 B.n547 B.n372 256.663
R522 B.n547 B.n373 256.663
R523 B.n547 B.n374 256.663
R524 B.n547 B.n375 256.663
R525 B.n547 B.n376 256.663
R526 B.n547 B.n377 256.663
R527 B.n548 B.n547 256.663
R528 B.n767 B.n766 256.663
R529 B.n115 B.n114 163.367
R530 B.n119 B.n118 163.367
R531 B.n123 B.n122 163.367
R532 B.n127 B.n126 163.367
R533 B.n131 B.n130 163.367
R534 B.n135 B.n134 163.367
R535 B.n139 B.n138 163.367
R536 B.n143 B.n142 163.367
R537 B.n147 B.n146 163.367
R538 B.n151 B.n150 163.367
R539 B.n155 B.n154 163.367
R540 B.n159 B.n158 163.367
R541 B.n163 B.n162 163.367
R542 B.n167 B.n166 163.367
R543 B.n171 B.n170 163.367
R544 B.n175 B.n174 163.367
R545 B.n179 B.n178 163.367
R546 B.n183 B.n182 163.367
R547 B.n188 B.n187 163.367
R548 B.n192 B.n191 163.367
R549 B.n196 B.n195 163.367
R550 B.n200 B.n199 163.367
R551 B.n204 B.n203 163.367
R552 B.n208 B.n207 163.367
R553 B.n212 B.n211 163.367
R554 B.n216 B.n215 163.367
R555 B.n220 B.n219 163.367
R556 B.n224 B.n223 163.367
R557 B.n228 B.n227 163.367
R558 B.n232 B.n231 163.367
R559 B.n236 B.n235 163.367
R560 B.n240 B.n239 163.367
R561 B.n244 B.n243 163.367
R562 B.n248 B.n247 163.367
R563 B.n252 B.n251 163.367
R564 B.n256 B.n255 163.367
R565 B.n260 B.n259 163.367
R566 B.n264 B.n263 163.367
R567 B.n268 B.n267 163.367
R568 B.n272 B.n271 163.367
R569 B.n696 B.n105 163.367
R570 B.n553 B.n336 163.367
R571 B.n553 B.n330 163.367
R572 B.n561 B.n330 163.367
R573 B.n561 B.n328 163.367
R574 B.n565 B.n328 163.367
R575 B.n565 B.n323 163.367
R576 B.n574 B.n323 163.367
R577 B.n574 B.n321 163.367
R578 B.n578 B.n321 163.367
R579 B.n578 B.n315 163.367
R580 B.n586 B.n315 163.367
R581 B.n586 B.n313 163.367
R582 B.n590 B.n313 163.367
R583 B.n590 B.n306 163.367
R584 B.n598 B.n306 163.367
R585 B.n598 B.n304 163.367
R586 B.n602 B.n304 163.367
R587 B.n602 B.n299 163.367
R588 B.n610 B.n299 163.367
R589 B.n610 B.n297 163.367
R590 B.n614 B.n297 163.367
R591 B.n614 B.n292 163.367
R592 B.n623 B.n292 163.367
R593 B.n623 B.n290 163.367
R594 B.n627 B.n290 163.367
R595 B.n627 B.n283 163.367
R596 B.n635 B.n283 163.367
R597 B.n635 B.n281 163.367
R598 B.n640 B.n281 163.367
R599 B.n640 B.n276 163.367
R600 B.n648 B.n276 163.367
R601 B.n649 B.n648 163.367
R602 B.n649 B.n5 163.367
R603 B.n6 B.n5 163.367
R604 B.n7 B.n6 163.367
R605 B.n655 B.n7 163.367
R606 B.n656 B.n655 163.367
R607 B.n656 B.n13 163.367
R608 B.n14 B.n13 163.367
R609 B.n15 B.n14 163.367
R610 B.n661 B.n15 163.367
R611 B.n661 B.n20 163.367
R612 B.n21 B.n20 163.367
R613 B.n22 B.n21 163.367
R614 B.n666 B.n22 163.367
R615 B.n666 B.n27 163.367
R616 B.n28 B.n27 163.367
R617 B.n29 B.n28 163.367
R618 B.n671 B.n29 163.367
R619 B.n671 B.n34 163.367
R620 B.n35 B.n34 163.367
R621 B.n36 B.n35 163.367
R622 B.n676 B.n36 163.367
R623 B.n676 B.n41 163.367
R624 B.n42 B.n41 163.367
R625 B.n43 B.n42 163.367
R626 B.n681 B.n43 163.367
R627 B.n681 B.n48 163.367
R628 B.n49 B.n48 163.367
R629 B.n50 B.n49 163.367
R630 B.n686 B.n50 163.367
R631 B.n686 B.n55 163.367
R632 B.n56 B.n55 163.367
R633 B.n57 B.n56 163.367
R634 B.n691 B.n57 163.367
R635 B.n691 B.n62 163.367
R636 B.n63 B.n62 163.367
R637 B.n379 B.n378 163.367
R638 B.n540 B.n378 163.367
R639 B.n538 B.n537 163.367
R640 B.n534 B.n533 163.367
R641 B.n530 B.n529 163.367
R642 B.n526 B.n525 163.367
R643 B.n522 B.n521 163.367
R644 B.n518 B.n517 163.367
R645 B.n514 B.n513 163.367
R646 B.n510 B.n509 163.367
R647 B.n506 B.n505 163.367
R648 B.n502 B.n501 163.367
R649 B.n498 B.n497 163.367
R650 B.n494 B.n493 163.367
R651 B.n490 B.n489 163.367
R652 B.n486 B.n485 163.367
R653 B.n482 B.n481 163.367
R654 B.n478 B.n477 163.367
R655 B.n474 B.n473 163.367
R656 B.n470 B.n469 163.367
R657 B.n466 B.n465 163.367
R658 B.n462 B.n461 163.367
R659 B.n458 B.n457 163.367
R660 B.n453 B.n452 163.367
R661 B.n449 B.n448 163.367
R662 B.n445 B.n444 163.367
R663 B.n441 B.n440 163.367
R664 B.n437 B.n436 163.367
R665 B.n433 B.n432 163.367
R666 B.n429 B.n428 163.367
R667 B.n425 B.n424 163.367
R668 B.n421 B.n420 163.367
R669 B.n417 B.n416 163.367
R670 B.n413 B.n412 163.367
R671 B.n409 B.n408 163.367
R672 B.n405 B.n404 163.367
R673 B.n401 B.n400 163.367
R674 B.n397 B.n396 163.367
R675 B.n393 B.n392 163.367
R676 B.n389 B.n388 163.367
R677 B.n385 B.n338 163.367
R678 B.n555 B.n334 163.367
R679 B.n555 B.n332 163.367
R680 B.n559 B.n332 163.367
R681 B.n559 B.n326 163.367
R682 B.n568 B.n326 163.367
R683 B.n568 B.n324 163.367
R684 B.n572 B.n324 163.367
R685 B.n572 B.n319 163.367
R686 B.n580 B.n319 163.367
R687 B.n580 B.n317 163.367
R688 B.n584 B.n317 163.367
R689 B.n584 B.n311 163.367
R690 B.n592 B.n311 163.367
R691 B.n592 B.n309 163.367
R692 B.n596 B.n309 163.367
R693 B.n596 B.n303 163.367
R694 B.n604 B.n303 163.367
R695 B.n604 B.n301 163.367
R696 B.n608 B.n301 163.367
R697 B.n608 B.n295 163.367
R698 B.n617 B.n295 163.367
R699 B.n617 B.n293 163.367
R700 B.n621 B.n293 163.367
R701 B.n621 B.n288 163.367
R702 B.n629 B.n288 163.367
R703 B.n629 B.n286 163.367
R704 B.n633 B.n286 163.367
R705 B.n633 B.n280 163.367
R706 B.n642 B.n280 163.367
R707 B.n642 B.n278 163.367
R708 B.n646 B.n278 163.367
R709 B.n646 B.n3 163.367
R710 B.n765 B.n3 163.367
R711 B.n761 B.n2 163.367
R712 B.n761 B.n760 163.367
R713 B.n760 B.n9 163.367
R714 B.n756 B.n9 163.367
R715 B.n756 B.n11 163.367
R716 B.n752 B.n11 163.367
R717 B.n752 B.n17 163.367
R718 B.n748 B.n17 163.367
R719 B.n748 B.n19 163.367
R720 B.n744 B.n19 163.367
R721 B.n744 B.n23 163.367
R722 B.n740 B.n23 163.367
R723 B.n740 B.n25 163.367
R724 B.n736 B.n25 163.367
R725 B.n736 B.n31 163.367
R726 B.n732 B.n31 163.367
R727 B.n732 B.n33 163.367
R728 B.n728 B.n33 163.367
R729 B.n728 B.n38 163.367
R730 B.n724 B.n38 163.367
R731 B.n724 B.n40 163.367
R732 B.n720 B.n40 163.367
R733 B.n720 B.n45 163.367
R734 B.n716 B.n45 163.367
R735 B.n716 B.n47 163.367
R736 B.n712 B.n47 163.367
R737 B.n712 B.n51 163.367
R738 B.n708 B.n51 163.367
R739 B.n708 B.n53 163.367
R740 B.n704 B.n53 163.367
R741 B.n704 B.n59 163.367
R742 B.n700 B.n59 163.367
R743 B.n700 B.n61 163.367
R744 B.n106 B.t15 111.505
R745 B.n383 B.t9 111.505
R746 B.n109 B.t18 111.493
R747 B.n380 B.t12 111.493
R748 B.n547 B.n335 88.3965
R749 B.n698 B.n697 88.3965
R750 B.n111 B.n64 71.676
R751 B.n115 B.n65 71.676
R752 B.n119 B.n66 71.676
R753 B.n123 B.n67 71.676
R754 B.n127 B.n68 71.676
R755 B.n131 B.n69 71.676
R756 B.n135 B.n70 71.676
R757 B.n139 B.n71 71.676
R758 B.n143 B.n72 71.676
R759 B.n147 B.n73 71.676
R760 B.n151 B.n74 71.676
R761 B.n155 B.n75 71.676
R762 B.n159 B.n76 71.676
R763 B.n163 B.n77 71.676
R764 B.n167 B.n78 71.676
R765 B.n171 B.n79 71.676
R766 B.n175 B.n80 71.676
R767 B.n179 B.n81 71.676
R768 B.n183 B.n82 71.676
R769 B.n188 B.n83 71.676
R770 B.n192 B.n84 71.676
R771 B.n196 B.n85 71.676
R772 B.n200 B.n86 71.676
R773 B.n204 B.n87 71.676
R774 B.n208 B.n88 71.676
R775 B.n212 B.n89 71.676
R776 B.n216 B.n90 71.676
R777 B.n220 B.n91 71.676
R778 B.n224 B.n92 71.676
R779 B.n228 B.n93 71.676
R780 B.n232 B.n94 71.676
R781 B.n236 B.n95 71.676
R782 B.n240 B.n96 71.676
R783 B.n244 B.n97 71.676
R784 B.n248 B.n98 71.676
R785 B.n252 B.n99 71.676
R786 B.n256 B.n100 71.676
R787 B.n260 B.n101 71.676
R788 B.n264 B.n102 71.676
R789 B.n268 B.n103 71.676
R790 B.n272 B.n104 71.676
R791 B.n105 B.n104 71.676
R792 B.n271 B.n103 71.676
R793 B.n267 B.n102 71.676
R794 B.n263 B.n101 71.676
R795 B.n259 B.n100 71.676
R796 B.n255 B.n99 71.676
R797 B.n251 B.n98 71.676
R798 B.n247 B.n97 71.676
R799 B.n243 B.n96 71.676
R800 B.n239 B.n95 71.676
R801 B.n235 B.n94 71.676
R802 B.n231 B.n93 71.676
R803 B.n227 B.n92 71.676
R804 B.n223 B.n91 71.676
R805 B.n219 B.n90 71.676
R806 B.n215 B.n89 71.676
R807 B.n211 B.n88 71.676
R808 B.n207 B.n87 71.676
R809 B.n203 B.n86 71.676
R810 B.n199 B.n85 71.676
R811 B.n195 B.n84 71.676
R812 B.n191 B.n83 71.676
R813 B.n187 B.n82 71.676
R814 B.n182 B.n81 71.676
R815 B.n178 B.n80 71.676
R816 B.n174 B.n79 71.676
R817 B.n170 B.n78 71.676
R818 B.n166 B.n77 71.676
R819 B.n162 B.n76 71.676
R820 B.n158 B.n75 71.676
R821 B.n154 B.n74 71.676
R822 B.n150 B.n73 71.676
R823 B.n146 B.n72 71.676
R824 B.n142 B.n71 71.676
R825 B.n138 B.n70 71.676
R826 B.n134 B.n69 71.676
R827 B.n130 B.n68 71.676
R828 B.n126 B.n67 71.676
R829 B.n122 B.n66 71.676
R830 B.n118 B.n65 71.676
R831 B.n114 B.n64 71.676
R832 B.n546 B.n545 71.676
R833 B.n540 B.n339 71.676
R834 B.n537 B.n340 71.676
R835 B.n533 B.n341 71.676
R836 B.n529 B.n342 71.676
R837 B.n525 B.n343 71.676
R838 B.n521 B.n344 71.676
R839 B.n517 B.n345 71.676
R840 B.n513 B.n346 71.676
R841 B.n509 B.n347 71.676
R842 B.n505 B.n348 71.676
R843 B.n501 B.n349 71.676
R844 B.n497 B.n350 71.676
R845 B.n493 B.n351 71.676
R846 B.n489 B.n352 71.676
R847 B.n485 B.n353 71.676
R848 B.n481 B.n354 71.676
R849 B.n477 B.n355 71.676
R850 B.n473 B.n356 71.676
R851 B.n469 B.n357 71.676
R852 B.n465 B.n358 71.676
R853 B.n461 B.n359 71.676
R854 B.n457 B.n360 71.676
R855 B.n452 B.n361 71.676
R856 B.n448 B.n362 71.676
R857 B.n444 B.n363 71.676
R858 B.n440 B.n364 71.676
R859 B.n436 B.n365 71.676
R860 B.n432 B.n366 71.676
R861 B.n428 B.n367 71.676
R862 B.n424 B.n368 71.676
R863 B.n420 B.n369 71.676
R864 B.n416 B.n370 71.676
R865 B.n412 B.n371 71.676
R866 B.n408 B.n372 71.676
R867 B.n404 B.n373 71.676
R868 B.n400 B.n374 71.676
R869 B.n396 B.n375 71.676
R870 B.n392 B.n376 71.676
R871 B.n388 B.n377 71.676
R872 B.n548 B.n338 71.676
R873 B.n546 B.n379 71.676
R874 B.n538 B.n339 71.676
R875 B.n534 B.n340 71.676
R876 B.n530 B.n341 71.676
R877 B.n526 B.n342 71.676
R878 B.n522 B.n343 71.676
R879 B.n518 B.n344 71.676
R880 B.n514 B.n345 71.676
R881 B.n510 B.n346 71.676
R882 B.n506 B.n347 71.676
R883 B.n502 B.n348 71.676
R884 B.n498 B.n349 71.676
R885 B.n494 B.n350 71.676
R886 B.n490 B.n351 71.676
R887 B.n486 B.n352 71.676
R888 B.n482 B.n353 71.676
R889 B.n478 B.n354 71.676
R890 B.n474 B.n355 71.676
R891 B.n470 B.n356 71.676
R892 B.n466 B.n357 71.676
R893 B.n462 B.n358 71.676
R894 B.n458 B.n359 71.676
R895 B.n453 B.n360 71.676
R896 B.n449 B.n361 71.676
R897 B.n445 B.n362 71.676
R898 B.n441 B.n363 71.676
R899 B.n437 B.n364 71.676
R900 B.n433 B.n365 71.676
R901 B.n429 B.n366 71.676
R902 B.n425 B.n367 71.676
R903 B.n421 B.n368 71.676
R904 B.n417 B.n369 71.676
R905 B.n413 B.n370 71.676
R906 B.n409 B.n371 71.676
R907 B.n405 B.n372 71.676
R908 B.n401 B.n373 71.676
R909 B.n397 B.n374 71.676
R910 B.n393 B.n375 71.676
R911 B.n389 B.n376 71.676
R912 B.n385 B.n377 71.676
R913 B.n549 B.n548 71.676
R914 B.n766 B.n765 71.676
R915 B.n766 B.n2 71.676
R916 B.n107 B.t16 69.615
R917 B.n384 B.t8 69.615
R918 B.n110 B.t19 69.6023
R919 B.n381 B.t11 69.6023
R920 B.n185 B.n110 59.5399
R921 B.n108 B.n107 59.5399
R922 B.n455 B.n384 59.5399
R923 B.n382 B.n381 59.5399
R924 B.n554 B.n335 48.0879
R925 B.n554 B.n331 48.0879
R926 B.n560 B.n331 48.0879
R927 B.n560 B.n327 48.0879
R928 B.n567 B.n327 48.0879
R929 B.n567 B.n566 48.0879
R930 B.n573 B.n320 48.0879
R931 B.n579 B.n320 48.0879
R932 B.n579 B.n316 48.0879
R933 B.n585 B.n316 48.0879
R934 B.n585 B.n312 48.0879
R935 B.n591 B.n312 48.0879
R936 B.n591 B.n307 48.0879
R937 B.n597 B.n307 48.0879
R938 B.n597 B.n308 48.0879
R939 B.n603 B.n300 48.0879
R940 B.n609 B.n300 48.0879
R941 B.n609 B.n296 48.0879
R942 B.n616 B.n296 48.0879
R943 B.n616 B.n615 48.0879
R944 B.n622 B.n289 48.0879
R945 B.n628 B.n289 48.0879
R946 B.n628 B.n284 48.0879
R947 B.n634 B.n284 48.0879
R948 B.n634 B.n285 48.0879
R949 B.n641 B.n277 48.0879
R950 B.n647 B.n277 48.0879
R951 B.n647 B.n4 48.0879
R952 B.n764 B.n4 48.0879
R953 B.n764 B.n763 48.0879
R954 B.n763 B.n762 48.0879
R955 B.n762 B.n8 48.0879
R956 B.n12 B.n8 48.0879
R957 B.n755 B.n12 48.0879
R958 B.n754 B.n753 48.0879
R959 B.n753 B.n16 48.0879
R960 B.n747 B.n16 48.0879
R961 B.n747 B.n746 48.0879
R962 B.n746 B.n745 48.0879
R963 B.n739 B.n26 48.0879
R964 B.n739 B.n738 48.0879
R965 B.n738 B.n737 48.0879
R966 B.n737 B.n30 48.0879
R967 B.n731 B.n30 48.0879
R968 B.n730 B.n729 48.0879
R969 B.n729 B.n37 48.0879
R970 B.n723 B.n37 48.0879
R971 B.n723 B.n722 48.0879
R972 B.n722 B.n721 48.0879
R973 B.n721 B.n44 48.0879
R974 B.n715 B.n44 48.0879
R975 B.n715 B.n714 48.0879
R976 B.n714 B.n713 48.0879
R977 B.n707 B.n54 48.0879
R978 B.n707 B.n706 48.0879
R979 B.n706 B.n705 48.0879
R980 B.n705 B.n58 48.0879
R981 B.n699 B.n58 48.0879
R982 B.n699 B.n698 48.0879
R983 B.n603 B.t1 47.3808
R984 B.n731 B.t0 47.3808
R985 B.n110 B.n109 41.8914
R986 B.n107 B.n106 41.8914
R987 B.n384 B.n383 41.8914
R988 B.n381 B.n380 41.8914
R989 B.n285 B.t2 34.6517
R990 B.t4 B.n754 34.6517
R991 B.n544 B.n333 31.0639
R992 B.n551 B.n550 31.0639
R993 B.n695 B.n694 31.0639
R994 B.n112 B.n60 31.0639
R995 B.n622 B.t3 30.4087
R996 B.n745 B.t5 30.4087
R997 B.n573 B.t7 26.1657
R998 B.n713 B.t14 26.1657
R999 B.n566 B.t7 21.9227
R1000 B.n54 B.t14 21.9227
R1001 B B.n767 18.0485
R1002 B.n615 B.t3 17.6797
R1003 B.n26 B.t5 17.6797
R1004 B.n641 B.t2 13.4367
R1005 B.n755 B.t4 13.4367
R1006 B.n556 B.n333 10.6151
R1007 B.n557 B.n556 10.6151
R1008 B.n558 B.n557 10.6151
R1009 B.n558 B.n325 10.6151
R1010 B.n569 B.n325 10.6151
R1011 B.n570 B.n569 10.6151
R1012 B.n571 B.n570 10.6151
R1013 B.n571 B.n318 10.6151
R1014 B.n581 B.n318 10.6151
R1015 B.n582 B.n581 10.6151
R1016 B.n583 B.n582 10.6151
R1017 B.n583 B.n310 10.6151
R1018 B.n593 B.n310 10.6151
R1019 B.n594 B.n593 10.6151
R1020 B.n595 B.n594 10.6151
R1021 B.n595 B.n302 10.6151
R1022 B.n605 B.n302 10.6151
R1023 B.n606 B.n605 10.6151
R1024 B.n607 B.n606 10.6151
R1025 B.n607 B.n294 10.6151
R1026 B.n618 B.n294 10.6151
R1027 B.n619 B.n618 10.6151
R1028 B.n620 B.n619 10.6151
R1029 B.n620 B.n287 10.6151
R1030 B.n630 B.n287 10.6151
R1031 B.n631 B.n630 10.6151
R1032 B.n632 B.n631 10.6151
R1033 B.n632 B.n279 10.6151
R1034 B.n643 B.n279 10.6151
R1035 B.n644 B.n643 10.6151
R1036 B.n645 B.n644 10.6151
R1037 B.n645 B.n0 10.6151
R1038 B.n544 B.n543 10.6151
R1039 B.n543 B.n542 10.6151
R1040 B.n542 B.n541 10.6151
R1041 B.n541 B.n539 10.6151
R1042 B.n539 B.n536 10.6151
R1043 B.n536 B.n535 10.6151
R1044 B.n535 B.n532 10.6151
R1045 B.n532 B.n531 10.6151
R1046 B.n531 B.n528 10.6151
R1047 B.n528 B.n527 10.6151
R1048 B.n527 B.n524 10.6151
R1049 B.n524 B.n523 10.6151
R1050 B.n523 B.n520 10.6151
R1051 B.n520 B.n519 10.6151
R1052 B.n519 B.n516 10.6151
R1053 B.n516 B.n515 10.6151
R1054 B.n515 B.n512 10.6151
R1055 B.n512 B.n511 10.6151
R1056 B.n511 B.n508 10.6151
R1057 B.n508 B.n507 10.6151
R1058 B.n507 B.n504 10.6151
R1059 B.n504 B.n503 10.6151
R1060 B.n503 B.n500 10.6151
R1061 B.n500 B.n499 10.6151
R1062 B.n499 B.n496 10.6151
R1063 B.n496 B.n495 10.6151
R1064 B.n495 B.n492 10.6151
R1065 B.n492 B.n491 10.6151
R1066 B.n491 B.n488 10.6151
R1067 B.n488 B.n487 10.6151
R1068 B.n487 B.n484 10.6151
R1069 B.n484 B.n483 10.6151
R1070 B.n483 B.n480 10.6151
R1071 B.n480 B.n479 10.6151
R1072 B.n479 B.n476 10.6151
R1073 B.n476 B.n475 10.6151
R1074 B.n472 B.n471 10.6151
R1075 B.n471 B.n468 10.6151
R1076 B.n468 B.n467 10.6151
R1077 B.n467 B.n464 10.6151
R1078 B.n464 B.n463 10.6151
R1079 B.n463 B.n460 10.6151
R1080 B.n460 B.n459 10.6151
R1081 B.n459 B.n456 10.6151
R1082 B.n454 B.n451 10.6151
R1083 B.n451 B.n450 10.6151
R1084 B.n450 B.n447 10.6151
R1085 B.n447 B.n446 10.6151
R1086 B.n446 B.n443 10.6151
R1087 B.n443 B.n442 10.6151
R1088 B.n442 B.n439 10.6151
R1089 B.n439 B.n438 10.6151
R1090 B.n438 B.n435 10.6151
R1091 B.n435 B.n434 10.6151
R1092 B.n434 B.n431 10.6151
R1093 B.n431 B.n430 10.6151
R1094 B.n430 B.n427 10.6151
R1095 B.n427 B.n426 10.6151
R1096 B.n426 B.n423 10.6151
R1097 B.n423 B.n422 10.6151
R1098 B.n422 B.n419 10.6151
R1099 B.n419 B.n418 10.6151
R1100 B.n418 B.n415 10.6151
R1101 B.n415 B.n414 10.6151
R1102 B.n414 B.n411 10.6151
R1103 B.n411 B.n410 10.6151
R1104 B.n410 B.n407 10.6151
R1105 B.n407 B.n406 10.6151
R1106 B.n406 B.n403 10.6151
R1107 B.n403 B.n402 10.6151
R1108 B.n402 B.n399 10.6151
R1109 B.n399 B.n398 10.6151
R1110 B.n398 B.n395 10.6151
R1111 B.n395 B.n394 10.6151
R1112 B.n394 B.n391 10.6151
R1113 B.n391 B.n390 10.6151
R1114 B.n390 B.n387 10.6151
R1115 B.n387 B.n386 10.6151
R1116 B.n386 B.n337 10.6151
R1117 B.n550 B.n337 10.6151
R1118 B.n552 B.n551 10.6151
R1119 B.n552 B.n329 10.6151
R1120 B.n562 B.n329 10.6151
R1121 B.n563 B.n562 10.6151
R1122 B.n564 B.n563 10.6151
R1123 B.n564 B.n322 10.6151
R1124 B.n575 B.n322 10.6151
R1125 B.n576 B.n575 10.6151
R1126 B.n577 B.n576 10.6151
R1127 B.n577 B.n314 10.6151
R1128 B.n587 B.n314 10.6151
R1129 B.n588 B.n587 10.6151
R1130 B.n589 B.n588 10.6151
R1131 B.n589 B.n305 10.6151
R1132 B.n599 B.n305 10.6151
R1133 B.n600 B.n599 10.6151
R1134 B.n601 B.n600 10.6151
R1135 B.n601 B.n298 10.6151
R1136 B.n611 B.n298 10.6151
R1137 B.n612 B.n611 10.6151
R1138 B.n613 B.n612 10.6151
R1139 B.n613 B.n291 10.6151
R1140 B.n624 B.n291 10.6151
R1141 B.n625 B.n624 10.6151
R1142 B.n626 B.n625 10.6151
R1143 B.n626 B.n282 10.6151
R1144 B.n636 B.n282 10.6151
R1145 B.n637 B.n636 10.6151
R1146 B.n639 B.n637 10.6151
R1147 B.n639 B.n638 10.6151
R1148 B.n638 B.n275 10.6151
R1149 B.n650 B.n275 10.6151
R1150 B.n651 B.n650 10.6151
R1151 B.n652 B.n651 10.6151
R1152 B.n653 B.n652 10.6151
R1153 B.n654 B.n653 10.6151
R1154 B.n657 B.n654 10.6151
R1155 B.n658 B.n657 10.6151
R1156 B.n659 B.n658 10.6151
R1157 B.n660 B.n659 10.6151
R1158 B.n662 B.n660 10.6151
R1159 B.n663 B.n662 10.6151
R1160 B.n664 B.n663 10.6151
R1161 B.n665 B.n664 10.6151
R1162 B.n667 B.n665 10.6151
R1163 B.n668 B.n667 10.6151
R1164 B.n669 B.n668 10.6151
R1165 B.n670 B.n669 10.6151
R1166 B.n672 B.n670 10.6151
R1167 B.n673 B.n672 10.6151
R1168 B.n674 B.n673 10.6151
R1169 B.n675 B.n674 10.6151
R1170 B.n677 B.n675 10.6151
R1171 B.n678 B.n677 10.6151
R1172 B.n679 B.n678 10.6151
R1173 B.n680 B.n679 10.6151
R1174 B.n682 B.n680 10.6151
R1175 B.n683 B.n682 10.6151
R1176 B.n684 B.n683 10.6151
R1177 B.n685 B.n684 10.6151
R1178 B.n687 B.n685 10.6151
R1179 B.n688 B.n687 10.6151
R1180 B.n689 B.n688 10.6151
R1181 B.n690 B.n689 10.6151
R1182 B.n692 B.n690 10.6151
R1183 B.n693 B.n692 10.6151
R1184 B.n694 B.n693 10.6151
R1185 B.n759 B.n1 10.6151
R1186 B.n759 B.n758 10.6151
R1187 B.n758 B.n757 10.6151
R1188 B.n757 B.n10 10.6151
R1189 B.n751 B.n10 10.6151
R1190 B.n751 B.n750 10.6151
R1191 B.n750 B.n749 10.6151
R1192 B.n749 B.n18 10.6151
R1193 B.n743 B.n18 10.6151
R1194 B.n743 B.n742 10.6151
R1195 B.n742 B.n741 10.6151
R1196 B.n741 B.n24 10.6151
R1197 B.n735 B.n24 10.6151
R1198 B.n735 B.n734 10.6151
R1199 B.n734 B.n733 10.6151
R1200 B.n733 B.n32 10.6151
R1201 B.n727 B.n32 10.6151
R1202 B.n727 B.n726 10.6151
R1203 B.n726 B.n725 10.6151
R1204 B.n725 B.n39 10.6151
R1205 B.n719 B.n39 10.6151
R1206 B.n719 B.n718 10.6151
R1207 B.n718 B.n717 10.6151
R1208 B.n717 B.n46 10.6151
R1209 B.n711 B.n46 10.6151
R1210 B.n711 B.n710 10.6151
R1211 B.n710 B.n709 10.6151
R1212 B.n709 B.n52 10.6151
R1213 B.n703 B.n52 10.6151
R1214 B.n703 B.n702 10.6151
R1215 B.n702 B.n701 10.6151
R1216 B.n701 B.n60 10.6151
R1217 B.n113 B.n112 10.6151
R1218 B.n116 B.n113 10.6151
R1219 B.n117 B.n116 10.6151
R1220 B.n120 B.n117 10.6151
R1221 B.n121 B.n120 10.6151
R1222 B.n124 B.n121 10.6151
R1223 B.n125 B.n124 10.6151
R1224 B.n128 B.n125 10.6151
R1225 B.n129 B.n128 10.6151
R1226 B.n132 B.n129 10.6151
R1227 B.n133 B.n132 10.6151
R1228 B.n136 B.n133 10.6151
R1229 B.n137 B.n136 10.6151
R1230 B.n140 B.n137 10.6151
R1231 B.n141 B.n140 10.6151
R1232 B.n144 B.n141 10.6151
R1233 B.n145 B.n144 10.6151
R1234 B.n148 B.n145 10.6151
R1235 B.n149 B.n148 10.6151
R1236 B.n152 B.n149 10.6151
R1237 B.n153 B.n152 10.6151
R1238 B.n156 B.n153 10.6151
R1239 B.n157 B.n156 10.6151
R1240 B.n160 B.n157 10.6151
R1241 B.n161 B.n160 10.6151
R1242 B.n164 B.n161 10.6151
R1243 B.n165 B.n164 10.6151
R1244 B.n168 B.n165 10.6151
R1245 B.n169 B.n168 10.6151
R1246 B.n172 B.n169 10.6151
R1247 B.n173 B.n172 10.6151
R1248 B.n176 B.n173 10.6151
R1249 B.n177 B.n176 10.6151
R1250 B.n180 B.n177 10.6151
R1251 B.n181 B.n180 10.6151
R1252 B.n184 B.n181 10.6151
R1253 B.n189 B.n186 10.6151
R1254 B.n190 B.n189 10.6151
R1255 B.n193 B.n190 10.6151
R1256 B.n194 B.n193 10.6151
R1257 B.n197 B.n194 10.6151
R1258 B.n198 B.n197 10.6151
R1259 B.n201 B.n198 10.6151
R1260 B.n202 B.n201 10.6151
R1261 B.n206 B.n205 10.6151
R1262 B.n209 B.n206 10.6151
R1263 B.n210 B.n209 10.6151
R1264 B.n213 B.n210 10.6151
R1265 B.n214 B.n213 10.6151
R1266 B.n217 B.n214 10.6151
R1267 B.n218 B.n217 10.6151
R1268 B.n221 B.n218 10.6151
R1269 B.n222 B.n221 10.6151
R1270 B.n225 B.n222 10.6151
R1271 B.n226 B.n225 10.6151
R1272 B.n229 B.n226 10.6151
R1273 B.n230 B.n229 10.6151
R1274 B.n233 B.n230 10.6151
R1275 B.n234 B.n233 10.6151
R1276 B.n237 B.n234 10.6151
R1277 B.n238 B.n237 10.6151
R1278 B.n241 B.n238 10.6151
R1279 B.n242 B.n241 10.6151
R1280 B.n245 B.n242 10.6151
R1281 B.n246 B.n245 10.6151
R1282 B.n249 B.n246 10.6151
R1283 B.n250 B.n249 10.6151
R1284 B.n253 B.n250 10.6151
R1285 B.n254 B.n253 10.6151
R1286 B.n257 B.n254 10.6151
R1287 B.n258 B.n257 10.6151
R1288 B.n261 B.n258 10.6151
R1289 B.n262 B.n261 10.6151
R1290 B.n265 B.n262 10.6151
R1291 B.n266 B.n265 10.6151
R1292 B.n269 B.n266 10.6151
R1293 B.n270 B.n269 10.6151
R1294 B.n273 B.n270 10.6151
R1295 B.n274 B.n273 10.6151
R1296 B.n695 B.n274 10.6151
R1297 B.n767 B.n0 8.11757
R1298 B.n767 B.n1 8.11757
R1299 B.n472 B.n382 6.5566
R1300 B.n456 B.n455 6.5566
R1301 B.n186 B.n185 6.5566
R1302 B.n202 B.n108 6.5566
R1303 B.n475 B.n382 4.05904
R1304 B.n455 B.n454 4.05904
R1305 B.n185 B.n184 4.05904
R1306 B.n205 B.n108 4.05904
R1307 B.n308 B.t1 0.707668
R1308 B.t0 B.n730 0.707668
R1309 VN.n2 VN.t5 165.827
R1310 VN.n14 VN.t3 165.827
R1311 VN.n21 VN.n12 161.3
R1312 VN.n20 VN.n19 161.3
R1313 VN.n18 VN.n13 161.3
R1314 VN.n17 VN.n16 161.3
R1315 VN.n9 VN.n0 161.3
R1316 VN.n8 VN.n7 161.3
R1317 VN.n6 VN.n1 161.3
R1318 VN.n5 VN.n4 161.3
R1319 VN.n3 VN.t1 135.381
R1320 VN.n10 VN.t2 135.381
R1321 VN.n15 VN.t0 135.381
R1322 VN.n22 VN.t4 135.381
R1323 VN.n11 VN.n10 90.7429
R1324 VN.n23 VN.n22 90.7429
R1325 VN.n3 VN.n2 57.7341
R1326 VN.n15 VN.n14 57.7341
R1327 VN.n8 VN.n1 56.5617
R1328 VN.n20 VN.n13 56.5617
R1329 VN VN.n23 44.6194
R1330 VN.n4 VN.n1 24.5923
R1331 VN.n9 VN.n8 24.5923
R1332 VN.n16 VN.n13 24.5923
R1333 VN.n21 VN.n20 24.5923
R1334 VN.n10 VN.n9 20.1658
R1335 VN.n22 VN.n21 20.1658
R1336 VN.n17 VN.n14 13.2724
R1337 VN.n5 VN.n2 13.2724
R1338 VN.n4 VN.n3 12.2964
R1339 VN.n16 VN.n15 12.2964
R1340 VN.n23 VN.n12 0.278335
R1341 VN.n11 VN.n0 0.278335
R1342 VN.n19 VN.n12 0.189894
R1343 VN.n19 VN.n18 0.189894
R1344 VN.n18 VN.n17 0.189894
R1345 VN.n6 VN.n5 0.189894
R1346 VN.n7 VN.n6 0.189894
R1347 VN.n7 VN.n0 0.189894
R1348 VN VN.n11 0.153485
R1349 VDD2.n1 VDD2.t5 64.9743
R1350 VDD2.n2 VDD2.t0 63.6333
R1351 VDD2.n1 VDD2.n0 62.1172
R1352 VDD2 VDD2.n3 62.1144
R1353 VDD2.n2 VDD2.n1 38.6291
R1354 VDD2.n3 VDD2.t1 1.92657
R1355 VDD2.n3 VDD2.t4 1.92657
R1356 VDD2.n0 VDD2.t2 1.92657
R1357 VDD2.n0 VDD2.t3 1.92657
R1358 VDD2 VDD2.n2 1.45524
R1359 VTAIL.n7 VTAIL.t8 46.9545
R1360 VTAIL.n11 VTAIL.t9 46.9543
R1361 VTAIL.n2 VTAIL.t2 46.9543
R1362 VTAIL.n10 VTAIL.t0 46.9543
R1363 VTAIL.n9 VTAIL.n8 45.0285
R1364 VTAIL.n6 VTAIL.n5 45.0285
R1365 VTAIL.n1 VTAIL.n0 45.0282
R1366 VTAIL.n4 VTAIL.n3 45.0282
R1367 VTAIL.n6 VTAIL.n4 24.9531
R1368 VTAIL.n11 VTAIL.n10 23.091
R1369 VTAIL.n0 VTAIL.t6 1.92657
R1370 VTAIL.n0 VTAIL.t10 1.92657
R1371 VTAIL.n3 VTAIL.t4 1.92657
R1372 VTAIL.n3 VTAIL.t1 1.92657
R1373 VTAIL.n8 VTAIL.t5 1.92657
R1374 VTAIL.n8 VTAIL.t3 1.92657
R1375 VTAIL.n5 VTAIL.t7 1.92657
R1376 VTAIL.n5 VTAIL.t11 1.92657
R1377 VTAIL.n7 VTAIL.n6 1.86257
R1378 VTAIL.n10 VTAIL.n9 1.86257
R1379 VTAIL.n4 VTAIL.n2 1.86257
R1380 VTAIL.n9 VTAIL.n7 1.40136
R1381 VTAIL.n2 VTAIL.n1 1.40136
R1382 VTAIL VTAIL.n11 1.33886
R1383 VTAIL VTAIL.n1 0.524207
R1384 VP.n6 VP.t1 165.827
R1385 VP.n9 VP.n8 161.3
R1386 VP.n10 VP.n5 161.3
R1387 VP.n12 VP.n11 161.3
R1388 VP.n13 VP.n4 161.3
R1389 VP.n30 VP.n0 161.3
R1390 VP.n29 VP.n28 161.3
R1391 VP.n27 VP.n1 161.3
R1392 VP.n26 VP.n25 161.3
R1393 VP.n23 VP.n2 161.3
R1394 VP.n22 VP.n21 161.3
R1395 VP.n20 VP.n3 161.3
R1396 VP.n19 VP.n18 161.3
R1397 VP.n17 VP.t2 135.381
R1398 VP.n24 VP.t5 135.381
R1399 VP.n31 VP.t3 135.381
R1400 VP.n14 VP.t0 135.381
R1401 VP.n7 VP.t4 135.381
R1402 VP.n17 VP.n16 90.7429
R1403 VP.n32 VP.n31 90.7429
R1404 VP.n15 VP.n14 90.7429
R1405 VP.n7 VP.n6 57.7341
R1406 VP.n22 VP.n3 56.5617
R1407 VP.n29 VP.n1 56.5617
R1408 VP.n12 VP.n5 56.5617
R1409 VP.n16 VP.n15 44.3406
R1410 VP.n18 VP.n3 24.5923
R1411 VP.n23 VP.n22 24.5923
R1412 VP.n25 VP.n1 24.5923
R1413 VP.n30 VP.n29 24.5923
R1414 VP.n13 VP.n12 24.5923
R1415 VP.n8 VP.n5 24.5923
R1416 VP.n18 VP.n17 20.1658
R1417 VP.n31 VP.n30 20.1658
R1418 VP.n14 VP.n13 20.1658
R1419 VP.n9 VP.n6 13.2724
R1420 VP.n24 VP.n23 12.2964
R1421 VP.n25 VP.n24 12.2964
R1422 VP.n8 VP.n7 12.2964
R1423 VP.n15 VP.n4 0.278335
R1424 VP.n19 VP.n16 0.278335
R1425 VP.n32 VP.n0 0.278335
R1426 VP.n10 VP.n9 0.189894
R1427 VP.n11 VP.n10 0.189894
R1428 VP.n11 VP.n4 0.189894
R1429 VP.n20 VP.n19 0.189894
R1430 VP.n21 VP.n20 0.189894
R1431 VP.n21 VP.n2 0.189894
R1432 VP.n26 VP.n2 0.189894
R1433 VP.n27 VP.n26 0.189894
R1434 VP.n28 VP.n27 0.189894
R1435 VP.n28 VP.n0 0.189894
R1436 VP VP.n32 0.153485
R1437 VDD1 VDD1.t4 65.088
R1438 VDD1.n1 VDD1.t3 64.9743
R1439 VDD1.n1 VDD1.n0 62.1172
R1440 VDD1.n3 VDD1.n2 61.7071
R1441 VDD1.n3 VDD1.n1 40.1431
R1442 VDD1.n2 VDD1.t1 1.92657
R1443 VDD1.n2 VDD1.t5 1.92657
R1444 VDD1.n0 VDD1.t0 1.92657
R1445 VDD1.n0 VDD1.t2 1.92657
R1446 VDD1 VDD1.n3 0.407828
C0 VDD2 VP 0.393332f
C1 VN VTAIL 5.42943f
C2 VDD2 VTAIL 7.10854f
C3 VN VDD1 0.15009f
C4 VDD2 VDD1 1.13232f
C5 VP VTAIL 5.443759f
C6 VP VDD1 5.61542f
C7 VTAIL VDD1 7.06337f
C8 VDD2 VN 5.37528f
C9 VP VN 5.86002f
C10 VDD2 B 5.064343f
C11 VDD1 B 5.350252f
C12 VTAIL B 6.620835f
C13 VN B 10.550051f
C14 VP B 9.07796f
C15 VDD1.t4 B 2.00174f
C16 VDD1.t3 B 2.00098f
C17 VDD1.t0 B 0.177616f
C18 VDD1.t2 B 0.177616f
C19 VDD1.n0 B 1.56857f
C20 VDD1.n1 B 2.24792f
C21 VDD1.t1 B 0.177616f
C22 VDD1.t5 B 0.177616f
C23 VDD1.n2 B 1.56625f
C24 VDD1.n3 B 2.13323f
C25 VP.n0 B 0.039331f
C26 VP.t3 B 1.5219f
C27 VP.n1 B 0.049972f
C28 VP.n2 B 0.029834f
C29 VP.t5 B 1.5219f
C30 VP.n3 B 0.036765f
C31 VP.n4 B 0.039331f
C32 VP.t0 B 1.5219f
C33 VP.n5 B 0.049972f
C34 VP.t1 B 1.648f
C35 VP.n6 B 0.627022f
C36 VP.t4 B 1.5219f
C37 VP.n7 B 0.618204f
C38 VP.n8 B 0.041669f
C39 VP.n9 B 0.218758f
C40 VP.n10 B 0.029834f
C41 VP.n11 B 0.029834f
C42 VP.n12 B 0.036765f
C43 VP.n13 B 0.050409f
C44 VP.n14 B 0.635362f
C45 VP.n15 B 1.36891f
C46 VP.n16 B 1.39317f
C47 VP.t2 B 1.5219f
C48 VP.n17 B 0.635362f
C49 VP.n18 B 0.050409f
C50 VP.n19 B 0.039331f
C51 VP.n20 B 0.029834f
C52 VP.n21 B 0.029834f
C53 VP.n22 B 0.049972f
C54 VP.n23 B 0.041669f
C55 VP.n24 B 0.551613f
C56 VP.n25 B 0.041669f
C57 VP.n26 B 0.029834f
C58 VP.n27 B 0.029834f
C59 VP.n28 B 0.029834f
C60 VP.n29 B 0.036765f
C61 VP.n30 B 0.050409f
C62 VP.n31 B 0.635362f
C63 VP.n32 B 0.035169f
C64 VTAIL.t6 B 0.193036f
C65 VTAIL.t10 B 0.193036f
C66 VTAIL.n0 B 1.63167f
C67 VTAIL.n1 B 0.380618f
C68 VTAIL.t2 B 2.07752f
C69 VTAIL.n2 B 0.563703f
C70 VTAIL.t4 B 0.193036f
C71 VTAIL.t1 B 0.193036f
C72 VTAIL.n3 B 1.63167f
C73 VTAIL.n4 B 1.66232f
C74 VTAIL.t7 B 0.193036f
C75 VTAIL.t11 B 0.193036f
C76 VTAIL.n5 B 1.63168f
C77 VTAIL.n6 B 1.66231f
C78 VTAIL.t8 B 2.07753f
C79 VTAIL.n7 B 0.563697f
C80 VTAIL.t5 B 0.193036f
C81 VTAIL.t3 B 0.193036f
C82 VTAIL.n8 B 1.63168f
C83 VTAIL.n9 B 0.483088f
C84 VTAIL.t0 B 2.07752f
C85 VTAIL.n10 B 1.60035f
C86 VTAIL.t9 B 2.07752f
C87 VTAIL.n11 B 1.56025f
C88 VDD2.t5 B 1.98208f
C89 VDD2.t2 B 0.175938f
C90 VDD2.t3 B 0.175938f
C91 VDD2.n0 B 1.55374f
C92 VDD2.n1 B 2.13719f
C93 VDD2.t0 B 1.97513f
C94 VDD2.n2 B 2.12187f
C95 VDD2.t1 B 0.175938f
C96 VDD2.t4 B 0.175938f
C97 VDD2.n3 B 1.55371f
C98 VN.n0 B 0.03877f
C99 VN.t2 B 1.50017f
C100 VN.n1 B 0.049259f
C101 VN.t5 B 1.62447f
C102 VN.n2 B 0.618068f
C103 VN.t1 B 1.50017f
C104 VN.n3 B 0.609375f
C105 VN.n4 B 0.041074f
C106 VN.n5 B 0.215634f
C107 VN.n6 B 0.029408f
C108 VN.n7 B 0.029408f
C109 VN.n8 B 0.03624f
C110 VN.n9 B 0.049689f
C111 VN.n10 B 0.626289f
C112 VN.n11 B 0.034667f
C113 VN.n12 B 0.03877f
C114 VN.t4 B 1.50017f
C115 VN.n13 B 0.049259f
C116 VN.t3 B 1.62447f
C117 VN.n14 B 0.618068f
C118 VN.t0 B 1.50017f
C119 VN.n15 B 0.609375f
C120 VN.n16 B 0.041074f
C121 VN.n17 B 0.215634f
C122 VN.n18 B 0.029408f
C123 VN.n19 B 0.029408f
C124 VN.n20 B 0.03624f
C125 VN.n21 B 0.049689f
C126 VN.n22 B 0.626289f
C127 VN.n23 B 1.36549f
.ends

