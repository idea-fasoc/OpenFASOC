* NGSPICE file created from diff_pair_sample_0686.ext - technology: sky130A

.subckt diff_pair_sample_0686 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t7 VN.t0 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=3.9975 ps=21.28 w=10.25 l=1.39
X1 VDD1.t7 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=3.9975 ps=21.28 w=10.25 l=1.39
X2 VTAIL.t15 VN.t1 VDD2.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=1.69125 ps=10.58 w=10.25 l=1.39
X3 VDD1.t6 VP.t1 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=3.9975 ps=21.28 w=10.25 l=1.39
X4 VTAIL.t14 VN.t2 VDD2.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
X5 VDD2.t4 VN.t3 VTAIL.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
X6 VDD1.t5 VP.t2 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
X7 VTAIL.t0 VP.t3 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
X8 VDD1.t3 VP.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
X9 B.t21 B.t19 B.t20 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=0 ps=0 w=10.25 l=1.39
X10 VDD2.t3 VN.t4 VTAIL.t12 B.t5 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=3.9975 ps=21.28 w=10.25 l=1.39
X11 VTAIL.t13 VN.t5 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=1.69125 ps=10.58 w=10.25 l=1.39
X12 B.t18 B.t16 B.t17 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=0 ps=0 w=10.25 l=1.39
X13 VTAIL.t4 VP.t5 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=1.69125 ps=10.58 w=10.25 l=1.39
X14 VTAIL.t9 VN.t6 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
X15 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=0 ps=0 w=10.25 l=1.39
X16 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=0 ps=0 w=10.25 l=1.39
X17 VTAIL.t3 VP.t6 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
X18 VTAIL.t2 VP.t7 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=3.9975 pd=21.28 as=1.69125 ps=10.58 w=10.25 l=1.39
X19 VDD2.t0 VN.t7 VTAIL.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.69125 pd=10.58 as=1.69125 ps=10.58 w=10.25 l=1.39
R0 VN.n5 VN.t5 209.338
R1 VN.n25 VN.t4 209.338
R2 VN.n4 VN.t7 177.716
R3 VN.n10 VN.t6 177.716
R4 VN.n17 VN.t0 177.716
R5 VN.n24 VN.t2 177.716
R6 VN.n22 VN.t3 177.716
R7 VN.n36 VN.t1 177.716
R8 VN.n18 VN.n17 169.619
R9 VN.n37 VN.n36 169.619
R10 VN.n35 VN.n19 161.3
R11 VN.n34 VN.n33 161.3
R12 VN.n32 VN.n20 161.3
R13 VN.n31 VN.n30 161.3
R14 VN.n29 VN.n21 161.3
R15 VN.n28 VN.n27 161.3
R16 VN.n26 VN.n23 161.3
R17 VN.n16 VN.n0 161.3
R18 VN.n15 VN.n14 161.3
R19 VN.n13 VN.n1 161.3
R20 VN.n12 VN.n11 161.3
R21 VN.n9 VN.n2 161.3
R22 VN.n8 VN.n7 161.3
R23 VN.n6 VN.n3 161.3
R24 VN.n5 VN.n4 59.48
R25 VN.n25 VN.n24 59.48
R26 VN.n9 VN.n8 56.5193
R27 VN.n29 VN.n28 56.5193
R28 VN VN.n37 44.2827
R29 VN.n15 VN.n1 43.4072
R30 VN.n34 VN.n20 43.4072
R31 VN.n16 VN.n15 37.5796
R32 VN.n35 VN.n34 37.5796
R33 VN.n26 VN.n25 26.5029
R34 VN.n6 VN.n5 26.5029
R35 VN.n8 VN.n3 24.4675
R36 VN.n11 VN.n9 24.4675
R37 VN.n28 VN.n23 24.4675
R38 VN.n30 VN.n29 24.4675
R39 VN.n10 VN.n1 19.0848
R40 VN.n22 VN.n20 19.0848
R41 VN.n17 VN.n16 16.1487
R42 VN.n36 VN.n35 16.1487
R43 VN.n4 VN.n3 5.38324
R44 VN.n11 VN.n10 5.38324
R45 VN.n24 VN.n23 5.38324
R46 VN.n30 VN.n22 5.38324
R47 VN.n37 VN.n19 0.189894
R48 VN.n33 VN.n19 0.189894
R49 VN.n33 VN.n32 0.189894
R50 VN.n32 VN.n31 0.189894
R51 VN.n31 VN.n21 0.189894
R52 VN.n27 VN.n21 0.189894
R53 VN.n27 VN.n26 0.189894
R54 VN.n7 VN.n6 0.189894
R55 VN.n7 VN.n2 0.189894
R56 VN.n12 VN.n2 0.189894
R57 VN.n13 VN.n12 0.189894
R58 VN.n14 VN.n13 0.189894
R59 VN.n14 VN.n0 0.189894
R60 VN.n18 VN.n0 0.189894
R61 VN VN.n18 0.0516364
R62 VTAIL.n11 VTAIL.t4 46.3783
R63 VTAIL.n10 VTAIL.t12 46.3783
R64 VTAIL.n7 VTAIL.t15 46.3783
R65 VTAIL.n15 VTAIL.t10 46.3781
R66 VTAIL.n2 VTAIL.t13 46.3781
R67 VTAIL.n3 VTAIL.t5 46.3781
R68 VTAIL.n6 VTAIL.t2 46.3781
R69 VTAIL.n14 VTAIL.t1 46.3781
R70 VTAIL.n13 VTAIL.n12 44.4466
R71 VTAIL.n9 VTAIL.n8 44.4466
R72 VTAIL.n1 VTAIL.n0 44.4464
R73 VTAIL.n5 VTAIL.n4 44.4464
R74 VTAIL.n15 VTAIL.n14 22.6858
R75 VTAIL.n7 VTAIL.n6 22.6858
R76 VTAIL.n0 VTAIL.t8 1.93221
R77 VTAIL.n0 VTAIL.t9 1.93221
R78 VTAIL.n4 VTAIL.t7 1.93221
R79 VTAIL.n4 VTAIL.t3 1.93221
R80 VTAIL.n12 VTAIL.t6 1.93221
R81 VTAIL.n12 VTAIL.t0 1.93221
R82 VTAIL.n8 VTAIL.t11 1.93221
R83 VTAIL.n8 VTAIL.t14 1.93221
R84 VTAIL.n9 VTAIL.n7 1.48326
R85 VTAIL.n10 VTAIL.n9 1.48326
R86 VTAIL.n13 VTAIL.n11 1.48326
R87 VTAIL.n14 VTAIL.n13 1.48326
R88 VTAIL.n6 VTAIL.n5 1.48326
R89 VTAIL.n5 VTAIL.n3 1.48326
R90 VTAIL.n2 VTAIL.n1 1.48326
R91 VTAIL VTAIL.n15 1.42507
R92 VTAIL.n11 VTAIL.n10 0.470328
R93 VTAIL.n3 VTAIL.n2 0.470328
R94 VTAIL VTAIL.n1 0.0586897
R95 VDD2.n2 VDD2.n1 61.8112
R96 VDD2.n2 VDD2.n0 61.8112
R97 VDD2 VDD2.n5 61.8084
R98 VDD2.n4 VDD2.n3 61.1254
R99 VDD2.n4 VDD2.n2 39.2239
R100 VDD2.n5 VDD2.t5 1.93221
R101 VDD2.n5 VDD2.t3 1.93221
R102 VDD2.n3 VDD2.t6 1.93221
R103 VDD2.n3 VDD2.t4 1.93221
R104 VDD2.n1 VDD2.t1 1.93221
R105 VDD2.n1 VDD2.t7 1.93221
R106 VDD2.n0 VDD2.t2 1.93221
R107 VDD2.n0 VDD2.t0 1.93221
R108 VDD2 VDD2.n4 0.800069
R109 B.n690 B.n689 585
R110 B.n270 B.n103 585
R111 B.n269 B.n268 585
R112 B.n267 B.n266 585
R113 B.n265 B.n264 585
R114 B.n263 B.n262 585
R115 B.n261 B.n260 585
R116 B.n259 B.n258 585
R117 B.n257 B.n256 585
R118 B.n255 B.n254 585
R119 B.n253 B.n252 585
R120 B.n251 B.n250 585
R121 B.n249 B.n248 585
R122 B.n247 B.n246 585
R123 B.n245 B.n244 585
R124 B.n243 B.n242 585
R125 B.n241 B.n240 585
R126 B.n239 B.n238 585
R127 B.n237 B.n236 585
R128 B.n235 B.n234 585
R129 B.n233 B.n232 585
R130 B.n231 B.n230 585
R131 B.n229 B.n228 585
R132 B.n227 B.n226 585
R133 B.n225 B.n224 585
R134 B.n223 B.n222 585
R135 B.n221 B.n220 585
R136 B.n219 B.n218 585
R137 B.n217 B.n216 585
R138 B.n215 B.n214 585
R139 B.n213 B.n212 585
R140 B.n211 B.n210 585
R141 B.n209 B.n208 585
R142 B.n207 B.n206 585
R143 B.n205 B.n204 585
R144 B.n203 B.n202 585
R145 B.n201 B.n200 585
R146 B.n199 B.n198 585
R147 B.n197 B.n196 585
R148 B.n195 B.n194 585
R149 B.n193 B.n192 585
R150 B.n191 B.n190 585
R151 B.n189 B.n188 585
R152 B.n187 B.n186 585
R153 B.n185 B.n184 585
R154 B.n183 B.n182 585
R155 B.n181 B.n180 585
R156 B.n179 B.n178 585
R157 B.n177 B.n176 585
R158 B.n175 B.n174 585
R159 B.n173 B.n172 585
R160 B.n171 B.n170 585
R161 B.n169 B.n168 585
R162 B.n167 B.n166 585
R163 B.n165 B.n164 585
R164 B.n163 B.n162 585
R165 B.n161 B.n160 585
R166 B.n159 B.n158 585
R167 B.n157 B.n156 585
R168 B.n155 B.n154 585
R169 B.n153 B.n152 585
R170 B.n151 B.n150 585
R171 B.n149 B.n148 585
R172 B.n147 B.n146 585
R173 B.n145 B.n144 585
R174 B.n143 B.n142 585
R175 B.n141 B.n140 585
R176 B.n139 B.n138 585
R177 B.n137 B.n136 585
R178 B.n135 B.n134 585
R179 B.n133 B.n132 585
R180 B.n131 B.n130 585
R181 B.n129 B.n128 585
R182 B.n127 B.n126 585
R183 B.n125 B.n124 585
R184 B.n123 B.n122 585
R185 B.n121 B.n120 585
R186 B.n119 B.n118 585
R187 B.n117 B.n116 585
R188 B.n115 B.n114 585
R189 B.n113 B.n112 585
R190 B.n111 B.n110 585
R191 B.n688 B.n62 585
R192 B.n693 B.n62 585
R193 B.n687 B.n61 585
R194 B.n694 B.n61 585
R195 B.n686 B.n685 585
R196 B.n685 B.n57 585
R197 B.n684 B.n56 585
R198 B.n700 B.n56 585
R199 B.n683 B.n55 585
R200 B.n701 B.n55 585
R201 B.n682 B.n54 585
R202 B.n702 B.n54 585
R203 B.n681 B.n680 585
R204 B.n680 B.n50 585
R205 B.n679 B.n49 585
R206 B.n708 B.n49 585
R207 B.n678 B.n48 585
R208 B.n709 B.n48 585
R209 B.n677 B.n47 585
R210 B.n710 B.n47 585
R211 B.n676 B.n675 585
R212 B.n675 B.n43 585
R213 B.n674 B.n42 585
R214 B.n716 B.n42 585
R215 B.n673 B.n41 585
R216 B.n717 B.n41 585
R217 B.n672 B.n40 585
R218 B.n718 B.n40 585
R219 B.n671 B.n670 585
R220 B.n670 B.n39 585
R221 B.n669 B.n35 585
R222 B.n724 B.n35 585
R223 B.n668 B.n34 585
R224 B.n725 B.n34 585
R225 B.n667 B.n33 585
R226 B.n726 B.n33 585
R227 B.n666 B.n665 585
R228 B.n665 B.n29 585
R229 B.n664 B.n28 585
R230 B.n732 B.n28 585
R231 B.n663 B.n27 585
R232 B.n733 B.n27 585
R233 B.n662 B.n26 585
R234 B.n734 B.n26 585
R235 B.n661 B.n660 585
R236 B.n660 B.n22 585
R237 B.n659 B.n21 585
R238 B.n740 B.n21 585
R239 B.n658 B.n20 585
R240 B.n741 B.n20 585
R241 B.n657 B.n19 585
R242 B.n742 B.n19 585
R243 B.n656 B.n655 585
R244 B.n655 B.n15 585
R245 B.n654 B.n14 585
R246 B.n748 B.n14 585
R247 B.n653 B.n13 585
R248 B.n749 B.n13 585
R249 B.n652 B.n12 585
R250 B.n750 B.n12 585
R251 B.n651 B.n650 585
R252 B.n650 B.n649 585
R253 B.n648 B.n647 585
R254 B.n648 B.n8 585
R255 B.n646 B.n7 585
R256 B.n757 B.n7 585
R257 B.n645 B.n6 585
R258 B.n758 B.n6 585
R259 B.n644 B.n5 585
R260 B.n759 B.n5 585
R261 B.n643 B.n642 585
R262 B.n642 B.n4 585
R263 B.n641 B.n271 585
R264 B.n641 B.n640 585
R265 B.n631 B.n272 585
R266 B.n273 B.n272 585
R267 B.n633 B.n632 585
R268 B.n634 B.n633 585
R269 B.n630 B.n278 585
R270 B.n278 B.n277 585
R271 B.n629 B.n628 585
R272 B.n628 B.n627 585
R273 B.n280 B.n279 585
R274 B.n281 B.n280 585
R275 B.n620 B.n619 585
R276 B.n621 B.n620 585
R277 B.n618 B.n285 585
R278 B.n289 B.n285 585
R279 B.n617 B.n616 585
R280 B.n616 B.n615 585
R281 B.n287 B.n286 585
R282 B.n288 B.n287 585
R283 B.n608 B.n607 585
R284 B.n609 B.n608 585
R285 B.n606 B.n294 585
R286 B.n294 B.n293 585
R287 B.n605 B.n604 585
R288 B.n604 B.n603 585
R289 B.n296 B.n295 585
R290 B.n297 B.n296 585
R291 B.n596 B.n595 585
R292 B.n597 B.n596 585
R293 B.n594 B.n302 585
R294 B.n302 B.n301 585
R295 B.n593 B.n592 585
R296 B.n592 B.n591 585
R297 B.n304 B.n303 585
R298 B.n584 B.n304 585
R299 B.n583 B.n582 585
R300 B.n585 B.n583 585
R301 B.n581 B.n309 585
R302 B.n309 B.n308 585
R303 B.n580 B.n579 585
R304 B.n579 B.n578 585
R305 B.n311 B.n310 585
R306 B.n312 B.n311 585
R307 B.n571 B.n570 585
R308 B.n572 B.n571 585
R309 B.n569 B.n317 585
R310 B.n317 B.n316 585
R311 B.n568 B.n567 585
R312 B.n567 B.n566 585
R313 B.n319 B.n318 585
R314 B.n320 B.n319 585
R315 B.n559 B.n558 585
R316 B.n560 B.n559 585
R317 B.n557 B.n325 585
R318 B.n325 B.n324 585
R319 B.n556 B.n555 585
R320 B.n555 B.n554 585
R321 B.n327 B.n326 585
R322 B.n328 B.n327 585
R323 B.n547 B.n546 585
R324 B.n548 B.n547 585
R325 B.n545 B.n333 585
R326 B.n333 B.n332 585
R327 B.n540 B.n539 585
R328 B.n538 B.n376 585
R329 B.n537 B.n375 585
R330 B.n542 B.n375 585
R331 B.n536 B.n535 585
R332 B.n534 B.n533 585
R333 B.n532 B.n531 585
R334 B.n530 B.n529 585
R335 B.n528 B.n527 585
R336 B.n526 B.n525 585
R337 B.n524 B.n523 585
R338 B.n522 B.n521 585
R339 B.n520 B.n519 585
R340 B.n518 B.n517 585
R341 B.n516 B.n515 585
R342 B.n514 B.n513 585
R343 B.n512 B.n511 585
R344 B.n510 B.n509 585
R345 B.n508 B.n507 585
R346 B.n506 B.n505 585
R347 B.n504 B.n503 585
R348 B.n502 B.n501 585
R349 B.n500 B.n499 585
R350 B.n498 B.n497 585
R351 B.n496 B.n495 585
R352 B.n494 B.n493 585
R353 B.n492 B.n491 585
R354 B.n490 B.n489 585
R355 B.n488 B.n487 585
R356 B.n486 B.n485 585
R357 B.n484 B.n483 585
R358 B.n482 B.n481 585
R359 B.n480 B.n479 585
R360 B.n478 B.n477 585
R361 B.n476 B.n475 585
R362 B.n474 B.n473 585
R363 B.n472 B.n471 585
R364 B.n469 B.n468 585
R365 B.n467 B.n466 585
R366 B.n465 B.n464 585
R367 B.n463 B.n462 585
R368 B.n461 B.n460 585
R369 B.n459 B.n458 585
R370 B.n457 B.n456 585
R371 B.n455 B.n454 585
R372 B.n453 B.n452 585
R373 B.n451 B.n450 585
R374 B.n448 B.n447 585
R375 B.n446 B.n445 585
R376 B.n444 B.n443 585
R377 B.n442 B.n441 585
R378 B.n440 B.n439 585
R379 B.n438 B.n437 585
R380 B.n436 B.n435 585
R381 B.n434 B.n433 585
R382 B.n432 B.n431 585
R383 B.n430 B.n429 585
R384 B.n428 B.n427 585
R385 B.n426 B.n425 585
R386 B.n424 B.n423 585
R387 B.n422 B.n421 585
R388 B.n420 B.n419 585
R389 B.n418 B.n417 585
R390 B.n416 B.n415 585
R391 B.n414 B.n413 585
R392 B.n412 B.n411 585
R393 B.n410 B.n409 585
R394 B.n408 B.n407 585
R395 B.n406 B.n405 585
R396 B.n404 B.n403 585
R397 B.n402 B.n401 585
R398 B.n400 B.n399 585
R399 B.n398 B.n397 585
R400 B.n396 B.n395 585
R401 B.n394 B.n393 585
R402 B.n392 B.n391 585
R403 B.n390 B.n389 585
R404 B.n388 B.n387 585
R405 B.n386 B.n385 585
R406 B.n384 B.n383 585
R407 B.n382 B.n381 585
R408 B.n335 B.n334 585
R409 B.n544 B.n543 585
R410 B.n543 B.n542 585
R411 B.n331 B.n330 585
R412 B.n332 B.n331 585
R413 B.n550 B.n549 585
R414 B.n549 B.n548 585
R415 B.n551 B.n329 585
R416 B.n329 B.n328 585
R417 B.n553 B.n552 585
R418 B.n554 B.n553 585
R419 B.n323 B.n322 585
R420 B.n324 B.n323 585
R421 B.n562 B.n561 585
R422 B.n561 B.n560 585
R423 B.n563 B.n321 585
R424 B.n321 B.n320 585
R425 B.n565 B.n564 585
R426 B.n566 B.n565 585
R427 B.n315 B.n314 585
R428 B.n316 B.n315 585
R429 B.n574 B.n573 585
R430 B.n573 B.n572 585
R431 B.n575 B.n313 585
R432 B.n313 B.n312 585
R433 B.n577 B.n576 585
R434 B.n578 B.n577 585
R435 B.n307 B.n306 585
R436 B.n308 B.n307 585
R437 B.n587 B.n586 585
R438 B.n586 B.n585 585
R439 B.n588 B.n305 585
R440 B.n584 B.n305 585
R441 B.n590 B.n589 585
R442 B.n591 B.n590 585
R443 B.n300 B.n299 585
R444 B.n301 B.n300 585
R445 B.n599 B.n598 585
R446 B.n598 B.n597 585
R447 B.n600 B.n298 585
R448 B.n298 B.n297 585
R449 B.n602 B.n601 585
R450 B.n603 B.n602 585
R451 B.n292 B.n291 585
R452 B.n293 B.n292 585
R453 B.n611 B.n610 585
R454 B.n610 B.n609 585
R455 B.n612 B.n290 585
R456 B.n290 B.n288 585
R457 B.n614 B.n613 585
R458 B.n615 B.n614 585
R459 B.n284 B.n283 585
R460 B.n289 B.n284 585
R461 B.n623 B.n622 585
R462 B.n622 B.n621 585
R463 B.n624 B.n282 585
R464 B.n282 B.n281 585
R465 B.n626 B.n625 585
R466 B.n627 B.n626 585
R467 B.n276 B.n275 585
R468 B.n277 B.n276 585
R469 B.n636 B.n635 585
R470 B.n635 B.n634 585
R471 B.n637 B.n274 585
R472 B.n274 B.n273 585
R473 B.n639 B.n638 585
R474 B.n640 B.n639 585
R475 B.n3 B.n0 585
R476 B.n4 B.n3 585
R477 B.n756 B.n1 585
R478 B.n757 B.n756 585
R479 B.n755 B.n754 585
R480 B.n755 B.n8 585
R481 B.n753 B.n9 585
R482 B.n649 B.n9 585
R483 B.n752 B.n751 585
R484 B.n751 B.n750 585
R485 B.n11 B.n10 585
R486 B.n749 B.n11 585
R487 B.n747 B.n746 585
R488 B.n748 B.n747 585
R489 B.n745 B.n16 585
R490 B.n16 B.n15 585
R491 B.n744 B.n743 585
R492 B.n743 B.n742 585
R493 B.n18 B.n17 585
R494 B.n741 B.n18 585
R495 B.n739 B.n738 585
R496 B.n740 B.n739 585
R497 B.n737 B.n23 585
R498 B.n23 B.n22 585
R499 B.n736 B.n735 585
R500 B.n735 B.n734 585
R501 B.n25 B.n24 585
R502 B.n733 B.n25 585
R503 B.n731 B.n730 585
R504 B.n732 B.n731 585
R505 B.n729 B.n30 585
R506 B.n30 B.n29 585
R507 B.n728 B.n727 585
R508 B.n727 B.n726 585
R509 B.n32 B.n31 585
R510 B.n725 B.n32 585
R511 B.n723 B.n722 585
R512 B.n724 B.n723 585
R513 B.n721 B.n36 585
R514 B.n39 B.n36 585
R515 B.n720 B.n719 585
R516 B.n719 B.n718 585
R517 B.n38 B.n37 585
R518 B.n717 B.n38 585
R519 B.n715 B.n714 585
R520 B.n716 B.n715 585
R521 B.n713 B.n44 585
R522 B.n44 B.n43 585
R523 B.n712 B.n711 585
R524 B.n711 B.n710 585
R525 B.n46 B.n45 585
R526 B.n709 B.n46 585
R527 B.n707 B.n706 585
R528 B.n708 B.n707 585
R529 B.n705 B.n51 585
R530 B.n51 B.n50 585
R531 B.n704 B.n703 585
R532 B.n703 B.n702 585
R533 B.n53 B.n52 585
R534 B.n701 B.n53 585
R535 B.n699 B.n698 585
R536 B.n700 B.n699 585
R537 B.n697 B.n58 585
R538 B.n58 B.n57 585
R539 B.n696 B.n695 585
R540 B.n695 B.n694 585
R541 B.n60 B.n59 585
R542 B.n693 B.n60 585
R543 B.n760 B.n759 585
R544 B.n758 B.n2 585
R545 B.n110 B.n60 526.135
R546 B.n690 B.n62 526.135
R547 B.n543 B.n333 526.135
R548 B.n540 B.n331 526.135
R549 B.n107 B.t19 382.721
R550 B.n104 B.t8 382.721
R551 B.n379 B.t16 382.721
R552 B.n377 B.t12 382.721
R553 B.n692 B.n691 256.663
R554 B.n692 B.n102 256.663
R555 B.n692 B.n101 256.663
R556 B.n692 B.n100 256.663
R557 B.n692 B.n99 256.663
R558 B.n692 B.n98 256.663
R559 B.n692 B.n97 256.663
R560 B.n692 B.n96 256.663
R561 B.n692 B.n95 256.663
R562 B.n692 B.n94 256.663
R563 B.n692 B.n93 256.663
R564 B.n692 B.n92 256.663
R565 B.n692 B.n91 256.663
R566 B.n692 B.n90 256.663
R567 B.n692 B.n89 256.663
R568 B.n692 B.n88 256.663
R569 B.n692 B.n87 256.663
R570 B.n692 B.n86 256.663
R571 B.n692 B.n85 256.663
R572 B.n692 B.n84 256.663
R573 B.n692 B.n83 256.663
R574 B.n692 B.n82 256.663
R575 B.n692 B.n81 256.663
R576 B.n692 B.n80 256.663
R577 B.n692 B.n79 256.663
R578 B.n692 B.n78 256.663
R579 B.n692 B.n77 256.663
R580 B.n692 B.n76 256.663
R581 B.n692 B.n75 256.663
R582 B.n692 B.n74 256.663
R583 B.n692 B.n73 256.663
R584 B.n692 B.n72 256.663
R585 B.n692 B.n71 256.663
R586 B.n692 B.n70 256.663
R587 B.n692 B.n69 256.663
R588 B.n692 B.n68 256.663
R589 B.n692 B.n67 256.663
R590 B.n692 B.n66 256.663
R591 B.n692 B.n65 256.663
R592 B.n692 B.n64 256.663
R593 B.n692 B.n63 256.663
R594 B.n542 B.n541 256.663
R595 B.n542 B.n336 256.663
R596 B.n542 B.n337 256.663
R597 B.n542 B.n338 256.663
R598 B.n542 B.n339 256.663
R599 B.n542 B.n340 256.663
R600 B.n542 B.n341 256.663
R601 B.n542 B.n342 256.663
R602 B.n542 B.n343 256.663
R603 B.n542 B.n344 256.663
R604 B.n542 B.n345 256.663
R605 B.n542 B.n346 256.663
R606 B.n542 B.n347 256.663
R607 B.n542 B.n348 256.663
R608 B.n542 B.n349 256.663
R609 B.n542 B.n350 256.663
R610 B.n542 B.n351 256.663
R611 B.n542 B.n352 256.663
R612 B.n542 B.n353 256.663
R613 B.n542 B.n354 256.663
R614 B.n542 B.n355 256.663
R615 B.n542 B.n356 256.663
R616 B.n542 B.n357 256.663
R617 B.n542 B.n358 256.663
R618 B.n542 B.n359 256.663
R619 B.n542 B.n360 256.663
R620 B.n542 B.n361 256.663
R621 B.n542 B.n362 256.663
R622 B.n542 B.n363 256.663
R623 B.n542 B.n364 256.663
R624 B.n542 B.n365 256.663
R625 B.n542 B.n366 256.663
R626 B.n542 B.n367 256.663
R627 B.n542 B.n368 256.663
R628 B.n542 B.n369 256.663
R629 B.n542 B.n370 256.663
R630 B.n542 B.n371 256.663
R631 B.n542 B.n372 256.663
R632 B.n542 B.n373 256.663
R633 B.n542 B.n374 256.663
R634 B.n762 B.n761 256.663
R635 B.n114 B.n113 163.367
R636 B.n118 B.n117 163.367
R637 B.n122 B.n121 163.367
R638 B.n126 B.n125 163.367
R639 B.n130 B.n129 163.367
R640 B.n134 B.n133 163.367
R641 B.n138 B.n137 163.367
R642 B.n142 B.n141 163.367
R643 B.n146 B.n145 163.367
R644 B.n150 B.n149 163.367
R645 B.n154 B.n153 163.367
R646 B.n158 B.n157 163.367
R647 B.n162 B.n161 163.367
R648 B.n166 B.n165 163.367
R649 B.n170 B.n169 163.367
R650 B.n174 B.n173 163.367
R651 B.n178 B.n177 163.367
R652 B.n182 B.n181 163.367
R653 B.n186 B.n185 163.367
R654 B.n190 B.n189 163.367
R655 B.n194 B.n193 163.367
R656 B.n198 B.n197 163.367
R657 B.n202 B.n201 163.367
R658 B.n206 B.n205 163.367
R659 B.n210 B.n209 163.367
R660 B.n214 B.n213 163.367
R661 B.n218 B.n217 163.367
R662 B.n222 B.n221 163.367
R663 B.n226 B.n225 163.367
R664 B.n230 B.n229 163.367
R665 B.n234 B.n233 163.367
R666 B.n238 B.n237 163.367
R667 B.n242 B.n241 163.367
R668 B.n246 B.n245 163.367
R669 B.n250 B.n249 163.367
R670 B.n254 B.n253 163.367
R671 B.n258 B.n257 163.367
R672 B.n262 B.n261 163.367
R673 B.n266 B.n265 163.367
R674 B.n268 B.n103 163.367
R675 B.n547 B.n333 163.367
R676 B.n547 B.n327 163.367
R677 B.n555 B.n327 163.367
R678 B.n555 B.n325 163.367
R679 B.n559 B.n325 163.367
R680 B.n559 B.n319 163.367
R681 B.n567 B.n319 163.367
R682 B.n567 B.n317 163.367
R683 B.n571 B.n317 163.367
R684 B.n571 B.n311 163.367
R685 B.n579 B.n311 163.367
R686 B.n579 B.n309 163.367
R687 B.n583 B.n309 163.367
R688 B.n583 B.n304 163.367
R689 B.n592 B.n304 163.367
R690 B.n592 B.n302 163.367
R691 B.n596 B.n302 163.367
R692 B.n596 B.n296 163.367
R693 B.n604 B.n296 163.367
R694 B.n604 B.n294 163.367
R695 B.n608 B.n294 163.367
R696 B.n608 B.n287 163.367
R697 B.n616 B.n287 163.367
R698 B.n616 B.n285 163.367
R699 B.n620 B.n285 163.367
R700 B.n620 B.n280 163.367
R701 B.n628 B.n280 163.367
R702 B.n628 B.n278 163.367
R703 B.n633 B.n278 163.367
R704 B.n633 B.n272 163.367
R705 B.n641 B.n272 163.367
R706 B.n642 B.n641 163.367
R707 B.n642 B.n5 163.367
R708 B.n6 B.n5 163.367
R709 B.n7 B.n6 163.367
R710 B.n648 B.n7 163.367
R711 B.n650 B.n648 163.367
R712 B.n650 B.n12 163.367
R713 B.n13 B.n12 163.367
R714 B.n14 B.n13 163.367
R715 B.n655 B.n14 163.367
R716 B.n655 B.n19 163.367
R717 B.n20 B.n19 163.367
R718 B.n21 B.n20 163.367
R719 B.n660 B.n21 163.367
R720 B.n660 B.n26 163.367
R721 B.n27 B.n26 163.367
R722 B.n28 B.n27 163.367
R723 B.n665 B.n28 163.367
R724 B.n665 B.n33 163.367
R725 B.n34 B.n33 163.367
R726 B.n35 B.n34 163.367
R727 B.n670 B.n35 163.367
R728 B.n670 B.n40 163.367
R729 B.n41 B.n40 163.367
R730 B.n42 B.n41 163.367
R731 B.n675 B.n42 163.367
R732 B.n675 B.n47 163.367
R733 B.n48 B.n47 163.367
R734 B.n49 B.n48 163.367
R735 B.n680 B.n49 163.367
R736 B.n680 B.n54 163.367
R737 B.n55 B.n54 163.367
R738 B.n56 B.n55 163.367
R739 B.n685 B.n56 163.367
R740 B.n685 B.n61 163.367
R741 B.n62 B.n61 163.367
R742 B.n376 B.n375 163.367
R743 B.n535 B.n375 163.367
R744 B.n533 B.n532 163.367
R745 B.n529 B.n528 163.367
R746 B.n525 B.n524 163.367
R747 B.n521 B.n520 163.367
R748 B.n517 B.n516 163.367
R749 B.n513 B.n512 163.367
R750 B.n509 B.n508 163.367
R751 B.n505 B.n504 163.367
R752 B.n501 B.n500 163.367
R753 B.n497 B.n496 163.367
R754 B.n493 B.n492 163.367
R755 B.n489 B.n488 163.367
R756 B.n485 B.n484 163.367
R757 B.n481 B.n480 163.367
R758 B.n477 B.n476 163.367
R759 B.n473 B.n472 163.367
R760 B.n468 B.n467 163.367
R761 B.n464 B.n463 163.367
R762 B.n460 B.n459 163.367
R763 B.n456 B.n455 163.367
R764 B.n452 B.n451 163.367
R765 B.n447 B.n446 163.367
R766 B.n443 B.n442 163.367
R767 B.n439 B.n438 163.367
R768 B.n435 B.n434 163.367
R769 B.n431 B.n430 163.367
R770 B.n427 B.n426 163.367
R771 B.n423 B.n422 163.367
R772 B.n419 B.n418 163.367
R773 B.n415 B.n414 163.367
R774 B.n411 B.n410 163.367
R775 B.n407 B.n406 163.367
R776 B.n403 B.n402 163.367
R777 B.n399 B.n398 163.367
R778 B.n395 B.n394 163.367
R779 B.n391 B.n390 163.367
R780 B.n387 B.n386 163.367
R781 B.n383 B.n382 163.367
R782 B.n543 B.n335 163.367
R783 B.n549 B.n331 163.367
R784 B.n549 B.n329 163.367
R785 B.n553 B.n329 163.367
R786 B.n553 B.n323 163.367
R787 B.n561 B.n323 163.367
R788 B.n561 B.n321 163.367
R789 B.n565 B.n321 163.367
R790 B.n565 B.n315 163.367
R791 B.n573 B.n315 163.367
R792 B.n573 B.n313 163.367
R793 B.n577 B.n313 163.367
R794 B.n577 B.n307 163.367
R795 B.n586 B.n307 163.367
R796 B.n586 B.n305 163.367
R797 B.n590 B.n305 163.367
R798 B.n590 B.n300 163.367
R799 B.n598 B.n300 163.367
R800 B.n598 B.n298 163.367
R801 B.n602 B.n298 163.367
R802 B.n602 B.n292 163.367
R803 B.n610 B.n292 163.367
R804 B.n610 B.n290 163.367
R805 B.n614 B.n290 163.367
R806 B.n614 B.n284 163.367
R807 B.n622 B.n284 163.367
R808 B.n622 B.n282 163.367
R809 B.n626 B.n282 163.367
R810 B.n626 B.n276 163.367
R811 B.n635 B.n276 163.367
R812 B.n635 B.n274 163.367
R813 B.n639 B.n274 163.367
R814 B.n639 B.n3 163.367
R815 B.n760 B.n3 163.367
R816 B.n756 B.n2 163.367
R817 B.n756 B.n755 163.367
R818 B.n755 B.n9 163.367
R819 B.n751 B.n9 163.367
R820 B.n751 B.n11 163.367
R821 B.n747 B.n11 163.367
R822 B.n747 B.n16 163.367
R823 B.n743 B.n16 163.367
R824 B.n743 B.n18 163.367
R825 B.n739 B.n18 163.367
R826 B.n739 B.n23 163.367
R827 B.n735 B.n23 163.367
R828 B.n735 B.n25 163.367
R829 B.n731 B.n25 163.367
R830 B.n731 B.n30 163.367
R831 B.n727 B.n30 163.367
R832 B.n727 B.n32 163.367
R833 B.n723 B.n32 163.367
R834 B.n723 B.n36 163.367
R835 B.n719 B.n36 163.367
R836 B.n719 B.n38 163.367
R837 B.n715 B.n38 163.367
R838 B.n715 B.n44 163.367
R839 B.n711 B.n44 163.367
R840 B.n711 B.n46 163.367
R841 B.n707 B.n46 163.367
R842 B.n707 B.n51 163.367
R843 B.n703 B.n51 163.367
R844 B.n703 B.n53 163.367
R845 B.n699 B.n53 163.367
R846 B.n699 B.n58 163.367
R847 B.n695 B.n58 163.367
R848 B.n695 B.n60 163.367
R849 B.n104 B.t10 102.397
R850 B.n379 B.t18 102.397
R851 B.n107 B.t20 102.383
R852 B.n377 B.t15 102.383
R853 B.n542 B.n332 82.899
R854 B.n693 B.n692 82.899
R855 B.n110 B.n63 71.676
R856 B.n114 B.n64 71.676
R857 B.n118 B.n65 71.676
R858 B.n122 B.n66 71.676
R859 B.n126 B.n67 71.676
R860 B.n130 B.n68 71.676
R861 B.n134 B.n69 71.676
R862 B.n138 B.n70 71.676
R863 B.n142 B.n71 71.676
R864 B.n146 B.n72 71.676
R865 B.n150 B.n73 71.676
R866 B.n154 B.n74 71.676
R867 B.n158 B.n75 71.676
R868 B.n162 B.n76 71.676
R869 B.n166 B.n77 71.676
R870 B.n170 B.n78 71.676
R871 B.n174 B.n79 71.676
R872 B.n178 B.n80 71.676
R873 B.n182 B.n81 71.676
R874 B.n186 B.n82 71.676
R875 B.n190 B.n83 71.676
R876 B.n194 B.n84 71.676
R877 B.n198 B.n85 71.676
R878 B.n202 B.n86 71.676
R879 B.n206 B.n87 71.676
R880 B.n210 B.n88 71.676
R881 B.n214 B.n89 71.676
R882 B.n218 B.n90 71.676
R883 B.n222 B.n91 71.676
R884 B.n226 B.n92 71.676
R885 B.n230 B.n93 71.676
R886 B.n234 B.n94 71.676
R887 B.n238 B.n95 71.676
R888 B.n242 B.n96 71.676
R889 B.n246 B.n97 71.676
R890 B.n250 B.n98 71.676
R891 B.n254 B.n99 71.676
R892 B.n258 B.n100 71.676
R893 B.n262 B.n101 71.676
R894 B.n266 B.n102 71.676
R895 B.n691 B.n103 71.676
R896 B.n691 B.n690 71.676
R897 B.n268 B.n102 71.676
R898 B.n265 B.n101 71.676
R899 B.n261 B.n100 71.676
R900 B.n257 B.n99 71.676
R901 B.n253 B.n98 71.676
R902 B.n249 B.n97 71.676
R903 B.n245 B.n96 71.676
R904 B.n241 B.n95 71.676
R905 B.n237 B.n94 71.676
R906 B.n233 B.n93 71.676
R907 B.n229 B.n92 71.676
R908 B.n225 B.n91 71.676
R909 B.n221 B.n90 71.676
R910 B.n217 B.n89 71.676
R911 B.n213 B.n88 71.676
R912 B.n209 B.n87 71.676
R913 B.n205 B.n86 71.676
R914 B.n201 B.n85 71.676
R915 B.n197 B.n84 71.676
R916 B.n193 B.n83 71.676
R917 B.n189 B.n82 71.676
R918 B.n185 B.n81 71.676
R919 B.n181 B.n80 71.676
R920 B.n177 B.n79 71.676
R921 B.n173 B.n78 71.676
R922 B.n169 B.n77 71.676
R923 B.n165 B.n76 71.676
R924 B.n161 B.n75 71.676
R925 B.n157 B.n74 71.676
R926 B.n153 B.n73 71.676
R927 B.n149 B.n72 71.676
R928 B.n145 B.n71 71.676
R929 B.n141 B.n70 71.676
R930 B.n137 B.n69 71.676
R931 B.n133 B.n68 71.676
R932 B.n129 B.n67 71.676
R933 B.n125 B.n66 71.676
R934 B.n121 B.n65 71.676
R935 B.n117 B.n64 71.676
R936 B.n113 B.n63 71.676
R937 B.n541 B.n540 71.676
R938 B.n535 B.n336 71.676
R939 B.n532 B.n337 71.676
R940 B.n528 B.n338 71.676
R941 B.n524 B.n339 71.676
R942 B.n520 B.n340 71.676
R943 B.n516 B.n341 71.676
R944 B.n512 B.n342 71.676
R945 B.n508 B.n343 71.676
R946 B.n504 B.n344 71.676
R947 B.n500 B.n345 71.676
R948 B.n496 B.n346 71.676
R949 B.n492 B.n347 71.676
R950 B.n488 B.n348 71.676
R951 B.n484 B.n349 71.676
R952 B.n480 B.n350 71.676
R953 B.n476 B.n351 71.676
R954 B.n472 B.n352 71.676
R955 B.n467 B.n353 71.676
R956 B.n463 B.n354 71.676
R957 B.n459 B.n355 71.676
R958 B.n455 B.n356 71.676
R959 B.n451 B.n357 71.676
R960 B.n446 B.n358 71.676
R961 B.n442 B.n359 71.676
R962 B.n438 B.n360 71.676
R963 B.n434 B.n361 71.676
R964 B.n430 B.n362 71.676
R965 B.n426 B.n363 71.676
R966 B.n422 B.n364 71.676
R967 B.n418 B.n365 71.676
R968 B.n414 B.n366 71.676
R969 B.n410 B.n367 71.676
R970 B.n406 B.n368 71.676
R971 B.n402 B.n369 71.676
R972 B.n398 B.n370 71.676
R973 B.n394 B.n371 71.676
R974 B.n390 B.n372 71.676
R975 B.n386 B.n373 71.676
R976 B.n382 B.n374 71.676
R977 B.n541 B.n376 71.676
R978 B.n533 B.n336 71.676
R979 B.n529 B.n337 71.676
R980 B.n525 B.n338 71.676
R981 B.n521 B.n339 71.676
R982 B.n517 B.n340 71.676
R983 B.n513 B.n341 71.676
R984 B.n509 B.n342 71.676
R985 B.n505 B.n343 71.676
R986 B.n501 B.n344 71.676
R987 B.n497 B.n345 71.676
R988 B.n493 B.n346 71.676
R989 B.n489 B.n347 71.676
R990 B.n485 B.n348 71.676
R991 B.n481 B.n349 71.676
R992 B.n477 B.n350 71.676
R993 B.n473 B.n351 71.676
R994 B.n468 B.n352 71.676
R995 B.n464 B.n353 71.676
R996 B.n460 B.n354 71.676
R997 B.n456 B.n355 71.676
R998 B.n452 B.n356 71.676
R999 B.n447 B.n357 71.676
R1000 B.n443 B.n358 71.676
R1001 B.n439 B.n359 71.676
R1002 B.n435 B.n360 71.676
R1003 B.n431 B.n361 71.676
R1004 B.n427 B.n362 71.676
R1005 B.n423 B.n363 71.676
R1006 B.n419 B.n364 71.676
R1007 B.n415 B.n365 71.676
R1008 B.n411 B.n366 71.676
R1009 B.n407 B.n367 71.676
R1010 B.n403 B.n368 71.676
R1011 B.n399 B.n369 71.676
R1012 B.n395 B.n370 71.676
R1013 B.n391 B.n371 71.676
R1014 B.n387 B.n372 71.676
R1015 B.n383 B.n373 71.676
R1016 B.n374 B.n335 71.676
R1017 B.n761 B.n760 71.676
R1018 B.n761 B.n2 71.676
R1019 B.n105 B.t11 69.0388
R1020 B.n380 B.t17 69.0388
R1021 B.n108 B.t21 69.0261
R1022 B.n378 B.t14 69.0261
R1023 B.n109 B.n108 59.5399
R1024 B.n106 B.n105 59.5399
R1025 B.n449 B.n380 59.5399
R1026 B.n470 B.n378 59.5399
R1027 B.n548 B.n332 48.1809
R1028 B.n548 B.n328 48.1809
R1029 B.n554 B.n328 48.1809
R1030 B.n554 B.n324 48.1809
R1031 B.n560 B.n324 48.1809
R1032 B.n566 B.n320 48.1809
R1033 B.n566 B.n316 48.1809
R1034 B.n572 B.n316 48.1809
R1035 B.n572 B.n312 48.1809
R1036 B.n578 B.n312 48.1809
R1037 B.n578 B.n308 48.1809
R1038 B.n585 B.n308 48.1809
R1039 B.n585 B.n584 48.1809
R1040 B.n591 B.n301 48.1809
R1041 B.n597 B.n301 48.1809
R1042 B.n597 B.n297 48.1809
R1043 B.n603 B.n297 48.1809
R1044 B.n609 B.n293 48.1809
R1045 B.n609 B.n288 48.1809
R1046 B.n615 B.n288 48.1809
R1047 B.n615 B.n289 48.1809
R1048 B.n621 B.n281 48.1809
R1049 B.n627 B.n281 48.1809
R1050 B.n627 B.n277 48.1809
R1051 B.n634 B.n277 48.1809
R1052 B.n640 B.n273 48.1809
R1053 B.n640 B.n4 48.1809
R1054 B.n759 B.n4 48.1809
R1055 B.n759 B.n758 48.1809
R1056 B.n758 B.n757 48.1809
R1057 B.n757 B.n8 48.1809
R1058 B.n649 B.n8 48.1809
R1059 B.n750 B.n749 48.1809
R1060 B.n749 B.n748 48.1809
R1061 B.n748 B.n15 48.1809
R1062 B.n742 B.n15 48.1809
R1063 B.n741 B.n740 48.1809
R1064 B.n740 B.n22 48.1809
R1065 B.n734 B.n22 48.1809
R1066 B.n734 B.n733 48.1809
R1067 B.n732 B.n29 48.1809
R1068 B.n726 B.n29 48.1809
R1069 B.n726 B.n725 48.1809
R1070 B.n725 B.n724 48.1809
R1071 B.n718 B.n39 48.1809
R1072 B.n718 B.n717 48.1809
R1073 B.n717 B.n716 48.1809
R1074 B.n716 B.n43 48.1809
R1075 B.n710 B.n43 48.1809
R1076 B.n710 B.n709 48.1809
R1077 B.n709 B.n708 48.1809
R1078 B.n708 B.n50 48.1809
R1079 B.n702 B.n701 48.1809
R1080 B.n701 B.n700 48.1809
R1081 B.n700 B.n57 48.1809
R1082 B.n694 B.n57 48.1809
R1083 B.n694 B.n693 48.1809
R1084 B.n560 B.t13 44.6382
R1085 B.n702 B.t9 44.6382
R1086 B.n591 B.t2 38.9699
R1087 B.n724 B.t1 38.9699
R1088 B.t7 B.n293 36.1358
R1089 B.n733 B.t0 36.1358
R1090 B.n539 B.n330 34.1859
R1091 B.n545 B.n544 34.1859
R1092 B.n689 B.n688 34.1859
R1093 B.n111 B.n59 34.1859
R1094 B.n108 B.n107 33.3581
R1095 B.n105 B.n104 33.3581
R1096 B.n380 B.n379 33.3581
R1097 B.n378 B.n377 33.3581
R1098 B.n621 B.t3 33.3016
R1099 B.n742 B.t6 33.3016
R1100 B.t5 B.n273 30.4675
R1101 B.n649 B.t4 30.4675
R1102 B B.n762 18.0485
R1103 B.n634 B.t5 17.7139
R1104 B.n750 B.t4 17.7139
R1105 B.n289 B.t3 14.8797
R1106 B.t6 B.n741 14.8797
R1107 B.n603 B.t7 12.0456
R1108 B.t0 B.n732 12.0456
R1109 B.n550 B.n330 10.6151
R1110 B.n551 B.n550 10.6151
R1111 B.n552 B.n551 10.6151
R1112 B.n552 B.n322 10.6151
R1113 B.n562 B.n322 10.6151
R1114 B.n563 B.n562 10.6151
R1115 B.n564 B.n563 10.6151
R1116 B.n564 B.n314 10.6151
R1117 B.n574 B.n314 10.6151
R1118 B.n575 B.n574 10.6151
R1119 B.n576 B.n575 10.6151
R1120 B.n576 B.n306 10.6151
R1121 B.n587 B.n306 10.6151
R1122 B.n588 B.n587 10.6151
R1123 B.n589 B.n588 10.6151
R1124 B.n589 B.n299 10.6151
R1125 B.n599 B.n299 10.6151
R1126 B.n600 B.n599 10.6151
R1127 B.n601 B.n600 10.6151
R1128 B.n601 B.n291 10.6151
R1129 B.n611 B.n291 10.6151
R1130 B.n612 B.n611 10.6151
R1131 B.n613 B.n612 10.6151
R1132 B.n613 B.n283 10.6151
R1133 B.n623 B.n283 10.6151
R1134 B.n624 B.n623 10.6151
R1135 B.n625 B.n624 10.6151
R1136 B.n625 B.n275 10.6151
R1137 B.n636 B.n275 10.6151
R1138 B.n637 B.n636 10.6151
R1139 B.n638 B.n637 10.6151
R1140 B.n638 B.n0 10.6151
R1141 B.n539 B.n538 10.6151
R1142 B.n538 B.n537 10.6151
R1143 B.n537 B.n536 10.6151
R1144 B.n536 B.n534 10.6151
R1145 B.n534 B.n531 10.6151
R1146 B.n531 B.n530 10.6151
R1147 B.n530 B.n527 10.6151
R1148 B.n527 B.n526 10.6151
R1149 B.n526 B.n523 10.6151
R1150 B.n523 B.n522 10.6151
R1151 B.n522 B.n519 10.6151
R1152 B.n519 B.n518 10.6151
R1153 B.n518 B.n515 10.6151
R1154 B.n515 B.n514 10.6151
R1155 B.n514 B.n511 10.6151
R1156 B.n511 B.n510 10.6151
R1157 B.n510 B.n507 10.6151
R1158 B.n507 B.n506 10.6151
R1159 B.n506 B.n503 10.6151
R1160 B.n503 B.n502 10.6151
R1161 B.n502 B.n499 10.6151
R1162 B.n499 B.n498 10.6151
R1163 B.n498 B.n495 10.6151
R1164 B.n495 B.n494 10.6151
R1165 B.n494 B.n491 10.6151
R1166 B.n491 B.n490 10.6151
R1167 B.n490 B.n487 10.6151
R1168 B.n487 B.n486 10.6151
R1169 B.n486 B.n483 10.6151
R1170 B.n483 B.n482 10.6151
R1171 B.n482 B.n479 10.6151
R1172 B.n479 B.n478 10.6151
R1173 B.n478 B.n475 10.6151
R1174 B.n475 B.n474 10.6151
R1175 B.n474 B.n471 10.6151
R1176 B.n469 B.n466 10.6151
R1177 B.n466 B.n465 10.6151
R1178 B.n465 B.n462 10.6151
R1179 B.n462 B.n461 10.6151
R1180 B.n461 B.n458 10.6151
R1181 B.n458 B.n457 10.6151
R1182 B.n457 B.n454 10.6151
R1183 B.n454 B.n453 10.6151
R1184 B.n453 B.n450 10.6151
R1185 B.n448 B.n445 10.6151
R1186 B.n445 B.n444 10.6151
R1187 B.n444 B.n441 10.6151
R1188 B.n441 B.n440 10.6151
R1189 B.n440 B.n437 10.6151
R1190 B.n437 B.n436 10.6151
R1191 B.n436 B.n433 10.6151
R1192 B.n433 B.n432 10.6151
R1193 B.n432 B.n429 10.6151
R1194 B.n429 B.n428 10.6151
R1195 B.n428 B.n425 10.6151
R1196 B.n425 B.n424 10.6151
R1197 B.n424 B.n421 10.6151
R1198 B.n421 B.n420 10.6151
R1199 B.n420 B.n417 10.6151
R1200 B.n417 B.n416 10.6151
R1201 B.n416 B.n413 10.6151
R1202 B.n413 B.n412 10.6151
R1203 B.n412 B.n409 10.6151
R1204 B.n409 B.n408 10.6151
R1205 B.n408 B.n405 10.6151
R1206 B.n405 B.n404 10.6151
R1207 B.n404 B.n401 10.6151
R1208 B.n401 B.n400 10.6151
R1209 B.n400 B.n397 10.6151
R1210 B.n397 B.n396 10.6151
R1211 B.n396 B.n393 10.6151
R1212 B.n393 B.n392 10.6151
R1213 B.n392 B.n389 10.6151
R1214 B.n389 B.n388 10.6151
R1215 B.n388 B.n385 10.6151
R1216 B.n385 B.n384 10.6151
R1217 B.n384 B.n381 10.6151
R1218 B.n381 B.n334 10.6151
R1219 B.n544 B.n334 10.6151
R1220 B.n546 B.n545 10.6151
R1221 B.n546 B.n326 10.6151
R1222 B.n556 B.n326 10.6151
R1223 B.n557 B.n556 10.6151
R1224 B.n558 B.n557 10.6151
R1225 B.n558 B.n318 10.6151
R1226 B.n568 B.n318 10.6151
R1227 B.n569 B.n568 10.6151
R1228 B.n570 B.n569 10.6151
R1229 B.n570 B.n310 10.6151
R1230 B.n580 B.n310 10.6151
R1231 B.n581 B.n580 10.6151
R1232 B.n582 B.n581 10.6151
R1233 B.n582 B.n303 10.6151
R1234 B.n593 B.n303 10.6151
R1235 B.n594 B.n593 10.6151
R1236 B.n595 B.n594 10.6151
R1237 B.n595 B.n295 10.6151
R1238 B.n605 B.n295 10.6151
R1239 B.n606 B.n605 10.6151
R1240 B.n607 B.n606 10.6151
R1241 B.n607 B.n286 10.6151
R1242 B.n617 B.n286 10.6151
R1243 B.n618 B.n617 10.6151
R1244 B.n619 B.n618 10.6151
R1245 B.n619 B.n279 10.6151
R1246 B.n629 B.n279 10.6151
R1247 B.n630 B.n629 10.6151
R1248 B.n632 B.n630 10.6151
R1249 B.n632 B.n631 10.6151
R1250 B.n631 B.n271 10.6151
R1251 B.n643 B.n271 10.6151
R1252 B.n644 B.n643 10.6151
R1253 B.n645 B.n644 10.6151
R1254 B.n646 B.n645 10.6151
R1255 B.n647 B.n646 10.6151
R1256 B.n651 B.n647 10.6151
R1257 B.n652 B.n651 10.6151
R1258 B.n653 B.n652 10.6151
R1259 B.n654 B.n653 10.6151
R1260 B.n656 B.n654 10.6151
R1261 B.n657 B.n656 10.6151
R1262 B.n658 B.n657 10.6151
R1263 B.n659 B.n658 10.6151
R1264 B.n661 B.n659 10.6151
R1265 B.n662 B.n661 10.6151
R1266 B.n663 B.n662 10.6151
R1267 B.n664 B.n663 10.6151
R1268 B.n666 B.n664 10.6151
R1269 B.n667 B.n666 10.6151
R1270 B.n668 B.n667 10.6151
R1271 B.n669 B.n668 10.6151
R1272 B.n671 B.n669 10.6151
R1273 B.n672 B.n671 10.6151
R1274 B.n673 B.n672 10.6151
R1275 B.n674 B.n673 10.6151
R1276 B.n676 B.n674 10.6151
R1277 B.n677 B.n676 10.6151
R1278 B.n678 B.n677 10.6151
R1279 B.n679 B.n678 10.6151
R1280 B.n681 B.n679 10.6151
R1281 B.n682 B.n681 10.6151
R1282 B.n683 B.n682 10.6151
R1283 B.n684 B.n683 10.6151
R1284 B.n686 B.n684 10.6151
R1285 B.n687 B.n686 10.6151
R1286 B.n688 B.n687 10.6151
R1287 B.n754 B.n1 10.6151
R1288 B.n754 B.n753 10.6151
R1289 B.n753 B.n752 10.6151
R1290 B.n752 B.n10 10.6151
R1291 B.n746 B.n10 10.6151
R1292 B.n746 B.n745 10.6151
R1293 B.n745 B.n744 10.6151
R1294 B.n744 B.n17 10.6151
R1295 B.n738 B.n17 10.6151
R1296 B.n738 B.n737 10.6151
R1297 B.n737 B.n736 10.6151
R1298 B.n736 B.n24 10.6151
R1299 B.n730 B.n24 10.6151
R1300 B.n730 B.n729 10.6151
R1301 B.n729 B.n728 10.6151
R1302 B.n728 B.n31 10.6151
R1303 B.n722 B.n31 10.6151
R1304 B.n722 B.n721 10.6151
R1305 B.n721 B.n720 10.6151
R1306 B.n720 B.n37 10.6151
R1307 B.n714 B.n37 10.6151
R1308 B.n714 B.n713 10.6151
R1309 B.n713 B.n712 10.6151
R1310 B.n712 B.n45 10.6151
R1311 B.n706 B.n45 10.6151
R1312 B.n706 B.n705 10.6151
R1313 B.n705 B.n704 10.6151
R1314 B.n704 B.n52 10.6151
R1315 B.n698 B.n52 10.6151
R1316 B.n698 B.n697 10.6151
R1317 B.n697 B.n696 10.6151
R1318 B.n696 B.n59 10.6151
R1319 B.n112 B.n111 10.6151
R1320 B.n115 B.n112 10.6151
R1321 B.n116 B.n115 10.6151
R1322 B.n119 B.n116 10.6151
R1323 B.n120 B.n119 10.6151
R1324 B.n123 B.n120 10.6151
R1325 B.n124 B.n123 10.6151
R1326 B.n127 B.n124 10.6151
R1327 B.n128 B.n127 10.6151
R1328 B.n131 B.n128 10.6151
R1329 B.n132 B.n131 10.6151
R1330 B.n135 B.n132 10.6151
R1331 B.n136 B.n135 10.6151
R1332 B.n139 B.n136 10.6151
R1333 B.n140 B.n139 10.6151
R1334 B.n143 B.n140 10.6151
R1335 B.n144 B.n143 10.6151
R1336 B.n147 B.n144 10.6151
R1337 B.n148 B.n147 10.6151
R1338 B.n151 B.n148 10.6151
R1339 B.n152 B.n151 10.6151
R1340 B.n155 B.n152 10.6151
R1341 B.n156 B.n155 10.6151
R1342 B.n159 B.n156 10.6151
R1343 B.n160 B.n159 10.6151
R1344 B.n163 B.n160 10.6151
R1345 B.n164 B.n163 10.6151
R1346 B.n167 B.n164 10.6151
R1347 B.n168 B.n167 10.6151
R1348 B.n171 B.n168 10.6151
R1349 B.n172 B.n171 10.6151
R1350 B.n175 B.n172 10.6151
R1351 B.n176 B.n175 10.6151
R1352 B.n179 B.n176 10.6151
R1353 B.n180 B.n179 10.6151
R1354 B.n184 B.n183 10.6151
R1355 B.n187 B.n184 10.6151
R1356 B.n188 B.n187 10.6151
R1357 B.n191 B.n188 10.6151
R1358 B.n192 B.n191 10.6151
R1359 B.n195 B.n192 10.6151
R1360 B.n196 B.n195 10.6151
R1361 B.n199 B.n196 10.6151
R1362 B.n200 B.n199 10.6151
R1363 B.n204 B.n203 10.6151
R1364 B.n207 B.n204 10.6151
R1365 B.n208 B.n207 10.6151
R1366 B.n211 B.n208 10.6151
R1367 B.n212 B.n211 10.6151
R1368 B.n215 B.n212 10.6151
R1369 B.n216 B.n215 10.6151
R1370 B.n219 B.n216 10.6151
R1371 B.n220 B.n219 10.6151
R1372 B.n223 B.n220 10.6151
R1373 B.n224 B.n223 10.6151
R1374 B.n227 B.n224 10.6151
R1375 B.n228 B.n227 10.6151
R1376 B.n231 B.n228 10.6151
R1377 B.n232 B.n231 10.6151
R1378 B.n235 B.n232 10.6151
R1379 B.n236 B.n235 10.6151
R1380 B.n239 B.n236 10.6151
R1381 B.n240 B.n239 10.6151
R1382 B.n243 B.n240 10.6151
R1383 B.n244 B.n243 10.6151
R1384 B.n247 B.n244 10.6151
R1385 B.n248 B.n247 10.6151
R1386 B.n251 B.n248 10.6151
R1387 B.n252 B.n251 10.6151
R1388 B.n255 B.n252 10.6151
R1389 B.n256 B.n255 10.6151
R1390 B.n259 B.n256 10.6151
R1391 B.n260 B.n259 10.6151
R1392 B.n263 B.n260 10.6151
R1393 B.n264 B.n263 10.6151
R1394 B.n267 B.n264 10.6151
R1395 B.n269 B.n267 10.6151
R1396 B.n270 B.n269 10.6151
R1397 B.n689 B.n270 10.6151
R1398 B.n471 B.n470 9.36635
R1399 B.n449 B.n448 9.36635
R1400 B.n180 B.n109 9.36635
R1401 B.n203 B.n106 9.36635
R1402 B.n584 B.t2 9.21145
R1403 B.n39 B.t1 9.21145
R1404 B.n762 B.n0 8.11757
R1405 B.n762 B.n1 8.11757
R1406 B.t13 B.n320 3.54317
R1407 B.t9 B.n50 3.54317
R1408 B.n470 B.n469 1.24928
R1409 B.n450 B.n449 1.24928
R1410 B.n183 B.n109 1.24928
R1411 B.n200 B.n106 1.24928
R1412 VP.n11 VP.t5 209.338
R1413 VP.n5 VP.t7 177.716
R1414 VP.n29 VP.t2 177.716
R1415 VP.n36 VP.t6 177.716
R1416 VP.n43 VP.t1 177.716
R1417 VP.n23 VP.t0 177.716
R1418 VP.n16 VP.t3 177.716
R1419 VP.n10 VP.t4 177.716
R1420 VP.n25 VP.n5 169.619
R1421 VP.n44 VP.n43 169.619
R1422 VP.n24 VP.n23 169.619
R1423 VP.n12 VP.n9 161.3
R1424 VP.n14 VP.n13 161.3
R1425 VP.n15 VP.n8 161.3
R1426 VP.n18 VP.n17 161.3
R1427 VP.n19 VP.n7 161.3
R1428 VP.n21 VP.n20 161.3
R1429 VP.n22 VP.n6 161.3
R1430 VP.n42 VP.n0 161.3
R1431 VP.n41 VP.n40 161.3
R1432 VP.n39 VP.n1 161.3
R1433 VP.n38 VP.n37 161.3
R1434 VP.n35 VP.n2 161.3
R1435 VP.n34 VP.n33 161.3
R1436 VP.n32 VP.n3 161.3
R1437 VP.n31 VP.n30 161.3
R1438 VP.n28 VP.n4 161.3
R1439 VP.n27 VP.n26 161.3
R1440 VP.n11 VP.n10 59.48
R1441 VP.n35 VP.n34 56.5193
R1442 VP.n15 VP.n14 56.5193
R1443 VP.n25 VP.n24 43.902
R1444 VP.n30 VP.n28 43.4072
R1445 VP.n41 VP.n1 43.4072
R1446 VP.n21 VP.n7 43.4072
R1447 VP.n28 VP.n27 37.5796
R1448 VP.n42 VP.n41 37.5796
R1449 VP.n22 VP.n21 37.5796
R1450 VP.n12 VP.n11 26.5029
R1451 VP.n34 VP.n3 24.4675
R1452 VP.n37 VP.n35 24.4675
R1453 VP.n17 VP.n15 24.4675
R1454 VP.n14 VP.n9 24.4675
R1455 VP.n30 VP.n29 19.0848
R1456 VP.n36 VP.n1 19.0848
R1457 VP.n16 VP.n7 19.0848
R1458 VP.n27 VP.n5 16.1487
R1459 VP.n43 VP.n42 16.1487
R1460 VP.n23 VP.n22 16.1487
R1461 VP.n29 VP.n3 5.38324
R1462 VP.n37 VP.n36 5.38324
R1463 VP.n17 VP.n16 5.38324
R1464 VP.n10 VP.n9 5.38324
R1465 VP.n13 VP.n12 0.189894
R1466 VP.n13 VP.n8 0.189894
R1467 VP.n18 VP.n8 0.189894
R1468 VP.n19 VP.n18 0.189894
R1469 VP.n20 VP.n19 0.189894
R1470 VP.n20 VP.n6 0.189894
R1471 VP.n24 VP.n6 0.189894
R1472 VP.n26 VP.n25 0.189894
R1473 VP.n26 VP.n4 0.189894
R1474 VP.n31 VP.n4 0.189894
R1475 VP.n32 VP.n31 0.189894
R1476 VP.n33 VP.n32 0.189894
R1477 VP.n33 VP.n2 0.189894
R1478 VP.n38 VP.n2 0.189894
R1479 VP.n39 VP.n38 0.189894
R1480 VP.n40 VP.n39 0.189894
R1481 VP.n40 VP.n0 0.189894
R1482 VP.n44 VP.n0 0.189894
R1483 VP VP.n44 0.0516364
R1484 VDD1 VDD1.n0 61.925
R1485 VDD1.n3 VDD1.n2 61.8112
R1486 VDD1.n3 VDD1.n1 61.8112
R1487 VDD1.n5 VDD1.n4 61.1252
R1488 VDD1.n5 VDD1.n3 39.8069
R1489 VDD1.n4 VDD1.t4 1.93221
R1490 VDD1.n4 VDD1.t7 1.93221
R1491 VDD1.n0 VDD1.t2 1.93221
R1492 VDD1.n0 VDD1.t3 1.93221
R1493 VDD1.n2 VDD1.t1 1.93221
R1494 VDD1.n2 VDD1.t6 1.93221
R1495 VDD1.n1 VDD1.t0 1.93221
R1496 VDD1.n1 VDD1.t5 1.93221
R1497 VDD1 VDD1.n5 0.68369
C0 VN VDD1 0.14911f
C1 VDD2 VP 0.390484f
C2 VDD2 VTAIL 7.82344f
C3 VTAIL VP 6.44965f
C4 VDD2 VN 6.36995f
C5 VN VP 5.85598f
C6 VDD2 VDD1 1.16999f
C7 VDD1 VP 6.61054f
C8 VN VTAIL 6.43555f
C9 VTAIL VDD1 7.77713f
C10 VDD2 B 4.014982f
C11 VDD1 B 4.322824f
C12 VTAIL B 8.5462f
C13 VN B 10.80582f
C14 VP B 9.21159f
C15 VDD1.t2 B 0.204907f
C16 VDD1.t3 B 0.204907f
C17 VDD1.n0 B 1.81117f
C18 VDD1.t0 B 0.204907f
C19 VDD1.t5 B 0.204907f
C20 VDD1.n1 B 1.81034f
C21 VDD1.t1 B 0.204907f
C22 VDD1.t6 B 0.204907f
C23 VDD1.n2 B 1.81034f
C24 VDD1.n3 B 2.54979f
C25 VDD1.t4 B 0.204907f
C26 VDD1.t7 B 0.204907f
C27 VDD1.n4 B 1.80595f
C28 VDD1.n5 B 2.45313f
C29 VP.n0 B 0.033058f
C30 VP.t1 B 1.27702f
C31 VP.n1 B 0.057837f
C32 VP.n2 B 0.033058f
C33 VP.n3 B 0.037886f
C34 VP.n4 B 0.033058f
C35 VP.t7 B 1.27702f
C36 VP.n5 B 0.541716f
C37 VP.n6 B 0.033058f
C38 VP.t0 B 1.27702f
C39 VP.n7 B 0.057837f
C40 VP.n8 B 0.033058f
C41 VP.n9 B 0.037886f
C42 VP.t5 B 1.36544f
C43 VP.t4 B 1.27702f
C44 VP.n10 B 0.518834f
C45 VP.n11 B 0.547728f
C46 VP.n12 B 0.178404f
C47 VP.n13 B 0.033058f
C48 VP.n14 B 0.048259f
C49 VP.n15 B 0.048259f
C50 VP.t3 B 1.27702f
C51 VP.n16 B 0.470399f
C52 VP.n17 B 0.037886f
C53 VP.n18 B 0.033058f
C54 VP.n19 B 0.033058f
C55 VP.n20 B 0.033058f
C56 VP.n21 B 0.027108f
C57 VP.n22 B 0.056149f
C58 VP.n23 B 0.541716f
C59 VP.n24 B 1.47116f
C60 VP.n25 B 1.49823f
C61 VP.n26 B 0.033058f
C62 VP.n27 B 0.056149f
C63 VP.n28 B 0.027108f
C64 VP.t2 B 1.27702f
C65 VP.n29 B 0.470399f
C66 VP.n30 B 0.057837f
C67 VP.n31 B 0.033058f
C68 VP.n32 B 0.033058f
C69 VP.n33 B 0.033058f
C70 VP.n34 B 0.048259f
C71 VP.n35 B 0.048259f
C72 VP.t6 B 1.27702f
C73 VP.n36 B 0.470399f
C74 VP.n37 B 0.037886f
C75 VP.n38 B 0.033058f
C76 VP.n39 B 0.033058f
C77 VP.n40 B 0.033058f
C78 VP.n41 B 0.027108f
C79 VP.n42 B 0.056149f
C80 VP.n43 B 0.541716f
C81 VP.n44 B 0.029297f
C82 VDD2.t2 B 0.203381f
C83 VDD2.t0 B 0.203381f
C84 VDD2.n0 B 1.79686f
C85 VDD2.t1 B 0.203381f
C86 VDD2.t7 B 0.203381f
C87 VDD2.n1 B 1.79686f
C88 VDD2.n2 B 2.47765f
C89 VDD2.t6 B 0.203381f
C90 VDD2.t4 B 0.203381f
C91 VDD2.n3 B 1.7925f
C92 VDD2.n4 B 2.40467f
C93 VDD2.t5 B 0.203381f
C94 VDD2.t3 B 0.203381f
C95 VDD2.n5 B 1.79683f
C96 VTAIL.t8 B 0.158597f
C97 VTAIL.t9 B 0.158597f
C98 VTAIL.n0 B 1.33875f
C99 VTAIL.n1 B 0.290764f
C100 VTAIL.t13 B 1.70411f
C101 VTAIL.n2 B 0.383906f
C102 VTAIL.t5 B 1.70411f
C103 VTAIL.n3 B 0.383906f
C104 VTAIL.t7 B 0.158597f
C105 VTAIL.t3 B 0.158597f
C106 VTAIL.n4 B 1.33875f
C107 VTAIL.n5 B 0.380643f
C108 VTAIL.t2 B 1.70411f
C109 VTAIL.n6 B 1.27128f
C110 VTAIL.t15 B 1.70412f
C111 VTAIL.n7 B 1.27128f
C112 VTAIL.t11 B 0.158597f
C113 VTAIL.t14 B 0.158597f
C114 VTAIL.n8 B 1.33875f
C115 VTAIL.n9 B 0.380639f
C116 VTAIL.t12 B 1.70412f
C117 VTAIL.n10 B 0.383902f
C118 VTAIL.t4 B 1.70412f
C119 VTAIL.n11 B 0.383902f
C120 VTAIL.t6 B 0.158597f
C121 VTAIL.t0 B 0.158597f
C122 VTAIL.n12 B 1.33875f
C123 VTAIL.n13 B 0.380639f
C124 VTAIL.t1 B 1.70411f
C125 VTAIL.n14 B 1.27128f
C126 VTAIL.t10 B 1.70411f
C127 VTAIL.n15 B 1.26761f
C128 VN.n0 B 0.032628f
C129 VN.t0 B 1.26041f
C130 VN.n1 B 0.057085f
C131 VN.n2 B 0.032628f
C132 VN.n3 B 0.037393f
C133 VN.t5 B 1.34768f
C134 VN.t7 B 1.26041f
C135 VN.n4 B 0.512085f
C136 VN.n5 B 0.540603f
C137 VN.n6 B 0.176083f
C138 VN.n7 B 0.032628f
C139 VN.n8 B 0.047631f
C140 VN.n9 B 0.047631f
C141 VN.t6 B 1.26041f
C142 VN.n10 B 0.46428f
C143 VN.n11 B 0.037393f
C144 VN.n12 B 0.032628f
C145 VN.n13 B 0.032628f
C146 VN.n14 B 0.032628f
C147 VN.n15 B 0.026756f
C148 VN.n16 B 0.055419f
C149 VN.n17 B 0.534669f
C150 VN.n18 B 0.028916f
C151 VN.n19 B 0.032628f
C152 VN.t1 B 1.26041f
C153 VN.n20 B 0.057085f
C154 VN.n21 B 0.032628f
C155 VN.t3 B 1.26041f
C156 VN.n22 B 0.46428f
C157 VN.n23 B 0.037393f
C158 VN.t4 B 1.34768f
C159 VN.t2 B 1.26041f
C160 VN.n24 B 0.512085f
C161 VN.n25 B 0.540603f
C162 VN.n26 B 0.176083f
C163 VN.n27 B 0.032628f
C164 VN.n28 B 0.047631f
C165 VN.n29 B 0.047631f
C166 VN.n30 B 0.037393f
C167 VN.n31 B 0.032628f
C168 VN.n32 B 0.032628f
C169 VN.n33 B 0.032628f
C170 VN.n34 B 0.026756f
C171 VN.n35 B 0.055419f
C172 VN.n36 B 0.534669f
C173 VN.n37 B 1.47339f
.ends

