* NGSPICE file created from diff_pair_sample_0446.ext - technology: sky130A

.subckt diff_pair_sample_0446 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=2.1957 ps=12.04 w=5.63 l=1.07
X1 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=0 ps=0 w=5.63 l=1.07
X2 VDD2.t0 VN.t1 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=2.1957 ps=12.04 w=5.63 l=1.07
X3 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=0 ps=0 w=5.63 l=1.07
X4 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=2.1957 ps=12.04 w=5.63 l=1.07
X5 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=2.1957 ps=12.04 w=5.63 l=1.07
X6 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=0 ps=0 w=5.63 l=1.07
X7 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1957 pd=12.04 as=0 ps=0 w=5.63 l=1.07
R0 VN VN.t0 361.214
R1 VN VN.t1 325.096
R2 VTAIL.n1 VTAIL.t2 54.5142
R3 VTAIL.n3 VTAIL.t3 54.514
R4 VTAIL.n0 VTAIL.t0 54.514
R5 VTAIL.n2 VTAIL.t1 54.514
R6 VTAIL.n1 VTAIL.n0 19.6514
R7 VTAIL.n3 VTAIL.n2 18.4445
R8 VTAIL.n2 VTAIL.n1 1.07378
R9 VTAIL VTAIL.n0 0.830241
R10 VTAIL VTAIL.n3 0.244034
R11 VDD2.n0 VDD2.t0 102.136
R12 VDD2.n0 VDD2.t1 71.1927
R13 VDD2 VDD2.n0 0.360414
R14 B.n419 B.n418 585
R15 B.n420 B.n419 585
R16 B.n172 B.n61 585
R17 B.n171 B.n170 585
R18 B.n169 B.n168 585
R19 B.n167 B.n166 585
R20 B.n165 B.n164 585
R21 B.n163 B.n162 585
R22 B.n161 B.n160 585
R23 B.n159 B.n158 585
R24 B.n157 B.n156 585
R25 B.n155 B.n154 585
R26 B.n153 B.n152 585
R27 B.n151 B.n150 585
R28 B.n149 B.n148 585
R29 B.n147 B.n146 585
R30 B.n145 B.n144 585
R31 B.n143 B.n142 585
R32 B.n141 B.n140 585
R33 B.n139 B.n138 585
R34 B.n137 B.n136 585
R35 B.n135 B.n134 585
R36 B.n133 B.n132 585
R37 B.n131 B.n130 585
R38 B.n129 B.n128 585
R39 B.n127 B.n126 585
R40 B.n125 B.n124 585
R41 B.n123 B.n122 585
R42 B.n121 B.n120 585
R43 B.n119 B.n118 585
R44 B.n117 B.n116 585
R45 B.n115 B.n114 585
R46 B.n113 B.n112 585
R47 B.n110 B.n109 585
R48 B.n108 B.n107 585
R49 B.n106 B.n105 585
R50 B.n104 B.n103 585
R51 B.n102 B.n101 585
R52 B.n100 B.n99 585
R53 B.n98 B.n97 585
R54 B.n96 B.n95 585
R55 B.n94 B.n93 585
R56 B.n92 B.n91 585
R57 B.n90 B.n89 585
R58 B.n88 B.n87 585
R59 B.n86 B.n85 585
R60 B.n84 B.n83 585
R61 B.n82 B.n81 585
R62 B.n80 B.n79 585
R63 B.n78 B.n77 585
R64 B.n76 B.n75 585
R65 B.n74 B.n73 585
R66 B.n72 B.n71 585
R67 B.n70 B.n69 585
R68 B.n68 B.n67 585
R69 B.n32 B.n31 585
R70 B.n417 B.n33 585
R71 B.n421 B.n33 585
R72 B.n416 B.n415 585
R73 B.n415 B.n29 585
R74 B.n414 B.n28 585
R75 B.n427 B.n28 585
R76 B.n413 B.n27 585
R77 B.n428 B.n27 585
R78 B.n412 B.n26 585
R79 B.n429 B.n26 585
R80 B.n411 B.n410 585
R81 B.n410 B.n25 585
R82 B.n409 B.n21 585
R83 B.n435 B.n21 585
R84 B.n408 B.n20 585
R85 B.n436 B.n20 585
R86 B.n407 B.n19 585
R87 B.n437 B.n19 585
R88 B.n406 B.n405 585
R89 B.n405 B.n15 585
R90 B.n404 B.n14 585
R91 B.n443 B.n14 585
R92 B.n403 B.n13 585
R93 B.n444 B.n13 585
R94 B.n402 B.n12 585
R95 B.n445 B.n12 585
R96 B.n401 B.n400 585
R97 B.n400 B.n399 585
R98 B.n398 B.n397 585
R99 B.n398 B.n8 585
R100 B.n396 B.n7 585
R101 B.n452 B.n7 585
R102 B.n395 B.n6 585
R103 B.n453 B.n6 585
R104 B.n394 B.n5 585
R105 B.n454 B.n5 585
R106 B.n393 B.n392 585
R107 B.n392 B.n4 585
R108 B.n391 B.n173 585
R109 B.n391 B.n390 585
R110 B.n381 B.n174 585
R111 B.n175 B.n174 585
R112 B.n383 B.n382 585
R113 B.n384 B.n383 585
R114 B.n380 B.n180 585
R115 B.n180 B.n179 585
R116 B.n379 B.n378 585
R117 B.n378 B.n377 585
R118 B.n182 B.n181 585
R119 B.n183 B.n182 585
R120 B.n370 B.n369 585
R121 B.n371 B.n370 585
R122 B.n368 B.n188 585
R123 B.n188 B.n187 585
R124 B.n367 B.n366 585
R125 B.n366 B.n365 585
R126 B.n190 B.n189 585
R127 B.n358 B.n190 585
R128 B.n357 B.n356 585
R129 B.n359 B.n357 585
R130 B.n355 B.n195 585
R131 B.n195 B.n194 585
R132 B.n354 B.n353 585
R133 B.n353 B.n352 585
R134 B.n197 B.n196 585
R135 B.n198 B.n197 585
R136 B.n345 B.n344 585
R137 B.n346 B.n345 585
R138 B.n201 B.n200 585
R139 B.n234 B.n233 585
R140 B.n235 B.n231 585
R141 B.n231 B.n202 585
R142 B.n237 B.n236 585
R143 B.n239 B.n230 585
R144 B.n242 B.n241 585
R145 B.n243 B.n229 585
R146 B.n245 B.n244 585
R147 B.n247 B.n228 585
R148 B.n250 B.n249 585
R149 B.n251 B.n227 585
R150 B.n253 B.n252 585
R151 B.n255 B.n226 585
R152 B.n258 B.n257 585
R153 B.n259 B.n225 585
R154 B.n261 B.n260 585
R155 B.n263 B.n224 585
R156 B.n266 B.n265 585
R157 B.n267 B.n223 585
R158 B.n269 B.n268 585
R159 B.n271 B.n222 585
R160 B.n274 B.n273 585
R161 B.n275 B.n219 585
R162 B.n278 B.n277 585
R163 B.n280 B.n218 585
R164 B.n283 B.n282 585
R165 B.n284 B.n217 585
R166 B.n286 B.n285 585
R167 B.n288 B.n216 585
R168 B.n291 B.n290 585
R169 B.n292 B.n215 585
R170 B.n297 B.n296 585
R171 B.n299 B.n214 585
R172 B.n302 B.n301 585
R173 B.n303 B.n213 585
R174 B.n305 B.n304 585
R175 B.n307 B.n212 585
R176 B.n310 B.n309 585
R177 B.n311 B.n211 585
R178 B.n313 B.n312 585
R179 B.n315 B.n210 585
R180 B.n318 B.n317 585
R181 B.n319 B.n209 585
R182 B.n321 B.n320 585
R183 B.n323 B.n208 585
R184 B.n326 B.n325 585
R185 B.n327 B.n207 585
R186 B.n329 B.n328 585
R187 B.n331 B.n206 585
R188 B.n334 B.n333 585
R189 B.n335 B.n205 585
R190 B.n337 B.n336 585
R191 B.n339 B.n204 585
R192 B.n342 B.n341 585
R193 B.n343 B.n203 585
R194 B.n348 B.n347 585
R195 B.n347 B.n346 585
R196 B.n349 B.n199 585
R197 B.n199 B.n198 585
R198 B.n351 B.n350 585
R199 B.n352 B.n351 585
R200 B.n193 B.n192 585
R201 B.n194 B.n193 585
R202 B.n361 B.n360 585
R203 B.n360 B.n359 585
R204 B.n362 B.n191 585
R205 B.n358 B.n191 585
R206 B.n364 B.n363 585
R207 B.n365 B.n364 585
R208 B.n186 B.n185 585
R209 B.n187 B.n186 585
R210 B.n373 B.n372 585
R211 B.n372 B.n371 585
R212 B.n374 B.n184 585
R213 B.n184 B.n183 585
R214 B.n376 B.n375 585
R215 B.n377 B.n376 585
R216 B.n178 B.n177 585
R217 B.n179 B.n178 585
R218 B.n386 B.n385 585
R219 B.n385 B.n384 585
R220 B.n387 B.n176 585
R221 B.n176 B.n175 585
R222 B.n389 B.n388 585
R223 B.n390 B.n389 585
R224 B.n3 B.n0 585
R225 B.n4 B.n3 585
R226 B.n451 B.n1 585
R227 B.n452 B.n451 585
R228 B.n450 B.n449 585
R229 B.n450 B.n8 585
R230 B.n448 B.n9 585
R231 B.n399 B.n9 585
R232 B.n447 B.n446 585
R233 B.n446 B.n445 585
R234 B.n11 B.n10 585
R235 B.n444 B.n11 585
R236 B.n442 B.n441 585
R237 B.n443 B.n442 585
R238 B.n440 B.n16 585
R239 B.n16 B.n15 585
R240 B.n439 B.n438 585
R241 B.n438 B.n437 585
R242 B.n18 B.n17 585
R243 B.n436 B.n18 585
R244 B.n434 B.n433 585
R245 B.n435 B.n434 585
R246 B.n432 B.n22 585
R247 B.n25 B.n22 585
R248 B.n431 B.n430 585
R249 B.n430 B.n429 585
R250 B.n24 B.n23 585
R251 B.n428 B.n24 585
R252 B.n426 B.n425 585
R253 B.n427 B.n426 585
R254 B.n424 B.n30 585
R255 B.n30 B.n29 585
R256 B.n423 B.n422 585
R257 B.n422 B.n421 585
R258 B.n455 B.n454 585
R259 B.n453 B.n2 585
R260 B.n422 B.n32 511.721
R261 B.n419 B.n33 511.721
R262 B.n345 B.n203 511.721
R263 B.n347 B.n201 511.721
R264 B.n65 B.t2 330.187
R265 B.n62 B.t10 330.187
R266 B.n293 B.t6 330.187
R267 B.n220 B.t13 330.187
R268 B.n420 B.n60 256.663
R269 B.n420 B.n59 256.663
R270 B.n420 B.n58 256.663
R271 B.n420 B.n57 256.663
R272 B.n420 B.n56 256.663
R273 B.n420 B.n55 256.663
R274 B.n420 B.n54 256.663
R275 B.n420 B.n53 256.663
R276 B.n420 B.n52 256.663
R277 B.n420 B.n51 256.663
R278 B.n420 B.n50 256.663
R279 B.n420 B.n49 256.663
R280 B.n420 B.n48 256.663
R281 B.n420 B.n47 256.663
R282 B.n420 B.n46 256.663
R283 B.n420 B.n45 256.663
R284 B.n420 B.n44 256.663
R285 B.n420 B.n43 256.663
R286 B.n420 B.n42 256.663
R287 B.n420 B.n41 256.663
R288 B.n420 B.n40 256.663
R289 B.n420 B.n39 256.663
R290 B.n420 B.n38 256.663
R291 B.n420 B.n37 256.663
R292 B.n420 B.n36 256.663
R293 B.n420 B.n35 256.663
R294 B.n420 B.n34 256.663
R295 B.n232 B.n202 256.663
R296 B.n238 B.n202 256.663
R297 B.n240 B.n202 256.663
R298 B.n246 B.n202 256.663
R299 B.n248 B.n202 256.663
R300 B.n254 B.n202 256.663
R301 B.n256 B.n202 256.663
R302 B.n262 B.n202 256.663
R303 B.n264 B.n202 256.663
R304 B.n270 B.n202 256.663
R305 B.n272 B.n202 256.663
R306 B.n279 B.n202 256.663
R307 B.n281 B.n202 256.663
R308 B.n287 B.n202 256.663
R309 B.n289 B.n202 256.663
R310 B.n298 B.n202 256.663
R311 B.n300 B.n202 256.663
R312 B.n306 B.n202 256.663
R313 B.n308 B.n202 256.663
R314 B.n314 B.n202 256.663
R315 B.n316 B.n202 256.663
R316 B.n322 B.n202 256.663
R317 B.n324 B.n202 256.663
R318 B.n330 B.n202 256.663
R319 B.n332 B.n202 256.663
R320 B.n338 B.n202 256.663
R321 B.n340 B.n202 256.663
R322 B.n457 B.n456 256.663
R323 B.n69 B.n68 163.367
R324 B.n73 B.n72 163.367
R325 B.n77 B.n76 163.367
R326 B.n81 B.n80 163.367
R327 B.n85 B.n84 163.367
R328 B.n89 B.n88 163.367
R329 B.n93 B.n92 163.367
R330 B.n97 B.n96 163.367
R331 B.n101 B.n100 163.367
R332 B.n105 B.n104 163.367
R333 B.n109 B.n108 163.367
R334 B.n114 B.n113 163.367
R335 B.n118 B.n117 163.367
R336 B.n122 B.n121 163.367
R337 B.n126 B.n125 163.367
R338 B.n130 B.n129 163.367
R339 B.n134 B.n133 163.367
R340 B.n138 B.n137 163.367
R341 B.n142 B.n141 163.367
R342 B.n146 B.n145 163.367
R343 B.n150 B.n149 163.367
R344 B.n154 B.n153 163.367
R345 B.n158 B.n157 163.367
R346 B.n162 B.n161 163.367
R347 B.n166 B.n165 163.367
R348 B.n170 B.n169 163.367
R349 B.n419 B.n61 163.367
R350 B.n345 B.n197 163.367
R351 B.n353 B.n197 163.367
R352 B.n353 B.n195 163.367
R353 B.n357 B.n195 163.367
R354 B.n357 B.n190 163.367
R355 B.n366 B.n190 163.367
R356 B.n366 B.n188 163.367
R357 B.n370 B.n188 163.367
R358 B.n370 B.n182 163.367
R359 B.n378 B.n182 163.367
R360 B.n378 B.n180 163.367
R361 B.n383 B.n180 163.367
R362 B.n383 B.n174 163.367
R363 B.n391 B.n174 163.367
R364 B.n392 B.n391 163.367
R365 B.n392 B.n5 163.367
R366 B.n6 B.n5 163.367
R367 B.n7 B.n6 163.367
R368 B.n398 B.n7 163.367
R369 B.n400 B.n398 163.367
R370 B.n400 B.n12 163.367
R371 B.n13 B.n12 163.367
R372 B.n14 B.n13 163.367
R373 B.n405 B.n14 163.367
R374 B.n405 B.n19 163.367
R375 B.n20 B.n19 163.367
R376 B.n21 B.n20 163.367
R377 B.n410 B.n21 163.367
R378 B.n410 B.n26 163.367
R379 B.n27 B.n26 163.367
R380 B.n28 B.n27 163.367
R381 B.n415 B.n28 163.367
R382 B.n415 B.n33 163.367
R383 B.n233 B.n231 163.367
R384 B.n237 B.n231 163.367
R385 B.n241 B.n239 163.367
R386 B.n245 B.n229 163.367
R387 B.n249 B.n247 163.367
R388 B.n253 B.n227 163.367
R389 B.n257 B.n255 163.367
R390 B.n261 B.n225 163.367
R391 B.n265 B.n263 163.367
R392 B.n269 B.n223 163.367
R393 B.n273 B.n271 163.367
R394 B.n278 B.n219 163.367
R395 B.n282 B.n280 163.367
R396 B.n286 B.n217 163.367
R397 B.n290 B.n288 163.367
R398 B.n297 B.n215 163.367
R399 B.n301 B.n299 163.367
R400 B.n305 B.n213 163.367
R401 B.n309 B.n307 163.367
R402 B.n313 B.n211 163.367
R403 B.n317 B.n315 163.367
R404 B.n321 B.n209 163.367
R405 B.n325 B.n323 163.367
R406 B.n329 B.n207 163.367
R407 B.n333 B.n331 163.367
R408 B.n337 B.n205 163.367
R409 B.n341 B.n339 163.367
R410 B.n347 B.n199 163.367
R411 B.n351 B.n199 163.367
R412 B.n351 B.n193 163.367
R413 B.n360 B.n193 163.367
R414 B.n360 B.n191 163.367
R415 B.n364 B.n191 163.367
R416 B.n364 B.n186 163.367
R417 B.n372 B.n186 163.367
R418 B.n372 B.n184 163.367
R419 B.n376 B.n184 163.367
R420 B.n376 B.n178 163.367
R421 B.n385 B.n178 163.367
R422 B.n385 B.n176 163.367
R423 B.n389 B.n176 163.367
R424 B.n389 B.n3 163.367
R425 B.n455 B.n3 163.367
R426 B.n451 B.n2 163.367
R427 B.n451 B.n450 163.367
R428 B.n450 B.n9 163.367
R429 B.n446 B.n9 163.367
R430 B.n446 B.n11 163.367
R431 B.n442 B.n11 163.367
R432 B.n442 B.n16 163.367
R433 B.n438 B.n16 163.367
R434 B.n438 B.n18 163.367
R435 B.n434 B.n18 163.367
R436 B.n434 B.n22 163.367
R437 B.n430 B.n22 163.367
R438 B.n430 B.n24 163.367
R439 B.n426 B.n24 163.367
R440 B.n426 B.n30 163.367
R441 B.n422 B.n30 163.367
R442 B.n346 B.n202 113.776
R443 B.n421 B.n420 113.776
R444 B.n62 B.t11 100.517
R445 B.n293 B.t9 100.517
R446 B.n65 B.t4 100.511
R447 B.n220 B.t15 100.511
R448 B.n63 B.t12 73.3661
R449 B.n294 B.t8 73.3661
R450 B.n66 B.t5 73.3603
R451 B.n221 B.t14 73.3603
R452 B.n34 B.n32 71.676
R453 B.n69 B.n35 71.676
R454 B.n73 B.n36 71.676
R455 B.n77 B.n37 71.676
R456 B.n81 B.n38 71.676
R457 B.n85 B.n39 71.676
R458 B.n89 B.n40 71.676
R459 B.n93 B.n41 71.676
R460 B.n97 B.n42 71.676
R461 B.n101 B.n43 71.676
R462 B.n105 B.n44 71.676
R463 B.n109 B.n45 71.676
R464 B.n114 B.n46 71.676
R465 B.n118 B.n47 71.676
R466 B.n122 B.n48 71.676
R467 B.n126 B.n49 71.676
R468 B.n130 B.n50 71.676
R469 B.n134 B.n51 71.676
R470 B.n138 B.n52 71.676
R471 B.n142 B.n53 71.676
R472 B.n146 B.n54 71.676
R473 B.n150 B.n55 71.676
R474 B.n154 B.n56 71.676
R475 B.n158 B.n57 71.676
R476 B.n162 B.n58 71.676
R477 B.n166 B.n59 71.676
R478 B.n170 B.n60 71.676
R479 B.n61 B.n60 71.676
R480 B.n169 B.n59 71.676
R481 B.n165 B.n58 71.676
R482 B.n161 B.n57 71.676
R483 B.n157 B.n56 71.676
R484 B.n153 B.n55 71.676
R485 B.n149 B.n54 71.676
R486 B.n145 B.n53 71.676
R487 B.n141 B.n52 71.676
R488 B.n137 B.n51 71.676
R489 B.n133 B.n50 71.676
R490 B.n129 B.n49 71.676
R491 B.n125 B.n48 71.676
R492 B.n121 B.n47 71.676
R493 B.n117 B.n46 71.676
R494 B.n113 B.n45 71.676
R495 B.n108 B.n44 71.676
R496 B.n104 B.n43 71.676
R497 B.n100 B.n42 71.676
R498 B.n96 B.n41 71.676
R499 B.n92 B.n40 71.676
R500 B.n88 B.n39 71.676
R501 B.n84 B.n38 71.676
R502 B.n80 B.n37 71.676
R503 B.n76 B.n36 71.676
R504 B.n72 B.n35 71.676
R505 B.n68 B.n34 71.676
R506 B.n232 B.n201 71.676
R507 B.n238 B.n237 71.676
R508 B.n241 B.n240 71.676
R509 B.n246 B.n245 71.676
R510 B.n249 B.n248 71.676
R511 B.n254 B.n253 71.676
R512 B.n257 B.n256 71.676
R513 B.n262 B.n261 71.676
R514 B.n265 B.n264 71.676
R515 B.n270 B.n269 71.676
R516 B.n273 B.n272 71.676
R517 B.n279 B.n278 71.676
R518 B.n282 B.n281 71.676
R519 B.n287 B.n286 71.676
R520 B.n290 B.n289 71.676
R521 B.n298 B.n297 71.676
R522 B.n301 B.n300 71.676
R523 B.n306 B.n305 71.676
R524 B.n309 B.n308 71.676
R525 B.n314 B.n313 71.676
R526 B.n317 B.n316 71.676
R527 B.n322 B.n321 71.676
R528 B.n325 B.n324 71.676
R529 B.n330 B.n329 71.676
R530 B.n333 B.n332 71.676
R531 B.n338 B.n337 71.676
R532 B.n341 B.n340 71.676
R533 B.n233 B.n232 71.676
R534 B.n239 B.n238 71.676
R535 B.n240 B.n229 71.676
R536 B.n247 B.n246 71.676
R537 B.n248 B.n227 71.676
R538 B.n255 B.n254 71.676
R539 B.n256 B.n225 71.676
R540 B.n263 B.n262 71.676
R541 B.n264 B.n223 71.676
R542 B.n271 B.n270 71.676
R543 B.n272 B.n219 71.676
R544 B.n280 B.n279 71.676
R545 B.n281 B.n217 71.676
R546 B.n288 B.n287 71.676
R547 B.n289 B.n215 71.676
R548 B.n299 B.n298 71.676
R549 B.n300 B.n213 71.676
R550 B.n307 B.n306 71.676
R551 B.n308 B.n211 71.676
R552 B.n315 B.n314 71.676
R553 B.n316 B.n209 71.676
R554 B.n323 B.n322 71.676
R555 B.n324 B.n207 71.676
R556 B.n331 B.n330 71.676
R557 B.n332 B.n205 71.676
R558 B.n339 B.n338 71.676
R559 B.n340 B.n203 71.676
R560 B.n456 B.n455 71.676
R561 B.n456 B.n2 71.676
R562 B.n346 B.n198 68.4673
R563 B.n352 B.n198 68.4673
R564 B.n352 B.n194 68.4673
R565 B.n359 B.n194 68.4673
R566 B.n359 B.n358 68.4673
R567 B.n365 B.n187 68.4673
R568 B.n371 B.n187 68.4673
R569 B.n371 B.n183 68.4673
R570 B.n377 B.n183 68.4673
R571 B.n377 B.n179 68.4673
R572 B.n384 B.n179 68.4673
R573 B.n390 B.n175 68.4673
R574 B.n390 B.n4 68.4673
R575 B.n454 B.n4 68.4673
R576 B.n454 B.n453 68.4673
R577 B.n453 B.n452 68.4673
R578 B.n452 B.n8 68.4673
R579 B.n399 B.n8 68.4673
R580 B.n445 B.n444 68.4673
R581 B.n444 B.n443 68.4673
R582 B.n443 B.n15 68.4673
R583 B.n437 B.n15 68.4673
R584 B.n437 B.n436 68.4673
R585 B.n436 B.n435 68.4673
R586 B.n429 B.n25 68.4673
R587 B.n429 B.n428 68.4673
R588 B.n428 B.n427 68.4673
R589 B.n427 B.n29 68.4673
R590 B.n421 B.n29 68.4673
R591 B.n111 B.n66 59.5399
R592 B.n64 B.n63 59.5399
R593 B.n295 B.n294 59.5399
R594 B.n276 B.n221 59.5399
R595 B.n384 B.t0 57.3918
R596 B.n445 B.t1 57.3918
R597 B.n358 B.t7 35.2408
R598 B.n25 B.t3 35.2408
R599 B.n348 B.n200 33.2493
R600 B.n344 B.n343 33.2493
R601 B.n418 B.n417 33.2493
R602 B.n423 B.n31 33.2493
R603 B.n365 B.t7 33.227
R604 B.n435 B.t3 33.227
R605 B.n66 B.n65 27.152
R606 B.n63 B.n62 27.152
R607 B.n294 B.n293 27.152
R608 B.n221 B.n220 27.152
R609 B B.n457 18.0485
R610 B.t0 B.n175 11.076
R611 B.n399 B.t1 11.076
R612 B.n349 B.n348 10.6151
R613 B.n350 B.n349 10.6151
R614 B.n350 B.n192 10.6151
R615 B.n361 B.n192 10.6151
R616 B.n362 B.n361 10.6151
R617 B.n363 B.n362 10.6151
R618 B.n363 B.n185 10.6151
R619 B.n373 B.n185 10.6151
R620 B.n374 B.n373 10.6151
R621 B.n375 B.n374 10.6151
R622 B.n375 B.n177 10.6151
R623 B.n386 B.n177 10.6151
R624 B.n387 B.n386 10.6151
R625 B.n388 B.n387 10.6151
R626 B.n388 B.n0 10.6151
R627 B.n234 B.n200 10.6151
R628 B.n235 B.n234 10.6151
R629 B.n236 B.n235 10.6151
R630 B.n236 B.n230 10.6151
R631 B.n242 B.n230 10.6151
R632 B.n243 B.n242 10.6151
R633 B.n244 B.n243 10.6151
R634 B.n244 B.n228 10.6151
R635 B.n250 B.n228 10.6151
R636 B.n251 B.n250 10.6151
R637 B.n252 B.n251 10.6151
R638 B.n252 B.n226 10.6151
R639 B.n258 B.n226 10.6151
R640 B.n259 B.n258 10.6151
R641 B.n260 B.n259 10.6151
R642 B.n260 B.n224 10.6151
R643 B.n266 B.n224 10.6151
R644 B.n267 B.n266 10.6151
R645 B.n268 B.n267 10.6151
R646 B.n268 B.n222 10.6151
R647 B.n274 B.n222 10.6151
R648 B.n275 B.n274 10.6151
R649 B.n277 B.n218 10.6151
R650 B.n283 B.n218 10.6151
R651 B.n284 B.n283 10.6151
R652 B.n285 B.n284 10.6151
R653 B.n285 B.n216 10.6151
R654 B.n291 B.n216 10.6151
R655 B.n292 B.n291 10.6151
R656 B.n296 B.n292 10.6151
R657 B.n302 B.n214 10.6151
R658 B.n303 B.n302 10.6151
R659 B.n304 B.n303 10.6151
R660 B.n304 B.n212 10.6151
R661 B.n310 B.n212 10.6151
R662 B.n311 B.n310 10.6151
R663 B.n312 B.n311 10.6151
R664 B.n312 B.n210 10.6151
R665 B.n318 B.n210 10.6151
R666 B.n319 B.n318 10.6151
R667 B.n320 B.n319 10.6151
R668 B.n320 B.n208 10.6151
R669 B.n326 B.n208 10.6151
R670 B.n327 B.n326 10.6151
R671 B.n328 B.n327 10.6151
R672 B.n328 B.n206 10.6151
R673 B.n334 B.n206 10.6151
R674 B.n335 B.n334 10.6151
R675 B.n336 B.n335 10.6151
R676 B.n336 B.n204 10.6151
R677 B.n342 B.n204 10.6151
R678 B.n343 B.n342 10.6151
R679 B.n344 B.n196 10.6151
R680 B.n354 B.n196 10.6151
R681 B.n355 B.n354 10.6151
R682 B.n356 B.n355 10.6151
R683 B.n356 B.n189 10.6151
R684 B.n367 B.n189 10.6151
R685 B.n368 B.n367 10.6151
R686 B.n369 B.n368 10.6151
R687 B.n369 B.n181 10.6151
R688 B.n379 B.n181 10.6151
R689 B.n380 B.n379 10.6151
R690 B.n382 B.n380 10.6151
R691 B.n382 B.n381 10.6151
R692 B.n381 B.n173 10.6151
R693 B.n393 B.n173 10.6151
R694 B.n394 B.n393 10.6151
R695 B.n395 B.n394 10.6151
R696 B.n396 B.n395 10.6151
R697 B.n397 B.n396 10.6151
R698 B.n401 B.n397 10.6151
R699 B.n402 B.n401 10.6151
R700 B.n403 B.n402 10.6151
R701 B.n404 B.n403 10.6151
R702 B.n406 B.n404 10.6151
R703 B.n407 B.n406 10.6151
R704 B.n408 B.n407 10.6151
R705 B.n409 B.n408 10.6151
R706 B.n411 B.n409 10.6151
R707 B.n412 B.n411 10.6151
R708 B.n413 B.n412 10.6151
R709 B.n414 B.n413 10.6151
R710 B.n416 B.n414 10.6151
R711 B.n417 B.n416 10.6151
R712 B.n449 B.n1 10.6151
R713 B.n449 B.n448 10.6151
R714 B.n448 B.n447 10.6151
R715 B.n447 B.n10 10.6151
R716 B.n441 B.n10 10.6151
R717 B.n441 B.n440 10.6151
R718 B.n440 B.n439 10.6151
R719 B.n439 B.n17 10.6151
R720 B.n433 B.n17 10.6151
R721 B.n433 B.n432 10.6151
R722 B.n432 B.n431 10.6151
R723 B.n431 B.n23 10.6151
R724 B.n425 B.n23 10.6151
R725 B.n425 B.n424 10.6151
R726 B.n424 B.n423 10.6151
R727 B.n67 B.n31 10.6151
R728 B.n70 B.n67 10.6151
R729 B.n71 B.n70 10.6151
R730 B.n74 B.n71 10.6151
R731 B.n75 B.n74 10.6151
R732 B.n78 B.n75 10.6151
R733 B.n79 B.n78 10.6151
R734 B.n82 B.n79 10.6151
R735 B.n83 B.n82 10.6151
R736 B.n86 B.n83 10.6151
R737 B.n87 B.n86 10.6151
R738 B.n90 B.n87 10.6151
R739 B.n91 B.n90 10.6151
R740 B.n94 B.n91 10.6151
R741 B.n95 B.n94 10.6151
R742 B.n98 B.n95 10.6151
R743 B.n99 B.n98 10.6151
R744 B.n102 B.n99 10.6151
R745 B.n103 B.n102 10.6151
R746 B.n106 B.n103 10.6151
R747 B.n107 B.n106 10.6151
R748 B.n110 B.n107 10.6151
R749 B.n115 B.n112 10.6151
R750 B.n116 B.n115 10.6151
R751 B.n119 B.n116 10.6151
R752 B.n120 B.n119 10.6151
R753 B.n123 B.n120 10.6151
R754 B.n124 B.n123 10.6151
R755 B.n127 B.n124 10.6151
R756 B.n128 B.n127 10.6151
R757 B.n132 B.n131 10.6151
R758 B.n135 B.n132 10.6151
R759 B.n136 B.n135 10.6151
R760 B.n139 B.n136 10.6151
R761 B.n140 B.n139 10.6151
R762 B.n143 B.n140 10.6151
R763 B.n144 B.n143 10.6151
R764 B.n147 B.n144 10.6151
R765 B.n148 B.n147 10.6151
R766 B.n151 B.n148 10.6151
R767 B.n152 B.n151 10.6151
R768 B.n155 B.n152 10.6151
R769 B.n156 B.n155 10.6151
R770 B.n159 B.n156 10.6151
R771 B.n160 B.n159 10.6151
R772 B.n163 B.n160 10.6151
R773 B.n164 B.n163 10.6151
R774 B.n167 B.n164 10.6151
R775 B.n168 B.n167 10.6151
R776 B.n171 B.n168 10.6151
R777 B.n172 B.n171 10.6151
R778 B.n418 B.n172 10.6151
R779 B.n457 B.n0 8.11757
R780 B.n457 B.n1 8.11757
R781 B.n277 B.n276 7.18099
R782 B.n296 B.n295 7.18099
R783 B.n112 B.n111 7.18099
R784 B.n128 B.n64 7.18099
R785 B.n276 B.n275 3.43465
R786 B.n295 B.n214 3.43465
R787 B.n111 B.n110 3.43465
R788 B.n131 B.n64 3.43465
R789 VP.n0 VP.t1 360.834
R790 VP.n0 VP.t0 325.046
R791 VP VP.n0 0.0516364
R792 VDD1 VDD1.t1 102.963
R793 VDD1 VDD1.t0 71.5527
C0 VDD1 VTAIL 3.18385f
C1 VDD2 VTAIL 3.22434f
C2 VTAIL VN 1.07408f
C3 VTAIL VP 1.08838f
C4 VDD1 VDD2 0.497961f
C5 VDD1 VN 0.148757f
C6 VDD1 VP 1.31901f
C7 VDD2 VN 1.20013f
C8 VDD2 VP 0.269547f
C9 VP VN 3.54919f
C10 VDD2 B 2.721385f
C11 VDD1 B 4.39816f
C12 VTAIL B 3.978227f
C13 VN B 6.15285f
C14 VP B 3.97049f
C15 VDD1.t0 B 0.693815f
C16 VDD1.t1 B 0.9251f
C17 VP.t1 B 0.761422f
C18 VP.t0 B 0.654283f
C19 VP.n0 B 2.06673f
C20 VDD2.t0 B 0.92504f
C21 VDD2.t1 B 0.704996f
C22 VDD2.n0 B 1.52273f
C23 VTAIL.t0 B 0.741448f
C24 VTAIL.n0 B 0.878245f
C25 VTAIL.t2 B 0.741451f
C26 VTAIL.n1 B 0.891568f
C27 VTAIL.t1 B 0.741448f
C28 VTAIL.n2 B 0.825533f
C29 VTAIL.t3 B 0.741448f
C30 VTAIL.n3 B 0.780132f
C31 VN.t1 B 0.646395f
C32 VN.t0 B 0.755228f
.ends

