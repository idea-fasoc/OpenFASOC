* NGSPICE file created from diff_pair_sample_0031.ext - technology: sky130A

.subckt diff_pair_sample_0031 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t7 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=3.37
X1 VDD2.t7 VN.t0 VTAIL.t0 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X2 VTAIL.t12 VP.t1 VDD1.t6 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X3 VTAIL.t1 VN.t1 VDD2.t6 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=3.37
X4 B.t11 B.t9 B.t10 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=3.37
X5 VTAIL.t2 VN.t2 VDD2.t5 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X6 B.t8 B.t6 B.t7 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=3.37
X7 VTAIL.t14 VN.t3 VDD2.t4 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X8 VDD2.t3 VN.t4 VTAIL.t13 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=3.37
X9 B.t5 B.t3 B.t4 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=3.37
X10 VDD1.t5 VP.t2 VTAIL.t9 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X11 VDD1.t4 VP.t3 VTAIL.t6 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X12 VDD2.t2 VN.t5 VTAIL.t4 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X13 VDD1.t3 VP.t4 VTAIL.t10 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=3.37
X14 B.t2 B.t0 B.t1 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=0 ps=0 w=10.43 l=3.37
X15 VTAIL.t5 VP.t5 VDD1.t2 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=3.37
X16 VTAIL.t15 VN.t6 VDD2.t1 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=3.37
X17 VTAIL.t8 VP.t6 VDD1.t1 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=4.0677 pd=21.64 as=1.72095 ps=10.76 w=10.43 l=3.37
X18 VTAIL.t11 VP.t7 VDD1.t0 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=1.72095 ps=10.76 w=10.43 l=3.37
X19 VDD2.t0 VN.t7 VTAIL.t3 w_n4670_n3054# sky130_fd_pr__pfet_01v8 ad=1.72095 pd=10.76 as=4.0677 ps=21.64 w=10.43 l=3.37
R0 VP.n24 VP.n21 161.3
R1 VP.n26 VP.n25 161.3
R2 VP.n27 VP.n20 161.3
R3 VP.n29 VP.n28 161.3
R4 VP.n30 VP.n19 161.3
R5 VP.n32 VP.n31 161.3
R6 VP.n33 VP.n18 161.3
R7 VP.n35 VP.n34 161.3
R8 VP.n37 VP.n36 161.3
R9 VP.n38 VP.n16 161.3
R10 VP.n40 VP.n39 161.3
R11 VP.n41 VP.n15 161.3
R12 VP.n43 VP.n42 161.3
R13 VP.n44 VP.n14 161.3
R14 VP.n46 VP.n45 161.3
R15 VP.n83 VP.n82 161.3
R16 VP.n81 VP.n1 161.3
R17 VP.n80 VP.n79 161.3
R18 VP.n78 VP.n2 161.3
R19 VP.n77 VP.n76 161.3
R20 VP.n75 VP.n3 161.3
R21 VP.n74 VP.n73 161.3
R22 VP.n72 VP.n71 161.3
R23 VP.n70 VP.n5 161.3
R24 VP.n69 VP.n68 161.3
R25 VP.n67 VP.n6 161.3
R26 VP.n66 VP.n65 161.3
R27 VP.n64 VP.n7 161.3
R28 VP.n63 VP.n62 161.3
R29 VP.n61 VP.n8 161.3
R30 VP.n60 VP.n59 161.3
R31 VP.n57 VP.n9 161.3
R32 VP.n56 VP.n55 161.3
R33 VP.n54 VP.n10 161.3
R34 VP.n53 VP.n52 161.3
R35 VP.n51 VP.n11 161.3
R36 VP.n50 VP.n49 161.3
R37 VP.n23 VP.t5 107.442
R38 VP.n48 VP.n12 75.3872
R39 VP.n84 VP.n0 75.3872
R40 VP.n47 VP.n13 75.3872
R41 VP.n12 VP.t6 74.5889
R42 VP.n58 VP.t2 74.5889
R43 VP.n4 VP.t7 74.5889
R44 VP.n0 VP.t4 74.5889
R45 VP.n13 VP.t0 74.5889
R46 VP.n17 VP.t1 74.5889
R47 VP.n22 VP.t3 74.5889
R48 VP.n23 VP.n22 69.6868
R49 VP.n65 VP.n6 56.5193
R50 VP.n28 VP.n19 56.5193
R51 VP.n48 VP.n47 53.4387
R52 VP.n56 VP.n10 45.3497
R53 VP.n76 VP.n2 45.3497
R54 VP.n39 VP.n15 45.3497
R55 VP.n52 VP.n10 35.6371
R56 VP.n80 VP.n2 35.6371
R57 VP.n43 VP.n15 35.6371
R58 VP.n51 VP.n50 24.4675
R59 VP.n52 VP.n51 24.4675
R60 VP.n57 VP.n56 24.4675
R61 VP.n59 VP.n57 24.4675
R62 VP.n63 VP.n8 24.4675
R63 VP.n64 VP.n63 24.4675
R64 VP.n65 VP.n64 24.4675
R65 VP.n69 VP.n6 24.4675
R66 VP.n70 VP.n69 24.4675
R67 VP.n71 VP.n70 24.4675
R68 VP.n75 VP.n74 24.4675
R69 VP.n76 VP.n75 24.4675
R70 VP.n81 VP.n80 24.4675
R71 VP.n82 VP.n81 24.4675
R72 VP.n44 VP.n43 24.4675
R73 VP.n45 VP.n44 24.4675
R74 VP.n32 VP.n19 24.4675
R75 VP.n33 VP.n32 24.4675
R76 VP.n34 VP.n33 24.4675
R77 VP.n38 VP.n37 24.4675
R78 VP.n39 VP.n38 24.4675
R79 VP.n26 VP.n21 24.4675
R80 VP.n27 VP.n26 24.4675
R81 VP.n28 VP.n27 24.4675
R82 VP.n59 VP.n58 19.5741
R83 VP.n74 VP.n4 19.5741
R84 VP.n37 VP.n17 19.5741
R85 VP.n50 VP.n12 14.6807
R86 VP.n82 VP.n0 14.6807
R87 VP.n45 VP.n13 14.6807
R88 VP.n58 VP.n8 4.8939
R89 VP.n71 VP.n4 4.8939
R90 VP.n34 VP.n17 4.8939
R91 VP.n22 VP.n21 4.8939
R92 VP.n24 VP.n23 4.16574
R93 VP.n47 VP.n46 0.354971
R94 VP.n49 VP.n48 0.354971
R95 VP.n84 VP.n83 0.354971
R96 VP VP.n84 0.26696
R97 VP.n25 VP.n24 0.189894
R98 VP.n25 VP.n20 0.189894
R99 VP.n29 VP.n20 0.189894
R100 VP.n30 VP.n29 0.189894
R101 VP.n31 VP.n30 0.189894
R102 VP.n31 VP.n18 0.189894
R103 VP.n35 VP.n18 0.189894
R104 VP.n36 VP.n35 0.189894
R105 VP.n36 VP.n16 0.189894
R106 VP.n40 VP.n16 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n14 0.189894
R110 VP.n46 VP.n14 0.189894
R111 VP.n49 VP.n11 0.189894
R112 VP.n53 VP.n11 0.189894
R113 VP.n54 VP.n53 0.189894
R114 VP.n55 VP.n54 0.189894
R115 VP.n55 VP.n9 0.189894
R116 VP.n60 VP.n9 0.189894
R117 VP.n61 VP.n60 0.189894
R118 VP.n62 VP.n61 0.189894
R119 VP.n62 VP.n7 0.189894
R120 VP.n66 VP.n7 0.189894
R121 VP.n67 VP.n66 0.189894
R122 VP.n68 VP.n67 0.189894
R123 VP.n68 VP.n5 0.189894
R124 VP.n72 VP.n5 0.189894
R125 VP.n73 VP.n72 0.189894
R126 VP.n73 VP.n3 0.189894
R127 VP.n77 VP.n3 0.189894
R128 VP.n78 VP.n77 0.189894
R129 VP.n79 VP.n78 0.189894
R130 VP.n79 VP.n1 0.189894
R131 VP.n83 VP.n1 0.189894
R132 VTAIL.n11 VTAIL.t5 65.0397
R133 VTAIL.n10 VTAIL.t13 65.0397
R134 VTAIL.n7 VTAIL.t1 65.0397
R135 VTAIL.n14 VTAIL.t7 65.0395
R136 VTAIL.n15 VTAIL.t3 65.0395
R137 VTAIL.n2 VTAIL.t15 65.0395
R138 VTAIL.n3 VTAIL.t10 65.0395
R139 VTAIL.n6 VTAIL.t8 65.0395
R140 VTAIL.n13 VTAIL.n12 61.9232
R141 VTAIL.n9 VTAIL.n8 61.9232
R142 VTAIL.n1 VTAIL.n0 61.923
R143 VTAIL.n5 VTAIL.n4 61.923
R144 VTAIL.n15 VTAIL.n14 24.5479
R145 VTAIL.n7 VTAIL.n6 24.5479
R146 VTAIL.n9 VTAIL.n7 3.19016
R147 VTAIL.n10 VTAIL.n9 3.19016
R148 VTAIL.n13 VTAIL.n11 3.19016
R149 VTAIL.n14 VTAIL.n13 3.19016
R150 VTAIL.n6 VTAIL.n5 3.19016
R151 VTAIL.n5 VTAIL.n3 3.19016
R152 VTAIL.n2 VTAIL.n1 3.19016
R153 VTAIL VTAIL.n15 3.13197
R154 VTAIL.n0 VTAIL.t0 3.11699
R155 VTAIL.n0 VTAIL.t14 3.11699
R156 VTAIL.n4 VTAIL.t9 3.11699
R157 VTAIL.n4 VTAIL.t11 3.11699
R158 VTAIL.n12 VTAIL.t6 3.11699
R159 VTAIL.n12 VTAIL.t12 3.11699
R160 VTAIL.n8 VTAIL.t4 3.11699
R161 VTAIL.n8 VTAIL.t2 3.11699
R162 VTAIL.n11 VTAIL.n10 0.470328
R163 VTAIL.n3 VTAIL.n2 0.470328
R164 VTAIL VTAIL.n1 0.0586897
R165 VDD1 VDD1.n0 80.255
R166 VDD1.n3 VDD1.n2 80.1413
R167 VDD1.n3 VDD1.n1 80.1413
R168 VDD1.n5 VDD1.n4 78.6018
R169 VDD1.n5 VDD1.n3 47.6431
R170 VDD1.n4 VDD1.t6 3.11699
R171 VDD1.n4 VDD1.t7 3.11699
R172 VDD1.n0 VDD1.t2 3.11699
R173 VDD1.n0 VDD1.t4 3.11699
R174 VDD1.n2 VDD1.t0 3.11699
R175 VDD1.n2 VDD1.t3 3.11699
R176 VDD1.n1 VDD1.t1 3.11699
R177 VDD1.n1 VDD1.t5 3.11699
R178 VDD1 VDD1.n5 1.53714
R179 VN.n68 VN.n67 161.3
R180 VN.n66 VN.n36 161.3
R181 VN.n65 VN.n64 161.3
R182 VN.n63 VN.n37 161.3
R183 VN.n62 VN.n61 161.3
R184 VN.n60 VN.n38 161.3
R185 VN.n59 VN.n58 161.3
R186 VN.n57 VN.n56 161.3
R187 VN.n55 VN.n40 161.3
R188 VN.n54 VN.n53 161.3
R189 VN.n52 VN.n41 161.3
R190 VN.n51 VN.n50 161.3
R191 VN.n49 VN.n42 161.3
R192 VN.n48 VN.n47 161.3
R193 VN.n46 VN.n43 161.3
R194 VN.n33 VN.n32 161.3
R195 VN.n31 VN.n1 161.3
R196 VN.n30 VN.n29 161.3
R197 VN.n28 VN.n2 161.3
R198 VN.n27 VN.n26 161.3
R199 VN.n25 VN.n3 161.3
R200 VN.n24 VN.n23 161.3
R201 VN.n22 VN.n21 161.3
R202 VN.n20 VN.n5 161.3
R203 VN.n19 VN.n18 161.3
R204 VN.n17 VN.n6 161.3
R205 VN.n16 VN.n15 161.3
R206 VN.n14 VN.n7 161.3
R207 VN.n13 VN.n12 161.3
R208 VN.n11 VN.n8 161.3
R209 VN.n10 VN.t6 107.444
R210 VN.n45 VN.t4 107.444
R211 VN.n34 VN.n0 75.3872
R212 VN.n69 VN.n35 75.3872
R213 VN.n9 VN.t0 74.5889
R214 VN.n4 VN.t3 74.5889
R215 VN.n0 VN.t7 74.5889
R216 VN.n44 VN.t2 74.5889
R217 VN.n39 VN.t5 74.5889
R218 VN.n35 VN.t1 74.5889
R219 VN.n10 VN.n9 69.6868
R220 VN.n45 VN.n44 69.6868
R221 VN.n15 VN.n6 56.5193
R222 VN.n50 VN.n41 56.5193
R223 VN VN.n69 53.6041
R224 VN.n26 VN.n2 45.3497
R225 VN.n61 VN.n37 45.3497
R226 VN.n30 VN.n2 35.6371
R227 VN.n65 VN.n37 35.6371
R228 VN.n13 VN.n8 24.4675
R229 VN.n14 VN.n13 24.4675
R230 VN.n15 VN.n14 24.4675
R231 VN.n19 VN.n6 24.4675
R232 VN.n20 VN.n19 24.4675
R233 VN.n21 VN.n20 24.4675
R234 VN.n25 VN.n24 24.4675
R235 VN.n26 VN.n25 24.4675
R236 VN.n31 VN.n30 24.4675
R237 VN.n32 VN.n31 24.4675
R238 VN.n50 VN.n49 24.4675
R239 VN.n49 VN.n48 24.4675
R240 VN.n48 VN.n43 24.4675
R241 VN.n61 VN.n60 24.4675
R242 VN.n60 VN.n59 24.4675
R243 VN.n56 VN.n55 24.4675
R244 VN.n55 VN.n54 24.4675
R245 VN.n54 VN.n41 24.4675
R246 VN.n67 VN.n66 24.4675
R247 VN.n66 VN.n65 24.4675
R248 VN.n24 VN.n4 19.5741
R249 VN.n59 VN.n39 19.5741
R250 VN.n32 VN.n0 14.6807
R251 VN.n67 VN.n35 14.6807
R252 VN.n9 VN.n8 4.8939
R253 VN.n21 VN.n4 4.8939
R254 VN.n44 VN.n43 4.8939
R255 VN.n56 VN.n39 4.8939
R256 VN.n11 VN.n10 4.16576
R257 VN.n46 VN.n45 4.16576
R258 VN.n69 VN.n68 0.354971
R259 VN.n34 VN.n33 0.354971
R260 VN VN.n34 0.26696
R261 VN.n68 VN.n36 0.189894
R262 VN.n64 VN.n36 0.189894
R263 VN.n64 VN.n63 0.189894
R264 VN.n63 VN.n62 0.189894
R265 VN.n62 VN.n38 0.189894
R266 VN.n58 VN.n38 0.189894
R267 VN.n58 VN.n57 0.189894
R268 VN.n57 VN.n40 0.189894
R269 VN.n53 VN.n40 0.189894
R270 VN.n53 VN.n52 0.189894
R271 VN.n52 VN.n51 0.189894
R272 VN.n51 VN.n42 0.189894
R273 VN.n47 VN.n42 0.189894
R274 VN.n47 VN.n46 0.189894
R275 VN.n12 VN.n11 0.189894
R276 VN.n12 VN.n7 0.189894
R277 VN.n16 VN.n7 0.189894
R278 VN.n17 VN.n16 0.189894
R279 VN.n18 VN.n17 0.189894
R280 VN.n18 VN.n5 0.189894
R281 VN.n22 VN.n5 0.189894
R282 VN.n23 VN.n22 0.189894
R283 VN.n23 VN.n3 0.189894
R284 VN.n27 VN.n3 0.189894
R285 VN.n28 VN.n27 0.189894
R286 VN.n29 VN.n28 0.189894
R287 VN.n29 VN.n1 0.189894
R288 VN.n33 VN.n1 0.189894
R289 VDD2.n2 VDD2.n1 80.1413
R290 VDD2.n2 VDD2.n0 80.1413
R291 VDD2 VDD2.n5 80.1385
R292 VDD2.n4 VDD2.n3 78.602
R293 VDD2.n4 VDD2.n2 47.0601
R294 VDD2.n5 VDD2.t5 3.11699
R295 VDD2.n5 VDD2.t3 3.11699
R296 VDD2.n3 VDD2.t6 3.11699
R297 VDD2.n3 VDD2.t2 3.11699
R298 VDD2.n1 VDD2.t4 3.11699
R299 VDD2.n1 VDD2.t0 3.11699
R300 VDD2.n0 VDD2.t1 3.11699
R301 VDD2.n0 VDD2.t7 3.11699
R302 VDD2 VDD2.n4 1.65352
R303 B.n438 B.n143 585
R304 B.n437 B.n436 585
R305 B.n435 B.n144 585
R306 B.n434 B.n433 585
R307 B.n432 B.n145 585
R308 B.n431 B.n430 585
R309 B.n429 B.n146 585
R310 B.n428 B.n427 585
R311 B.n426 B.n147 585
R312 B.n425 B.n424 585
R313 B.n423 B.n148 585
R314 B.n422 B.n421 585
R315 B.n420 B.n149 585
R316 B.n419 B.n418 585
R317 B.n417 B.n150 585
R318 B.n416 B.n415 585
R319 B.n414 B.n151 585
R320 B.n413 B.n412 585
R321 B.n411 B.n152 585
R322 B.n410 B.n409 585
R323 B.n408 B.n153 585
R324 B.n407 B.n406 585
R325 B.n405 B.n154 585
R326 B.n404 B.n403 585
R327 B.n402 B.n155 585
R328 B.n401 B.n400 585
R329 B.n399 B.n156 585
R330 B.n398 B.n397 585
R331 B.n396 B.n157 585
R332 B.n395 B.n394 585
R333 B.n393 B.n158 585
R334 B.n392 B.n391 585
R335 B.n390 B.n159 585
R336 B.n389 B.n388 585
R337 B.n387 B.n160 585
R338 B.n386 B.n385 585
R339 B.n384 B.n161 585
R340 B.n383 B.n382 585
R341 B.n378 B.n162 585
R342 B.n377 B.n376 585
R343 B.n375 B.n163 585
R344 B.n374 B.n373 585
R345 B.n372 B.n164 585
R346 B.n371 B.n370 585
R347 B.n369 B.n165 585
R348 B.n368 B.n367 585
R349 B.n366 B.n166 585
R350 B.n364 B.n363 585
R351 B.n362 B.n169 585
R352 B.n361 B.n360 585
R353 B.n359 B.n170 585
R354 B.n358 B.n357 585
R355 B.n356 B.n171 585
R356 B.n355 B.n354 585
R357 B.n353 B.n172 585
R358 B.n352 B.n351 585
R359 B.n350 B.n173 585
R360 B.n349 B.n348 585
R361 B.n347 B.n174 585
R362 B.n346 B.n345 585
R363 B.n344 B.n175 585
R364 B.n343 B.n342 585
R365 B.n341 B.n176 585
R366 B.n340 B.n339 585
R367 B.n338 B.n177 585
R368 B.n337 B.n336 585
R369 B.n335 B.n178 585
R370 B.n334 B.n333 585
R371 B.n332 B.n179 585
R372 B.n331 B.n330 585
R373 B.n329 B.n180 585
R374 B.n328 B.n327 585
R375 B.n326 B.n181 585
R376 B.n325 B.n324 585
R377 B.n323 B.n182 585
R378 B.n322 B.n321 585
R379 B.n320 B.n183 585
R380 B.n319 B.n318 585
R381 B.n317 B.n184 585
R382 B.n316 B.n315 585
R383 B.n314 B.n185 585
R384 B.n313 B.n312 585
R385 B.n311 B.n186 585
R386 B.n310 B.n309 585
R387 B.n440 B.n439 585
R388 B.n441 B.n142 585
R389 B.n443 B.n442 585
R390 B.n444 B.n141 585
R391 B.n446 B.n445 585
R392 B.n447 B.n140 585
R393 B.n449 B.n448 585
R394 B.n450 B.n139 585
R395 B.n452 B.n451 585
R396 B.n453 B.n138 585
R397 B.n455 B.n454 585
R398 B.n456 B.n137 585
R399 B.n458 B.n457 585
R400 B.n459 B.n136 585
R401 B.n461 B.n460 585
R402 B.n462 B.n135 585
R403 B.n464 B.n463 585
R404 B.n465 B.n134 585
R405 B.n467 B.n466 585
R406 B.n468 B.n133 585
R407 B.n470 B.n469 585
R408 B.n471 B.n132 585
R409 B.n473 B.n472 585
R410 B.n474 B.n131 585
R411 B.n476 B.n475 585
R412 B.n477 B.n130 585
R413 B.n479 B.n478 585
R414 B.n480 B.n129 585
R415 B.n482 B.n481 585
R416 B.n483 B.n128 585
R417 B.n485 B.n484 585
R418 B.n486 B.n127 585
R419 B.n488 B.n487 585
R420 B.n489 B.n126 585
R421 B.n491 B.n490 585
R422 B.n492 B.n125 585
R423 B.n494 B.n493 585
R424 B.n495 B.n124 585
R425 B.n497 B.n496 585
R426 B.n498 B.n123 585
R427 B.n500 B.n499 585
R428 B.n501 B.n122 585
R429 B.n503 B.n502 585
R430 B.n504 B.n121 585
R431 B.n506 B.n505 585
R432 B.n507 B.n120 585
R433 B.n509 B.n508 585
R434 B.n510 B.n119 585
R435 B.n512 B.n511 585
R436 B.n513 B.n118 585
R437 B.n515 B.n514 585
R438 B.n516 B.n117 585
R439 B.n518 B.n517 585
R440 B.n519 B.n116 585
R441 B.n521 B.n520 585
R442 B.n522 B.n115 585
R443 B.n524 B.n523 585
R444 B.n525 B.n114 585
R445 B.n527 B.n526 585
R446 B.n528 B.n113 585
R447 B.n530 B.n529 585
R448 B.n531 B.n112 585
R449 B.n533 B.n532 585
R450 B.n534 B.n111 585
R451 B.n536 B.n535 585
R452 B.n537 B.n110 585
R453 B.n539 B.n538 585
R454 B.n540 B.n109 585
R455 B.n542 B.n541 585
R456 B.n543 B.n108 585
R457 B.n545 B.n544 585
R458 B.n546 B.n107 585
R459 B.n548 B.n547 585
R460 B.n549 B.n106 585
R461 B.n551 B.n550 585
R462 B.n552 B.n105 585
R463 B.n554 B.n553 585
R464 B.n555 B.n104 585
R465 B.n557 B.n556 585
R466 B.n558 B.n103 585
R467 B.n560 B.n559 585
R468 B.n561 B.n102 585
R469 B.n563 B.n562 585
R470 B.n564 B.n101 585
R471 B.n566 B.n565 585
R472 B.n567 B.n100 585
R473 B.n569 B.n568 585
R474 B.n570 B.n99 585
R475 B.n572 B.n571 585
R476 B.n573 B.n98 585
R477 B.n575 B.n574 585
R478 B.n576 B.n97 585
R479 B.n578 B.n577 585
R480 B.n579 B.n96 585
R481 B.n581 B.n580 585
R482 B.n582 B.n95 585
R483 B.n584 B.n583 585
R484 B.n585 B.n94 585
R485 B.n587 B.n586 585
R486 B.n588 B.n93 585
R487 B.n590 B.n589 585
R488 B.n591 B.n92 585
R489 B.n593 B.n592 585
R490 B.n594 B.n91 585
R491 B.n596 B.n595 585
R492 B.n597 B.n90 585
R493 B.n599 B.n598 585
R494 B.n600 B.n89 585
R495 B.n602 B.n601 585
R496 B.n603 B.n88 585
R497 B.n605 B.n604 585
R498 B.n606 B.n87 585
R499 B.n608 B.n607 585
R500 B.n609 B.n86 585
R501 B.n611 B.n610 585
R502 B.n612 B.n85 585
R503 B.n614 B.n613 585
R504 B.n615 B.n84 585
R505 B.n617 B.n616 585
R506 B.n618 B.n83 585
R507 B.n620 B.n619 585
R508 B.n621 B.n82 585
R509 B.n623 B.n622 585
R510 B.n624 B.n81 585
R511 B.n626 B.n625 585
R512 B.n627 B.n80 585
R513 B.n754 B.n33 585
R514 B.n753 B.n752 585
R515 B.n751 B.n34 585
R516 B.n750 B.n749 585
R517 B.n748 B.n35 585
R518 B.n747 B.n746 585
R519 B.n745 B.n36 585
R520 B.n744 B.n743 585
R521 B.n742 B.n37 585
R522 B.n741 B.n740 585
R523 B.n739 B.n38 585
R524 B.n738 B.n737 585
R525 B.n736 B.n39 585
R526 B.n735 B.n734 585
R527 B.n733 B.n40 585
R528 B.n732 B.n731 585
R529 B.n730 B.n41 585
R530 B.n729 B.n728 585
R531 B.n727 B.n42 585
R532 B.n726 B.n725 585
R533 B.n724 B.n43 585
R534 B.n723 B.n722 585
R535 B.n721 B.n44 585
R536 B.n720 B.n719 585
R537 B.n718 B.n45 585
R538 B.n717 B.n716 585
R539 B.n715 B.n46 585
R540 B.n714 B.n713 585
R541 B.n712 B.n47 585
R542 B.n711 B.n710 585
R543 B.n709 B.n48 585
R544 B.n708 B.n707 585
R545 B.n706 B.n49 585
R546 B.n705 B.n704 585
R547 B.n703 B.n50 585
R548 B.n702 B.n701 585
R549 B.n700 B.n51 585
R550 B.n698 B.n697 585
R551 B.n696 B.n54 585
R552 B.n695 B.n694 585
R553 B.n693 B.n55 585
R554 B.n692 B.n691 585
R555 B.n690 B.n56 585
R556 B.n689 B.n688 585
R557 B.n687 B.n57 585
R558 B.n686 B.n685 585
R559 B.n684 B.n58 585
R560 B.n683 B.n682 585
R561 B.n681 B.n59 585
R562 B.n680 B.n679 585
R563 B.n678 B.n63 585
R564 B.n677 B.n676 585
R565 B.n675 B.n64 585
R566 B.n674 B.n673 585
R567 B.n672 B.n65 585
R568 B.n671 B.n670 585
R569 B.n669 B.n66 585
R570 B.n668 B.n667 585
R571 B.n666 B.n67 585
R572 B.n665 B.n664 585
R573 B.n663 B.n68 585
R574 B.n662 B.n661 585
R575 B.n660 B.n69 585
R576 B.n659 B.n658 585
R577 B.n657 B.n70 585
R578 B.n656 B.n655 585
R579 B.n654 B.n71 585
R580 B.n653 B.n652 585
R581 B.n651 B.n72 585
R582 B.n650 B.n649 585
R583 B.n648 B.n73 585
R584 B.n647 B.n646 585
R585 B.n645 B.n74 585
R586 B.n644 B.n643 585
R587 B.n642 B.n75 585
R588 B.n641 B.n640 585
R589 B.n639 B.n76 585
R590 B.n638 B.n637 585
R591 B.n636 B.n77 585
R592 B.n635 B.n634 585
R593 B.n633 B.n78 585
R594 B.n632 B.n631 585
R595 B.n630 B.n79 585
R596 B.n629 B.n628 585
R597 B.n756 B.n755 585
R598 B.n757 B.n32 585
R599 B.n759 B.n758 585
R600 B.n760 B.n31 585
R601 B.n762 B.n761 585
R602 B.n763 B.n30 585
R603 B.n765 B.n764 585
R604 B.n766 B.n29 585
R605 B.n768 B.n767 585
R606 B.n769 B.n28 585
R607 B.n771 B.n770 585
R608 B.n772 B.n27 585
R609 B.n774 B.n773 585
R610 B.n775 B.n26 585
R611 B.n777 B.n776 585
R612 B.n778 B.n25 585
R613 B.n780 B.n779 585
R614 B.n781 B.n24 585
R615 B.n783 B.n782 585
R616 B.n784 B.n23 585
R617 B.n786 B.n785 585
R618 B.n787 B.n22 585
R619 B.n789 B.n788 585
R620 B.n790 B.n21 585
R621 B.n792 B.n791 585
R622 B.n793 B.n20 585
R623 B.n795 B.n794 585
R624 B.n796 B.n19 585
R625 B.n798 B.n797 585
R626 B.n799 B.n18 585
R627 B.n801 B.n800 585
R628 B.n802 B.n17 585
R629 B.n804 B.n803 585
R630 B.n805 B.n16 585
R631 B.n807 B.n806 585
R632 B.n808 B.n15 585
R633 B.n810 B.n809 585
R634 B.n811 B.n14 585
R635 B.n813 B.n812 585
R636 B.n814 B.n13 585
R637 B.n816 B.n815 585
R638 B.n817 B.n12 585
R639 B.n819 B.n818 585
R640 B.n820 B.n11 585
R641 B.n822 B.n821 585
R642 B.n823 B.n10 585
R643 B.n825 B.n824 585
R644 B.n826 B.n9 585
R645 B.n828 B.n827 585
R646 B.n829 B.n8 585
R647 B.n831 B.n830 585
R648 B.n832 B.n7 585
R649 B.n834 B.n833 585
R650 B.n835 B.n6 585
R651 B.n837 B.n836 585
R652 B.n838 B.n5 585
R653 B.n840 B.n839 585
R654 B.n841 B.n4 585
R655 B.n843 B.n842 585
R656 B.n844 B.n3 585
R657 B.n846 B.n845 585
R658 B.n847 B.n0 585
R659 B.n2 B.n1 585
R660 B.n218 B.n217 585
R661 B.n220 B.n219 585
R662 B.n221 B.n216 585
R663 B.n223 B.n222 585
R664 B.n224 B.n215 585
R665 B.n226 B.n225 585
R666 B.n227 B.n214 585
R667 B.n229 B.n228 585
R668 B.n230 B.n213 585
R669 B.n232 B.n231 585
R670 B.n233 B.n212 585
R671 B.n235 B.n234 585
R672 B.n236 B.n211 585
R673 B.n238 B.n237 585
R674 B.n239 B.n210 585
R675 B.n241 B.n240 585
R676 B.n242 B.n209 585
R677 B.n244 B.n243 585
R678 B.n245 B.n208 585
R679 B.n247 B.n246 585
R680 B.n248 B.n207 585
R681 B.n250 B.n249 585
R682 B.n251 B.n206 585
R683 B.n253 B.n252 585
R684 B.n254 B.n205 585
R685 B.n256 B.n255 585
R686 B.n257 B.n204 585
R687 B.n259 B.n258 585
R688 B.n260 B.n203 585
R689 B.n262 B.n261 585
R690 B.n263 B.n202 585
R691 B.n265 B.n264 585
R692 B.n266 B.n201 585
R693 B.n268 B.n267 585
R694 B.n269 B.n200 585
R695 B.n271 B.n270 585
R696 B.n272 B.n199 585
R697 B.n274 B.n273 585
R698 B.n275 B.n198 585
R699 B.n277 B.n276 585
R700 B.n278 B.n197 585
R701 B.n280 B.n279 585
R702 B.n281 B.n196 585
R703 B.n283 B.n282 585
R704 B.n284 B.n195 585
R705 B.n286 B.n285 585
R706 B.n287 B.n194 585
R707 B.n289 B.n288 585
R708 B.n290 B.n193 585
R709 B.n292 B.n291 585
R710 B.n293 B.n192 585
R711 B.n295 B.n294 585
R712 B.n296 B.n191 585
R713 B.n298 B.n297 585
R714 B.n299 B.n190 585
R715 B.n301 B.n300 585
R716 B.n302 B.n189 585
R717 B.n304 B.n303 585
R718 B.n305 B.n188 585
R719 B.n307 B.n306 585
R720 B.n308 B.n187 585
R721 B.n309 B.n308 468.476
R722 B.n439 B.n438 468.476
R723 B.n629 B.n80 468.476
R724 B.n756 B.n33 468.476
R725 B.n167 B.t3 283.562
R726 B.n379 B.t6 283.562
R727 B.n60 B.t9 283.562
R728 B.n52 B.t0 283.562
R729 B.n849 B.n848 256.663
R730 B.n848 B.n847 235.042
R731 B.n848 B.n2 235.042
R732 B.n379 B.t7 183.751
R733 B.n60 B.t11 183.751
R734 B.n167 B.t4 183.738
R735 B.n52 B.t2 183.738
R736 B.n309 B.n186 163.367
R737 B.n313 B.n186 163.367
R738 B.n314 B.n313 163.367
R739 B.n315 B.n314 163.367
R740 B.n315 B.n184 163.367
R741 B.n319 B.n184 163.367
R742 B.n320 B.n319 163.367
R743 B.n321 B.n320 163.367
R744 B.n321 B.n182 163.367
R745 B.n325 B.n182 163.367
R746 B.n326 B.n325 163.367
R747 B.n327 B.n326 163.367
R748 B.n327 B.n180 163.367
R749 B.n331 B.n180 163.367
R750 B.n332 B.n331 163.367
R751 B.n333 B.n332 163.367
R752 B.n333 B.n178 163.367
R753 B.n337 B.n178 163.367
R754 B.n338 B.n337 163.367
R755 B.n339 B.n338 163.367
R756 B.n339 B.n176 163.367
R757 B.n343 B.n176 163.367
R758 B.n344 B.n343 163.367
R759 B.n345 B.n344 163.367
R760 B.n345 B.n174 163.367
R761 B.n349 B.n174 163.367
R762 B.n350 B.n349 163.367
R763 B.n351 B.n350 163.367
R764 B.n351 B.n172 163.367
R765 B.n355 B.n172 163.367
R766 B.n356 B.n355 163.367
R767 B.n357 B.n356 163.367
R768 B.n357 B.n170 163.367
R769 B.n361 B.n170 163.367
R770 B.n362 B.n361 163.367
R771 B.n363 B.n362 163.367
R772 B.n363 B.n166 163.367
R773 B.n368 B.n166 163.367
R774 B.n369 B.n368 163.367
R775 B.n370 B.n369 163.367
R776 B.n370 B.n164 163.367
R777 B.n374 B.n164 163.367
R778 B.n375 B.n374 163.367
R779 B.n376 B.n375 163.367
R780 B.n376 B.n162 163.367
R781 B.n383 B.n162 163.367
R782 B.n384 B.n383 163.367
R783 B.n385 B.n384 163.367
R784 B.n385 B.n160 163.367
R785 B.n389 B.n160 163.367
R786 B.n390 B.n389 163.367
R787 B.n391 B.n390 163.367
R788 B.n391 B.n158 163.367
R789 B.n395 B.n158 163.367
R790 B.n396 B.n395 163.367
R791 B.n397 B.n396 163.367
R792 B.n397 B.n156 163.367
R793 B.n401 B.n156 163.367
R794 B.n402 B.n401 163.367
R795 B.n403 B.n402 163.367
R796 B.n403 B.n154 163.367
R797 B.n407 B.n154 163.367
R798 B.n408 B.n407 163.367
R799 B.n409 B.n408 163.367
R800 B.n409 B.n152 163.367
R801 B.n413 B.n152 163.367
R802 B.n414 B.n413 163.367
R803 B.n415 B.n414 163.367
R804 B.n415 B.n150 163.367
R805 B.n419 B.n150 163.367
R806 B.n420 B.n419 163.367
R807 B.n421 B.n420 163.367
R808 B.n421 B.n148 163.367
R809 B.n425 B.n148 163.367
R810 B.n426 B.n425 163.367
R811 B.n427 B.n426 163.367
R812 B.n427 B.n146 163.367
R813 B.n431 B.n146 163.367
R814 B.n432 B.n431 163.367
R815 B.n433 B.n432 163.367
R816 B.n433 B.n144 163.367
R817 B.n437 B.n144 163.367
R818 B.n438 B.n437 163.367
R819 B.n625 B.n80 163.367
R820 B.n625 B.n624 163.367
R821 B.n624 B.n623 163.367
R822 B.n623 B.n82 163.367
R823 B.n619 B.n82 163.367
R824 B.n619 B.n618 163.367
R825 B.n618 B.n617 163.367
R826 B.n617 B.n84 163.367
R827 B.n613 B.n84 163.367
R828 B.n613 B.n612 163.367
R829 B.n612 B.n611 163.367
R830 B.n611 B.n86 163.367
R831 B.n607 B.n86 163.367
R832 B.n607 B.n606 163.367
R833 B.n606 B.n605 163.367
R834 B.n605 B.n88 163.367
R835 B.n601 B.n88 163.367
R836 B.n601 B.n600 163.367
R837 B.n600 B.n599 163.367
R838 B.n599 B.n90 163.367
R839 B.n595 B.n90 163.367
R840 B.n595 B.n594 163.367
R841 B.n594 B.n593 163.367
R842 B.n593 B.n92 163.367
R843 B.n589 B.n92 163.367
R844 B.n589 B.n588 163.367
R845 B.n588 B.n587 163.367
R846 B.n587 B.n94 163.367
R847 B.n583 B.n94 163.367
R848 B.n583 B.n582 163.367
R849 B.n582 B.n581 163.367
R850 B.n581 B.n96 163.367
R851 B.n577 B.n96 163.367
R852 B.n577 B.n576 163.367
R853 B.n576 B.n575 163.367
R854 B.n575 B.n98 163.367
R855 B.n571 B.n98 163.367
R856 B.n571 B.n570 163.367
R857 B.n570 B.n569 163.367
R858 B.n569 B.n100 163.367
R859 B.n565 B.n100 163.367
R860 B.n565 B.n564 163.367
R861 B.n564 B.n563 163.367
R862 B.n563 B.n102 163.367
R863 B.n559 B.n102 163.367
R864 B.n559 B.n558 163.367
R865 B.n558 B.n557 163.367
R866 B.n557 B.n104 163.367
R867 B.n553 B.n104 163.367
R868 B.n553 B.n552 163.367
R869 B.n552 B.n551 163.367
R870 B.n551 B.n106 163.367
R871 B.n547 B.n106 163.367
R872 B.n547 B.n546 163.367
R873 B.n546 B.n545 163.367
R874 B.n545 B.n108 163.367
R875 B.n541 B.n108 163.367
R876 B.n541 B.n540 163.367
R877 B.n540 B.n539 163.367
R878 B.n539 B.n110 163.367
R879 B.n535 B.n110 163.367
R880 B.n535 B.n534 163.367
R881 B.n534 B.n533 163.367
R882 B.n533 B.n112 163.367
R883 B.n529 B.n112 163.367
R884 B.n529 B.n528 163.367
R885 B.n528 B.n527 163.367
R886 B.n527 B.n114 163.367
R887 B.n523 B.n114 163.367
R888 B.n523 B.n522 163.367
R889 B.n522 B.n521 163.367
R890 B.n521 B.n116 163.367
R891 B.n517 B.n116 163.367
R892 B.n517 B.n516 163.367
R893 B.n516 B.n515 163.367
R894 B.n515 B.n118 163.367
R895 B.n511 B.n118 163.367
R896 B.n511 B.n510 163.367
R897 B.n510 B.n509 163.367
R898 B.n509 B.n120 163.367
R899 B.n505 B.n120 163.367
R900 B.n505 B.n504 163.367
R901 B.n504 B.n503 163.367
R902 B.n503 B.n122 163.367
R903 B.n499 B.n122 163.367
R904 B.n499 B.n498 163.367
R905 B.n498 B.n497 163.367
R906 B.n497 B.n124 163.367
R907 B.n493 B.n124 163.367
R908 B.n493 B.n492 163.367
R909 B.n492 B.n491 163.367
R910 B.n491 B.n126 163.367
R911 B.n487 B.n126 163.367
R912 B.n487 B.n486 163.367
R913 B.n486 B.n485 163.367
R914 B.n485 B.n128 163.367
R915 B.n481 B.n128 163.367
R916 B.n481 B.n480 163.367
R917 B.n480 B.n479 163.367
R918 B.n479 B.n130 163.367
R919 B.n475 B.n130 163.367
R920 B.n475 B.n474 163.367
R921 B.n474 B.n473 163.367
R922 B.n473 B.n132 163.367
R923 B.n469 B.n132 163.367
R924 B.n469 B.n468 163.367
R925 B.n468 B.n467 163.367
R926 B.n467 B.n134 163.367
R927 B.n463 B.n134 163.367
R928 B.n463 B.n462 163.367
R929 B.n462 B.n461 163.367
R930 B.n461 B.n136 163.367
R931 B.n457 B.n136 163.367
R932 B.n457 B.n456 163.367
R933 B.n456 B.n455 163.367
R934 B.n455 B.n138 163.367
R935 B.n451 B.n138 163.367
R936 B.n451 B.n450 163.367
R937 B.n450 B.n449 163.367
R938 B.n449 B.n140 163.367
R939 B.n445 B.n140 163.367
R940 B.n445 B.n444 163.367
R941 B.n444 B.n443 163.367
R942 B.n443 B.n142 163.367
R943 B.n439 B.n142 163.367
R944 B.n752 B.n33 163.367
R945 B.n752 B.n751 163.367
R946 B.n751 B.n750 163.367
R947 B.n750 B.n35 163.367
R948 B.n746 B.n35 163.367
R949 B.n746 B.n745 163.367
R950 B.n745 B.n744 163.367
R951 B.n744 B.n37 163.367
R952 B.n740 B.n37 163.367
R953 B.n740 B.n739 163.367
R954 B.n739 B.n738 163.367
R955 B.n738 B.n39 163.367
R956 B.n734 B.n39 163.367
R957 B.n734 B.n733 163.367
R958 B.n733 B.n732 163.367
R959 B.n732 B.n41 163.367
R960 B.n728 B.n41 163.367
R961 B.n728 B.n727 163.367
R962 B.n727 B.n726 163.367
R963 B.n726 B.n43 163.367
R964 B.n722 B.n43 163.367
R965 B.n722 B.n721 163.367
R966 B.n721 B.n720 163.367
R967 B.n720 B.n45 163.367
R968 B.n716 B.n45 163.367
R969 B.n716 B.n715 163.367
R970 B.n715 B.n714 163.367
R971 B.n714 B.n47 163.367
R972 B.n710 B.n47 163.367
R973 B.n710 B.n709 163.367
R974 B.n709 B.n708 163.367
R975 B.n708 B.n49 163.367
R976 B.n704 B.n49 163.367
R977 B.n704 B.n703 163.367
R978 B.n703 B.n702 163.367
R979 B.n702 B.n51 163.367
R980 B.n697 B.n51 163.367
R981 B.n697 B.n696 163.367
R982 B.n696 B.n695 163.367
R983 B.n695 B.n55 163.367
R984 B.n691 B.n55 163.367
R985 B.n691 B.n690 163.367
R986 B.n690 B.n689 163.367
R987 B.n689 B.n57 163.367
R988 B.n685 B.n57 163.367
R989 B.n685 B.n684 163.367
R990 B.n684 B.n683 163.367
R991 B.n683 B.n59 163.367
R992 B.n679 B.n59 163.367
R993 B.n679 B.n678 163.367
R994 B.n678 B.n677 163.367
R995 B.n677 B.n64 163.367
R996 B.n673 B.n64 163.367
R997 B.n673 B.n672 163.367
R998 B.n672 B.n671 163.367
R999 B.n671 B.n66 163.367
R1000 B.n667 B.n66 163.367
R1001 B.n667 B.n666 163.367
R1002 B.n666 B.n665 163.367
R1003 B.n665 B.n68 163.367
R1004 B.n661 B.n68 163.367
R1005 B.n661 B.n660 163.367
R1006 B.n660 B.n659 163.367
R1007 B.n659 B.n70 163.367
R1008 B.n655 B.n70 163.367
R1009 B.n655 B.n654 163.367
R1010 B.n654 B.n653 163.367
R1011 B.n653 B.n72 163.367
R1012 B.n649 B.n72 163.367
R1013 B.n649 B.n648 163.367
R1014 B.n648 B.n647 163.367
R1015 B.n647 B.n74 163.367
R1016 B.n643 B.n74 163.367
R1017 B.n643 B.n642 163.367
R1018 B.n642 B.n641 163.367
R1019 B.n641 B.n76 163.367
R1020 B.n637 B.n76 163.367
R1021 B.n637 B.n636 163.367
R1022 B.n636 B.n635 163.367
R1023 B.n635 B.n78 163.367
R1024 B.n631 B.n78 163.367
R1025 B.n631 B.n630 163.367
R1026 B.n630 B.n629 163.367
R1027 B.n757 B.n756 163.367
R1028 B.n758 B.n757 163.367
R1029 B.n758 B.n31 163.367
R1030 B.n762 B.n31 163.367
R1031 B.n763 B.n762 163.367
R1032 B.n764 B.n763 163.367
R1033 B.n764 B.n29 163.367
R1034 B.n768 B.n29 163.367
R1035 B.n769 B.n768 163.367
R1036 B.n770 B.n769 163.367
R1037 B.n770 B.n27 163.367
R1038 B.n774 B.n27 163.367
R1039 B.n775 B.n774 163.367
R1040 B.n776 B.n775 163.367
R1041 B.n776 B.n25 163.367
R1042 B.n780 B.n25 163.367
R1043 B.n781 B.n780 163.367
R1044 B.n782 B.n781 163.367
R1045 B.n782 B.n23 163.367
R1046 B.n786 B.n23 163.367
R1047 B.n787 B.n786 163.367
R1048 B.n788 B.n787 163.367
R1049 B.n788 B.n21 163.367
R1050 B.n792 B.n21 163.367
R1051 B.n793 B.n792 163.367
R1052 B.n794 B.n793 163.367
R1053 B.n794 B.n19 163.367
R1054 B.n798 B.n19 163.367
R1055 B.n799 B.n798 163.367
R1056 B.n800 B.n799 163.367
R1057 B.n800 B.n17 163.367
R1058 B.n804 B.n17 163.367
R1059 B.n805 B.n804 163.367
R1060 B.n806 B.n805 163.367
R1061 B.n806 B.n15 163.367
R1062 B.n810 B.n15 163.367
R1063 B.n811 B.n810 163.367
R1064 B.n812 B.n811 163.367
R1065 B.n812 B.n13 163.367
R1066 B.n816 B.n13 163.367
R1067 B.n817 B.n816 163.367
R1068 B.n818 B.n817 163.367
R1069 B.n818 B.n11 163.367
R1070 B.n822 B.n11 163.367
R1071 B.n823 B.n822 163.367
R1072 B.n824 B.n823 163.367
R1073 B.n824 B.n9 163.367
R1074 B.n828 B.n9 163.367
R1075 B.n829 B.n828 163.367
R1076 B.n830 B.n829 163.367
R1077 B.n830 B.n7 163.367
R1078 B.n834 B.n7 163.367
R1079 B.n835 B.n834 163.367
R1080 B.n836 B.n835 163.367
R1081 B.n836 B.n5 163.367
R1082 B.n840 B.n5 163.367
R1083 B.n841 B.n840 163.367
R1084 B.n842 B.n841 163.367
R1085 B.n842 B.n3 163.367
R1086 B.n846 B.n3 163.367
R1087 B.n847 B.n846 163.367
R1088 B.n218 B.n2 163.367
R1089 B.n219 B.n218 163.367
R1090 B.n219 B.n216 163.367
R1091 B.n223 B.n216 163.367
R1092 B.n224 B.n223 163.367
R1093 B.n225 B.n224 163.367
R1094 B.n225 B.n214 163.367
R1095 B.n229 B.n214 163.367
R1096 B.n230 B.n229 163.367
R1097 B.n231 B.n230 163.367
R1098 B.n231 B.n212 163.367
R1099 B.n235 B.n212 163.367
R1100 B.n236 B.n235 163.367
R1101 B.n237 B.n236 163.367
R1102 B.n237 B.n210 163.367
R1103 B.n241 B.n210 163.367
R1104 B.n242 B.n241 163.367
R1105 B.n243 B.n242 163.367
R1106 B.n243 B.n208 163.367
R1107 B.n247 B.n208 163.367
R1108 B.n248 B.n247 163.367
R1109 B.n249 B.n248 163.367
R1110 B.n249 B.n206 163.367
R1111 B.n253 B.n206 163.367
R1112 B.n254 B.n253 163.367
R1113 B.n255 B.n254 163.367
R1114 B.n255 B.n204 163.367
R1115 B.n259 B.n204 163.367
R1116 B.n260 B.n259 163.367
R1117 B.n261 B.n260 163.367
R1118 B.n261 B.n202 163.367
R1119 B.n265 B.n202 163.367
R1120 B.n266 B.n265 163.367
R1121 B.n267 B.n266 163.367
R1122 B.n267 B.n200 163.367
R1123 B.n271 B.n200 163.367
R1124 B.n272 B.n271 163.367
R1125 B.n273 B.n272 163.367
R1126 B.n273 B.n198 163.367
R1127 B.n277 B.n198 163.367
R1128 B.n278 B.n277 163.367
R1129 B.n279 B.n278 163.367
R1130 B.n279 B.n196 163.367
R1131 B.n283 B.n196 163.367
R1132 B.n284 B.n283 163.367
R1133 B.n285 B.n284 163.367
R1134 B.n285 B.n194 163.367
R1135 B.n289 B.n194 163.367
R1136 B.n290 B.n289 163.367
R1137 B.n291 B.n290 163.367
R1138 B.n291 B.n192 163.367
R1139 B.n295 B.n192 163.367
R1140 B.n296 B.n295 163.367
R1141 B.n297 B.n296 163.367
R1142 B.n297 B.n190 163.367
R1143 B.n301 B.n190 163.367
R1144 B.n302 B.n301 163.367
R1145 B.n303 B.n302 163.367
R1146 B.n303 B.n188 163.367
R1147 B.n307 B.n188 163.367
R1148 B.n308 B.n307 163.367
R1149 B.n380 B.t8 111.993
R1150 B.n61 B.t10 111.993
R1151 B.n168 B.t5 111.981
R1152 B.n53 B.t1 111.981
R1153 B.n168 B.n167 71.7581
R1154 B.n380 B.n379 71.7581
R1155 B.n61 B.n60 71.7581
R1156 B.n53 B.n52 71.7581
R1157 B.n365 B.n168 59.5399
R1158 B.n381 B.n380 59.5399
R1159 B.n62 B.n61 59.5399
R1160 B.n699 B.n53 59.5399
R1161 B.n440 B.n143 30.4395
R1162 B.n755 B.n754 30.4395
R1163 B.n628 B.n627 30.4395
R1164 B.n310 B.n187 30.4395
R1165 B B.n849 18.0485
R1166 B.n755 B.n32 10.6151
R1167 B.n759 B.n32 10.6151
R1168 B.n760 B.n759 10.6151
R1169 B.n761 B.n760 10.6151
R1170 B.n761 B.n30 10.6151
R1171 B.n765 B.n30 10.6151
R1172 B.n766 B.n765 10.6151
R1173 B.n767 B.n766 10.6151
R1174 B.n767 B.n28 10.6151
R1175 B.n771 B.n28 10.6151
R1176 B.n772 B.n771 10.6151
R1177 B.n773 B.n772 10.6151
R1178 B.n773 B.n26 10.6151
R1179 B.n777 B.n26 10.6151
R1180 B.n778 B.n777 10.6151
R1181 B.n779 B.n778 10.6151
R1182 B.n779 B.n24 10.6151
R1183 B.n783 B.n24 10.6151
R1184 B.n784 B.n783 10.6151
R1185 B.n785 B.n784 10.6151
R1186 B.n785 B.n22 10.6151
R1187 B.n789 B.n22 10.6151
R1188 B.n790 B.n789 10.6151
R1189 B.n791 B.n790 10.6151
R1190 B.n791 B.n20 10.6151
R1191 B.n795 B.n20 10.6151
R1192 B.n796 B.n795 10.6151
R1193 B.n797 B.n796 10.6151
R1194 B.n797 B.n18 10.6151
R1195 B.n801 B.n18 10.6151
R1196 B.n802 B.n801 10.6151
R1197 B.n803 B.n802 10.6151
R1198 B.n803 B.n16 10.6151
R1199 B.n807 B.n16 10.6151
R1200 B.n808 B.n807 10.6151
R1201 B.n809 B.n808 10.6151
R1202 B.n809 B.n14 10.6151
R1203 B.n813 B.n14 10.6151
R1204 B.n814 B.n813 10.6151
R1205 B.n815 B.n814 10.6151
R1206 B.n815 B.n12 10.6151
R1207 B.n819 B.n12 10.6151
R1208 B.n820 B.n819 10.6151
R1209 B.n821 B.n820 10.6151
R1210 B.n821 B.n10 10.6151
R1211 B.n825 B.n10 10.6151
R1212 B.n826 B.n825 10.6151
R1213 B.n827 B.n826 10.6151
R1214 B.n827 B.n8 10.6151
R1215 B.n831 B.n8 10.6151
R1216 B.n832 B.n831 10.6151
R1217 B.n833 B.n832 10.6151
R1218 B.n833 B.n6 10.6151
R1219 B.n837 B.n6 10.6151
R1220 B.n838 B.n837 10.6151
R1221 B.n839 B.n838 10.6151
R1222 B.n839 B.n4 10.6151
R1223 B.n843 B.n4 10.6151
R1224 B.n844 B.n843 10.6151
R1225 B.n845 B.n844 10.6151
R1226 B.n845 B.n0 10.6151
R1227 B.n754 B.n753 10.6151
R1228 B.n753 B.n34 10.6151
R1229 B.n749 B.n34 10.6151
R1230 B.n749 B.n748 10.6151
R1231 B.n748 B.n747 10.6151
R1232 B.n747 B.n36 10.6151
R1233 B.n743 B.n36 10.6151
R1234 B.n743 B.n742 10.6151
R1235 B.n742 B.n741 10.6151
R1236 B.n741 B.n38 10.6151
R1237 B.n737 B.n38 10.6151
R1238 B.n737 B.n736 10.6151
R1239 B.n736 B.n735 10.6151
R1240 B.n735 B.n40 10.6151
R1241 B.n731 B.n40 10.6151
R1242 B.n731 B.n730 10.6151
R1243 B.n730 B.n729 10.6151
R1244 B.n729 B.n42 10.6151
R1245 B.n725 B.n42 10.6151
R1246 B.n725 B.n724 10.6151
R1247 B.n724 B.n723 10.6151
R1248 B.n723 B.n44 10.6151
R1249 B.n719 B.n44 10.6151
R1250 B.n719 B.n718 10.6151
R1251 B.n718 B.n717 10.6151
R1252 B.n717 B.n46 10.6151
R1253 B.n713 B.n46 10.6151
R1254 B.n713 B.n712 10.6151
R1255 B.n712 B.n711 10.6151
R1256 B.n711 B.n48 10.6151
R1257 B.n707 B.n48 10.6151
R1258 B.n707 B.n706 10.6151
R1259 B.n706 B.n705 10.6151
R1260 B.n705 B.n50 10.6151
R1261 B.n701 B.n50 10.6151
R1262 B.n701 B.n700 10.6151
R1263 B.n698 B.n54 10.6151
R1264 B.n694 B.n54 10.6151
R1265 B.n694 B.n693 10.6151
R1266 B.n693 B.n692 10.6151
R1267 B.n692 B.n56 10.6151
R1268 B.n688 B.n56 10.6151
R1269 B.n688 B.n687 10.6151
R1270 B.n687 B.n686 10.6151
R1271 B.n686 B.n58 10.6151
R1272 B.n682 B.n681 10.6151
R1273 B.n681 B.n680 10.6151
R1274 B.n680 B.n63 10.6151
R1275 B.n676 B.n63 10.6151
R1276 B.n676 B.n675 10.6151
R1277 B.n675 B.n674 10.6151
R1278 B.n674 B.n65 10.6151
R1279 B.n670 B.n65 10.6151
R1280 B.n670 B.n669 10.6151
R1281 B.n669 B.n668 10.6151
R1282 B.n668 B.n67 10.6151
R1283 B.n664 B.n67 10.6151
R1284 B.n664 B.n663 10.6151
R1285 B.n663 B.n662 10.6151
R1286 B.n662 B.n69 10.6151
R1287 B.n658 B.n69 10.6151
R1288 B.n658 B.n657 10.6151
R1289 B.n657 B.n656 10.6151
R1290 B.n656 B.n71 10.6151
R1291 B.n652 B.n71 10.6151
R1292 B.n652 B.n651 10.6151
R1293 B.n651 B.n650 10.6151
R1294 B.n650 B.n73 10.6151
R1295 B.n646 B.n73 10.6151
R1296 B.n646 B.n645 10.6151
R1297 B.n645 B.n644 10.6151
R1298 B.n644 B.n75 10.6151
R1299 B.n640 B.n75 10.6151
R1300 B.n640 B.n639 10.6151
R1301 B.n639 B.n638 10.6151
R1302 B.n638 B.n77 10.6151
R1303 B.n634 B.n77 10.6151
R1304 B.n634 B.n633 10.6151
R1305 B.n633 B.n632 10.6151
R1306 B.n632 B.n79 10.6151
R1307 B.n628 B.n79 10.6151
R1308 B.n627 B.n626 10.6151
R1309 B.n626 B.n81 10.6151
R1310 B.n622 B.n81 10.6151
R1311 B.n622 B.n621 10.6151
R1312 B.n621 B.n620 10.6151
R1313 B.n620 B.n83 10.6151
R1314 B.n616 B.n83 10.6151
R1315 B.n616 B.n615 10.6151
R1316 B.n615 B.n614 10.6151
R1317 B.n614 B.n85 10.6151
R1318 B.n610 B.n85 10.6151
R1319 B.n610 B.n609 10.6151
R1320 B.n609 B.n608 10.6151
R1321 B.n608 B.n87 10.6151
R1322 B.n604 B.n87 10.6151
R1323 B.n604 B.n603 10.6151
R1324 B.n603 B.n602 10.6151
R1325 B.n602 B.n89 10.6151
R1326 B.n598 B.n89 10.6151
R1327 B.n598 B.n597 10.6151
R1328 B.n597 B.n596 10.6151
R1329 B.n596 B.n91 10.6151
R1330 B.n592 B.n91 10.6151
R1331 B.n592 B.n591 10.6151
R1332 B.n591 B.n590 10.6151
R1333 B.n590 B.n93 10.6151
R1334 B.n586 B.n93 10.6151
R1335 B.n586 B.n585 10.6151
R1336 B.n585 B.n584 10.6151
R1337 B.n584 B.n95 10.6151
R1338 B.n580 B.n95 10.6151
R1339 B.n580 B.n579 10.6151
R1340 B.n579 B.n578 10.6151
R1341 B.n578 B.n97 10.6151
R1342 B.n574 B.n97 10.6151
R1343 B.n574 B.n573 10.6151
R1344 B.n573 B.n572 10.6151
R1345 B.n572 B.n99 10.6151
R1346 B.n568 B.n99 10.6151
R1347 B.n568 B.n567 10.6151
R1348 B.n567 B.n566 10.6151
R1349 B.n566 B.n101 10.6151
R1350 B.n562 B.n101 10.6151
R1351 B.n562 B.n561 10.6151
R1352 B.n561 B.n560 10.6151
R1353 B.n560 B.n103 10.6151
R1354 B.n556 B.n103 10.6151
R1355 B.n556 B.n555 10.6151
R1356 B.n555 B.n554 10.6151
R1357 B.n554 B.n105 10.6151
R1358 B.n550 B.n105 10.6151
R1359 B.n550 B.n549 10.6151
R1360 B.n549 B.n548 10.6151
R1361 B.n548 B.n107 10.6151
R1362 B.n544 B.n107 10.6151
R1363 B.n544 B.n543 10.6151
R1364 B.n543 B.n542 10.6151
R1365 B.n542 B.n109 10.6151
R1366 B.n538 B.n109 10.6151
R1367 B.n538 B.n537 10.6151
R1368 B.n537 B.n536 10.6151
R1369 B.n536 B.n111 10.6151
R1370 B.n532 B.n111 10.6151
R1371 B.n532 B.n531 10.6151
R1372 B.n531 B.n530 10.6151
R1373 B.n530 B.n113 10.6151
R1374 B.n526 B.n113 10.6151
R1375 B.n526 B.n525 10.6151
R1376 B.n525 B.n524 10.6151
R1377 B.n524 B.n115 10.6151
R1378 B.n520 B.n115 10.6151
R1379 B.n520 B.n519 10.6151
R1380 B.n519 B.n518 10.6151
R1381 B.n518 B.n117 10.6151
R1382 B.n514 B.n117 10.6151
R1383 B.n514 B.n513 10.6151
R1384 B.n513 B.n512 10.6151
R1385 B.n512 B.n119 10.6151
R1386 B.n508 B.n119 10.6151
R1387 B.n508 B.n507 10.6151
R1388 B.n507 B.n506 10.6151
R1389 B.n506 B.n121 10.6151
R1390 B.n502 B.n121 10.6151
R1391 B.n502 B.n501 10.6151
R1392 B.n501 B.n500 10.6151
R1393 B.n500 B.n123 10.6151
R1394 B.n496 B.n123 10.6151
R1395 B.n496 B.n495 10.6151
R1396 B.n495 B.n494 10.6151
R1397 B.n494 B.n125 10.6151
R1398 B.n490 B.n125 10.6151
R1399 B.n490 B.n489 10.6151
R1400 B.n489 B.n488 10.6151
R1401 B.n488 B.n127 10.6151
R1402 B.n484 B.n127 10.6151
R1403 B.n484 B.n483 10.6151
R1404 B.n483 B.n482 10.6151
R1405 B.n482 B.n129 10.6151
R1406 B.n478 B.n129 10.6151
R1407 B.n478 B.n477 10.6151
R1408 B.n477 B.n476 10.6151
R1409 B.n476 B.n131 10.6151
R1410 B.n472 B.n131 10.6151
R1411 B.n472 B.n471 10.6151
R1412 B.n471 B.n470 10.6151
R1413 B.n470 B.n133 10.6151
R1414 B.n466 B.n133 10.6151
R1415 B.n466 B.n465 10.6151
R1416 B.n465 B.n464 10.6151
R1417 B.n464 B.n135 10.6151
R1418 B.n460 B.n135 10.6151
R1419 B.n460 B.n459 10.6151
R1420 B.n459 B.n458 10.6151
R1421 B.n458 B.n137 10.6151
R1422 B.n454 B.n137 10.6151
R1423 B.n454 B.n453 10.6151
R1424 B.n453 B.n452 10.6151
R1425 B.n452 B.n139 10.6151
R1426 B.n448 B.n139 10.6151
R1427 B.n448 B.n447 10.6151
R1428 B.n447 B.n446 10.6151
R1429 B.n446 B.n141 10.6151
R1430 B.n442 B.n141 10.6151
R1431 B.n442 B.n441 10.6151
R1432 B.n441 B.n440 10.6151
R1433 B.n217 B.n1 10.6151
R1434 B.n220 B.n217 10.6151
R1435 B.n221 B.n220 10.6151
R1436 B.n222 B.n221 10.6151
R1437 B.n222 B.n215 10.6151
R1438 B.n226 B.n215 10.6151
R1439 B.n227 B.n226 10.6151
R1440 B.n228 B.n227 10.6151
R1441 B.n228 B.n213 10.6151
R1442 B.n232 B.n213 10.6151
R1443 B.n233 B.n232 10.6151
R1444 B.n234 B.n233 10.6151
R1445 B.n234 B.n211 10.6151
R1446 B.n238 B.n211 10.6151
R1447 B.n239 B.n238 10.6151
R1448 B.n240 B.n239 10.6151
R1449 B.n240 B.n209 10.6151
R1450 B.n244 B.n209 10.6151
R1451 B.n245 B.n244 10.6151
R1452 B.n246 B.n245 10.6151
R1453 B.n246 B.n207 10.6151
R1454 B.n250 B.n207 10.6151
R1455 B.n251 B.n250 10.6151
R1456 B.n252 B.n251 10.6151
R1457 B.n252 B.n205 10.6151
R1458 B.n256 B.n205 10.6151
R1459 B.n257 B.n256 10.6151
R1460 B.n258 B.n257 10.6151
R1461 B.n258 B.n203 10.6151
R1462 B.n262 B.n203 10.6151
R1463 B.n263 B.n262 10.6151
R1464 B.n264 B.n263 10.6151
R1465 B.n264 B.n201 10.6151
R1466 B.n268 B.n201 10.6151
R1467 B.n269 B.n268 10.6151
R1468 B.n270 B.n269 10.6151
R1469 B.n270 B.n199 10.6151
R1470 B.n274 B.n199 10.6151
R1471 B.n275 B.n274 10.6151
R1472 B.n276 B.n275 10.6151
R1473 B.n276 B.n197 10.6151
R1474 B.n280 B.n197 10.6151
R1475 B.n281 B.n280 10.6151
R1476 B.n282 B.n281 10.6151
R1477 B.n282 B.n195 10.6151
R1478 B.n286 B.n195 10.6151
R1479 B.n287 B.n286 10.6151
R1480 B.n288 B.n287 10.6151
R1481 B.n288 B.n193 10.6151
R1482 B.n292 B.n193 10.6151
R1483 B.n293 B.n292 10.6151
R1484 B.n294 B.n293 10.6151
R1485 B.n294 B.n191 10.6151
R1486 B.n298 B.n191 10.6151
R1487 B.n299 B.n298 10.6151
R1488 B.n300 B.n299 10.6151
R1489 B.n300 B.n189 10.6151
R1490 B.n304 B.n189 10.6151
R1491 B.n305 B.n304 10.6151
R1492 B.n306 B.n305 10.6151
R1493 B.n306 B.n187 10.6151
R1494 B.n311 B.n310 10.6151
R1495 B.n312 B.n311 10.6151
R1496 B.n312 B.n185 10.6151
R1497 B.n316 B.n185 10.6151
R1498 B.n317 B.n316 10.6151
R1499 B.n318 B.n317 10.6151
R1500 B.n318 B.n183 10.6151
R1501 B.n322 B.n183 10.6151
R1502 B.n323 B.n322 10.6151
R1503 B.n324 B.n323 10.6151
R1504 B.n324 B.n181 10.6151
R1505 B.n328 B.n181 10.6151
R1506 B.n329 B.n328 10.6151
R1507 B.n330 B.n329 10.6151
R1508 B.n330 B.n179 10.6151
R1509 B.n334 B.n179 10.6151
R1510 B.n335 B.n334 10.6151
R1511 B.n336 B.n335 10.6151
R1512 B.n336 B.n177 10.6151
R1513 B.n340 B.n177 10.6151
R1514 B.n341 B.n340 10.6151
R1515 B.n342 B.n341 10.6151
R1516 B.n342 B.n175 10.6151
R1517 B.n346 B.n175 10.6151
R1518 B.n347 B.n346 10.6151
R1519 B.n348 B.n347 10.6151
R1520 B.n348 B.n173 10.6151
R1521 B.n352 B.n173 10.6151
R1522 B.n353 B.n352 10.6151
R1523 B.n354 B.n353 10.6151
R1524 B.n354 B.n171 10.6151
R1525 B.n358 B.n171 10.6151
R1526 B.n359 B.n358 10.6151
R1527 B.n360 B.n359 10.6151
R1528 B.n360 B.n169 10.6151
R1529 B.n364 B.n169 10.6151
R1530 B.n367 B.n366 10.6151
R1531 B.n367 B.n165 10.6151
R1532 B.n371 B.n165 10.6151
R1533 B.n372 B.n371 10.6151
R1534 B.n373 B.n372 10.6151
R1535 B.n373 B.n163 10.6151
R1536 B.n377 B.n163 10.6151
R1537 B.n378 B.n377 10.6151
R1538 B.n382 B.n378 10.6151
R1539 B.n386 B.n161 10.6151
R1540 B.n387 B.n386 10.6151
R1541 B.n388 B.n387 10.6151
R1542 B.n388 B.n159 10.6151
R1543 B.n392 B.n159 10.6151
R1544 B.n393 B.n392 10.6151
R1545 B.n394 B.n393 10.6151
R1546 B.n394 B.n157 10.6151
R1547 B.n398 B.n157 10.6151
R1548 B.n399 B.n398 10.6151
R1549 B.n400 B.n399 10.6151
R1550 B.n400 B.n155 10.6151
R1551 B.n404 B.n155 10.6151
R1552 B.n405 B.n404 10.6151
R1553 B.n406 B.n405 10.6151
R1554 B.n406 B.n153 10.6151
R1555 B.n410 B.n153 10.6151
R1556 B.n411 B.n410 10.6151
R1557 B.n412 B.n411 10.6151
R1558 B.n412 B.n151 10.6151
R1559 B.n416 B.n151 10.6151
R1560 B.n417 B.n416 10.6151
R1561 B.n418 B.n417 10.6151
R1562 B.n418 B.n149 10.6151
R1563 B.n422 B.n149 10.6151
R1564 B.n423 B.n422 10.6151
R1565 B.n424 B.n423 10.6151
R1566 B.n424 B.n147 10.6151
R1567 B.n428 B.n147 10.6151
R1568 B.n429 B.n428 10.6151
R1569 B.n430 B.n429 10.6151
R1570 B.n430 B.n145 10.6151
R1571 B.n434 B.n145 10.6151
R1572 B.n435 B.n434 10.6151
R1573 B.n436 B.n435 10.6151
R1574 B.n436 B.n143 10.6151
R1575 B.n700 B.n699 9.36635
R1576 B.n682 B.n62 9.36635
R1577 B.n365 B.n364 9.36635
R1578 B.n381 B.n161 9.36635
R1579 B.n849 B.n0 8.11757
R1580 B.n849 B.n1 8.11757
R1581 B.n699 B.n698 1.24928
R1582 B.n62 B.n58 1.24928
R1583 B.n366 B.n365 1.24928
R1584 B.n382 B.n381 1.24928
C0 VTAIL B 4.77381f
C1 VN w_n4670_n3054# 9.689151f
C2 VDD2 VP 0.601315f
C3 VDD1 VN 0.152828f
C4 VN VTAIL 8.69117f
C5 VDD2 w_n4670_n3054# 2.30313f
C6 VDD1 VDD2 2.17389f
C7 VN B 1.38604f
C8 VDD2 VTAIL 7.95858f
C9 VDD2 B 1.96217f
C10 VDD2 VN 7.97254f
C11 VP w_n4670_n3054# 10.297701f
C12 VDD1 VP 8.41924f
C13 VTAIL VP 8.70528f
C14 VDD1 w_n4670_n3054# 2.15612f
C15 VP B 2.41025f
C16 VTAIL w_n4670_n3054# 3.9377f
C17 VDD1 VTAIL 7.899f
C18 B w_n4670_n3054# 10.853901f
C19 VN VP 8.31351f
C20 VDD1 B 1.84192f
C21 VDD2 VSUBS 2.222635f
C22 VDD1 VSUBS 3.00486f
C23 VTAIL VSUBS 1.410293f
C24 VN VSUBS 7.74318f
C25 VP VSUBS 4.326365f
C26 B VSUBS 5.729547f
C27 w_n4670_n3054# VSUBS 0.176022p
C28 B.n0 VSUBS 0.006767f
C29 B.n1 VSUBS 0.006767f
C30 B.n2 VSUBS 0.010008f
C31 B.n3 VSUBS 0.007669f
C32 B.n4 VSUBS 0.007669f
C33 B.n5 VSUBS 0.007669f
C34 B.n6 VSUBS 0.007669f
C35 B.n7 VSUBS 0.007669f
C36 B.n8 VSUBS 0.007669f
C37 B.n9 VSUBS 0.007669f
C38 B.n10 VSUBS 0.007669f
C39 B.n11 VSUBS 0.007669f
C40 B.n12 VSUBS 0.007669f
C41 B.n13 VSUBS 0.007669f
C42 B.n14 VSUBS 0.007669f
C43 B.n15 VSUBS 0.007669f
C44 B.n16 VSUBS 0.007669f
C45 B.n17 VSUBS 0.007669f
C46 B.n18 VSUBS 0.007669f
C47 B.n19 VSUBS 0.007669f
C48 B.n20 VSUBS 0.007669f
C49 B.n21 VSUBS 0.007669f
C50 B.n22 VSUBS 0.007669f
C51 B.n23 VSUBS 0.007669f
C52 B.n24 VSUBS 0.007669f
C53 B.n25 VSUBS 0.007669f
C54 B.n26 VSUBS 0.007669f
C55 B.n27 VSUBS 0.007669f
C56 B.n28 VSUBS 0.007669f
C57 B.n29 VSUBS 0.007669f
C58 B.n30 VSUBS 0.007669f
C59 B.n31 VSUBS 0.007669f
C60 B.n32 VSUBS 0.007669f
C61 B.n33 VSUBS 0.017795f
C62 B.n34 VSUBS 0.007669f
C63 B.n35 VSUBS 0.007669f
C64 B.n36 VSUBS 0.007669f
C65 B.n37 VSUBS 0.007669f
C66 B.n38 VSUBS 0.007669f
C67 B.n39 VSUBS 0.007669f
C68 B.n40 VSUBS 0.007669f
C69 B.n41 VSUBS 0.007669f
C70 B.n42 VSUBS 0.007669f
C71 B.n43 VSUBS 0.007669f
C72 B.n44 VSUBS 0.007669f
C73 B.n45 VSUBS 0.007669f
C74 B.n46 VSUBS 0.007669f
C75 B.n47 VSUBS 0.007669f
C76 B.n48 VSUBS 0.007669f
C77 B.n49 VSUBS 0.007669f
C78 B.n50 VSUBS 0.007669f
C79 B.n51 VSUBS 0.007669f
C80 B.t1 VSUBS 0.366391f
C81 B.t2 VSUBS 0.394151f
C82 B.t0 VSUBS 1.79694f
C83 B.n52 VSUBS 0.219704f
C84 B.n53 VSUBS 0.08202f
C85 B.n54 VSUBS 0.007669f
C86 B.n55 VSUBS 0.007669f
C87 B.n56 VSUBS 0.007669f
C88 B.n57 VSUBS 0.007669f
C89 B.n58 VSUBS 0.004286f
C90 B.n59 VSUBS 0.007669f
C91 B.t10 VSUBS 0.366385f
C92 B.t11 VSUBS 0.394146f
C93 B.t9 VSUBS 1.79694f
C94 B.n60 VSUBS 0.219709f
C95 B.n61 VSUBS 0.082025f
C96 B.n62 VSUBS 0.017769f
C97 B.n63 VSUBS 0.007669f
C98 B.n64 VSUBS 0.007669f
C99 B.n65 VSUBS 0.007669f
C100 B.n66 VSUBS 0.007669f
C101 B.n67 VSUBS 0.007669f
C102 B.n68 VSUBS 0.007669f
C103 B.n69 VSUBS 0.007669f
C104 B.n70 VSUBS 0.007669f
C105 B.n71 VSUBS 0.007669f
C106 B.n72 VSUBS 0.007669f
C107 B.n73 VSUBS 0.007669f
C108 B.n74 VSUBS 0.007669f
C109 B.n75 VSUBS 0.007669f
C110 B.n76 VSUBS 0.007669f
C111 B.n77 VSUBS 0.007669f
C112 B.n78 VSUBS 0.007669f
C113 B.n79 VSUBS 0.007669f
C114 B.n80 VSUBS 0.016491f
C115 B.n81 VSUBS 0.007669f
C116 B.n82 VSUBS 0.007669f
C117 B.n83 VSUBS 0.007669f
C118 B.n84 VSUBS 0.007669f
C119 B.n85 VSUBS 0.007669f
C120 B.n86 VSUBS 0.007669f
C121 B.n87 VSUBS 0.007669f
C122 B.n88 VSUBS 0.007669f
C123 B.n89 VSUBS 0.007669f
C124 B.n90 VSUBS 0.007669f
C125 B.n91 VSUBS 0.007669f
C126 B.n92 VSUBS 0.007669f
C127 B.n93 VSUBS 0.007669f
C128 B.n94 VSUBS 0.007669f
C129 B.n95 VSUBS 0.007669f
C130 B.n96 VSUBS 0.007669f
C131 B.n97 VSUBS 0.007669f
C132 B.n98 VSUBS 0.007669f
C133 B.n99 VSUBS 0.007669f
C134 B.n100 VSUBS 0.007669f
C135 B.n101 VSUBS 0.007669f
C136 B.n102 VSUBS 0.007669f
C137 B.n103 VSUBS 0.007669f
C138 B.n104 VSUBS 0.007669f
C139 B.n105 VSUBS 0.007669f
C140 B.n106 VSUBS 0.007669f
C141 B.n107 VSUBS 0.007669f
C142 B.n108 VSUBS 0.007669f
C143 B.n109 VSUBS 0.007669f
C144 B.n110 VSUBS 0.007669f
C145 B.n111 VSUBS 0.007669f
C146 B.n112 VSUBS 0.007669f
C147 B.n113 VSUBS 0.007669f
C148 B.n114 VSUBS 0.007669f
C149 B.n115 VSUBS 0.007669f
C150 B.n116 VSUBS 0.007669f
C151 B.n117 VSUBS 0.007669f
C152 B.n118 VSUBS 0.007669f
C153 B.n119 VSUBS 0.007669f
C154 B.n120 VSUBS 0.007669f
C155 B.n121 VSUBS 0.007669f
C156 B.n122 VSUBS 0.007669f
C157 B.n123 VSUBS 0.007669f
C158 B.n124 VSUBS 0.007669f
C159 B.n125 VSUBS 0.007669f
C160 B.n126 VSUBS 0.007669f
C161 B.n127 VSUBS 0.007669f
C162 B.n128 VSUBS 0.007669f
C163 B.n129 VSUBS 0.007669f
C164 B.n130 VSUBS 0.007669f
C165 B.n131 VSUBS 0.007669f
C166 B.n132 VSUBS 0.007669f
C167 B.n133 VSUBS 0.007669f
C168 B.n134 VSUBS 0.007669f
C169 B.n135 VSUBS 0.007669f
C170 B.n136 VSUBS 0.007669f
C171 B.n137 VSUBS 0.007669f
C172 B.n138 VSUBS 0.007669f
C173 B.n139 VSUBS 0.007669f
C174 B.n140 VSUBS 0.007669f
C175 B.n141 VSUBS 0.007669f
C176 B.n142 VSUBS 0.007669f
C177 B.n143 VSUBS 0.016823f
C178 B.n144 VSUBS 0.007669f
C179 B.n145 VSUBS 0.007669f
C180 B.n146 VSUBS 0.007669f
C181 B.n147 VSUBS 0.007669f
C182 B.n148 VSUBS 0.007669f
C183 B.n149 VSUBS 0.007669f
C184 B.n150 VSUBS 0.007669f
C185 B.n151 VSUBS 0.007669f
C186 B.n152 VSUBS 0.007669f
C187 B.n153 VSUBS 0.007669f
C188 B.n154 VSUBS 0.007669f
C189 B.n155 VSUBS 0.007669f
C190 B.n156 VSUBS 0.007669f
C191 B.n157 VSUBS 0.007669f
C192 B.n158 VSUBS 0.007669f
C193 B.n159 VSUBS 0.007669f
C194 B.n160 VSUBS 0.007669f
C195 B.n161 VSUBS 0.007218f
C196 B.n162 VSUBS 0.007669f
C197 B.n163 VSUBS 0.007669f
C198 B.n164 VSUBS 0.007669f
C199 B.n165 VSUBS 0.007669f
C200 B.n166 VSUBS 0.007669f
C201 B.t5 VSUBS 0.366391f
C202 B.t4 VSUBS 0.394151f
C203 B.t3 VSUBS 1.79694f
C204 B.n167 VSUBS 0.219704f
C205 B.n168 VSUBS 0.08202f
C206 B.n169 VSUBS 0.007669f
C207 B.n170 VSUBS 0.007669f
C208 B.n171 VSUBS 0.007669f
C209 B.n172 VSUBS 0.007669f
C210 B.n173 VSUBS 0.007669f
C211 B.n174 VSUBS 0.007669f
C212 B.n175 VSUBS 0.007669f
C213 B.n176 VSUBS 0.007669f
C214 B.n177 VSUBS 0.007669f
C215 B.n178 VSUBS 0.007669f
C216 B.n179 VSUBS 0.007669f
C217 B.n180 VSUBS 0.007669f
C218 B.n181 VSUBS 0.007669f
C219 B.n182 VSUBS 0.007669f
C220 B.n183 VSUBS 0.007669f
C221 B.n184 VSUBS 0.007669f
C222 B.n185 VSUBS 0.007669f
C223 B.n186 VSUBS 0.007669f
C224 B.n187 VSUBS 0.016491f
C225 B.n188 VSUBS 0.007669f
C226 B.n189 VSUBS 0.007669f
C227 B.n190 VSUBS 0.007669f
C228 B.n191 VSUBS 0.007669f
C229 B.n192 VSUBS 0.007669f
C230 B.n193 VSUBS 0.007669f
C231 B.n194 VSUBS 0.007669f
C232 B.n195 VSUBS 0.007669f
C233 B.n196 VSUBS 0.007669f
C234 B.n197 VSUBS 0.007669f
C235 B.n198 VSUBS 0.007669f
C236 B.n199 VSUBS 0.007669f
C237 B.n200 VSUBS 0.007669f
C238 B.n201 VSUBS 0.007669f
C239 B.n202 VSUBS 0.007669f
C240 B.n203 VSUBS 0.007669f
C241 B.n204 VSUBS 0.007669f
C242 B.n205 VSUBS 0.007669f
C243 B.n206 VSUBS 0.007669f
C244 B.n207 VSUBS 0.007669f
C245 B.n208 VSUBS 0.007669f
C246 B.n209 VSUBS 0.007669f
C247 B.n210 VSUBS 0.007669f
C248 B.n211 VSUBS 0.007669f
C249 B.n212 VSUBS 0.007669f
C250 B.n213 VSUBS 0.007669f
C251 B.n214 VSUBS 0.007669f
C252 B.n215 VSUBS 0.007669f
C253 B.n216 VSUBS 0.007669f
C254 B.n217 VSUBS 0.007669f
C255 B.n218 VSUBS 0.007669f
C256 B.n219 VSUBS 0.007669f
C257 B.n220 VSUBS 0.007669f
C258 B.n221 VSUBS 0.007669f
C259 B.n222 VSUBS 0.007669f
C260 B.n223 VSUBS 0.007669f
C261 B.n224 VSUBS 0.007669f
C262 B.n225 VSUBS 0.007669f
C263 B.n226 VSUBS 0.007669f
C264 B.n227 VSUBS 0.007669f
C265 B.n228 VSUBS 0.007669f
C266 B.n229 VSUBS 0.007669f
C267 B.n230 VSUBS 0.007669f
C268 B.n231 VSUBS 0.007669f
C269 B.n232 VSUBS 0.007669f
C270 B.n233 VSUBS 0.007669f
C271 B.n234 VSUBS 0.007669f
C272 B.n235 VSUBS 0.007669f
C273 B.n236 VSUBS 0.007669f
C274 B.n237 VSUBS 0.007669f
C275 B.n238 VSUBS 0.007669f
C276 B.n239 VSUBS 0.007669f
C277 B.n240 VSUBS 0.007669f
C278 B.n241 VSUBS 0.007669f
C279 B.n242 VSUBS 0.007669f
C280 B.n243 VSUBS 0.007669f
C281 B.n244 VSUBS 0.007669f
C282 B.n245 VSUBS 0.007669f
C283 B.n246 VSUBS 0.007669f
C284 B.n247 VSUBS 0.007669f
C285 B.n248 VSUBS 0.007669f
C286 B.n249 VSUBS 0.007669f
C287 B.n250 VSUBS 0.007669f
C288 B.n251 VSUBS 0.007669f
C289 B.n252 VSUBS 0.007669f
C290 B.n253 VSUBS 0.007669f
C291 B.n254 VSUBS 0.007669f
C292 B.n255 VSUBS 0.007669f
C293 B.n256 VSUBS 0.007669f
C294 B.n257 VSUBS 0.007669f
C295 B.n258 VSUBS 0.007669f
C296 B.n259 VSUBS 0.007669f
C297 B.n260 VSUBS 0.007669f
C298 B.n261 VSUBS 0.007669f
C299 B.n262 VSUBS 0.007669f
C300 B.n263 VSUBS 0.007669f
C301 B.n264 VSUBS 0.007669f
C302 B.n265 VSUBS 0.007669f
C303 B.n266 VSUBS 0.007669f
C304 B.n267 VSUBS 0.007669f
C305 B.n268 VSUBS 0.007669f
C306 B.n269 VSUBS 0.007669f
C307 B.n270 VSUBS 0.007669f
C308 B.n271 VSUBS 0.007669f
C309 B.n272 VSUBS 0.007669f
C310 B.n273 VSUBS 0.007669f
C311 B.n274 VSUBS 0.007669f
C312 B.n275 VSUBS 0.007669f
C313 B.n276 VSUBS 0.007669f
C314 B.n277 VSUBS 0.007669f
C315 B.n278 VSUBS 0.007669f
C316 B.n279 VSUBS 0.007669f
C317 B.n280 VSUBS 0.007669f
C318 B.n281 VSUBS 0.007669f
C319 B.n282 VSUBS 0.007669f
C320 B.n283 VSUBS 0.007669f
C321 B.n284 VSUBS 0.007669f
C322 B.n285 VSUBS 0.007669f
C323 B.n286 VSUBS 0.007669f
C324 B.n287 VSUBS 0.007669f
C325 B.n288 VSUBS 0.007669f
C326 B.n289 VSUBS 0.007669f
C327 B.n290 VSUBS 0.007669f
C328 B.n291 VSUBS 0.007669f
C329 B.n292 VSUBS 0.007669f
C330 B.n293 VSUBS 0.007669f
C331 B.n294 VSUBS 0.007669f
C332 B.n295 VSUBS 0.007669f
C333 B.n296 VSUBS 0.007669f
C334 B.n297 VSUBS 0.007669f
C335 B.n298 VSUBS 0.007669f
C336 B.n299 VSUBS 0.007669f
C337 B.n300 VSUBS 0.007669f
C338 B.n301 VSUBS 0.007669f
C339 B.n302 VSUBS 0.007669f
C340 B.n303 VSUBS 0.007669f
C341 B.n304 VSUBS 0.007669f
C342 B.n305 VSUBS 0.007669f
C343 B.n306 VSUBS 0.007669f
C344 B.n307 VSUBS 0.007669f
C345 B.n308 VSUBS 0.016491f
C346 B.n309 VSUBS 0.017795f
C347 B.n310 VSUBS 0.017795f
C348 B.n311 VSUBS 0.007669f
C349 B.n312 VSUBS 0.007669f
C350 B.n313 VSUBS 0.007669f
C351 B.n314 VSUBS 0.007669f
C352 B.n315 VSUBS 0.007669f
C353 B.n316 VSUBS 0.007669f
C354 B.n317 VSUBS 0.007669f
C355 B.n318 VSUBS 0.007669f
C356 B.n319 VSUBS 0.007669f
C357 B.n320 VSUBS 0.007669f
C358 B.n321 VSUBS 0.007669f
C359 B.n322 VSUBS 0.007669f
C360 B.n323 VSUBS 0.007669f
C361 B.n324 VSUBS 0.007669f
C362 B.n325 VSUBS 0.007669f
C363 B.n326 VSUBS 0.007669f
C364 B.n327 VSUBS 0.007669f
C365 B.n328 VSUBS 0.007669f
C366 B.n329 VSUBS 0.007669f
C367 B.n330 VSUBS 0.007669f
C368 B.n331 VSUBS 0.007669f
C369 B.n332 VSUBS 0.007669f
C370 B.n333 VSUBS 0.007669f
C371 B.n334 VSUBS 0.007669f
C372 B.n335 VSUBS 0.007669f
C373 B.n336 VSUBS 0.007669f
C374 B.n337 VSUBS 0.007669f
C375 B.n338 VSUBS 0.007669f
C376 B.n339 VSUBS 0.007669f
C377 B.n340 VSUBS 0.007669f
C378 B.n341 VSUBS 0.007669f
C379 B.n342 VSUBS 0.007669f
C380 B.n343 VSUBS 0.007669f
C381 B.n344 VSUBS 0.007669f
C382 B.n345 VSUBS 0.007669f
C383 B.n346 VSUBS 0.007669f
C384 B.n347 VSUBS 0.007669f
C385 B.n348 VSUBS 0.007669f
C386 B.n349 VSUBS 0.007669f
C387 B.n350 VSUBS 0.007669f
C388 B.n351 VSUBS 0.007669f
C389 B.n352 VSUBS 0.007669f
C390 B.n353 VSUBS 0.007669f
C391 B.n354 VSUBS 0.007669f
C392 B.n355 VSUBS 0.007669f
C393 B.n356 VSUBS 0.007669f
C394 B.n357 VSUBS 0.007669f
C395 B.n358 VSUBS 0.007669f
C396 B.n359 VSUBS 0.007669f
C397 B.n360 VSUBS 0.007669f
C398 B.n361 VSUBS 0.007669f
C399 B.n362 VSUBS 0.007669f
C400 B.n363 VSUBS 0.007669f
C401 B.n364 VSUBS 0.007218f
C402 B.n365 VSUBS 0.017769f
C403 B.n366 VSUBS 0.004286f
C404 B.n367 VSUBS 0.007669f
C405 B.n368 VSUBS 0.007669f
C406 B.n369 VSUBS 0.007669f
C407 B.n370 VSUBS 0.007669f
C408 B.n371 VSUBS 0.007669f
C409 B.n372 VSUBS 0.007669f
C410 B.n373 VSUBS 0.007669f
C411 B.n374 VSUBS 0.007669f
C412 B.n375 VSUBS 0.007669f
C413 B.n376 VSUBS 0.007669f
C414 B.n377 VSUBS 0.007669f
C415 B.n378 VSUBS 0.007669f
C416 B.t8 VSUBS 0.366385f
C417 B.t7 VSUBS 0.394146f
C418 B.t6 VSUBS 1.79694f
C419 B.n379 VSUBS 0.219709f
C420 B.n380 VSUBS 0.082025f
C421 B.n381 VSUBS 0.017769f
C422 B.n382 VSUBS 0.004286f
C423 B.n383 VSUBS 0.007669f
C424 B.n384 VSUBS 0.007669f
C425 B.n385 VSUBS 0.007669f
C426 B.n386 VSUBS 0.007669f
C427 B.n387 VSUBS 0.007669f
C428 B.n388 VSUBS 0.007669f
C429 B.n389 VSUBS 0.007669f
C430 B.n390 VSUBS 0.007669f
C431 B.n391 VSUBS 0.007669f
C432 B.n392 VSUBS 0.007669f
C433 B.n393 VSUBS 0.007669f
C434 B.n394 VSUBS 0.007669f
C435 B.n395 VSUBS 0.007669f
C436 B.n396 VSUBS 0.007669f
C437 B.n397 VSUBS 0.007669f
C438 B.n398 VSUBS 0.007669f
C439 B.n399 VSUBS 0.007669f
C440 B.n400 VSUBS 0.007669f
C441 B.n401 VSUBS 0.007669f
C442 B.n402 VSUBS 0.007669f
C443 B.n403 VSUBS 0.007669f
C444 B.n404 VSUBS 0.007669f
C445 B.n405 VSUBS 0.007669f
C446 B.n406 VSUBS 0.007669f
C447 B.n407 VSUBS 0.007669f
C448 B.n408 VSUBS 0.007669f
C449 B.n409 VSUBS 0.007669f
C450 B.n410 VSUBS 0.007669f
C451 B.n411 VSUBS 0.007669f
C452 B.n412 VSUBS 0.007669f
C453 B.n413 VSUBS 0.007669f
C454 B.n414 VSUBS 0.007669f
C455 B.n415 VSUBS 0.007669f
C456 B.n416 VSUBS 0.007669f
C457 B.n417 VSUBS 0.007669f
C458 B.n418 VSUBS 0.007669f
C459 B.n419 VSUBS 0.007669f
C460 B.n420 VSUBS 0.007669f
C461 B.n421 VSUBS 0.007669f
C462 B.n422 VSUBS 0.007669f
C463 B.n423 VSUBS 0.007669f
C464 B.n424 VSUBS 0.007669f
C465 B.n425 VSUBS 0.007669f
C466 B.n426 VSUBS 0.007669f
C467 B.n427 VSUBS 0.007669f
C468 B.n428 VSUBS 0.007669f
C469 B.n429 VSUBS 0.007669f
C470 B.n430 VSUBS 0.007669f
C471 B.n431 VSUBS 0.007669f
C472 B.n432 VSUBS 0.007669f
C473 B.n433 VSUBS 0.007669f
C474 B.n434 VSUBS 0.007669f
C475 B.n435 VSUBS 0.007669f
C476 B.n436 VSUBS 0.007669f
C477 B.n437 VSUBS 0.007669f
C478 B.n438 VSUBS 0.017795f
C479 B.n439 VSUBS 0.016491f
C480 B.n440 VSUBS 0.017463f
C481 B.n441 VSUBS 0.007669f
C482 B.n442 VSUBS 0.007669f
C483 B.n443 VSUBS 0.007669f
C484 B.n444 VSUBS 0.007669f
C485 B.n445 VSUBS 0.007669f
C486 B.n446 VSUBS 0.007669f
C487 B.n447 VSUBS 0.007669f
C488 B.n448 VSUBS 0.007669f
C489 B.n449 VSUBS 0.007669f
C490 B.n450 VSUBS 0.007669f
C491 B.n451 VSUBS 0.007669f
C492 B.n452 VSUBS 0.007669f
C493 B.n453 VSUBS 0.007669f
C494 B.n454 VSUBS 0.007669f
C495 B.n455 VSUBS 0.007669f
C496 B.n456 VSUBS 0.007669f
C497 B.n457 VSUBS 0.007669f
C498 B.n458 VSUBS 0.007669f
C499 B.n459 VSUBS 0.007669f
C500 B.n460 VSUBS 0.007669f
C501 B.n461 VSUBS 0.007669f
C502 B.n462 VSUBS 0.007669f
C503 B.n463 VSUBS 0.007669f
C504 B.n464 VSUBS 0.007669f
C505 B.n465 VSUBS 0.007669f
C506 B.n466 VSUBS 0.007669f
C507 B.n467 VSUBS 0.007669f
C508 B.n468 VSUBS 0.007669f
C509 B.n469 VSUBS 0.007669f
C510 B.n470 VSUBS 0.007669f
C511 B.n471 VSUBS 0.007669f
C512 B.n472 VSUBS 0.007669f
C513 B.n473 VSUBS 0.007669f
C514 B.n474 VSUBS 0.007669f
C515 B.n475 VSUBS 0.007669f
C516 B.n476 VSUBS 0.007669f
C517 B.n477 VSUBS 0.007669f
C518 B.n478 VSUBS 0.007669f
C519 B.n479 VSUBS 0.007669f
C520 B.n480 VSUBS 0.007669f
C521 B.n481 VSUBS 0.007669f
C522 B.n482 VSUBS 0.007669f
C523 B.n483 VSUBS 0.007669f
C524 B.n484 VSUBS 0.007669f
C525 B.n485 VSUBS 0.007669f
C526 B.n486 VSUBS 0.007669f
C527 B.n487 VSUBS 0.007669f
C528 B.n488 VSUBS 0.007669f
C529 B.n489 VSUBS 0.007669f
C530 B.n490 VSUBS 0.007669f
C531 B.n491 VSUBS 0.007669f
C532 B.n492 VSUBS 0.007669f
C533 B.n493 VSUBS 0.007669f
C534 B.n494 VSUBS 0.007669f
C535 B.n495 VSUBS 0.007669f
C536 B.n496 VSUBS 0.007669f
C537 B.n497 VSUBS 0.007669f
C538 B.n498 VSUBS 0.007669f
C539 B.n499 VSUBS 0.007669f
C540 B.n500 VSUBS 0.007669f
C541 B.n501 VSUBS 0.007669f
C542 B.n502 VSUBS 0.007669f
C543 B.n503 VSUBS 0.007669f
C544 B.n504 VSUBS 0.007669f
C545 B.n505 VSUBS 0.007669f
C546 B.n506 VSUBS 0.007669f
C547 B.n507 VSUBS 0.007669f
C548 B.n508 VSUBS 0.007669f
C549 B.n509 VSUBS 0.007669f
C550 B.n510 VSUBS 0.007669f
C551 B.n511 VSUBS 0.007669f
C552 B.n512 VSUBS 0.007669f
C553 B.n513 VSUBS 0.007669f
C554 B.n514 VSUBS 0.007669f
C555 B.n515 VSUBS 0.007669f
C556 B.n516 VSUBS 0.007669f
C557 B.n517 VSUBS 0.007669f
C558 B.n518 VSUBS 0.007669f
C559 B.n519 VSUBS 0.007669f
C560 B.n520 VSUBS 0.007669f
C561 B.n521 VSUBS 0.007669f
C562 B.n522 VSUBS 0.007669f
C563 B.n523 VSUBS 0.007669f
C564 B.n524 VSUBS 0.007669f
C565 B.n525 VSUBS 0.007669f
C566 B.n526 VSUBS 0.007669f
C567 B.n527 VSUBS 0.007669f
C568 B.n528 VSUBS 0.007669f
C569 B.n529 VSUBS 0.007669f
C570 B.n530 VSUBS 0.007669f
C571 B.n531 VSUBS 0.007669f
C572 B.n532 VSUBS 0.007669f
C573 B.n533 VSUBS 0.007669f
C574 B.n534 VSUBS 0.007669f
C575 B.n535 VSUBS 0.007669f
C576 B.n536 VSUBS 0.007669f
C577 B.n537 VSUBS 0.007669f
C578 B.n538 VSUBS 0.007669f
C579 B.n539 VSUBS 0.007669f
C580 B.n540 VSUBS 0.007669f
C581 B.n541 VSUBS 0.007669f
C582 B.n542 VSUBS 0.007669f
C583 B.n543 VSUBS 0.007669f
C584 B.n544 VSUBS 0.007669f
C585 B.n545 VSUBS 0.007669f
C586 B.n546 VSUBS 0.007669f
C587 B.n547 VSUBS 0.007669f
C588 B.n548 VSUBS 0.007669f
C589 B.n549 VSUBS 0.007669f
C590 B.n550 VSUBS 0.007669f
C591 B.n551 VSUBS 0.007669f
C592 B.n552 VSUBS 0.007669f
C593 B.n553 VSUBS 0.007669f
C594 B.n554 VSUBS 0.007669f
C595 B.n555 VSUBS 0.007669f
C596 B.n556 VSUBS 0.007669f
C597 B.n557 VSUBS 0.007669f
C598 B.n558 VSUBS 0.007669f
C599 B.n559 VSUBS 0.007669f
C600 B.n560 VSUBS 0.007669f
C601 B.n561 VSUBS 0.007669f
C602 B.n562 VSUBS 0.007669f
C603 B.n563 VSUBS 0.007669f
C604 B.n564 VSUBS 0.007669f
C605 B.n565 VSUBS 0.007669f
C606 B.n566 VSUBS 0.007669f
C607 B.n567 VSUBS 0.007669f
C608 B.n568 VSUBS 0.007669f
C609 B.n569 VSUBS 0.007669f
C610 B.n570 VSUBS 0.007669f
C611 B.n571 VSUBS 0.007669f
C612 B.n572 VSUBS 0.007669f
C613 B.n573 VSUBS 0.007669f
C614 B.n574 VSUBS 0.007669f
C615 B.n575 VSUBS 0.007669f
C616 B.n576 VSUBS 0.007669f
C617 B.n577 VSUBS 0.007669f
C618 B.n578 VSUBS 0.007669f
C619 B.n579 VSUBS 0.007669f
C620 B.n580 VSUBS 0.007669f
C621 B.n581 VSUBS 0.007669f
C622 B.n582 VSUBS 0.007669f
C623 B.n583 VSUBS 0.007669f
C624 B.n584 VSUBS 0.007669f
C625 B.n585 VSUBS 0.007669f
C626 B.n586 VSUBS 0.007669f
C627 B.n587 VSUBS 0.007669f
C628 B.n588 VSUBS 0.007669f
C629 B.n589 VSUBS 0.007669f
C630 B.n590 VSUBS 0.007669f
C631 B.n591 VSUBS 0.007669f
C632 B.n592 VSUBS 0.007669f
C633 B.n593 VSUBS 0.007669f
C634 B.n594 VSUBS 0.007669f
C635 B.n595 VSUBS 0.007669f
C636 B.n596 VSUBS 0.007669f
C637 B.n597 VSUBS 0.007669f
C638 B.n598 VSUBS 0.007669f
C639 B.n599 VSUBS 0.007669f
C640 B.n600 VSUBS 0.007669f
C641 B.n601 VSUBS 0.007669f
C642 B.n602 VSUBS 0.007669f
C643 B.n603 VSUBS 0.007669f
C644 B.n604 VSUBS 0.007669f
C645 B.n605 VSUBS 0.007669f
C646 B.n606 VSUBS 0.007669f
C647 B.n607 VSUBS 0.007669f
C648 B.n608 VSUBS 0.007669f
C649 B.n609 VSUBS 0.007669f
C650 B.n610 VSUBS 0.007669f
C651 B.n611 VSUBS 0.007669f
C652 B.n612 VSUBS 0.007669f
C653 B.n613 VSUBS 0.007669f
C654 B.n614 VSUBS 0.007669f
C655 B.n615 VSUBS 0.007669f
C656 B.n616 VSUBS 0.007669f
C657 B.n617 VSUBS 0.007669f
C658 B.n618 VSUBS 0.007669f
C659 B.n619 VSUBS 0.007669f
C660 B.n620 VSUBS 0.007669f
C661 B.n621 VSUBS 0.007669f
C662 B.n622 VSUBS 0.007669f
C663 B.n623 VSUBS 0.007669f
C664 B.n624 VSUBS 0.007669f
C665 B.n625 VSUBS 0.007669f
C666 B.n626 VSUBS 0.007669f
C667 B.n627 VSUBS 0.016491f
C668 B.n628 VSUBS 0.017795f
C669 B.n629 VSUBS 0.017795f
C670 B.n630 VSUBS 0.007669f
C671 B.n631 VSUBS 0.007669f
C672 B.n632 VSUBS 0.007669f
C673 B.n633 VSUBS 0.007669f
C674 B.n634 VSUBS 0.007669f
C675 B.n635 VSUBS 0.007669f
C676 B.n636 VSUBS 0.007669f
C677 B.n637 VSUBS 0.007669f
C678 B.n638 VSUBS 0.007669f
C679 B.n639 VSUBS 0.007669f
C680 B.n640 VSUBS 0.007669f
C681 B.n641 VSUBS 0.007669f
C682 B.n642 VSUBS 0.007669f
C683 B.n643 VSUBS 0.007669f
C684 B.n644 VSUBS 0.007669f
C685 B.n645 VSUBS 0.007669f
C686 B.n646 VSUBS 0.007669f
C687 B.n647 VSUBS 0.007669f
C688 B.n648 VSUBS 0.007669f
C689 B.n649 VSUBS 0.007669f
C690 B.n650 VSUBS 0.007669f
C691 B.n651 VSUBS 0.007669f
C692 B.n652 VSUBS 0.007669f
C693 B.n653 VSUBS 0.007669f
C694 B.n654 VSUBS 0.007669f
C695 B.n655 VSUBS 0.007669f
C696 B.n656 VSUBS 0.007669f
C697 B.n657 VSUBS 0.007669f
C698 B.n658 VSUBS 0.007669f
C699 B.n659 VSUBS 0.007669f
C700 B.n660 VSUBS 0.007669f
C701 B.n661 VSUBS 0.007669f
C702 B.n662 VSUBS 0.007669f
C703 B.n663 VSUBS 0.007669f
C704 B.n664 VSUBS 0.007669f
C705 B.n665 VSUBS 0.007669f
C706 B.n666 VSUBS 0.007669f
C707 B.n667 VSUBS 0.007669f
C708 B.n668 VSUBS 0.007669f
C709 B.n669 VSUBS 0.007669f
C710 B.n670 VSUBS 0.007669f
C711 B.n671 VSUBS 0.007669f
C712 B.n672 VSUBS 0.007669f
C713 B.n673 VSUBS 0.007669f
C714 B.n674 VSUBS 0.007669f
C715 B.n675 VSUBS 0.007669f
C716 B.n676 VSUBS 0.007669f
C717 B.n677 VSUBS 0.007669f
C718 B.n678 VSUBS 0.007669f
C719 B.n679 VSUBS 0.007669f
C720 B.n680 VSUBS 0.007669f
C721 B.n681 VSUBS 0.007669f
C722 B.n682 VSUBS 0.007218f
C723 B.n683 VSUBS 0.007669f
C724 B.n684 VSUBS 0.007669f
C725 B.n685 VSUBS 0.007669f
C726 B.n686 VSUBS 0.007669f
C727 B.n687 VSUBS 0.007669f
C728 B.n688 VSUBS 0.007669f
C729 B.n689 VSUBS 0.007669f
C730 B.n690 VSUBS 0.007669f
C731 B.n691 VSUBS 0.007669f
C732 B.n692 VSUBS 0.007669f
C733 B.n693 VSUBS 0.007669f
C734 B.n694 VSUBS 0.007669f
C735 B.n695 VSUBS 0.007669f
C736 B.n696 VSUBS 0.007669f
C737 B.n697 VSUBS 0.007669f
C738 B.n698 VSUBS 0.004286f
C739 B.n699 VSUBS 0.017769f
C740 B.n700 VSUBS 0.007218f
C741 B.n701 VSUBS 0.007669f
C742 B.n702 VSUBS 0.007669f
C743 B.n703 VSUBS 0.007669f
C744 B.n704 VSUBS 0.007669f
C745 B.n705 VSUBS 0.007669f
C746 B.n706 VSUBS 0.007669f
C747 B.n707 VSUBS 0.007669f
C748 B.n708 VSUBS 0.007669f
C749 B.n709 VSUBS 0.007669f
C750 B.n710 VSUBS 0.007669f
C751 B.n711 VSUBS 0.007669f
C752 B.n712 VSUBS 0.007669f
C753 B.n713 VSUBS 0.007669f
C754 B.n714 VSUBS 0.007669f
C755 B.n715 VSUBS 0.007669f
C756 B.n716 VSUBS 0.007669f
C757 B.n717 VSUBS 0.007669f
C758 B.n718 VSUBS 0.007669f
C759 B.n719 VSUBS 0.007669f
C760 B.n720 VSUBS 0.007669f
C761 B.n721 VSUBS 0.007669f
C762 B.n722 VSUBS 0.007669f
C763 B.n723 VSUBS 0.007669f
C764 B.n724 VSUBS 0.007669f
C765 B.n725 VSUBS 0.007669f
C766 B.n726 VSUBS 0.007669f
C767 B.n727 VSUBS 0.007669f
C768 B.n728 VSUBS 0.007669f
C769 B.n729 VSUBS 0.007669f
C770 B.n730 VSUBS 0.007669f
C771 B.n731 VSUBS 0.007669f
C772 B.n732 VSUBS 0.007669f
C773 B.n733 VSUBS 0.007669f
C774 B.n734 VSUBS 0.007669f
C775 B.n735 VSUBS 0.007669f
C776 B.n736 VSUBS 0.007669f
C777 B.n737 VSUBS 0.007669f
C778 B.n738 VSUBS 0.007669f
C779 B.n739 VSUBS 0.007669f
C780 B.n740 VSUBS 0.007669f
C781 B.n741 VSUBS 0.007669f
C782 B.n742 VSUBS 0.007669f
C783 B.n743 VSUBS 0.007669f
C784 B.n744 VSUBS 0.007669f
C785 B.n745 VSUBS 0.007669f
C786 B.n746 VSUBS 0.007669f
C787 B.n747 VSUBS 0.007669f
C788 B.n748 VSUBS 0.007669f
C789 B.n749 VSUBS 0.007669f
C790 B.n750 VSUBS 0.007669f
C791 B.n751 VSUBS 0.007669f
C792 B.n752 VSUBS 0.007669f
C793 B.n753 VSUBS 0.007669f
C794 B.n754 VSUBS 0.017795f
C795 B.n755 VSUBS 0.016491f
C796 B.n756 VSUBS 0.016491f
C797 B.n757 VSUBS 0.007669f
C798 B.n758 VSUBS 0.007669f
C799 B.n759 VSUBS 0.007669f
C800 B.n760 VSUBS 0.007669f
C801 B.n761 VSUBS 0.007669f
C802 B.n762 VSUBS 0.007669f
C803 B.n763 VSUBS 0.007669f
C804 B.n764 VSUBS 0.007669f
C805 B.n765 VSUBS 0.007669f
C806 B.n766 VSUBS 0.007669f
C807 B.n767 VSUBS 0.007669f
C808 B.n768 VSUBS 0.007669f
C809 B.n769 VSUBS 0.007669f
C810 B.n770 VSUBS 0.007669f
C811 B.n771 VSUBS 0.007669f
C812 B.n772 VSUBS 0.007669f
C813 B.n773 VSUBS 0.007669f
C814 B.n774 VSUBS 0.007669f
C815 B.n775 VSUBS 0.007669f
C816 B.n776 VSUBS 0.007669f
C817 B.n777 VSUBS 0.007669f
C818 B.n778 VSUBS 0.007669f
C819 B.n779 VSUBS 0.007669f
C820 B.n780 VSUBS 0.007669f
C821 B.n781 VSUBS 0.007669f
C822 B.n782 VSUBS 0.007669f
C823 B.n783 VSUBS 0.007669f
C824 B.n784 VSUBS 0.007669f
C825 B.n785 VSUBS 0.007669f
C826 B.n786 VSUBS 0.007669f
C827 B.n787 VSUBS 0.007669f
C828 B.n788 VSUBS 0.007669f
C829 B.n789 VSUBS 0.007669f
C830 B.n790 VSUBS 0.007669f
C831 B.n791 VSUBS 0.007669f
C832 B.n792 VSUBS 0.007669f
C833 B.n793 VSUBS 0.007669f
C834 B.n794 VSUBS 0.007669f
C835 B.n795 VSUBS 0.007669f
C836 B.n796 VSUBS 0.007669f
C837 B.n797 VSUBS 0.007669f
C838 B.n798 VSUBS 0.007669f
C839 B.n799 VSUBS 0.007669f
C840 B.n800 VSUBS 0.007669f
C841 B.n801 VSUBS 0.007669f
C842 B.n802 VSUBS 0.007669f
C843 B.n803 VSUBS 0.007669f
C844 B.n804 VSUBS 0.007669f
C845 B.n805 VSUBS 0.007669f
C846 B.n806 VSUBS 0.007669f
C847 B.n807 VSUBS 0.007669f
C848 B.n808 VSUBS 0.007669f
C849 B.n809 VSUBS 0.007669f
C850 B.n810 VSUBS 0.007669f
C851 B.n811 VSUBS 0.007669f
C852 B.n812 VSUBS 0.007669f
C853 B.n813 VSUBS 0.007669f
C854 B.n814 VSUBS 0.007669f
C855 B.n815 VSUBS 0.007669f
C856 B.n816 VSUBS 0.007669f
C857 B.n817 VSUBS 0.007669f
C858 B.n818 VSUBS 0.007669f
C859 B.n819 VSUBS 0.007669f
C860 B.n820 VSUBS 0.007669f
C861 B.n821 VSUBS 0.007669f
C862 B.n822 VSUBS 0.007669f
C863 B.n823 VSUBS 0.007669f
C864 B.n824 VSUBS 0.007669f
C865 B.n825 VSUBS 0.007669f
C866 B.n826 VSUBS 0.007669f
C867 B.n827 VSUBS 0.007669f
C868 B.n828 VSUBS 0.007669f
C869 B.n829 VSUBS 0.007669f
C870 B.n830 VSUBS 0.007669f
C871 B.n831 VSUBS 0.007669f
C872 B.n832 VSUBS 0.007669f
C873 B.n833 VSUBS 0.007669f
C874 B.n834 VSUBS 0.007669f
C875 B.n835 VSUBS 0.007669f
C876 B.n836 VSUBS 0.007669f
C877 B.n837 VSUBS 0.007669f
C878 B.n838 VSUBS 0.007669f
C879 B.n839 VSUBS 0.007669f
C880 B.n840 VSUBS 0.007669f
C881 B.n841 VSUBS 0.007669f
C882 B.n842 VSUBS 0.007669f
C883 B.n843 VSUBS 0.007669f
C884 B.n844 VSUBS 0.007669f
C885 B.n845 VSUBS 0.007669f
C886 B.n846 VSUBS 0.007669f
C887 B.n847 VSUBS 0.010008f
C888 B.n848 VSUBS 0.010661f
C889 B.n849 VSUBS 0.0212f
C890 VDD2.t1 VSUBS 0.255585f
C891 VDD2.t7 VSUBS 0.255585f
C892 VDD2.n0 VSUBS 1.97291f
C893 VDD2.t4 VSUBS 0.255585f
C894 VDD2.t0 VSUBS 0.255585f
C895 VDD2.n1 VSUBS 1.97291f
C896 VDD2.n2 VSUBS 5.09704f
C897 VDD2.t6 VSUBS 0.255585f
C898 VDD2.t2 VSUBS 0.255585f
C899 VDD2.n3 VSUBS 1.95287f
C900 VDD2.n4 VSUBS 4.14529f
C901 VDD2.t5 VSUBS 0.255585f
C902 VDD2.t3 VSUBS 0.255585f
C903 VDD2.n5 VSUBS 1.97285f
C904 VN.t7 VSUBS 2.53797f
C905 VN.n0 VSUBS 1.00517f
C906 VN.n1 VSUBS 0.026616f
C907 VN.n2 VSUBS 0.022383f
C908 VN.n3 VSUBS 0.026616f
C909 VN.t3 VSUBS 2.53797f
C910 VN.n4 VSUBS 0.898412f
C911 VN.n5 VSUBS 0.026616f
C912 VN.n6 VSUBS 0.038854f
C913 VN.n7 VSUBS 0.026616f
C914 VN.n8 VSUBS 0.030013f
C915 VN.t0 VSUBS 2.53797f
C916 VN.n9 VSUBS 0.981754f
C917 VN.t6 VSUBS 2.87158f
C918 VN.n10 VSUBS 0.934966f
C919 VN.n11 VSUBS 0.31516f
C920 VN.n12 VSUBS 0.026616f
C921 VN.n13 VSUBS 0.049605f
C922 VN.n14 VSUBS 0.049605f
C923 VN.n15 VSUBS 0.038854f
C924 VN.n16 VSUBS 0.026616f
C925 VN.n17 VSUBS 0.026616f
C926 VN.n18 VSUBS 0.026616f
C927 VN.n19 VSUBS 0.049605f
C928 VN.n20 VSUBS 0.049605f
C929 VN.n21 VSUBS 0.030013f
C930 VN.n22 VSUBS 0.026616f
C931 VN.n23 VSUBS 0.026616f
C932 VN.n24 VSUBS 0.044707f
C933 VN.n25 VSUBS 0.049605f
C934 VN.n26 VSUBS 0.051182f
C935 VN.n27 VSUBS 0.026616f
C936 VN.n28 VSUBS 0.026616f
C937 VN.n29 VSUBS 0.026616f
C938 VN.n30 VSUBS 0.053748f
C939 VN.n31 VSUBS 0.049605f
C940 VN.n32 VSUBS 0.039809f
C941 VN.n33 VSUBS 0.042957f
C942 VN.n34 VSUBS 0.065171f
C943 VN.t1 VSUBS 2.53797f
C944 VN.n35 VSUBS 1.00517f
C945 VN.n36 VSUBS 0.026616f
C946 VN.n37 VSUBS 0.022383f
C947 VN.n38 VSUBS 0.026616f
C948 VN.t5 VSUBS 2.53797f
C949 VN.n39 VSUBS 0.898412f
C950 VN.n40 VSUBS 0.026616f
C951 VN.n41 VSUBS 0.038854f
C952 VN.n42 VSUBS 0.026616f
C953 VN.n43 VSUBS 0.030013f
C954 VN.t4 VSUBS 2.87158f
C955 VN.t2 VSUBS 2.53797f
C956 VN.n44 VSUBS 0.981754f
C957 VN.n45 VSUBS 0.934966f
C958 VN.n46 VSUBS 0.31516f
C959 VN.n47 VSUBS 0.026616f
C960 VN.n48 VSUBS 0.049605f
C961 VN.n49 VSUBS 0.049605f
C962 VN.n50 VSUBS 0.038854f
C963 VN.n51 VSUBS 0.026616f
C964 VN.n52 VSUBS 0.026616f
C965 VN.n53 VSUBS 0.026616f
C966 VN.n54 VSUBS 0.049605f
C967 VN.n55 VSUBS 0.049605f
C968 VN.n56 VSUBS 0.030013f
C969 VN.n57 VSUBS 0.026616f
C970 VN.n58 VSUBS 0.026616f
C971 VN.n59 VSUBS 0.044707f
C972 VN.n60 VSUBS 0.049605f
C973 VN.n61 VSUBS 0.051182f
C974 VN.n62 VSUBS 0.026616f
C975 VN.n63 VSUBS 0.026616f
C976 VN.n64 VSUBS 0.026616f
C977 VN.n65 VSUBS 0.053748f
C978 VN.n66 VSUBS 0.049605f
C979 VN.n67 VSUBS 0.039809f
C980 VN.n68 VSUBS 0.042957f
C981 VN.n69 VSUBS 1.67586f
C982 VDD1.t2 VSUBS 0.256645f
C983 VDD1.t4 VSUBS 0.256645f
C984 VDD1.n0 VSUBS 1.98277f
C985 VDD1.t1 VSUBS 0.256645f
C986 VDD1.t5 VSUBS 0.256645f
C987 VDD1.n1 VSUBS 1.98109f
C988 VDD1.t0 VSUBS 0.256645f
C989 VDD1.t3 VSUBS 0.256645f
C990 VDD1.n2 VSUBS 1.98109f
C991 VDD1.n3 VSUBS 5.18258f
C992 VDD1.t6 VSUBS 0.256645f
C993 VDD1.t7 VSUBS 0.256645f
C994 VDD1.n4 VSUBS 1.96096f
C995 VDD1.n5 VSUBS 4.20141f
C996 VTAIL.t0 VSUBS 0.218689f
C997 VTAIL.t14 VSUBS 0.218689f
C998 VTAIL.n0 VSUBS 1.54372f
C999 VTAIL.n1 VSUBS 0.846274f
C1000 VTAIL.t15 VSUBS 2.04807f
C1001 VTAIL.n2 VSUBS 0.973538f
C1002 VTAIL.t10 VSUBS 2.04807f
C1003 VTAIL.n3 VSUBS 0.973538f
C1004 VTAIL.t9 VSUBS 0.218689f
C1005 VTAIL.t11 VSUBS 0.218689f
C1006 VTAIL.n4 VSUBS 1.54372f
C1007 VTAIL.n5 VSUBS 1.114f
C1008 VTAIL.t8 VSUBS 2.04807f
C1009 VTAIL.n6 VSUBS 2.33522f
C1010 VTAIL.t1 VSUBS 2.04808f
C1011 VTAIL.n7 VSUBS 2.33521f
C1012 VTAIL.t4 VSUBS 0.218689f
C1013 VTAIL.t2 VSUBS 0.218689f
C1014 VTAIL.n8 VSUBS 1.54372f
C1015 VTAIL.n9 VSUBS 1.114f
C1016 VTAIL.t13 VSUBS 2.04808f
C1017 VTAIL.n10 VSUBS 0.973532f
C1018 VTAIL.t5 VSUBS 2.04808f
C1019 VTAIL.n11 VSUBS 0.973532f
C1020 VTAIL.t6 VSUBS 0.218689f
C1021 VTAIL.t12 VSUBS 0.218689f
C1022 VTAIL.n12 VSUBS 1.54372f
C1023 VTAIL.n13 VSUBS 1.114f
C1024 VTAIL.t7 VSUBS 2.04807f
C1025 VTAIL.n14 VSUBS 2.33522f
C1026 VTAIL.t3 VSUBS 2.04807f
C1027 VTAIL.n15 VSUBS 2.33025f
C1028 VP.t4 VSUBS 2.78966f
C1029 VP.n0 VSUBS 1.10485f
C1030 VP.n1 VSUBS 0.029255f
C1031 VP.n2 VSUBS 0.024603f
C1032 VP.n3 VSUBS 0.029255f
C1033 VP.t7 VSUBS 2.78966f
C1034 VP.n4 VSUBS 0.987505f
C1035 VP.n5 VSUBS 0.029255f
C1036 VP.n6 VSUBS 0.042707f
C1037 VP.n7 VSUBS 0.029255f
C1038 VP.n8 VSUBS 0.032989f
C1039 VP.n9 VSUBS 0.029255f
C1040 VP.n10 VSUBS 0.024603f
C1041 VP.n11 VSUBS 0.029255f
C1042 VP.t6 VSUBS 2.78966f
C1043 VP.n12 VSUBS 1.10485f
C1044 VP.t0 VSUBS 2.78966f
C1045 VP.n13 VSUBS 1.10485f
C1046 VP.n14 VSUBS 0.029255f
C1047 VP.n15 VSUBS 0.024603f
C1048 VP.n16 VSUBS 0.029255f
C1049 VP.t1 VSUBS 2.78966f
C1050 VP.n17 VSUBS 0.987505f
C1051 VP.n18 VSUBS 0.029255f
C1052 VP.n19 VSUBS 0.042707f
C1053 VP.n20 VSUBS 0.029255f
C1054 VP.n21 VSUBS 0.032989f
C1055 VP.t5 VSUBS 3.15635f
C1056 VP.t3 VSUBS 2.78966f
C1057 VP.n22 VSUBS 1.07911f
C1058 VP.n23 VSUBS 1.02769f
C1059 VP.n24 VSUBS 0.346415f
C1060 VP.n25 VSUBS 0.029255f
C1061 VP.n26 VSUBS 0.054524f
C1062 VP.n27 VSUBS 0.054524f
C1063 VP.n28 VSUBS 0.042707f
C1064 VP.n29 VSUBS 0.029255f
C1065 VP.n30 VSUBS 0.029255f
C1066 VP.n31 VSUBS 0.029255f
C1067 VP.n32 VSUBS 0.054524f
C1068 VP.n33 VSUBS 0.054524f
C1069 VP.n34 VSUBS 0.032989f
C1070 VP.n35 VSUBS 0.029255f
C1071 VP.n36 VSUBS 0.029255f
C1072 VP.n37 VSUBS 0.049141f
C1073 VP.n38 VSUBS 0.054524f
C1074 VP.n39 VSUBS 0.056257f
C1075 VP.n40 VSUBS 0.029255f
C1076 VP.n41 VSUBS 0.029255f
C1077 VP.n42 VSUBS 0.029255f
C1078 VP.n43 VSUBS 0.059078f
C1079 VP.n44 VSUBS 0.054524f
C1080 VP.n45 VSUBS 0.043757f
C1081 VP.n46 VSUBS 0.047217f
C1082 VP.n47 VSUBS 1.83035f
C1083 VP.n48 VSUBS 1.85003f
C1084 VP.n49 VSUBS 0.047217f
C1085 VP.n50 VSUBS 0.043757f
C1086 VP.n51 VSUBS 0.054524f
C1087 VP.n52 VSUBS 0.059078f
C1088 VP.n53 VSUBS 0.029255f
C1089 VP.n54 VSUBS 0.029255f
C1090 VP.n55 VSUBS 0.029255f
C1091 VP.n56 VSUBS 0.056257f
C1092 VP.n57 VSUBS 0.054524f
C1093 VP.t2 VSUBS 2.78966f
C1094 VP.n58 VSUBS 0.987505f
C1095 VP.n59 VSUBS 0.049141f
C1096 VP.n60 VSUBS 0.029255f
C1097 VP.n61 VSUBS 0.029255f
C1098 VP.n62 VSUBS 0.029255f
C1099 VP.n63 VSUBS 0.054524f
C1100 VP.n64 VSUBS 0.054524f
C1101 VP.n65 VSUBS 0.042707f
C1102 VP.n66 VSUBS 0.029255f
C1103 VP.n67 VSUBS 0.029255f
C1104 VP.n68 VSUBS 0.029255f
C1105 VP.n69 VSUBS 0.054524f
C1106 VP.n70 VSUBS 0.054524f
C1107 VP.n71 VSUBS 0.032989f
C1108 VP.n72 VSUBS 0.029255f
C1109 VP.n73 VSUBS 0.029255f
C1110 VP.n74 VSUBS 0.049141f
C1111 VP.n75 VSUBS 0.054524f
C1112 VP.n76 VSUBS 0.056257f
C1113 VP.n77 VSUBS 0.029255f
C1114 VP.n78 VSUBS 0.029255f
C1115 VP.n79 VSUBS 0.029255f
C1116 VP.n80 VSUBS 0.059078f
C1117 VP.n81 VSUBS 0.054524f
C1118 VP.n82 VSUBS 0.043757f
C1119 VP.n83 VSUBS 0.047217f
C1120 VP.n84 VSUBS 0.071633f
.ends

