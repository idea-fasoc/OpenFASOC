* NGSPICE file created from diff_pair_sample_1422.ext - technology: sky130A

.subckt diff_pair_sample_1422 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=0 ps=0 w=14.58 l=2.28
X1 VDD2.t5 VN.t0 VTAIL.t5 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=2.4057 ps=14.91 w=14.58 l=2.28
X2 B.t8 B.t6 B.t7 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=0 ps=0 w=14.58 l=2.28
X3 B.t5 B.t3 B.t4 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=0 ps=0 w=14.58 l=2.28
X4 VDD2.t4 VN.t1 VTAIL.t6 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=5.6862 ps=29.94 w=14.58 l=2.28
X5 VTAIL.t3 VP.t0 VDD1.t5 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=2.4057 ps=14.91 w=14.58 l=2.28
X6 B.t2 B.t0 B.t1 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=0 ps=0 w=14.58 l=2.28
X7 VTAIL.t4 VP.t1 VDD1.t4 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=2.4057 ps=14.91 w=14.58 l=2.28
X8 VTAIL.t10 VN.t2 VDD2.t3 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=2.4057 ps=14.91 w=14.58 l=2.28
X9 VDD1.t3 VP.t2 VTAIL.t2 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=2.4057 ps=14.91 w=14.58 l=2.28
X10 VDD1.t2 VP.t3 VTAIL.t11 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=5.6862 ps=29.94 w=14.58 l=2.28
X11 VTAIL.t8 VN.t3 VDD2.t2 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=2.4057 ps=14.91 w=14.58 l=2.28
X12 VDD2.t1 VN.t4 VTAIL.t7 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=5.6862 ps=29.94 w=14.58 l=2.28
X13 VDD2.t0 VN.t5 VTAIL.t9 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=2.4057 ps=14.91 w=14.58 l=2.28
X14 VDD1.t1 VP.t4 VTAIL.t1 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=5.6862 pd=29.94 as=2.4057 ps=14.91 w=14.58 l=2.28
X15 VDD1.t0 VP.t5 VTAIL.t0 w_n3058_n3884# sky130_fd_pr__pfet_01v8 ad=2.4057 pd=14.91 as=5.6862 ps=29.94 w=14.58 l=2.28
R0 B.n537 B.n536 585
R1 B.n538 B.n79 585
R2 B.n540 B.n539 585
R3 B.n541 B.n78 585
R4 B.n543 B.n542 585
R5 B.n544 B.n77 585
R6 B.n546 B.n545 585
R7 B.n547 B.n76 585
R8 B.n549 B.n548 585
R9 B.n550 B.n75 585
R10 B.n552 B.n551 585
R11 B.n553 B.n74 585
R12 B.n555 B.n554 585
R13 B.n556 B.n73 585
R14 B.n558 B.n557 585
R15 B.n559 B.n72 585
R16 B.n561 B.n560 585
R17 B.n562 B.n71 585
R18 B.n564 B.n563 585
R19 B.n565 B.n70 585
R20 B.n567 B.n566 585
R21 B.n568 B.n69 585
R22 B.n570 B.n569 585
R23 B.n571 B.n68 585
R24 B.n573 B.n572 585
R25 B.n574 B.n67 585
R26 B.n576 B.n575 585
R27 B.n577 B.n66 585
R28 B.n579 B.n578 585
R29 B.n580 B.n65 585
R30 B.n582 B.n581 585
R31 B.n583 B.n64 585
R32 B.n585 B.n584 585
R33 B.n586 B.n63 585
R34 B.n588 B.n587 585
R35 B.n589 B.n62 585
R36 B.n591 B.n590 585
R37 B.n592 B.n61 585
R38 B.n594 B.n593 585
R39 B.n595 B.n60 585
R40 B.n597 B.n596 585
R41 B.n598 B.n59 585
R42 B.n600 B.n599 585
R43 B.n601 B.n58 585
R44 B.n603 B.n602 585
R45 B.n604 B.n57 585
R46 B.n606 B.n605 585
R47 B.n607 B.n56 585
R48 B.n609 B.n608 585
R49 B.n611 B.n53 585
R50 B.n613 B.n612 585
R51 B.n614 B.n52 585
R52 B.n616 B.n615 585
R53 B.n617 B.n51 585
R54 B.n619 B.n618 585
R55 B.n620 B.n50 585
R56 B.n622 B.n621 585
R57 B.n623 B.n49 585
R58 B.n625 B.n624 585
R59 B.n627 B.n626 585
R60 B.n628 B.n45 585
R61 B.n630 B.n629 585
R62 B.n631 B.n44 585
R63 B.n633 B.n632 585
R64 B.n634 B.n43 585
R65 B.n636 B.n635 585
R66 B.n637 B.n42 585
R67 B.n639 B.n638 585
R68 B.n640 B.n41 585
R69 B.n642 B.n641 585
R70 B.n643 B.n40 585
R71 B.n645 B.n644 585
R72 B.n646 B.n39 585
R73 B.n648 B.n647 585
R74 B.n649 B.n38 585
R75 B.n651 B.n650 585
R76 B.n652 B.n37 585
R77 B.n654 B.n653 585
R78 B.n655 B.n36 585
R79 B.n657 B.n656 585
R80 B.n658 B.n35 585
R81 B.n660 B.n659 585
R82 B.n661 B.n34 585
R83 B.n663 B.n662 585
R84 B.n664 B.n33 585
R85 B.n666 B.n665 585
R86 B.n667 B.n32 585
R87 B.n669 B.n668 585
R88 B.n670 B.n31 585
R89 B.n672 B.n671 585
R90 B.n673 B.n30 585
R91 B.n675 B.n674 585
R92 B.n676 B.n29 585
R93 B.n678 B.n677 585
R94 B.n679 B.n28 585
R95 B.n681 B.n680 585
R96 B.n682 B.n27 585
R97 B.n684 B.n683 585
R98 B.n685 B.n26 585
R99 B.n687 B.n686 585
R100 B.n688 B.n25 585
R101 B.n690 B.n689 585
R102 B.n691 B.n24 585
R103 B.n693 B.n692 585
R104 B.n694 B.n23 585
R105 B.n696 B.n695 585
R106 B.n697 B.n22 585
R107 B.n699 B.n698 585
R108 B.n535 B.n80 585
R109 B.n534 B.n533 585
R110 B.n532 B.n81 585
R111 B.n531 B.n530 585
R112 B.n529 B.n82 585
R113 B.n528 B.n527 585
R114 B.n526 B.n83 585
R115 B.n525 B.n524 585
R116 B.n523 B.n84 585
R117 B.n522 B.n521 585
R118 B.n520 B.n85 585
R119 B.n519 B.n518 585
R120 B.n517 B.n86 585
R121 B.n516 B.n515 585
R122 B.n514 B.n87 585
R123 B.n513 B.n512 585
R124 B.n511 B.n88 585
R125 B.n510 B.n509 585
R126 B.n508 B.n89 585
R127 B.n507 B.n506 585
R128 B.n505 B.n90 585
R129 B.n504 B.n503 585
R130 B.n502 B.n91 585
R131 B.n501 B.n500 585
R132 B.n499 B.n92 585
R133 B.n498 B.n497 585
R134 B.n496 B.n93 585
R135 B.n495 B.n494 585
R136 B.n493 B.n94 585
R137 B.n492 B.n491 585
R138 B.n490 B.n95 585
R139 B.n489 B.n488 585
R140 B.n487 B.n96 585
R141 B.n486 B.n485 585
R142 B.n484 B.n97 585
R143 B.n483 B.n482 585
R144 B.n481 B.n98 585
R145 B.n480 B.n479 585
R146 B.n478 B.n99 585
R147 B.n477 B.n476 585
R148 B.n475 B.n100 585
R149 B.n474 B.n473 585
R150 B.n472 B.n101 585
R151 B.n471 B.n470 585
R152 B.n469 B.n102 585
R153 B.n468 B.n467 585
R154 B.n466 B.n103 585
R155 B.n465 B.n464 585
R156 B.n463 B.n104 585
R157 B.n462 B.n461 585
R158 B.n460 B.n105 585
R159 B.n459 B.n458 585
R160 B.n457 B.n106 585
R161 B.n456 B.n455 585
R162 B.n454 B.n107 585
R163 B.n453 B.n452 585
R164 B.n451 B.n108 585
R165 B.n450 B.n449 585
R166 B.n448 B.n109 585
R167 B.n447 B.n446 585
R168 B.n445 B.n110 585
R169 B.n444 B.n443 585
R170 B.n442 B.n111 585
R171 B.n441 B.n440 585
R172 B.n439 B.n112 585
R173 B.n438 B.n437 585
R174 B.n436 B.n113 585
R175 B.n435 B.n434 585
R176 B.n433 B.n114 585
R177 B.n432 B.n431 585
R178 B.n430 B.n115 585
R179 B.n429 B.n428 585
R180 B.n427 B.n116 585
R181 B.n426 B.n425 585
R182 B.n424 B.n117 585
R183 B.n423 B.n422 585
R184 B.n421 B.n118 585
R185 B.n420 B.n419 585
R186 B.n418 B.n119 585
R187 B.n255 B.n254 585
R188 B.n256 B.n177 585
R189 B.n258 B.n257 585
R190 B.n259 B.n176 585
R191 B.n261 B.n260 585
R192 B.n262 B.n175 585
R193 B.n264 B.n263 585
R194 B.n265 B.n174 585
R195 B.n267 B.n266 585
R196 B.n268 B.n173 585
R197 B.n270 B.n269 585
R198 B.n271 B.n172 585
R199 B.n273 B.n272 585
R200 B.n274 B.n171 585
R201 B.n276 B.n275 585
R202 B.n277 B.n170 585
R203 B.n279 B.n278 585
R204 B.n280 B.n169 585
R205 B.n282 B.n281 585
R206 B.n283 B.n168 585
R207 B.n285 B.n284 585
R208 B.n286 B.n167 585
R209 B.n288 B.n287 585
R210 B.n289 B.n166 585
R211 B.n291 B.n290 585
R212 B.n292 B.n165 585
R213 B.n294 B.n293 585
R214 B.n295 B.n164 585
R215 B.n297 B.n296 585
R216 B.n298 B.n163 585
R217 B.n300 B.n299 585
R218 B.n301 B.n162 585
R219 B.n303 B.n302 585
R220 B.n304 B.n161 585
R221 B.n306 B.n305 585
R222 B.n307 B.n160 585
R223 B.n309 B.n308 585
R224 B.n310 B.n159 585
R225 B.n312 B.n311 585
R226 B.n313 B.n158 585
R227 B.n315 B.n314 585
R228 B.n316 B.n157 585
R229 B.n318 B.n317 585
R230 B.n319 B.n156 585
R231 B.n321 B.n320 585
R232 B.n322 B.n155 585
R233 B.n324 B.n323 585
R234 B.n325 B.n154 585
R235 B.n327 B.n326 585
R236 B.n329 B.n151 585
R237 B.n331 B.n330 585
R238 B.n332 B.n150 585
R239 B.n334 B.n333 585
R240 B.n335 B.n149 585
R241 B.n337 B.n336 585
R242 B.n338 B.n148 585
R243 B.n340 B.n339 585
R244 B.n341 B.n147 585
R245 B.n343 B.n342 585
R246 B.n345 B.n344 585
R247 B.n346 B.n143 585
R248 B.n348 B.n347 585
R249 B.n349 B.n142 585
R250 B.n351 B.n350 585
R251 B.n352 B.n141 585
R252 B.n354 B.n353 585
R253 B.n355 B.n140 585
R254 B.n357 B.n356 585
R255 B.n358 B.n139 585
R256 B.n360 B.n359 585
R257 B.n361 B.n138 585
R258 B.n363 B.n362 585
R259 B.n364 B.n137 585
R260 B.n366 B.n365 585
R261 B.n367 B.n136 585
R262 B.n369 B.n368 585
R263 B.n370 B.n135 585
R264 B.n372 B.n371 585
R265 B.n373 B.n134 585
R266 B.n375 B.n374 585
R267 B.n376 B.n133 585
R268 B.n378 B.n377 585
R269 B.n379 B.n132 585
R270 B.n381 B.n380 585
R271 B.n382 B.n131 585
R272 B.n384 B.n383 585
R273 B.n385 B.n130 585
R274 B.n387 B.n386 585
R275 B.n388 B.n129 585
R276 B.n390 B.n389 585
R277 B.n391 B.n128 585
R278 B.n393 B.n392 585
R279 B.n394 B.n127 585
R280 B.n396 B.n395 585
R281 B.n397 B.n126 585
R282 B.n399 B.n398 585
R283 B.n400 B.n125 585
R284 B.n402 B.n401 585
R285 B.n403 B.n124 585
R286 B.n405 B.n404 585
R287 B.n406 B.n123 585
R288 B.n408 B.n407 585
R289 B.n409 B.n122 585
R290 B.n411 B.n410 585
R291 B.n412 B.n121 585
R292 B.n414 B.n413 585
R293 B.n415 B.n120 585
R294 B.n417 B.n416 585
R295 B.n253 B.n178 585
R296 B.n252 B.n251 585
R297 B.n250 B.n179 585
R298 B.n249 B.n248 585
R299 B.n247 B.n180 585
R300 B.n246 B.n245 585
R301 B.n244 B.n181 585
R302 B.n243 B.n242 585
R303 B.n241 B.n182 585
R304 B.n240 B.n239 585
R305 B.n238 B.n183 585
R306 B.n237 B.n236 585
R307 B.n235 B.n184 585
R308 B.n234 B.n233 585
R309 B.n232 B.n185 585
R310 B.n231 B.n230 585
R311 B.n229 B.n186 585
R312 B.n228 B.n227 585
R313 B.n226 B.n187 585
R314 B.n225 B.n224 585
R315 B.n223 B.n188 585
R316 B.n222 B.n221 585
R317 B.n220 B.n189 585
R318 B.n219 B.n218 585
R319 B.n217 B.n190 585
R320 B.n216 B.n215 585
R321 B.n214 B.n191 585
R322 B.n213 B.n212 585
R323 B.n211 B.n192 585
R324 B.n210 B.n209 585
R325 B.n208 B.n193 585
R326 B.n207 B.n206 585
R327 B.n205 B.n194 585
R328 B.n204 B.n203 585
R329 B.n202 B.n195 585
R330 B.n201 B.n200 585
R331 B.n199 B.n196 585
R332 B.n198 B.n197 585
R333 B.n2 B.n0 585
R334 B.n757 B.n1 585
R335 B.n756 B.n755 585
R336 B.n754 B.n3 585
R337 B.n753 B.n752 585
R338 B.n751 B.n4 585
R339 B.n750 B.n749 585
R340 B.n748 B.n5 585
R341 B.n747 B.n746 585
R342 B.n745 B.n6 585
R343 B.n744 B.n743 585
R344 B.n742 B.n7 585
R345 B.n741 B.n740 585
R346 B.n739 B.n8 585
R347 B.n738 B.n737 585
R348 B.n736 B.n9 585
R349 B.n735 B.n734 585
R350 B.n733 B.n10 585
R351 B.n732 B.n731 585
R352 B.n730 B.n11 585
R353 B.n729 B.n728 585
R354 B.n727 B.n12 585
R355 B.n726 B.n725 585
R356 B.n724 B.n13 585
R357 B.n723 B.n722 585
R358 B.n721 B.n14 585
R359 B.n720 B.n719 585
R360 B.n718 B.n15 585
R361 B.n717 B.n716 585
R362 B.n715 B.n16 585
R363 B.n714 B.n713 585
R364 B.n712 B.n17 585
R365 B.n711 B.n710 585
R366 B.n709 B.n18 585
R367 B.n708 B.n707 585
R368 B.n706 B.n19 585
R369 B.n705 B.n704 585
R370 B.n703 B.n20 585
R371 B.n702 B.n701 585
R372 B.n700 B.n21 585
R373 B.n759 B.n758 585
R374 B.n254 B.n253 468.476
R375 B.n698 B.n21 468.476
R376 B.n416 B.n119 468.476
R377 B.n536 B.n535 468.476
R378 B.n144 B.t0 361.62
R379 B.n152 B.t6 361.62
R380 B.n46 B.t3 361.62
R381 B.n54 B.t9 361.62
R382 B.n253 B.n252 163.367
R383 B.n252 B.n179 163.367
R384 B.n248 B.n179 163.367
R385 B.n248 B.n247 163.367
R386 B.n247 B.n246 163.367
R387 B.n246 B.n181 163.367
R388 B.n242 B.n181 163.367
R389 B.n242 B.n241 163.367
R390 B.n241 B.n240 163.367
R391 B.n240 B.n183 163.367
R392 B.n236 B.n183 163.367
R393 B.n236 B.n235 163.367
R394 B.n235 B.n234 163.367
R395 B.n234 B.n185 163.367
R396 B.n230 B.n185 163.367
R397 B.n230 B.n229 163.367
R398 B.n229 B.n228 163.367
R399 B.n228 B.n187 163.367
R400 B.n224 B.n187 163.367
R401 B.n224 B.n223 163.367
R402 B.n223 B.n222 163.367
R403 B.n222 B.n189 163.367
R404 B.n218 B.n189 163.367
R405 B.n218 B.n217 163.367
R406 B.n217 B.n216 163.367
R407 B.n216 B.n191 163.367
R408 B.n212 B.n191 163.367
R409 B.n212 B.n211 163.367
R410 B.n211 B.n210 163.367
R411 B.n210 B.n193 163.367
R412 B.n206 B.n193 163.367
R413 B.n206 B.n205 163.367
R414 B.n205 B.n204 163.367
R415 B.n204 B.n195 163.367
R416 B.n200 B.n195 163.367
R417 B.n200 B.n199 163.367
R418 B.n199 B.n198 163.367
R419 B.n198 B.n2 163.367
R420 B.n758 B.n2 163.367
R421 B.n758 B.n757 163.367
R422 B.n757 B.n756 163.367
R423 B.n756 B.n3 163.367
R424 B.n752 B.n3 163.367
R425 B.n752 B.n751 163.367
R426 B.n751 B.n750 163.367
R427 B.n750 B.n5 163.367
R428 B.n746 B.n5 163.367
R429 B.n746 B.n745 163.367
R430 B.n745 B.n744 163.367
R431 B.n744 B.n7 163.367
R432 B.n740 B.n7 163.367
R433 B.n740 B.n739 163.367
R434 B.n739 B.n738 163.367
R435 B.n738 B.n9 163.367
R436 B.n734 B.n9 163.367
R437 B.n734 B.n733 163.367
R438 B.n733 B.n732 163.367
R439 B.n732 B.n11 163.367
R440 B.n728 B.n11 163.367
R441 B.n728 B.n727 163.367
R442 B.n727 B.n726 163.367
R443 B.n726 B.n13 163.367
R444 B.n722 B.n13 163.367
R445 B.n722 B.n721 163.367
R446 B.n721 B.n720 163.367
R447 B.n720 B.n15 163.367
R448 B.n716 B.n15 163.367
R449 B.n716 B.n715 163.367
R450 B.n715 B.n714 163.367
R451 B.n714 B.n17 163.367
R452 B.n710 B.n17 163.367
R453 B.n710 B.n709 163.367
R454 B.n709 B.n708 163.367
R455 B.n708 B.n19 163.367
R456 B.n704 B.n19 163.367
R457 B.n704 B.n703 163.367
R458 B.n703 B.n702 163.367
R459 B.n702 B.n21 163.367
R460 B.n254 B.n177 163.367
R461 B.n258 B.n177 163.367
R462 B.n259 B.n258 163.367
R463 B.n260 B.n259 163.367
R464 B.n260 B.n175 163.367
R465 B.n264 B.n175 163.367
R466 B.n265 B.n264 163.367
R467 B.n266 B.n265 163.367
R468 B.n266 B.n173 163.367
R469 B.n270 B.n173 163.367
R470 B.n271 B.n270 163.367
R471 B.n272 B.n271 163.367
R472 B.n272 B.n171 163.367
R473 B.n276 B.n171 163.367
R474 B.n277 B.n276 163.367
R475 B.n278 B.n277 163.367
R476 B.n278 B.n169 163.367
R477 B.n282 B.n169 163.367
R478 B.n283 B.n282 163.367
R479 B.n284 B.n283 163.367
R480 B.n284 B.n167 163.367
R481 B.n288 B.n167 163.367
R482 B.n289 B.n288 163.367
R483 B.n290 B.n289 163.367
R484 B.n290 B.n165 163.367
R485 B.n294 B.n165 163.367
R486 B.n295 B.n294 163.367
R487 B.n296 B.n295 163.367
R488 B.n296 B.n163 163.367
R489 B.n300 B.n163 163.367
R490 B.n301 B.n300 163.367
R491 B.n302 B.n301 163.367
R492 B.n302 B.n161 163.367
R493 B.n306 B.n161 163.367
R494 B.n307 B.n306 163.367
R495 B.n308 B.n307 163.367
R496 B.n308 B.n159 163.367
R497 B.n312 B.n159 163.367
R498 B.n313 B.n312 163.367
R499 B.n314 B.n313 163.367
R500 B.n314 B.n157 163.367
R501 B.n318 B.n157 163.367
R502 B.n319 B.n318 163.367
R503 B.n320 B.n319 163.367
R504 B.n320 B.n155 163.367
R505 B.n324 B.n155 163.367
R506 B.n325 B.n324 163.367
R507 B.n326 B.n325 163.367
R508 B.n326 B.n151 163.367
R509 B.n331 B.n151 163.367
R510 B.n332 B.n331 163.367
R511 B.n333 B.n332 163.367
R512 B.n333 B.n149 163.367
R513 B.n337 B.n149 163.367
R514 B.n338 B.n337 163.367
R515 B.n339 B.n338 163.367
R516 B.n339 B.n147 163.367
R517 B.n343 B.n147 163.367
R518 B.n344 B.n343 163.367
R519 B.n344 B.n143 163.367
R520 B.n348 B.n143 163.367
R521 B.n349 B.n348 163.367
R522 B.n350 B.n349 163.367
R523 B.n350 B.n141 163.367
R524 B.n354 B.n141 163.367
R525 B.n355 B.n354 163.367
R526 B.n356 B.n355 163.367
R527 B.n356 B.n139 163.367
R528 B.n360 B.n139 163.367
R529 B.n361 B.n360 163.367
R530 B.n362 B.n361 163.367
R531 B.n362 B.n137 163.367
R532 B.n366 B.n137 163.367
R533 B.n367 B.n366 163.367
R534 B.n368 B.n367 163.367
R535 B.n368 B.n135 163.367
R536 B.n372 B.n135 163.367
R537 B.n373 B.n372 163.367
R538 B.n374 B.n373 163.367
R539 B.n374 B.n133 163.367
R540 B.n378 B.n133 163.367
R541 B.n379 B.n378 163.367
R542 B.n380 B.n379 163.367
R543 B.n380 B.n131 163.367
R544 B.n384 B.n131 163.367
R545 B.n385 B.n384 163.367
R546 B.n386 B.n385 163.367
R547 B.n386 B.n129 163.367
R548 B.n390 B.n129 163.367
R549 B.n391 B.n390 163.367
R550 B.n392 B.n391 163.367
R551 B.n392 B.n127 163.367
R552 B.n396 B.n127 163.367
R553 B.n397 B.n396 163.367
R554 B.n398 B.n397 163.367
R555 B.n398 B.n125 163.367
R556 B.n402 B.n125 163.367
R557 B.n403 B.n402 163.367
R558 B.n404 B.n403 163.367
R559 B.n404 B.n123 163.367
R560 B.n408 B.n123 163.367
R561 B.n409 B.n408 163.367
R562 B.n410 B.n409 163.367
R563 B.n410 B.n121 163.367
R564 B.n414 B.n121 163.367
R565 B.n415 B.n414 163.367
R566 B.n416 B.n415 163.367
R567 B.n420 B.n119 163.367
R568 B.n421 B.n420 163.367
R569 B.n422 B.n421 163.367
R570 B.n422 B.n117 163.367
R571 B.n426 B.n117 163.367
R572 B.n427 B.n426 163.367
R573 B.n428 B.n427 163.367
R574 B.n428 B.n115 163.367
R575 B.n432 B.n115 163.367
R576 B.n433 B.n432 163.367
R577 B.n434 B.n433 163.367
R578 B.n434 B.n113 163.367
R579 B.n438 B.n113 163.367
R580 B.n439 B.n438 163.367
R581 B.n440 B.n439 163.367
R582 B.n440 B.n111 163.367
R583 B.n444 B.n111 163.367
R584 B.n445 B.n444 163.367
R585 B.n446 B.n445 163.367
R586 B.n446 B.n109 163.367
R587 B.n450 B.n109 163.367
R588 B.n451 B.n450 163.367
R589 B.n452 B.n451 163.367
R590 B.n452 B.n107 163.367
R591 B.n456 B.n107 163.367
R592 B.n457 B.n456 163.367
R593 B.n458 B.n457 163.367
R594 B.n458 B.n105 163.367
R595 B.n462 B.n105 163.367
R596 B.n463 B.n462 163.367
R597 B.n464 B.n463 163.367
R598 B.n464 B.n103 163.367
R599 B.n468 B.n103 163.367
R600 B.n469 B.n468 163.367
R601 B.n470 B.n469 163.367
R602 B.n470 B.n101 163.367
R603 B.n474 B.n101 163.367
R604 B.n475 B.n474 163.367
R605 B.n476 B.n475 163.367
R606 B.n476 B.n99 163.367
R607 B.n480 B.n99 163.367
R608 B.n481 B.n480 163.367
R609 B.n482 B.n481 163.367
R610 B.n482 B.n97 163.367
R611 B.n486 B.n97 163.367
R612 B.n487 B.n486 163.367
R613 B.n488 B.n487 163.367
R614 B.n488 B.n95 163.367
R615 B.n492 B.n95 163.367
R616 B.n493 B.n492 163.367
R617 B.n494 B.n493 163.367
R618 B.n494 B.n93 163.367
R619 B.n498 B.n93 163.367
R620 B.n499 B.n498 163.367
R621 B.n500 B.n499 163.367
R622 B.n500 B.n91 163.367
R623 B.n504 B.n91 163.367
R624 B.n505 B.n504 163.367
R625 B.n506 B.n505 163.367
R626 B.n506 B.n89 163.367
R627 B.n510 B.n89 163.367
R628 B.n511 B.n510 163.367
R629 B.n512 B.n511 163.367
R630 B.n512 B.n87 163.367
R631 B.n516 B.n87 163.367
R632 B.n517 B.n516 163.367
R633 B.n518 B.n517 163.367
R634 B.n518 B.n85 163.367
R635 B.n522 B.n85 163.367
R636 B.n523 B.n522 163.367
R637 B.n524 B.n523 163.367
R638 B.n524 B.n83 163.367
R639 B.n528 B.n83 163.367
R640 B.n529 B.n528 163.367
R641 B.n530 B.n529 163.367
R642 B.n530 B.n81 163.367
R643 B.n534 B.n81 163.367
R644 B.n535 B.n534 163.367
R645 B.n698 B.n697 163.367
R646 B.n697 B.n696 163.367
R647 B.n696 B.n23 163.367
R648 B.n692 B.n23 163.367
R649 B.n692 B.n691 163.367
R650 B.n691 B.n690 163.367
R651 B.n690 B.n25 163.367
R652 B.n686 B.n25 163.367
R653 B.n686 B.n685 163.367
R654 B.n685 B.n684 163.367
R655 B.n684 B.n27 163.367
R656 B.n680 B.n27 163.367
R657 B.n680 B.n679 163.367
R658 B.n679 B.n678 163.367
R659 B.n678 B.n29 163.367
R660 B.n674 B.n29 163.367
R661 B.n674 B.n673 163.367
R662 B.n673 B.n672 163.367
R663 B.n672 B.n31 163.367
R664 B.n668 B.n31 163.367
R665 B.n668 B.n667 163.367
R666 B.n667 B.n666 163.367
R667 B.n666 B.n33 163.367
R668 B.n662 B.n33 163.367
R669 B.n662 B.n661 163.367
R670 B.n661 B.n660 163.367
R671 B.n660 B.n35 163.367
R672 B.n656 B.n35 163.367
R673 B.n656 B.n655 163.367
R674 B.n655 B.n654 163.367
R675 B.n654 B.n37 163.367
R676 B.n650 B.n37 163.367
R677 B.n650 B.n649 163.367
R678 B.n649 B.n648 163.367
R679 B.n648 B.n39 163.367
R680 B.n644 B.n39 163.367
R681 B.n644 B.n643 163.367
R682 B.n643 B.n642 163.367
R683 B.n642 B.n41 163.367
R684 B.n638 B.n41 163.367
R685 B.n638 B.n637 163.367
R686 B.n637 B.n636 163.367
R687 B.n636 B.n43 163.367
R688 B.n632 B.n43 163.367
R689 B.n632 B.n631 163.367
R690 B.n631 B.n630 163.367
R691 B.n630 B.n45 163.367
R692 B.n626 B.n45 163.367
R693 B.n626 B.n625 163.367
R694 B.n625 B.n49 163.367
R695 B.n621 B.n49 163.367
R696 B.n621 B.n620 163.367
R697 B.n620 B.n619 163.367
R698 B.n619 B.n51 163.367
R699 B.n615 B.n51 163.367
R700 B.n615 B.n614 163.367
R701 B.n614 B.n613 163.367
R702 B.n613 B.n53 163.367
R703 B.n608 B.n53 163.367
R704 B.n608 B.n607 163.367
R705 B.n607 B.n606 163.367
R706 B.n606 B.n57 163.367
R707 B.n602 B.n57 163.367
R708 B.n602 B.n601 163.367
R709 B.n601 B.n600 163.367
R710 B.n600 B.n59 163.367
R711 B.n596 B.n59 163.367
R712 B.n596 B.n595 163.367
R713 B.n595 B.n594 163.367
R714 B.n594 B.n61 163.367
R715 B.n590 B.n61 163.367
R716 B.n590 B.n589 163.367
R717 B.n589 B.n588 163.367
R718 B.n588 B.n63 163.367
R719 B.n584 B.n63 163.367
R720 B.n584 B.n583 163.367
R721 B.n583 B.n582 163.367
R722 B.n582 B.n65 163.367
R723 B.n578 B.n65 163.367
R724 B.n578 B.n577 163.367
R725 B.n577 B.n576 163.367
R726 B.n576 B.n67 163.367
R727 B.n572 B.n67 163.367
R728 B.n572 B.n571 163.367
R729 B.n571 B.n570 163.367
R730 B.n570 B.n69 163.367
R731 B.n566 B.n69 163.367
R732 B.n566 B.n565 163.367
R733 B.n565 B.n564 163.367
R734 B.n564 B.n71 163.367
R735 B.n560 B.n71 163.367
R736 B.n560 B.n559 163.367
R737 B.n559 B.n558 163.367
R738 B.n558 B.n73 163.367
R739 B.n554 B.n73 163.367
R740 B.n554 B.n553 163.367
R741 B.n553 B.n552 163.367
R742 B.n552 B.n75 163.367
R743 B.n548 B.n75 163.367
R744 B.n548 B.n547 163.367
R745 B.n547 B.n546 163.367
R746 B.n546 B.n77 163.367
R747 B.n542 B.n77 163.367
R748 B.n542 B.n541 163.367
R749 B.n541 B.n540 163.367
R750 B.n540 B.n79 163.367
R751 B.n536 B.n79 163.367
R752 B.n144 B.t2 163.06
R753 B.n54 B.t10 163.06
R754 B.n152 B.t8 163.042
R755 B.n46 B.t4 163.042
R756 B.n145 B.t1 112.442
R757 B.n55 B.t11 112.442
R758 B.n153 B.t7 112.424
R759 B.n47 B.t5 112.424
R760 B.n146 B.n145 59.5399
R761 B.n328 B.n153 59.5399
R762 B.n48 B.n47 59.5399
R763 B.n610 B.n55 59.5399
R764 B.n145 B.n144 50.6187
R765 B.n153 B.n152 50.6187
R766 B.n47 B.n46 50.6187
R767 B.n55 B.n54 50.6187
R768 B.n700 B.n699 30.4395
R769 B.n418 B.n417 30.4395
R770 B.n255 B.n178 30.4395
R771 B.n537 B.n80 30.4395
R772 B B.n759 18.0485
R773 B.n699 B.n22 10.6151
R774 B.n695 B.n22 10.6151
R775 B.n695 B.n694 10.6151
R776 B.n694 B.n693 10.6151
R777 B.n693 B.n24 10.6151
R778 B.n689 B.n24 10.6151
R779 B.n689 B.n688 10.6151
R780 B.n688 B.n687 10.6151
R781 B.n687 B.n26 10.6151
R782 B.n683 B.n26 10.6151
R783 B.n683 B.n682 10.6151
R784 B.n682 B.n681 10.6151
R785 B.n681 B.n28 10.6151
R786 B.n677 B.n28 10.6151
R787 B.n677 B.n676 10.6151
R788 B.n676 B.n675 10.6151
R789 B.n675 B.n30 10.6151
R790 B.n671 B.n30 10.6151
R791 B.n671 B.n670 10.6151
R792 B.n670 B.n669 10.6151
R793 B.n669 B.n32 10.6151
R794 B.n665 B.n32 10.6151
R795 B.n665 B.n664 10.6151
R796 B.n664 B.n663 10.6151
R797 B.n663 B.n34 10.6151
R798 B.n659 B.n34 10.6151
R799 B.n659 B.n658 10.6151
R800 B.n658 B.n657 10.6151
R801 B.n657 B.n36 10.6151
R802 B.n653 B.n36 10.6151
R803 B.n653 B.n652 10.6151
R804 B.n652 B.n651 10.6151
R805 B.n651 B.n38 10.6151
R806 B.n647 B.n38 10.6151
R807 B.n647 B.n646 10.6151
R808 B.n646 B.n645 10.6151
R809 B.n645 B.n40 10.6151
R810 B.n641 B.n40 10.6151
R811 B.n641 B.n640 10.6151
R812 B.n640 B.n639 10.6151
R813 B.n639 B.n42 10.6151
R814 B.n635 B.n42 10.6151
R815 B.n635 B.n634 10.6151
R816 B.n634 B.n633 10.6151
R817 B.n633 B.n44 10.6151
R818 B.n629 B.n44 10.6151
R819 B.n629 B.n628 10.6151
R820 B.n628 B.n627 10.6151
R821 B.n624 B.n623 10.6151
R822 B.n623 B.n622 10.6151
R823 B.n622 B.n50 10.6151
R824 B.n618 B.n50 10.6151
R825 B.n618 B.n617 10.6151
R826 B.n617 B.n616 10.6151
R827 B.n616 B.n52 10.6151
R828 B.n612 B.n52 10.6151
R829 B.n612 B.n611 10.6151
R830 B.n609 B.n56 10.6151
R831 B.n605 B.n56 10.6151
R832 B.n605 B.n604 10.6151
R833 B.n604 B.n603 10.6151
R834 B.n603 B.n58 10.6151
R835 B.n599 B.n58 10.6151
R836 B.n599 B.n598 10.6151
R837 B.n598 B.n597 10.6151
R838 B.n597 B.n60 10.6151
R839 B.n593 B.n60 10.6151
R840 B.n593 B.n592 10.6151
R841 B.n592 B.n591 10.6151
R842 B.n591 B.n62 10.6151
R843 B.n587 B.n62 10.6151
R844 B.n587 B.n586 10.6151
R845 B.n586 B.n585 10.6151
R846 B.n585 B.n64 10.6151
R847 B.n581 B.n64 10.6151
R848 B.n581 B.n580 10.6151
R849 B.n580 B.n579 10.6151
R850 B.n579 B.n66 10.6151
R851 B.n575 B.n66 10.6151
R852 B.n575 B.n574 10.6151
R853 B.n574 B.n573 10.6151
R854 B.n573 B.n68 10.6151
R855 B.n569 B.n68 10.6151
R856 B.n569 B.n568 10.6151
R857 B.n568 B.n567 10.6151
R858 B.n567 B.n70 10.6151
R859 B.n563 B.n70 10.6151
R860 B.n563 B.n562 10.6151
R861 B.n562 B.n561 10.6151
R862 B.n561 B.n72 10.6151
R863 B.n557 B.n72 10.6151
R864 B.n557 B.n556 10.6151
R865 B.n556 B.n555 10.6151
R866 B.n555 B.n74 10.6151
R867 B.n551 B.n74 10.6151
R868 B.n551 B.n550 10.6151
R869 B.n550 B.n549 10.6151
R870 B.n549 B.n76 10.6151
R871 B.n545 B.n76 10.6151
R872 B.n545 B.n544 10.6151
R873 B.n544 B.n543 10.6151
R874 B.n543 B.n78 10.6151
R875 B.n539 B.n78 10.6151
R876 B.n539 B.n538 10.6151
R877 B.n538 B.n537 10.6151
R878 B.n419 B.n418 10.6151
R879 B.n419 B.n118 10.6151
R880 B.n423 B.n118 10.6151
R881 B.n424 B.n423 10.6151
R882 B.n425 B.n424 10.6151
R883 B.n425 B.n116 10.6151
R884 B.n429 B.n116 10.6151
R885 B.n430 B.n429 10.6151
R886 B.n431 B.n430 10.6151
R887 B.n431 B.n114 10.6151
R888 B.n435 B.n114 10.6151
R889 B.n436 B.n435 10.6151
R890 B.n437 B.n436 10.6151
R891 B.n437 B.n112 10.6151
R892 B.n441 B.n112 10.6151
R893 B.n442 B.n441 10.6151
R894 B.n443 B.n442 10.6151
R895 B.n443 B.n110 10.6151
R896 B.n447 B.n110 10.6151
R897 B.n448 B.n447 10.6151
R898 B.n449 B.n448 10.6151
R899 B.n449 B.n108 10.6151
R900 B.n453 B.n108 10.6151
R901 B.n454 B.n453 10.6151
R902 B.n455 B.n454 10.6151
R903 B.n455 B.n106 10.6151
R904 B.n459 B.n106 10.6151
R905 B.n460 B.n459 10.6151
R906 B.n461 B.n460 10.6151
R907 B.n461 B.n104 10.6151
R908 B.n465 B.n104 10.6151
R909 B.n466 B.n465 10.6151
R910 B.n467 B.n466 10.6151
R911 B.n467 B.n102 10.6151
R912 B.n471 B.n102 10.6151
R913 B.n472 B.n471 10.6151
R914 B.n473 B.n472 10.6151
R915 B.n473 B.n100 10.6151
R916 B.n477 B.n100 10.6151
R917 B.n478 B.n477 10.6151
R918 B.n479 B.n478 10.6151
R919 B.n479 B.n98 10.6151
R920 B.n483 B.n98 10.6151
R921 B.n484 B.n483 10.6151
R922 B.n485 B.n484 10.6151
R923 B.n485 B.n96 10.6151
R924 B.n489 B.n96 10.6151
R925 B.n490 B.n489 10.6151
R926 B.n491 B.n490 10.6151
R927 B.n491 B.n94 10.6151
R928 B.n495 B.n94 10.6151
R929 B.n496 B.n495 10.6151
R930 B.n497 B.n496 10.6151
R931 B.n497 B.n92 10.6151
R932 B.n501 B.n92 10.6151
R933 B.n502 B.n501 10.6151
R934 B.n503 B.n502 10.6151
R935 B.n503 B.n90 10.6151
R936 B.n507 B.n90 10.6151
R937 B.n508 B.n507 10.6151
R938 B.n509 B.n508 10.6151
R939 B.n509 B.n88 10.6151
R940 B.n513 B.n88 10.6151
R941 B.n514 B.n513 10.6151
R942 B.n515 B.n514 10.6151
R943 B.n515 B.n86 10.6151
R944 B.n519 B.n86 10.6151
R945 B.n520 B.n519 10.6151
R946 B.n521 B.n520 10.6151
R947 B.n521 B.n84 10.6151
R948 B.n525 B.n84 10.6151
R949 B.n526 B.n525 10.6151
R950 B.n527 B.n526 10.6151
R951 B.n527 B.n82 10.6151
R952 B.n531 B.n82 10.6151
R953 B.n532 B.n531 10.6151
R954 B.n533 B.n532 10.6151
R955 B.n533 B.n80 10.6151
R956 B.n256 B.n255 10.6151
R957 B.n257 B.n256 10.6151
R958 B.n257 B.n176 10.6151
R959 B.n261 B.n176 10.6151
R960 B.n262 B.n261 10.6151
R961 B.n263 B.n262 10.6151
R962 B.n263 B.n174 10.6151
R963 B.n267 B.n174 10.6151
R964 B.n268 B.n267 10.6151
R965 B.n269 B.n268 10.6151
R966 B.n269 B.n172 10.6151
R967 B.n273 B.n172 10.6151
R968 B.n274 B.n273 10.6151
R969 B.n275 B.n274 10.6151
R970 B.n275 B.n170 10.6151
R971 B.n279 B.n170 10.6151
R972 B.n280 B.n279 10.6151
R973 B.n281 B.n280 10.6151
R974 B.n281 B.n168 10.6151
R975 B.n285 B.n168 10.6151
R976 B.n286 B.n285 10.6151
R977 B.n287 B.n286 10.6151
R978 B.n287 B.n166 10.6151
R979 B.n291 B.n166 10.6151
R980 B.n292 B.n291 10.6151
R981 B.n293 B.n292 10.6151
R982 B.n293 B.n164 10.6151
R983 B.n297 B.n164 10.6151
R984 B.n298 B.n297 10.6151
R985 B.n299 B.n298 10.6151
R986 B.n299 B.n162 10.6151
R987 B.n303 B.n162 10.6151
R988 B.n304 B.n303 10.6151
R989 B.n305 B.n304 10.6151
R990 B.n305 B.n160 10.6151
R991 B.n309 B.n160 10.6151
R992 B.n310 B.n309 10.6151
R993 B.n311 B.n310 10.6151
R994 B.n311 B.n158 10.6151
R995 B.n315 B.n158 10.6151
R996 B.n316 B.n315 10.6151
R997 B.n317 B.n316 10.6151
R998 B.n317 B.n156 10.6151
R999 B.n321 B.n156 10.6151
R1000 B.n322 B.n321 10.6151
R1001 B.n323 B.n322 10.6151
R1002 B.n323 B.n154 10.6151
R1003 B.n327 B.n154 10.6151
R1004 B.n330 B.n329 10.6151
R1005 B.n330 B.n150 10.6151
R1006 B.n334 B.n150 10.6151
R1007 B.n335 B.n334 10.6151
R1008 B.n336 B.n335 10.6151
R1009 B.n336 B.n148 10.6151
R1010 B.n340 B.n148 10.6151
R1011 B.n341 B.n340 10.6151
R1012 B.n342 B.n341 10.6151
R1013 B.n346 B.n345 10.6151
R1014 B.n347 B.n346 10.6151
R1015 B.n347 B.n142 10.6151
R1016 B.n351 B.n142 10.6151
R1017 B.n352 B.n351 10.6151
R1018 B.n353 B.n352 10.6151
R1019 B.n353 B.n140 10.6151
R1020 B.n357 B.n140 10.6151
R1021 B.n358 B.n357 10.6151
R1022 B.n359 B.n358 10.6151
R1023 B.n359 B.n138 10.6151
R1024 B.n363 B.n138 10.6151
R1025 B.n364 B.n363 10.6151
R1026 B.n365 B.n364 10.6151
R1027 B.n365 B.n136 10.6151
R1028 B.n369 B.n136 10.6151
R1029 B.n370 B.n369 10.6151
R1030 B.n371 B.n370 10.6151
R1031 B.n371 B.n134 10.6151
R1032 B.n375 B.n134 10.6151
R1033 B.n376 B.n375 10.6151
R1034 B.n377 B.n376 10.6151
R1035 B.n377 B.n132 10.6151
R1036 B.n381 B.n132 10.6151
R1037 B.n382 B.n381 10.6151
R1038 B.n383 B.n382 10.6151
R1039 B.n383 B.n130 10.6151
R1040 B.n387 B.n130 10.6151
R1041 B.n388 B.n387 10.6151
R1042 B.n389 B.n388 10.6151
R1043 B.n389 B.n128 10.6151
R1044 B.n393 B.n128 10.6151
R1045 B.n394 B.n393 10.6151
R1046 B.n395 B.n394 10.6151
R1047 B.n395 B.n126 10.6151
R1048 B.n399 B.n126 10.6151
R1049 B.n400 B.n399 10.6151
R1050 B.n401 B.n400 10.6151
R1051 B.n401 B.n124 10.6151
R1052 B.n405 B.n124 10.6151
R1053 B.n406 B.n405 10.6151
R1054 B.n407 B.n406 10.6151
R1055 B.n407 B.n122 10.6151
R1056 B.n411 B.n122 10.6151
R1057 B.n412 B.n411 10.6151
R1058 B.n413 B.n412 10.6151
R1059 B.n413 B.n120 10.6151
R1060 B.n417 B.n120 10.6151
R1061 B.n251 B.n178 10.6151
R1062 B.n251 B.n250 10.6151
R1063 B.n250 B.n249 10.6151
R1064 B.n249 B.n180 10.6151
R1065 B.n245 B.n180 10.6151
R1066 B.n245 B.n244 10.6151
R1067 B.n244 B.n243 10.6151
R1068 B.n243 B.n182 10.6151
R1069 B.n239 B.n182 10.6151
R1070 B.n239 B.n238 10.6151
R1071 B.n238 B.n237 10.6151
R1072 B.n237 B.n184 10.6151
R1073 B.n233 B.n184 10.6151
R1074 B.n233 B.n232 10.6151
R1075 B.n232 B.n231 10.6151
R1076 B.n231 B.n186 10.6151
R1077 B.n227 B.n186 10.6151
R1078 B.n227 B.n226 10.6151
R1079 B.n226 B.n225 10.6151
R1080 B.n225 B.n188 10.6151
R1081 B.n221 B.n188 10.6151
R1082 B.n221 B.n220 10.6151
R1083 B.n220 B.n219 10.6151
R1084 B.n219 B.n190 10.6151
R1085 B.n215 B.n190 10.6151
R1086 B.n215 B.n214 10.6151
R1087 B.n214 B.n213 10.6151
R1088 B.n213 B.n192 10.6151
R1089 B.n209 B.n192 10.6151
R1090 B.n209 B.n208 10.6151
R1091 B.n208 B.n207 10.6151
R1092 B.n207 B.n194 10.6151
R1093 B.n203 B.n194 10.6151
R1094 B.n203 B.n202 10.6151
R1095 B.n202 B.n201 10.6151
R1096 B.n201 B.n196 10.6151
R1097 B.n197 B.n196 10.6151
R1098 B.n197 B.n0 10.6151
R1099 B.n755 B.n1 10.6151
R1100 B.n755 B.n754 10.6151
R1101 B.n754 B.n753 10.6151
R1102 B.n753 B.n4 10.6151
R1103 B.n749 B.n4 10.6151
R1104 B.n749 B.n748 10.6151
R1105 B.n748 B.n747 10.6151
R1106 B.n747 B.n6 10.6151
R1107 B.n743 B.n6 10.6151
R1108 B.n743 B.n742 10.6151
R1109 B.n742 B.n741 10.6151
R1110 B.n741 B.n8 10.6151
R1111 B.n737 B.n8 10.6151
R1112 B.n737 B.n736 10.6151
R1113 B.n736 B.n735 10.6151
R1114 B.n735 B.n10 10.6151
R1115 B.n731 B.n10 10.6151
R1116 B.n731 B.n730 10.6151
R1117 B.n730 B.n729 10.6151
R1118 B.n729 B.n12 10.6151
R1119 B.n725 B.n12 10.6151
R1120 B.n725 B.n724 10.6151
R1121 B.n724 B.n723 10.6151
R1122 B.n723 B.n14 10.6151
R1123 B.n719 B.n14 10.6151
R1124 B.n719 B.n718 10.6151
R1125 B.n718 B.n717 10.6151
R1126 B.n717 B.n16 10.6151
R1127 B.n713 B.n16 10.6151
R1128 B.n713 B.n712 10.6151
R1129 B.n712 B.n711 10.6151
R1130 B.n711 B.n18 10.6151
R1131 B.n707 B.n18 10.6151
R1132 B.n707 B.n706 10.6151
R1133 B.n706 B.n705 10.6151
R1134 B.n705 B.n20 10.6151
R1135 B.n701 B.n20 10.6151
R1136 B.n701 B.n700 10.6151
R1137 B.n627 B.n48 9.36635
R1138 B.n610 B.n609 9.36635
R1139 B.n328 B.n327 9.36635
R1140 B.n345 B.n146 9.36635
R1141 B.n759 B.n0 2.81026
R1142 B.n759 B.n1 2.81026
R1143 B.n624 B.n48 1.24928
R1144 B.n611 B.n610 1.24928
R1145 B.n329 B.n328 1.24928
R1146 B.n342 B.n146 1.24928
R1147 VN.n3 VN.t5 187.627
R1148 VN.n17 VN.t1 187.627
R1149 VN.n25 VN.n14 161.3
R1150 VN.n24 VN.n23 161.3
R1151 VN.n22 VN.n15 161.3
R1152 VN.n21 VN.n20 161.3
R1153 VN.n19 VN.n16 161.3
R1154 VN.n11 VN.n0 161.3
R1155 VN.n10 VN.n9 161.3
R1156 VN.n8 VN.n1 161.3
R1157 VN.n7 VN.n6 161.3
R1158 VN.n5 VN.n2 161.3
R1159 VN.n4 VN.t2 154.113
R1160 VN.n12 VN.t4 154.113
R1161 VN.n18 VN.t3 154.113
R1162 VN.n26 VN.t0 154.113
R1163 VN.n13 VN.n12 93.2021
R1164 VN.n27 VN.n26 93.2021
R1165 VN.n4 VN.n3 59.4076
R1166 VN.n18 VN.n17 59.4076
R1167 VN VN.n27 49.7141
R1168 VN.n10 VN.n1 45.9053
R1169 VN.n24 VN.n15 45.9053
R1170 VN.n6 VN.n1 35.2488
R1171 VN.n20 VN.n15 35.2488
R1172 VN.n6 VN.n5 24.5923
R1173 VN.n11 VN.n10 24.5923
R1174 VN.n20 VN.n19 24.5923
R1175 VN.n25 VN.n24 24.5923
R1176 VN.n12 VN.n11 17.7066
R1177 VN.n26 VN.n25 17.7066
R1178 VN.n5 VN.n4 12.2964
R1179 VN.n19 VN.n18 12.2964
R1180 VN.n17 VN.n16 9.18042
R1181 VN.n3 VN.n2 9.18042
R1182 VN.n27 VN.n14 0.278335
R1183 VN.n13 VN.n0 0.278335
R1184 VN.n23 VN.n14 0.189894
R1185 VN.n23 VN.n22 0.189894
R1186 VN.n22 VN.n21 0.189894
R1187 VN.n21 VN.n16 0.189894
R1188 VN.n7 VN.n2 0.189894
R1189 VN.n8 VN.n7 0.189894
R1190 VN.n9 VN.n8 0.189894
R1191 VN.n9 VN.n0 0.189894
R1192 VN VN.n13 0.153485
R1193 VTAIL.n7 VTAIL.t6 55.7229
R1194 VTAIL.n10 VTAIL.t11 55.7229
R1195 VTAIL.n11 VTAIL.t7 55.7227
R1196 VTAIL.n2 VTAIL.t0 55.7227
R1197 VTAIL.n9 VTAIL.n8 53.4935
R1198 VTAIL.n6 VTAIL.n5 53.4935
R1199 VTAIL.n1 VTAIL.n0 53.4934
R1200 VTAIL.n4 VTAIL.n3 53.4934
R1201 VTAIL.n6 VTAIL.n4 29.4358
R1202 VTAIL.n11 VTAIL.n10 27.1858
R1203 VTAIL.n7 VTAIL.n6 2.2505
R1204 VTAIL.n10 VTAIL.n9 2.2505
R1205 VTAIL.n4 VTAIL.n2 2.2505
R1206 VTAIL.n0 VTAIL.t9 2.22992
R1207 VTAIL.n0 VTAIL.t10 2.22992
R1208 VTAIL.n3 VTAIL.t2 2.22992
R1209 VTAIL.n3 VTAIL.t3 2.22992
R1210 VTAIL.n8 VTAIL.t1 2.22992
R1211 VTAIL.n8 VTAIL.t4 2.22992
R1212 VTAIL.n5 VTAIL.t5 2.22992
R1213 VTAIL.n5 VTAIL.t8 2.22992
R1214 VTAIL VTAIL.n11 1.62981
R1215 VTAIL.n9 VTAIL.n7 1.59533
R1216 VTAIL.n2 VTAIL.n1 1.59533
R1217 VTAIL VTAIL.n1 0.62119
R1218 VDD2.n1 VDD2.t0 74.0336
R1219 VDD2.n2 VDD2.t5 72.4017
R1220 VDD2.n1 VDD2.n0 70.6794
R1221 VDD2 VDD2.n3 70.6766
R1222 VDD2.n2 VDD2.n1 43.5968
R1223 VDD2.n3 VDD2.t2 2.22992
R1224 VDD2.n3 VDD2.t4 2.22992
R1225 VDD2.n0 VDD2.t3 2.22992
R1226 VDD2.n0 VDD2.t1 2.22992
R1227 VDD2 VDD2.n2 1.74619
R1228 VP.n9 VP.t4 187.627
R1229 VP.n11 VP.n8 161.3
R1230 VP.n13 VP.n12 161.3
R1231 VP.n14 VP.n7 161.3
R1232 VP.n16 VP.n15 161.3
R1233 VP.n17 VP.n6 161.3
R1234 VP.n36 VP.n0 161.3
R1235 VP.n35 VP.n34 161.3
R1236 VP.n33 VP.n1 161.3
R1237 VP.n32 VP.n31 161.3
R1238 VP.n30 VP.n2 161.3
R1239 VP.n28 VP.n27 161.3
R1240 VP.n26 VP.n3 161.3
R1241 VP.n25 VP.n24 161.3
R1242 VP.n23 VP.n4 161.3
R1243 VP.n22 VP.n21 161.3
R1244 VP.n5 VP.t2 154.113
R1245 VP.n29 VP.t0 154.113
R1246 VP.n37 VP.t5 154.113
R1247 VP.n18 VP.t3 154.113
R1248 VP.n10 VP.t1 154.113
R1249 VP.n20 VP.n5 93.2021
R1250 VP.n38 VP.n37 93.2021
R1251 VP.n19 VP.n18 93.2021
R1252 VP.n10 VP.n9 59.4076
R1253 VP.n20 VP.n19 49.4353
R1254 VP.n24 VP.n23 45.9053
R1255 VP.n35 VP.n1 45.9053
R1256 VP.n16 VP.n7 45.9053
R1257 VP.n24 VP.n3 35.2488
R1258 VP.n31 VP.n1 35.2488
R1259 VP.n12 VP.n7 35.2488
R1260 VP.n23 VP.n22 24.5923
R1261 VP.n28 VP.n3 24.5923
R1262 VP.n31 VP.n30 24.5923
R1263 VP.n36 VP.n35 24.5923
R1264 VP.n17 VP.n16 24.5923
R1265 VP.n12 VP.n11 24.5923
R1266 VP.n22 VP.n5 17.7066
R1267 VP.n37 VP.n36 17.7066
R1268 VP.n18 VP.n17 17.7066
R1269 VP.n29 VP.n28 12.2964
R1270 VP.n30 VP.n29 12.2964
R1271 VP.n11 VP.n10 12.2964
R1272 VP.n9 VP.n8 9.18042
R1273 VP.n19 VP.n6 0.278335
R1274 VP.n21 VP.n20 0.278335
R1275 VP.n38 VP.n0 0.278335
R1276 VP.n13 VP.n8 0.189894
R1277 VP.n14 VP.n13 0.189894
R1278 VP.n15 VP.n14 0.189894
R1279 VP.n15 VP.n6 0.189894
R1280 VP.n21 VP.n4 0.189894
R1281 VP.n25 VP.n4 0.189894
R1282 VP.n26 VP.n25 0.189894
R1283 VP.n27 VP.n26 0.189894
R1284 VP.n27 VP.n2 0.189894
R1285 VP.n32 VP.n2 0.189894
R1286 VP.n33 VP.n32 0.189894
R1287 VP.n34 VP.n33 0.189894
R1288 VP.n34 VP.n0 0.189894
R1289 VP VP.n38 0.153485
R1290 VDD1 VDD1.t1 74.1474
R1291 VDD1.n1 VDD1.t3 74.0336
R1292 VDD1.n1 VDD1.n0 70.6794
R1293 VDD1.n3 VDD1.n2 70.1723
R1294 VDD1.n3 VDD1.n1 45.3048
R1295 VDD1.n2 VDD1.t4 2.22992
R1296 VDD1.n2 VDD1.t2 2.22992
R1297 VDD1.n0 VDD1.t5 2.22992
R1298 VDD1.n0 VDD1.t0 2.22992
R1299 VDD1 VDD1.n3 0.50481
C0 VDD2 VP 0.43164f
C1 w_n3058_n3884# VP 6.15072f
C2 VN VTAIL 7.84884f
C3 VDD2 VTAIL 8.73367f
C4 VN VDD1 0.150509f
C5 VDD2 VDD1 1.28183f
C6 VN B 1.13342f
C7 w_n3058_n3884# VTAIL 3.31096f
C8 VDD2 B 2.27743f
C9 w_n3058_n3884# VDD1 2.39224f
C10 w_n3058_n3884# B 9.957231f
C11 VP VTAIL 7.8632f
C12 VP VDD1 8.155251f
C13 VP B 1.79041f
C14 VTAIL VDD1 8.68604f
C15 B VTAIL 4.12363f
C16 VDD2 VN 7.8779f
C17 B VDD1 2.21101f
C18 w_n3058_n3884# VN 5.75626f
C19 w_n3058_n3884# VDD2 2.46713f
C20 VP VN 7.08766f
C21 VDD2 VSUBS 1.921271f
C22 VDD1 VSUBS 2.37786f
C23 VTAIL VSUBS 1.222125f
C24 VN VSUBS 5.64501f
C25 VP VSUBS 2.784345f
C26 B VSUBS 4.538014f
C27 w_n3058_n3884# VSUBS 0.14572p
C28 VDD1.t1 VSUBS 3.33153f
C29 VDD1.t3 VSUBS 3.33011f
C30 VDD1.t5 VSUBS 0.31684f
C31 VDD1.t0 VSUBS 0.31684f
C32 VDD1.n0 VSUBS 2.54944f
C33 VDD1.n1 VSUBS 3.99467f
C34 VDD1.t4 VSUBS 0.31684f
C35 VDD1.t2 VSUBS 0.31684f
C36 VDD1.n2 VSUBS 2.54372f
C37 VDD1.n3 VSUBS 3.50069f
C38 VP.n0 VSUBS 0.0422f
C39 VP.t5 VSUBS 2.91393f
C40 VP.n1 VSUBS 0.02711f
C41 VP.n2 VSUBS 0.03201f
C42 VP.t0 VSUBS 2.91393f
C43 VP.n3 VSUBS 0.064322f
C44 VP.n4 VSUBS 0.03201f
C45 VP.t2 VSUBS 2.91393f
C46 VP.n5 VSUBS 1.13003f
C47 VP.n6 VSUBS 0.0422f
C48 VP.t3 VSUBS 2.91393f
C49 VP.n7 VSUBS 0.02711f
C50 VP.n8 VSUBS 0.274921f
C51 VP.t1 VSUBS 2.91393f
C52 VP.t4 VSUBS 3.12876f
C53 VP.n9 VSUBS 1.09089f
C54 VP.n10 VSUBS 1.1072f
C55 VP.n11 VSUBS 0.044708f
C56 VP.n12 VSUBS 0.064322f
C57 VP.n13 VSUBS 0.03201f
C58 VP.n14 VSUBS 0.03201f
C59 VP.n15 VSUBS 0.03201f
C60 VP.n16 VSUBS 0.060993f
C61 VP.n17 VSUBS 0.051155f
C62 VP.n18 VSUBS 1.13003f
C63 VP.n19 VSUBS 1.74216f
C64 VP.n20 VSUBS 1.7655f
C65 VP.n21 VSUBS 0.0422f
C66 VP.n22 VSUBS 0.051155f
C67 VP.n23 VSUBS 0.060993f
C68 VP.n24 VSUBS 0.02711f
C69 VP.n25 VSUBS 0.03201f
C70 VP.n26 VSUBS 0.03201f
C71 VP.n27 VSUBS 0.03201f
C72 VP.n28 VSUBS 0.044708f
C73 VP.n29 VSUBS 1.02334f
C74 VP.n30 VSUBS 0.044708f
C75 VP.n31 VSUBS 0.064322f
C76 VP.n32 VSUBS 0.03201f
C77 VP.n33 VSUBS 0.03201f
C78 VP.n34 VSUBS 0.03201f
C79 VP.n35 VSUBS 0.060993f
C80 VP.n36 VSUBS 0.051155f
C81 VP.n37 VSUBS 1.13003f
C82 VP.n38 VSUBS 0.042544f
C83 VDD2.t0 VSUBS 3.33036f
C84 VDD2.t3 VSUBS 0.316863f
C85 VDD2.t1 VSUBS 0.316863f
C86 VDD2.n0 VSUBS 2.54963f
C87 VDD2.n1 VSUBS 3.86563f
C88 VDD2.t5 VSUBS 3.31289f
C89 VDD2.n2 VSUBS 3.53451f
C90 VDD2.t2 VSUBS 0.316863f
C91 VDD2.t4 VSUBS 0.316863f
C92 VDD2.n3 VSUBS 2.54959f
C93 VTAIL.t9 VSUBS 0.323421f
C94 VTAIL.t10 VSUBS 0.323421f
C95 VTAIL.n0 VSUBS 2.42602f
C96 VTAIL.n1 VSUBS 0.88505f
C97 VTAIL.t0 VSUBS 3.18866f
C98 VTAIL.n2 VSUBS 1.15184f
C99 VTAIL.t2 VSUBS 0.323421f
C100 VTAIL.t3 VSUBS 0.323421f
C101 VTAIL.n3 VSUBS 2.42602f
C102 VTAIL.n4 VSUBS 2.81339f
C103 VTAIL.t5 VSUBS 0.323421f
C104 VTAIL.t8 VSUBS 0.323421f
C105 VTAIL.n5 VSUBS 2.42603f
C106 VTAIL.n6 VSUBS 2.81338f
C107 VTAIL.t6 VSUBS 3.18867f
C108 VTAIL.n7 VSUBS 1.15183f
C109 VTAIL.t1 VSUBS 0.323421f
C110 VTAIL.t4 VSUBS 0.323421f
C111 VTAIL.n8 VSUBS 2.42603f
C112 VTAIL.n9 VSUBS 1.03242f
C113 VTAIL.t11 VSUBS 3.18868f
C114 VTAIL.n10 VSUBS 2.72927f
C115 VTAIL.t7 VSUBS 3.18866f
C116 VTAIL.n11 VSUBS 2.67315f
C117 VN.n0 VSUBS 0.040989f
C118 VN.t4 VSUBS 2.83031f
C119 VN.n1 VSUBS 0.026332f
C120 VN.n2 VSUBS 0.267031f
C121 VN.t2 VSUBS 2.83031f
C122 VN.t5 VSUBS 3.03898f
C123 VN.n3 VSUBS 1.05958f
C124 VN.n4 VSUBS 1.07543f
C125 VN.n5 VSUBS 0.043425f
C126 VN.n6 VSUBS 0.062476f
C127 VN.n7 VSUBS 0.031092f
C128 VN.n8 VSUBS 0.031092f
C129 VN.n9 VSUBS 0.031092f
C130 VN.n10 VSUBS 0.059243f
C131 VN.n11 VSUBS 0.049687f
C132 VN.n12 VSUBS 1.0976f
C133 VN.n13 VSUBS 0.041323f
C134 VN.n14 VSUBS 0.040989f
C135 VN.t0 VSUBS 2.83031f
C136 VN.n15 VSUBS 0.026332f
C137 VN.n16 VSUBS 0.267031f
C138 VN.t3 VSUBS 2.83031f
C139 VN.t1 VSUBS 3.03898f
C140 VN.n17 VSUBS 1.05958f
C141 VN.n18 VSUBS 1.07543f
C142 VN.n19 VSUBS 0.043425f
C143 VN.n20 VSUBS 0.062476f
C144 VN.n21 VSUBS 0.031092f
C145 VN.n22 VSUBS 0.031092f
C146 VN.n23 VSUBS 0.031092f
C147 VN.n24 VSUBS 0.059243f
C148 VN.n25 VSUBS 0.049687f
C149 VN.n26 VSUBS 1.0976f
C150 VN.n27 VSUBS 1.7089f
C151 B.n0 VSUBS 0.004953f
C152 B.n1 VSUBS 0.004953f
C153 B.n2 VSUBS 0.007833f
C154 B.n3 VSUBS 0.007833f
C155 B.n4 VSUBS 0.007833f
C156 B.n5 VSUBS 0.007833f
C157 B.n6 VSUBS 0.007833f
C158 B.n7 VSUBS 0.007833f
C159 B.n8 VSUBS 0.007833f
C160 B.n9 VSUBS 0.007833f
C161 B.n10 VSUBS 0.007833f
C162 B.n11 VSUBS 0.007833f
C163 B.n12 VSUBS 0.007833f
C164 B.n13 VSUBS 0.007833f
C165 B.n14 VSUBS 0.007833f
C166 B.n15 VSUBS 0.007833f
C167 B.n16 VSUBS 0.007833f
C168 B.n17 VSUBS 0.007833f
C169 B.n18 VSUBS 0.007833f
C170 B.n19 VSUBS 0.007833f
C171 B.n20 VSUBS 0.007833f
C172 B.n21 VSUBS 0.017182f
C173 B.n22 VSUBS 0.007833f
C174 B.n23 VSUBS 0.007833f
C175 B.n24 VSUBS 0.007833f
C176 B.n25 VSUBS 0.007833f
C177 B.n26 VSUBS 0.007833f
C178 B.n27 VSUBS 0.007833f
C179 B.n28 VSUBS 0.007833f
C180 B.n29 VSUBS 0.007833f
C181 B.n30 VSUBS 0.007833f
C182 B.n31 VSUBS 0.007833f
C183 B.n32 VSUBS 0.007833f
C184 B.n33 VSUBS 0.007833f
C185 B.n34 VSUBS 0.007833f
C186 B.n35 VSUBS 0.007833f
C187 B.n36 VSUBS 0.007833f
C188 B.n37 VSUBS 0.007833f
C189 B.n38 VSUBS 0.007833f
C190 B.n39 VSUBS 0.007833f
C191 B.n40 VSUBS 0.007833f
C192 B.n41 VSUBS 0.007833f
C193 B.n42 VSUBS 0.007833f
C194 B.n43 VSUBS 0.007833f
C195 B.n44 VSUBS 0.007833f
C196 B.n45 VSUBS 0.007833f
C197 B.t5 VSUBS 0.541821f
C198 B.t4 VSUBS 0.562886f
C199 B.t3 VSUBS 1.65751f
C200 B.n46 VSUBS 0.287528f
C201 B.n47 VSUBS 0.07902f
C202 B.n48 VSUBS 0.018148f
C203 B.n49 VSUBS 0.007833f
C204 B.n50 VSUBS 0.007833f
C205 B.n51 VSUBS 0.007833f
C206 B.n52 VSUBS 0.007833f
C207 B.n53 VSUBS 0.007833f
C208 B.t11 VSUBS 0.541807f
C209 B.t10 VSUBS 0.562874f
C210 B.t9 VSUBS 1.65751f
C211 B.n54 VSUBS 0.28754f
C212 B.n55 VSUBS 0.079034f
C213 B.n56 VSUBS 0.007833f
C214 B.n57 VSUBS 0.007833f
C215 B.n58 VSUBS 0.007833f
C216 B.n59 VSUBS 0.007833f
C217 B.n60 VSUBS 0.007833f
C218 B.n61 VSUBS 0.007833f
C219 B.n62 VSUBS 0.007833f
C220 B.n63 VSUBS 0.007833f
C221 B.n64 VSUBS 0.007833f
C222 B.n65 VSUBS 0.007833f
C223 B.n66 VSUBS 0.007833f
C224 B.n67 VSUBS 0.007833f
C225 B.n68 VSUBS 0.007833f
C226 B.n69 VSUBS 0.007833f
C227 B.n70 VSUBS 0.007833f
C228 B.n71 VSUBS 0.007833f
C229 B.n72 VSUBS 0.007833f
C230 B.n73 VSUBS 0.007833f
C231 B.n74 VSUBS 0.007833f
C232 B.n75 VSUBS 0.007833f
C233 B.n76 VSUBS 0.007833f
C234 B.n77 VSUBS 0.007833f
C235 B.n78 VSUBS 0.007833f
C236 B.n79 VSUBS 0.007833f
C237 B.n80 VSUBS 0.018175f
C238 B.n81 VSUBS 0.007833f
C239 B.n82 VSUBS 0.007833f
C240 B.n83 VSUBS 0.007833f
C241 B.n84 VSUBS 0.007833f
C242 B.n85 VSUBS 0.007833f
C243 B.n86 VSUBS 0.007833f
C244 B.n87 VSUBS 0.007833f
C245 B.n88 VSUBS 0.007833f
C246 B.n89 VSUBS 0.007833f
C247 B.n90 VSUBS 0.007833f
C248 B.n91 VSUBS 0.007833f
C249 B.n92 VSUBS 0.007833f
C250 B.n93 VSUBS 0.007833f
C251 B.n94 VSUBS 0.007833f
C252 B.n95 VSUBS 0.007833f
C253 B.n96 VSUBS 0.007833f
C254 B.n97 VSUBS 0.007833f
C255 B.n98 VSUBS 0.007833f
C256 B.n99 VSUBS 0.007833f
C257 B.n100 VSUBS 0.007833f
C258 B.n101 VSUBS 0.007833f
C259 B.n102 VSUBS 0.007833f
C260 B.n103 VSUBS 0.007833f
C261 B.n104 VSUBS 0.007833f
C262 B.n105 VSUBS 0.007833f
C263 B.n106 VSUBS 0.007833f
C264 B.n107 VSUBS 0.007833f
C265 B.n108 VSUBS 0.007833f
C266 B.n109 VSUBS 0.007833f
C267 B.n110 VSUBS 0.007833f
C268 B.n111 VSUBS 0.007833f
C269 B.n112 VSUBS 0.007833f
C270 B.n113 VSUBS 0.007833f
C271 B.n114 VSUBS 0.007833f
C272 B.n115 VSUBS 0.007833f
C273 B.n116 VSUBS 0.007833f
C274 B.n117 VSUBS 0.007833f
C275 B.n118 VSUBS 0.007833f
C276 B.n119 VSUBS 0.017182f
C277 B.n120 VSUBS 0.007833f
C278 B.n121 VSUBS 0.007833f
C279 B.n122 VSUBS 0.007833f
C280 B.n123 VSUBS 0.007833f
C281 B.n124 VSUBS 0.007833f
C282 B.n125 VSUBS 0.007833f
C283 B.n126 VSUBS 0.007833f
C284 B.n127 VSUBS 0.007833f
C285 B.n128 VSUBS 0.007833f
C286 B.n129 VSUBS 0.007833f
C287 B.n130 VSUBS 0.007833f
C288 B.n131 VSUBS 0.007833f
C289 B.n132 VSUBS 0.007833f
C290 B.n133 VSUBS 0.007833f
C291 B.n134 VSUBS 0.007833f
C292 B.n135 VSUBS 0.007833f
C293 B.n136 VSUBS 0.007833f
C294 B.n137 VSUBS 0.007833f
C295 B.n138 VSUBS 0.007833f
C296 B.n139 VSUBS 0.007833f
C297 B.n140 VSUBS 0.007833f
C298 B.n141 VSUBS 0.007833f
C299 B.n142 VSUBS 0.007833f
C300 B.n143 VSUBS 0.007833f
C301 B.t1 VSUBS 0.541807f
C302 B.t2 VSUBS 0.562874f
C303 B.t0 VSUBS 1.65751f
C304 B.n144 VSUBS 0.28754f
C305 B.n145 VSUBS 0.079034f
C306 B.n146 VSUBS 0.018148f
C307 B.n147 VSUBS 0.007833f
C308 B.n148 VSUBS 0.007833f
C309 B.n149 VSUBS 0.007833f
C310 B.n150 VSUBS 0.007833f
C311 B.n151 VSUBS 0.007833f
C312 B.t7 VSUBS 0.541821f
C313 B.t8 VSUBS 0.562886f
C314 B.t6 VSUBS 1.65751f
C315 B.n152 VSUBS 0.287528f
C316 B.n153 VSUBS 0.07902f
C317 B.n154 VSUBS 0.007833f
C318 B.n155 VSUBS 0.007833f
C319 B.n156 VSUBS 0.007833f
C320 B.n157 VSUBS 0.007833f
C321 B.n158 VSUBS 0.007833f
C322 B.n159 VSUBS 0.007833f
C323 B.n160 VSUBS 0.007833f
C324 B.n161 VSUBS 0.007833f
C325 B.n162 VSUBS 0.007833f
C326 B.n163 VSUBS 0.007833f
C327 B.n164 VSUBS 0.007833f
C328 B.n165 VSUBS 0.007833f
C329 B.n166 VSUBS 0.007833f
C330 B.n167 VSUBS 0.007833f
C331 B.n168 VSUBS 0.007833f
C332 B.n169 VSUBS 0.007833f
C333 B.n170 VSUBS 0.007833f
C334 B.n171 VSUBS 0.007833f
C335 B.n172 VSUBS 0.007833f
C336 B.n173 VSUBS 0.007833f
C337 B.n174 VSUBS 0.007833f
C338 B.n175 VSUBS 0.007833f
C339 B.n176 VSUBS 0.007833f
C340 B.n177 VSUBS 0.007833f
C341 B.n178 VSUBS 0.017182f
C342 B.n179 VSUBS 0.007833f
C343 B.n180 VSUBS 0.007833f
C344 B.n181 VSUBS 0.007833f
C345 B.n182 VSUBS 0.007833f
C346 B.n183 VSUBS 0.007833f
C347 B.n184 VSUBS 0.007833f
C348 B.n185 VSUBS 0.007833f
C349 B.n186 VSUBS 0.007833f
C350 B.n187 VSUBS 0.007833f
C351 B.n188 VSUBS 0.007833f
C352 B.n189 VSUBS 0.007833f
C353 B.n190 VSUBS 0.007833f
C354 B.n191 VSUBS 0.007833f
C355 B.n192 VSUBS 0.007833f
C356 B.n193 VSUBS 0.007833f
C357 B.n194 VSUBS 0.007833f
C358 B.n195 VSUBS 0.007833f
C359 B.n196 VSUBS 0.007833f
C360 B.n197 VSUBS 0.007833f
C361 B.n198 VSUBS 0.007833f
C362 B.n199 VSUBS 0.007833f
C363 B.n200 VSUBS 0.007833f
C364 B.n201 VSUBS 0.007833f
C365 B.n202 VSUBS 0.007833f
C366 B.n203 VSUBS 0.007833f
C367 B.n204 VSUBS 0.007833f
C368 B.n205 VSUBS 0.007833f
C369 B.n206 VSUBS 0.007833f
C370 B.n207 VSUBS 0.007833f
C371 B.n208 VSUBS 0.007833f
C372 B.n209 VSUBS 0.007833f
C373 B.n210 VSUBS 0.007833f
C374 B.n211 VSUBS 0.007833f
C375 B.n212 VSUBS 0.007833f
C376 B.n213 VSUBS 0.007833f
C377 B.n214 VSUBS 0.007833f
C378 B.n215 VSUBS 0.007833f
C379 B.n216 VSUBS 0.007833f
C380 B.n217 VSUBS 0.007833f
C381 B.n218 VSUBS 0.007833f
C382 B.n219 VSUBS 0.007833f
C383 B.n220 VSUBS 0.007833f
C384 B.n221 VSUBS 0.007833f
C385 B.n222 VSUBS 0.007833f
C386 B.n223 VSUBS 0.007833f
C387 B.n224 VSUBS 0.007833f
C388 B.n225 VSUBS 0.007833f
C389 B.n226 VSUBS 0.007833f
C390 B.n227 VSUBS 0.007833f
C391 B.n228 VSUBS 0.007833f
C392 B.n229 VSUBS 0.007833f
C393 B.n230 VSUBS 0.007833f
C394 B.n231 VSUBS 0.007833f
C395 B.n232 VSUBS 0.007833f
C396 B.n233 VSUBS 0.007833f
C397 B.n234 VSUBS 0.007833f
C398 B.n235 VSUBS 0.007833f
C399 B.n236 VSUBS 0.007833f
C400 B.n237 VSUBS 0.007833f
C401 B.n238 VSUBS 0.007833f
C402 B.n239 VSUBS 0.007833f
C403 B.n240 VSUBS 0.007833f
C404 B.n241 VSUBS 0.007833f
C405 B.n242 VSUBS 0.007833f
C406 B.n243 VSUBS 0.007833f
C407 B.n244 VSUBS 0.007833f
C408 B.n245 VSUBS 0.007833f
C409 B.n246 VSUBS 0.007833f
C410 B.n247 VSUBS 0.007833f
C411 B.n248 VSUBS 0.007833f
C412 B.n249 VSUBS 0.007833f
C413 B.n250 VSUBS 0.007833f
C414 B.n251 VSUBS 0.007833f
C415 B.n252 VSUBS 0.007833f
C416 B.n253 VSUBS 0.017182f
C417 B.n254 VSUBS 0.017836f
C418 B.n255 VSUBS 0.017836f
C419 B.n256 VSUBS 0.007833f
C420 B.n257 VSUBS 0.007833f
C421 B.n258 VSUBS 0.007833f
C422 B.n259 VSUBS 0.007833f
C423 B.n260 VSUBS 0.007833f
C424 B.n261 VSUBS 0.007833f
C425 B.n262 VSUBS 0.007833f
C426 B.n263 VSUBS 0.007833f
C427 B.n264 VSUBS 0.007833f
C428 B.n265 VSUBS 0.007833f
C429 B.n266 VSUBS 0.007833f
C430 B.n267 VSUBS 0.007833f
C431 B.n268 VSUBS 0.007833f
C432 B.n269 VSUBS 0.007833f
C433 B.n270 VSUBS 0.007833f
C434 B.n271 VSUBS 0.007833f
C435 B.n272 VSUBS 0.007833f
C436 B.n273 VSUBS 0.007833f
C437 B.n274 VSUBS 0.007833f
C438 B.n275 VSUBS 0.007833f
C439 B.n276 VSUBS 0.007833f
C440 B.n277 VSUBS 0.007833f
C441 B.n278 VSUBS 0.007833f
C442 B.n279 VSUBS 0.007833f
C443 B.n280 VSUBS 0.007833f
C444 B.n281 VSUBS 0.007833f
C445 B.n282 VSUBS 0.007833f
C446 B.n283 VSUBS 0.007833f
C447 B.n284 VSUBS 0.007833f
C448 B.n285 VSUBS 0.007833f
C449 B.n286 VSUBS 0.007833f
C450 B.n287 VSUBS 0.007833f
C451 B.n288 VSUBS 0.007833f
C452 B.n289 VSUBS 0.007833f
C453 B.n290 VSUBS 0.007833f
C454 B.n291 VSUBS 0.007833f
C455 B.n292 VSUBS 0.007833f
C456 B.n293 VSUBS 0.007833f
C457 B.n294 VSUBS 0.007833f
C458 B.n295 VSUBS 0.007833f
C459 B.n296 VSUBS 0.007833f
C460 B.n297 VSUBS 0.007833f
C461 B.n298 VSUBS 0.007833f
C462 B.n299 VSUBS 0.007833f
C463 B.n300 VSUBS 0.007833f
C464 B.n301 VSUBS 0.007833f
C465 B.n302 VSUBS 0.007833f
C466 B.n303 VSUBS 0.007833f
C467 B.n304 VSUBS 0.007833f
C468 B.n305 VSUBS 0.007833f
C469 B.n306 VSUBS 0.007833f
C470 B.n307 VSUBS 0.007833f
C471 B.n308 VSUBS 0.007833f
C472 B.n309 VSUBS 0.007833f
C473 B.n310 VSUBS 0.007833f
C474 B.n311 VSUBS 0.007833f
C475 B.n312 VSUBS 0.007833f
C476 B.n313 VSUBS 0.007833f
C477 B.n314 VSUBS 0.007833f
C478 B.n315 VSUBS 0.007833f
C479 B.n316 VSUBS 0.007833f
C480 B.n317 VSUBS 0.007833f
C481 B.n318 VSUBS 0.007833f
C482 B.n319 VSUBS 0.007833f
C483 B.n320 VSUBS 0.007833f
C484 B.n321 VSUBS 0.007833f
C485 B.n322 VSUBS 0.007833f
C486 B.n323 VSUBS 0.007833f
C487 B.n324 VSUBS 0.007833f
C488 B.n325 VSUBS 0.007833f
C489 B.n326 VSUBS 0.007833f
C490 B.n327 VSUBS 0.007372f
C491 B.n328 VSUBS 0.018148f
C492 B.n329 VSUBS 0.004377f
C493 B.n330 VSUBS 0.007833f
C494 B.n331 VSUBS 0.007833f
C495 B.n332 VSUBS 0.007833f
C496 B.n333 VSUBS 0.007833f
C497 B.n334 VSUBS 0.007833f
C498 B.n335 VSUBS 0.007833f
C499 B.n336 VSUBS 0.007833f
C500 B.n337 VSUBS 0.007833f
C501 B.n338 VSUBS 0.007833f
C502 B.n339 VSUBS 0.007833f
C503 B.n340 VSUBS 0.007833f
C504 B.n341 VSUBS 0.007833f
C505 B.n342 VSUBS 0.004377f
C506 B.n343 VSUBS 0.007833f
C507 B.n344 VSUBS 0.007833f
C508 B.n345 VSUBS 0.007372f
C509 B.n346 VSUBS 0.007833f
C510 B.n347 VSUBS 0.007833f
C511 B.n348 VSUBS 0.007833f
C512 B.n349 VSUBS 0.007833f
C513 B.n350 VSUBS 0.007833f
C514 B.n351 VSUBS 0.007833f
C515 B.n352 VSUBS 0.007833f
C516 B.n353 VSUBS 0.007833f
C517 B.n354 VSUBS 0.007833f
C518 B.n355 VSUBS 0.007833f
C519 B.n356 VSUBS 0.007833f
C520 B.n357 VSUBS 0.007833f
C521 B.n358 VSUBS 0.007833f
C522 B.n359 VSUBS 0.007833f
C523 B.n360 VSUBS 0.007833f
C524 B.n361 VSUBS 0.007833f
C525 B.n362 VSUBS 0.007833f
C526 B.n363 VSUBS 0.007833f
C527 B.n364 VSUBS 0.007833f
C528 B.n365 VSUBS 0.007833f
C529 B.n366 VSUBS 0.007833f
C530 B.n367 VSUBS 0.007833f
C531 B.n368 VSUBS 0.007833f
C532 B.n369 VSUBS 0.007833f
C533 B.n370 VSUBS 0.007833f
C534 B.n371 VSUBS 0.007833f
C535 B.n372 VSUBS 0.007833f
C536 B.n373 VSUBS 0.007833f
C537 B.n374 VSUBS 0.007833f
C538 B.n375 VSUBS 0.007833f
C539 B.n376 VSUBS 0.007833f
C540 B.n377 VSUBS 0.007833f
C541 B.n378 VSUBS 0.007833f
C542 B.n379 VSUBS 0.007833f
C543 B.n380 VSUBS 0.007833f
C544 B.n381 VSUBS 0.007833f
C545 B.n382 VSUBS 0.007833f
C546 B.n383 VSUBS 0.007833f
C547 B.n384 VSUBS 0.007833f
C548 B.n385 VSUBS 0.007833f
C549 B.n386 VSUBS 0.007833f
C550 B.n387 VSUBS 0.007833f
C551 B.n388 VSUBS 0.007833f
C552 B.n389 VSUBS 0.007833f
C553 B.n390 VSUBS 0.007833f
C554 B.n391 VSUBS 0.007833f
C555 B.n392 VSUBS 0.007833f
C556 B.n393 VSUBS 0.007833f
C557 B.n394 VSUBS 0.007833f
C558 B.n395 VSUBS 0.007833f
C559 B.n396 VSUBS 0.007833f
C560 B.n397 VSUBS 0.007833f
C561 B.n398 VSUBS 0.007833f
C562 B.n399 VSUBS 0.007833f
C563 B.n400 VSUBS 0.007833f
C564 B.n401 VSUBS 0.007833f
C565 B.n402 VSUBS 0.007833f
C566 B.n403 VSUBS 0.007833f
C567 B.n404 VSUBS 0.007833f
C568 B.n405 VSUBS 0.007833f
C569 B.n406 VSUBS 0.007833f
C570 B.n407 VSUBS 0.007833f
C571 B.n408 VSUBS 0.007833f
C572 B.n409 VSUBS 0.007833f
C573 B.n410 VSUBS 0.007833f
C574 B.n411 VSUBS 0.007833f
C575 B.n412 VSUBS 0.007833f
C576 B.n413 VSUBS 0.007833f
C577 B.n414 VSUBS 0.007833f
C578 B.n415 VSUBS 0.007833f
C579 B.n416 VSUBS 0.017836f
C580 B.n417 VSUBS 0.017836f
C581 B.n418 VSUBS 0.017182f
C582 B.n419 VSUBS 0.007833f
C583 B.n420 VSUBS 0.007833f
C584 B.n421 VSUBS 0.007833f
C585 B.n422 VSUBS 0.007833f
C586 B.n423 VSUBS 0.007833f
C587 B.n424 VSUBS 0.007833f
C588 B.n425 VSUBS 0.007833f
C589 B.n426 VSUBS 0.007833f
C590 B.n427 VSUBS 0.007833f
C591 B.n428 VSUBS 0.007833f
C592 B.n429 VSUBS 0.007833f
C593 B.n430 VSUBS 0.007833f
C594 B.n431 VSUBS 0.007833f
C595 B.n432 VSUBS 0.007833f
C596 B.n433 VSUBS 0.007833f
C597 B.n434 VSUBS 0.007833f
C598 B.n435 VSUBS 0.007833f
C599 B.n436 VSUBS 0.007833f
C600 B.n437 VSUBS 0.007833f
C601 B.n438 VSUBS 0.007833f
C602 B.n439 VSUBS 0.007833f
C603 B.n440 VSUBS 0.007833f
C604 B.n441 VSUBS 0.007833f
C605 B.n442 VSUBS 0.007833f
C606 B.n443 VSUBS 0.007833f
C607 B.n444 VSUBS 0.007833f
C608 B.n445 VSUBS 0.007833f
C609 B.n446 VSUBS 0.007833f
C610 B.n447 VSUBS 0.007833f
C611 B.n448 VSUBS 0.007833f
C612 B.n449 VSUBS 0.007833f
C613 B.n450 VSUBS 0.007833f
C614 B.n451 VSUBS 0.007833f
C615 B.n452 VSUBS 0.007833f
C616 B.n453 VSUBS 0.007833f
C617 B.n454 VSUBS 0.007833f
C618 B.n455 VSUBS 0.007833f
C619 B.n456 VSUBS 0.007833f
C620 B.n457 VSUBS 0.007833f
C621 B.n458 VSUBS 0.007833f
C622 B.n459 VSUBS 0.007833f
C623 B.n460 VSUBS 0.007833f
C624 B.n461 VSUBS 0.007833f
C625 B.n462 VSUBS 0.007833f
C626 B.n463 VSUBS 0.007833f
C627 B.n464 VSUBS 0.007833f
C628 B.n465 VSUBS 0.007833f
C629 B.n466 VSUBS 0.007833f
C630 B.n467 VSUBS 0.007833f
C631 B.n468 VSUBS 0.007833f
C632 B.n469 VSUBS 0.007833f
C633 B.n470 VSUBS 0.007833f
C634 B.n471 VSUBS 0.007833f
C635 B.n472 VSUBS 0.007833f
C636 B.n473 VSUBS 0.007833f
C637 B.n474 VSUBS 0.007833f
C638 B.n475 VSUBS 0.007833f
C639 B.n476 VSUBS 0.007833f
C640 B.n477 VSUBS 0.007833f
C641 B.n478 VSUBS 0.007833f
C642 B.n479 VSUBS 0.007833f
C643 B.n480 VSUBS 0.007833f
C644 B.n481 VSUBS 0.007833f
C645 B.n482 VSUBS 0.007833f
C646 B.n483 VSUBS 0.007833f
C647 B.n484 VSUBS 0.007833f
C648 B.n485 VSUBS 0.007833f
C649 B.n486 VSUBS 0.007833f
C650 B.n487 VSUBS 0.007833f
C651 B.n488 VSUBS 0.007833f
C652 B.n489 VSUBS 0.007833f
C653 B.n490 VSUBS 0.007833f
C654 B.n491 VSUBS 0.007833f
C655 B.n492 VSUBS 0.007833f
C656 B.n493 VSUBS 0.007833f
C657 B.n494 VSUBS 0.007833f
C658 B.n495 VSUBS 0.007833f
C659 B.n496 VSUBS 0.007833f
C660 B.n497 VSUBS 0.007833f
C661 B.n498 VSUBS 0.007833f
C662 B.n499 VSUBS 0.007833f
C663 B.n500 VSUBS 0.007833f
C664 B.n501 VSUBS 0.007833f
C665 B.n502 VSUBS 0.007833f
C666 B.n503 VSUBS 0.007833f
C667 B.n504 VSUBS 0.007833f
C668 B.n505 VSUBS 0.007833f
C669 B.n506 VSUBS 0.007833f
C670 B.n507 VSUBS 0.007833f
C671 B.n508 VSUBS 0.007833f
C672 B.n509 VSUBS 0.007833f
C673 B.n510 VSUBS 0.007833f
C674 B.n511 VSUBS 0.007833f
C675 B.n512 VSUBS 0.007833f
C676 B.n513 VSUBS 0.007833f
C677 B.n514 VSUBS 0.007833f
C678 B.n515 VSUBS 0.007833f
C679 B.n516 VSUBS 0.007833f
C680 B.n517 VSUBS 0.007833f
C681 B.n518 VSUBS 0.007833f
C682 B.n519 VSUBS 0.007833f
C683 B.n520 VSUBS 0.007833f
C684 B.n521 VSUBS 0.007833f
C685 B.n522 VSUBS 0.007833f
C686 B.n523 VSUBS 0.007833f
C687 B.n524 VSUBS 0.007833f
C688 B.n525 VSUBS 0.007833f
C689 B.n526 VSUBS 0.007833f
C690 B.n527 VSUBS 0.007833f
C691 B.n528 VSUBS 0.007833f
C692 B.n529 VSUBS 0.007833f
C693 B.n530 VSUBS 0.007833f
C694 B.n531 VSUBS 0.007833f
C695 B.n532 VSUBS 0.007833f
C696 B.n533 VSUBS 0.007833f
C697 B.n534 VSUBS 0.007833f
C698 B.n535 VSUBS 0.017182f
C699 B.n536 VSUBS 0.017836f
C700 B.n537 VSUBS 0.016843f
C701 B.n538 VSUBS 0.007833f
C702 B.n539 VSUBS 0.007833f
C703 B.n540 VSUBS 0.007833f
C704 B.n541 VSUBS 0.007833f
C705 B.n542 VSUBS 0.007833f
C706 B.n543 VSUBS 0.007833f
C707 B.n544 VSUBS 0.007833f
C708 B.n545 VSUBS 0.007833f
C709 B.n546 VSUBS 0.007833f
C710 B.n547 VSUBS 0.007833f
C711 B.n548 VSUBS 0.007833f
C712 B.n549 VSUBS 0.007833f
C713 B.n550 VSUBS 0.007833f
C714 B.n551 VSUBS 0.007833f
C715 B.n552 VSUBS 0.007833f
C716 B.n553 VSUBS 0.007833f
C717 B.n554 VSUBS 0.007833f
C718 B.n555 VSUBS 0.007833f
C719 B.n556 VSUBS 0.007833f
C720 B.n557 VSUBS 0.007833f
C721 B.n558 VSUBS 0.007833f
C722 B.n559 VSUBS 0.007833f
C723 B.n560 VSUBS 0.007833f
C724 B.n561 VSUBS 0.007833f
C725 B.n562 VSUBS 0.007833f
C726 B.n563 VSUBS 0.007833f
C727 B.n564 VSUBS 0.007833f
C728 B.n565 VSUBS 0.007833f
C729 B.n566 VSUBS 0.007833f
C730 B.n567 VSUBS 0.007833f
C731 B.n568 VSUBS 0.007833f
C732 B.n569 VSUBS 0.007833f
C733 B.n570 VSUBS 0.007833f
C734 B.n571 VSUBS 0.007833f
C735 B.n572 VSUBS 0.007833f
C736 B.n573 VSUBS 0.007833f
C737 B.n574 VSUBS 0.007833f
C738 B.n575 VSUBS 0.007833f
C739 B.n576 VSUBS 0.007833f
C740 B.n577 VSUBS 0.007833f
C741 B.n578 VSUBS 0.007833f
C742 B.n579 VSUBS 0.007833f
C743 B.n580 VSUBS 0.007833f
C744 B.n581 VSUBS 0.007833f
C745 B.n582 VSUBS 0.007833f
C746 B.n583 VSUBS 0.007833f
C747 B.n584 VSUBS 0.007833f
C748 B.n585 VSUBS 0.007833f
C749 B.n586 VSUBS 0.007833f
C750 B.n587 VSUBS 0.007833f
C751 B.n588 VSUBS 0.007833f
C752 B.n589 VSUBS 0.007833f
C753 B.n590 VSUBS 0.007833f
C754 B.n591 VSUBS 0.007833f
C755 B.n592 VSUBS 0.007833f
C756 B.n593 VSUBS 0.007833f
C757 B.n594 VSUBS 0.007833f
C758 B.n595 VSUBS 0.007833f
C759 B.n596 VSUBS 0.007833f
C760 B.n597 VSUBS 0.007833f
C761 B.n598 VSUBS 0.007833f
C762 B.n599 VSUBS 0.007833f
C763 B.n600 VSUBS 0.007833f
C764 B.n601 VSUBS 0.007833f
C765 B.n602 VSUBS 0.007833f
C766 B.n603 VSUBS 0.007833f
C767 B.n604 VSUBS 0.007833f
C768 B.n605 VSUBS 0.007833f
C769 B.n606 VSUBS 0.007833f
C770 B.n607 VSUBS 0.007833f
C771 B.n608 VSUBS 0.007833f
C772 B.n609 VSUBS 0.007372f
C773 B.n610 VSUBS 0.018148f
C774 B.n611 VSUBS 0.004377f
C775 B.n612 VSUBS 0.007833f
C776 B.n613 VSUBS 0.007833f
C777 B.n614 VSUBS 0.007833f
C778 B.n615 VSUBS 0.007833f
C779 B.n616 VSUBS 0.007833f
C780 B.n617 VSUBS 0.007833f
C781 B.n618 VSUBS 0.007833f
C782 B.n619 VSUBS 0.007833f
C783 B.n620 VSUBS 0.007833f
C784 B.n621 VSUBS 0.007833f
C785 B.n622 VSUBS 0.007833f
C786 B.n623 VSUBS 0.007833f
C787 B.n624 VSUBS 0.004377f
C788 B.n625 VSUBS 0.007833f
C789 B.n626 VSUBS 0.007833f
C790 B.n627 VSUBS 0.007372f
C791 B.n628 VSUBS 0.007833f
C792 B.n629 VSUBS 0.007833f
C793 B.n630 VSUBS 0.007833f
C794 B.n631 VSUBS 0.007833f
C795 B.n632 VSUBS 0.007833f
C796 B.n633 VSUBS 0.007833f
C797 B.n634 VSUBS 0.007833f
C798 B.n635 VSUBS 0.007833f
C799 B.n636 VSUBS 0.007833f
C800 B.n637 VSUBS 0.007833f
C801 B.n638 VSUBS 0.007833f
C802 B.n639 VSUBS 0.007833f
C803 B.n640 VSUBS 0.007833f
C804 B.n641 VSUBS 0.007833f
C805 B.n642 VSUBS 0.007833f
C806 B.n643 VSUBS 0.007833f
C807 B.n644 VSUBS 0.007833f
C808 B.n645 VSUBS 0.007833f
C809 B.n646 VSUBS 0.007833f
C810 B.n647 VSUBS 0.007833f
C811 B.n648 VSUBS 0.007833f
C812 B.n649 VSUBS 0.007833f
C813 B.n650 VSUBS 0.007833f
C814 B.n651 VSUBS 0.007833f
C815 B.n652 VSUBS 0.007833f
C816 B.n653 VSUBS 0.007833f
C817 B.n654 VSUBS 0.007833f
C818 B.n655 VSUBS 0.007833f
C819 B.n656 VSUBS 0.007833f
C820 B.n657 VSUBS 0.007833f
C821 B.n658 VSUBS 0.007833f
C822 B.n659 VSUBS 0.007833f
C823 B.n660 VSUBS 0.007833f
C824 B.n661 VSUBS 0.007833f
C825 B.n662 VSUBS 0.007833f
C826 B.n663 VSUBS 0.007833f
C827 B.n664 VSUBS 0.007833f
C828 B.n665 VSUBS 0.007833f
C829 B.n666 VSUBS 0.007833f
C830 B.n667 VSUBS 0.007833f
C831 B.n668 VSUBS 0.007833f
C832 B.n669 VSUBS 0.007833f
C833 B.n670 VSUBS 0.007833f
C834 B.n671 VSUBS 0.007833f
C835 B.n672 VSUBS 0.007833f
C836 B.n673 VSUBS 0.007833f
C837 B.n674 VSUBS 0.007833f
C838 B.n675 VSUBS 0.007833f
C839 B.n676 VSUBS 0.007833f
C840 B.n677 VSUBS 0.007833f
C841 B.n678 VSUBS 0.007833f
C842 B.n679 VSUBS 0.007833f
C843 B.n680 VSUBS 0.007833f
C844 B.n681 VSUBS 0.007833f
C845 B.n682 VSUBS 0.007833f
C846 B.n683 VSUBS 0.007833f
C847 B.n684 VSUBS 0.007833f
C848 B.n685 VSUBS 0.007833f
C849 B.n686 VSUBS 0.007833f
C850 B.n687 VSUBS 0.007833f
C851 B.n688 VSUBS 0.007833f
C852 B.n689 VSUBS 0.007833f
C853 B.n690 VSUBS 0.007833f
C854 B.n691 VSUBS 0.007833f
C855 B.n692 VSUBS 0.007833f
C856 B.n693 VSUBS 0.007833f
C857 B.n694 VSUBS 0.007833f
C858 B.n695 VSUBS 0.007833f
C859 B.n696 VSUBS 0.007833f
C860 B.n697 VSUBS 0.007833f
C861 B.n698 VSUBS 0.017836f
C862 B.n699 VSUBS 0.017836f
C863 B.n700 VSUBS 0.017182f
C864 B.n701 VSUBS 0.007833f
C865 B.n702 VSUBS 0.007833f
C866 B.n703 VSUBS 0.007833f
C867 B.n704 VSUBS 0.007833f
C868 B.n705 VSUBS 0.007833f
C869 B.n706 VSUBS 0.007833f
C870 B.n707 VSUBS 0.007833f
C871 B.n708 VSUBS 0.007833f
C872 B.n709 VSUBS 0.007833f
C873 B.n710 VSUBS 0.007833f
C874 B.n711 VSUBS 0.007833f
C875 B.n712 VSUBS 0.007833f
C876 B.n713 VSUBS 0.007833f
C877 B.n714 VSUBS 0.007833f
C878 B.n715 VSUBS 0.007833f
C879 B.n716 VSUBS 0.007833f
C880 B.n717 VSUBS 0.007833f
C881 B.n718 VSUBS 0.007833f
C882 B.n719 VSUBS 0.007833f
C883 B.n720 VSUBS 0.007833f
C884 B.n721 VSUBS 0.007833f
C885 B.n722 VSUBS 0.007833f
C886 B.n723 VSUBS 0.007833f
C887 B.n724 VSUBS 0.007833f
C888 B.n725 VSUBS 0.007833f
C889 B.n726 VSUBS 0.007833f
C890 B.n727 VSUBS 0.007833f
C891 B.n728 VSUBS 0.007833f
C892 B.n729 VSUBS 0.007833f
C893 B.n730 VSUBS 0.007833f
C894 B.n731 VSUBS 0.007833f
C895 B.n732 VSUBS 0.007833f
C896 B.n733 VSUBS 0.007833f
C897 B.n734 VSUBS 0.007833f
C898 B.n735 VSUBS 0.007833f
C899 B.n736 VSUBS 0.007833f
C900 B.n737 VSUBS 0.007833f
C901 B.n738 VSUBS 0.007833f
C902 B.n739 VSUBS 0.007833f
C903 B.n740 VSUBS 0.007833f
C904 B.n741 VSUBS 0.007833f
C905 B.n742 VSUBS 0.007833f
C906 B.n743 VSUBS 0.007833f
C907 B.n744 VSUBS 0.007833f
C908 B.n745 VSUBS 0.007833f
C909 B.n746 VSUBS 0.007833f
C910 B.n747 VSUBS 0.007833f
C911 B.n748 VSUBS 0.007833f
C912 B.n749 VSUBS 0.007833f
C913 B.n750 VSUBS 0.007833f
C914 B.n751 VSUBS 0.007833f
C915 B.n752 VSUBS 0.007833f
C916 B.n753 VSUBS 0.007833f
C917 B.n754 VSUBS 0.007833f
C918 B.n755 VSUBS 0.007833f
C919 B.n756 VSUBS 0.007833f
C920 B.n757 VSUBS 0.007833f
C921 B.n758 VSUBS 0.007833f
C922 B.n759 VSUBS 0.017737f
.ends

