* NGSPICE file created from diff_pair_sample_0271.ext - technology: sky130A

.subckt diff_pair_sample_0271 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=0 ps=0 w=9.24 l=0.32
X1 VDD1.t3 VP.t0 VTAIL.t7 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=1.5246 pd=9.57 as=3.6036 ps=19.26 w=9.24 l=0.32
X2 VTAIL.t4 VP.t1 VDD1.t2 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=1.5246 ps=9.57 w=9.24 l=0.32
X3 VTAIL.t2 VN.t0 VDD2.t3 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=1.5246 ps=9.57 w=9.24 l=0.32
X4 VDD1.t1 VP.t2 VTAIL.t6 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=1.5246 pd=9.57 as=3.6036 ps=19.26 w=9.24 l=0.32
X5 B.t8 B.t6 B.t7 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=0 ps=0 w=9.24 l=0.32
X6 B.t5 B.t3 B.t4 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=0 ps=0 w=9.24 l=0.32
X7 VDD2.t2 VN.t1 VTAIL.t1 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=1.5246 pd=9.57 as=3.6036 ps=19.26 w=9.24 l=0.32
X8 VTAIL.t5 VP.t3 VDD1.t0 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=1.5246 ps=9.57 w=9.24 l=0.32
X9 B.t2 B.t0 B.t1 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=0 ps=0 w=9.24 l=0.32
X10 VTAIL.t0 VN.t2 VDD2.t1 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=3.6036 pd=19.26 as=1.5246 ps=9.57 w=9.24 l=0.32
X11 VDD2.t0 VN.t3 VTAIL.t3 w_n1360_n2820# sky130_fd_pr__pfet_01v8 ad=1.5246 pd=9.57 as=3.6036 ps=19.26 w=9.24 l=0.32
R0 B.n84 B.t9 909.644
R1 B.n90 B.t6 909.644
R2 B.n26 B.t3 909.644
R3 B.n34 B.t0 909.644
R4 B.n297 B.n296 585
R5 B.n298 B.n51 585
R6 B.n300 B.n299 585
R7 B.n301 B.n50 585
R8 B.n303 B.n302 585
R9 B.n304 B.n49 585
R10 B.n306 B.n305 585
R11 B.n307 B.n48 585
R12 B.n309 B.n308 585
R13 B.n310 B.n47 585
R14 B.n312 B.n311 585
R15 B.n313 B.n46 585
R16 B.n315 B.n314 585
R17 B.n316 B.n45 585
R18 B.n318 B.n317 585
R19 B.n319 B.n44 585
R20 B.n321 B.n320 585
R21 B.n322 B.n43 585
R22 B.n324 B.n323 585
R23 B.n325 B.n42 585
R24 B.n327 B.n326 585
R25 B.n328 B.n41 585
R26 B.n330 B.n329 585
R27 B.n331 B.n40 585
R28 B.n333 B.n332 585
R29 B.n334 B.n39 585
R30 B.n336 B.n335 585
R31 B.n337 B.n38 585
R32 B.n339 B.n338 585
R33 B.n340 B.n37 585
R34 B.n342 B.n341 585
R35 B.n343 B.n36 585
R36 B.n345 B.n344 585
R37 B.n346 B.n33 585
R38 B.n349 B.n348 585
R39 B.n350 B.n32 585
R40 B.n352 B.n351 585
R41 B.n353 B.n31 585
R42 B.n355 B.n354 585
R43 B.n356 B.n30 585
R44 B.n358 B.n357 585
R45 B.n359 B.n29 585
R46 B.n361 B.n360 585
R47 B.n363 B.n362 585
R48 B.n364 B.n25 585
R49 B.n366 B.n365 585
R50 B.n367 B.n24 585
R51 B.n369 B.n368 585
R52 B.n370 B.n23 585
R53 B.n372 B.n371 585
R54 B.n373 B.n22 585
R55 B.n375 B.n374 585
R56 B.n376 B.n21 585
R57 B.n378 B.n377 585
R58 B.n379 B.n20 585
R59 B.n381 B.n380 585
R60 B.n382 B.n19 585
R61 B.n384 B.n383 585
R62 B.n385 B.n18 585
R63 B.n387 B.n386 585
R64 B.n388 B.n17 585
R65 B.n390 B.n389 585
R66 B.n391 B.n16 585
R67 B.n393 B.n392 585
R68 B.n394 B.n15 585
R69 B.n396 B.n395 585
R70 B.n397 B.n14 585
R71 B.n399 B.n398 585
R72 B.n400 B.n13 585
R73 B.n402 B.n401 585
R74 B.n403 B.n12 585
R75 B.n405 B.n404 585
R76 B.n406 B.n11 585
R77 B.n408 B.n407 585
R78 B.n409 B.n10 585
R79 B.n411 B.n410 585
R80 B.n412 B.n9 585
R81 B.n295 B.n52 585
R82 B.n294 B.n293 585
R83 B.n292 B.n53 585
R84 B.n291 B.n290 585
R85 B.n289 B.n54 585
R86 B.n288 B.n287 585
R87 B.n286 B.n55 585
R88 B.n285 B.n284 585
R89 B.n283 B.n56 585
R90 B.n282 B.n281 585
R91 B.n280 B.n57 585
R92 B.n279 B.n278 585
R93 B.n277 B.n58 585
R94 B.n276 B.n275 585
R95 B.n274 B.n59 585
R96 B.n273 B.n272 585
R97 B.n271 B.n60 585
R98 B.n270 B.n269 585
R99 B.n268 B.n61 585
R100 B.n267 B.n266 585
R101 B.n265 B.n62 585
R102 B.n264 B.n263 585
R103 B.n262 B.n63 585
R104 B.n261 B.n260 585
R105 B.n259 B.n64 585
R106 B.n258 B.n257 585
R107 B.n256 B.n65 585
R108 B.n255 B.n254 585
R109 B.n253 B.n66 585
R110 B.n136 B.n109 585
R111 B.n138 B.n137 585
R112 B.n139 B.n108 585
R113 B.n141 B.n140 585
R114 B.n142 B.n107 585
R115 B.n144 B.n143 585
R116 B.n145 B.n106 585
R117 B.n147 B.n146 585
R118 B.n148 B.n105 585
R119 B.n150 B.n149 585
R120 B.n151 B.n104 585
R121 B.n153 B.n152 585
R122 B.n154 B.n103 585
R123 B.n156 B.n155 585
R124 B.n157 B.n102 585
R125 B.n159 B.n158 585
R126 B.n160 B.n101 585
R127 B.n162 B.n161 585
R128 B.n163 B.n100 585
R129 B.n165 B.n164 585
R130 B.n166 B.n99 585
R131 B.n168 B.n167 585
R132 B.n169 B.n98 585
R133 B.n171 B.n170 585
R134 B.n172 B.n97 585
R135 B.n174 B.n173 585
R136 B.n175 B.n96 585
R137 B.n177 B.n176 585
R138 B.n178 B.n95 585
R139 B.n180 B.n179 585
R140 B.n181 B.n94 585
R141 B.n183 B.n182 585
R142 B.n184 B.n93 585
R143 B.n186 B.n185 585
R144 B.n188 B.n187 585
R145 B.n189 B.n89 585
R146 B.n191 B.n190 585
R147 B.n192 B.n88 585
R148 B.n194 B.n193 585
R149 B.n195 B.n87 585
R150 B.n197 B.n196 585
R151 B.n198 B.n86 585
R152 B.n200 B.n199 585
R153 B.n202 B.n83 585
R154 B.n204 B.n203 585
R155 B.n205 B.n82 585
R156 B.n207 B.n206 585
R157 B.n208 B.n81 585
R158 B.n210 B.n209 585
R159 B.n211 B.n80 585
R160 B.n213 B.n212 585
R161 B.n214 B.n79 585
R162 B.n216 B.n215 585
R163 B.n217 B.n78 585
R164 B.n219 B.n218 585
R165 B.n220 B.n77 585
R166 B.n222 B.n221 585
R167 B.n223 B.n76 585
R168 B.n225 B.n224 585
R169 B.n226 B.n75 585
R170 B.n228 B.n227 585
R171 B.n229 B.n74 585
R172 B.n231 B.n230 585
R173 B.n232 B.n73 585
R174 B.n234 B.n233 585
R175 B.n235 B.n72 585
R176 B.n237 B.n236 585
R177 B.n238 B.n71 585
R178 B.n240 B.n239 585
R179 B.n241 B.n70 585
R180 B.n243 B.n242 585
R181 B.n244 B.n69 585
R182 B.n246 B.n245 585
R183 B.n247 B.n68 585
R184 B.n249 B.n248 585
R185 B.n250 B.n67 585
R186 B.n252 B.n251 585
R187 B.n135 B.n134 585
R188 B.n133 B.n110 585
R189 B.n132 B.n131 585
R190 B.n130 B.n111 585
R191 B.n129 B.n128 585
R192 B.n127 B.n112 585
R193 B.n126 B.n125 585
R194 B.n124 B.n113 585
R195 B.n123 B.n122 585
R196 B.n121 B.n114 585
R197 B.n120 B.n119 585
R198 B.n118 B.n115 585
R199 B.n117 B.n116 585
R200 B.n2 B.n0 585
R201 B.n433 B.n1 585
R202 B.n432 B.n431 585
R203 B.n430 B.n3 585
R204 B.n429 B.n428 585
R205 B.n427 B.n4 585
R206 B.n426 B.n425 585
R207 B.n424 B.n5 585
R208 B.n423 B.n422 585
R209 B.n421 B.n6 585
R210 B.n420 B.n419 585
R211 B.n418 B.n7 585
R212 B.n417 B.n416 585
R213 B.n415 B.n8 585
R214 B.n414 B.n413 585
R215 B.n435 B.n434 585
R216 B.n134 B.n109 449.257
R217 B.n414 B.n9 449.257
R218 B.n253 B.n252 449.257
R219 B.n296 B.n295 449.257
R220 B.n84 B.t11 338.397
R221 B.n34 B.t1 338.397
R222 B.n90 B.t8 338.397
R223 B.n26 B.t4 338.397
R224 B.n85 B.t10 325.791
R225 B.n35 B.t2 325.791
R226 B.n91 B.t7 325.791
R227 B.n27 B.t5 325.791
R228 B.n134 B.n133 163.367
R229 B.n133 B.n132 163.367
R230 B.n132 B.n111 163.367
R231 B.n128 B.n111 163.367
R232 B.n128 B.n127 163.367
R233 B.n127 B.n126 163.367
R234 B.n126 B.n113 163.367
R235 B.n122 B.n113 163.367
R236 B.n122 B.n121 163.367
R237 B.n121 B.n120 163.367
R238 B.n120 B.n115 163.367
R239 B.n116 B.n115 163.367
R240 B.n116 B.n2 163.367
R241 B.n434 B.n2 163.367
R242 B.n434 B.n433 163.367
R243 B.n433 B.n432 163.367
R244 B.n432 B.n3 163.367
R245 B.n428 B.n3 163.367
R246 B.n428 B.n427 163.367
R247 B.n427 B.n426 163.367
R248 B.n426 B.n5 163.367
R249 B.n422 B.n5 163.367
R250 B.n422 B.n421 163.367
R251 B.n421 B.n420 163.367
R252 B.n420 B.n7 163.367
R253 B.n416 B.n7 163.367
R254 B.n416 B.n415 163.367
R255 B.n415 B.n414 163.367
R256 B.n138 B.n109 163.367
R257 B.n139 B.n138 163.367
R258 B.n140 B.n139 163.367
R259 B.n140 B.n107 163.367
R260 B.n144 B.n107 163.367
R261 B.n145 B.n144 163.367
R262 B.n146 B.n145 163.367
R263 B.n146 B.n105 163.367
R264 B.n150 B.n105 163.367
R265 B.n151 B.n150 163.367
R266 B.n152 B.n151 163.367
R267 B.n152 B.n103 163.367
R268 B.n156 B.n103 163.367
R269 B.n157 B.n156 163.367
R270 B.n158 B.n157 163.367
R271 B.n158 B.n101 163.367
R272 B.n162 B.n101 163.367
R273 B.n163 B.n162 163.367
R274 B.n164 B.n163 163.367
R275 B.n164 B.n99 163.367
R276 B.n168 B.n99 163.367
R277 B.n169 B.n168 163.367
R278 B.n170 B.n169 163.367
R279 B.n170 B.n97 163.367
R280 B.n174 B.n97 163.367
R281 B.n175 B.n174 163.367
R282 B.n176 B.n175 163.367
R283 B.n176 B.n95 163.367
R284 B.n180 B.n95 163.367
R285 B.n181 B.n180 163.367
R286 B.n182 B.n181 163.367
R287 B.n182 B.n93 163.367
R288 B.n186 B.n93 163.367
R289 B.n187 B.n186 163.367
R290 B.n187 B.n89 163.367
R291 B.n191 B.n89 163.367
R292 B.n192 B.n191 163.367
R293 B.n193 B.n192 163.367
R294 B.n193 B.n87 163.367
R295 B.n197 B.n87 163.367
R296 B.n198 B.n197 163.367
R297 B.n199 B.n198 163.367
R298 B.n199 B.n83 163.367
R299 B.n204 B.n83 163.367
R300 B.n205 B.n204 163.367
R301 B.n206 B.n205 163.367
R302 B.n206 B.n81 163.367
R303 B.n210 B.n81 163.367
R304 B.n211 B.n210 163.367
R305 B.n212 B.n211 163.367
R306 B.n212 B.n79 163.367
R307 B.n216 B.n79 163.367
R308 B.n217 B.n216 163.367
R309 B.n218 B.n217 163.367
R310 B.n218 B.n77 163.367
R311 B.n222 B.n77 163.367
R312 B.n223 B.n222 163.367
R313 B.n224 B.n223 163.367
R314 B.n224 B.n75 163.367
R315 B.n228 B.n75 163.367
R316 B.n229 B.n228 163.367
R317 B.n230 B.n229 163.367
R318 B.n230 B.n73 163.367
R319 B.n234 B.n73 163.367
R320 B.n235 B.n234 163.367
R321 B.n236 B.n235 163.367
R322 B.n236 B.n71 163.367
R323 B.n240 B.n71 163.367
R324 B.n241 B.n240 163.367
R325 B.n242 B.n241 163.367
R326 B.n242 B.n69 163.367
R327 B.n246 B.n69 163.367
R328 B.n247 B.n246 163.367
R329 B.n248 B.n247 163.367
R330 B.n248 B.n67 163.367
R331 B.n252 B.n67 163.367
R332 B.n254 B.n253 163.367
R333 B.n254 B.n65 163.367
R334 B.n258 B.n65 163.367
R335 B.n259 B.n258 163.367
R336 B.n260 B.n259 163.367
R337 B.n260 B.n63 163.367
R338 B.n264 B.n63 163.367
R339 B.n265 B.n264 163.367
R340 B.n266 B.n265 163.367
R341 B.n266 B.n61 163.367
R342 B.n270 B.n61 163.367
R343 B.n271 B.n270 163.367
R344 B.n272 B.n271 163.367
R345 B.n272 B.n59 163.367
R346 B.n276 B.n59 163.367
R347 B.n277 B.n276 163.367
R348 B.n278 B.n277 163.367
R349 B.n278 B.n57 163.367
R350 B.n282 B.n57 163.367
R351 B.n283 B.n282 163.367
R352 B.n284 B.n283 163.367
R353 B.n284 B.n55 163.367
R354 B.n288 B.n55 163.367
R355 B.n289 B.n288 163.367
R356 B.n290 B.n289 163.367
R357 B.n290 B.n53 163.367
R358 B.n294 B.n53 163.367
R359 B.n295 B.n294 163.367
R360 B.n410 B.n9 163.367
R361 B.n410 B.n409 163.367
R362 B.n409 B.n408 163.367
R363 B.n408 B.n11 163.367
R364 B.n404 B.n11 163.367
R365 B.n404 B.n403 163.367
R366 B.n403 B.n402 163.367
R367 B.n402 B.n13 163.367
R368 B.n398 B.n13 163.367
R369 B.n398 B.n397 163.367
R370 B.n397 B.n396 163.367
R371 B.n396 B.n15 163.367
R372 B.n392 B.n15 163.367
R373 B.n392 B.n391 163.367
R374 B.n391 B.n390 163.367
R375 B.n390 B.n17 163.367
R376 B.n386 B.n17 163.367
R377 B.n386 B.n385 163.367
R378 B.n385 B.n384 163.367
R379 B.n384 B.n19 163.367
R380 B.n380 B.n19 163.367
R381 B.n380 B.n379 163.367
R382 B.n379 B.n378 163.367
R383 B.n378 B.n21 163.367
R384 B.n374 B.n21 163.367
R385 B.n374 B.n373 163.367
R386 B.n373 B.n372 163.367
R387 B.n372 B.n23 163.367
R388 B.n368 B.n23 163.367
R389 B.n368 B.n367 163.367
R390 B.n367 B.n366 163.367
R391 B.n366 B.n25 163.367
R392 B.n362 B.n25 163.367
R393 B.n362 B.n361 163.367
R394 B.n361 B.n29 163.367
R395 B.n357 B.n29 163.367
R396 B.n357 B.n356 163.367
R397 B.n356 B.n355 163.367
R398 B.n355 B.n31 163.367
R399 B.n351 B.n31 163.367
R400 B.n351 B.n350 163.367
R401 B.n350 B.n349 163.367
R402 B.n349 B.n33 163.367
R403 B.n344 B.n33 163.367
R404 B.n344 B.n343 163.367
R405 B.n343 B.n342 163.367
R406 B.n342 B.n37 163.367
R407 B.n338 B.n37 163.367
R408 B.n338 B.n337 163.367
R409 B.n337 B.n336 163.367
R410 B.n336 B.n39 163.367
R411 B.n332 B.n39 163.367
R412 B.n332 B.n331 163.367
R413 B.n331 B.n330 163.367
R414 B.n330 B.n41 163.367
R415 B.n326 B.n41 163.367
R416 B.n326 B.n325 163.367
R417 B.n325 B.n324 163.367
R418 B.n324 B.n43 163.367
R419 B.n320 B.n43 163.367
R420 B.n320 B.n319 163.367
R421 B.n319 B.n318 163.367
R422 B.n318 B.n45 163.367
R423 B.n314 B.n45 163.367
R424 B.n314 B.n313 163.367
R425 B.n313 B.n312 163.367
R426 B.n312 B.n47 163.367
R427 B.n308 B.n47 163.367
R428 B.n308 B.n307 163.367
R429 B.n307 B.n306 163.367
R430 B.n306 B.n49 163.367
R431 B.n302 B.n49 163.367
R432 B.n302 B.n301 163.367
R433 B.n301 B.n300 163.367
R434 B.n300 B.n51 163.367
R435 B.n296 B.n51 163.367
R436 B.n201 B.n85 59.5399
R437 B.n92 B.n91 59.5399
R438 B.n28 B.n27 59.5399
R439 B.n347 B.n35 59.5399
R440 B.n413 B.n412 29.1907
R441 B.n297 B.n52 29.1907
R442 B.n251 B.n66 29.1907
R443 B.n136 B.n135 29.1907
R444 B B.n435 18.0485
R445 B.n85 B.n84 12.6066
R446 B.n91 B.n90 12.6066
R447 B.n27 B.n26 12.6066
R448 B.n35 B.n34 12.6066
R449 B.n412 B.n411 10.6151
R450 B.n411 B.n10 10.6151
R451 B.n407 B.n10 10.6151
R452 B.n407 B.n406 10.6151
R453 B.n406 B.n405 10.6151
R454 B.n405 B.n12 10.6151
R455 B.n401 B.n12 10.6151
R456 B.n401 B.n400 10.6151
R457 B.n400 B.n399 10.6151
R458 B.n399 B.n14 10.6151
R459 B.n395 B.n14 10.6151
R460 B.n395 B.n394 10.6151
R461 B.n394 B.n393 10.6151
R462 B.n393 B.n16 10.6151
R463 B.n389 B.n16 10.6151
R464 B.n389 B.n388 10.6151
R465 B.n388 B.n387 10.6151
R466 B.n387 B.n18 10.6151
R467 B.n383 B.n18 10.6151
R468 B.n383 B.n382 10.6151
R469 B.n382 B.n381 10.6151
R470 B.n381 B.n20 10.6151
R471 B.n377 B.n20 10.6151
R472 B.n377 B.n376 10.6151
R473 B.n376 B.n375 10.6151
R474 B.n375 B.n22 10.6151
R475 B.n371 B.n22 10.6151
R476 B.n371 B.n370 10.6151
R477 B.n370 B.n369 10.6151
R478 B.n369 B.n24 10.6151
R479 B.n365 B.n24 10.6151
R480 B.n365 B.n364 10.6151
R481 B.n364 B.n363 10.6151
R482 B.n360 B.n359 10.6151
R483 B.n359 B.n358 10.6151
R484 B.n358 B.n30 10.6151
R485 B.n354 B.n30 10.6151
R486 B.n354 B.n353 10.6151
R487 B.n353 B.n352 10.6151
R488 B.n352 B.n32 10.6151
R489 B.n348 B.n32 10.6151
R490 B.n346 B.n345 10.6151
R491 B.n345 B.n36 10.6151
R492 B.n341 B.n36 10.6151
R493 B.n341 B.n340 10.6151
R494 B.n340 B.n339 10.6151
R495 B.n339 B.n38 10.6151
R496 B.n335 B.n38 10.6151
R497 B.n335 B.n334 10.6151
R498 B.n334 B.n333 10.6151
R499 B.n333 B.n40 10.6151
R500 B.n329 B.n40 10.6151
R501 B.n329 B.n328 10.6151
R502 B.n328 B.n327 10.6151
R503 B.n327 B.n42 10.6151
R504 B.n323 B.n42 10.6151
R505 B.n323 B.n322 10.6151
R506 B.n322 B.n321 10.6151
R507 B.n321 B.n44 10.6151
R508 B.n317 B.n44 10.6151
R509 B.n317 B.n316 10.6151
R510 B.n316 B.n315 10.6151
R511 B.n315 B.n46 10.6151
R512 B.n311 B.n46 10.6151
R513 B.n311 B.n310 10.6151
R514 B.n310 B.n309 10.6151
R515 B.n309 B.n48 10.6151
R516 B.n305 B.n48 10.6151
R517 B.n305 B.n304 10.6151
R518 B.n304 B.n303 10.6151
R519 B.n303 B.n50 10.6151
R520 B.n299 B.n50 10.6151
R521 B.n299 B.n298 10.6151
R522 B.n298 B.n297 10.6151
R523 B.n255 B.n66 10.6151
R524 B.n256 B.n255 10.6151
R525 B.n257 B.n256 10.6151
R526 B.n257 B.n64 10.6151
R527 B.n261 B.n64 10.6151
R528 B.n262 B.n261 10.6151
R529 B.n263 B.n262 10.6151
R530 B.n263 B.n62 10.6151
R531 B.n267 B.n62 10.6151
R532 B.n268 B.n267 10.6151
R533 B.n269 B.n268 10.6151
R534 B.n269 B.n60 10.6151
R535 B.n273 B.n60 10.6151
R536 B.n274 B.n273 10.6151
R537 B.n275 B.n274 10.6151
R538 B.n275 B.n58 10.6151
R539 B.n279 B.n58 10.6151
R540 B.n280 B.n279 10.6151
R541 B.n281 B.n280 10.6151
R542 B.n281 B.n56 10.6151
R543 B.n285 B.n56 10.6151
R544 B.n286 B.n285 10.6151
R545 B.n287 B.n286 10.6151
R546 B.n287 B.n54 10.6151
R547 B.n291 B.n54 10.6151
R548 B.n292 B.n291 10.6151
R549 B.n293 B.n292 10.6151
R550 B.n293 B.n52 10.6151
R551 B.n137 B.n136 10.6151
R552 B.n137 B.n108 10.6151
R553 B.n141 B.n108 10.6151
R554 B.n142 B.n141 10.6151
R555 B.n143 B.n142 10.6151
R556 B.n143 B.n106 10.6151
R557 B.n147 B.n106 10.6151
R558 B.n148 B.n147 10.6151
R559 B.n149 B.n148 10.6151
R560 B.n149 B.n104 10.6151
R561 B.n153 B.n104 10.6151
R562 B.n154 B.n153 10.6151
R563 B.n155 B.n154 10.6151
R564 B.n155 B.n102 10.6151
R565 B.n159 B.n102 10.6151
R566 B.n160 B.n159 10.6151
R567 B.n161 B.n160 10.6151
R568 B.n161 B.n100 10.6151
R569 B.n165 B.n100 10.6151
R570 B.n166 B.n165 10.6151
R571 B.n167 B.n166 10.6151
R572 B.n167 B.n98 10.6151
R573 B.n171 B.n98 10.6151
R574 B.n172 B.n171 10.6151
R575 B.n173 B.n172 10.6151
R576 B.n173 B.n96 10.6151
R577 B.n177 B.n96 10.6151
R578 B.n178 B.n177 10.6151
R579 B.n179 B.n178 10.6151
R580 B.n179 B.n94 10.6151
R581 B.n183 B.n94 10.6151
R582 B.n184 B.n183 10.6151
R583 B.n185 B.n184 10.6151
R584 B.n189 B.n188 10.6151
R585 B.n190 B.n189 10.6151
R586 B.n190 B.n88 10.6151
R587 B.n194 B.n88 10.6151
R588 B.n195 B.n194 10.6151
R589 B.n196 B.n195 10.6151
R590 B.n196 B.n86 10.6151
R591 B.n200 B.n86 10.6151
R592 B.n203 B.n202 10.6151
R593 B.n203 B.n82 10.6151
R594 B.n207 B.n82 10.6151
R595 B.n208 B.n207 10.6151
R596 B.n209 B.n208 10.6151
R597 B.n209 B.n80 10.6151
R598 B.n213 B.n80 10.6151
R599 B.n214 B.n213 10.6151
R600 B.n215 B.n214 10.6151
R601 B.n215 B.n78 10.6151
R602 B.n219 B.n78 10.6151
R603 B.n220 B.n219 10.6151
R604 B.n221 B.n220 10.6151
R605 B.n221 B.n76 10.6151
R606 B.n225 B.n76 10.6151
R607 B.n226 B.n225 10.6151
R608 B.n227 B.n226 10.6151
R609 B.n227 B.n74 10.6151
R610 B.n231 B.n74 10.6151
R611 B.n232 B.n231 10.6151
R612 B.n233 B.n232 10.6151
R613 B.n233 B.n72 10.6151
R614 B.n237 B.n72 10.6151
R615 B.n238 B.n237 10.6151
R616 B.n239 B.n238 10.6151
R617 B.n239 B.n70 10.6151
R618 B.n243 B.n70 10.6151
R619 B.n244 B.n243 10.6151
R620 B.n245 B.n244 10.6151
R621 B.n245 B.n68 10.6151
R622 B.n249 B.n68 10.6151
R623 B.n250 B.n249 10.6151
R624 B.n251 B.n250 10.6151
R625 B.n135 B.n110 10.6151
R626 B.n131 B.n110 10.6151
R627 B.n131 B.n130 10.6151
R628 B.n130 B.n129 10.6151
R629 B.n129 B.n112 10.6151
R630 B.n125 B.n112 10.6151
R631 B.n125 B.n124 10.6151
R632 B.n124 B.n123 10.6151
R633 B.n123 B.n114 10.6151
R634 B.n119 B.n114 10.6151
R635 B.n119 B.n118 10.6151
R636 B.n118 B.n117 10.6151
R637 B.n117 B.n0 10.6151
R638 B.n431 B.n1 10.6151
R639 B.n431 B.n430 10.6151
R640 B.n430 B.n429 10.6151
R641 B.n429 B.n4 10.6151
R642 B.n425 B.n4 10.6151
R643 B.n425 B.n424 10.6151
R644 B.n424 B.n423 10.6151
R645 B.n423 B.n6 10.6151
R646 B.n419 B.n6 10.6151
R647 B.n419 B.n418 10.6151
R648 B.n418 B.n417 10.6151
R649 B.n417 B.n8 10.6151
R650 B.n413 B.n8 10.6151
R651 B.n360 B.n28 7.18099
R652 B.n348 B.n347 7.18099
R653 B.n188 B.n92 7.18099
R654 B.n201 B.n200 7.18099
R655 B.n363 B.n28 3.43465
R656 B.n347 B.n346 3.43465
R657 B.n185 B.n92 3.43465
R658 B.n202 B.n201 3.43465
R659 B.n435 B.n0 2.81026
R660 B.n435 B.n1 2.81026
R661 VP.n1 VP.t2 842.77
R662 VP.n1 VP.t3 842.77
R663 VP.n0 VP.t1 842.77
R664 VP.n0 VP.t0 842.77
R665 VP.n2 VP.n0 198.573
R666 VP.n2 VP.n1 161.3
R667 VP VP.n2 0.0516364
R668 VTAIL.n394 VTAIL.n350 756.745
R669 VTAIL.n44 VTAIL.n0 756.745
R670 VTAIL.n94 VTAIL.n50 756.745
R671 VTAIL.n144 VTAIL.n100 756.745
R672 VTAIL.n344 VTAIL.n300 756.745
R673 VTAIL.n294 VTAIL.n250 756.745
R674 VTAIL.n244 VTAIL.n200 756.745
R675 VTAIL.n194 VTAIL.n150 756.745
R676 VTAIL.n367 VTAIL.n366 585
R677 VTAIL.n369 VTAIL.n368 585
R678 VTAIL.n362 VTAIL.n361 585
R679 VTAIL.n375 VTAIL.n374 585
R680 VTAIL.n377 VTAIL.n376 585
R681 VTAIL.n358 VTAIL.n357 585
R682 VTAIL.n384 VTAIL.n383 585
R683 VTAIL.n385 VTAIL.n356 585
R684 VTAIL.n387 VTAIL.n386 585
R685 VTAIL.n354 VTAIL.n353 585
R686 VTAIL.n393 VTAIL.n392 585
R687 VTAIL.n395 VTAIL.n394 585
R688 VTAIL.n17 VTAIL.n16 585
R689 VTAIL.n19 VTAIL.n18 585
R690 VTAIL.n12 VTAIL.n11 585
R691 VTAIL.n25 VTAIL.n24 585
R692 VTAIL.n27 VTAIL.n26 585
R693 VTAIL.n8 VTAIL.n7 585
R694 VTAIL.n34 VTAIL.n33 585
R695 VTAIL.n35 VTAIL.n6 585
R696 VTAIL.n37 VTAIL.n36 585
R697 VTAIL.n4 VTAIL.n3 585
R698 VTAIL.n43 VTAIL.n42 585
R699 VTAIL.n45 VTAIL.n44 585
R700 VTAIL.n67 VTAIL.n66 585
R701 VTAIL.n69 VTAIL.n68 585
R702 VTAIL.n62 VTAIL.n61 585
R703 VTAIL.n75 VTAIL.n74 585
R704 VTAIL.n77 VTAIL.n76 585
R705 VTAIL.n58 VTAIL.n57 585
R706 VTAIL.n84 VTAIL.n83 585
R707 VTAIL.n85 VTAIL.n56 585
R708 VTAIL.n87 VTAIL.n86 585
R709 VTAIL.n54 VTAIL.n53 585
R710 VTAIL.n93 VTAIL.n92 585
R711 VTAIL.n95 VTAIL.n94 585
R712 VTAIL.n117 VTAIL.n116 585
R713 VTAIL.n119 VTAIL.n118 585
R714 VTAIL.n112 VTAIL.n111 585
R715 VTAIL.n125 VTAIL.n124 585
R716 VTAIL.n127 VTAIL.n126 585
R717 VTAIL.n108 VTAIL.n107 585
R718 VTAIL.n134 VTAIL.n133 585
R719 VTAIL.n135 VTAIL.n106 585
R720 VTAIL.n137 VTAIL.n136 585
R721 VTAIL.n104 VTAIL.n103 585
R722 VTAIL.n143 VTAIL.n142 585
R723 VTAIL.n145 VTAIL.n144 585
R724 VTAIL.n345 VTAIL.n344 585
R725 VTAIL.n343 VTAIL.n342 585
R726 VTAIL.n304 VTAIL.n303 585
R727 VTAIL.n308 VTAIL.n306 585
R728 VTAIL.n337 VTAIL.n336 585
R729 VTAIL.n335 VTAIL.n334 585
R730 VTAIL.n310 VTAIL.n309 585
R731 VTAIL.n329 VTAIL.n328 585
R732 VTAIL.n327 VTAIL.n326 585
R733 VTAIL.n314 VTAIL.n313 585
R734 VTAIL.n321 VTAIL.n320 585
R735 VTAIL.n319 VTAIL.n318 585
R736 VTAIL.n295 VTAIL.n294 585
R737 VTAIL.n293 VTAIL.n292 585
R738 VTAIL.n254 VTAIL.n253 585
R739 VTAIL.n258 VTAIL.n256 585
R740 VTAIL.n287 VTAIL.n286 585
R741 VTAIL.n285 VTAIL.n284 585
R742 VTAIL.n260 VTAIL.n259 585
R743 VTAIL.n279 VTAIL.n278 585
R744 VTAIL.n277 VTAIL.n276 585
R745 VTAIL.n264 VTAIL.n263 585
R746 VTAIL.n271 VTAIL.n270 585
R747 VTAIL.n269 VTAIL.n268 585
R748 VTAIL.n245 VTAIL.n244 585
R749 VTAIL.n243 VTAIL.n242 585
R750 VTAIL.n204 VTAIL.n203 585
R751 VTAIL.n208 VTAIL.n206 585
R752 VTAIL.n237 VTAIL.n236 585
R753 VTAIL.n235 VTAIL.n234 585
R754 VTAIL.n210 VTAIL.n209 585
R755 VTAIL.n229 VTAIL.n228 585
R756 VTAIL.n227 VTAIL.n226 585
R757 VTAIL.n214 VTAIL.n213 585
R758 VTAIL.n221 VTAIL.n220 585
R759 VTAIL.n219 VTAIL.n218 585
R760 VTAIL.n195 VTAIL.n194 585
R761 VTAIL.n193 VTAIL.n192 585
R762 VTAIL.n154 VTAIL.n153 585
R763 VTAIL.n158 VTAIL.n156 585
R764 VTAIL.n187 VTAIL.n186 585
R765 VTAIL.n185 VTAIL.n184 585
R766 VTAIL.n160 VTAIL.n159 585
R767 VTAIL.n179 VTAIL.n178 585
R768 VTAIL.n177 VTAIL.n176 585
R769 VTAIL.n164 VTAIL.n163 585
R770 VTAIL.n171 VTAIL.n170 585
R771 VTAIL.n169 VTAIL.n168 585
R772 VTAIL.n365 VTAIL.t1 329.038
R773 VTAIL.n15 VTAIL.t2 329.038
R774 VTAIL.n65 VTAIL.t6 329.038
R775 VTAIL.n115 VTAIL.t5 329.038
R776 VTAIL.n317 VTAIL.t7 329.038
R777 VTAIL.n267 VTAIL.t4 329.038
R778 VTAIL.n217 VTAIL.t3 329.038
R779 VTAIL.n167 VTAIL.t0 329.038
R780 VTAIL.n368 VTAIL.n367 171.744
R781 VTAIL.n368 VTAIL.n361 171.744
R782 VTAIL.n375 VTAIL.n361 171.744
R783 VTAIL.n376 VTAIL.n375 171.744
R784 VTAIL.n376 VTAIL.n357 171.744
R785 VTAIL.n384 VTAIL.n357 171.744
R786 VTAIL.n385 VTAIL.n384 171.744
R787 VTAIL.n386 VTAIL.n385 171.744
R788 VTAIL.n386 VTAIL.n353 171.744
R789 VTAIL.n393 VTAIL.n353 171.744
R790 VTAIL.n394 VTAIL.n393 171.744
R791 VTAIL.n18 VTAIL.n17 171.744
R792 VTAIL.n18 VTAIL.n11 171.744
R793 VTAIL.n25 VTAIL.n11 171.744
R794 VTAIL.n26 VTAIL.n25 171.744
R795 VTAIL.n26 VTAIL.n7 171.744
R796 VTAIL.n34 VTAIL.n7 171.744
R797 VTAIL.n35 VTAIL.n34 171.744
R798 VTAIL.n36 VTAIL.n35 171.744
R799 VTAIL.n36 VTAIL.n3 171.744
R800 VTAIL.n43 VTAIL.n3 171.744
R801 VTAIL.n44 VTAIL.n43 171.744
R802 VTAIL.n68 VTAIL.n67 171.744
R803 VTAIL.n68 VTAIL.n61 171.744
R804 VTAIL.n75 VTAIL.n61 171.744
R805 VTAIL.n76 VTAIL.n75 171.744
R806 VTAIL.n76 VTAIL.n57 171.744
R807 VTAIL.n84 VTAIL.n57 171.744
R808 VTAIL.n85 VTAIL.n84 171.744
R809 VTAIL.n86 VTAIL.n85 171.744
R810 VTAIL.n86 VTAIL.n53 171.744
R811 VTAIL.n93 VTAIL.n53 171.744
R812 VTAIL.n94 VTAIL.n93 171.744
R813 VTAIL.n118 VTAIL.n117 171.744
R814 VTAIL.n118 VTAIL.n111 171.744
R815 VTAIL.n125 VTAIL.n111 171.744
R816 VTAIL.n126 VTAIL.n125 171.744
R817 VTAIL.n126 VTAIL.n107 171.744
R818 VTAIL.n134 VTAIL.n107 171.744
R819 VTAIL.n135 VTAIL.n134 171.744
R820 VTAIL.n136 VTAIL.n135 171.744
R821 VTAIL.n136 VTAIL.n103 171.744
R822 VTAIL.n143 VTAIL.n103 171.744
R823 VTAIL.n144 VTAIL.n143 171.744
R824 VTAIL.n344 VTAIL.n343 171.744
R825 VTAIL.n343 VTAIL.n303 171.744
R826 VTAIL.n308 VTAIL.n303 171.744
R827 VTAIL.n336 VTAIL.n308 171.744
R828 VTAIL.n336 VTAIL.n335 171.744
R829 VTAIL.n335 VTAIL.n309 171.744
R830 VTAIL.n328 VTAIL.n309 171.744
R831 VTAIL.n328 VTAIL.n327 171.744
R832 VTAIL.n327 VTAIL.n313 171.744
R833 VTAIL.n320 VTAIL.n313 171.744
R834 VTAIL.n320 VTAIL.n319 171.744
R835 VTAIL.n294 VTAIL.n293 171.744
R836 VTAIL.n293 VTAIL.n253 171.744
R837 VTAIL.n258 VTAIL.n253 171.744
R838 VTAIL.n286 VTAIL.n258 171.744
R839 VTAIL.n286 VTAIL.n285 171.744
R840 VTAIL.n285 VTAIL.n259 171.744
R841 VTAIL.n278 VTAIL.n259 171.744
R842 VTAIL.n278 VTAIL.n277 171.744
R843 VTAIL.n277 VTAIL.n263 171.744
R844 VTAIL.n270 VTAIL.n263 171.744
R845 VTAIL.n270 VTAIL.n269 171.744
R846 VTAIL.n244 VTAIL.n243 171.744
R847 VTAIL.n243 VTAIL.n203 171.744
R848 VTAIL.n208 VTAIL.n203 171.744
R849 VTAIL.n236 VTAIL.n208 171.744
R850 VTAIL.n236 VTAIL.n235 171.744
R851 VTAIL.n235 VTAIL.n209 171.744
R852 VTAIL.n228 VTAIL.n209 171.744
R853 VTAIL.n228 VTAIL.n227 171.744
R854 VTAIL.n227 VTAIL.n213 171.744
R855 VTAIL.n220 VTAIL.n213 171.744
R856 VTAIL.n220 VTAIL.n219 171.744
R857 VTAIL.n194 VTAIL.n193 171.744
R858 VTAIL.n193 VTAIL.n153 171.744
R859 VTAIL.n158 VTAIL.n153 171.744
R860 VTAIL.n186 VTAIL.n158 171.744
R861 VTAIL.n186 VTAIL.n185 171.744
R862 VTAIL.n185 VTAIL.n159 171.744
R863 VTAIL.n178 VTAIL.n159 171.744
R864 VTAIL.n178 VTAIL.n177 171.744
R865 VTAIL.n177 VTAIL.n163 171.744
R866 VTAIL.n170 VTAIL.n163 171.744
R867 VTAIL.n170 VTAIL.n169 171.744
R868 VTAIL.n367 VTAIL.t1 85.8723
R869 VTAIL.n17 VTAIL.t2 85.8723
R870 VTAIL.n67 VTAIL.t6 85.8723
R871 VTAIL.n117 VTAIL.t5 85.8723
R872 VTAIL.n319 VTAIL.t7 85.8723
R873 VTAIL.n269 VTAIL.t4 85.8723
R874 VTAIL.n219 VTAIL.t3 85.8723
R875 VTAIL.n169 VTAIL.t0 85.8723
R876 VTAIL.n399 VTAIL.n398 32.1853
R877 VTAIL.n49 VTAIL.n48 32.1853
R878 VTAIL.n99 VTAIL.n98 32.1853
R879 VTAIL.n149 VTAIL.n148 32.1853
R880 VTAIL.n349 VTAIL.n348 32.1853
R881 VTAIL.n299 VTAIL.n298 32.1853
R882 VTAIL.n249 VTAIL.n248 32.1853
R883 VTAIL.n199 VTAIL.n198 32.1853
R884 VTAIL.n399 VTAIL.n349 20.91
R885 VTAIL.n199 VTAIL.n149 20.91
R886 VTAIL.n387 VTAIL.n354 13.1884
R887 VTAIL.n37 VTAIL.n4 13.1884
R888 VTAIL.n87 VTAIL.n54 13.1884
R889 VTAIL.n137 VTAIL.n104 13.1884
R890 VTAIL.n306 VTAIL.n304 13.1884
R891 VTAIL.n256 VTAIL.n254 13.1884
R892 VTAIL.n206 VTAIL.n204 13.1884
R893 VTAIL.n156 VTAIL.n154 13.1884
R894 VTAIL.n388 VTAIL.n356 12.8005
R895 VTAIL.n392 VTAIL.n391 12.8005
R896 VTAIL.n38 VTAIL.n6 12.8005
R897 VTAIL.n42 VTAIL.n41 12.8005
R898 VTAIL.n88 VTAIL.n56 12.8005
R899 VTAIL.n92 VTAIL.n91 12.8005
R900 VTAIL.n138 VTAIL.n106 12.8005
R901 VTAIL.n142 VTAIL.n141 12.8005
R902 VTAIL.n342 VTAIL.n341 12.8005
R903 VTAIL.n338 VTAIL.n337 12.8005
R904 VTAIL.n292 VTAIL.n291 12.8005
R905 VTAIL.n288 VTAIL.n287 12.8005
R906 VTAIL.n242 VTAIL.n241 12.8005
R907 VTAIL.n238 VTAIL.n237 12.8005
R908 VTAIL.n192 VTAIL.n191 12.8005
R909 VTAIL.n188 VTAIL.n187 12.8005
R910 VTAIL.n383 VTAIL.n382 12.0247
R911 VTAIL.n395 VTAIL.n352 12.0247
R912 VTAIL.n33 VTAIL.n32 12.0247
R913 VTAIL.n45 VTAIL.n2 12.0247
R914 VTAIL.n83 VTAIL.n82 12.0247
R915 VTAIL.n95 VTAIL.n52 12.0247
R916 VTAIL.n133 VTAIL.n132 12.0247
R917 VTAIL.n145 VTAIL.n102 12.0247
R918 VTAIL.n345 VTAIL.n302 12.0247
R919 VTAIL.n334 VTAIL.n307 12.0247
R920 VTAIL.n295 VTAIL.n252 12.0247
R921 VTAIL.n284 VTAIL.n257 12.0247
R922 VTAIL.n245 VTAIL.n202 12.0247
R923 VTAIL.n234 VTAIL.n207 12.0247
R924 VTAIL.n195 VTAIL.n152 12.0247
R925 VTAIL.n184 VTAIL.n157 12.0247
R926 VTAIL.n381 VTAIL.n358 11.249
R927 VTAIL.n396 VTAIL.n350 11.249
R928 VTAIL.n31 VTAIL.n8 11.249
R929 VTAIL.n46 VTAIL.n0 11.249
R930 VTAIL.n81 VTAIL.n58 11.249
R931 VTAIL.n96 VTAIL.n50 11.249
R932 VTAIL.n131 VTAIL.n108 11.249
R933 VTAIL.n146 VTAIL.n100 11.249
R934 VTAIL.n346 VTAIL.n300 11.249
R935 VTAIL.n333 VTAIL.n310 11.249
R936 VTAIL.n296 VTAIL.n250 11.249
R937 VTAIL.n283 VTAIL.n260 11.249
R938 VTAIL.n246 VTAIL.n200 11.249
R939 VTAIL.n233 VTAIL.n210 11.249
R940 VTAIL.n196 VTAIL.n150 11.249
R941 VTAIL.n183 VTAIL.n160 11.249
R942 VTAIL.n366 VTAIL.n365 10.7239
R943 VTAIL.n16 VTAIL.n15 10.7239
R944 VTAIL.n66 VTAIL.n65 10.7239
R945 VTAIL.n116 VTAIL.n115 10.7239
R946 VTAIL.n318 VTAIL.n317 10.7239
R947 VTAIL.n268 VTAIL.n267 10.7239
R948 VTAIL.n218 VTAIL.n217 10.7239
R949 VTAIL.n168 VTAIL.n167 10.7239
R950 VTAIL.n378 VTAIL.n377 10.4732
R951 VTAIL.n28 VTAIL.n27 10.4732
R952 VTAIL.n78 VTAIL.n77 10.4732
R953 VTAIL.n128 VTAIL.n127 10.4732
R954 VTAIL.n330 VTAIL.n329 10.4732
R955 VTAIL.n280 VTAIL.n279 10.4732
R956 VTAIL.n230 VTAIL.n229 10.4732
R957 VTAIL.n180 VTAIL.n179 10.4732
R958 VTAIL.n374 VTAIL.n360 9.69747
R959 VTAIL.n24 VTAIL.n10 9.69747
R960 VTAIL.n74 VTAIL.n60 9.69747
R961 VTAIL.n124 VTAIL.n110 9.69747
R962 VTAIL.n326 VTAIL.n312 9.69747
R963 VTAIL.n276 VTAIL.n262 9.69747
R964 VTAIL.n226 VTAIL.n212 9.69747
R965 VTAIL.n176 VTAIL.n162 9.69747
R966 VTAIL.n398 VTAIL.n397 9.45567
R967 VTAIL.n48 VTAIL.n47 9.45567
R968 VTAIL.n98 VTAIL.n97 9.45567
R969 VTAIL.n148 VTAIL.n147 9.45567
R970 VTAIL.n348 VTAIL.n347 9.45567
R971 VTAIL.n298 VTAIL.n297 9.45567
R972 VTAIL.n248 VTAIL.n247 9.45567
R973 VTAIL.n198 VTAIL.n197 9.45567
R974 VTAIL.n397 VTAIL.n396 9.3005
R975 VTAIL.n352 VTAIL.n351 9.3005
R976 VTAIL.n391 VTAIL.n390 9.3005
R977 VTAIL.n364 VTAIL.n363 9.3005
R978 VTAIL.n371 VTAIL.n370 9.3005
R979 VTAIL.n373 VTAIL.n372 9.3005
R980 VTAIL.n360 VTAIL.n359 9.3005
R981 VTAIL.n379 VTAIL.n378 9.3005
R982 VTAIL.n381 VTAIL.n380 9.3005
R983 VTAIL.n382 VTAIL.n355 9.3005
R984 VTAIL.n389 VTAIL.n388 9.3005
R985 VTAIL.n47 VTAIL.n46 9.3005
R986 VTAIL.n2 VTAIL.n1 9.3005
R987 VTAIL.n41 VTAIL.n40 9.3005
R988 VTAIL.n14 VTAIL.n13 9.3005
R989 VTAIL.n21 VTAIL.n20 9.3005
R990 VTAIL.n23 VTAIL.n22 9.3005
R991 VTAIL.n10 VTAIL.n9 9.3005
R992 VTAIL.n29 VTAIL.n28 9.3005
R993 VTAIL.n31 VTAIL.n30 9.3005
R994 VTAIL.n32 VTAIL.n5 9.3005
R995 VTAIL.n39 VTAIL.n38 9.3005
R996 VTAIL.n97 VTAIL.n96 9.3005
R997 VTAIL.n52 VTAIL.n51 9.3005
R998 VTAIL.n91 VTAIL.n90 9.3005
R999 VTAIL.n64 VTAIL.n63 9.3005
R1000 VTAIL.n71 VTAIL.n70 9.3005
R1001 VTAIL.n73 VTAIL.n72 9.3005
R1002 VTAIL.n60 VTAIL.n59 9.3005
R1003 VTAIL.n79 VTAIL.n78 9.3005
R1004 VTAIL.n81 VTAIL.n80 9.3005
R1005 VTAIL.n82 VTAIL.n55 9.3005
R1006 VTAIL.n89 VTAIL.n88 9.3005
R1007 VTAIL.n147 VTAIL.n146 9.3005
R1008 VTAIL.n102 VTAIL.n101 9.3005
R1009 VTAIL.n141 VTAIL.n140 9.3005
R1010 VTAIL.n114 VTAIL.n113 9.3005
R1011 VTAIL.n121 VTAIL.n120 9.3005
R1012 VTAIL.n123 VTAIL.n122 9.3005
R1013 VTAIL.n110 VTAIL.n109 9.3005
R1014 VTAIL.n129 VTAIL.n128 9.3005
R1015 VTAIL.n131 VTAIL.n130 9.3005
R1016 VTAIL.n132 VTAIL.n105 9.3005
R1017 VTAIL.n139 VTAIL.n138 9.3005
R1018 VTAIL.n316 VTAIL.n315 9.3005
R1019 VTAIL.n323 VTAIL.n322 9.3005
R1020 VTAIL.n325 VTAIL.n324 9.3005
R1021 VTAIL.n312 VTAIL.n311 9.3005
R1022 VTAIL.n331 VTAIL.n330 9.3005
R1023 VTAIL.n333 VTAIL.n332 9.3005
R1024 VTAIL.n307 VTAIL.n305 9.3005
R1025 VTAIL.n339 VTAIL.n338 9.3005
R1026 VTAIL.n347 VTAIL.n346 9.3005
R1027 VTAIL.n302 VTAIL.n301 9.3005
R1028 VTAIL.n341 VTAIL.n340 9.3005
R1029 VTAIL.n266 VTAIL.n265 9.3005
R1030 VTAIL.n273 VTAIL.n272 9.3005
R1031 VTAIL.n275 VTAIL.n274 9.3005
R1032 VTAIL.n262 VTAIL.n261 9.3005
R1033 VTAIL.n281 VTAIL.n280 9.3005
R1034 VTAIL.n283 VTAIL.n282 9.3005
R1035 VTAIL.n257 VTAIL.n255 9.3005
R1036 VTAIL.n289 VTAIL.n288 9.3005
R1037 VTAIL.n297 VTAIL.n296 9.3005
R1038 VTAIL.n252 VTAIL.n251 9.3005
R1039 VTAIL.n291 VTAIL.n290 9.3005
R1040 VTAIL.n216 VTAIL.n215 9.3005
R1041 VTAIL.n223 VTAIL.n222 9.3005
R1042 VTAIL.n225 VTAIL.n224 9.3005
R1043 VTAIL.n212 VTAIL.n211 9.3005
R1044 VTAIL.n231 VTAIL.n230 9.3005
R1045 VTAIL.n233 VTAIL.n232 9.3005
R1046 VTAIL.n207 VTAIL.n205 9.3005
R1047 VTAIL.n239 VTAIL.n238 9.3005
R1048 VTAIL.n247 VTAIL.n246 9.3005
R1049 VTAIL.n202 VTAIL.n201 9.3005
R1050 VTAIL.n241 VTAIL.n240 9.3005
R1051 VTAIL.n166 VTAIL.n165 9.3005
R1052 VTAIL.n173 VTAIL.n172 9.3005
R1053 VTAIL.n175 VTAIL.n174 9.3005
R1054 VTAIL.n162 VTAIL.n161 9.3005
R1055 VTAIL.n181 VTAIL.n180 9.3005
R1056 VTAIL.n183 VTAIL.n182 9.3005
R1057 VTAIL.n157 VTAIL.n155 9.3005
R1058 VTAIL.n189 VTAIL.n188 9.3005
R1059 VTAIL.n197 VTAIL.n196 9.3005
R1060 VTAIL.n152 VTAIL.n151 9.3005
R1061 VTAIL.n191 VTAIL.n190 9.3005
R1062 VTAIL.n373 VTAIL.n362 8.92171
R1063 VTAIL.n23 VTAIL.n12 8.92171
R1064 VTAIL.n73 VTAIL.n62 8.92171
R1065 VTAIL.n123 VTAIL.n112 8.92171
R1066 VTAIL.n325 VTAIL.n314 8.92171
R1067 VTAIL.n275 VTAIL.n264 8.92171
R1068 VTAIL.n225 VTAIL.n214 8.92171
R1069 VTAIL.n175 VTAIL.n164 8.92171
R1070 VTAIL.n370 VTAIL.n369 8.14595
R1071 VTAIL.n20 VTAIL.n19 8.14595
R1072 VTAIL.n70 VTAIL.n69 8.14595
R1073 VTAIL.n120 VTAIL.n119 8.14595
R1074 VTAIL.n322 VTAIL.n321 8.14595
R1075 VTAIL.n272 VTAIL.n271 8.14595
R1076 VTAIL.n222 VTAIL.n221 8.14595
R1077 VTAIL.n172 VTAIL.n171 8.14595
R1078 VTAIL.n366 VTAIL.n364 7.3702
R1079 VTAIL.n16 VTAIL.n14 7.3702
R1080 VTAIL.n66 VTAIL.n64 7.3702
R1081 VTAIL.n116 VTAIL.n114 7.3702
R1082 VTAIL.n318 VTAIL.n316 7.3702
R1083 VTAIL.n268 VTAIL.n266 7.3702
R1084 VTAIL.n218 VTAIL.n216 7.3702
R1085 VTAIL.n168 VTAIL.n166 7.3702
R1086 VTAIL.n369 VTAIL.n364 5.81868
R1087 VTAIL.n19 VTAIL.n14 5.81868
R1088 VTAIL.n69 VTAIL.n64 5.81868
R1089 VTAIL.n119 VTAIL.n114 5.81868
R1090 VTAIL.n321 VTAIL.n316 5.81868
R1091 VTAIL.n271 VTAIL.n266 5.81868
R1092 VTAIL.n221 VTAIL.n216 5.81868
R1093 VTAIL.n171 VTAIL.n166 5.81868
R1094 VTAIL.n370 VTAIL.n362 5.04292
R1095 VTAIL.n20 VTAIL.n12 5.04292
R1096 VTAIL.n70 VTAIL.n62 5.04292
R1097 VTAIL.n120 VTAIL.n112 5.04292
R1098 VTAIL.n322 VTAIL.n314 5.04292
R1099 VTAIL.n272 VTAIL.n264 5.04292
R1100 VTAIL.n222 VTAIL.n214 5.04292
R1101 VTAIL.n172 VTAIL.n164 5.04292
R1102 VTAIL.n374 VTAIL.n373 4.26717
R1103 VTAIL.n24 VTAIL.n23 4.26717
R1104 VTAIL.n74 VTAIL.n73 4.26717
R1105 VTAIL.n124 VTAIL.n123 4.26717
R1106 VTAIL.n326 VTAIL.n325 4.26717
R1107 VTAIL.n276 VTAIL.n275 4.26717
R1108 VTAIL.n226 VTAIL.n225 4.26717
R1109 VTAIL.n176 VTAIL.n175 4.26717
R1110 VTAIL.n377 VTAIL.n360 3.49141
R1111 VTAIL.n27 VTAIL.n10 3.49141
R1112 VTAIL.n77 VTAIL.n60 3.49141
R1113 VTAIL.n127 VTAIL.n110 3.49141
R1114 VTAIL.n329 VTAIL.n312 3.49141
R1115 VTAIL.n279 VTAIL.n262 3.49141
R1116 VTAIL.n229 VTAIL.n212 3.49141
R1117 VTAIL.n179 VTAIL.n162 3.49141
R1118 VTAIL.n378 VTAIL.n358 2.71565
R1119 VTAIL.n398 VTAIL.n350 2.71565
R1120 VTAIL.n28 VTAIL.n8 2.71565
R1121 VTAIL.n48 VTAIL.n0 2.71565
R1122 VTAIL.n78 VTAIL.n58 2.71565
R1123 VTAIL.n98 VTAIL.n50 2.71565
R1124 VTAIL.n128 VTAIL.n108 2.71565
R1125 VTAIL.n148 VTAIL.n100 2.71565
R1126 VTAIL.n348 VTAIL.n300 2.71565
R1127 VTAIL.n330 VTAIL.n310 2.71565
R1128 VTAIL.n298 VTAIL.n250 2.71565
R1129 VTAIL.n280 VTAIL.n260 2.71565
R1130 VTAIL.n248 VTAIL.n200 2.71565
R1131 VTAIL.n230 VTAIL.n210 2.71565
R1132 VTAIL.n198 VTAIL.n150 2.71565
R1133 VTAIL.n180 VTAIL.n160 2.71565
R1134 VTAIL.n365 VTAIL.n363 2.41283
R1135 VTAIL.n15 VTAIL.n13 2.41283
R1136 VTAIL.n65 VTAIL.n63 2.41283
R1137 VTAIL.n115 VTAIL.n113 2.41283
R1138 VTAIL.n317 VTAIL.n315 2.41283
R1139 VTAIL.n267 VTAIL.n265 2.41283
R1140 VTAIL.n217 VTAIL.n215 2.41283
R1141 VTAIL.n167 VTAIL.n165 2.41283
R1142 VTAIL.n383 VTAIL.n381 1.93989
R1143 VTAIL.n396 VTAIL.n395 1.93989
R1144 VTAIL.n33 VTAIL.n31 1.93989
R1145 VTAIL.n46 VTAIL.n45 1.93989
R1146 VTAIL.n83 VTAIL.n81 1.93989
R1147 VTAIL.n96 VTAIL.n95 1.93989
R1148 VTAIL.n133 VTAIL.n131 1.93989
R1149 VTAIL.n146 VTAIL.n145 1.93989
R1150 VTAIL.n346 VTAIL.n345 1.93989
R1151 VTAIL.n334 VTAIL.n333 1.93989
R1152 VTAIL.n296 VTAIL.n295 1.93989
R1153 VTAIL.n284 VTAIL.n283 1.93989
R1154 VTAIL.n246 VTAIL.n245 1.93989
R1155 VTAIL.n234 VTAIL.n233 1.93989
R1156 VTAIL.n196 VTAIL.n195 1.93989
R1157 VTAIL.n184 VTAIL.n183 1.93989
R1158 VTAIL.n382 VTAIL.n356 1.16414
R1159 VTAIL.n392 VTAIL.n352 1.16414
R1160 VTAIL.n32 VTAIL.n6 1.16414
R1161 VTAIL.n42 VTAIL.n2 1.16414
R1162 VTAIL.n82 VTAIL.n56 1.16414
R1163 VTAIL.n92 VTAIL.n52 1.16414
R1164 VTAIL.n132 VTAIL.n106 1.16414
R1165 VTAIL.n142 VTAIL.n102 1.16414
R1166 VTAIL.n342 VTAIL.n302 1.16414
R1167 VTAIL.n337 VTAIL.n307 1.16414
R1168 VTAIL.n292 VTAIL.n252 1.16414
R1169 VTAIL.n287 VTAIL.n257 1.16414
R1170 VTAIL.n242 VTAIL.n202 1.16414
R1171 VTAIL.n237 VTAIL.n207 1.16414
R1172 VTAIL.n192 VTAIL.n152 1.16414
R1173 VTAIL.n187 VTAIL.n157 1.16414
R1174 VTAIL.n249 VTAIL.n199 0.560845
R1175 VTAIL.n349 VTAIL.n299 0.560845
R1176 VTAIL.n149 VTAIL.n99 0.560845
R1177 VTAIL.n299 VTAIL.n249 0.470328
R1178 VTAIL.n99 VTAIL.n49 0.470328
R1179 VTAIL.n388 VTAIL.n387 0.388379
R1180 VTAIL.n391 VTAIL.n354 0.388379
R1181 VTAIL.n38 VTAIL.n37 0.388379
R1182 VTAIL.n41 VTAIL.n4 0.388379
R1183 VTAIL.n88 VTAIL.n87 0.388379
R1184 VTAIL.n91 VTAIL.n54 0.388379
R1185 VTAIL.n138 VTAIL.n137 0.388379
R1186 VTAIL.n141 VTAIL.n104 0.388379
R1187 VTAIL.n341 VTAIL.n304 0.388379
R1188 VTAIL.n338 VTAIL.n306 0.388379
R1189 VTAIL.n291 VTAIL.n254 0.388379
R1190 VTAIL.n288 VTAIL.n256 0.388379
R1191 VTAIL.n241 VTAIL.n204 0.388379
R1192 VTAIL.n238 VTAIL.n206 0.388379
R1193 VTAIL.n191 VTAIL.n154 0.388379
R1194 VTAIL.n188 VTAIL.n156 0.388379
R1195 VTAIL VTAIL.n49 0.338862
R1196 VTAIL VTAIL.n399 0.222483
R1197 VTAIL.n371 VTAIL.n363 0.155672
R1198 VTAIL.n372 VTAIL.n371 0.155672
R1199 VTAIL.n372 VTAIL.n359 0.155672
R1200 VTAIL.n379 VTAIL.n359 0.155672
R1201 VTAIL.n380 VTAIL.n379 0.155672
R1202 VTAIL.n380 VTAIL.n355 0.155672
R1203 VTAIL.n389 VTAIL.n355 0.155672
R1204 VTAIL.n390 VTAIL.n389 0.155672
R1205 VTAIL.n390 VTAIL.n351 0.155672
R1206 VTAIL.n397 VTAIL.n351 0.155672
R1207 VTAIL.n21 VTAIL.n13 0.155672
R1208 VTAIL.n22 VTAIL.n21 0.155672
R1209 VTAIL.n22 VTAIL.n9 0.155672
R1210 VTAIL.n29 VTAIL.n9 0.155672
R1211 VTAIL.n30 VTAIL.n29 0.155672
R1212 VTAIL.n30 VTAIL.n5 0.155672
R1213 VTAIL.n39 VTAIL.n5 0.155672
R1214 VTAIL.n40 VTAIL.n39 0.155672
R1215 VTAIL.n40 VTAIL.n1 0.155672
R1216 VTAIL.n47 VTAIL.n1 0.155672
R1217 VTAIL.n71 VTAIL.n63 0.155672
R1218 VTAIL.n72 VTAIL.n71 0.155672
R1219 VTAIL.n72 VTAIL.n59 0.155672
R1220 VTAIL.n79 VTAIL.n59 0.155672
R1221 VTAIL.n80 VTAIL.n79 0.155672
R1222 VTAIL.n80 VTAIL.n55 0.155672
R1223 VTAIL.n89 VTAIL.n55 0.155672
R1224 VTAIL.n90 VTAIL.n89 0.155672
R1225 VTAIL.n90 VTAIL.n51 0.155672
R1226 VTAIL.n97 VTAIL.n51 0.155672
R1227 VTAIL.n121 VTAIL.n113 0.155672
R1228 VTAIL.n122 VTAIL.n121 0.155672
R1229 VTAIL.n122 VTAIL.n109 0.155672
R1230 VTAIL.n129 VTAIL.n109 0.155672
R1231 VTAIL.n130 VTAIL.n129 0.155672
R1232 VTAIL.n130 VTAIL.n105 0.155672
R1233 VTAIL.n139 VTAIL.n105 0.155672
R1234 VTAIL.n140 VTAIL.n139 0.155672
R1235 VTAIL.n140 VTAIL.n101 0.155672
R1236 VTAIL.n147 VTAIL.n101 0.155672
R1237 VTAIL.n347 VTAIL.n301 0.155672
R1238 VTAIL.n340 VTAIL.n301 0.155672
R1239 VTAIL.n340 VTAIL.n339 0.155672
R1240 VTAIL.n339 VTAIL.n305 0.155672
R1241 VTAIL.n332 VTAIL.n305 0.155672
R1242 VTAIL.n332 VTAIL.n331 0.155672
R1243 VTAIL.n331 VTAIL.n311 0.155672
R1244 VTAIL.n324 VTAIL.n311 0.155672
R1245 VTAIL.n324 VTAIL.n323 0.155672
R1246 VTAIL.n323 VTAIL.n315 0.155672
R1247 VTAIL.n297 VTAIL.n251 0.155672
R1248 VTAIL.n290 VTAIL.n251 0.155672
R1249 VTAIL.n290 VTAIL.n289 0.155672
R1250 VTAIL.n289 VTAIL.n255 0.155672
R1251 VTAIL.n282 VTAIL.n255 0.155672
R1252 VTAIL.n282 VTAIL.n281 0.155672
R1253 VTAIL.n281 VTAIL.n261 0.155672
R1254 VTAIL.n274 VTAIL.n261 0.155672
R1255 VTAIL.n274 VTAIL.n273 0.155672
R1256 VTAIL.n273 VTAIL.n265 0.155672
R1257 VTAIL.n247 VTAIL.n201 0.155672
R1258 VTAIL.n240 VTAIL.n201 0.155672
R1259 VTAIL.n240 VTAIL.n239 0.155672
R1260 VTAIL.n239 VTAIL.n205 0.155672
R1261 VTAIL.n232 VTAIL.n205 0.155672
R1262 VTAIL.n232 VTAIL.n231 0.155672
R1263 VTAIL.n231 VTAIL.n211 0.155672
R1264 VTAIL.n224 VTAIL.n211 0.155672
R1265 VTAIL.n224 VTAIL.n223 0.155672
R1266 VTAIL.n223 VTAIL.n215 0.155672
R1267 VTAIL.n197 VTAIL.n151 0.155672
R1268 VTAIL.n190 VTAIL.n151 0.155672
R1269 VTAIL.n190 VTAIL.n189 0.155672
R1270 VTAIL.n189 VTAIL.n155 0.155672
R1271 VTAIL.n182 VTAIL.n155 0.155672
R1272 VTAIL.n182 VTAIL.n181 0.155672
R1273 VTAIL.n181 VTAIL.n161 0.155672
R1274 VTAIL.n174 VTAIL.n161 0.155672
R1275 VTAIL.n174 VTAIL.n173 0.155672
R1276 VTAIL.n173 VTAIL.n165 0.155672
R1277 VDD1 VDD1.n1 112.484
R1278 VDD1 VDD1.n0 78.6389
R1279 VDD1.n0 VDD1.t2 3.51836
R1280 VDD1.n0 VDD1.t3 3.51836
R1281 VDD1.n1 VDD1.t0 3.51836
R1282 VDD1.n1 VDD1.t1 3.51836
R1283 VN.n0 VN.t1 842.77
R1284 VN.n0 VN.t0 842.77
R1285 VN.n1 VN.t2 842.77
R1286 VN.n1 VN.t3 842.77
R1287 VN VN.n1 198.953
R1288 VN VN.n0 161.351
R1289 VDD2.n2 VDD2.n0 111.96
R1290 VDD2.n2 VDD2.n1 78.5807
R1291 VDD2.n1 VDD2.t1 3.51836
R1292 VDD2.n1 VDD2.t0 3.51836
R1293 VDD2.n0 VDD2.t3 3.51836
R1294 VDD2.n0 VDD2.t2 3.51836
R1295 VDD2 VDD2.n2 0.0586897
C0 VDD2 w_n1360_n2820# 0.906202f
C1 B w_n1360_n2820# 5.67726f
C2 VP VDD1 1.81828f
C3 VN VTAIL 1.31937f
C4 VDD2 VDD1 0.482688f
C5 B VDD1 0.784329f
C6 VP VDD2 0.250032f
C7 VP B 0.907487f
C8 VN w_n1360_n2820# 1.83198f
C9 B VDD2 0.800606f
C10 VTAIL w_n1360_n2820# 3.5183f
C11 VN VDD1 0.147746f
C12 VN VP 4.03276f
C13 VN VDD2 1.71616f
C14 VN B 0.637539f
C15 VTAIL VDD1 7.37754f
C16 VTAIL VP 1.33347f
C17 VTAIL VDD2 7.41646f
C18 VTAIL B 2.83281f
C19 VDD1 w_n1360_n2820# 0.899004f
C20 VP w_n1360_n2820# 2.00105f
C21 VDD2 VSUBS 0.552299f
C22 VDD1 VSUBS 4.027284f
C23 VTAIL VSUBS 0.643667f
C24 VN VSUBS 3.64519f
C25 VP VSUBS 0.995225f
C26 B VSUBS 2.063126f
C27 w_n1360_n2820# VSUBS 47.4422f
C28 VDD2.t3 VSUBS 0.190673f
C29 VDD2.t2 VSUBS 0.190673f
C30 VDD2.n0 VSUBS 1.88225f
C31 VDD2.t1 VSUBS 0.190673f
C32 VDD2.t0 VSUBS 0.190673f
C33 VDD2.n1 VSUBS 1.41738f
C34 VDD2.n2 VSUBS 3.28491f
C35 VN.t0 VSUBS 0.289446f
C36 VN.t1 VSUBS 0.289446f
C37 VN.n0 VSUBS 0.240566f
C38 VN.t2 VSUBS 0.289446f
C39 VN.t3 VSUBS 0.289446f
C40 VN.n1 VSUBS 0.460616f
C41 VDD1.t2 VSUBS 0.18822f
C42 VDD1.t3 VSUBS 0.18822f
C43 VDD1.n0 VSUBS 1.39953f
C44 VDD1.t0 VSUBS 0.18822f
C45 VDD1.t1 VSUBS 0.18822f
C46 VDD1.n1 VSUBS 1.879f
C47 VTAIL.n0 VSUBS 0.023819f
C48 VTAIL.n1 VSUBS 0.023198f
C49 VTAIL.n2 VSUBS 0.012466f
C50 VTAIL.n3 VSUBS 0.029464f
C51 VTAIL.n4 VSUBS 0.012832f
C52 VTAIL.n5 VSUBS 0.023198f
C53 VTAIL.n6 VSUBS 0.013199f
C54 VTAIL.n7 VSUBS 0.029464f
C55 VTAIL.n8 VSUBS 0.013199f
C56 VTAIL.n9 VSUBS 0.023198f
C57 VTAIL.n10 VSUBS 0.012466f
C58 VTAIL.n11 VSUBS 0.029464f
C59 VTAIL.n12 VSUBS 0.013199f
C60 VTAIL.n13 VSUBS 0.859206f
C61 VTAIL.n14 VSUBS 0.012466f
C62 VTAIL.t2 VSUBS 0.063303f
C63 VTAIL.n15 VSUBS 0.153772f
C64 VTAIL.n16 VSUBS 0.022165f
C65 VTAIL.n17 VSUBS 0.022098f
C66 VTAIL.n18 VSUBS 0.029464f
C67 VTAIL.n19 VSUBS 0.013199f
C68 VTAIL.n20 VSUBS 0.012466f
C69 VTAIL.n21 VSUBS 0.023198f
C70 VTAIL.n22 VSUBS 0.023198f
C71 VTAIL.n23 VSUBS 0.012466f
C72 VTAIL.n24 VSUBS 0.013199f
C73 VTAIL.n25 VSUBS 0.029464f
C74 VTAIL.n26 VSUBS 0.029464f
C75 VTAIL.n27 VSUBS 0.013199f
C76 VTAIL.n28 VSUBS 0.012466f
C77 VTAIL.n29 VSUBS 0.023198f
C78 VTAIL.n30 VSUBS 0.023198f
C79 VTAIL.n31 VSUBS 0.012466f
C80 VTAIL.n32 VSUBS 0.012466f
C81 VTAIL.n33 VSUBS 0.013199f
C82 VTAIL.n34 VSUBS 0.029464f
C83 VTAIL.n35 VSUBS 0.029464f
C84 VTAIL.n36 VSUBS 0.029464f
C85 VTAIL.n37 VSUBS 0.012832f
C86 VTAIL.n38 VSUBS 0.012466f
C87 VTAIL.n39 VSUBS 0.023198f
C88 VTAIL.n40 VSUBS 0.023198f
C89 VTAIL.n41 VSUBS 0.012466f
C90 VTAIL.n42 VSUBS 0.013199f
C91 VTAIL.n43 VSUBS 0.029464f
C92 VTAIL.n44 VSUBS 0.06564f
C93 VTAIL.n45 VSUBS 0.013199f
C94 VTAIL.n46 VSUBS 0.012466f
C95 VTAIL.n47 VSUBS 0.053621f
C96 VTAIL.n48 VSUBS 0.032757f
C97 VTAIL.n49 VSUBS 0.080225f
C98 VTAIL.n50 VSUBS 0.023819f
C99 VTAIL.n51 VSUBS 0.023198f
C100 VTAIL.n52 VSUBS 0.012466f
C101 VTAIL.n53 VSUBS 0.029464f
C102 VTAIL.n54 VSUBS 0.012832f
C103 VTAIL.n55 VSUBS 0.023198f
C104 VTAIL.n56 VSUBS 0.013199f
C105 VTAIL.n57 VSUBS 0.029464f
C106 VTAIL.n58 VSUBS 0.013199f
C107 VTAIL.n59 VSUBS 0.023198f
C108 VTAIL.n60 VSUBS 0.012466f
C109 VTAIL.n61 VSUBS 0.029464f
C110 VTAIL.n62 VSUBS 0.013199f
C111 VTAIL.n63 VSUBS 0.859206f
C112 VTAIL.n64 VSUBS 0.012466f
C113 VTAIL.t6 VSUBS 0.063303f
C114 VTAIL.n65 VSUBS 0.153772f
C115 VTAIL.n66 VSUBS 0.022165f
C116 VTAIL.n67 VSUBS 0.022098f
C117 VTAIL.n68 VSUBS 0.029464f
C118 VTAIL.n69 VSUBS 0.013199f
C119 VTAIL.n70 VSUBS 0.012466f
C120 VTAIL.n71 VSUBS 0.023198f
C121 VTAIL.n72 VSUBS 0.023198f
C122 VTAIL.n73 VSUBS 0.012466f
C123 VTAIL.n74 VSUBS 0.013199f
C124 VTAIL.n75 VSUBS 0.029464f
C125 VTAIL.n76 VSUBS 0.029464f
C126 VTAIL.n77 VSUBS 0.013199f
C127 VTAIL.n78 VSUBS 0.012466f
C128 VTAIL.n79 VSUBS 0.023198f
C129 VTAIL.n80 VSUBS 0.023198f
C130 VTAIL.n81 VSUBS 0.012466f
C131 VTAIL.n82 VSUBS 0.012466f
C132 VTAIL.n83 VSUBS 0.013199f
C133 VTAIL.n84 VSUBS 0.029464f
C134 VTAIL.n85 VSUBS 0.029464f
C135 VTAIL.n86 VSUBS 0.029464f
C136 VTAIL.n87 VSUBS 0.012832f
C137 VTAIL.n88 VSUBS 0.012466f
C138 VTAIL.n89 VSUBS 0.023198f
C139 VTAIL.n90 VSUBS 0.023198f
C140 VTAIL.n91 VSUBS 0.012466f
C141 VTAIL.n92 VSUBS 0.013199f
C142 VTAIL.n93 VSUBS 0.029464f
C143 VTAIL.n94 VSUBS 0.06564f
C144 VTAIL.n95 VSUBS 0.013199f
C145 VTAIL.n96 VSUBS 0.012466f
C146 VTAIL.n97 VSUBS 0.053621f
C147 VTAIL.n98 VSUBS 0.032757f
C148 VTAIL.n99 VSUBS 0.096818f
C149 VTAIL.n100 VSUBS 0.023819f
C150 VTAIL.n101 VSUBS 0.023198f
C151 VTAIL.n102 VSUBS 0.012466f
C152 VTAIL.n103 VSUBS 0.029464f
C153 VTAIL.n104 VSUBS 0.012832f
C154 VTAIL.n105 VSUBS 0.023198f
C155 VTAIL.n106 VSUBS 0.013199f
C156 VTAIL.n107 VSUBS 0.029464f
C157 VTAIL.n108 VSUBS 0.013199f
C158 VTAIL.n109 VSUBS 0.023198f
C159 VTAIL.n110 VSUBS 0.012466f
C160 VTAIL.n111 VSUBS 0.029464f
C161 VTAIL.n112 VSUBS 0.013199f
C162 VTAIL.n113 VSUBS 0.859206f
C163 VTAIL.n114 VSUBS 0.012466f
C164 VTAIL.t5 VSUBS 0.063303f
C165 VTAIL.n115 VSUBS 0.153772f
C166 VTAIL.n116 VSUBS 0.022165f
C167 VTAIL.n117 VSUBS 0.022098f
C168 VTAIL.n118 VSUBS 0.029464f
C169 VTAIL.n119 VSUBS 0.013199f
C170 VTAIL.n120 VSUBS 0.012466f
C171 VTAIL.n121 VSUBS 0.023198f
C172 VTAIL.n122 VSUBS 0.023198f
C173 VTAIL.n123 VSUBS 0.012466f
C174 VTAIL.n124 VSUBS 0.013199f
C175 VTAIL.n125 VSUBS 0.029464f
C176 VTAIL.n126 VSUBS 0.029464f
C177 VTAIL.n127 VSUBS 0.013199f
C178 VTAIL.n128 VSUBS 0.012466f
C179 VTAIL.n129 VSUBS 0.023198f
C180 VTAIL.n130 VSUBS 0.023198f
C181 VTAIL.n131 VSUBS 0.012466f
C182 VTAIL.n132 VSUBS 0.012466f
C183 VTAIL.n133 VSUBS 0.013199f
C184 VTAIL.n134 VSUBS 0.029464f
C185 VTAIL.n135 VSUBS 0.029464f
C186 VTAIL.n136 VSUBS 0.029464f
C187 VTAIL.n137 VSUBS 0.012832f
C188 VTAIL.n138 VSUBS 0.012466f
C189 VTAIL.n139 VSUBS 0.023198f
C190 VTAIL.n140 VSUBS 0.023198f
C191 VTAIL.n141 VSUBS 0.012466f
C192 VTAIL.n142 VSUBS 0.013199f
C193 VTAIL.n143 VSUBS 0.029464f
C194 VTAIL.n144 VSUBS 0.06564f
C195 VTAIL.n145 VSUBS 0.013199f
C196 VTAIL.n146 VSUBS 0.012466f
C197 VTAIL.n147 VSUBS 0.053621f
C198 VTAIL.n148 VSUBS 0.032757f
C199 VTAIL.n149 VSUBS 1.01541f
C200 VTAIL.n150 VSUBS 0.023819f
C201 VTAIL.n151 VSUBS 0.023198f
C202 VTAIL.n152 VSUBS 0.012466f
C203 VTAIL.n153 VSUBS 0.029464f
C204 VTAIL.n154 VSUBS 0.012832f
C205 VTAIL.n155 VSUBS 0.023198f
C206 VTAIL.n156 VSUBS 0.012832f
C207 VTAIL.n157 VSUBS 0.012466f
C208 VTAIL.n158 VSUBS 0.029464f
C209 VTAIL.n159 VSUBS 0.029464f
C210 VTAIL.n160 VSUBS 0.013199f
C211 VTAIL.n161 VSUBS 0.023198f
C212 VTAIL.n162 VSUBS 0.012466f
C213 VTAIL.n163 VSUBS 0.029464f
C214 VTAIL.n164 VSUBS 0.013199f
C215 VTAIL.n165 VSUBS 0.859206f
C216 VTAIL.n166 VSUBS 0.012466f
C217 VTAIL.t0 VSUBS 0.063303f
C218 VTAIL.n167 VSUBS 0.153772f
C219 VTAIL.n168 VSUBS 0.022165f
C220 VTAIL.n169 VSUBS 0.022098f
C221 VTAIL.n170 VSUBS 0.029464f
C222 VTAIL.n171 VSUBS 0.013199f
C223 VTAIL.n172 VSUBS 0.012466f
C224 VTAIL.n173 VSUBS 0.023198f
C225 VTAIL.n174 VSUBS 0.023198f
C226 VTAIL.n175 VSUBS 0.012466f
C227 VTAIL.n176 VSUBS 0.013199f
C228 VTAIL.n177 VSUBS 0.029464f
C229 VTAIL.n178 VSUBS 0.029464f
C230 VTAIL.n179 VSUBS 0.013199f
C231 VTAIL.n180 VSUBS 0.012466f
C232 VTAIL.n181 VSUBS 0.023198f
C233 VTAIL.n182 VSUBS 0.023198f
C234 VTAIL.n183 VSUBS 0.012466f
C235 VTAIL.n184 VSUBS 0.013199f
C236 VTAIL.n185 VSUBS 0.029464f
C237 VTAIL.n186 VSUBS 0.029464f
C238 VTAIL.n187 VSUBS 0.013199f
C239 VTAIL.n188 VSUBS 0.012466f
C240 VTAIL.n189 VSUBS 0.023198f
C241 VTAIL.n190 VSUBS 0.023198f
C242 VTAIL.n191 VSUBS 0.012466f
C243 VTAIL.n192 VSUBS 0.013199f
C244 VTAIL.n193 VSUBS 0.029464f
C245 VTAIL.n194 VSUBS 0.06564f
C246 VTAIL.n195 VSUBS 0.013199f
C247 VTAIL.n196 VSUBS 0.012466f
C248 VTAIL.n197 VSUBS 0.053621f
C249 VTAIL.n198 VSUBS 0.032757f
C250 VTAIL.n199 VSUBS 1.01541f
C251 VTAIL.n200 VSUBS 0.023819f
C252 VTAIL.n201 VSUBS 0.023198f
C253 VTAIL.n202 VSUBS 0.012466f
C254 VTAIL.n203 VSUBS 0.029464f
C255 VTAIL.n204 VSUBS 0.012832f
C256 VTAIL.n205 VSUBS 0.023198f
C257 VTAIL.n206 VSUBS 0.012832f
C258 VTAIL.n207 VSUBS 0.012466f
C259 VTAIL.n208 VSUBS 0.029464f
C260 VTAIL.n209 VSUBS 0.029464f
C261 VTAIL.n210 VSUBS 0.013199f
C262 VTAIL.n211 VSUBS 0.023198f
C263 VTAIL.n212 VSUBS 0.012466f
C264 VTAIL.n213 VSUBS 0.029464f
C265 VTAIL.n214 VSUBS 0.013199f
C266 VTAIL.n215 VSUBS 0.859206f
C267 VTAIL.n216 VSUBS 0.012466f
C268 VTAIL.t3 VSUBS 0.063303f
C269 VTAIL.n217 VSUBS 0.153772f
C270 VTAIL.n218 VSUBS 0.022165f
C271 VTAIL.n219 VSUBS 0.022098f
C272 VTAIL.n220 VSUBS 0.029464f
C273 VTAIL.n221 VSUBS 0.013199f
C274 VTAIL.n222 VSUBS 0.012466f
C275 VTAIL.n223 VSUBS 0.023198f
C276 VTAIL.n224 VSUBS 0.023198f
C277 VTAIL.n225 VSUBS 0.012466f
C278 VTAIL.n226 VSUBS 0.013199f
C279 VTAIL.n227 VSUBS 0.029464f
C280 VTAIL.n228 VSUBS 0.029464f
C281 VTAIL.n229 VSUBS 0.013199f
C282 VTAIL.n230 VSUBS 0.012466f
C283 VTAIL.n231 VSUBS 0.023198f
C284 VTAIL.n232 VSUBS 0.023198f
C285 VTAIL.n233 VSUBS 0.012466f
C286 VTAIL.n234 VSUBS 0.013199f
C287 VTAIL.n235 VSUBS 0.029464f
C288 VTAIL.n236 VSUBS 0.029464f
C289 VTAIL.n237 VSUBS 0.013199f
C290 VTAIL.n238 VSUBS 0.012466f
C291 VTAIL.n239 VSUBS 0.023198f
C292 VTAIL.n240 VSUBS 0.023198f
C293 VTAIL.n241 VSUBS 0.012466f
C294 VTAIL.n242 VSUBS 0.013199f
C295 VTAIL.n243 VSUBS 0.029464f
C296 VTAIL.n244 VSUBS 0.06564f
C297 VTAIL.n245 VSUBS 0.013199f
C298 VTAIL.n246 VSUBS 0.012466f
C299 VTAIL.n247 VSUBS 0.053621f
C300 VTAIL.n248 VSUBS 0.032757f
C301 VTAIL.n249 VSUBS 0.096818f
C302 VTAIL.n250 VSUBS 0.023819f
C303 VTAIL.n251 VSUBS 0.023198f
C304 VTAIL.n252 VSUBS 0.012466f
C305 VTAIL.n253 VSUBS 0.029464f
C306 VTAIL.n254 VSUBS 0.012832f
C307 VTAIL.n255 VSUBS 0.023198f
C308 VTAIL.n256 VSUBS 0.012832f
C309 VTAIL.n257 VSUBS 0.012466f
C310 VTAIL.n258 VSUBS 0.029464f
C311 VTAIL.n259 VSUBS 0.029464f
C312 VTAIL.n260 VSUBS 0.013199f
C313 VTAIL.n261 VSUBS 0.023198f
C314 VTAIL.n262 VSUBS 0.012466f
C315 VTAIL.n263 VSUBS 0.029464f
C316 VTAIL.n264 VSUBS 0.013199f
C317 VTAIL.n265 VSUBS 0.859206f
C318 VTAIL.n266 VSUBS 0.012466f
C319 VTAIL.t4 VSUBS 0.063303f
C320 VTAIL.n267 VSUBS 0.153772f
C321 VTAIL.n268 VSUBS 0.022165f
C322 VTAIL.n269 VSUBS 0.022098f
C323 VTAIL.n270 VSUBS 0.029464f
C324 VTAIL.n271 VSUBS 0.013199f
C325 VTAIL.n272 VSUBS 0.012466f
C326 VTAIL.n273 VSUBS 0.023198f
C327 VTAIL.n274 VSUBS 0.023198f
C328 VTAIL.n275 VSUBS 0.012466f
C329 VTAIL.n276 VSUBS 0.013199f
C330 VTAIL.n277 VSUBS 0.029464f
C331 VTAIL.n278 VSUBS 0.029464f
C332 VTAIL.n279 VSUBS 0.013199f
C333 VTAIL.n280 VSUBS 0.012466f
C334 VTAIL.n281 VSUBS 0.023198f
C335 VTAIL.n282 VSUBS 0.023198f
C336 VTAIL.n283 VSUBS 0.012466f
C337 VTAIL.n284 VSUBS 0.013199f
C338 VTAIL.n285 VSUBS 0.029464f
C339 VTAIL.n286 VSUBS 0.029464f
C340 VTAIL.n287 VSUBS 0.013199f
C341 VTAIL.n288 VSUBS 0.012466f
C342 VTAIL.n289 VSUBS 0.023198f
C343 VTAIL.n290 VSUBS 0.023198f
C344 VTAIL.n291 VSUBS 0.012466f
C345 VTAIL.n292 VSUBS 0.013199f
C346 VTAIL.n293 VSUBS 0.029464f
C347 VTAIL.n294 VSUBS 0.06564f
C348 VTAIL.n295 VSUBS 0.013199f
C349 VTAIL.n296 VSUBS 0.012466f
C350 VTAIL.n297 VSUBS 0.053621f
C351 VTAIL.n298 VSUBS 0.032757f
C352 VTAIL.n299 VSUBS 0.096818f
C353 VTAIL.n300 VSUBS 0.023819f
C354 VTAIL.n301 VSUBS 0.023198f
C355 VTAIL.n302 VSUBS 0.012466f
C356 VTAIL.n303 VSUBS 0.029464f
C357 VTAIL.n304 VSUBS 0.012832f
C358 VTAIL.n305 VSUBS 0.023198f
C359 VTAIL.n306 VSUBS 0.012832f
C360 VTAIL.n307 VSUBS 0.012466f
C361 VTAIL.n308 VSUBS 0.029464f
C362 VTAIL.n309 VSUBS 0.029464f
C363 VTAIL.n310 VSUBS 0.013199f
C364 VTAIL.n311 VSUBS 0.023198f
C365 VTAIL.n312 VSUBS 0.012466f
C366 VTAIL.n313 VSUBS 0.029464f
C367 VTAIL.n314 VSUBS 0.013199f
C368 VTAIL.n315 VSUBS 0.859206f
C369 VTAIL.n316 VSUBS 0.012466f
C370 VTAIL.t7 VSUBS 0.063303f
C371 VTAIL.n317 VSUBS 0.153772f
C372 VTAIL.n318 VSUBS 0.022165f
C373 VTAIL.n319 VSUBS 0.022098f
C374 VTAIL.n320 VSUBS 0.029464f
C375 VTAIL.n321 VSUBS 0.013199f
C376 VTAIL.n322 VSUBS 0.012466f
C377 VTAIL.n323 VSUBS 0.023198f
C378 VTAIL.n324 VSUBS 0.023198f
C379 VTAIL.n325 VSUBS 0.012466f
C380 VTAIL.n326 VSUBS 0.013199f
C381 VTAIL.n327 VSUBS 0.029464f
C382 VTAIL.n328 VSUBS 0.029464f
C383 VTAIL.n329 VSUBS 0.013199f
C384 VTAIL.n330 VSUBS 0.012466f
C385 VTAIL.n331 VSUBS 0.023198f
C386 VTAIL.n332 VSUBS 0.023198f
C387 VTAIL.n333 VSUBS 0.012466f
C388 VTAIL.n334 VSUBS 0.013199f
C389 VTAIL.n335 VSUBS 0.029464f
C390 VTAIL.n336 VSUBS 0.029464f
C391 VTAIL.n337 VSUBS 0.013199f
C392 VTAIL.n338 VSUBS 0.012466f
C393 VTAIL.n339 VSUBS 0.023198f
C394 VTAIL.n340 VSUBS 0.023198f
C395 VTAIL.n341 VSUBS 0.012466f
C396 VTAIL.n342 VSUBS 0.013199f
C397 VTAIL.n343 VSUBS 0.029464f
C398 VTAIL.n344 VSUBS 0.06564f
C399 VTAIL.n345 VSUBS 0.013199f
C400 VTAIL.n346 VSUBS 0.012466f
C401 VTAIL.n347 VSUBS 0.053621f
C402 VTAIL.n348 VSUBS 0.032757f
C403 VTAIL.n349 VSUBS 1.01541f
C404 VTAIL.n350 VSUBS 0.023819f
C405 VTAIL.n351 VSUBS 0.023198f
C406 VTAIL.n352 VSUBS 0.012466f
C407 VTAIL.n353 VSUBS 0.029464f
C408 VTAIL.n354 VSUBS 0.012832f
C409 VTAIL.n355 VSUBS 0.023198f
C410 VTAIL.n356 VSUBS 0.013199f
C411 VTAIL.n357 VSUBS 0.029464f
C412 VTAIL.n358 VSUBS 0.013199f
C413 VTAIL.n359 VSUBS 0.023198f
C414 VTAIL.n360 VSUBS 0.012466f
C415 VTAIL.n361 VSUBS 0.029464f
C416 VTAIL.n362 VSUBS 0.013199f
C417 VTAIL.n363 VSUBS 0.859206f
C418 VTAIL.n364 VSUBS 0.012466f
C419 VTAIL.t1 VSUBS 0.063303f
C420 VTAIL.n365 VSUBS 0.153772f
C421 VTAIL.n366 VSUBS 0.022165f
C422 VTAIL.n367 VSUBS 0.022098f
C423 VTAIL.n368 VSUBS 0.029464f
C424 VTAIL.n369 VSUBS 0.013199f
C425 VTAIL.n370 VSUBS 0.012466f
C426 VTAIL.n371 VSUBS 0.023198f
C427 VTAIL.n372 VSUBS 0.023198f
C428 VTAIL.n373 VSUBS 0.012466f
C429 VTAIL.n374 VSUBS 0.013199f
C430 VTAIL.n375 VSUBS 0.029464f
C431 VTAIL.n376 VSUBS 0.029464f
C432 VTAIL.n377 VSUBS 0.013199f
C433 VTAIL.n378 VSUBS 0.012466f
C434 VTAIL.n379 VSUBS 0.023198f
C435 VTAIL.n380 VSUBS 0.023198f
C436 VTAIL.n381 VSUBS 0.012466f
C437 VTAIL.n382 VSUBS 0.012466f
C438 VTAIL.n383 VSUBS 0.013199f
C439 VTAIL.n384 VSUBS 0.029464f
C440 VTAIL.n385 VSUBS 0.029464f
C441 VTAIL.n386 VSUBS 0.029464f
C442 VTAIL.n387 VSUBS 0.012832f
C443 VTAIL.n388 VSUBS 0.012466f
C444 VTAIL.n389 VSUBS 0.023198f
C445 VTAIL.n390 VSUBS 0.023198f
C446 VTAIL.n391 VSUBS 0.012466f
C447 VTAIL.n392 VSUBS 0.013199f
C448 VTAIL.n393 VSUBS 0.029464f
C449 VTAIL.n394 VSUBS 0.06564f
C450 VTAIL.n395 VSUBS 0.013199f
C451 VTAIL.n396 VSUBS 0.012466f
C452 VTAIL.n397 VSUBS 0.053621f
C453 VTAIL.n398 VSUBS 0.032757f
C454 VTAIL.n399 VSUBS 0.990119f
C455 VP.t1 VSUBS 0.439377f
C456 VP.t0 VSUBS 0.439377f
C457 VP.n0 VSUBS 0.690109f
C458 VP.t3 VSUBS 0.439377f
C459 VP.t2 VSUBS 0.439377f
C460 VP.n1 VSUBS 0.36516f
C461 VP.n2 VSUBS 3.16086f
C462 B.n0 VSUBS 0.00571f
C463 B.n1 VSUBS 0.00571f
C464 B.n2 VSUBS 0.009029f
C465 B.n3 VSUBS 0.009029f
C466 B.n4 VSUBS 0.009029f
C467 B.n5 VSUBS 0.009029f
C468 B.n6 VSUBS 0.009029f
C469 B.n7 VSUBS 0.009029f
C470 B.n8 VSUBS 0.009029f
C471 B.n9 VSUBS 0.02022f
C472 B.n10 VSUBS 0.009029f
C473 B.n11 VSUBS 0.009029f
C474 B.n12 VSUBS 0.009029f
C475 B.n13 VSUBS 0.009029f
C476 B.n14 VSUBS 0.009029f
C477 B.n15 VSUBS 0.009029f
C478 B.n16 VSUBS 0.009029f
C479 B.n17 VSUBS 0.009029f
C480 B.n18 VSUBS 0.009029f
C481 B.n19 VSUBS 0.009029f
C482 B.n20 VSUBS 0.009029f
C483 B.n21 VSUBS 0.009029f
C484 B.n22 VSUBS 0.009029f
C485 B.n23 VSUBS 0.009029f
C486 B.n24 VSUBS 0.009029f
C487 B.n25 VSUBS 0.009029f
C488 B.t5 VSUBS 0.195368f
C489 B.t4 VSUBS 0.204603f
C490 B.t3 VSUBS 0.152047f
C491 B.n26 VSUBS 0.292141f
C492 B.n27 VSUBS 0.260779f
C493 B.n28 VSUBS 0.02092f
C494 B.n29 VSUBS 0.009029f
C495 B.n30 VSUBS 0.009029f
C496 B.n31 VSUBS 0.009029f
C497 B.n32 VSUBS 0.009029f
C498 B.n33 VSUBS 0.009029f
C499 B.t2 VSUBS 0.195372f
C500 B.t1 VSUBS 0.204606f
C501 B.t0 VSUBS 0.152047f
C502 B.n34 VSUBS 0.292138f
C503 B.n35 VSUBS 0.260775f
C504 B.n36 VSUBS 0.009029f
C505 B.n37 VSUBS 0.009029f
C506 B.n38 VSUBS 0.009029f
C507 B.n39 VSUBS 0.009029f
C508 B.n40 VSUBS 0.009029f
C509 B.n41 VSUBS 0.009029f
C510 B.n42 VSUBS 0.009029f
C511 B.n43 VSUBS 0.009029f
C512 B.n44 VSUBS 0.009029f
C513 B.n45 VSUBS 0.009029f
C514 B.n46 VSUBS 0.009029f
C515 B.n47 VSUBS 0.009029f
C516 B.n48 VSUBS 0.009029f
C517 B.n49 VSUBS 0.009029f
C518 B.n50 VSUBS 0.009029f
C519 B.n51 VSUBS 0.009029f
C520 B.n52 VSUBS 0.020278f
C521 B.n53 VSUBS 0.009029f
C522 B.n54 VSUBS 0.009029f
C523 B.n55 VSUBS 0.009029f
C524 B.n56 VSUBS 0.009029f
C525 B.n57 VSUBS 0.009029f
C526 B.n58 VSUBS 0.009029f
C527 B.n59 VSUBS 0.009029f
C528 B.n60 VSUBS 0.009029f
C529 B.n61 VSUBS 0.009029f
C530 B.n62 VSUBS 0.009029f
C531 B.n63 VSUBS 0.009029f
C532 B.n64 VSUBS 0.009029f
C533 B.n65 VSUBS 0.009029f
C534 B.n66 VSUBS 0.019085f
C535 B.n67 VSUBS 0.009029f
C536 B.n68 VSUBS 0.009029f
C537 B.n69 VSUBS 0.009029f
C538 B.n70 VSUBS 0.009029f
C539 B.n71 VSUBS 0.009029f
C540 B.n72 VSUBS 0.009029f
C541 B.n73 VSUBS 0.009029f
C542 B.n74 VSUBS 0.009029f
C543 B.n75 VSUBS 0.009029f
C544 B.n76 VSUBS 0.009029f
C545 B.n77 VSUBS 0.009029f
C546 B.n78 VSUBS 0.009029f
C547 B.n79 VSUBS 0.009029f
C548 B.n80 VSUBS 0.009029f
C549 B.n81 VSUBS 0.009029f
C550 B.n82 VSUBS 0.009029f
C551 B.n83 VSUBS 0.009029f
C552 B.t10 VSUBS 0.195372f
C553 B.t11 VSUBS 0.204606f
C554 B.t9 VSUBS 0.152047f
C555 B.n84 VSUBS 0.292138f
C556 B.n85 VSUBS 0.260775f
C557 B.n86 VSUBS 0.009029f
C558 B.n87 VSUBS 0.009029f
C559 B.n88 VSUBS 0.009029f
C560 B.n89 VSUBS 0.009029f
C561 B.t7 VSUBS 0.195368f
C562 B.t8 VSUBS 0.204603f
C563 B.t6 VSUBS 0.152047f
C564 B.n90 VSUBS 0.292141f
C565 B.n91 VSUBS 0.260779f
C566 B.n92 VSUBS 0.02092f
C567 B.n93 VSUBS 0.009029f
C568 B.n94 VSUBS 0.009029f
C569 B.n95 VSUBS 0.009029f
C570 B.n96 VSUBS 0.009029f
C571 B.n97 VSUBS 0.009029f
C572 B.n98 VSUBS 0.009029f
C573 B.n99 VSUBS 0.009029f
C574 B.n100 VSUBS 0.009029f
C575 B.n101 VSUBS 0.009029f
C576 B.n102 VSUBS 0.009029f
C577 B.n103 VSUBS 0.009029f
C578 B.n104 VSUBS 0.009029f
C579 B.n105 VSUBS 0.009029f
C580 B.n106 VSUBS 0.009029f
C581 B.n107 VSUBS 0.009029f
C582 B.n108 VSUBS 0.009029f
C583 B.n109 VSUBS 0.02022f
C584 B.n110 VSUBS 0.009029f
C585 B.n111 VSUBS 0.009029f
C586 B.n112 VSUBS 0.009029f
C587 B.n113 VSUBS 0.009029f
C588 B.n114 VSUBS 0.009029f
C589 B.n115 VSUBS 0.009029f
C590 B.n116 VSUBS 0.009029f
C591 B.n117 VSUBS 0.009029f
C592 B.n118 VSUBS 0.009029f
C593 B.n119 VSUBS 0.009029f
C594 B.n120 VSUBS 0.009029f
C595 B.n121 VSUBS 0.009029f
C596 B.n122 VSUBS 0.009029f
C597 B.n123 VSUBS 0.009029f
C598 B.n124 VSUBS 0.009029f
C599 B.n125 VSUBS 0.009029f
C600 B.n126 VSUBS 0.009029f
C601 B.n127 VSUBS 0.009029f
C602 B.n128 VSUBS 0.009029f
C603 B.n129 VSUBS 0.009029f
C604 B.n130 VSUBS 0.009029f
C605 B.n131 VSUBS 0.009029f
C606 B.n132 VSUBS 0.009029f
C607 B.n133 VSUBS 0.009029f
C608 B.n134 VSUBS 0.019085f
C609 B.n135 VSUBS 0.019085f
C610 B.n136 VSUBS 0.02022f
C611 B.n137 VSUBS 0.009029f
C612 B.n138 VSUBS 0.009029f
C613 B.n139 VSUBS 0.009029f
C614 B.n140 VSUBS 0.009029f
C615 B.n141 VSUBS 0.009029f
C616 B.n142 VSUBS 0.009029f
C617 B.n143 VSUBS 0.009029f
C618 B.n144 VSUBS 0.009029f
C619 B.n145 VSUBS 0.009029f
C620 B.n146 VSUBS 0.009029f
C621 B.n147 VSUBS 0.009029f
C622 B.n148 VSUBS 0.009029f
C623 B.n149 VSUBS 0.009029f
C624 B.n150 VSUBS 0.009029f
C625 B.n151 VSUBS 0.009029f
C626 B.n152 VSUBS 0.009029f
C627 B.n153 VSUBS 0.009029f
C628 B.n154 VSUBS 0.009029f
C629 B.n155 VSUBS 0.009029f
C630 B.n156 VSUBS 0.009029f
C631 B.n157 VSUBS 0.009029f
C632 B.n158 VSUBS 0.009029f
C633 B.n159 VSUBS 0.009029f
C634 B.n160 VSUBS 0.009029f
C635 B.n161 VSUBS 0.009029f
C636 B.n162 VSUBS 0.009029f
C637 B.n163 VSUBS 0.009029f
C638 B.n164 VSUBS 0.009029f
C639 B.n165 VSUBS 0.009029f
C640 B.n166 VSUBS 0.009029f
C641 B.n167 VSUBS 0.009029f
C642 B.n168 VSUBS 0.009029f
C643 B.n169 VSUBS 0.009029f
C644 B.n170 VSUBS 0.009029f
C645 B.n171 VSUBS 0.009029f
C646 B.n172 VSUBS 0.009029f
C647 B.n173 VSUBS 0.009029f
C648 B.n174 VSUBS 0.009029f
C649 B.n175 VSUBS 0.009029f
C650 B.n176 VSUBS 0.009029f
C651 B.n177 VSUBS 0.009029f
C652 B.n178 VSUBS 0.009029f
C653 B.n179 VSUBS 0.009029f
C654 B.n180 VSUBS 0.009029f
C655 B.n181 VSUBS 0.009029f
C656 B.n182 VSUBS 0.009029f
C657 B.n183 VSUBS 0.009029f
C658 B.n184 VSUBS 0.009029f
C659 B.n185 VSUBS 0.005975f
C660 B.n186 VSUBS 0.009029f
C661 B.n187 VSUBS 0.009029f
C662 B.n188 VSUBS 0.007569f
C663 B.n189 VSUBS 0.009029f
C664 B.n190 VSUBS 0.009029f
C665 B.n191 VSUBS 0.009029f
C666 B.n192 VSUBS 0.009029f
C667 B.n193 VSUBS 0.009029f
C668 B.n194 VSUBS 0.009029f
C669 B.n195 VSUBS 0.009029f
C670 B.n196 VSUBS 0.009029f
C671 B.n197 VSUBS 0.009029f
C672 B.n198 VSUBS 0.009029f
C673 B.n199 VSUBS 0.009029f
C674 B.n200 VSUBS 0.007569f
C675 B.n201 VSUBS 0.02092f
C676 B.n202 VSUBS 0.005975f
C677 B.n203 VSUBS 0.009029f
C678 B.n204 VSUBS 0.009029f
C679 B.n205 VSUBS 0.009029f
C680 B.n206 VSUBS 0.009029f
C681 B.n207 VSUBS 0.009029f
C682 B.n208 VSUBS 0.009029f
C683 B.n209 VSUBS 0.009029f
C684 B.n210 VSUBS 0.009029f
C685 B.n211 VSUBS 0.009029f
C686 B.n212 VSUBS 0.009029f
C687 B.n213 VSUBS 0.009029f
C688 B.n214 VSUBS 0.009029f
C689 B.n215 VSUBS 0.009029f
C690 B.n216 VSUBS 0.009029f
C691 B.n217 VSUBS 0.009029f
C692 B.n218 VSUBS 0.009029f
C693 B.n219 VSUBS 0.009029f
C694 B.n220 VSUBS 0.009029f
C695 B.n221 VSUBS 0.009029f
C696 B.n222 VSUBS 0.009029f
C697 B.n223 VSUBS 0.009029f
C698 B.n224 VSUBS 0.009029f
C699 B.n225 VSUBS 0.009029f
C700 B.n226 VSUBS 0.009029f
C701 B.n227 VSUBS 0.009029f
C702 B.n228 VSUBS 0.009029f
C703 B.n229 VSUBS 0.009029f
C704 B.n230 VSUBS 0.009029f
C705 B.n231 VSUBS 0.009029f
C706 B.n232 VSUBS 0.009029f
C707 B.n233 VSUBS 0.009029f
C708 B.n234 VSUBS 0.009029f
C709 B.n235 VSUBS 0.009029f
C710 B.n236 VSUBS 0.009029f
C711 B.n237 VSUBS 0.009029f
C712 B.n238 VSUBS 0.009029f
C713 B.n239 VSUBS 0.009029f
C714 B.n240 VSUBS 0.009029f
C715 B.n241 VSUBS 0.009029f
C716 B.n242 VSUBS 0.009029f
C717 B.n243 VSUBS 0.009029f
C718 B.n244 VSUBS 0.009029f
C719 B.n245 VSUBS 0.009029f
C720 B.n246 VSUBS 0.009029f
C721 B.n247 VSUBS 0.009029f
C722 B.n248 VSUBS 0.009029f
C723 B.n249 VSUBS 0.009029f
C724 B.n250 VSUBS 0.009029f
C725 B.n251 VSUBS 0.02022f
C726 B.n252 VSUBS 0.02022f
C727 B.n253 VSUBS 0.019085f
C728 B.n254 VSUBS 0.009029f
C729 B.n255 VSUBS 0.009029f
C730 B.n256 VSUBS 0.009029f
C731 B.n257 VSUBS 0.009029f
C732 B.n258 VSUBS 0.009029f
C733 B.n259 VSUBS 0.009029f
C734 B.n260 VSUBS 0.009029f
C735 B.n261 VSUBS 0.009029f
C736 B.n262 VSUBS 0.009029f
C737 B.n263 VSUBS 0.009029f
C738 B.n264 VSUBS 0.009029f
C739 B.n265 VSUBS 0.009029f
C740 B.n266 VSUBS 0.009029f
C741 B.n267 VSUBS 0.009029f
C742 B.n268 VSUBS 0.009029f
C743 B.n269 VSUBS 0.009029f
C744 B.n270 VSUBS 0.009029f
C745 B.n271 VSUBS 0.009029f
C746 B.n272 VSUBS 0.009029f
C747 B.n273 VSUBS 0.009029f
C748 B.n274 VSUBS 0.009029f
C749 B.n275 VSUBS 0.009029f
C750 B.n276 VSUBS 0.009029f
C751 B.n277 VSUBS 0.009029f
C752 B.n278 VSUBS 0.009029f
C753 B.n279 VSUBS 0.009029f
C754 B.n280 VSUBS 0.009029f
C755 B.n281 VSUBS 0.009029f
C756 B.n282 VSUBS 0.009029f
C757 B.n283 VSUBS 0.009029f
C758 B.n284 VSUBS 0.009029f
C759 B.n285 VSUBS 0.009029f
C760 B.n286 VSUBS 0.009029f
C761 B.n287 VSUBS 0.009029f
C762 B.n288 VSUBS 0.009029f
C763 B.n289 VSUBS 0.009029f
C764 B.n290 VSUBS 0.009029f
C765 B.n291 VSUBS 0.009029f
C766 B.n292 VSUBS 0.009029f
C767 B.n293 VSUBS 0.009029f
C768 B.n294 VSUBS 0.009029f
C769 B.n295 VSUBS 0.019085f
C770 B.n296 VSUBS 0.02022f
C771 B.n297 VSUBS 0.019026f
C772 B.n298 VSUBS 0.009029f
C773 B.n299 VSUBS 0.009029f
C774 B.n300 VSUBS 0.009029f
C775 B.n301 VSUBS 0.009029f
C776 B.n302 VSUBS 0.009029f
C777 B.n303 VSUBS 0.009029f
C778 B.n304 VSUBS 0.009029f
C779 B.n305 VSUBS 0.009029f
C780 B.n306 VSUBS 0.009029f
C781 B.n307 VSUBS 0.009029f
C782 B.n308 VSUBS 0.009029f
C783 B.n309 VSUBS 0.009029f
C784 B.n310 VSUBS 0.009029f
C785 B.n311 VSUBS 0.009029f
C786 B.n312 VSUBS 0.009029f
C787 B.n313 VSUBS 0.009029f
C788 B.n314 VSUBS 0.009029f
C789 B.n315 VSUBS 0.009029f
C790 B.n316 VSUBS 0.009029f
C791 B.n317 VSUBS 0.009029f
C792 B.n318 VSUBS 0.009029f
C793 B.n319 VSUBS 0.009029f
C794 B.n320 VSUBS 0.009029f
C795 B.n321 VSUBS 0.009029f
C796 B.n322 VSUBS 0.009029f
C797 B.n323 VSUBS 0.009029f
C798 B.n324 VSUBS 0.009029f
C799 B.n325 VSUBS 0.009029f
C800 B.n326 VSUBS 0.009029f
C801 B.n327 VSUBS 0.009029f
C802 B.n328 VSUBS 0.009029f
C803 B.n329 VSUBS 0.009029f
C804 B.n330 VSUBS 0.009029f
C805 B.n331 VSUBS 0.009029f
C806 B.n332 VSUBS 0.009029f
C807 B.n333 VSUBS 0.009029f
C808 B.n334 VSUBS 0.009029f
C809 B.n335 VSUBS 0.009029f
C810 B.n336 VSUBS 0.009029f
C811 B.n337 VSUBS 0.009029f
C812 B.n338 VSUBS 0.009029f
C813 B.n339 VSUBS 0.009029f
C814 B.n340 VSUBS 0.009029f
C815 B.n341 VSUBS 0.009029f
C816 B.n342 VSUBS 0.009029f
C817 B.n343 VSUBS 0.009029f
C818 B.n344 VSUBS 0.009029f
C819 B.n345 VSUBS 0.009029f
C820 B.n346 VSUBS 0.005975f
C821 B.n347 VSUBS 0.02092f
C822 B.n348 VSUBS 0.007569f
C823 B.n349 VSUBS 0.009029f
C824 B.n350 VSUBS 0.009029f
C825 B.n351 VSUBS 0.009029f
C826 B.n352 VSUBS 0.009029f
C827 B.n353 VSUBS 0.009029f
C828 B.n354 VSUBS 0.009029f
C829 B.n355 VSUBS 0.009029f
C830 B.n356 VSUBS 0.009029f
C831 B.n357 VSUBS 0.009029f
C832 B.n358 VSUBS 0.009029f
C833 B.n359 VSUBS 0.009029f
C834 B.n360 VSUBS 0.007569f
C835 B.n361 VSUBS 0.009029f
C836 B.n362 VSUBS 0.009029f
C837 B.n363 VSUBS 0.005975f
C838 B.n364 VSUBS 0.009029f
C839 B.n365 VSUBS 0.009029f
C840 B.n366 VSUBS 0.009029f
C841 B.n367 VSUBS 0.009029f
C842 B.n368 VSUBS 0.009029f
C843 B.n369 VSUBS 0.009029f
C844 B.n370 VSUBS 0.009029f
C845 B.n371 VSUBS 0.009029f
C846 B.n372 VSUBS 0.009029f
C847 B.n373 VSUBS 0.009029f
C848 B.n374 VSUBS 0.009029f
C849 B.n375 VSUBS 0.009029f
C850 B.n376 VSUBS 0.009029f
C851 B.n377 VSUBS 0.009029f
C852 B.n378 VSUBS 0.009029f
C853 B.n379 VSUBS 0.009029f
C854 B.n380 VSUBS 0.009029f
C855 B.n381 VSUBS 0.009029f
C856 B.n382 VSUBS 0.009029f
C857 B.n383 VSUBS 0.009029f
C858 B.n384 VSUBS 0.009029f
C859 B.n385 VSUBS 0.009029f
C860 B.n386 VSUBS 0.009029f
C861 B.n387 VSUBS 0.009029f
C862 B.n388 VSUBS 0.009029f
C863 B.n389 VSUBS 0.009029f
C864 B.n390 VSUBS 0.009029f
C865 B.n391 VSUBS 0.009029f
C866 B.n392 VSUBS 0.009029f
C867 B.n393 VSUBS 0.009029f
C868 B.n394 VSUBS 0.009029f
C869 B.n395 VSUBS 0.009029f
C870 B.n396 VSUBS 0.009029f
C871 B.n397 VSUBS 0.009029f
C872 B.n398 VSUBS 0.009029f
C873 B.n399 VSUBS 0.009029f
C874 B.n400 VSUBS 0.009029f
C875 B.n401 VSUBS 0.009029f
C876 B.n402 VSUBS 0.009029f
C877 B.n403 VSUBS 0.009029f
C878 B.n404 VSUBS 0.009029f
C879 B.n405 VSUBS 0.009029f
C880 B.n406 VSUBS 0.009029f
C881 B.n407 VSUBS 0.009029f
C882 B.n408 VSUBS 0.009029f
C883 B.n409 VSUBS 0.009029f
C884 B.n410 VSUBS 0.009029f
C885 B.n411 VSUBS 0.009029f
C886 B.n412 VSUBS 0.02022f
C887 B.n413 VSUBS 0.019085f
C888 B.n414 VSUBS 0.019085f
C889 B.n415 VSUBS 0.009029f
C890 B.n416 VSUBS 0.009029f
C891 B.n417 VSUBS 0.009029f
C892 B.n418 VSUBS 0.009029f
C893 B.n419 VSUBS 0.009029f
C894 B.n420 VSUBS 0.009029f
C895 B.n421 VSUBS 0.009029f
C896 B.n422 VSUBS 0.009029f
C897 B.n423 VSUBS 0.009029f
C898 B.n424 VSUBS 0.009029f
C899 B.n425 VSUBS 0.009029f
C900 B.n426 VSUBS 0.009029f
C901 B.n427 VSUBS 0.009029f
C902 B.n428 VSUBS 0.009029f
C903 B.n429 VSUBS 0.009029f
C904 B.n430 VSUBS 0.009029f
C905 B.n431 VSUBS 0.009029f
C906 B.n432 VSUBS 0.009029f
C907 B.n433 VSUBS 0.009029f
C908 B.n434 VSUBS 0.009029f
C909 B.n435 VSUBS 0.020446f
.ends

