* NGSPICE file created from diff_pair_sample_0567.ext - technology: sky130A

.subckt diff_pair_sample_0567 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t5 VN.t0 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=1.94535 ps=12.12 w=11.79 l=3.11
X1 VTAIL.t7 VN.t1 VDD2.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=1.94535 ps=12.12 w=11.79 l=3.11
X2 VTAIL.t3 VP.t0 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=1.94535 ps=12.12 w=11.79 l=3.11
X3 VDD2.t3 VN.t2 VTAIL.t10 B.t4 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=1.94535 ps=12.12 w=11.79 l=3.11
X4 VTAIL.t8 VN.t3 VDD2.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=1.94535 ps=12.12 w=11.79 l=3.11
X5 VDD1.t4 VP.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=4.5981 ps=24.36 w=11.79 l=3.11
X6 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=0 ps=0 w=11.79 l=3.11
X7 VDD1.t3 VP.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=1.94535 ps=12.12 w=11.79 l=3.11
X8 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=0 ps=0 w=11.79 l=3.11
X9 VDD2.t1 VN.t4 VTAIL.t11 B.t5 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=4.5981 ps=24.36 w=11.79 l=3.11
X10 VTAIL.t1 VP.t3 VDD1.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=1.94535 ps=12.12 w=11.79 l=3.11
X11 VDD2.t0 VN.t5 VTAIL.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=4.5981 ps=24.36 w=11.79 l=3.11
X12 VDD1.t1 VP.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.94535 pd=12.12 as=4.5981 ps=24.36 w=11.79 l=3.11
X13 VDD1.t0 VP.t5 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=1.94535 ps=12.12 w=11.79 l=3.11
X14 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=0 ps=0 w=11.79 l=3.11
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=4.5981 pd=24.36 as=0 ps=0 w=11.79 l=3.11
R0 VN.n30 VN.n29 161.3
R1 VN.n28 VN.n17 161.3
R2 VN.n27 VN.n26 161.3
R3 VN.n25 VN.n18 161.3
R4 VN.n24 VN.n23 161.3
R5 VN.n22 VN.n19 161.3
R6 VN.n14 VN.n13 161.3
R7 VN.n12 VN.n1 161.3
R8 VN.n11 VN.n10 161.3
R9 VN.n9 VN.n2 161.3
R10 VN.n8 VN.n7 161.3
R11 VN.n6 VN.n3 161.3
R12 VN.n20 VN.t5 124.781
R13 VN.n4 VN.t0 124.781
R14 VN.n5 VN.t1 91.3635
R15 VN.n0 VN.t4 91.3635
R16 VN.n21 VN.t3 91.3635
R17 VN.n16 VN.t2 91.3635
R18 VN.n15 VN.n0 68.5364
R19 VN.n31 VN.n16 68.5364
R20 VN.n11 VN.n2 56.5193
R21 VN.n27 VN.n18 56.5193
R22 VN VN.n31 50.8541
R23 VN.n5 VN.n4 49.4728
R24 VN.n21 VN.n20 49.4728
R25 VN.n6 VN.n5 24.4675
R26 VN.n7 VN.n6 24.4675
R27 VN.n7 VN.n2 24.4675
R28 VN.n12 VN.n11 24.4675
R29 VN.n13 VN.n12 24.4675
R30 VN.n23 VN.n18 24.4675
R31 VN.n23 VN.n22 24.4675
R32 VN.n22 VN.n21 24.4675
R33 VN.n29 VN.n28 24.4675
R34 VN.n28 VN.n27 24.4675
R35 VN.n13 VN.n0 21.5315
R36 VN.n29 VN.n16 21.5315
R37 VN.n20 VN.n19 3.84099
R38 VN.n4 VN.n3 3.84099
R39 VN.n31 VN.n30 0.354971
R40 VN.n15 VN.n14 0.354971
R41 VN VN.n15 0.26696
R42 VN.n30 VN.n17 0.189894
R43 VN.n26 VN.n17 0.189894
R44 VN.n26 VN.n25 0.189894
R45 VN.n25 VN.n24 0.189894
R46 VN.n24 VN.n19 0.189894
R47 VN.n8 VN.n3 0.189894
R48 VN.n9 VN.n8 0.189894
R49 VN.n10 VN.n9 0.189894
R50 VN.n10 VN.n1 0.189894
R51 VN.n14 VN.n1 0.189894
R52 VTAIL.n7 VTAIL.t6 47.5624
R53 VTAIL.n11 VTAIL.t11 47.5622
R54 VTAIL.n2 VTAIL.t0 47.5622
R55 VTAIL.n10 VTAIL.t5 47.5622
R56 VTAIL.n9 VTAIL.n8 45.8831
R57 VTAIL.n6 VTAIL.n5 45.8831
R58 VTAIL.n1 VTAIL.n0 45.8828
R59 VTAIL.n4 VTAIL.n3 45.8828
R60 VTAIL.n6 VTAIL.n4 28.4617
R61 VTAIL.n11 VTAIL.n10 25.4962
R62 VTAIL.n7 VTAIL.n6 2.96602
R63 VTAIL.n10 VTAIL.n9 2.96602
R64 VTAIL.n4 VTAIL.n2 2.96602
R65 VTAIL VTAIL.n11 2.16645
R66 VTAIL.n9 VTAIL.n7 1.95309
R67 VTAIL.n2 VTAIL.n1 1.95309
R68 VTAIL.n0 VTAIL.t9 1.67989
R69 VTAIL.n0 VTAIL.t7 1.67989
R70 VTAIL.n3 VTAIL.t4 1.67989
R71 VTAIL.n3 VTAIL.t1 1.67989
R72 VTAIL.n8 VTAIL.t2 1.67989
R73 VTAIL.n8 VTAIL.t3 1.67989
R74 VTAIL.n5 VTAIL.t10 1.67989
R75 VTAIL.n5 VTAIL.t8 1.67989
R76 VTAIL VTAIL.n1 0.800069
R77 VDD2.n1 VDD2.t5 66.4098
R78 VDD2.n2 VDD2.t3 64.2412
R79 VDD2.n1 VDD2.n0 63.2476
R80 VDD2 VDD2.n3 63.2449
R81 VDD2.n2 VDD2.n1 43.517
R82 VDD2 VDD2.n2 2.28283
R83 VDD2.n3 VDD2.t2 1.67989
R84 VDD2.n3 VDD2.t0 1.67989
R85 VDD2.n0 VDD2.t4 1.67989
R86 VDD2.n0 VDD2.t1 1.67989
R87 B.n859 B.n858 585
R88 B.n321 B.n136 585
R89 B.n320 B.n319 585
R90 B.n318 B.n317 585
R91 B.n316 B.n315 585
R92 B.n314 B.n313 585
R93 B.n312 B.n311 585
R94 B.n310 B.n309 585
R95 B.n308 B.n307 585
R96 B.n306 B.n305 585
R97 B.n304 B.n303 585
R98 B.n302 B.n301 585
R99 B.n300 B.n299 585
R100 B.n298 B.n297 585
R101 B.n296 B.n295 585
R102 B.n294 B.n293 585
R103 B.n292 B.n291 585
R104 B.n290 B.n289 585
R105 B.n288 B.n287 585
R106 B.n286 B.n285 585
R107 B.n284 B.n283 585
R108 B.n282 B.n281 585
R109 B.n280 B.n279 585
R110 B.n278 B.n277 585
R111 B.n276 B.n275 585
R112 B.n274 B.n273 585
R113 B.n272 B.n271 585
R114 B.n270 B.n269 585
R115 B.n268 B.n267 585
R116 B.n266 B.n265 585
R117 B.n264 B.n263 585
R118 B.n262 B.n261 585
R119 B.n260 B.n259 585
R120 B.n258 B.n257 585
R121 B.n256 B.n255 585
R122 B.n254 B.n253 585
R123 B.n252 B.n251 585
R124 B.n250 B.n249 585
R125 B.n248 B.n247 585
R126 B.n246 B.n245 585
R127 B.n244 B.n243 585
R128 B.n241 B.n240 585
R129 B.n239 B.n238 585
R130 B.n237 B.n236 585
R131 B.n235 B.n234 585
R132 B.n233 B.n232 585
R133 B.n231 B.n230 585
R134 B.n229 B.n228 585
R135 B.n227 B.n226 585
R136 B.n225 B.n224 585
R137 B.n223 B.n222 585
R138 B.n220 B.n219 585
R139 B.n218 B.n217 585
R140 B.n216 B.n215 585
R141 B.n214 B.n213 585
R142 B.n212 B.n211 585
R143 B.n210 B.n209 585
R144 B.n208 B.n207 585
R145 B.n206 B.n205 585
R146 B.n204 B.n203 585
R147 B.n202 B.n201 585
R148 B.n200 B.n199 585
R149 B.n198 B.n197 585
R150 B.n196 B.n195 585
R151 B.n194 B.n193 585
R152 B.n192 B.n191 585
R153 B.n190 B.n189 585
R154 B.n188 B.n187 585
R155 B.n186 B.n185 585
R156 B.n184 B.n183 585
R157 B.n182 B.n181 585
R158 B.n180 B.n179 585
R159 B.n178 B.n177 585
R160 B.n176 B.n175 585
R161 B.n174 B.n173 585
R162 B.n172 B.n171 585
R163 B.n170 B.n169 585
R164 B.n168 B.n167 585
R165 B.n166 B.n165 585
R166 B.n164 B.n163 585
R167 B.n162 B.n161 585
R168 B.n160 B.n159 585
R169 B.n158 B.n157 585
R170 B.n156 B.n155 585
R171 B.n154 B.n153 585
R172 B.n152 B.n151 585
R173 B.n150 B.n149 585
R174 B.n148 B.n147 585
R175 B.n146 B.n145 585
R176 B.n144 B.n143 585
R177 B.n142 B.n141 585
R178 B.n89 B.n88 585
R179 B.n857 B.n90 585
R180 B.n862 B.n90 585
R181 B.n856 B.n855 585
R182 B.n855 B.n86 585
R183 B.n854 B.n85 585
R184 B.n868 B.n85 585
R185 B.n853 B.n84 585
R186 B.n869 B.n84 585
R187 B.n852 B.n83 585
R188 B.n870 B.n83 585
R189 B.n851 B.n850 585
R190 B.n850 B.n79 585
R191 B.n849 B.n78 585
R192 B.n876 B.n78 585
R193 B.n848 B.n77 585
R194 B.n877 B.n77 585
R195 B.n847 B.n76 585
R196 B.n878 B.n76 585
R197 B.n846 B.n845 585
R198 B.n845 B.n72 585
R199 B.n844 B.n71 585
R200 B.n884 B.n71 585
R201 B.n843 B.n70 585
R202 B.n885 B.n70 585
R203 B.n842 B.n69 585
R204 B.n886 B.n69 585
R205 B.n841 B.n840 585
R206 B.n840 B.n65 585
R207 B.n839 B.n64 585
R208 B.n892 B.n64 585
R209 B.n838 B.n63 585
R210 B.n893 B.n63 585
R211 B.n837 B.n62 585
R212 B.n894 B.n62 585
R213 B.n836 B.n835 585
R214 B.n835 B.n58 585
R215 B.n834 B.n57 585
R216 B.n900 B.n57 585
R217 B.n833 B.n56 585
R218 B.n901 B.n56 585
R219 B.n832 B.n55 585
R220 B.n902 B.n55 585
R221 B.n831 B.n830 585
R222 B.n830 B.n54 585
R223 B.n829 B.n50 585
R224 B.n908 B.n50 585
R225 B.n828 B.n49 585
R226 B.n909 B.n49 585
R227 B.n827 B.n48 585
R228 B.n910 B.n48 585
R229 B.n826 B.n825 585
R230 B.n825 B.n44 585
R231 B.n824 B.n43 585
R232 B.n916 B.n43 585
R233 B.n823 B.n42 585
R234 B.n917 B.n42 585
R235 B.n822 B.n41 585
R236 B.n918 B.n41 585
R237 B.n821 B.n820 585
R238 B.n820 B.n37 585
R239 B.n819 B.n36 585
R240 B.n924 B.n36 585
R241 B.n818 B.n35 585
R242 B.n925 B.n35 585
R243 B.n817 B.n34 585
R244 B.n926 B.n34 585
R245 B.n816 B.n815 585
R246 B.n815 B.n30 585
R247 B.n814 B.n29 585
R248 B.n932 B.n29 585
R249 B.n813 B.n28 585
R250 B.n933 B.n28 585
R251 B.n812 B.n27 585
R252 B.n934 B.n27 585
R253 B.n811 B.n810 585
R254 B.n810 B.n23 585
R255 B.n809 B.n22 585
R256 B.n940 B.n22 585
R257 B.n808 B.n21 585
R258 B.n941 B.n21 585
R259 B.n807 B.n20 585
R260 B.n942 B.n20 585
R261 B.n806 B.n805 585
R262 B.n805 B.n19 585
R263 B.n804 B.n15 585
R264 B.n948 B.n15 585
R265 B.n803 B.n14 585
R266 B.n949 B.n14 585
R267 B.n802 B.n13 585
R268 B.n950 B.n13 585
R269 B.n801 B.n800 585
R270 B.n800 B.n12 585
R271 B.n799 B.n798 585
R272 B.n799 B.n8 585
R273 B.n797 B.n7 585
R274 B.n957 B.n7 585
R275 B.n796 B.n6 585
R276 B.n958 B.n6 585
R277 B.n795 B.n5 585
R278 B.n959 B.n5 585
R279 B.n794 B.n793 585
R280 B.n793 B.n4 585
R281 B.n792 B.n322 585
R282 B.n792 B.n791 585
R283 B.n782 B.n323 585
R284 B.n324 B.n323 585
R285 B.n784 B.n783 585
R286 B.n785 B.n784 585
R287 B.n781 B.n329 585
R288 B.n329 B.n328 585
R289 B.n780 B.n779 585
R290 B.n779 B.n778 585
R291 B.n331 B.n330 585
R292 B.n771 B.n331 585
R293 B.n770 B.n769 585
R294 B.n772 B.n770 585
R295 B.n768 B.n336 585
R296 B.n336 B.n335 585
R297 B.n767 B.n766 585
R298 B.n766 B.n765 585
R299 B.n338 B.n337 585
R300 B.n339 B.n338 585
R301 B.n758 B.n757 585
R302 B.n759 B.n758 585
R303 B.n756 B.n344 585
R304 B.n344 B.n343 585
R305 B.n755 B.n754 585
R306 B.n754 B.n753 585
R307 B.n346 B.n345 585
R308 B.n347 B.n346 585
R309 B.n746 B.n745 585
R310 B.n747 B.n746 585
R311 B.n744 B.n351 585
R312 B.n355 B.n351 585
R313 B.n743 B.n742 585
R314 B.n742 B.n741 585
R315 B.n353 B.n352 585
R316 B.n354 B.n353 585
R317 B.n734 B.n733 585
R318 B.n735 B.n734 585
R319 B.n732 B.n360 585
R320 B.n360 B.n359 585
R321 B.n731 B.n730 585
R322 B.n730 B.n729 585
R323 B.n362 B.n361 585
R324 B.n363 B.n362 585
R325 B.n722 B.n721 585
R326 B.n723 B.n722 585
R327 B.n720 B.n368 585
R328 B.n368 B.n367 585
R329 B.n719 B.n718 585
R330 B.n718 B.n717 585
R331 B.n370 B.n369 585
R332 B.n710 B.n370 585
R333 B.n709 B.n708 585
R334 B.n711 B.n709 585
R335 B.n707 B.n375 585
R336 B.n375 B.n374 585
R337 B.n706 B.n705 585
R338 B.n705 B.n704 585
R339 B.n377 B.n376 585
R340 B.n378 B.n377 585
R341 B.n697 B.n696 585
R342 B.n698 B.n697 585
R343 B.n695 B.n383 585
R344 B.n383 B.n382 585
R345 B.n694 B.n693 585
R346 B.n693 B.n692 585
R347 B.n385 B.n384 585
R348 B.n386 B.n385 585
R349 B.n685 B.n684 585
R350 B.n686 B.n685 585
R351 B.n683 B.n391 585
R352 B.n391 B.n390 585
R353 B.n682 B.n681 585
R354 B.n681 B.n680 585
R355 B.n393 B.n392 585
R356 B.n394 B.n393 585
R357 B.n673 B.n672 585
R358 B.n674 B.n673 585
R359 B.n671 B.n399 585
R360 B.n399 B.n398 585
R361 B.n670 B.n669 585
R362 B.n669 B.n668 585
R363 B.n401 B.n400 585
R364 B.n402 B.n401 585
R365 B.n661 B.n660 585
R366 B.n662 B.n661 585
R367 B.n659 B.n407 585
R368 B.n407 B.n406 585
R369 B.n658 B.n657 585
R370 B.n657 B.n656 585
R371 B.n409 B.n408 585
R372 B.n410 B.n409 585
R373 B.n649 B.n648 585
R374 B.n650 B.n649 585
R375 B.n413 B.n412 585
R376 B.n468 B.n467 585
R377 B.n469 B.n465 585
R378 B.n465 B.n414 585
R379 B.n471 B.n470 585
R380 B.n473 B.n464 585
R381 B.n476 B.n475 585
R382 B.n477 B.n463 585
R383 B.n479 B.n478 585
R384 B.n481 B.n462 585
R385 B.n484 B.n483 585
R386 B.n485 B.n461 585
R387 B.n487 B.n486 585
R388 B.n489 B.n460 585
R389 B.n492 B.n491 585
R390 B.n493 B.n459 585
R391 B.n495 B.n494 585
R392 B.n497 B.n458 585
R393 B.n500 B.n499 585
R394 B.n501 B.n457 585
R395 B.n503 B.n502 585
R396 B.n505 B.n456 585
R397 B.n508 B.n507 585
R398 B.n509 B.n455 585
R399 B.n511 B.n510 585
R400 B.n513 B.n454 585
R401 B.n516 B.n515 585
R402 B.n517 B.n453 585
R403 B.n519 B.n518 585
R404 B.n521 B.n452 585
R405 B.n524 B.n523 585
R406 B.n525 B.n451 585
R407 B.n527 B.n526 585
R408 B.n529 B.n450 585
R409 B.n532 B.n531 585
R410 B.n533 B.n449 585
R411 B.n535 B.n534 585
R412 B.n537 B.n448 585
R413 B.n540 B.n539 585
R414 B.n541 B.n447 585
R415 B.n543 B.n542 585
R416 B.n545 B.n446 585
R417 B.n548 B.n547 585
R418 B.n549 B.n442 585
R419 B.n551 B.n550 585
R420 B.n553 B.n441 585
R421 B.n556 B.n555 585
R422 B.n557 B.n440 585
R423 B.n559 B.n558 585
R424 B.n561 B.n439 585
R425 B.n564 B.n563 585
R426 B.n565 B.n436 585
R427 B.n568 B.n567 585
R428 B.n570 B.n435 585
R429 B.n573 B.n572 585
R430 B.n574 B.n434 585
R431 B.n576 B.n575 585
R432 B.n578 B.n433 585
R433 B.n581 B.n580 585
R434 B.n582 B.n432 585
R435 B.n584 B.n583 585
R436 B.n586 B.n431 585
R437 B.n589 B.n588 585
R438 B.n590 B.n430 585
R439 B.n592 B.n591 585
R440 B.n594 B.n429 585
R441 B.n597 B.n596 585
R442 B.n598 B.n428 585
R443 B.n600 B.n599 585
R444 B.n602 B.n427 585
R445 B.n605 B.n604 585
R446 B.n606 B.n426 585
R447 B.n608 B.n607 585
R448 B.n610 B.n425 585
R449 B.n613 B.n612 585
R450 B.n614 B.n424 585
R451 B.n616 B.n615 585
R452 B.n618 B.n423 585
R453 B.n621 B.n620 585
R454 B.n622 B.n422 585
R455 B.n624 B.n623 585
R456 B.n626 B.n421 585
R457 B.n629 B.n628 585
R458 B.n630 B.n420 585
R459 B.n632 B.n631 585
R460 B.n634 B.n419 585
R461 B.n637 B.n636 585
R462 B.n638 B.n418 585
R463 B.n640 B.n639 585
R464 B.n642 B.n417 585
R465 B.n643 B.n416 585
R466 B.n646 B.n645 585
R467 B.n647 B.n415 585
R468 B.n415 B.n414 585
R469 B.n652 B.n651 585
R470 B.n651 B.n650 585
R471 B.n653 B.n411 585
R472 B.n411 B.n410 585
R473 B.n655 B.n654 585
R474 B.n656 B.n655 585
R475 B.n405 B.n404 585
R476 B.n406 B.n405 585
R477 B.n664 B.n663 585
R478 B.n663 B.n662 585
R479 B.n665 B.n403 585
R480 B.n403 B.n402 585
R481 B.n667 B.n666 585
R482 B.n668 B.n667 585
R483 B.n397 B.n396 585
R484 B.n398 B.n397 585
R485 B.n676 B.n675 585
R486 B.n675 B.n674 585
R487 B.n677 B.n395 585
R488 B.n395 B.n394 585
R489 B.n679 B.n678 585
R490 B.n680 B.n679 585
R491 B.n389 B.n388 585
R492 B.n390 B.n389 585
R493 B.n688 B.n687 585
R494 B.n687 B.n686 585
R495 B.n689 B.n387 585
R496 B.n387 B.n386 585
R497 B.n691 B.n690 585
R498 B.n692 B.n691 585
R499 B.n381 B.n380 585
R500 B.n382 B.n381 585
R501 B.n700 B.n699 585
R502 B.n699 B.n698 585
R503 B.n701 B.n379 585
R504 B.n379 B.n378 585
R505 B.n703 B.n702 585
R506 B.n704 B.n703 585
R507 B.n373 B.n372 585
R508 B.n374 B.n373 585
R509 B.n713 B.n712 585
R510 B.n712 B.n711 585
R511 B.n714 B.n371 585
R512 B.n710 B.n371 585
R513 B.n716 B.n715 585
R514 B.n717 B.n716 585
R515 B.n366 B.n365 585
R516 B.n367 B.n366 585
R517 B.n725 B.n724 585
R518 B.n724 B.n723 585
R519 B.n726 B.n364 585
R520 B.n364 B.n363 585
R521 B.n728 B.n727 585
R522 B.n729 B.n728 585
R523 B.n358 B.n357 585
R524 B.n359 B.n358 585
R525 B.n737 B.n736 585
R526 B.n736 B.n735 585
R527 B.n738 B.n356 585
R528 B.n356 B.n354 585
R529 B.n740 B.n739 585
R530 B.n741 B.n740 585
R531 B.n350 B.n349 585
R532 B.n355 B.n350 585
R533 B.n749 B.n748 585
R534 B.n748 B.n747 585
R535 B.n750 B.n348 585
R536 B.n348 B.n347 585
R537 B.n752 B.n751 585
R538 B.n753 B.n752 585
R539 B.n342 B.n341 585
R540 B.n343 B.n342 585
R541 B.n761 B.n760 585
R542 B.n760 B.n759 585
R543 B.n762 B.n340 585
R544 B.n340 B.n339 585
R545 B.n764 B.n763 585
R546 B.n765 B.n764 585
R547 B.n334 B.n333 585
R548 B.n335 B.n334 585
R549 B.n774 B.n773 585
R550 B.n773 B.n772 585
R551 B.n775 B.n332 585
R552 B.n771 B.n332 585
R553 B.n777 B.n776 585
R554 B.n778 B.n777 585
R555 B.n327 B.n326 585
R556 B.n328 B.n327 585
R557 B.n787 B.n786 585
R558 B.n786 B.n785 585
R559 B.n788 B.n325 585
R560 B.n325 B.n324 585
R561 B.n790 B.n789 585
R562 B.n791 B.n790 585
R563 B.n3 B.n0 585
R564 B.n4 B.n3 585
R565 B.n956 B.n1 585
R566 B.n957 B.n956 585
R567 B.n955 B.n954 585
R568 B.n955 B.n8 585
R569 B.n953 B.n9 585
R570 B.n12 B.n9 585
R571 B.n952 B.n951 585
R572 B.n951 B.n950 585
R573 B.n11 B.n10 585
R574 B.n949 B.n11 585
R575 B.n947 B.n946 585
R576 B.n948 B.n947 585
R577 B.n945 B.n16 585
R578 B.n19 B.n16 585
R579 B.n944 B.n943 585
R580 B.n943 B.n942 585
R581 B.n18 B.n17 585
R582 B.n941 B.n18 585
R583 B.n939 B.n938 585
R584 B.n940 B.n939 585
R585 B.n937 B.n24 585
R586 B.n24 B.n23 585
R587 B.n936 B.n935 585
R588 B.n935 B.n934 585
R589 B.n26 B.n25 585
R590 B.n933 B.n26 585
R591 B.n931 B.n930 585
R592 B.n932 B.n931 585
R593 B.n929 B.n31 585
R594 B.n31 B.n30 585
R595 B.n928 B.n927 585
R596 B.n927 B.n926 585
R597 B.n33 B.n32 585
R598 B.n925 B.n33 585
R599 B.n923 B.n922 585
R600 B.n924 B.n923 585
R601 B.n921 B.n38 585
R602 B.n38 B.n37 585
R603 B.n920 B.n919 585
R604 B.n919 B.n918 585
R605 B.n40 B.n39 585
R606 B.n917 B.n40 585
R607 B.n915 B.n914 585
R608 B.n916 B.n915 585
R609 B.n913 B.n45 585
R610 B.n45 B.n44 585
R611 B.n912 B.n911 585
R612 B.n911 B.n910 585
R613 B.n47 B.n46 585
R614 B.n909 B.n47 585
R615 B.n907 B.n906 585
R616 B.n908 B.n907 585
R617 B.n905 B.n51 585
R618 B.n54 B.n51 585
R619 B.n904 B.n903 585
R620 B.n903 B.n902 585
R621 B.n53 B.n52 585
R622 B.n901 B.n53 585
R623 B.n899 B.n898 585
R624 B.n900 B.n899 585
R625 B.n897 B.n59 585
R626 B.n59 B.n58 585
R627 B.n896 B.n895 585
R628 B.n895 B.n894 585
R629 B.n61 B.n60 585
R630 B.n893 B.n61 585
R631 B.n891 B.n890 585
R632 B.n892 B.n891 585
R633 B.n889 B.n66 585
R634 B.n66 B.n65 585
R635 B.n888 B.n887 585
R636 B.n887 B.n886 585
R637 B.n68 B.n67 585
R638 B.n885 B.n68 585
R639 B.n883 B.n882 585
R640 B.n884 B.n883 585
R641 B.n881 B.n73 585
R642 B.n73 B.n72 585
R643 B.n880 B.n879 585
R644 B.n879 B.n878 585
R645 B.n75 B.n74 585
R646 B.n877 B.n75 585
R647 B.n875 B.n874 585
R648 B.n876 B.n875 585
R649 B.n873 B.n80 585
R650 B.n80 B.n79 585
R651 B.n872 B.n871 585
R652 B.n871 B.n870 585
R653 B.n82 B.n81 585
R654 B.n869 B.n82 585
R655 B.n867 B.n866 585
R656 B.n868 B.n867 585
R657 B.n865 B.n87 585
R658 B.n87 B.n86 585
R659 B.n864 B.n863 585
R660 B.n863 B.n862 585
R661 B.n960 B.n959 585
R662 B.n958 B.n2 585
R663 B.n863 B.n89 478.086
R664 B.n859 B.n90 478.086
R665 B.n649 B.n415 478.086
R666 B.n651 B.n413 478.086
R667 B.n139 B.t6 300.068
R668 B.n137 B.t14 300.068
R669 B.n437 B.t10 300.068
R670 B.n443 B.t17 300.068
R671 B.n861 B.n860 256.663
R672 B.n861 B.n135 256.663
R673 B.n861 B.n134 256.663
R674 B.n861 B.n133 256.663
R675 B.n861 B.n132 256.663
R676 B.n861 B.n131 256.663
R677 B.n861 B.n130 256.663
R678 B.n861 B.n129 256.663
R679 B.n861 B.n128 256.663
R680 B.n861 B.n127 256.663
R681 B.n861 B.n126 256.663
R682 B.n861 B.n125 256.663
R683 B.n861 B.n124 256.663
R684 B.n861 B.n123 256.663
R685 B.n861 B.n122 256.663
R686 B.n861 B.n121 256.663
R687 B.n861 B.n120 256.663
R688 B.n861 B.n119 256.663
R689 B.n861 B.n118 256.663
R690 B.n861 B.n117 256.663
R691 B.n861 B.n116 256.663
R692 B.n861 B.n115 256.663
R693 B.n861 B.n114 256.663
R694 B.n861 B.n113 256.663
R695 B.n861 B.n112 256.663
R696 B.n861 B.n111 256.663
R697 B.n861 B.n110 256.663
R698 B.n861 B.n109 256.663
R699 B.n861 B.n108 256.663
R700 B.n861 B.n107 256.663
R701 B.n861 B.n106 256.663
R702 B.n861 B.n105 256.663
R703 B.n861 B.n104 256.663
R704 B.n861 B.n103 256.663
R705 B.n861 B.n102 256.663
R706 B.n861 B.n101 256.663
R707 B.n861 B.n100 256.663
R708 B.n861 B.n99 256.663
R709 B.n861 B.n98 256.663
R710 B.n861 B.n97 256.663
R711 B.n861 B.n96 256.663
R712 B.n861 B.n95 256.663
R713 B.n861 B.n94 256.663
R714 B.n861 B.n93 256.663
R715 B.n861 B.n92 256.663
R716 B.n861 B.n91 256.663
R717 B.n466 B.n414 256.663
R718 B.n472 B.n414 256.663
R719 B.n474 B.n414 256.663
R720 B.n480 B.n414 256.663
R721 B.n482 B.n414 256.663
R722 B.n488 B.n414 256.663
R723 B.n490 B.n414 256.663
R724 B.n496 B.n414 256.663
R725 B.n498 B.n414 256.663
R726 B.n504 B.n414 256.663
R727 B.n506 B.n414 256.663
R728 B.n512 B.n414 256.663
R729 B.n514 B.n414 256.663
R730 B.n520 B.n414 256.663
R731 B.n522 B.n414 256.663
R732 B.n528 B.n414 256.663
R733 B.n530 B.n414 256.663
R734 B.n536 B.n414 256.663
R735 B.n538 B.n414 256.663
R736 B.n544 B.n414 256.663
R737 B.n546 B.n414 256.663
R738 B.n552 B.n414 256.663
R739 B.n554 B.n414 256.663
R740 B.n560 B.n414 256.663
R741 B.n562 B.n414 256.663
R742 B.n569 B.n414 256.663
R743 B.n571 B.n414 256.663
R744 B.n577 B.n414 256.663
R745 B.n579 B.n414 256.663
R746 B.n585 B.n414 256.663
R747 B.n587 B.n414 256.663
R748 B.n593 B.n414 256.663
R749 B.n595 B.n414 256.663
R750 B.n601 B.n414 256.663
R751 B.n603 B.n414 256.663
R752 B.n609 B.n414 256.663
R753 B.n611 B.n414 256.663
R754 B.n617 B.n414 256.663
R755 B.n619 B.n414 256.663
R756 B.n625 B.n414 256.663
R757 B.n627 B.n414 256.663
R758 B.n633 B.n414 256.663
R759 B.n635 B.n414 256.663
R760 B.n641 B.n414 256.663
R761 B.n644 B.n414 256.663
R762 B.n962 B.n961 256.663
R763 B.n143 B.n142 163.367
R764 B.n147 B.n146 163.367
R765 B.n151 B.n150 163.367
R766 B.n155 B.n154 163.367
R767 B.n159 B.n158 163.367
R768 B.n163 B.n162 163.367
R769 B.n167 B.n166 163.367
R770 B.n171 B.n170 163.367
R771 B.n175 B.n174 163.367
R772 B.n179 B.n178 163.367
R773 B.n183 B.n182 163.367
R774 B.n187 B.n186 163.367
R775 B.n191 B.n190 163.367
R776 B.n195 B.n194 163.367
R777 B.n199 B.n198 163.367
R778 B.n203 B.n202 163.367
R779 B.n207 B.n206 163.367
R780 B.n211 B.n210 163.367
R781 B.n215 B.n214 163.367
R782 B.n219 B.n218 163.367
R783 B.n224 B.n223 163.367
R784 B.n228 B.n227 163.367
R785 B.n232 B.n231 163.367
R786 B.n236 B.n235 163.367
R787 B.n240 B.n239 163.367
R788 B.n245 B.n244 163.367
R789 B.n249 B.n248 163.367
R790 B.n253 B.n252 163.367
R791 B.n257 B.n256 163.367
R792 B.n261 B.n260 163.367
R793 B.n265 B.n264 163.367
R794 B.n269 B.n268 163.367
R795 B.n273 B.n272 163.367
R796 B.n277 B.n276 163.367
R797 B.n281 B.n280 163.367
R798 B.n285 B.n284 163.367
R799 B.n289 B.n288 163.367
R800 B.n293 B.n292 163.367
R801 B.n297 B.n296 163.367
R802 B.n301 B.n300 163.367
R803 B.n305 B.n304 163.367
R804 B.n309 B.n308 163.367
R805 B.n313 B.n312 163.367
R806 B.n317 B.n316 163.367
R807 B.n319 B.n136 163.367
R808 B.n649 B.n409 163.367
R809 B.n657 B.n409 163.367
R810 B.n657 B.n407 163.367
R811 B.n661 B.n407 163.367
R812 B.n661 B.n401 163.367
R813 B.n669 B.n401 163.367
R814 B.n669 B.n399 163.367
R815 B.n673 B.n399 163.367
R816 B.n673 B.n393 163.367
R817 B.n681 B.n393 163.367
R818 B.n681 B.n391 163.367
R819 B.n685 B.n391 163.367
R820 B.n685 B.n385 163.367
R821 B.n693 B.n385 163.367
R822 B.n693 B.n383 163.367
R823 B.n697 B.n383 163.367
R824 B.n697 B.n377 163.367
R825 B.n705 B.n377 163.367
R826 B.n705 B.n375 163.367
R827 B.n709 B.n375 163.367
R828 B.n709 B.n370 163.367
R829 B.n718 B.n370 163.367
R830 B.n718 B.n368 163.367
R831 B.n722 B.n368 163.367
R832 B.n722 B.n362 163.367
R833 B.n730 B.n362 163.367
R834 B.n730 B.n360 163.367
R835 B.n734 B.n360 163.367
R836 B.n734 B.n353 163.367
R837 B.n742 B.n353 163.367
R838 B.n742 B.n351 163.367
R839 B.n746 B.n351 163.367
R840 B.n746 B.n346 163.367
R841 B.n754 B.n346 163.367
R842 B.n754 B.n344 163.367
R843 B.n758 B.n344 163.367
R844 B.n758 B.n338 163.367
R845 B.n766 B.n338 163.367
R846 B.n766 B.n336 163.367
R847 B.n770 B.n336 163.367
R848 B.n770 B.n331 163.367
R849 B.n779 B.n331 163.367
R850 B.n779 B.n329 163.367
R851 B.n784 B.n329 163.367
R852 B.n784 B.n323 163.367
R853 B.n792 B.n323 163.367
R854 B.n793 B.n792 163.367
R855 B.n793 B.n5 163.367
R856 B.n6 B.n5 163.367
R857 B.n7 B.n6 163.367
R858 B.n799 B.n7 163.367
R859 B.n800 B.n799 163.367
R860 B.n800 B.n13 163.367
R861 B.n14 B.n13 163.367
R862 B.n15 B.n14 163.367
R863 B.n805 B.n15 163.367
R864 B.n805 B.n20 163.367
R865 B.n21 B.n20 163.367
R866 B.n22 B.n21 163.367
R867 B.n810 B.n22 163.367
R868 B.n810 B.n27 163.367
R869 B.n28 B.n27 163.367
R870 B.n29 B.n28 163.367
R871 B.n815 B.n29 163.367
R872 B.n815 B.n34 163.367
R873 B.n35 B.n34 163.367
R874 B.n36 B.n35 163.367
R875 B.n820 B.n36 163.367
R876 B.n820 B.n41 163.367
R877 B.n42 B.n41 163.367
R878 B.n43 B.n42 163.367
R879 B.n825 B.n43 163.367
R880 B.n825 B.n48 163.367
R881 B.n49 B.n48 163.367
R882 B.n50 B.n49 163.367
R883 B.n830 B.n50 163.367
R884 B.n830 B.n55 163.367
R885 B.n56 B.n55 163.367
R886 B.n57 B.n56 163.367
R887 B.n835 B.n57 163.367
R888 B.n835 B.n62 163.367
R889 B.n63 B.n62 163.367
R890 B.n64 B.n63 163.367
R891 B.n840 B.n64 163.367
R892 B.n840 B.n69 163.367
R893 B.n70 B.n69 163.367
R894 B.n71 B.n70 163.367
R895 B.n845 B.n71 163.367
R896 B.n845 B.n76 163.367
R897 B.n77 B.n76 163.367
R898 B.n78 B.n77 163.367
R899 B.n850 B.n78 163.367
R900 B.n850 B.n83 163.367
R901 B.n84 B.n83 163.367
R902 B.n85 B.n84 163.367
R903 B.n855 B.n85 163.367
R904 B.n855 B.n90 163.367
R905 B.n467 B.n465 163.367
R906 B.n471 B.n465 163.367
R907 B.n475 B.n473 163.367
R908 B.n479 B.n463 163.367
R909 B.n483 B.n481 163.367
R910 B.n487 B.n461 163.367
R911 B.n491 B.n489 163.367
R912 B.n495 B.n459 163.367
R913 B.n499 B.n497 163.367
R914 B.n503 B.n457 163.367
R915 B.n507 B.n505 163.367
R916 B.n511 B.n455 163.367
R917 B.n515 B.n513 163.367
R918 B.n519 B.n453 163.367
R919 B.n523 B.n521 163.367
R920 B.n527 B.n451 163.367
R921 B.n531 B.n529 163.367
R922 B.n535 B.n449 163.367
R923 B.n539 B.n537 163.367
R924 B.n543 B.n447 163.367
R925 B.n547 B.n545 163.367
R926 B.n551 B.n442 163.367
R927 B.n555 B.n553 163.367
R928 B.n559 B.n440 163.367
R929 B.n563 B.n561 163.367
R930 B.n568 B.n436 163.367
R931 B.n572 B.n570 163.367
R932 B.n576 B.n434 163.367
R933 B.n580 B.n578 163.367
R934 B.n584 B.n432 163.367
R935 B.n588 B.n586 163.367
R936 B.n592 B.n430 163.367
R937 B.n596 B.n594 163.367
R938 B.n600 B.n428 163.367
R939 B.n604 B.n602 163.367
R940 B.n608 B.n426 163.367
R941 B.n612 B.n610 163.367
R942 B.n616 B.n424 163.367
R943 B.n620 B.n618 163.367
R944 B.n624 B.n422 163.367
R945 B.n628 B.n626 163.367
R946 B.n632 B.n420 163.367
R947 B.n636 B.n634 163.367
R948 B.n640 B.n418 163.367
R949 B.n643 B.n642 163.367
R950 B.n645 B.n415 163.367
R951 B.n651 B.n411 163.367
R952 B.n655 B.n411 163.367
R953 B.n655 B.n405 163.367
R954 B.n663 B.n405 163.367
R955 B.n663 B.n403 163.367
R956 B.n667 B.n403 163.367
R957 B.n667 B.n397 163.367
R958 B.n675 B.n397 163.367
R959 B.n675 B.n395 163.367
R960 B.n679 B.n395 163.367
R961 B.n679 B.n389 163.367
R962 B.n687 B.n389 163.367
R963 B.n687 B.n387 163.367
R964 B.n691 B.n387 163.367
R965 B.n691 B.n381 163.367
R966 B.n699 B.n381 163.367
R967 B.n699 B.n379 163.367
R968 B.n703 B.n379 163.367
R969 B.n703 B.n373 163.367
R970 B.n712 B.n373 163.367
R971 B.n712 B.n371 163.367
R972 B.n716 B.n371 163.367
R973 B.n716 B.n366 163.367
R974 B.n724 B.n366 163.367
R975 B.n724 B.n364 163.367
R976 B.n728 B.n364 163.367
R977 B.n728 B.n358 163.367
R978 B.n736 B.n358 163.367
R979 B.n736 B.n356 163.367
R980 B.n740 B.n356 163.367
R981 B.n740 B.n350 163.367
R982 B.n748 B.n350 163.367
R983 B.n748 B.n348 163.367
R984 B.n752 B.n348 163.367
R985 B.n752 B.n342 163.367
R986 B.n760 B.n342 163.367
R987 B.n760 B.n340 163.367
R988 B.n764 B.n340 163.367
R989 B.n764 B.n334 163.367
R990 B.n773 B.n334 163.367
R991 B.n773 B.n332 163.367
R992 B.n777 B.n332 163.367
R993 B.n777 B.n327 163.367
R994 B.n786 B.n327 163.367
R995 B.n786 B.n325 163.367
R996 B.n790 B.n325 163.367
R997 B.n790 B.n3 163.367
R998 B.n960 B.n3 163.367
R999 B.n956 B.n2 163.367
R1000 B.n956 B.n955 163.367
R1001 B.n955 B.n9 163.367
R1002 B.n951 B.n9 163.367
R1003 B.n951 B.n11 163.367
R1004 B.n947 B.n11 163.367
R1005 B.n947 B.n16 163.367
R1006 B.n943 B.n16 163.367
R1007 B.n943 B.n18 163.367
R1008 B.n939 B.n18 163.367
R1009 B.n939 B.n24 163.367
R1010 B.n935 B.n24 163.367
R1011 B.n935 B.n26 163.367
R1012 B.n931 B.n26 163.367
R1013 B.n931 B.n31 163.367
R1014 B.n927 B.n31 163.367
R1015 B.n927 B.n33 163.367
R1016 B.n923 B.n33 163.367
R1017 B.n923 B.n38 163.367
R1018 B.n919 B.n38 163.367
R1019 B.n919 B.n40 163.367
R1020 B.n915 B.n40 163.367
R1021 B.n915 B.n45 163.367
R1022 B.n911 B.n45 163.367
R1023 B.n911 B.n47 163.367
R1024 B.n907 B.n47 163.367
R1025 B.n907 B.n51 163.367
R1026 B.n903 B.n51 163.367
R1027 B.n903 B.n53 163.367
R1028 B.n899 B.n53 163.367
R1029 B.n899 B.n59 163.367
R1030 B.n895 B.n59 163.367
R1031 B.n895 B.n61 163.367
R1032 B.n891 B.n61 163.367
R1033 B.n891 B.n66 163.367
R1034 B.n887 B.n66 163.367
R1035 B.n887 B.n68 163.367
R1036 B.n883 B.n68 163.367
R1037 B.n883 B.n73 163.367
R1038 B.n879 B.n73 163.367
R1039 B.n879 B.n75 163.367
R1040 B.n875 B.n75 163.367
R1041 B.n875 B.n80 163.367
R1042 B.n871 B.n80 163.367
R1043 B.n871 B.n82 163.367
R1044 B.n867 B.n82 163.367
R1045 B.n867 B.n87 163.367
R1046 B.n863 B.n87 163.367
R1047 B.n137 B.t15 138.994
R1048 B.n437 B.t13 138.994
R1049 B.n139 B.t8 138.98
R1050 B.n443 B.t19 138.98
R1051 B.n650 B.n414 83.1531
R1052 B.n862 B.n861 83.1531
R1053 B.n138 B.t16 72.2794
R1054 B.n438 B.t12 72.2794
R1055 B.n140 B.t9 72.2647
R1056 B.n444 B.t18 72.2647
R1057 B.n91 B.n89 71.676
R1058 B.n143 B.n92 71.676
R1059 B.n147 B.n93 71.676
R1060 B.n151 B.n94 71.676
R1061 B.n155 B.n95 71.676
R1062 B.n159 B.n96 71.676
R1063 B.n163 B.n97 71.676
R1064 B.n167 B.n98 71.676
R1065 B.n171 B.n99 71.676
R1066 B.n175 B.n100 71.676
R1067 B.n179 B.n101 71.676
R1068 B.n183 B.n102 71.676
R1069 B.n187 B.n103 71.676
R1070 B.n191 B.n104 71.676
R1071 B.n195 B.n105 71.676
R1072 B.n199 B.n106 71.676
R1073 B.n203 B.n107 71.676
R1074 B.n207 B.n108 71.676
R1075 B.n211 B.n109 71.676
R1076 B.n215 B.n110 71.676
R1077 B.n219 B.n111 71.676
R1078 B.n224 B.n112 71.676
R1079 B.n228 B.n113 71.676
R1080 B.n232 B.n114 71.676
R1081 B.n236 B.n115 71.676
R1082 B.n240 B.n116 71.676
R1083 B.n245 B.n117 71.676
R1084 B.n249 B.n118 71.676
R1085 B.n253 B.n119 71.676
R1086 B.n257 B.n120 71.676
R1087 B.n261 B.n121 71.676
R1088 B.n265 B.n122 71.676
R1089 B.n269 B.n123 71.676
R1090 B.n273 B.n124 71.676
R1091 B.n277 B.n125 71.676
R1092 B.n281 B.n126 71.676
R1093 B.n285 B.n127 71.676
R1094 B.n289 B.n128 71.676
R1095 B.n293 B.n129 71.676
R1096 B.n297 B.n130 71.676
R1097 B.n301 B.n131 71.676
R1098 B.n305 B.n132 71.676
R1099 B.n309 B.n133 71.676
R1100 B.n313 B.n134 71.676
R1101 B.n317 B.n135 71.676
R1102 B.n860 B.n136 71.676
R1103 B.n860 B.n859 71.676
R1104 B.n319 B.n135 71.676
R1105 B.n316 B.n134 71.676
R1106 B.n312 B.n133 71.676
R1107 B.n308 B.n132 71.676
R1108 B.n304 B.n131 71.676
R1109 B.n300 B.n130 71.676
R1110 B.n296 B.n129 71.676
R1111 B.n292 B.n128 71.676
R1112 B.n288 B.n127 71.676
R1113 B.n284 B.n126 71.676
R1114 B.n280 B.n125 71.676
R1115 B.n276 B.n124 71.676
R1116 B.n272 B.n123 71.676
R1117 B.n268 B.n122 71.676
R1118 B.n264 B.n121 71.676
R1119 B.n260 B.n120 71.676
R1120 B.n256 B.n119 71.676
R1121 B.n252 B.n118 71.676
R1122 B.n248 B.n117 71.676
R1123 B.n244 B.n116 71.676
R1124 B.n239 B.n115 71.676
R1125 B.n235 B.n114 71.676
R1126 B.n231 B.n113 71.676
R1127 B.n227 B.n112 71.676
R1128 B.n223 B.n111 71.676
R1129 B.n218 B.n110 71.676
R1130 B.n214 B.n109 71.676
R1131 B.n210 B.n108 71.676
R1132 B.n206 B.n107 71.676
R1133 B.n202 B.n106 71.676
R1134 B.n198 B.n105 71.676
R1135 B.n194 B.n104 71.676
R1136 B.n190 B.n103 71.676
R1137 B.n186 B.n102 71.676
R1138 B.n182 B.n101 71.676
R1139 B.n178 B.n100 71.676
R1140 B.n174 B.n99 71.676
R1141 B.n170 B.n98 71.676
R1142 B.n166 B.n97 71.676
R1143 B.n162 B.n96 71.676
R1144 B.n158 B.n95 71.676
R1145 B.n154 B.n94 71.676
R1146 B.n150 B.n93 71.676
R1147 B.n146 B.n92 71.676
R1148 B.n142 B.n91 71.676
R1149 B.n466 B.n413 71.676
R1150 B.n472 B.n471 71.676
R1151 B.n475 B.n474 71.676
R1152 B.n480 B.n479 71.676
R1153 B.n483 B.n482 71.676
R1154 B.n488 B.n487 71.676
R1155 B.n491 B.n490 71.676
R1156 B.n496 B.n495 71.676
R1157 B.n499 B.n498 71.676
R1158 B.n504 B.n503 71.676
R1159 B.n507 B.n506 71.676
R1160 B.n512 B.n511 71.676
R1161 B.n515 B.n514 71.676
R1162 B.n520 B.n519 71.676
R1163 B.n523 B.n522 71.676
R1164 B.n528 B.n527 71.676
R1165 B.n531 B.n530 71.676
R1166 B.n536 B.n535 71.676
R1167 B.n539 B.n538 71.676
R1168 B.n544 B.n543 71.676
R1169 B.n547 B.n546 71.676
R1170 B.n552 B.n551 71.676
R1171 B.n555 B.n554 71.676
R1172 B.n560 B.n559 71.676
R1173 B.n563 B.n562 71.676
R1174 B.n569 B.n568 71.676
R1175 B.n572 B.n571 71.676
R1176 B.n577 B.n576 71.676
R1177 B.n580 B.n579 71.676
R1178 B.n585 B.n584 71.676
R1179 B.n588 B.n587 71.676
R1180 B.n593 B.n592 71.676
R1181 B.n596 B.n595 71.676
R1182 B.n601 B.n600 71.676
R1183 B.n604 B.n603 71.676
R1184 B.n609 B.n608 71.676
R1185 B.n612 B.n611 71.676
R1186 B.n617 B.n616 71.676
R1187 B.n620 B.n619 71.676
R1188 B.n625 B.n624 71.676
R1189 B.n628 B.n627 71.676
R1190 B.n633 B.n632 71.676
R1191 B.n636 B.n635 71.676
R1192 B.n641 B.n640 71.676
R1193 B.n644 B.n643 71.676
R1194 B.n467 B.n466 71.676
R1195 B.n473 B.n472 71.676
R1196 B.n474 B.n463 71.676
R1197 B.n481 B.n480 71.676
R1198 B.n482 B.n461 71.676
R1199 B.n489 B.n488 71.676
R1200 B.n490 B.n459 71.676
R1201 B.n497 B.n496 71.676
R1202 B.n498 B.n457 71.676
R1203 B.n505 B.n504 71.676
R1204 B.n506 B.n455 71.676
R1205 B.n513 B.n512 71.676
R1206 B.n514 B.n453 71.676
R1207 B.n521 B.n520 71.676
R1208 B.n522 B.n451 71.676
R1209 B.n529 B.n528 71.676
R1210 B.n530 B.n449 71.676
R1211 B.n537 B.n536 71.676
R1212 B.n538 B.n447 71.676
R1213 B.n545 B.n544 71.676
R1214 B.n546 B.n442 71.676
R1215 B.n553 B.n552 71.676
R1216 B.n554 B.n440 71.676
R1217 B.n561 B.n560 71.676
R1218 B.n562 B.n436 71.676
R1219 B.n570 B.n569 71.676
R1220 B.n571 B.n434 71.676
R1221 B.n578 B.n577 71.676
R1222 B.n579 B.n432 71.676
R1223 B.n586 B.n585 71.676
R1224 B.n587 B.n430 71.676
R1225 B.n594 B.n593 71.676
R1226 B.n595 B.n428 71.676
R1227 B.n602 B.n601 71.676
R1228 B.n603 B.n426 71.676
R1229 B.n610 B.n609 71.676
R1230 B.n611 B.n424 71.676
R1231 B.n618 B.n617 71.676
R1232 B.n619 B.n422 71.676
R1233 B.n626 B.n625 71.676
R1234 B.n627 B.n420 71.676
R1235 B.n634 B.n633 71.676
R1236 B.n635 B.n418 71.676
R1237 B.n642 B.n641 71.676
R1238 B.n645 B.n644 71.676
R1239 B.n961 B.n960 71.676
R1240 B.n961 B.n2 71.676
R1241 B.n140 B.n139 66.7156
R1242 B.n138 B.n137 66.7156
R1243 B.n438 B.n437 66.7156
R1244 B.n444 B.n443 66.7156
R1245 B.n221 B.n140 59.5399
R1246 B.n242 B.n138 59.5399
R1247 B.n566 B.n438 59.5399
R1248 B.n445 B.n444 59.5399
R1249 B.n650 B.n410 43.8329
R1250 B.n656 B.n410 43.8329
R1251 B.n656 B.n406 43.8329
R1252 B.n662 B.n406 43.8329
R1253 B.n662 B.n402 43.8329
R1254 B.n668 B.n402 43.8329
R1255 B.n668 B.n398 43.8329
R1256 B.n674 B.n398 43.8329
R1257 B.n680 B.n394 43.8329
R1258 B.n680 B.n390 43.8329
R1259 B.n686 B.n390 43.8329
R1260 B.n686 B.n386 43.8329
R1261 B.n692 B.n386 43.8329
R1262 B.n692 B.n382 43.8329
R1263 B.n698 B.n382 43.8329
R1264 B.n698 B.n378 43.8329
R1265 B.n704 B.n378 43.8329
R1266 B.n704 B.n374 43.8329
R1267 B.n711 B.n374 43.8329
R1268 B.n711 B.n710 43.8329
R1269 B.n717 B.n367 43.8329
R1270 B.n723 B.n367 43.8329
R1271 B.n723 B.n363 43.8329
R1272 B.n729 B.n363 43.8329
R1273 B.n729 B.n359 43.8329
R1274 B.n735 B.n359 43.8329
R1275 B.n735 B.n354 43.8329
R1276 B.n741 B.n354 43.8329
R1277 B.n741 B.n355 43.8329
R1278 B.n747 B.n347 43.8329
R1279 B.n753 B.n347 43.8329
R1280 B.n753 B.n343 43.8329
R1281 B.n759 B.n343 43.8329
R1282 B.n759 B.n339 43.8329
R1283 B.n765 B.n339 43.8329
R1284 B.n765 B.n335 43.8329
R1285 B.n772 B.n335 43.8329
R1286 B.n772 B.n771 43.8329
R1287 B.n778 B.n328 43.8329
R1288 B.n785 B.n328 43.8329
R1289 B.n785 B.n324 43.8329
R1290 B.n791 B.n324 43.8329
R1291 B.n791 B.n4 43.8329
R1292 B.n959 B.n4 43.8329
R1293 B.n959 B.n958 43.8329
R1294 B.n958 B.n957 43.8329
R1295 B.n957 B.n8 43.8329
R1296 B.n12 B.n8 43.8329
R1297 B.n950 B.n12 43.8329
R1298 B.n950 B.n949 43.8329
R1299 B.n949 B.n948 43.8329
R1300 B.n942 B.n19 43.8329
R1301 B.n942 B.n941 43.8329
R1302 B.n941 B.n940 43.8329
R1303 B.n940 B.n23 43.8329
R1304 B.n934 B.n23 43.8329
R1305 B.n934 B.n933 43.8329
R1306 B.n933 B.n932 43.8329
R1307 B.n932 B.n30 43.8329
R1308 B.n926 B.n30 43.8329
R1309 B.n925 B.n924 43.8329
R1310 B.n924 B.n37 43.8329
R1311 B.n918 B.n37 43.8329
R1312 B.n918 B.n917 43.8329
R1313 B.n917 B.n916 43.8329
R1314 B.n916 B.n44 43.8329
R1315 B.n910 B.n44 43.8329
R1316 B.n910 B.n909 43.8329
R1317 B.n909 B.n908 43.8329
R1318 B.n902 B.n54 43.8329
R1319 B.n902 B.n901 43.8329
R1320 B.n901 B.n900 43.8329
R1321 B.n900 B.n58 43.8329
R1322 B.n894 B.n58 43.8329
R1323 B.n894 B.n893 43.8329
R1324 B.n893 B.n892 43.8329
R1325 B.n892 B.n65 43.8329
R1326 B.n886 B.n65 43.8329
R1327 B.n886 B.n885 43.8329
R1328 B.n885 B.n884 43.8329
R1329 B.n884 B.n72 43.8329
R1330 B.n878 B.n877 43.8329
R1331 B.n877 B.n876 43.8329
R1332 B.n876 B.n79 43.8329
R1333 B.n870 B.n79 43.8329
R1334 B.n870 B.n869 43.8329
R1335 B.n869 B.n868 43.8329
R1336 B.n868 B.n86 43.8329
R1337 B.n862 B.n86 43.8329
R1338 B.n771 B.t0 36.7424
R1339 B.n19 B.t2 36.7424
R1340 B.t11 B.n394 31.5856
R1341 B.n355 B.t1 31.5856
R1342 B.t3 B.n925 31.5856
R1343 B.t7 B.n72 31.5856
R1344 B.n652 B.n412 31.0639
R1345 B.n648 B.n647 31.0639
R1346 B.n858 B.n857 31.0639
R1347 B.n864 B.n88 31.0639
R1348 B.n710 B.t4 26.4289
R1349 B.n54 B.t5 26.4289
R1350 B B.n962 18.0485
R1351 B.n717 B.t4 17.4045
R1352 B.n908 B.t5 17.4045
R1353 B.n674 B.t11 12.2478
R1354 B.n747 B.t1 12.2478
R1355 B.n926 B.t3 12.2478
R1356 B.n878 B.t7 12.2478
R1357 B.n653 B.n652 10.6151
R1358 B.n654 B.n653 10.6151
R1359 B.n654 B.n404 10.6151
R1360 B.n664 B.n404 10.6151
R1361 B.n665 B.n664 10.6151
R1362 B.n666 B.n665 10.6151
R1363 B.n666 B.n396 10.6151
R1364 B.n676 B.n396 10.6151
R1365 B.n677 B.n676 10.6151
R1366 B.n678 B.n677 10.6151
R1367 B.n678 B.n388 10.6151
R1368 B.n688 B.n388 10.6151
R1369 B.n689 B.n688 10.6151
R1370 B.n690 B.n689 10.6151
R1371 B.n690 B.n380 10.6151
R1372 B.n700 B.n380 10.6151
R1373 B.n701 B.n700 10.6151
R1374 B.n702 B.n701 10.6151
R1375 B.n702 B.n372 10.6151
R1376 B.n713 B.n372 10.6151
R1377 B.n714 B.n713 10.6151
R1378 B.n715 B.n714 10.6151
R1379 B.n715 B.n365 10.6151
R1380 B.n725 B.n365 10.6151
R1381 B.n726 B.n725 10.6151
R1382 B.n727 B.n726 10.6151
R1383 B.n727 B.n357 10.6151
R1384 B.n737 B.n357 10.6151
R1385 B.n738 B.n737 10.6151
R1386 B.n739 B.n738 10.6151
R1387 B.n739 B.n349 10.6151
R1388 B.n749 B.n349 10.6151
R1389 B.n750 B.n749 10.6151
R1390 B.n751 B.n750 10.6151
R1391 B.n751 B.n341 10.6151
R1392 B.n761 B.n341 10.6151
R1393 B.n762 B.n761 10.6151
R1394 B.n763 B.n762 10.6151
R1395 B.n763 B.n333 10.6151
R1396 B.n774 B.n333 10.6151
R1397 B.n775 B.n774 10.6151
R1398 B.n776 B.n775 10.6151
R1399 B.n776 B.n326 10.6151
R1400 B.n787 B.n326 10.6151
R1401 B.n788 B.n787 10.6151
R1402 B.n789 B.n788 10.6151
R1403 B.n789 B.n0 10.6151
R1404 B.n468 B.n412 10.6151
R1405 B.n469 B.n468 10.6151
R1406 B.n470 B.n469 10.6151
R1407 B.n470 B.n464 10.6151
R1408 B.n476 B.n464 10.6151
R1409 B.n477 B.n476 10.6151
R1410 B.n478 B.n477 10.6151
R1411 B.n478 B.n462 10.6151
R1412 B.n484 B.n462 10.6151
R1413 B.n485 B.n484 10.6151
R1414 B.n486 B.n485 10.6151
R1415 B.n486 B.n460 10.6151
R1416 B.n492 B.n460 10.6151
R1417 B.n493 B.n492 10.6151
R1418 B.n494 B.n493 10.6151
R1419 B.n494 B.n458 10.6151
R1420 B.n500 B.n458 10.6151
R1421 B.n501 B.n500 10.6151
R1422 B.n502 B.n501 10.6151
R1423 B.n502 B.n456 10.6151
R1424 B.n508 B.n456 10.6151
R1425 B.n509 B.n508 10.6151
R1426 B.n510 B.n509 10.6151
R1427 B.n510 B.n454 10.6151
R1428 B.n516 B.n454 10.6151
R1429 B.n517 B.n516 10.6151
R1430 B.n518 B.n517 10.6151
R1431 B.n518 B.n452 10.6151
R1432 B.n524 B.n452 10.6151
R1433 B.n525 B.n524 10.6151
R1434 B.n526 B.n525 10.6151
R1435 B.n526 B.n450 10.6151
R1436 B.n532 B.n450 10.6151
R1437 B.n533 B.n532 10.6151
R1438 B.n534 B.n533 10.6151
R1439 B.n534 B.n448 10.6151
R1440 B.n540 B.n448 10.6151
R1441 B.n541 B.n540 10.6151
R1442 B.n542 B.n541 10.6151
R1443 B.n542 B.n446 10.6151
R1444 B.n549 B.n548 10.6151
R1445 B.n550 B.n549 10.6151
R1446 B.n550 B.n441 10.6151
R1447 B.n556 B.n441 10.6151
R1448 B.n557 B.n556 10.6151
R1449 B.n558 B.n557 10.6151
R1450 B.n558 B.n439 10.6151
R1451 B.n564 B.n439 10.6151
R1452 B.n565 B.n564 10.6151
R1453 B.n567 B.n435 10.6151
R1454 B.n573 B.n435 10.6151
R1455 B.n574 B.n573 10.6151
R1456 B.n575 B.n574 10.6151
R1457 B.n575 B.n433 10.6151
R1458 B.n581 B.n433 10.6151
R1459 B.n582 B.n581 10.6151
R1460 B.n583 B.n582 10.6151
R1461 B.n583 B.n431 10.6151
R1462 B.n589 B.n431 10.6151
R1463 B.n590 B.n589 10.6151
R1464 B.n591 B.n590 10.6151
R1465 B.n591 B.n429 10.6151
R1466 B.n597 B.n429 10.6151
R1467 B.n598 B.n597 10.6151
R1468 B.n599 B.n598 10.6151
R1469 B.n599 B.n427 10.6151
R1470 B.n605 B.n427 10.6151
R1471 B.n606 B.n605 10.6151
R1472 B.n607 B.n606 10.6151
R1473 B.n607 B.n425 10.6151
R1474 B.n613 B.n425 10.6151
R1475 B.n614 B.n613 10.6151
R1476 B.n615 B.n614 10.6151
R1477 B.n615 B.n423 10.6151
R1478 B.n621 B.n423 10.6151
R1479 B.n622 B.n621 10.6151
R1480 B.n623 B.n622 10.6151
R1481 B.n623 B.n421 10.6151
R1482 B.n629 B.n421 10.6151
R1483 B.n630 B.n629 10.6151
R1484 B.n631 B.n630 10.6151
R1485 B.n631 B.n419 10.6151
R1486 B.n637 B.n419 10.6151
R1487 B.n638 B.n637 10.6151
R1488 B.n639 B.n638 10.6151
R1489 B.n639 B.n417 10.6151
R1490 B.n417 B.n416 10.6151
R1491 B.n646 B.n416 10.6151
R1492 B.n647 B.n646 10.6151
R1493 B.n648 B.n408 10.6151
R1494 B.n658 B.n408 10.6151
R1495 B.n659 B.n658 10.6151
R1496 B.n660 B.n659 10.6151
R1497 B.n660 B.n400 10.6151
R1498 B.n670 B.n400 10.6151
R1499 B.n671 B.n670 10.6151
R1500 B.n672 B.n671 10.6151
R1501 B.n672 B.n392 10.6151
R1502 B.n682 B.n392 10.6151
R1503 B.n683 B.n682 10.6151
R1504 B.n684 B.n683 10.6151
R1505 B.n684 B.n384 10.6151
R1506 B.n694 B.n384 10.6151
R1507 B.n695 B.n694 10.6151
R1508 B.n696 B.n695 10.6151
R1509 B.n696 B.n376 10.6151
R1510 B.n706 B.n376 10.6151
R1511 B.n707 B.n706 10.6151
R1512 B.n708 B.n707 10.6151
R1513 B.n708 B.n369 10.6151
R1514 B.n719 B.n369 10.6151
R1515 B.n720 B.n719 10.6151
R1516 B.n721 B.n720 10.6151
R1517 B.n721 B.n361 10.6151
R1518 B.n731 B.n361 10.6151
R1519 B.n732 B.n731 10.6151
R1520 B.n733 B.n732 10.6151
R1521 B.n733 B.n352 10.6151
R1522 B.n743 B.n352 10.6151
R1523 B.n744 B.n743 10.6151
R1524 B.n745 B.n744 10.6151
R1525 B.n745 B.n345 10.6151
R1526 B.n755 B.n345 10.6151
R1527 B.n756 B.n755 10.6151
R1528 B.n757 B.n756 10.6151
R1529 B.n757 B.n337 10.6151
R1530 B.n767 B.n337 10.6151
R1531 B.n768 B.n767 10.6151
R1532 B.n769 B.n768 10.6151
R1533 B.n769 B.n330 10.6151
R1534 B.n780 B.n330 10.6151
R1535 B.n781 B.n780 10.6151
R1536 B.n783 B.n781 10.6151
R1537 B.n783 B.n782 10.6151
R1538 B.n782 B.n322 10.6151
R1539 B.n794 B.n322 10.6151
R1540 B.n795 B.n794 10.6151
R1541 B.n796 B.n795 10.6151
R1542 B.n797 B.n796 10.6151
R1543 B.n798 B.n797 10.6151
R1544 B.n801 B.n798 10.6151
R1545 B.n802 B.n801 10.6151
R1546 B.n803 B.n802 10.6151
R1547 B.n804 B.n803 10.6151
R1548 B.n806 B.n804 10.6151
R1549 B.n807 B.n806 10.6151
R1550 B.n808 B.n807 10.6151
R1551 B.n809 B.n808 10.6151
R1552 B.n811 B.n809 10.6151
R1553 B.n812 B.n811 10.6151
R1554 B.n813 B.n812 10.6151
R1555 B.n814 B.n813 10.6151
R1556 B.n816 B.n814 10.6151
R1557 B.n817 B.n816 10.6151
R1558 B.n818 B.n817 10.6151
R1559 B.n819 B.n818 10.6151
R1560 B.n821 B.n819 10.6151
R1561 B.n822 B.n821 10.6151
R1562 B.n823 B.n822 10.6151
R1563 B.n824 B.n823 10.6151
R1564 B.n826 B.n824 10.6151
R1565 B.n827 B.n826 10.6151
R1566 B.n828 B.n827 10.6151
R1567 B.n829 B.n828 10.6151
R1568 B.n831 B.n829 10.6151
R1569 B.n832 B.n831 10.6151
R1570 B.n833 B.n832 10.6151
R1571 B.n834 B.n833 10.6151
R1572 B.n836 B.n834 10.6151
R1573 B.n837 B.n836 10.6151
R1574 B.n838 B.n837 10.6151
R1575 B.n839 B.n838 10.6151
R1576 B.n841 B.n839 10.6151
R1577 B.n842 B.n841 10.6151
R1578 B.n843 B.n842 10.6151
R1579 B.n844 B.n843 10.6151
R1580 B.n846 B.n844 10.6151
R1581 B.n847 B.n846 10.6151
R1582 B.n848 B.n847 10.6151
R1583 B.n849 B.n848 10.6151
R1584 B.n851 B.n849 10.6151
R1585 B.n852 B.n851 10.6151
R1586 B.n853 B.n852 10.6151
R1587 B.n854 B.n853 10.6151
R1588 B.n856 B.n854 10.6151
R1589 B.n857 B.n856 10.6151
R1590 B.n954 B.n1 10.6151
R1591 B.n954 B.n953 10.6151
R1592 B.n953 B.n952 10.6151
R1593 B.n952 B.n10 10.6151
R1594 B.n946 B.n10 10.6151
R1595 B.n946 B.n945 10.6151
R1596 B.n945 B.n944 10.6151
R1597 B.n944 B.n17 10.6151
R1598 B.n938 B.n17 10.6151
R1599 B.n938 B.n937 10.6151
R1600 B.n937 B.n936 10.6151
R1601 B.n936 B.n25 10.6151
R1602 B.n930 B.n25 10.6151
R1603 B.n930 B.n929 10.6151
R1604 B.n929 B.n928 10.6151
R1605 B.n928 B.n32 10.6151
R1606 B.n922 B.n32 10.6151
R1607 B.n922 B.n921 10.6151
R1608 B.n921 B.n920 10.6151
R1609 B.n920 B.n39 10.6151
R1610 B.n914 B.n39 10.6151
R1611 B.n914 B.n913 10.6151
R1612 B.n913 B.n912 10.6151
R1613 B.n912 B.n46 10.6151
R1614 B.n906 B.n46 10.6151
R1615 B.n906 B.n905 10.6151
R1616 B.n905 B.n904 10.6151
R1617 B.n904 B.n52 10.6151
R1618 B.n898 B.n52 10.6151
R1619 B.n898 B.n897 10.6151
R1620 B.n897 B.n896 10.6151
R1621 B.n896 B.n60 10.6151
R1622 B.n890 B.n60 10.6151
R1623 B.n890 B.n889 10.6151
R1624 B.n889 B.n888 10.6151
R1625 B.n888 B.n67 10.6151
R1626 B.n882 B.n67 10.6151
R1627 B.n882 B.n881 10.6151
R1628 B.n881 B.n880 10.6151
R1629 B.n880 B.n74 10.6151
R1630 B.n874 B.n74 10.6151
R1631 B.n874 B.n873 10.6151
R1632 B.n873 B.n872 10.6151
R1633 B.n872 B.n81 10.6151
R1634 B.n866 B.n81 10.6151
R1635 B.n866 B.n865 10.6151
R1636 B.n865 B.n864 10.6151
R1637 B.n141 B.n88 10.6151
R1638 B.n144 B.n141 10.6151
R1639 B.n145 B.n144 10.6151
R1640 B.n148 B.n145 10.6151
R1641 B.n149 B.n148 10.6151
R1642 B.n152 B.n149 10.6151
R1643 B.n153 B.n152 10.6151
R1644 B.n156 B.n153 10.6151
R1645 B.n157 B.n156 10.6151
R1646 B.n160 B.n157 10.6151
R1647 B.n161 B.n160 10.6151
R1648 B.n164 B.n161 10.6151
R1649 B.n165 B.n164 10.6151
R1650 B.n168 B.n165 10.6151
R1651 B.n169 B.n168 10.6151
R1652 B.n172 B.n169 10.6151
R1653 B.n173 B.n172 10.6151
R1654 B.n176 B.n173 10.6151
R1655 B.n177 B.n176 10.6151
R1656 B.n180 B.n177 10.6151
R1657 B.n181 B.n180 10.6151
R1658 B.n184 B.n181 10.6151
R1659 B.n185 B.n184 10.6151
R1660 B.n188 B.n185 10.6151
R1661 B.n189 B.n188 10.6151
R1662 B.n192 B.n189 10.6151
R1663 B.n193 B.n192 10.6151
R1664 B.n196 B.n193 10.6151
R1665 B.n197 B.n196 10.6151
R1666 B.n200 B.n197 10.6151
R1667 B.n201 B.n200 10.6151
R1668 B.n204 B.n201 10.6151
R1669 B.n205 B.n204 10.6151
R1670 B.n208 B.n205 10.6151
R1671 B.n209 B.n208 10.6151
R1672 B.n212 B.n209 10.6151
R1673 B.n213 B.n212 10.6151
R1674 B.n216 B.n213 10.6151
R1675 B.n217 B.n216 10.6151
R1676 B.n220 B.n217 10.6151
R1677 B.n225 B.n222 10.6151
R1678 B.n226 B.n225 10.6151
R1679 B.n229 B.n226 10.6151
R1680 B.n230 B.n229 10.6151
R1681 B.n233 B.n230 10.6151
R1682 B.n234 B.n233 10.6151
R1683 B.n237 B.n234 10.6151
R1684 B.n238 B.n237 10.6151
R1685 B.n241 B.n238 10.6151
R1686 B.n246 B.n243 10.6151
R1687 B.n247 B.n246 10.6151
R1688 B.n250 B.n247 10.6151
R1689 B.n251 B.n250 10.6151
R1690 B.n254 B.n251 10.6151
R1691 B.n255 B.n254 10.6151
R1692 B.n258 B.n255 10.6151
R1693 B.n259 B.n258 10.6151
R1694 B.n262 B.n259 10.6151
R1695 B.n263 B.n262 10.6151
R1696 B.n266 B.n263 10.6151
R1697 B.n267 B.n266 10.6151
R1698 B.n270 B.n267 10.6151
R1699 B.n271 B.n270 10.6151
R1700 B.n274 B.n271 10.6151
R1701 B.n275 B.n274 10.6151
R1702 B.n278 B.n275 10.6151
R1703 B.n279 B.n278 10.6151
R1704 B.n282 B.n279 10.6151
R1705 B.n283 B.n282 10.6151
R1706 B.n286 B.n283 10.6151
R1707 B.n287 B.n286 10.6151
R1708 B.n290 B.n287 10.6151
R1709 B.n291 B.n290 10.6151
R1710 B.n294 B.n291 10.6151
R1711 B.n295 B.n294 10.6151
R1712 B.n298 B.n295 10.6151
R1713 B.n299 B.n298 10.6151
R1714 B.n302 B.n299 10.6151
R1715 B.n303 B.n302 10.6151
R1716 B.n306 B.n303 10.6151
R1717 B.n307 B.n306 10.6151
R1718 B.n310 B.n307 10.6151
R1719 B.n311 B.n310 10.6151
R1720 B.n314 B.n311 10.6151
R1721 B.n315 B.n314 10.6151
R1722 B.n318 B.n315 10.6151
R1723 B.n320 B.n318 10.6151
R1724 B.n321 B.n320 10.6151
R1725 B.n858 B.n321 10.6151
R1726 B.n446 B.n445 9.36635
R1727 B.n567 B.n566 9.36635
R1728 B.n221 B.n220 9.36635
R1729 B.n243 B.n242 9.36635
R1730 B.n962 B.n0 8.11757
R1731 B.n962 B.n1 8.11757
R1732 B.n778 B.t0 7.09104
R1733 B.n948 B.t2 7.09104
R1734 B.n548 B.n445 1.24928
R1735 B.n566 B.n565 1.24928
R1736 B.n222 B.n221 1.24928
R1737 B.n242 B.n241 1.24928
R1738 VP.n13 VP.n10 161.3
R1739 VP.n15 VP.n14 161.3
R1740 VP.n16 VP.n9 161.3
R1741 VP.n18 VP.n17 161.3
R1742 VP.n19 VP.n8 161.3
R1743 VP.n21 VP.n20 161.3
R1744 VP.n44 VP.n43 161.3
R1745 VP.n42 VP.n1 161.3
R1746 VP.n41 VP.n40 161.3
R1747 VP.n39 VP.n2 161.3
R1748 VP.n38 VP.n37 161.3
R1749 VP.n36 VP.n3 161.3
R1750 VP.n35 VP.n34 161.3
R1751 VP.n33 VP.n4 161.3
R1752 VP.n32 VP.n31 161.3
R1753 VP.n30 VP.n5 161.3
R1754 VP.n29 VP.n28 161.3
R1755 VP.n27 VP.n6 161.3
R1756 VP.n26 VP.n25 161.3
R1757 VP.n11 VP.t2 124.781
R1758 VP.n35 VP.t3 91.3635
R1759 VP.n24 VP.t5 91.3635
R1760 VP.n0 VP.t1 91.3635
R1761 VP.n12 VP.t0 91.3635
R1762 VP.n7 VP.t4 91.3635
R1763 VP.n24 VP.n23 68.5364
R1764 VP.n45 VP.n0 68.5364
R1765 VP.n22 VP.n7 68.5364
R1766 VP.n30 VP.n29 56.5193
R1767 VP.n41 VP.n2 56.5193
R1768 VP.n18 VP.n9 56.5193
R1769 VP.n23 VP.n22 50.6887
R1770 VP.n12 VP.n11 49.4728
R1771 VP.n25 VP.n6 24.4675
R1772 VP.n29 VP.n6 24.4675
R1773 VP.n31 VP.n30 24.4675
R1774 VP.n31 VP.n4 24.4675
R1775 VP.n35 VP.n4 24.4675
R1776 VP.n36 VP.n35 24.4675
R1777 VP.n37 VP.n36 24.4675
R1778 VP.n37 VP.n2 24.4675
R1779 VP.n42 VP.n41 24.4675
R1780 VP.n43 VP.n42 24.4675
R1781 VP.n19 VP.n18 24.4675
R1782 VP.n20 VP.n19 24.4675
R1783 VP.n13 VP.n12 24.4675
R1784 VP.n14 VP.n13 24.4675
R1785 VP.n14 VP.n9 24.4675
R1786 VP.n25 VP.n24 21.5315
R1787 VP.n43 VP.n0 21.5315
R1788 VP.n20 VP.n7 21.5315
R1789 VP.n11 VP.n10 3.84097
R1790 VP.n22 VP.n21 0.354971
R1791 VP.n26 VP.n23 0.354971
R1792 VP.n45 VP.n44 0.354971
R1793 VP VP.n45 0.26696
R1794 VP.n15 VP.n10 0.189894
R1795 VP.n16 VP.n15 0.189894
R1796 VP.n17 VP.n16 0.189894
R1797 VP.n17 VP.n8 0.189894
R1798 VP.n21 VP.n8 0.189894
R1799 VP.n27 VP.n26 0.189894
R1800 VP.n28 VP.n27 0.189894
R1801 VP.n28 VP.n5 0.189894
R1802 VP.n32 VP.n5 0.189894
R1803 VP.n33 VP.n32 0.189894
R1804 VP.n34 VP.n33 0.189894
R1805 VP.n34 VP.n3 0.189894
R1806 VP.n38 VP.n3 0.189894
R1807 VP.n39 VP.n38 0.189894
R1808 VP.n40 VP.n39 0.189894
R1809 VP.n40 VP.n1 0.189894
R1810 VP.n44 VP.n1 0.189894
R1811 VDD1 VDD1.t3 66.5236
R1812 VDD1.n1 VDD1.t0 66.4098
R1813 VDD1.n1 VDD1.n0 63.2476
R1814 VDD1.n3 VDD1.n2 62.5617
R1815 VDD1.n3 VDD1.n1 45.5828
R1816 VDD1.n2 VDD1.t5 1.67989
R1817 VDD1.n2 VDD1.t1 1.67989
R1818 VDD1.n0 VDD1.t2 1.67989
R1819 VDD1.n0 VDD1.t4 1.67989
R1820 VDD1 VDD1.n3 0.68369
C0 VTAIL VP 7.12796f
C1 VN VP 7.382871f
C2 VP VDD2 0.501634f
C3 VTAIL VN 7.113709f
C4 VTAIL VDD2 7.84893f
C5 VN VDD2 6.82153f
C6 VDD1 VP 7.168581f
C7 VTAIL VDD1 7.79416f
C8 VN VDD1 0.151525f
C9 VDD1 VDD2 1.60648f
C10 VDD2 B 6.336493f
C11 VDD1 B 6.68961f
C12 VTAIL B 8.067971f
C13 VN B 14.365701f
C14 VP B 13.047493f
C15 VDD1.t3 B 2.31188f
C16 VDD1.t0 B 2.31096f
C17 VDD1.t2 B 0.202426f
C18 VDD1.t4 B 0.202426f
C19 VDD1.n0 B 1.80702f
C20 VDD1.n1 B 2.8248f
C21 VDD1.t5 B 0.202426f
C22 VDD1.t1 B 0.202426f
C23 VDD1.n2 B 1.8022f
C24 VDD1.n3 B 2.53569f
C25 VP.t1 B 2.11865f
C26 VP.n0 B 0.835177f
C27 VP.n1 B 0.021218f
C28 VP.n2 B 0.0292f
C29 VP.n3 B 0.021218f
C30 VP.t3 B 2.11865f
C31 VP.n4 B 0.039545f
C32 VP.n5 B 0.021218f
C33 VP.n6 B 0.039545f
C34 VP.t4 B 2.11865f
C35 VP.n7 B 0.835177f
C36 VP.n8 B 0.021218f
C37 VP.n9 B 0.0292f
C38 VP.n10 B 0.241369f
C39 VP.t0 B 2.11865f
C40 VP.t2 B 2.35943f
C41 VP.n11 B 0.782325f
C42 VP.n12 B 0.826298f
C43 VP.n13 B 0.039545f
C44 VP.n14 B 0.039545f
C45 VP.n15 B 0.021218f
C46 VP.n16 B 0.021218f
C47 VP.n17 B 0.021218f
C48 VP.n18 B 0.032748f
C49 VP.n19 B 0.039545f
C50 VP.n20 B 0.037202f
C51 VP.n21 B 0.034245f
C52 VP.n22 B 1.22367f
C53 VP.n23 B 1.23871f
C54 VP.t5 B 2.11865f
C55 VP.n24 B 0.835177f
C56 VP.n25 B 0.037202f
C57 VP.n26 B 0.034245f
C58 VP.n27 B 0.021218f
C59 VP.n28 B 0.021218f
C60 VP.n29 B 0.032748f
C61 VP.n30 B 0.0292f
C62 VP.n31 B 0.039545f
C63 VP.n32 B 0.021218f
C64 VP.n33 B 0.021218f
C65 VP.n34 B 0.021218f
C66 VP.n35 B 0.76631f
C67 VP.n36 B 0.039545f
C68 VP.n37 B 0.039545f
C69 VP.n38 B 0.021218f
C70 VP.n39 B 0.021218f
C71 VP.n40 B 0.021218f
C72 VP.n41 B 0.032748f
C73 VP.n42 B 0.039545f
C74 VP.n43 B 0.037202f
C75 VP.n44 B 0.034245f
C76 VP.n45 B 0.04334f
C77 VDD2.t5 B 2.26143f
C78 VDD2.t4 B 0.198088f
C79 VDD2.t1 B 0.198088f
C80 VDD2.n0 B 1.76829f
C81 VDD2.n1 B 2.64742f
C82 VDD2.t3 B 2.24877f
C83 VDD2.n2 B 2.48109f
C84 VDD2.t2 B 0.198088f
C85 VDD2.t0 B 0.198088f
C86 VDD2.n3 B 1.76826f
C87 VTAIL.t9 B 0.224059f
C88 VTAIL.t7 B 0.224059f
C89 VTAIL.n0 B 1.92436f
C90 VTAIL.n1 B 0.44937f
C91 VTAIL.t0 B 2.45382f
C92 VTAIL.n2 B 0.698825f
C93 VTAIL.t4 B 0.224059f
C94 VTAIL.t1 B 0.224059f
C95 VTAIL.n3 B 1.92436f
C96 VTAIL.n4 B 2.03978f
C97 VTAIL.t10 B 0.224059f
C98 VTAIL.t8 B 0.224059f
C99 VTAIL.n5 B 1.92437f
C100 VTAIL.n6 B 2.03978f
C101 VTAIL.t6 B 2.45382f
C102 VTAIL.n7 B 0.698819f
C103 VTAIL.t2 B 0.224059f
C104 VTAIL.t3 B 0.224059f
C105 VTAIL.n8 B 1.92437f
C106 VTAIL.n9 B 0.617205f
C107 VTAIL.t5 B 2.45382f
C108 VTAIL.n10 B 1.8916f
C109 VTAIL.t11 B 2.45382f
C110 VTAIL.n11 B 1.82964f
C111 VN.t4 B 2.07675f
C112 VN.n0 B 0.818657f
C113 VN.n1 B 0.020798f
C114 VN.n2 B 0.028623f
C115 VN.n3 B 0.236595f
C116 VN.t1 B 2.07675f
C117 VN.t0 B 2.31277f
C118 VN.n4 B 0.76685f
C119 VN.n5 B 0.809954f
C120 VN.n6 B 0.038763f
C121 VN.n7 B 0.038763f
C122 VN.n8 B 0.020798f
C123 VN.n9 B 0.020798f
C124 VN.n10 B 0.020798f
C125 VN.n11 B 0.0321f
C126 VN.n12 B 0.038763f
C127 VN.n13 B 0.036466f
C128 VN.n14 B 0.033568f
C129 VN.n15 B 0.042483f
C130 VN.t2 B 2.07675f
C131 VN.n16 B 0.818657f
C132 VN.n17 B 0.020798f
C133 VN.n18 B 0.028623f
C134 VN.n19 B 0.236595f
C135 VN.t3 B 2.07675f
C136 VN.t5 B 2.31277f
C137 VN.n20 B 0.76685f
C138 VN.n21 B 0.809954f
C139 VN.n22 B 0.038763f
C140 VN.n23 B 0.038763f
C141 VN.n24 B 0.020798f
C142 VN.n25 B 0.020798f
C143 VN.n26 B 0.020798f
C144 VN.n27 B 0.0321f
C145 VN.n28 B 0.038763f
C146 VN.n29 B 0.036466f
C147 VN.n30 B 0.033568f
C148 VN.n31 B 1.20793f
.ends

