* NGSPICE file created from diff_pair_sample_1263.ext - technology: sky130A

.subckt diff_pair_sample_1263 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t12 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=1.9968 ps=11.02 w=5.12 l=2.16
X1 VTAIL.t0 VN.t0 VDD2.t9 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X2 VDD2.t8 VN.t1 VTAIL.t3 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=1.9968 ps=11.02 w=5.12 l=2.16
X3 VDD1.t8 VP.t1 VTAIL.t10 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X4 VTAIL.t14 VP.t2 VDD1.t7 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X5 VDD1.t6 VP.t3 VTAIL.t15 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0.8448 ps=5.45 w=5.12 l=2.16
X6 VDD2.t7 VN.t2 VTAIL.t1 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0.8448 ps=5.45 w=5.12 l=2.16
X7 B.t11 B.t9 B.t10 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0 ps=0 w=5.12 l=2.16
X8 VDD2.t6 VN.t3 VTAIL.t17 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=1.9968 ps=11.02 w=5.12 l=2.16
X9 B.t8 B.t6 B.t7 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0 ps=0 w=5.12 l=2.16
X10 VTAIL.t2 VN.t4 VDD2.t5 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X11 VTAIL.t5 VN.t5 VDD2.t4 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X12 B.t5 B.t3 B.t4 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0 ps=0 w=5.12 l=2.16
X13 VDD1.t5 VP.t4 VTAIL.t11 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0.8448 ps=5.45 w=5.12 l=2.16
X14 VDD1.t4 VP.t5 VTAIL.t7 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=1.9968 ps=11.02 w=5.12 l=2.16
X15 VTAIL.t13 VP.t6 VDD1.t3 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X16 VTAIL.t8 VP.t7 VDD1.t2 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X17 VDD2.t3 VN.t6 VTAIL.t4 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X18 VDD2.t2 VN.t7 VTAIL.t6 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X19 VDD2.t1 VN.t8 VTAIL.t18 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0.8448 ps=5.45 w=5.12 l=2.16
X20 VTAIL.t19 VN.t9 VDD2.t0 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X21 VTAIL.t9 VP.t8 VDD1.t1 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X22 VDD1.t0 VP.t9 VTAIL.t16 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=0.8448 pd=5.45 as=0.8448 ps=5.45 w=5.12 l=2.16
X23 B.t2 B.t0 B.t1 w_n3958_n1992# sky130_fd_pr__pfet_01v8 ad=1.9968 pd=11.02 as=0 ps=0 w=5.12 l=2.16
R0 VP.n22 VP.n21 161.3
R1 VP.n23 VP.n18 161.3
R2 VP.n25 VP.n24 161.3
R3 VP.n26 VP.n17 161.3
R4 VP.n28 VP.n27 161.3
R5 VP.n30 VP.n29 161.3
R6 VP.n31 VP.n15 161.3
R7 VP.n33 VP.n32 161.3
R8 VP.n34 VP.n14 161.3
R9 VP.n36 VP.n35 161.3
R10 VP.n38 VP.n13 161.3
R11 VP.n40 VP.n39 161.3
R12 VP.n41 VP.n12 161.3
R13 VP.n43 VP.n42 161.3
R14 VP.n44 VP.n11 161.3
R15 VP.n80 VP.n0 161.3
R16 VP.n79 VP.n78 161.3
R17 VP.n77 VP.n1 161.3
R18 VP.n76 VP.n75 161.3
R19 VP.n74 VP.n2 161.3
R20 VP.n72 VP.n71 161.3
R21 VP.n70 VP.n3 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n67 VP.n4 161.3
R24 VP.n66 VP.n65 161.3
R25 VP.n64 VP.n63 161.3
R26 VP.n62 VP.n6 161.3
R27 VP.n61 VP.n60 161.3
R28 VP.n59 VP.n7 161.3
R29 VP.n58 VP.n57 161.3
R30 VP.n55 VP.n8 161.3
R31 VP.n54 VP.n53 161.3
R32 VP.n52 VP.n9 161.3
R33 VP.n51 VP.n50 161.3
R34 VP.n49 VP.n10 161.3
R35 VP.n48 VP.n47 99.596
R36 VP.n82 VP.n81 99.596
R37 VP.n46 VP.n45 99.596
R38 VP.n19 VP.t4 88.8788
R39 VP.n20 VP.n19 59.9481
R40 VP.n48 VP.t3 57.1264
R41 VP.n56 VP.t2 57.1264
R42 VP.n5 VP.t1 57.1264
R43 VP.n73 VP.t8 57.1264
R44 VP.n81 VP.t5 57.1264
R45 VP.n45 VP.t0 57.1264
R46 VP.n37 VP.t7 57.1264
R47 VP.n16 VP.t9 57.1264
R48 VP.n20 VP.t6 57.1264
R49 VP.n47 VP.n46 45.4428
R50 VP.n54 VP.n9 42.0302
R51 VP.n75 VP.n1 42.0302
R52 VP.n39 VP.n12 42.0302
R53 VP.n62 VP.n61 41.0614
R54 VP.n68 VP.n67 41.0614
R55 VP.n32 VP.n31 41.0614
R56 VP.n26 VP.n25 41.0614
R57 VP.n61 VP.n7 40.0926
R58 VP.n68 VP.n3 40.0926
R59 VP.n32 VP.n14 40.0926
R60 VP.n25 VP.n18 40.0926
R61 VP.n50 VP.n9 39.1239
R62 VP.n79 VP.n1 39.1239
R63 VP.n43 VP.n12 39.1239
R64 VP.n50 VP.n49 24.5923
R65 VP.n55 VP.n54 24.5923
R66 VP.n57 VP.n7 24.5923
R67 VP.n63 VP.n62 24.5923
R68 VP.n67 VP.n66 24.5923
R69 VP.n72 VP.n3 24.5923
R70 VP.n75 VP.n74 24.5923
R71 VP.n80 VP.n79 24.5923
R72 VP.n44 VP.n43 24.5923
R73 VP.n36 VP.n14 24.5923
R74 VP.n39 VP.n38 24.5923
R75 VP.n27 VP.n26 24.5923
R76 VP.n31 VP.n30 24.5923
R77 VP.n21 VP.n18 24.5923
R78 VP.n56 VP.n55 12.7883
R79 VP.n74 VP.n73 12.7883
R80 VP.n38 VP.n37 12.7883
R81 VP.n63 VP.n5 12.2964
R82 VP.n66 VP.n5 12.2964
R83 VP.n27 VP.n16 12.2964
R84 VP.n30 VP.n16 12.2964
R85 VP.n57 VP.n56 11.8046
R86 VP.n73 VP.n72 11.8046
R87 VP.n37 VP.n36 11.8046
R88 VP.n21 VP.n20 11.8046
R89 VP.n49 VP.n48 11.3127
R90 VP.n81 VP.n80 11.3127
R91 VP.n45 VP.n44 11.3127
R92 VP.n22 VP.n19 9.80572
R93 VP.n46 VP.n11 0.278335
R94 VP.n47 VP.n10 0.278335
R95 VP.n82 VP.n0 0.278335
R96 VP.n23 VP.n22 0.189894
R97 VP.n24 VP.n23 0.189894
R98 VP.n24 VP.n17 0.189894
R99 VP.n28 VP.n17 0.189894
R100 VP.n29 VP.n28 0.189894
R101 VP.n29 VP.n15 0.189894
R102 VP.n33 VP.n15 0.189894
R103 VP.n34 VP.n33 0.189894
R104 VP.n35 VP.n34 0.189894
R105 VP.n35 VP.n13 0.189894
R106 VP.n40 VP.n13 0.189894
R107 VP.n41 VP.n40 0.189894
R108 VP.n42 VP.n41 0.189894
R109 VP.n42 VP.n11 0.189894
R110 VP.n51 VP.n10 0.189894
R111 VP.n52 VP.n51 0.189894
R112 VP.n53 VP.n52 0.189894
R113 VP.n53 VP.n8 0.189894
R114 VP.n58 VP.n8 0.189894
R115 VP.n59 VP.n58 0.189894
R116 VP.n60 VP.n59 0.189894
R117 VP.n60 VP.n6 0.189894
R118 VP.n64 VP.n6 0.189894
R119 VP.n65 VP.n64 0.189894
R120 VP.n65 VP.n4 0.189894
R121 VP.n69 VP.n4 0.189894
R122 VP.n70 VP.n69 0.189894
R123 VP.n71 VP.n70 0.189894
R124 VP.n71 VP.n2 0.189894
R125 VP.n76 VP.n2 0.189894
R126 VP.n77 VP.n76 0.189894
R127 VP.n78 VP.n77 0.189894
R128 VP.n78 VP.n0 0.189894
R129 VP VP.n82 0.153485
R130 VTAIL.n116 VTAIL.n115 756.745
R131 VTAIL.n26 VTAIL.n25 756.745
R132 VTAIL.n90 VTAIL.n89 756.745
R133 VTAIL.n60 VTAIL.n59 756.745
R134 VTAIL.n101 VTAIL.n100 585
R135 VTAIL.n98 VTAIL.n97 585
R136 VTAIL.n107 VTAIL.n106 585
R137 VTAIL.n109 VTAIL.n108 585
R138 VTAIL.n94 VTAIL.n93 585
R139 VTAIL.n115 VTAIL.n114 585
R140 VTAIL.n11 VTAIL.n10 585
R141 VTAIL.n8 VTAIL.n7 585
R142 VTAIL.n17 VTAIL.n16 585
R143 VTAIL.n19 VTAIL.n18 585
R144 VTAIL.n4 VTAIL.n3 585
R145 VTAIL.n25 VTAIL.n24 585
R146 VTAIL.n89 VTAIL.n88 585
R147 VTAIL.n68 VTAIL.n67 585
R148 VTAIL.n83 VTAIL.n82 585
R149 VTAIL.n81 VTAIL.n80 585
R150 VTAIL.n72 VTAIL.n71 585
R151 VTAIL.n75 VTAIL.n74 585
R152 VTAIL.n59 VTAIL.n58 585
R153 VTAIL.n38 VTAIL.n37 585
R154 VTAIL.n53 VTAIL.n52 585
R155 VTAIL.n51 VTAIL.n50 585
R156 VTAIL.n42 VTAIL.n41 585
R157 VTAIL.n45 VTAIL.n44 585
R158 VTAIL.t12 VTAIL.n73 329.435
R159 VTAIL.t3 VTAIL.n99 329.435
R160 VTAIL.t7 VTAIL.n9 329.435
R161 VTAIL.t17 VTAIL.n43 329.435
R162 VTAIL.n100 VTAIL.n97 171.744
R163 VTAIL.n107 VTAIL.n97 171.744
R164 VTAIL.n108 VTAIL.n107 171.744
R165 VTAIL.n108 VTAIL.n93 171.744
R166 VTAIL.n115 VTAIL.n93 171.744
R167 VTAIL.n10 VTAIL.n7 171.744
R168 VTAIL.n17 VTAIL.n7 171.744
R169 VTAIL.n18 VTAIL.n17 171.744
R170 VTAIL.n18 VTAIL.n3 171.744
R171 VTAIL.n25 VTAIL.n3 171.744
R172 VTAIL.n89 VTAIL.n67 171.744
R173 VTAIL.n82 VTAIL.n67 171.744
R174 VTAIL.n82 VTAIL.n81 171.744
R175 VTAIL.n81 VTAIL.n71 171.744
R176 VTAIL.n74 VTAIL.n71 171.744
R177 VTAIL.n59 VTAIL.n37 171.744
R178 VTAIL.n52 VTAIL.n37 171.744
R179 VTAIL.n52 VTAIL.n51 171.744
R180 VTAIL.n51 VTAIL.n41 171.744
R181 VTAIL.n44 VTAIL.n41 171.744
R182 VTAIL.n100 VTAIL.t3 85.8723
R183 VTAIL.n10 VTAIL.t7 85.8723
R184 VTAIL.n74 VTAIL.t12 85.8723
R185 VTAIL.n44 VTAIL.t17 85.8723
R186 VTAIL.n65 VTAIL.n64 83.699
R187 VTAIL.n63 VTAIL.n62 83.699
R188 VTAIL.n35 VTAIL.n34 83.699
R189 VTAIL.n33 VTAIL.n32 83.699
R190 VTAIL.n119 VTAIL.n118 83.6989
R191 VTAIL.n1 VTAIL.n0 83.6989
R192 VTAIL.n29 VTAIL.n28 83.6989
R193 VTAIL.n31 VTAIL.n30 83.6989
R194 VTAIL.n117 VTAIL.n116 34.1247
R195 VTAIL.n27 VTAIL.n26 34.1247
R196 VTAIL.n91 VTAIL.n90 34.1247
R197 VTAIL.n61 VTAIL.n60 34.1247
R198 VTAIL.n33 VTAIL.n31 21.0738
R199 VTAIL.n117 VTAIL.n91 18.9272
R200 VTAIL.n114 VTAIL.n92 11.249
R201 VTAIL.n24 VTAIL.n2 11.249
R202 VTAIL.n88 VTAIL.n66 11.249
R203 VTAIL.n58 VTAIL.n36 11.249
R204 VTAIL.n101 VTAIL.n99 10.7185
R205 VTAIL.n11 VTAIL.n9 10.7185
R206 VTAIL.n75 VTAIL.n73 10.7185
R207 VTAIL.n45 VTAIL.n43 10.7185
R208 VTAIL.n113 VTAIL.n94 10.4732
R209 VTAIL.n23 VTAIL.n4 10.4732
R210 VTAIL.n87 VTAIL.n68 10.4732
R211 VTAIL.n57 VTAIL.n38 10.4732
R212 VTAIL.n110 VTAIL.n109 9.69747
R213 VTAIL.n20 VTAIL.n19 9.69747
R214 VTAIL.n84 VTAIL.n83 9.69747
R215 VTAIL.n54 VTAIL.n53 9.69747
R216 VTAIL.n112 VTAIL.n92 9.45567
R217 VTAIL.n22 VTAIL.n2 9.45567
R218 VTAIL.n86 VTAIL.n66 9.45567
R219 VTAIL.n56 VTAIL.n36 9.45567
R220 VTAIL.n103 VTAIL.n102 9.3005
R221 VTAIL.n105 VTAIL.n104 9.3005
R222 VTAIL.n96 VTAIL.n95 9.3005
R223 VTAIL.n111 VTAIL.n110 9.3005
R224 VTAIL.n113 VTAIL.n112 9.3005
R225 VTAIL.n13 VTAIL.n12 9.3005
R226 VTAIL.n15 VTAIL.n14 9.3005
R227 VTAIL.n6 VTAIL.n5 9.3005
R228 VTAIL.n21 VTAIL.n20 9.3005
R229 VTAIL.n23 VTAIL.n22 9.3005
R230 VTAIL.n87 VTAIL.n86 9.3005
R231 VTAIL.n85 VTAIL.n84 9.3005
R232 VTAIL.n70 VTAIL.n69 9.3005
R233 VTAIL.n79 VTAIL.n78 9.3005
R234 VTAIL.n77 VTAIL.n76 9.3005
R235 VTAIL.n49 VTAIL.n48 9.3005
R236 VTAIL.n40 VTAIL.n39 9.3005
R237 VTAIL.n55 VTAIL.n54 9.3005
R238 VTAIL.n57 VTAIL.n56 9.3005
R239 VTAIL.n47 VTAIL.n46 9.3005
R240 VTAIL.n106 VTAIL.n96 8.92171
R241 VTAIL.n16 VTAIL.n6 8.92171
R242 VTAIL.n80 VTAIL.n70 8.92171
R243 VTAIL.n50 VTAIL.n40 8.92171
R244 VTAIL.n105 VTAIL.n98 8.14595
R245 VTAIL.n15 VTAIL.n8 8.14595
R246 VTAIL.n79 VTAIL.n72 8.14595
R247 VTAIL.n49 VTAIL.n42 8.14595
R248 VTAIL.n102 VTAIL.n101 7.3702
R249 VTAIL.n12 VTAIL.n11 7.3702
R250 VTAIL.n76 VTAIL.n75 7.3702
R251 VTAIL.n46 VTAIL.n45 7.3702
R252 VTAIL.n118 VTAIL.t6 6.34913
R253 VTAIL.n118 VTAIL.t19 6.34913
R254 VTAIL.n0 VTAIL.t1 6.34913
R255 VTAIL.n0 VTAIL.t2 6.34913
R256 VTAIL.n28 VTAIL.t10 6.34913
R257 VTAIL.n28 VTAIL.t9 6.34913
R258 VTAIL.n30 VTAIL.t15 6.34913
R259 VTAIL.n30 VTAIL.t14 6.34913
R260 VTAIL.n64 VTAIL.t16 6.34913
R261 VTAIL.n64 VTAIL.t8 6.34913
R262 VTAIL.n62 VTAIL.t11 6.34913
R263 VTAIL.n62 VTAIL.t13 6.34913
R264 VTAIL.n34 VTAIL.t4 6.34913
R265 VTAIL.n34 VTAIL.t5 6.34913
R266 VTAIL.n32 VTAIL.t18 6.34913
R267 VTAIL.n32 VTAIL.t0 6.34913
R268 VTAIL.n102 VTAIL.n98 5.81868
R269 VTAIL.n12 VTAIL.n8 5.81868
R270 VTAIL.n76 VTAIL.n72 5.81868
R271 VTAIL.n46 VTAIL.n42 5.81868
R272 VTAIL.n106 VTAIL.n105 5.04292
R273 VTAIL.n16 VTAIL.n15 5.04292
R274 VTAIL.n80 VTAIL.n79 5.04292
R275 VTAIL.n50 VTAIL.n49 5.04292
R276 VTAIL.n109 VTAIL.n96 4.26717
R277 VTAIL.n19 VTAIL.n6 4.26717
R278 VTAIL.n83 VTAIL.n70 4.26717
R279 VTAIL.n53 VTAIL.n40 4.26717
R280 VTAIL.n110 VTAIL.n94 3.49141
R281 VTAIL.n20 VTAIL.n4 3.49141
R282 VTAIL.n84 VTAIL.n68 3.49141
R283 VTAIL.n54 VTAIL.n38 3.49141
R284 VTAIL.n114 VTAIL.n113 2.71565
R285 VTAIL.n24 VTAIL.n23 2.71565
R286 VTAIL.n88 VTAIL.n87 2.71565
R287 VTAIL.n58 VTAIL.n57 2.71565
R288 VTAIL.n103 VTAIL.n99 2.41827
R289 VTAIL.n13 VTAIL.n9 2.41827
R290 VTAIL.n77 VTAIL.n73 2.41827
R291 VTAIL.n47 VTAIL.n43 2.41827
R292 VTAIL.n35 VTAIL.n33 2.14705
R293 VTAIL.n61 VTAIL.n35 2.14705
R294 VTAIL.n65 VTAIL.n63 2.14705
R295 VTAIL.n91 VTAIL.n65 2.14705
R296 VTAIL.n31 VTAIL.n29 2.14705
R297 VTAIL.n29 VTAIL.n27 2.14705
R298 VTAIL.n119 VTAIL.n117 2.14705
R299 VTAIL.n116 VTAIL.n92 1.93989
R300 VTAIL.n26 VTAIL.n2 1.93989
R301 VTAIL.n90 VTAIL.n66 1.93989
R302 VTAIL.n60 VTAIL.n36 1.93989
R303 VTAIL VTAIL.n1 1.6686
R304 VTAIL.n63 VTAIL.n61 1.5436
R305 VTAIL.n27 VTAIL.n1 1.5436
R306 VTAIL VTAIL.n119 0.478948
R307 VTAIL.n104 VTAIL.n103 0.155672
R308 VTAIL.n104 VTAIL.n95 0.155672
R309 VTAIL.n111 VTAIL.n95 0.155672
R310 VTAIL.n112 VTAIL.n111 0.155672
R311 VTAIL.n14 VTAIL.n13 0.155672
R312 VTAIL.n14 VTAIL.n5 0.155672
R313 VTAIL.n21 VTAIL.n5 0.155672
R314 VTAIL.n22 VTAIL.n21 0.155672
R315 VTAIL.n86 VTAIL.n85 0.155672
R316 VTAIL.n85 VTAIL.n69 0.155672
R317 VTAIL.n78 VTAIL.n69 0.155672
R318 VTAIL.n78 VTAIL.n77 0.155672
R319 VTAIL.n56 VTAIL.n55 0.155672
R320 VTAIL.n55 VTAIL.n39 0.155672
R321 VTAIL.n48 VTAIL.n39 0.155672
R322 VTAIL.n48 VTAIL.n47 0.155672
R323 VDD1.n24 VDD1.n23 756.745
R324 VDD1.n51 VDD1.n50 756.745
R325 VDD1.n23 VDD1.n22 585
R326 VDD1.n2 VDD1.n1 585
R327 VDD1.n17 VDD1.n16 585
R328 VDD1.n15 VDD1.n14 585
R329 VDD1.n6 VDD1.n5 585
R330 VDD1.n9 VDD1.n8 585
R331 VDD1.n36 VDD1.n35 585
R332 VDD1.n33 VDD1.n32 585
R333 VDD1.n42 VDD1.n41 585
R334 VDD1.n44 VDD1.n43 585
R335 VDD1.n29 VDD1.n28 585
R336 VDD1.n50 VDD1.n49 585
R337 VDD1.t5 VDD1.n7 329.435
R338 VDD1.t6 VDD1.n34 329.435
R339 VDD1.n23 VDD1.n1 171.744
R340 VDD1.n16 VDD1.n1 171.744
R341 VDD1.n16 VDD1.n15 171.744
R342 VDD1.n15 VDD1.n5 171.744
R343 VDD1.n8 VDD1.n5 171.744
R344 VDD1.n35 VDD1.n32 171.744
R345 VDD1.n42 VDD1.n32 171.744
R346 VDD1.n43 VDD1.n42 171.744
R347 VDD1.n43 VDD1.n28 171.744
R348 VDD1.n50 VDD1.n28 171.744
R349 VDD1.n55 VDD1.n54 101.933
R350 VDD1.n26 VDD1.n25 100.377
R351 VDD1.n53 VDD1.n52 100.377
R352 VDD1.n57 VDD1.n56 100.376
R353 VDD1.n8 VDD1.t5 85.8723
R354 VDD1.n35 VDD1.t6 85.8723
R355 VDD1.n26 VDD1.n24 52.9501
R356 VDD1.n53 VDD1.n51 52.9501
R357 VDD1.n57 VDD1.n55 39.9815
R358 VDD1.n22 VDD1.n0 11.249
R359 VDD1.n49 VDD1.n27 11.249
R360 VDD1.n9 VDD1.n7 10.7185
R361 VDD1.n36 VDD1.n34 10.7185
R362 VDD1.n21 VDD1.n2 10.4732
R363 VDD1.n48 VDD1.n29 10.4732
R364 VDD1.n18 VDD1.n17 9.69747
R365 VDD1.n45 VDD1.n44 9.69747
R366 VDD1.n20 VDD1.n0 9.45567
R367 VDD1.n47 VDD1.n27 9.45567
R368 VDD1.n13 VDD1.n12 9.3005
R369 VDD1.n4 VDD1.n3 9.3005
R370 VDD1.n19 VDD1.n18 9.3005
R371 VDD1.n21 VDD1.n20 9.3005
R372 VDD1.n11 VDD1.n10 9.3005
R373 VDD1.n38 VDD1.n37 9.3005
R374 VDD1.n40 VDD1.n39 9.3005
R375 VDD1.n31 VDD1.n30 9.3005
R376 VDD1.n46 VDD1.n45 9.3005
R377 VDD1.n48 VDD1.n47 9.3005
R378 VDD1.n14 VDD1.n4 8.92171
R379 VDD1.n41 VDD1.n31 8.92171
R380 VDD1.n13 VDD1.n6 8.14595
R381 VDD1.n40 VDD1.n33 8.14595
R382 VDD1.n10 VDD1.n9 7.3702
R383 VDD1.n37 VDD1.n36 7.3702
R384 VDD1.n56 VDD1.t2 6.34913
R385 VDD1.n56 VDD1.t9 6.34913
R386 VDD1.n25 VDD1.t3 6.34913
R387 VDD1.n25 VDD1.t0 6.34913
R388 VDD1.n54 VDD1.t1 6.34913
R389 VDD1.n54 VDD1.t4 6.34913
R390 VDD1.n52 VDD1.t7 6.34913
R391 VDD1.n52 VDD1.t8 6.34913
R392 VDD1.n10 VDD1.n6 5.81868
R393 VDD1.n37 VDD1.n33 5.81868
R394 VDD1.n14 VDD1.n13 5.04292
R395 VDD1.n41 VDD1.n40 5.04292
R396 VDD1.n17 VDD1.n4 4.26717
R397 VDD1.n44 VDD1.n31 4.26717
R398 VDD1.n18 VDD1.n2 3.49141
R399 VDD1.n45 VDD1.n29 3.49141
R400 VDD1.n22 VDD1.n21 2.71565
R401 VDD1.n49 VDD1.n48 2.71565
R402 VDD1.n11 VDD1.n7 2.41827
R403 VDD1.n38 VDD1.n34 2.41827
R404 VDD1.n24 VDD1.n0 1.93989
R405 VDD1.n51 VDD1.n27 1.93989
R406 VDD1 VDD1.n57 1.55222
R407 VDD1 VDD1.n26 0.595328
R408 VDD1.n55 VDD1.n53 0.481792
R409 VDD1.n20 VDD1.n19 0.155672
R410 VDD1.n19 VDD1.n3 0.155672
R411 VDD1.n12 VDD1.n3 0.155672
R412 VDD1.n12 VDD1.n11 0.155672
R413 VDD1.n39 VDD1.n38 0.155672
R414 VDD1.n39 VDD1.n30 0.155672
R415 VDD1.n46 VDD1.n30 0.155672
R416 VDD1.n47 VDD1.n46 0.155672
R417 VN.n69 VN.n36 161.3
R418 VN.n68 VN.n67 161.3
R419 VN.n66 VN.n37 161.3
R420 VN.n65 VN.n64 161.3
R421 VN.n63 VN.n38 161.3
R422 VN.n61 VN.n60 161.3
R423 VN.n59 VN.n39 161.3
R424 VN.n58 VN.n57 161.3
R425 VN.n56 VN.n40 161.3
R426 VN.n55 VN.n54 161.3
R427 VN.n53 VN.n52 161.3
R428 VN.n51 VN.n42 161.3
R429 VN.n50 VN.n49 161.3
R430 VN.n48 VN.n43 161.3
R431 VN.n47 VN.n46 161.3
R432 VN.n33 VN.n0 161.3
R433 VN.n32 VN.n31 161.3
R434 VN.n30 VN.n1 161.3
R435 VN.n29 VN.n28 161.3
R436 VN.n27 VN.n2 161.3
R437 VN.n25 VN.n24 161.3
R438 VN.n23 VN.n3 161.3
R439 VN.n22 VN.n21 161.3
R440 VN.n20 VN.n4 161.3
R441 VN.n19 VN.n18 161.3
R442 VN.n17 VN.n16 161.3
R443 VN.n15 VN.n6 161.3
R444 VN.n14 VN.n13 161.3
R445 VN.n12 VN.n7 161.3
R446 VN.n11 VN.n10 161.3
R447 VN.n35 VN.n34 99.596
R448 VN.n71 VN.n70 99.596
R449 VN.n8 VN.t2 88.8788
R450 VN.n44 VN.t3 88.8788
R451 VN.n9 VN.n8 59.9481
R452 VN.n45 VN.n44 59.9481
R453 VN.n9 VN.t4 57.1264
R454 VN.n5 VN.t7 57.1264
R455 VN.n26 VN.t9 57.1264
R456 VN.n34 VN.t1 57.1264
R457 VN.n45 VN.t5 57.1264
R458 VN.n41 VN.t6 57.1264
R459 VN.n62 VN.t0 57.1264
R460 VN.n70 VN.t8 57.1264
R461 VN VN.n71 45.7217
R462 VN.n28 VN.n1 42.0302
R463 VN.n64 VN.n37 42.0302
R464 VN.n15 VN.n14 41.0614
R465 VN.n21 VN.n20 41.0614
R466 VN.n51 VN.n50 41.0614
R467 VN.n57 VN.n56 41.0614
R468 VN.n14 VN.n7 40.0926
R469 VN.n21 VN.n3 40.0926
R470 VN.n50 VN.n43 40.0926
R471 VN.n57 VN.n39 40.0926
R472 VN.n32 VN.n1 39.1239
R473 VN.n68 VN.n37 39.1239
R474 VN.n10 VN.n7 24.5923
R475 VN.n16 VN.n15 24.5923
R476 VN.n20 VN.n19 24.5923
R477 VN.n25 VN.n3 24.5923
R478 VN.n28 VN.n27 24.5923
R479 VN.n33 VN.n32 24.5923
R480 VN.n46 VN.n43 24.5923
R481 VN.n56 VN.n55 24.5923
R482 VN.n52 VN.n51 24.5923
R483 VN.n64 VN.n63 24.5923
R484 VN.n61 VN.n39 24.5923
R485 VN.n69 VN.n68 24.5923
R486 VN.n27 VN.n26 12.7883
R487 VN.n63 VN.n62 12.7883
R488 VN.n16 VN.n5 12.2964
R489 VN.n19 VN.n5 12.2964
R490 VN.n55 VN.n41 12.2964
R491 VN.n52 VN.n41 12.2964
R492 VN.n10 VN.n9 11.8046
R493 VN.n26 VN.n25 11.8046
R494 VN.n46 VN.n45 11.8046
R495 VN.n62 VN.n61 11.8046
R496 VN.n34 VN.n33 11.3127
R497 VN.n70 VN.n69 11.3127
R498 VN.n47 VN.n44 9.80572
R499 VN.n11 VN.n8 9.80572
R500 VN.n71 VN.n36 0.278335
R501 VN.n35 VN.n0 0.278335
R502 VN.n67 VN.n36 0.189894
R503 VN.n67 VN.n66 0.189894
R504 VN.n66 VN.n65 0.189894
R505 VN.n65 VN.n38 0.189894
R506 VN.n60 VN.n38 0.189894
R507 VN.n60 VN.n59 0.189894
R508 VN.n59 VN.n58 0.189894
R509 VN.n58 VN.n40 0.189894
R510 VN.n54 VN.n40 0.189894
R511 VN.n54 VN.n53 0.189894
R512 VN.n53 VN.n42 0.189894
R513 VN.n49 VN.n42 0.189894
R514 VN.n49 VN.n48 0.189894
R515 VN.n48 VN.n47 0.189894
R516 VN.n12 VN.n11 0.189894
R517 VN.n13 VN.n12 0.189894
R518 VN.n13 VN.n6 0.189894
R519 VN.n17 VN.n6 0.189894
R520 VN.n18 VN.n17 0.189894
R521 VN.n18 VN.n4 0.189894
R522 VN.n22 VN.n4 0.189894
R523 VN.n23 VN.n22 0.189894
R524 VN.n24 VN.n23 0.189894
R525 VN.n24 VN.n2 0.189894
R526 VN.n29 VN.n2 0.189894
R527 VN.n30 VN.n29 0.189894
R528 VN.n31 VN.n30 0.189894
R529 VN.n31 VN.n0 0.189894
R530 VN VN.n35 0.153485
R531 VDD2.n53 VDD2.n52 756.745
R532 VDD2.n24 VDD2.n23 756.745
R533 VDD2.n52 VDD2.n51 585
R534 VDD2.n31 VDD2.n30 585
R535 VDD2.n46 VDD2.n45 585
R536 VDD2.n44 VDD2.n43 585
R537 VDD2.n35 VDD2.n34 585
R538 VDD2.n38 VDD2.n37 585
R539 VDD2.n9 VDD2.n8 585
R540 VDD2.n6 VDD2.n5 585
R541 VDD2.n15 VDD2.n14 585
R542 VDD2.n17 VDD2.n16 585
R543 VDD2.n2 VDD2.n1 585
R544 VDD2.n23 VDD2.n22 585
R545 VDD2.t1 VDD2.n36 329.435
R546 VDD2.t7 VDD2.n7 329.435
R547 VDD2.n52 VDD2.n30 171.744
R548 VDD2.n45 VDD2.n30 171.744
R549 VDD2.n45 VDD2.n44 171.744
R550 VDD2.n44 VDD2.n34 171.744
R551 VDD2.n37 VDD2.n34 171.744
R552 VDD2.n8 VDD2.n5 171.744
R553 VDD2.n15 VDD2.n5 171.744
R554 VDD2.n16 VDD2.n15 171.744
R555 VDD2.n16 VDD2.n1 171.744
R556 VDD2.n23 VDD2.n1 171.744
R557 VDD2.n28 VDD2.n27 101.933
R558 VDD2 VDD2.n57 101.928
R559 VDD2.n56 VDD2.n55 100.377
R560 VDD2.n26 VDD2.n25 100.377
R561 VDD2.n37 VDD2.t1 85.8723
R562 VDD2.n8 VDD2.t7 85.8723
R563 VDD2.n26 VDD2.n24 52.9501
R564 VDD2.n54 VDD2.n53 50.8035
R565 VDD2.n54 VDD2.n28 38.3252
R566 VDD2.n51 VDD2.n29 11.249
R567 VDD2.n22 VDD2.n0 11.249
R568 VDD2.n38 VDD2.n36 10.7185
R569 VDD2.n9 VDD2.n7 10.7185
R570 VDD2.n50 VDD2.n31 10.4732
R571 VDD2.n21 VDD2.n2 10.4732
R572 VDD2.n47 VDD2.n46 9.69747
R573 VDD2.n18 VDD2.n17 9.69747
R574 VDD2.n49 VDD2.n29 9.45567
R575 VDD2.n20 VDD2.n0 9.45567
R576 VDD2.n42 VDD2.n41 9.3005
R577 VDD2.n33 VDD2.n32 9.3005
R578 VDD2.n48 VDD2.n47 9.3005
R579 VDD2.n50 VDD2.n49 9.3005
R580 VDD2.n40 VDD2.n39 9.3005
R581 VDD2.n11 VDD2.n10 9.3005
R582 VDD2.n13 VDD2.n12 9.3005
R583 VDD2.n4 VDD2.n3 9.3005
R584 VDD2.n19 VDD2.n18 9.3005
R585 VDD2.n21 VDD2.n20 9.3005
R586 VDD2.n43 VDD2.n33 8.92171
R587 VDD2.n14 VDD2.n4 8.92171
R588 VDD2.n42 VDD2.n35 8.14595
R589 VDD2.n13 VDD2.n6 8.14595
R590 VDD2.n39 VDD2.n38 7.3702
R591 VDD2.n10 VDD2.n9 7.3702
R592 VDD2.n57 VDD2.t4 6.34913
R593 VDD2.n57 VDD2.t6 6.34913
R594 VDD2.n55 VDD2.t9 6.34913
R595 VDD2.n55 VDD2.t3 6.34913
R596 VDD2.n27 VDD2.t0 6.34913
R597 VDD2.n27 VDD2.t8 6.34913
R598 VDD2.n25 VDD2.t5 6.34913
R599 VDD2.n25 VDD2.t2 6.34913
R600 VDD2.n39 VDD2.n35 5.81868
R601 VDD2.n10 VDD2.n6 5.81868
R602 VDD2.n43 VDD2.n42 5.04292
R603 VDD2.n14 VDD2.n13 5.04292
R604 VDD2.n46 VDD2.n33 4.26717
R605 VDD2.n17 VDD2.n4 4.26717
R606 VDD2.n47 VDD2.n31 3.49141
R607 VDD2.n18 VDD2.n2 3.49141
R608 VDD2.n51 VDD2.n50 2.71565
R609 VDD2.n22 VDD2.n21 2.71565
R610 VDD2.n40 VDD2.n36 2.41827
R611 VDD2.n11 VDD2.n7 2.41827
R612 VDD2.n56 VDD2.n54 2.14705
R613 VDD2.n53 VDD2.n29 1.93989
R614 VDD2.n24 VDD2.n0 1.93989
R615 VDD2 VDD2.n56 0.595328
R616 VDD2.n28 VDD2.n26 0.481792
R617 VDD2.n49 VDD2.n48 0.155672
R618 VDD2.n48 VDD2.n32 0.155672
R619 VDD2.n41 VDD2.n32 0.155672
R620 VDD2.n41 VDD2.n40 0.155672
R621 VDD2.n12 VDD2.n11 0.155672
R622 VDD2.n12 VDD2.n3 0.155672
R623 VDD2.n19 VDD2.n3 0.155672
R624 VDD2.n20 VDD2.n19 0.155672
R625 B.n482 B.n481 585
R626 B.n483 B.n58 585
R627 B.n485 B.n484 585
R628 B.n486 B.n57 585
R629 B.n488 B.n487 585
R630 B.n489 B.n56 585
R631 B.n491 B.n490 585
R632 B.n492 B.n55 585
R633 B.n494 B.n493 585
R634 B.n495 B.n54 585
R635 B.n497 B.n496 585
R636 B.n498 B.n53 585
R637 B.n500 B.n499 585
R638 B.n501 B.n52 585
R639 B.n503 B.n502 585
R640 B.n504 B.n51 585
R641 B.n506 B.n505 585
R642 B.n507 B.n50 585
R643 B.n509 B.n508 585
R644 B.n510 B.n49 585
R645 B.n512 B.n511 585
R646 B.n514 B.n46 585
R647 B.n516 B.n515 585
R648 B.n517 B.n45 585
R649 B.n519 B.n518 585
R650 B.n520 B.n44 585
R651 B.n522 B.n521 585
R652 B.n523 B.n43 585
R653 B.n525 B.n524 585
R654 B.n526 B.n39 585
R655 B.n528 B.n527 585
R656 B.n529 B.n38 585
R657 B.n531 B.n530 585
R658 B.n532 B.n37 585
R659 B.n534 B.n533 585
R660 B.n535 B.n36 585
R661 B.n537 B.n536 585
R662 B.n538 B.n35 585
R663 B.n540 B.n539 585
R664 B.n541 B.n34 585
R665 B.n543 B.n542 585
R666 B.n544 B.n33 585
R667 B.n546 B.n545 585
R668 B.n547 B.n32 585
R669 B.n549 B.n548 585
R670 B.n550 B.n31 585
R671 B.n552 B.n551 585
R672 B.n553 B.n30 585
R673 B.n555 B.n554 585
R674 B.n556 B.n29 585
R675 B.n558 B.n557 585
R676 B.n559 B.n28 585
R677 B.n480 B.n59 585
R678 B.n479 B.n478 585
R679 B.n477 B.n60 585
R680 B.n476 B.n475 585
R681 B.n474 B.n61 585
R682 B.n473 B.n472 585
R683 B.n471 B.n62 585
R684 B.n470 B.n469 585
R685 B.n468 B.n63 585
R686 B.n467 B.n466 585
R687 B.n465 B.n64 585
R688 B.n464 B.n463 585
R689 B.n462 B.n65 585
R690 B.n461 B.n460 585
R691 B.n459 B.n66 585
R692 B.n458 B.n457 585
R693 B.n456 B.n67 585
R694 B.n455 B.n454 585
R695 B.n453 B.n68 585
R696 B.n452 B.n451 585
R697 B.n450 B.n69 585
R698 B.n449 B.n448 585
R699 B.n447 B.n70 585
R700 B.n446 B.n445 585
R701 B.n444 B.n71 585
R702 B.n443 B.n442 585
R703 B.n441 B.n72 585
R704 B.n440 B.n439 585
R705 B.n438 B.n73 585
R706 B.n437 B.n436 585
R707 B.n435 B.n74 585
R708 B.n434 B.n433 585
R709 B.n432 B.n75 585
R710 B.n431 B.n430 585
R711 B.n429 B.n76 585
R712 B.n428 B.n427 585
R713 B.n426 B.n77 585
R714 B.n425 B.n424 585
R715 B.n423 B.n78 585
R716 B.n422 B.n421 585
R717 B.n420 B.n79 585
R718 B.n419 B.n418 585
R719 B.n417 B.n80 585
R720 B.n416 B.n415 585
R721 B.n414 B.n81 585
R722 B.n413 B.n412 585
R723 B.n411 B.n82 585
R724 B.n410 B.n409 585
R725 B.n408 B.n83 585
R726 B.n407 B.n406 585
R727 B.n405 B.n84 585
R728 B.n404 B.n403 585
R729 B.n402 B.n85 585
R730 B.n401 B.n400 585
R731 B.n399 B.n86 585
R732 B.n398 B.n397 585
R733 B.n396 B.n87 585
R734 B.n395 B.n394 585
R735 B.n393 B.n88 585
R736 B.n392 B.n391 585
R737 B.n390 B.n89 585
R738 B.n389 B.n388 585
R739 B.n387 B.n90 585
R740 B.n386 B.n385 585
R741 B.n384 B.n91 585
R742 B.n383 B.n382 585
R743 B.n381 B.n92 585
R744 B.n380 B.n379 585
R745 B.n378 B.n93 585
R746 B.n377 B.n376 585
R747 B.n375 B.n94 585
R748 B.n374 B.n373 585
R749 B.n372 B.n95 585
R750 B.n371 B.n370 585
R751 B.n369 B.n96 585
R752 B.n368 B.n367 585
R753 B.n366 B.n97 585
R754 B.n365 B.n364 585
R755 B.n363 B.n98 585
R756 B.n362 B.n361 585
R757 B.n360 B.n99 585
R758 B.n359 B.n358 585
R759 B.n357 B.n100 585
R760 B.n356 B.n355 585
R761 B.n354 B.n101 585
R762 B.n353 B.n352 585
R763 B.n351 B.n102 585
R764 B.n350 B.n349 585
R765 B.n348 B.n103 585
R766 B.n347 B.n346 585
R767 B.n345 B.n104 585
R768 B.n344 B.n343 585
R769 B.n342 B.n105 585
R770 B.n341 B.n340 585
R771 B.n339 B.n106 585
R772 B.n338 B.n337 585
R773 B.n336 B.n107 585
R774 B.n335 B.n334 585
R775 B.n333 B.n108 585
R776 B.n332 B.n331 585
R777 B.n330 B.n109 585
R778 B.n329 B.n328 585
R779 B.n327 B.n110 585
R780 B.n326 B.n325 585
R781 B.n324 B.n111 585
R782 B.n245 B.n244 585
R783 B.n246 B.n141 585
R784 B.n248 B.n247 585
R785 B.n249 B.n140 585
R786 B.n251 B.n250 585
R787 B.n252 B.n139 585
R788 B.n254 B.n253 585
R789 B.n255 B.n138 585
R790 B.n257 B.n256 585
R791 B.n258 B.n137 585
R792 B.n260 B.n259 585
R793 B.n261 B.n136 585
R794 B.n263 B.n262 585
R795 B.n264 B.n135 585
R796 B.n266 B.n265 585
R797 B.n267 B.n134 585
R798 B.n269 B.n268 585
R799 B.n270 B.n133 585
R800 B.n272 B.n271 585
R801 B.n273 B.n132 585
R802 B.n275 B.n274 585
R803 B.n277 B.n276 585
R804 B.n278 B.n128 585
R805 B.n280 B.n279 585
R806 B.n281 B.n127 585
R807 B.n283 B.n282 585
R808 B.n284 B.n126 585
R809 B.n286 B.n285 585
R810 B.n287 B.n125 585
R811 B.n289 B.n288 585
R812 B.n290 B.n122 585
R813 B.n293 B.n292 585
R814 B.n294 B.n121 585
R815 B.n296 B.n295 585
R816 B.n297 B.n120 585
R817 B.n299 B.n298 585
R818 B.n300 B.n119 585
R819 B.n302 B.n301 585
R820 B.n303 B.n118 585
R821 B.n305 B.n304 585
R822 B.n306 B.n117 585
R823 B.n308 B.n307 585
R824 B.n309 B.n116 585
R825 B.n311 B.n310 585
R826 B.n312 B.n115 585
R827 B.n314 B.n313 585
R828 B.n315 B.n114 585
R829 B.n317 B.n316 585
R830 B.n318 B.n113 585
R831 B.n320 B.n319 585
R832 B.n321 B.n112 585
R833 B.n323 B.n322 585
R834 B.n243 B.n142 585
R835 B.n242 B.n241 585
R836 B.n240 B.n143 585
R837 B.n239 B.n238 585
R838 B.n237 B.n144 585
R839 B.n236 B.n235 585
R840 B.n234 B.n145 585
R841 B.n233 B.n232 585
R842 B.n231 B.n146 585
R843 B.n230 B.n229 585
R844 B.n228 B.n147 585
R845 B.n227 B.n226 585
R846 B.n225 B.n148 585
R847 B.n224 B.n223 585
R848 B.n222 B.n149 585
R849 B.n221 B.n220 585
R850 B.n219 B.n150 585
R851 B.n218 B.n217 585
R852 B.n216 B.n151 585
R853 B.n215 B.n214 585
R854 B.n213 B.n152 585
R855 B.n212 B.n211 585
R856 B.n210 B.n153 585
R857 B.n209 B.n208 585
R858 B.n207 B.n154 585
R859 B.n206 B.n205 585
R860 B.n204 B.n155 585
R861 B.n203 B.n202 585
R862 B.n201 B.n156 585
R863 B.n200 B.n199 585
R864 B.n198 B.n157 585
R865 B.n197 B.n196 585
R866 B.n195 B.n158 585
R867 B.n194 B.n193 585
R868 B.n192 B.n159 585
R869 B.n191 B.n190 585
R870 B.n189 B.n160 585
R871 B.n188 B.n187 585
R872 B.n186 B.n161 585
R873 B.n185 B.n184 585
R874 B.n183 B.n162 585
R875 B.n182 B.n181 585
R876 B.n180 B.n163 585
R877 B.n179 B.n178 585
R878 B.n177 B.n164 585
R879 B.n176 B.n175 585
R880 B.n174 B.n165 585
R881 B.n173 B.n172 585
R882 B.n171 B.n166 585
R883 B.n170 B.n169 585
R884 B.n168 B.n167 585
R885 B.n2 B.n0 585
R886 B.n637 B.n1 585
R887 B.n636 B.n635 585
R888 B.n634 B.n3 585
R889 B.n633 B.n632 585
R890 B.n631 B.n4 585
R891 B.n630 B.n629 585
R892 B.n628 B.n5 585
R893 B.n627 B.n626 585
R894 B.n625 B.n6 585
R895 B.n624 B.n623 585
R896 B.n622 B.n7 585
R897 B.n621 B.n620 585
R898 B.n619 B.n8 585
R899 B.n618 B.n617 585
R900 B.n616 B.n9 585
R901 B.n615 B.n614 585
R902 B.n613 B.n10 585
R903 B.n612 B.n611 585
R904 B.n610 B.n11 585
R905 B.n609 B.n608 585
R906 B.n607 B.n12 585
R907 B.n606 B.n605 585
R908 B.n604 B.n13 585
R909 B.n603 B.n602 585
R910 B.n601 B.n14 585
R911 B.n600 B.n599 585
R912 B.n598 B.n15 585
R913 B.n597 B.n596 585
R914 B.n595 B.n16 585
R915 B.n594 B.n593 585
R916 B.n592 B.n17 585
R917 B.n591 B.n590 585
R918 B.n589 B.n18 585
R919 B.n588 B.n587 585
R920 B.n586 B.n19 585
R921 B.n585 B.n584 585
R922 B.n583 B.n20 585
R923 B.n582 B.n581 585
R924 B.n580 B.n21 585
R925 B.n579 B.n578 585
R926 B.n577 B.n22 585
R927 B.n576 B.n575 585
R928 B.n574 B.n23 585
R929 B.n573 B.n572 585
R930 B.n571 B.n24 585
R931 B.n570 B.n569 585
R932 B.n568 B.n25 585
R933 B.n567 B.n566 585
R934 B.n565 B.n26 585
R935 B.n564 B.n563 585
R936 B.n562 B.n27 585
R937 B.n561 B.n560 585
R938 B.n639 B.n638 585
R939 B.n245 B.n142 535.745
R940 B.n560 B.n559 535.745
R941 B.n324 B.n323 535.745
R942 B.n481 B.n480 535.745
R943 B.n123 B.t11 300.837
R944 B.n47 B.t1 300.837
R945 B.n129 B.t5 300.837
R946 B.n40 B.t7 300.837
R947 B.n123 B.t9 264.397
R948 B.n129 B.t3 264.397
R949 B.n40 B.t6 264.397
R950 B.n47 B.t0 264.397
R951 B.n124 B.t10 252.546
R952 B.n48 B.t2 252.546
R953 B.n130 B.t4 252.546
R954 B.n41 B.t8 252.546
R955 B.n241 B.n142 163.367
R956 B.n241 B.n240 163.367
R957 B.n240 B.n239 163.367
R958 B.n239 B.n144 163.367
R959 B.n235 B.n144 163.367
R960 B.n235 B.n234 163.367
R961 B.n234 B.n233 163.367
R962 B.n233 B.n146 163.367
R963 B.n229 B.n146 163.367
R964 B.n229 B.n228 163.367
R965 B.n228 B.n227 163.367
R966 B.n227 B.n148 163.367
R967 B.n223 B.n148 163.367
R968 B.n223 B.n222 163.367
R969 B.n222 B.n221 163.367
R970 B.n221 B.n150 163.367
R971 B.n217 B.n150 163.367
R972 B.n217 B.n216 163.367
R973 B.n216 B.n215 163.367
R974 B.n215 B.n152 163.367
R975 B.n211 B.n152 163.367
R976 B.n211 B.n210 163.367
R977 B.n210 B.n209 163.367
R978 B.n209 B.n154 163.367
R979 B.n205 B.n154 163.367
R980 B.n205 B.n204 163.367
R981 B.n204 B.n203 163.367
R982 B.n203 B.n156 163.367
R983 B.n199 B.n156 163.367
R984 B.n199 B.n198 163.367
R985 B.n198 B.n197 163.367
R986 B.n197 B.n158 163.367
R987 B.n193 B.n158 163.367
R988 B.n193 B.n192 163.367
R989 B.n192 B.n191 163.367
R990 B.n191 B.n160 163.367
R991 B.n187 B.n160 163.367
R992 B.n187 B.n186 163.367
R993 B.n186 B.n185 163.367
R994 B.n185 B.n162 163.367
R995 B.n181 B.n162 163.367
R996 B.n181 B.n180 163.367
R997 B.n180 B.n179 163.367
R998 B.n179 B.n164 163.367
R999 B.n175 B.n164 163.367
R1000 B.n175 B.n174 163.367
R1001 B.n174 B.n173 163.367
R1002 B.n173 B.n166 163.367
R1003 B.n169 B.n166 163.367
R1004 B.n169 B.n168 163.367
R1005 B.n168 B.n2 163.367
R1006 B.n638 B.n2 163.367
R1007 B.n638 B.n637 163.367
R1008 B.n637 B.n636 163.367
R1009 B.n636 B.n3 163.367
R1010 B.n632 B.n3 163.367
R1011 B.n632 B.n631 163.367
R1012 B.n631 B.n630 163.367
R1013 B.n630 B.n5 163.367
R1014 B.n626 B.n5 163.367
R1015 B.n626 B.n625 163.367
R1016 B.n625 B.n624 163.367
R1017 B.n624 B.n7 163.367
R1018 B.n620 B.n7 163.367
R1019 B.n620 B.n619 163.367
R1020 B.n619 B.n618 163.367
R1021 B.n618 B.n9 163.367
R1022 B.n614 B.n9 163.367
R1023 B.n614 B.n613 163.367
R1024 B.n613 B.n612 163.367
R1025 B.n612 B.n11 163.367
R1026 B.n608 B.n11 163.367
R1027 B.n608 B.n607 163.367
R1028 B.n607 B.n606 163.367
R1029 B.n606 B.n13 163.367
R1030 B.n602 B.n13 163.367
R1031 B.n602 B.n601 163.367
R1032 B.n601 B.n600 163.367
R1033 B.n600 B.n15 163.367
R1034 B.n596 B.n15 163.367
R1035 B.n596 B.n595 163.367
R1036 B.n595 B.n594 163.367
R1037 B.n594 B.n17 163.367
R1038 B.n590 B.n17 163.367
R1039 B.n590 B.n589 163.367
R1040 B.n589 B.n588 163.367
R1041 B.n588 B.n19 163.367
R1042 B.n584 B.n19 163.367
R1043 B.n584 B.n583 163.367
R1044 B.n583 B.n582 163.367
R1045 B.n582 B.n21 163.367
R1046 B.n578 B.n21 163.367
R1047 B.n578 B.n577 163.367
R1048 B.n577 B.n576 163.367
R1049 B.n576 B.n23 163.367
R1050 B.n572 B.n23 163.367
R1051 B.n572 B.n571 163.367
R1052 B.n571 B.n570 163.367
R1053 B.n570 B.n25 163.367
R1054 B.n566 B.n25 163.367
R1055 B.n566 B.n565 163.367
R1056 B.n565 B.n564 163.367
R1057 B.n564 B.n27 163.367
R1058 B.n560 B.n27 163.367
R1059 B.n246 B.n245 163.367
R1060 B.n247 B.n246 163.367
R1061 B.n247 B.n140 163.367
R1062 B.n251 B.n140 163.367
R1063 B.n252 B.n251 163.367
R1064 B.n253 B.n252 163.367
R1065 B.n253 B.n138 163.367
R1066 B.n257 B.n138 163.367
R1067 B.n258 B.n257 163.367
R1068 B.n259 B.n258 163.367
R1069 B.n259 B.n136 163.367
R1070 B.n263 B.n136 163.367
R1071 B.n264 B.n263 163.367
R1072 B.n265 B.n264 163.367
R1073 B.n265 B.n134 163.367
R1074 B.n269 B.n134 163.367
R1075 B.n270 B.n269 163.367
R1076 B.n271 B.n270 163.367
R1077 B.n271 B.n132 163.367
R1078 B.n275 B.n132 163.367
R1079 B.n276 B.n275 163.367
R1080 B.n276 B.n128 163.367
R1081 B.n280 B.n128 163.367
R1082 B.n281 B.n280 163.367
R1083 B.n282 B.n281 163.367
R1084 B.n282 B.n126 163.367
R1085 B.n286 B.n126 163.367
R1086 B.n287 B.n286 163.367
R1087 B.n288 B.n287 163.367
R1088 B.n288 B.n122 163.367
R1089 B.n293 B.n122 163.367
R1090 B.n294 B.n293 163.367
R1091 B.n295 B.n294 163.367
R1092 B.n295 B.n120 163.367
R1093 B.n299 B.n120 163.367
R1094 B.n300 B.n299 163.367
R1095 B.n301 B.n300 163.367
R1096 B.n301 B.n118 163.367
R1097 B.n305 B.n118 163.367
R1098 B.n306 B.n305 163.367
R1099 B.n307 B.n306 163.367
R1100 B.n307 B.n116 163.367
R1101 B.n311 B.n116 163.367
R1102 B.n312 B.n311 163.367
R1103 B.n313 B.n312 163.367
R1104 B.n313 B.n114 163.367
R1105 B.n317 B.n114 163.367
R1106 B.n318 B.n317 163.367
R1107 B.n319 B.n318 163.367
R1108 B.n319 B.n112 163.367
R1109 B.n323 B.n112 163.367
R1110 B.n325 B.n324 163.367
R1111 B.n325 B.n110 163.367
R1112 B.n329 B.n110 163.367
R1113 B.n330 B.n329 163.367
R1114 B.n331 B.n330 163.367
R1115 B.n331 B.n108 163.367
R1116 B.n335 B.n108 163.367
R1117 B.n336 B.n335 163.367
R1118 B.n337 B.n336 163.367
R1119 B.n337 B.n106 163.367
R1120 B.n341 B.n106 163.367
R1121 B.n342 B.n341 163.367
R1122 B.n343 B.n342 163.367
R1123 B.n343 B.n104 163.367
R1124 B.n347 B.n104 163.367
R1125 B.n348 B.n347 163.367
R1126 B.n349 B.n348 163.367
R1127 B.n349 B.n102 163.367
R1128 B.n353 B.n102 163.367
R1129 B.n354 B.n353 163.367
R1130 B.n355 B.n354 163.367
R1131 B.n355 B.n100 163.367
R1132 B.n359 B.n100 163.367
R1133 B.n360 B.n359 163.367
R1134 B.n361 B.n360 163.367
R1135 B.n361 B.n98 163.367
R1136 B.n365 B.n98 163.367
R1137 B.n366 B.n365 163.367
R1138 B.n367 B.n366 163.367
R1139 B.n367 B.n96 163.367
R1140 B.n371 B.n96 163.367
R1141 B.n372 B.n371 163.367
R1142 B.n373 B.n372 163.367
R1143 B.n373 B.n94 163.367
R1144 B.n377 B.n94 163.367
R1145 B.n378 B.n377 163.367
R1146 B.n379 B.n378 163.367
R1147 B.n379 B.n92 163.367
R1148 B.n383 B.n92 163.367
R1149 B.n384 B.n383 163.367
R1150 B.n385 B.n384 163.367
R1151 B.n385 B.n90 163.367
R1152 B.n389 B.n90 163.367
R1153 B.n390 B.n389 163.367
R1154 B.n391 B.n390 163.367
R1155 B.n391 B.n88 163.367
R1156 B.n395 B.n88 163.367
R1157 B.n396 B.n395 163.367
R1158 B.n397 B.n396 163.367
R1159 B.n397 B.n86 163.367
R1160 B.n401 B.n86 163.367
R1161 B.n402 B.n401 163.367
R1162 B.n403 B.n402 163.367
R1163 B.n403 B.n84 163.367
R1164 B.n407 B.n84 163.367
R1165 B.n408 B.n407 163.367
R1166 B.n409 B.n408 163.367
R1167 B.n409 B.n82 163.367
R1168 B.n413 B.n82 163.367
R1169 B.n414 B.n413 163.367
R1170 B.n415 B.n414 163.367
R1171 B.n415 B.n80 163.367
R1172 B.n419 B.n80 163.367
R1173 B.n420 B.n419 163.367
R1174 B.n421 B.n420 163.367
R1175 B.n421 B.n78 163.367
R1176 B.n425 B.n78 163.367
R1177 B.n426 B.n425 163.367
R1178 B.n427 B.n426 163.367
R1179 B.n427 B.n76 163.367
R1180 B.n431 B.n76 163.367
R1181 B.n432 B.n431 163.367
R1182 B.n433 B.n432 163.367
R1183 B.n433 B.n74 163.367
R1184 B.n437 B.n74 163.367
R1185 B.n438 B.n437 163.367
R1186 B.n439 B.n438 163.367
R1187 B.n439 B.n72 163.367
R1188 B.n443 B.n72 163.367
R1189 B.n444 B.n443 163.367
R1190 B.n445 B.n444 163.367
R1191 B.n445 B.n70 163.367
R1192 B.n449 B.n70 163.367
R1193 B.n450 B.n449 163.367
R1194 B.n451 B.n450 163.367
R1195 B.n451 B.n68 163.367
R1196 B.n455 B.n68 163.367
R1197 B.n456 B.n455 163.367
R1198 B.n457 B.n456 163.367
R1199 B.n457 B.n66 163.367
R1200 B.n461 B.n66 163.367
R1201 B.n462 B.n461 163.367
R1202 B.n463 B.n462 163.367
R1203 B.n463 B.n64 163.367
R1204 B.n467 B.n64 163.367
R1205 B.n468 B.n467 163.367
R1206 B.n469 B.n468 163.367
R1207 B.n469 B.n62 163.367
R1208 B.n473 B.n62 163.367
R1209 B.n474 B.n473 163.367
R1210 B.n475 B.n474 163.367
R1211 B.n475 B.n60 163.367
R1212 B.n479 B.n60 163.367
R1213 B.n480 B.n479 163.367
R1214 B.n559 B.n558 163.367
R1215 B.n558 B.n29 163.367
R1216 B.n554 B.n29 163.367
R1217 B.n554 B.n553 163.367
R1218 B.n553 B.n552 163.367
R1219 B.n552 B.n31 163.367
R1220 B.n548 B.n31 163.367
R1221 B.n548 B.n547 163.367
R1222 B.n547 B.n546 163.367
R1223 B.n546 B.n33 163.367
R1224 B.n542 B.n33 163.367
R1225 B.n542 B.n541 163.367
R1226 B.n541 B.n540 163.367
R1227 B.n540 B.n35 163.367
R1228 B.n536 B.n35 163.367
R1229 B.n536 B.n535 163.367
R1230 B.n535 B.n534 163.367
R1231 B.n534 B.n37 163.367
R1232 B.n530 B.n37 163.367
R1233 B.n530 B.n529 163.367
R1234 B.n529 B.n528 163.367
R1235 B.n528 B.n39 163.367
R1236 B.n524 B.n39 163.367
R1237 B.n524 B.n523 163.367
R1238 B.n523 B.n522 163.367
R1239 B.n522 B.n44 163.367
R1240 B.n518 B.n44 163.367
R1241 B.n518 B.n517 163.367
R1242 B.n517 B.n516 163.367
R1243 B.n516 B.n46 163.367
R1244 B.n511 B.n46 163.367
R1245 B.n511 B.n510 163.367
R1246 B.n510 B.n509 163.367
R1247 B.n509 B.n50 163.367
R1248 B.n505 B.n50 163.367
R1249 B.n505 B.n504 163.367
R1250 B.n504 B.n503 163.367
R1251 B.n503 B.n52 163.367
R1252 B.n499 B.n52 163.367
R1253 B.n499 B.n498 163.367
R1254 B.n498 B.n497 163.367
R1255 B.n497 B.n54 163.367
R1256 B.n493 B.n54 163.367
R1257 B.n493 B.n492 163.367
R1258 B.n492 B.n491 163.367
R1259 B.n491 B.n56 163.367
R1260 B.n487 B.n56 163.367
R1261 B.n487 B.n486 163.367
R1262 B.n486 B.n485 163.367
R1263 B.n485 B.n58 163.367
R1264 B.n481 B.n58 163.367
R1265 B.n291 B.n124 59.5399
R1266 B.n131 B.n130 59.5399
R1267 B.n42 B.n41 59.5399
R1268 B.n513 B.n48 59.5399
R1269 B.n124 B.n123 48.2914
R1270 B.n130 B.n129 48.2914
R1271 B.n41 B.n40 48.2914
R1272 B.n48 B.n47 48.2914
R1273 B.n561 B.n28 34.8103
R1274 B.n482 B.n59 34.8103
R1275 B.n322 B.n111 34.8103
R1276 B.n244 B.n243 34.8103
R1277 B B.n639 18.0485
R1278 B.n557 B.n28 10.6151
R1279 B.n557 B.n556 10.6151
R1280 B.n556 B.n555 10.6151
R1281 B.n555 B.n30 10.6151
R1282 B.n551 B.n30 10.6151
R1283 B.n551 B.n550 10.6151
R1284 B.n550 B.n549 10.6151
R1285 B.n549 B.n32 10.6151
R1286 B.n545 B.n32 10.6151
R1287 B.n545 B.n544 10.6151
R1288 B.n544 B.n543 10.6151
R1289 B.n543 B.n34 10.6151
R1290 B.n539 B.n34 10.6151
R1291 B.n539 B.n538 10.6151
R1292 B.n538 B.n537 10.6151
R1293 B.n537 B.n36 10.6151
R1294 B.n533 B.n36 10.6151
R1295 B.n533 B.n532 10.6151
R1296 B.n532 B.n531 10.6151
R1297 B.n531 B.n38 10.6151
R1298 B.n527 B.n526 10.6151
R1299 B.n526 B.n525 10.6151
R1300 B.n525 B.n43 10.6151
R1301 B.n521 B.n43 10.6151
R1302 B.n521 B.n520 10.6151
R1303 B.n520 B.n519 10.6151
R1304 B.n519 B.n45 10.6151
R1305 B.n515 B.n45 10.6151
R1306 B.n515 B.n514 10.6151
R1307 B.n512 B.n49 10.6151
R1308 B.n508 B.n49 10.6151
R1309 B.n508 B.n507 10.6151
R1310 B.n507 B.n506 10.6151
R1311 B.n506 B.n51 10.6151
R1312 B.n502 B.n51 10.6151
R1313 B.n502 B.n501 10.6151
R1314 B.n501 B.n500 10.6151
R1315 B.n500 B.n53 10.6151
R1316 B.n496 B.n53 10.6151
R1317 B.n496 B.n495 10.6151
R1318 B.n495 B.n494 10.6151
R1319 B.n494 B.n55 10.6151
R1320 B.n490 B.n55 10.6151
R1321 B.n490 B.n489 10.6151
R1322 B.n489 B.n488 10.6151
R1323 B.n488 B.n57 10.6151
R1324 B.n484 B.n57 10.6151
R1325 B.n484 B.n483 10.6151
R1326 B.n483 B.n482 10.6151
R1327 B.n326 B.n111 10.6151
R1328 B.n327 B.n326 10.6151
R1329 B.n328 B.n327 10.6151
R1330 B.n328 B.n109 10.6151
R1331 B.n332 B.n109 10.6151
R1332 B.n333 B.n332 10.6151
R1333 B.n334 B.n333 10.6151
R1334 B.n334 B.n107 10.6151
R1335 B.n338 B.n107 10.6151
R1336 B.n339 B.n338 10.6151
R1337 B.n340 B.n339 10.6151
R1338 B.n340 B.n105 10.6151
R1339 B.n344 B.n105 10.6151
R1340 B.n345 B.n344 10.6151
R1341 B.n346 B.n345 10.6151
R1342 B.n346 B.n103 10.6151
R1343 B.n350 B.n103 10.6151
R1344 B.n351 B.n350 10.6151
R1345 B.n352 B.n351 10.6151
R1346 B.n352 B.n101 10.6151
R1347 B.n356 B.n101 10.6151
R1348 B.n357 B.n356 10.6151
R1349 B.n358 B.n357 10.6151
R1350 B.n358 B.n99 10.6151
R1351 B.n362 B.n99 10.6151
R1352 B.n363 B.n362 10.6151
R1353 B.n364 B.n363 10.6151
R1354 B.n364 B.n97 10.6151
R1355 B.n368 B.n97 10.6151
R1356 B.n369 B.n368 10.6151
R1357 B.n370 B.n369 10.6151
R1358 B.n370 B.n95 10.6151
R1359 B.n374 B.n95 10.6151
R1360 B.n375 B.n374 10.6151
R1361 B.n376 B.n375 10.6151
R1362 B.n376 B.n93 10.6151
R1363 B.n380 B.n93 10.6151
R1364 B.n381 B.n380 10.6151
R1365 B.n382 B.n381 10.6151
R1366 B.n382 B.n91 10.6151
R1367 B.n386 B.n91 10.6151
R1368 B.n387 B.n386 10.6151
R1369 B.n388 B.n387 10.6151
R1370 B.n388 B.n89 10.6151
R1371 B.n392 B.n89 10.6151
R1372 B.n393 B.n392 10.6151
R1373 B.n394 B.n393 10.6151
R1374 B.n394 B.n87 10.6151
R1375 B.n398 B.n87 10.6151
R1376 B.n399 B.n398 10.6151
R1377 B.n400 B.n399 10.6151
R1378 B.n400 B.n85 10.6151
R1379 B.n404 B.n85 10.6151
R1380 B.n405 B.n404 10.6151
R1381 B.n406 B.n405 10.6151
R1382 B.n406 B.n83 10.6151
R1383 B.n410 B.n83 10.6151
R1384 B.n411 B.n410 10.6151
R1385 B.n412 B.n411 10.6151
R1386 B.n412 B.n81 10.6151
R1387 B.n416 B.n81 10.6151
R1388 B.n417 B.n416 10.6151
R1389 B.n418 B.n417 10.6151
R1390 B.n418 B.n79 10.6151
R1391 B.n422 B.n79 10.6151
R1392 B.n423 B.n422 10.6151
R1393 B.n424 B.n423 10.6151
R1394 B.n424 B.n77 10.6151
R1395 B.n428 B.n77 10.6151
R1396 B.n429 B.n428 10.6151
R1397 B.n430 B.n429 10.6151
R1398 B.n430 B.n75 10.6151
R1399 B.n434 B.n75 10.6151
R1400 B.n435 B.n434 10.6151
R1401 B.n436 B.n435 10.6151
R1402 B.n436 B.n73 10.6151
R1403 B.n440 B.n73 10.6151
R1404 B.n441 B.n440 10.6151
R1405 B.n442 B.n441 10.6151
R1406 B.n442 B.n71 10.6151
R1407 B.n446 B.n71 10.6151
R1408 B.n447 B.n446 10.6151
R1409 B.n448 B.n447 10.6151
R1410 B.n448 B.n69 10.6151
R1411 B.n452 B.n69 10.6151
R1412 B.n453 B.n452 10.6151
R1413 B.n454 B.n453 10.6151
R1414 B.n454 B.n67 10.6151
R1415 B.n458 B.n67 10.6151
R1416 B.n459 B.n458 10.6151
R1417 B.n460 B.n459 10.6151
R1418 B.n460 B.n65 10.6151
R1419 B.n464 B.n65 10.6151
R1420 B.n465 B.n464 10.6151
R1421 B.n466 B.n465 10.6151
R1422 B.n466 B.n63 10.6151
R1423 B.n470 B.n63 10.6151
R1424 B.n471 B.n470 10.6151
R1425 B.n472 B.n471 10.6151
R1426 B.n472 B.n61 10.6151
R1427 B.n476 B.n61 10.6151
R1428 B.n477 B.n476 10.6151
R1429 B.n478 B.n477 10.6151
R1430 B.n478 B.n59 10.6151
R1431 B.n244 B.n141 10.6151
R1432 B.n248 B.n141 10.6151
R1433 B.n249 B.n248 10.6151
R1434 B.n250 B.n249 10.6151
R1435 B.n250 B.n139 10.6151
R1436 B.n254 B.n139 10.6151
R1437 B.n255 B.n254 10.6151
R1438 B.n256 B.n255 10.6151
R1439 B.n256 B.n137 10.6151
R1440 B.n260 B.n137 10.6151
R1441 B.n261 B.n260 10.6151
R1442 B.n262 B.n261 10.6151
R1443 B.n262 B.n135 10.6151
R1444 B.n266 B.n135 10.6151
R1445 B.n267 B.n266 10.6151
R1446 B.n268 B.n267 10.6151
R1447 B.n268 B.n133 10.6151
R1448 B.n272 B.n133 10.6151
R1449 B.n273 B.n272 10.6151
R1450 B.n274 B.n273 10.6151
R1451 B.n278 B.n277 10.6151
R1452 B.n279 B.n278 10.6151
R1453 B.n279 B.n127 10.6151
R1454 B.n283 B.n127 10.6151
R1455 B.n284 B.n283 10.6151
R1456 B.n285 B.n284 10.6151
R1457 B.n285 B.n125 10.6151
R1458 B.n289 B.n125 10.6151
R1459 B.n290 B.n289 10.6151
R1460 B.n292 B.n121 10.6151
R1461 B.n296 B.n121 10.6151
R1462 B.n297 B.n296 10.6151
R1463 B.n298 B.n297 10.6151
R1464 B.n298 B.n119 10.6151
R1465 B.n302 B.n119 10.6151
R1466 B.n303 B.n302 10.6151
R1467 B.n304 B.n303 10.6151
R1468 B.n304 B.n117 10.6151
R1469 B.n308 B.n117 10.6151
R1470 B.n309 B.n308 10.6151
R1471 B.n310 B.n309 10.6151
R1472 B.n310 B.n115 10.6151
R1473 B.n314 B.n115 10.6151
R1474 B.n315 B.n314 10.6151
R1475 B.n316 B.n315 10.6151
R1476 B.n316 B.n113 10.6151
R1477 B.n320 B.n113 10.6151
R1478 B.n321 B.n320 10.6151
R1479 B.n322 B.n321 10.6151
R1480 B.n243 B.n242 10.6151
R1481 B.n242 B.n143 10.6151
R1482 B.n238 B.n143 10.6151
R1483 B.n238 B.n237 10.6151
R1484 B.n237 B.n236 10.6151
R1485 B.n236 B.n145 10.6151
R1486 B.n232 B.n145 10.6151
R1487 B.n232 B.n231 10.6151
R1488 B.n231 B.n230 10.6151
R1489 B.n230 B.n147 10.6151
R1490 B.n226 B.n147 10.6151
R1491 B.n226 B.n225 10.6151
R1492 B.n225 B.n224 10.6151
R1493 B.n224 B.n149 10.6151
R1494 B.n220 B.n149 10.6151
R1495 B.n220 B.n219 10.6151
R1496 B.n219 B.n218 10.6151
R1497 B.n218 B.n151 10.6151
R1498 B.n214 B.n151 10.6151
R1499 B.n214 B.n213 10.6151
R1500 B.n213 B.n212 10.6151
R1501 B.n212 B.n153 10.6151
R1502 B.n208 B.n153 10.6151
R1503 B.n208 B.n207 10.6151
R1504 B.n207 B.n206 10.6151
R1505 B.n206 B.n155 10.6151
R1506 B.n202 B.n155 10.6151
R1507 B.n202 B.n201 10.6151
R1508 B.n201 B.n200 10.6151
R1509 B.n200 B.n157 10.6151
R1510 B.n196 B.n157 10.6151
R1511 B.n196 B.n195 10.6151
R1512 B.n195 B.n194 10.6151
R1513 B.n194 B.n159 10.6151
R1514 B.n190 B.n159 10.6151
R1515 B.n190 B.n189 10.6151
R1516 B.n189 B.n188 10.6151
R1517 B.n188 B.n161 10.6151
R1518 B.n184 B.n161 10.6151
R1519 B.n184 B.n183 10.6151
R1520 B.n183 B.n182 10.6151
R1521 B.n182 B.n163 10.6151
R1522 B.n178 B.n163 10.6151
R1523 B.n178 B.n177 10.6151
R1524 B.n177 B.n176 10.6151
R1525 B.n176 B.n165 10.6151
R1526 B.n172 B.n165 10.6151
R1527 B.n172 B.n171 10.6151
R1528 B.n171 B.n170 10.6151
R1529 B.n170 B.n167 10.6151
R1530 B.n167 B.n0 10.6151
R1531 B.n635 B.n1 10.6151
R1532 B.n635 B.n634 10.6151
R1533 B.n634 B.n633 10.6151
R1534 B.n633 B.n4 10.6151
R1535 B.n629 B.n4 10.6151
R1536 B.n629 B.n628 10.6151
R1537 B.n628 B.n627 10.6151
R1538 B.n627 B.n6 10.6151
R1539 B.n623 B.n6 10.6151
R1540 B.n623 B.n622 10.6151
R1541 B.n622 B.n621 10.6151
R1542 B.n621 B.n8 10.6151
R1543 B.n617 B.n8 10.6151
R1544 B.n617 B.n616 10.6151
R1545 B.n616 B.n615 10.6151
R1546 B.n615 B.n10 10.6151
R1547 B.n611 B.n10 10.6151
R1548 B.n611 B.n610 10.6151
R1549 B.n610 B.n609 10.6151
R1550 B.n609 B.n12 10.6151
R1551 B.n605 B.n12 10.6151
R1552 B.n605 B.n604 10.6151
R1553 B.n604 B.n603 10.6151
R1554 B.n603 B.n14 10.6151
R1555 B.n599 B.n14 10.6151
R1556 B.n599 B.n598 10.6151
R1557 B.n598 B.n597 10.6151
R1558 B.n597 B.n16 10.6151
R1559 B.n593 B.n16 10.6151
R1560 B.n593 B.n592 10.6151
R1561 B.n592 B.n591 10.6151
R1562 B.n591 B.n18 10.6151
R1563 B.n587 B.n18 10.6151
R1564 B.n587 B.n586 10.6151
R1565 B.n586 B.n585 10.6151
R1566 B.n585 B.n20 10.6151
R1567 B.n581 B.n20 10.6151
R1568 B.n581 B.n580 10.6151
R1569 B.n580 B.n579 10.6151
R1570 B.n579 B.n22 10.6151
R1571 B.n575 B.n22 10.6151
R1572 B.n575 B.n574 10.6151
R1573 B.n574 B.n573 10.6151
R1574 B.n573 B.n24 10.6151
R1575 B.n569 B.n24 10.6151
R1576 B.n569 B.n568 10.6151
R1577 B.n568 B.n567 10.6151
R1578 B.n567 B.n26 10.6151
R1579 B.n563 B.n26 10.6151
R1580 B.n563 B.n562 10.6151
R1581 B.n562 B.n561 10.6151
R1582 B.n42 B.n38 9.36635
R1583 B.n513 B.n512 9.36635
R1584 B.n274 B.n131 9.36635
R1585 B.n292 B.n291 9.36635
R1586 B.n639 B.n0 2.81026
R1587 B.n639 B.n1 2.81026
R1588 B.n527 B.n42 1.24928
R1589 B.n514 B.n513 1.24928
R1590 B.n277 B.n131 1.24928
R1591 B.n291 B.n290 1.24928
C0 VDD2 VN 4.6718f
C1 VP VDD2 0.530975f
C2 VTAIL VDD2 6.95349f
C3 B w_n3958_n1992# 7.88783f
C4 VDD1 B 1.77033f
C5 VDD1 w_n3958_n1992# 2.13146f
C6 VP VN 6.47452f
C7 VTAIL VN 5.60928f
C8 VP VTAIL 5.62348f
C9 B VDD2 1.87123f
C10 VDD2 w_n3958_n1992# 2.25196f
C11 VDD1 VDD2 1.88426f
C12 B VN 1.12859f
C13 VN w_n3958_n1992# 8.22544f
C14 VDD1 VN 0.152273f
C15 VP B 1.99036f
C16 B VTAIL 2.03296f
C17 VP w_n3958_n1992# 8.73931f
C18 VTAIL w_n3958_n1992# 2.15402f
C19 VP VDD1 5.04366f
C20 VDD1 VTAIL 6.90413f
C21 VDD2 VSUBS 1.620329f
C22 VDD1 VSUBS 1.553789f
C23 VTAIL VSUBS 0.604824f
C24 VN VSUBS 6.63387f
C25 VP VSUBS 3.16856f
C26 B VSUBS 3.998492f
C27 w_n3958_n1992# VSUBS 98.7442f
C28 B.n0 VSUBS 0.005093f
C29 B.n1 VSUBS 0.005093f
C30 B.n2 VSUBS 0.008053f
C31 B.n3 VSUBS 0.008053f
C32 B.n4 VSUBS 0.008053f
C33 B.n5 VSUBS 0.008053f
C34 B.n6 VSUBS 0.008053f
C35 B.n7 VSUBS 0.008053f
C36 B.n8 VSUBS 0.008053f
C37 B.n9 VSUBS 0.008053f
C38 B.n10 VSUBS 0.008053f
C39 B.n11 VSUBS 0.008053f
C40 B.n12 VSUBS 0.008053f
C41 B.n13 VSUBS 0.008053f
C42 B.n14 VSUBS 0.008053f
C43 B.n15 VSUBS 0.008053f
C44 B.n16 VSUBS 0.008053f
C45 B.n17 VSUBS 0.008053f
C46 B.n18 VSUBS 0.008053f
C47 B.n19 VSUBS 0.008053f
C48 B.n20 VSUBS 0.008053f
C49 B.n21 VSUBS 0.008053f
C50 B.n22 VSUBS 0.008053f
C51 B.n23 VSUBS 0.008053f
C52 B.n24 VSUBS 0.008053f
C53 B.n25 VSUBS 0.008053f
C54 B.n26 VSUBS 0.008053f
C55 B.n27 VSUBS 0.008053f
C56 B.n28 VSUBS 0.019997f
C57 B.n29 VSUBS 0.008053f
C58 B.n30 VSUBS 0.008053f
C59 B.n31 VSUBS 0.008053f
C60 B.n32 VSUBS 0.008053f
C61 B.n33 VSUBS 0.008053f
C62 B.n34 VSUBS 0.008053f
C63 B.n35 VSUBS 0.008053f
C64 B.n36 VSUBS 0.008053f
C65 B.n37 VSUBS 0.008053f
C66 B.n38 VSUBS 0.00758f
C67 B.n39 VSUBS 0.008053f
C68 B.t8 VSUBS 0.085461f
C69 B.t7 VSUBS 0.109105f
C70 B.t6 VSUBS 0.600846f
C71 B.n40 VSUBS 0.191746f
C72 B.n41 VSUBS 0.158778f
C73 B.n42 VSUBS 0.018659f
C74 B.n43 VSUBS 0.008053f
C75 B.n44 VSUBS 0.008053f
C76 B.n45 VSUBS 0.008053f
C77 B.n46 VSUBS 0.008053f
C78 B.t2 VSUBS 0.085463f
C79 B.t1 VSUBS 0.109106f
C80 B.t0 VSUBS 0.600846f
C81 B.n47 VSUBS 0.191744f
C82 B.n48 VSUBS 0.158776f
C83 B.n49 VSUBS 0.008053f
C84 B.n50 VSUBS 0.008053f
C85 B.n51 VSUBS 0.008053f
C86 B.n52 VSUBS 0.008053f
C87 B.n53 VSUBS 0.008053f
C88 B.n54 VSUBS 0.008053f
C89 B.n55 VSUBS 0.008053f
C90 B.n56 VSUBS 0.008053f
C91 B.n57 VSUBS 0.008053f
C92 B.n58 VSUBS 0.008053f
C93 B.n59 VSUBS 0.020215f
C94 B.n60 VSUBS 0.008053f
C95 B.n61 VSUBS 0.008053f
C96 B.n62 VSUBS 0.008053f
C97 B.n63 VSUBS 0.008053f
C98 B.n64 VSUBS 0.008053f
C99 B.n65 VSUBS 0.008053f
C100 B.n66 VSUBS 0.008053f
C101 B.n67 VSUBS 0.008053f
C102 B.n68 VSUBS 0.008053f
C103 B.n69 VSUBS 0.008053f
C104 B.n70 VSUBS 0.008053f
C105 B.n71 VSUBS 0.008053f
C106 B.n72 VSUBS 0.008053f
C107 B.n73 VSUBS 0.008053f
C108 B.n74 VSUBS 0.008053f
C109 B.n75 VSUBS 0.008053f
C110 B.n76 VSUBS 0.008053f
C111 B.n77 VSUBS 0.008053f
C112 B.n78 VSUBS 0.008053f
C113 B.n79 VSUBS 0.008053f
C114 B.n80 VSUBS 0.008053f
C115 B.n81 VSUBS 0.008053f
C116 B.n82 VSUBS 0.008053f
C117 B.n83 VSUBS 0.008053f
C118 B.n84 VSUBS 0.008053f
C119 B.n85 VSUBS 0.008053f
C120 B.n86 VSUBS 0.008053f
C121 B.n87 VSUBS 0.008053f
C122 B.n88 VSUBS 0.008053f
C123 B.n89 VSUBS 0.008053f
C124 B.n90 VSUBS 0.008053f
C125 B.n91 VSUBS 0.008053f
C126 B.n92 VSUBS 0.008053f
C127 B.n93 VSUBS 0.008053f
C128 B.n94 VSUBS 0.008053f
C129 B.n95 VSUBS 0.008053f
C130 B.n96 VSUBS 0.008053f
C131 B.n97 VSUBS 0.008053f
C132 B.n98 VSUBS 0.008053f
C133 B.n99 VSUBS 0.008053f
C134 B.n100 VSUBS 0.008053f
C135 B.n101 VSUBS 0.008053f
C136 B.n102 VSUBS 0.008053f
C137 B.n103 VSUBS 0.008053f
C138 B.n104 VSUBS 0.008053f
C139 B.n105 VSUBS 0.008053f
C140 B.n106 VSUBS 0.008053f
C141 B.n107 VSUBS 0.008053f
C142 B.n108 VSUBS 0.008053f
C143 B.n109 VSUBS 0.008053f
C144 B.n110 VSUBS 0.008053f
C145 B.n111 VSUBS 0.019323f
C146 B.n112 VSUBS 0.008053f
C147 B.n113 VSUBS 0.008053f
C148 B.n114 VSUBS 0.008053f
C149 B.n115 VSUBS 0.008053f
C150 B.n116 VSUBS 0.008053f
C151 B.n117 VSUBS 0.008053f
C152 B.n118 VSUBS 0.008053f
C153 B.n119 VSUBS 0.008053f
C154 B.n120 VSUBS 0.008053f
C155 B.n121 VSUBS 0.008053f
C156 B.n122 VSUBS 0.008053f
C157 B.t10 VSUBS 0.085463f
C158 B.t11 VSUBS 0.109106f
C159 B.t9 VSUBS 0.600846f
C160 B.n123 VSUBS 0.191744f
C161 B.n124 VSUBS 0.158776f
C162 B.n125 VSUBS 0.008053f
C163 B.n126 VSUBS 0.008053f
C164 B.n127 VSUBS 0.008053f
C165 B.n128 VSUBS 0.008053f
C166 B.t4 VSUBS 0.085461f
C167 B.t5 VSUBS 0.109105f
C168 B.t3 VSUBS 0.600846f
C169 B.n129 VSUBS 0.191746f
C170 B.n130 VSUBS 0.158778f
C171 B.n131 VSUBS 0.018659f
C172 B.n132 VSUBS 0.008053f
C173 B.n133 VSUBS 0.008053f
C174 B.n134 VSUBS 0.008053f
C175 B.n135 VSUBS 0.008053f
C176 B.n136 VSUBS 0.008053f
C177 B.n137 VSUBS 0.008053f
C178 B.n138 VSUBS 0.008053f
C179 B.n139 VSUBS 0.008053f
C180 B.n140 VSUBS 0.008053f
C181 B.n141 VSUBS 0.008053f
C182 B.n142 VSUBS 0.019323f
C183 B.n143 VSUBS 0.008053f
C184 B.n144 VSUBS 0.008053f
C185 B.n145 VSUBS 0.008053f
C186 B.n146 VSUBS 0.008053f
C187 B.n147 VSUBS 0.008053f
C188 B.n148 VSUBS 0.008053f
C189 B.n149 VSUBS 0.008053f
C190 B.n150 VSUBS 0.008053f
C191 B.n151 VSUBS 0.008053f
C192 B.n152 VSUBS 0.008053f
C193 B.n153 VSUBS 0.008053f
C194 B.n154 VSUBS 0.008053f
C195 B.n155 VSUBS 0.008053f
C196 B.n156 VSUBS 0.008053f
C197 B.n157 VSUBS 0.008053f
C198 B.n158 VSUBS 0.008053f
C199 B.n159 VSUBS 0.008053f
C200 B.n160 VSUBS 0.008053f
C201 B.n161 VSUBS 0.008053f
C202 B.n162 VSUBS 0.008053f
C203 B.n163 VSUBS 0.008053f
C204 B.n164 VSUBS 0.008053f
C205 B.n165 VSUBS 0.008053f
C206 B.n166 VSUBS 0.008053f
C207 B.n167 VSUBS 0.008053f
C208 B.n168 VSUBS 0.008053f
C209 B.n169 VSUBS 0.008053f
C210 B.n170 VSUBS 0.008053f
C211 B.n171 VSUBS 0.008053f
C212 B.n172 VSUBS 0.008053f
C213 B.n173 VSUBS 0.008053f
C214 B.n174 VSUBS 0.008053f
C215 B.n175 VSUBS 0.008053f
C216 B.n176 VSUBS 0.008053f
C217 B.n177 VSUBS 0.008053f
C218 B.n178 VSUBS 0.008053f
C219 B.n179 VSUBS 0.008053f
C220 B.n180 VSUBS 0.008053f
C221 B.n181 VSUBS 0.008053f
C222 B.n182 VSUBS 0.008053f
C223 B.n183 VSUBS 0.008053f
C224 B.n184 VSUBS 0.008053f
C225 B.n185 VSUBS 0.008053f
C226 B.n186 VSUBS 0.008053f
C227 B.n187 VSUBS 0.008053f
C228 B.n188 VSUBS 0.008053f
C229 B.n189 VSUBS 0.008053f
C230 B.n190 VSUBS 0.008053f
C231 B.n191 VSUBS 0.008053f
C232 B.n192 VSUBS 0.008053f
C233 B.n193 VSUBS 0.008053f
C234 B.n194 VSUBS 0.008053f
C235 B.n195 VSUBS 0.008053f
C236 B.n196 VSUBS 0.008053f
C237 B.n197 VSUBS 0.008053f
C238 B.n198 VSUBS 0.008053f
C239 B.n199 VSUBS 0.008053f
C240 B.n200 VSUBS 0.008053f
C241 B.n201 VSUBS 0.008053f
C242 B.n202 VSUBS 0.008053f
C243 B.n203 VSUBS 0.008053f
C244 B.n204 VSUBS 0.008053f
C245 B.n205 VSUBS 0.008053f
C246 B.n206 VSUBS 0.008053f
C247 B.n207 VSUBS 0.008053f
C248 B.n208 VSUBS 0.008053f
C249 B.n209 VSUBS 0.008053f
C250 B.n210 VSUBS 0.008053f
C251 B.n211 VSUBS 0.008053f
C252 B.n212 VSUBS 0.008053f
C253 B.n213 VSUBS 0.008053f
C254 B.n214 VSUBS 0.008053f
C255 B.n215 VSUBS 0.008053f
C256 B.n216 VSUBS 0.008053f
C257 B.n217 VSUBS 0.008053f
C258 B.n218 VSUBS 0.008053f
C259 B.n219 VSUBS 0.008053f
C260 B.n220 VSUBS 0.008053f
C261 B.n221 VSUBS 0.008053f
C262 B.n222 VSUBS 0.008053f
C263 B.n223 VSUBS 0.008053f
C264 B.n224 VSUBS 0.008053f
C265 B.n225 VSUBS 0.008053f
C266 B.n226 VSUBS 0.008053f
C267 B.n227 VSUBS 0.008053f
C268 B.n228 VSUBS 0.008053f
C269 B.n229 VSUBS 0.008053f
C270 B.n230 VSUBS 0.008053f
C271 B.n231 VSUBS 0.008053f
C272 B.n232 VSUBS 0.008053f
C273 B.n233 VSUBS 0.008053f
C274 B.n234 VSUBS 0.008053f
C275 B.n235 VSUBS 0.008053f
C276 B.n236 VSUBS 0.008053f
C277 B.n237 VSUBS 0.008053f
C278 B.n238 VSUBS 0.008053f
C279 B.n239 VSUBS 0.008053f
C280 B.n240 VSUBS 0.008053f
C281 B.n241 VSUBS 0.008053f
C282 B.n242 VSUBS 0.008053f
C283 B.n243 VSUBS 0.019323f
C284 B.n244 VSUBS 0.019997f
C285 B.n245 VSUBS 0.019997f
C286 B.n246 VSUBS 0.008053f
C287 B.n247 VSUBS 0.008053f
C288 B.n248 VSUBS 0.008053f
C289 B.n249 VSUBS 0.008053f
C290 B.n250 VSUBS 0.008053f
C291 B.n251 VSUBS 0.008053f
C292 B.n252 VSUBS 0.008053f
C293 B.n253 VSUBS 0.008053f
C294 B.n254 VSUBS 0.008053f
C295 B.n255 VSUBS 0.008053f
C296 B.n256 VSUBS 0.008053f
C297 B.n257 VSUBS 0.008053f
C298 B.n258 VSUBS 0.008053f
C299 B.n259 VSUBS 0.008053f
C300 B.n260 VSUBS 0.008053f
C301 B.n261 VSUBS 0.008053f
C302 B.n262 VSUBS 0.008053f
C303 B.n263 VSUBS 0.008053f
C304 B.n264 VSUBS 0.008053f
C305 B.n265 VSUBS 0.008053f
C306 B.n266 VSUBS 0.008053f
C307 B.n267 VSUBS 0.008053f
C308 B.n268 VSUBS 0.008053f
C309 B.n269 VSUBS 0.008053f
C310 B.n270 VSUBS 0.008053f
C311 B.n271 VSUBS 0.008053f
C312 B.n272 VSUBS 0.008053f
C313 B.n273 VSUBS 0.008053f
C314 B.n274 VSUBS 0.00758f
C315 B.n275 VSUBS 0.008053f
C316 B.n276 VSUBS 0.008053f
C317 B.n277 VSUBS 0.0045f
C318 B.n278 VSUBS 0.008053f
C319 B.n279 VSUBS 0.008053f
C320 B.n280 VSUBS 0.008053f
C321 B.n281 VSUBS 0.008053f
C322 B.n282 VSUBS 0.008053f
C323 B.n283 VSUBS 0.008053f
C324 B.n284 VSUBS 0.008053f
C325 B.n285 VSUBS 0.008053f
C326 B.n286 VSUBS 0.008053f
C327 B.n287 VSUBS 0.008053f
C328 B.n288 VSUBS 0.008053f
C329 B.n289 VSUBS 0.008053f
C330 B.n290 VSUBS 0.0045f
C331 B.n291 VSUBS 0.018659f
C332 B.n292 VSUBS 0.00758f
C333 B.n293 VSUBS 0.008053f
C334 B.n294 VSUBS 0.008053f
C335 B.n295 VSUBS 0.008053f
C336 B.n296 VSUBS 0.008053f
C337 B.n297 VSUBS 0.008053f
C338 B.n298 VSUBS 0.008053f
C339 B.n299 VSUBS 0.008053f
C340 B.n300 VSUBS 0.008053f
C341 B.n301 VSUBS 0.008053f
C342 B.n302 VSUBS 0.008053f
C343 B.n303 VSUBS 0.008053f
C344 B.n304 VSUBS 0.008053f
C345 B.n305 VSUBS 0.008053f
C346 B.n306 VSUBS 0.008053f
C347 B.n307 VSUBS 0.008053f
C348 B.n308 VSUBS 0.008053f
C349 B.n309 VSUBS 0.008053f
C350 B.n310 VSUBS 0.008053f
C351 B.n311 VSUBS 0.008053f
C352 B.n312 VSUBS 0.008053f
C353 B.n313 VSUBS 0.008053f
C354 B.n314 VSUBS 0.008053f
C355 B.n315 VSUBS 0.008053f
C356 B.n316 VSUBS 0.008053f
C357 B.n317 VSUBS 0.008053f
C358 B.n318 VSUBS 0.008053f
C359 B.n319 VSUBS 0.008053f
C360 B.n320 VSUBS 0.008053f
C361 B.n321 VSUBS 0.008053f
C362 B.n322 VSUBS 0.019997f
C363 B.n323 VSUBS 0.019997f
C364 B.n324 VSUBS 0.019323f
C365 B.n325 VSUBS 0.008053f
C366 B.n326 VSUBS 0.008053f
C367 B.n327 VSUBS 0.008053f
C368 B.n328 VSUBS 0.008053f
C369 B.n329 VSUBS 0.008053f
C370 B.n330 VSUBS 0.008053f
C371 B.n331 VSUBS 0.008053f
C372 B.n332 VSUBS 0.008053f
C373 B.n333 VSUBS 0.008053f
C374 B.n334 VSUBS 0.008053f
C375 B.n335 VSUBS 0.008053f
C376 B.n336 VSUBS 0.008053f
C377 B.n337 VSUBS 0.008053f
C378 B.n338 VSUBS 0.008053f
C379 B.n339 VSUBS 0.008053f
C380 B.n340 VSUBS 0.008053f
C381 B.n341 VSUBS 0.008053f
C382 B.n342 VSUBS 0.008053f
C383 B.n343 VSUBS 0.008053f
C384 B.n344 VSUBS 0.008053f
C385 B.n345 VSUBS 0.008053f
C386 B.n346 VSUBS 0.008053f
C387 B.n347 VSUBS 0.008053f
C388 B.n348 VSUBS 0.008053f
C389 B.n349 VSUBS 0.008053f
C390 B.n350 VSUBS 0.008053f
C391 B.n351 VSUBS 0.008053f
C392 B.n352 VSUBS 0.008053f
C393 B.n353 VSUBS 0.008053f
C394 B.n354 VSUBS 0.008053f
C395 B.n355 VSUBS 0.008053f
C396 B.n356 VSUBS 0.008053f
C397 B.n357 VSUBS 0.008053f
C398 B.n358 VSUBS 0.008053f
C399 B.n359 VSUBS 0.008053f
C400 B.n360 VSUBS 0.008053f
C401 B.n361 VSUBS 0.008053f
C402 B.n362 VSUBS 0.008053f
C403 B.n363 VSUBS 0.008053f
C404 B.n364 VSUBS 0.008053f
C405 B.n365 VSUBS 0.008053f
C406 B.n366 VSUBS 0.008053f
C407 B.n367 VSUBS 0.008053f
C408 B.n368 VSUBS 0.008053f
C409 B.n369 VSUBS 0.008053f
C410 B.n370 VSUBS 0.008053f
C411 B.n371 VSUBS 0.008053f
C412 B.n372 VSUBS 0.008053f
C413 B.n373 VSUBS 0.008053f
C414 B.n374 VSUBS 0.008053f
C415 B.n375 VSUBS 0.008053f
C416 B.n376 VSUBS 0.008053f
C417 B.n377 VSUBS 0.008053f
C418 B.n378 VSUBS 0.008053f
C419 B.n379 VSUBS 0.008053f
C420 B.n380 VSUBS 0.008053f
C421 B.n381 VSUBS 0.008053f
C422 B.n382 VSUBS 0.008053f
C423 B.n383 VSUBS 0.008053f
C424 B.n384 VSUBS 0.008053f
C425 B.n385 VSUBS 0.008053f
C426 B.n386 VSUBS 0.008053f
C427 B.n387 VSUBS 0.008053f
C428 B.n388 VSUBS 0.008053f
C429 B.n389 VSUBS 0.008053f
C430 B.n390 VSUBS 0.008053f
C431 B.n391 VSUBS 0.008053f
C432 B.n392 VSUBS 0.008053f
C433 B.n393 VSUBS 0.008053f
C434 B.n394 VSUBS 0.008053f
C435 B.n395 VSUBS 0.008053f
C436 B.n396 VSUBS 0.008053f
C437 B.n397 VSUBS 0.008053f
C438 B.n398 VSUBS 0.008053f
C439 B.n399 VSUBS 0.008053f
C440 B.n400 VSUBS 0.008053f
C441 B.n401 VSUBS 0.008053f
C442 B.n402 VSUBS 0.008053f
C443 B.n403 VSUBS 0.008053f
C444 B.n404 VSUBS 0.008053f
C445 B.n405 VSUBS 0.008053f
C446 B.n406 VSUBS 0.008053f
C447 B.n407 VSUBS 0.008053f
C448 B.n408 VSUBS 0.008053f
C449 B.n409 VSUBS 0.008053f
C450 B.n410 VSUBS 0.008053f
C451 B.n411 VSUBS 0.008053f
C452 B.n412 VSUBS 0.008053f
C453 B.n413 VSUBS 0.008053f
C454 B.n414 VSUBS 0.008053f
C455 B.n415 VSUBS 0.008053f
C456 B.n416 VSUBS 0.008053f
C457 B.n417 VSUBS 0.008053f
C458 B.n418 VSUBS 0.008053f
C459 B.n419 VSUBS 0.008053f
C460 B.n420 VSUBS 0.008053f
C461 B.n421 VSUBS 0.008053f
C462 B.n422 VSUBS 0.008053f
C463 B.n423 VSUBS 0.008053f
C464 B.n424 VSUBS 0.008053f
C465 B.n425 VSUBS 0.008053f
C466 B.n426 VSUBS 0.008053f
C467 B.n427 VSUBS 0.008053f
C468 B.n428 VSUBS 0.008053f
C469 B.n429 VSUBS 0.008053f
C470 B.n430 VSUBS 0.008053f
C471 B.n431 VSUBS 0.008053f
C472 B.n432 VSUBS 0.008053f
C473 B.n433 VSUBS 0.008053f
C474 B.n434 VSUBS 0.008053f
C475 B.n435 VSUBS 0.008053f
C476 B.n436 VSUBS 0.008053f
C477 B.n437 VSUBS 0.008053f
C478 B.n438 VSUBS 0.008053f
C479 B.n439 VSUBS 0.008053f
C480 B.n440 VSUBS 0.008053f
C481 B.n441 VSUBS 0.008053f
C482 B.n442 VSUBS 0.008053f
C483 B.n443 VSUBS 0.008053f
C484 B.n444 VSUBS 0.008053f
C485 B.n445 VSUBS 0.008053f
C486 B.n446 VSUBS 0.008053f
C487 B.n447 VSUBS 0.008053f
C488 B.n448 VSUBS 0.008053f
C489 B.n449 VSUBS 0.008053f
C490 B.n450 VSUBS 0.008053f
C491 B.n451 VSUBS 0.008053f
C492 B.n452 VSUBS 0.008053f
C493 B.n453 VSUBS 0.008053f
C494 B.n454 VSUBS 0.008053f
C495 B.n455 VSUBS 0.008053f
C496 B.n456 VSUBS 0.008053f
C497 B.n457 VSUBS 0.008053f
C498 B.n458 VSUBS 0.008053f
C499 B.n459 VSUBS 0.008053f
C500 B.n460 VSUBS 0.008053f
C501 B.n461 VSUBS 0.008053f
C502 B.n462 VSUBS 0.008053f
C503 B.n463 VSUBS 0.008053f
C504 B.n464 VSUBS 0.008053f
C505 B.n465 VSUBS 0.008053f
C506 B.n466 VSUBS 0.008053f
C507 B.n467 VSUBS 0.008053f
C508 B.n468 VSUBS 0.008053f
C509 B.n469 VSUBS 0.008053f
C510 B.n470 VSUBS 0.008053f
C511 B.n471 VSUBS 0.008053f
C512 B.n472 VSUBS 0.008053f
C513 B.n473 VSUBS 0.008053f
C514 B.n474 VSUBS 0.008053f
C515 B.n475 VSUBS 0.008053f
C516 B.n476 VSUBS 0.008053f
C517 B.n477 VSUBS 0.008053f
C518 B.n478 VSUBS 0.008053f
C519 B.n479 VSUBS 0.008053f
C520 B.n480 VSUBS 0.019323f
C521 B.n481 VSUBS 0.019997f
C522 B.n482 VSUBS 0.019105f
C523 B.n483 VSUBS 0.008053f
C524 B.n484 VSUBS 0.008053f
C525 B.n485 VSUBS 0.008053f
C526 B.n486 VSUBS 0.008053f
C527 B.n487 VSUBS 0.008053f
C528 B.n488 VSUBS 0.008053f
C529 B.n489 VSUBS 0.008053f
C530 B.n490 VSUBS 0.008053f
C531 B.n491 VSUBS 0.008053f
C532 B.n492 VSUBS 0.008053f
C533 B.n493 VSUBS 0.008053f
C534 B.n494 VSUBS 0.008053f
C535 B.n495 VSUBS 0.008053f
C536 B.n496 VSUBS 0.008053f
C537 B.n497 VSUBS 0.008053f
C538 B.n498 VSUBS 0.008053f
C539 B.n499 VSUBS 0.008053f
C540 B.n500 VSUBS 0.008053f
C541 B.n501 VSUBS 0.008053f
C542 B.n502 VSUBS 0.008053f
C543 B.n503 VSUBS 0.008053f
C544 B.n504 VSUBS 0.008053f
C545 B.n505 VSUBS 0.008053f
C546 B.n506 VSUBS 0.008053f
C547 B.n507 VSUBS 0.008053f
C548 B.n508 VSUBS 0.008053f
C549 B.n509 VSUBS 0.008053f
C550 B.n510 VSUBS 0.008053f
C551 B.n511 VSUBS 0.008053f
C552 B.n512 VSUBS 0.00758f
C553 B.n513 VSUBS 0.018659f
C554 B.n514 VSUBS 0.0045f
C555 B.n515 VSUBS 0.008053f
C556 B.n516 VSUBS 0.008053f
C557 B.n517 VSUBS 0.008053f
C558 B.n518 VSUBS 0.008053f
C559 B.n519 VSUBS 0.008053f
C560 B.n520 VSUBS 0.008053f
C561 B.n521 VSUBS 0.008053f
C562 B.n522 VSUBS 0.008053f
C563 B.n523 VSUBS 0.008053f
C564 B.n524 VSUBS 0.008053f
C565 B.n525 VSUBS 0.008053f
C566 B.n526 VSUBS 0.008053f
C567 B.n527 VSUBS 0.0045f
C568 B.n528 VSUBS 0.008053f
C569 B.n529 VSUBS 0.008053f
C570 B.n530 VSUBS 0.008053f
C571 B.n531 VSUBS 0.008053f
C572 B.n532 VSUBS 0.008053f
C573 B.n533 VSUBS 0.008053f
C574 B.n534 VSUBS 0.008053f
C575 B.n535 VSUBS 0.008053f
C576 B.n536 VSUBS 0.008053f
C577 B.n537 VSUBS 0.008053f
C578 B.n538 VSUBS 0.008053f
C579 B.n539 VSUBS 0.008053f
C580 B.n540 VSUBS 0.008053f
C581 B.n541 VSUBS 0.008053f
C582 B.n542 VSUBS 0.008053f
C583 B.n543 VSUBS 0.008053f
C584 B.n544 VSUBS 0.008053f
C585 B.n545 VSUBS 0.008053f
C586 B.n546 VSUBS 0.008053f
C587 B.n547 VSUBS 0.008053f
C588 B.n548 VSUBS 0.008053f
C589 B.n549 VSUBS 0.008053f
C590 B.n550 VSUBS 0.008053f
C591 B.n551 VSUBS 0.008053f
C592 B.n552 VSUBS 0.008053f
C593 B.n553 VSUBS 0.008053f
C594 B.n554 VSUBS 0.008053f
C595 B.n555 VSUBS 0.008053f
C596 B.n556 VSUBS 0.008053f
C597 B.n557 VSUBS 0.008053f
C598 B.n558 VSUBS 0.008053f
C599 B.n559 VSUBS 0.019997f
C600 B.n560 VSUBS 0.019323f
C601 B.n561 VSUBS 0.019323f
C602 B.n562 VSUBS 0.008053f
C603 B.n563 VSUBS 0.008053f
C604 B.n564 VSUBS 0.008053f
C605 B.n565 VSUBS 0.008053f
C606 B.n566 VSUBS 0.008053f
C607 B.n567 VSUBS 0.008053f
C608 B.n568 VSUBS 0.008053f
C609 B.n569 VSUBS 0.008053f
C610 B.n570 VSUBS 0.008053f
C611 B.n571 VSUBS 0.008053f
C612 B.n572 VSUBS 0.008053f
C613 B.n573 VSUBS 0.008053f
C614 B.n574 VSUBS 0.008053f
C615 B.n575 VSUBS 0.008053f
C616 B.n576 VSUBS 0.008053f
C617 B.n577 VSUBS 0.008053f
C618 B.n578 VSUBS 0.008053f
C619 B.n579 VSUBS 0.008053f
C620 B.n580 VSUBS 0.008053f
C621 B.n581 VSUBS 0.008053f
C622 B.n582 VSUBS 0.008053f
C623 B.n583 VSUBS 0.008053f
C624 B.n584 VSUBS 0.008053f
C625 B.n585 VSUBS 0.008053f
C626 B.n586 VSUBS 0.008053f
C627 B.n587 VSUBS 0.008053f
C628 B.n588 VSUBS 0.008053f
C629 B.n589 VSUBS 0.008053f
C630 B.n590 VSUBS 0.008053f
C631 B.n591 VSUBS 0.008053f
C632 B.n592 VSUBS 0.008053f
C633 B.n593 VSUBS 0.008053f
C634 B.n594 VSUBS 0.008053f
C635 B.n595 VSUBS 0.008053f
C636 B.n596 VSUBS 0.008053f
C637 B.n597 VSUBS 0.008053f
C638 B.n598 VSUBS 0.008053f
C639 B.n599 VSUBS 0.008053f
C640 B.n600 VSUBS 0.008053f
C641 B.n601 VSUBS 0.008053f
C642 B.n602 VSUBS 0.008053f
C643 B.n603 VSUBS 0.008053f
C644 B.n604 VSUBS 0.008053f
C645 B.n605 VSUBS 0.008053f
C646 B.n606 VSUBS 0.008053f
C647 B.n607 VSUBS 0.008053f
C648 B.n608 VSUBS 0.008053f
C649 B.n609 VSUBS 0.008053f
C650 B.n610 VSUBS 0.008053f
C651 B.n611 VSUBS 0.008053f
C652 B.n612 VSUBS 0.008053f
C653 B.n613 VSUBS 0.008053f
C654 B.n614 VSUBS 0.008053f
C655 B.n615 VSUBS 0.008053f
C656 B.n616 VSUBS 0.008053f
C657 B.n617 VSUBS 0.008053f
C658 B.n618 VSUBS 0.008053f
C659 B.n619 VSUBS 0.008053f
C660 B.n620 VSUBS 0.008053f
C661 B.n621 VSUBS 0.008053f
C662 B.n622 VSUBS 0.008053f
C663 B.n623 VSUBS 0.008053f
C664 B.n624 VSUBS 0.008053f
C665 B.n625 VSUBS 0.008053f
C666 B.n626 VSUBS 0.008053f
C667 B.n627 VSUBS 0.008053f
C668 B.n628 VSUBS 0.008053f
C669 B.n629 VSUBS 0.008053f
C670 B.n630 VSUBS 0.008053f
C671 B.n631 VSUBS 0.008053f
C672 B.n632 VSUBS 0.008053f
C673 B.n633 VSUBS 0.008053f
C674 B.n634 VSUBS 0.008053f
C675 B.n635 VSUBS 0.008053f
C676 B.n636 VSUBS 0.008053f
C677 B.n637 VSUBS 0.008053f
C678 B.n638 VSUBS 0.008053f
C679 B.n639 VSUBS 0.018236f
C680 VDD2.n0 VSUBS 0.01539f
C681 VDD2.n1 VSUBS 0.034669f
C682 VDD2.n2 VSUBS 0.015531f
C683 VDD2.n3 VSUBS 0.027296f
C684 VDD2.n4 VSUBS 0.014668f
C685 VDD2.n5 VSUBS 0.034669f
C686 VDD2.n6 VSUBS 0.015531f
C687 VDD2.n7 VSUBS 0.130712f
C688 VDD2.t7 VSUBS 0.074909f
C689 VDD2.n8 VSUBS 0.026002f
C690 VDD2.n9 VSUBS 0.026048f
C691 VDD2.n10 VSUBS 0.014668f
C692 VDD2.n11 VSUBS 0.516833f
C693 VDD2.n12 VSUBS 0.027296f
C694 VDD2.n13 VSUBS 0.014668f
C695 VDD2.n14 VSUBS 0.015531f
C696 VDD2.n15 VSUBS 0.034669f
C697 VDD2.n16 VSUBS 0.034669f
C698 VDD2.n17 VSUBS 0.015531f
C699 VDD2.n18 VSUBS 0.014668f
C700 VDD2.n19 VSUBS 0.027296f
C701 VDD2.n20 VSUBS 0.070552f
C702 VDD2.n21 VSUBS 0.014668f
C703 VDD2.n22 VSUBS 0.015531f
C704 VDD2.n23 VSUBS 0.075659f
C705 VDD2.n24 VSUBS 0.080015f
C706 VDD2.t5 VSUBS 0.11044f
C707 VDD2.t2 VSUBS 0.11044f
C708 VDD2.n25 VSUBS 0.717107f
C709 VDD2.n26 VSUBS 0.869271f
C710 VDD2.t0 VSUBS 0.11044f
C711 VDD2.t8 VSUBS 0.11044f
C712 VDD2.n27 VSUBS 0.728395f
C713 VDD2.n28 VSUBS 2.64768f
C714 VDD2.n29 VSUBS 0.01539f
C715 VDD2.n30 VSUBS 0.034669f
C716 VDD2.n31 VSUBS 0.015531f
C717 VDD2.n32 VSUBS 0.027296f
C718 VDD2.n33 VSUBS 0.014668f
C719 VDD2.n34 VSUBS 0.034669f
C720 VDD2.n35 VSUBS 0.015531f
C721 VDD2.n36 VSUBS 0.130712f
C722 VDD2.t1 VSUBS 0.074909f
C723 VDD2.n37 VSUBS 0.026002f
C724 VDD2.n38 VSUBS 0.026048f
C725 VDD2.n39 VSUBS 0.014668f
C726 VDD2.n40 VSUBS 0.516833f
C727 VDD2.n41 VSUBS 0.027296f
C728 VDD2.n42 VSUBS 0.014668f
C729 VDD2.n43 VSUBS 0.015531f
C730 VDD2.n44 VSUBS 0.034669f
C731 VDD2.n45 VSUBS 0.034669f
C732 VDD2.n46 VSUBS 0.015531f
C733 VDD2.n47 VSUBS 0.014668f
C734 VDD2.n48 VSUBS 0.027296f
C735 VDD2.n49 VSUBS 0.070552f
C736 VDD2.n50 VSUBS 0.014668f
C737 VDD2.n51 VSUBS 0.015531f
C738 VDD2.n52 VSUBS 0.075659f
C739 VDD2.n53 VSUBS 0.070144f
C740 VDD2.n54 VSUBS 2.38174f
C741 VDD2.t9 VSUBS 0.11044f
C742 VDD2.t3 VSUBS 0.11044f
C743 VDD2.n55 VSUBS 0.71711f
C744 VDD2.n56 VSUBS 0.644316f
C745 VDD2.t4 VSUBS 0.11044f
C746 VDD2.t6 VSUBS 0.11044f
C747 VDD2.n57 VSUBS 0.728364f
C748 VN.n0 VSUBS 0.053326f
C749 VN.t1 VSUBS 1.17205f
C750 VN.n1 VSUBS 0.032786f
C751 VN.n2 VSUBS 0.04045f
C752 VN.t9 VSUBS 1.17205f
C753 VN.n3 VSUBS 0.080165f
C754 VN.n4 VSUBS 0.04045f
C755 VN.t7 VSUBS 1.17205f
C756 VN.n5 VSUBS 0.454919f
C757 VN.n6 VSUBS 0.04045f
C758 VN.n7 VSUBS 0.080165f
C759 VN.t2 VSUBS 1.40948f
C760 VN.n8 VSUBS 0.546705f
C761 VN.t4 VSUBS 1.17205f
C762 VN.n9 VSUBS 0.556849f
C763 VN.n10 VSUBS 0.055755f
C764 VN.n11 VSUBS 0.342178f
C765 VN.n12 VSUBS 0.04045f
C766 VN.n13 VSUBS 0.04045f
C767 VN.n14 VSUBS 0.032683f
C768 VN.n15 VSUBS 0.079763f
C769 VN.n16 VSUBS 0.056495f
C770 VN.n17 VSUBS 0.04045f
C771 VN.n18 VSUBS 0.04045f
C772 VN.n19 VSUBS 0.056495f
C773 VN.n20 VSUBS 0.079763f
C774 VN.n21 VSUBS 0.032683f
C775 VN.n22 VSUBS 0.04045f
C776 VN.n23 VSUBS 0.04045f
C777 VN.n24 VSUBS 0.04045f
C778 VN.n25 VSUBS 0.055755f
C779 VN.n26 VSUBS 0.454919f
C780 VN.n27 VSUBS 0.057236f
C781 VN.n28 VSUBS 0.079312f
C782 VN.n29 VSUBS 0.04045f
C783 VN.n30 VSUBS 0.04045f
C784 VN.n31 VSUBS 0.04045f
C785 VN.n32 VSUBS 0.080512f
C786 VN.n33 VSUBS 0.055014f
C787 VN.n34 VSUBS 0.568257f
C788 VN.n35 VSUBS 0.059199f
C789 VN.n36 VSUBS 0.053326f
C790 VN.t8 VSUBS 1.17205f
C791 VN.n37 VSUBS 0.032786f
C792 VN.n38 VSUBS 0.04045f
C793 VN.t0 VSUBS 1.17205f
C794 VN.n39 VSUBS 0.080165f
C795 VN.n40 VSUBS 0.04045f
C796 VN.t6 VSUBS 1.17205f
C797 VN.n41 VSUBS 0.454919f
C798 VN.n42 VSUBS 0.04045f
C799 VN.n43 VSUBS 0.080165f
C800 VN.t3 VSUBS 1.40948f
C801 VN.n44 VSUBS 0.546705f
C802 VN.t5 VSUBS 1.17205f
C803 VN.n45 VSUBS 0.556849f
C804 VN.n46 VSUBS 0.055755f
C805 VN.n47 VSUBS 0.342178f
C806 VN.n48 VSUBS 0.04045f
C807 VN.n49 VSUBS 0.04045f
C808 VN.n50 VSUBS 0.032683f
C809 VN.n51 VSUBS 0.079763f
C810 VN.n52 VSUBS 0.056495f
C811 VN.n53 VSUBS 0.04045f
C812 VN.n54 VSUBS 0.04045f
C813 VN.n55 VSUBS 0.056495f
C814 VN.n56 VSUBS 0.079763f
C815 VN.n57 VSUBS 0.032683f
C816 VN.n58 VSUBS 0.04045f
C817 VN.n59 VSUBS 0.04045f
C818 VN.n60 VSUBS 0.04045f
C819 VN.n61 VSUBS 0.055755f
C820 VN.n62 VSUBS 0.454919f
C821 VN.n63 VSUBS 0.057236f
C822 VN.n64 VSUBS 0.079312f
C823 VN.n65 VSUBS 0.04045f
C824 VN.n66 VSUBS 0.04045f
C825 VN.n67 VSUBS 0.04045f
C826 VN.n68 VSUBS 0.080512f
C827 VN.n69 VSUBS 0.055014f
C828 VN.n70 VSUBS 0.568257f
C829 VN.n71 VSUBS 1.96237f
C830 VDD1.n0 VSUBS 0.015279f
C831 VDD1.n1 VSUBS 0.034421f
C832 VDD1.n2 VSUBS 0.01542f
C833 VDD1.n3 VSUBS 0.027101f
C834 VDD1.n4 VSUBS 0.014563f
C835 VDD1.n5 VSUBS 0.034421f
C836 VDD1.n6 VSUBS 0.01542f
C837 VDD1.n7 VSUBS 0.129777f
C838 VDD1.t5 VSUBS 0.074374f
C839 VDD1.n8 VSUBS 0.025816f
C840 VDD1.n9 VSUBS 0.025862f
C841 VDD1.n10 VSUBS 0.014563f
C842 VDD1.n11 VSUBS 0.513138f
C843 VDD1.n12 VSUBS 0.027101f
C844 VDD1.n13 VSUBS 0.014563f
C845 VDD1.n14 VSUBS 0.01542f
C846 VDD1.n15 VSUBS 0.034421f
C847 VDD1.n16 VSUBS 0.034421f
C848 VDD1.n17 VSUBS 0.01542f
C849 VDD1.n18 VSUBS 0.014563f
C850 VDD1.n19 VSUBS 0.027101f
C851 VDD1.n20 VSUBS 0.070047f
C852 VDD1.n21 VSUBS 0.014563f
C853 VDD1.n22 VSUBS 0.01542f
C854 VDD1.n23 VSUBS 0.075118f
C855 VDD1.n24 VSUBS 0.079443f
C856 VDD1.t3 VSUBS 0.10965f
C857 VDD1.t0 VSUBS 0.10965f
C858 VDD1.n25 VSUBS 0.711983f
C859 VDD1.n26 VSUBS 0.871662f
C860 VDD1.n27 VSUBS 0.015279f
C861 VDD1.n28 VSUBS 0.034421f
C862 VDD1.n29 VSUBS 0.01542f
C863 VDD1.n30 VSUBS 0.027101f
C864 VDD1.n31 VSUBS 0.014563f
C865 VDD1.n32 VSUBS 0.034421f
C866 VDD1.n33 VSUBS 0.01542f
C867 VDD1.n34 VSUBS 0.129777f
C868 VDD1.t6 VSUBS 0.074374f
C869 VDD1.n35 VSUBS 0.025816f
C870 VDD1.n36 VSUBS 0.025862f
C871 VDD1.n37 VSUBS 0.014563f
C872 VDD1.n38 VSUBS 0.513138f
C873 VDD1.n39 VSUBS 0.027101f
C874 VDD1.n40 VSUBS 0.014563f
C875 VDD1.n41 VSUBS 0.01542f
C876 VDD1.n42 VSUBS 0.034421f
C877 VDD1.n43 VSUBS 0.034421f
C878 VDD1.n44 VSUBS 0.01542f
C879 VDD1.n45 VSUBS 0.014563f
C880 VDD1.n46 VSUBS 0.027101f
C881 VDD1.n47 VSUBS 0.070047f
C882 VDD1.n48 VSUBS 0.014563f
C883 VDD1.n49 VSUBS 0.01542f
C884 VDD1.n50 VSUBS 0.075118f
C885 VDD1.n51 VSUBS 0.079443f
C886 VDD1.t7 VSUBS 0.10965f
C887 VDD1.t8 VSUBS 0.10965f
C888 VDD1.n52 VSUBS 0.71198f
C889 VDD1.n53 VSUBS 0.863056f
C890 VDD1.t1 VSUBS 0.10965f
C891 VDD1.t4 VSUBS 0.10965f
C892 VDD1.n54 VSUBS 0.723187f
C893 VDD1.n55 VSUBS 2.74592f
C894 VDD1.t2 VSUBS 0.10965f
C895 VDD1.t9 VSUBS 0.10965f
C896 VDD1.n56 VSUBS 0.711979f
C897 VDD1.n57 VSUBS 2.84007f
C898 VTAIL.t1 VSUBS 0.136519f
C899 VTAIL.t2 VSUBS 0.136519f
C900 VTAIL.n0 VSUBS 0.788405f
C901 VTAIL.n1 VSUBS 0.899728f
C902 VTAIL.n2 VSUBS 0.019024f
C903 VTAIL.n3 VSUBS 0.042856f
C904 VTAIL.n4 VSUBS 0.019198f
C905 VTAIL.n5 VSUBS 0.033742f
C906 VTAIL.n6 VSUBS 0.018132f
C907 VTAIL.n7 VSUBS 0.042856f
C908 VTAIL.n8 VSUBS 0.019198f
C909 VTAIL.n9 VSUBS 0.161578f
C910 VTAIL.t7 VSUBS 0.092598f
C911 VTAIL.n10 VSUBS 0.032142f
C912 VTAIL.n11 VSUBS 0.032199f
C913 VTAIL.n12 VSUBS 0.018132f
C914 VTAIL.n13 VSUBS 0.638879f
C915 VTAIL.n14 VSUBS 0.033742f
C916 VTAIL.n15 VSUBS 0.018132f
C917 VTAIL.n16 VSUBS 0.019198f
C918 VTAIL.n17 VSUBS 0.042856f
C919 VTAIL.n18 VSUBS 0.042856f
C920 VTAIL.n19 VSUBS 0.019198f
C921 VTAIL.n20 VSUBS 0.018132f
C922 VTAIL.n21 VSUBS 0.033742f
C923 VTAIL.n22 VSUBS 0.087212f
C924 VTAIL.n23 VSUBS 0.018132f
C925 VTAIL.n24 VSUBS 0.019198f
C926 VTAIL.n25 VSUBS 0.093525f
C927 VTAIL.n26 VSUBS 0.063444f
C928 VTAIL.n27 VSUBS 0.432578f
C929 VTAIL.t10 VSUBS 0.136519f
C930 VTAIL.t9 VSUBS 0.136519f
C931 VTAIL.n28 VSUBS 0.788405f
C932 VTAIL.n29 VSUBS 1.01736f
C933 VTAIL.t15 VSUBS 0.136519f
C934 VTAIL.t14 VSUBS 0.136519f
C935 VTAIL.n30 VSUBS 0.788405f
C936 VTAIL.n31 VSUBS 2.18897f
C937 VTAIL.t18 VSUBS 0.136519f
C938 VTAIL.t0 VSUBS 0.136519f
C939 VTAIL.n32 VSUBS 0.78841f
C940 VTAIL.n33 VSUBS 2.18896f
C941 VTAIL.t4 VSUBS 0.136519f
C942 VTAIL.t5 VSUBS 0.136519f
C943 VTAIL.n34 VSUBS 0.78841f
C944 VTAIL.n35 VSUBS 1.01735f
C945 VTAIL.n36 VSUBS 0.019024f
C946 VTAIL.n37 VSUBS 0.042856f
C947 VTAIL.n38 VSUBS 0.019198f
C948 VTAIL.n39 VSUBS 0.033742f
C949 VTAIL.n40 VSUBS 0.018132f
C950 VTAIL.n41 VSUBS 0.042856f
C951 VTAIL.n42 VSUBS 0.019198f
C952 VTAIL.n43 VSUBS 0.161578f
C953 VTAIL.t17 VSUBS 0.092598f
C954 VTAIL.n44 VSUBS 0.032142f
C955 VTAIL.n45 VSUBS 0.032199f
C956 VTAIL.n46 VSUBS 0.018132f
C957 VTAIL.n47 VSUBS 0.638879f
C958 VTAIL.n48 VSUBS 0.033742f
C959 VTAIL.n49 VSUBS 0.018132f
C960 VTAIL.n50 VSUBS 0.019198f
C961 VTAIL.n51 VSUBS 0.042856f
C962 VTAIL.n52 VSUBS 0.042856f
C963 VTAIL.n53 VSUBS 0.019198f
C964 VTAIL.n54 VSUBS 0.018132f
C965 VTAIL.n55 VSUBS 0.033742f
C966 VTAIL.n56 VSUBS 0.087212f
C967 VTAIL.n57 VSUBS 0.018132f
C968 VTAIL.n58 VSUBS 0.019198f
C969 VTAIL.n59 VSUBS 0.093525f
C970 VTAIL.n60 VSUBS 0.063444f
C971 VTAIL.n61 VSUBS 0.432578f
C972 VTAIL.t11 VSUBS 0.136519f
C973 VTAIL.t13 VSUBS 0.136519f
C974 VTAIL.n62 VSUBS 0.78841f
C975 VTAIL.n63 VSUBS 0.951743f
C976 VTAIL.t16 VSUBS 0.136519f
C977 VTAIL.t8 VSUBS 0.136519f
C978 VTAIL.n64 VSUBS 0.78841f
C979 VTAIL.n65 VSUBS 1.01735f
C980 VTAIL.n66 VSUBS 0.019024f
C981 VTAIL.n67 VSUBS 0.042856f
C982 VTAIL.n68 VSUBS 0.019198f
C983 VTAIL.n69 VSUBS 0.033742f
C984 VTAIL.n70 VSUBS 0.018132f
C985 VTAIL.n71 VSUBS 0.042856f
C986 VTAIL.n72 VSUBS 0.019198f
C987 VTAIL.n73 VSUBS 0.161578f
C988 VTAIL.t12 VSUBS 0.092598f
C989 VTAIL.n74 VSUBS 0.032142f
C990 VTAIL.n75 VSUBS 0.032199f
C991 VTAIL.n76 VSUBS 0.018132f
C992 VTAIL.n77 VSUBS 0.638879f
C993 VTAIL.n78 VSUBS 0.033742f
C994 VTAIL.n79 VSUBS 0.018132f
C995 VTAIL.n80 VSUBS 0.019198f
C996 VTAIL.n81 VSUBS 0.042856f
C997 VTAIL.n82 VSUBS 0.042856f
C998 VTAIL.n83 VSUBS 0.019198f
C999 VTAIL.n84 VSUBS 0.018132f
C1000 VTAIL.n85 VSUBS 0.033742f
C1001 VTAIL.n86 VSUBS 0.087212f
C1002 VTAIL.n87 VSUBS 0.018132f
C1003 VTAIL.n88 VSUBS 0.019198f
C1004 VTAIL.n89 VSUBS 0.093525f
C1005 VTAIL.n90 VSUBS 0.063444f
C1006 VTAIL.n91 VSUBS 1.43642f
C1007 VTAIL.n92 VSUBS 0.019024f
C1008 VTAIL.n93 VSUBS 0.042856f
C1009 VTAIL.n94 VSUBS 0.019198f
C1010 VTAIL.n95 VSUBS 0.033742f
C1011 VTAIL.n96 VSUBS 0.018132f
C1012 VTAIL.n97 VSUBS 0.042856f
C1013 VTAIL.n98 VSUBS 0.019198f
C1014 VTAIL.n99 VSUBS 0.161578f
C1015 VTAIL.t3 VSUBS 0.092598f
C1016 VTAIL.n100 VSUBS 0.032142f
C1017 VTAIL.n101 VSUBS 0.032199f
C1018 VTAIL.n102 VSUBS 0.018132f
C1019 VTAIL.n103 VSUBS 0.638879f
C1020 VTAIL.n104 VSUBS 0.033742f
C1021 VTAIL.n105 VSUBS 0.018132f
C1022 VTAIL.n106 VSUBS 0.019198f
C1023 VTAIL.n107 VSUBS 0.042856f
C1024 VTAIL.n108 VSUBS 0.042856f
C1025 VTAIL.n109 VSUBS 0.019198f
C1026 VTAIL.n110 VSUBS 0.018132f
C1027 VTAIL.n111 VSUBS 0.033742f
C1028 VTAIL.n112 VSUBS 0.087212f
C1029 VTAIL.n113 VSUBS 0.018132f
C1030 VTAIL.n114 VSUBS 0.019198f
C1031 VTAIL.n115 VSUBS 0.093525f
C1032 VTAIL.n116 VSUBS 0.063444f
C1033 VTAIL.n117 VSUBS 1.43642f
C1034 VTAIL.t6 VSUBS 0.136519f
C1035 VTAIL.t19 VSUBS 0.136519f
C1036 VTAIL.n118 VSUBS 0.788405f
C1037 VTAIL.n119 VSUBS 0.835993f
C1038 VP.n0 VSUBS 0.055158f
C1039 VP.t5 VSUBS 1.21231f
C1040 VP.n1 VSUBS 0.033912f
C1041 VP.n2 VSUBS 0.041839f
C1042 VP.t8 VSUBS 1.21231f
C1043 VP.n3 VSUBS 0.082918f
C1044 VP.n4 VSUBS 0.041839f
C1045 VP.t1 VSUBS 1.21231f
C1046 VP.n5 VSUBS 0.470547f
C1047 VP.n6 VSUBS 0.041839f
C1048 VP.n7 VSUBS 0.082918f
C1049 VP.n8 VSUBS 0.041839f
C1050 VP.t2 VSUBS 1.21231f
C1051 VP.n9 VSUBS 0.033912f
C1052 VP.n10 VSUBS 0.055158f
C1053 VP.t3 VSUBS 1.21231f
C1054 VP.n11 VSUBS 0.055158f
C1055 VP.t0 VSUBS 1.21231f
C1056 VP.n12 VSUBS 0.033912f
C1057 VP.n13 VSUBS 0.041839f
C1058 VP.t7 VSUBS 1.21231f
C1059 VP.n14 VSUBS 0.082918f
C1060 VP.n15 VSUBS 0.041839f
C1061 VP.t9 VSUBS 1.21231f
C1062 VP.n16 VSUBS 0.470547f
C1063 VP.n17 VSUBS 0.041839f
C1064 VP.n18 VSUBS 0.082918f
C1065 VP.t4 VSUBS 1.4579f
C1066 VP.n19 VSUBS 0.565486f
C1067 VP.t6 VSUBS 1.21231f
C1068 VP.n20 VSUBS 0.575978f
C1069 VP.n21 VSUBS 0.05767f
C1070 VP.n22 VSUBS 0.353933f
C1071 VP.n23 VSUBS 0.041839f
C1072 VP.n24 VSUBS 0.041839f
C1073 VP.n25 VSUBS 0.033806f
C1074 VP.n26 VSUBS 0.082503f
C1075 VP.n27 VSUBS 0.058436f
C1076 VP.n28 VSUBS 0.041839f
C1077 VP.n29 VSUBS 0.041839f
C1078 VP.n30 VSUBS 0.058436f
C1079 VP.n31 VSUBS 0.082503f
C1080 VP.n32 VSUBS 0.033806f
C1081 VP.n33 VSUBS 0.041839f
C1082 VP.n34 VSUBS 0.041839f
C1083 VP.n35 VSUBS 0.041839f
C1084 VP.n36 VSUBS 0.05767f
C1085 VP.n37 VSUBS 0.470547f
C1086 VP.n38 VSUBS 0.059202f
C1087 VP.n39 VSUBS 0.082037f
C1088 VP.n40 VSUBS 0.041839f
C1089 VP.n41 VSUBS 0.041839f
C1090 VP.n42 VSUBS 0.041839f
C1091 VP.n43 VSUBS 0.083278f
C1092 VP.n44 VSUBS 0.056904f
C1093 VP.n45 VSUBS 0.587779f
C1094 VP.n46 VSUBS 2.00694f
C1095 VP.n47 VSUBS 2.04013f
C1096 VP.n48 VSUBS 0.587779f
C1097 VP.n49 VSUBS 0.056904f
C1098 VP.n50 VSUBS 0.083278f
C1099 VP.n51 VSUBS 0.041839f
C1100 VP.n52 VSUBS 0.041839f
C1101 VP.n53 VSUBS 0.041839f
C1102 VP.n54 VSUBS 0.082037f
C1103 VP.n55 VSUBS 0.059202f
C1104 VP.n56 VSUBS 0.470547f
C1105 VP.n57 VSUBS 0.05767f
C1106 VP.n58 VSUBS 0.041839f
C1107 VP.n59 VSUBS 0.041839f
C1108 VP.n60 VSUBS 0.041839f
C1109 VP.n61 VSUBS 0.033806f
C1110 VP.n62 VSUBS 0.082503f
C1111 VP.n63 VSUBS 0.058436f
C1112 VP.n64 VSUBS 0.041839f
C1113 VP.n65 VSUBS 0.041839f
C1114 VP.n66 VSUBS 0.058436f
C1115 VP.n67 VSUBS 0.082503f
C1116 VP.n68 VSUBS 0.033806f
C1117 VP.n69 VSUBS 0.041839f
C1118 VP.n70 VSUBS 0.041839f
C1119 VP.n71 VSUBS 0.041839f
C1120 VP.n72 VSUBS 0.05767f
C1121 VP.n73 VSUBS 0.470547f
C1122 VP.n74 VSUBS 0.059202f
C1123 VP.n75 VSUBS 0.082037f
C1124 VP.n76 VSUBS 0.041839f
C1125 VP.n77 VSUBS 0.041839f
C1126 VP.n78 VSUBS 0.041839f
C1127 VP.n79 VSUBS 0.083278f
C1128 VP.n80 VSUBS 0.056904f
C1129 VP.n81 VSUBS 0.587779f
C1130 VP.n82 VSUBS 0.061232f
.ends

