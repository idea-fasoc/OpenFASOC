* NGSPICE file created from diff_pair_sample_0077.ext - technology: sky130A

.subckt diff_pair_sample_0077 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t3 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
X1 VTAIL.t4 VN.t0 VDD2.t7 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=2.8908 ps=17.85 w=17.52 l=2.49
X2 VDD2.t6 VN.t1 VTAIL.t2 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
X3 VDD2.t5 VN.t2 VTAIL.t1 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=6.8328 ps=35.82 w=17.52 l=2.49
X4 B.t11 B.t9 B.t10 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=0 ps=0 w=17.52 l=2.49
X5 B.t8 B.t6 B.t7 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=0 ps=0 w=17.52 l=2.49
X6 VTAIL.t0 VN.t3 VDD2.t4 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
X7 VDD1.t2 VP.t1 VTAIL.t14 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
X8 VTAIL.t5 VN.t4 VDD2.t3 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
X9 VDD2.t2 VN.t5 VTAIL.t6 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
X10 VDD2.t1 VN.t6 VTAIL.t3 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=6.8328 ps=35.82 w=17.52 l=2.49
X11 VTAIL.t7 VN.t7 VDD2.t0 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=2.8908 ps=17.85 w=17.52 l=2.49
X12 VDD1.t1 VP.t2 VTAIL.t13 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
X13 VTAIL.t12 VP.t3 VDD1.t0 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=2.8908 ps=17.85 w=17.52 l=2.49
X14 VTAIL.t11 VP.t4 VDD1.t7 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=2.8908 ps=17.85 w=17.52 l=2.49
X15 VDD1.t6 VP.t5 VTAIL.t10 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=6.8328 ps=35.82 w=17.52 l=2.49
X16 B.t5 B.t3 B.t4 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=0 ps=0 w=17.52 l=2.49
X17 VDD1.t5 VP.t6 VTAIL.t9 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=6.8328 ps=35.82 w=17.52 l=2.49
X18 B.t2 B.t0 B.t1 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=6.8328 pd=35.82 as=0 ps=0 w=17.52 l=2.49
X19 VTAIL.t8 VP.t7 VDD1.t4 w_n3790_n4472# sky130_fd_pr__pfet_01v8 ad=2.8908 pd=17.85 as=2.8908 ps=17.85 w=17.52 l=2.49
R0 VP.n16 VP.t3 203.607
R1 VP.n9 VP.t4 169.571
R2 VP.n47 VP.t2 169.571
R3 VP.n3 VP.t7 169.571
R4 VP.n65 VP.t6 169.571
R5 VP.n35 VP.t5 169.571
R6 VP.n13 VP.t0 169.571
R7 VP.n17 VP.t1 169.571
R8 VP.n19 VP.n18 161.3
R9 VP.n20 VP.n15 161.3
R10 VP.n22 VP.n21 161.3
R11 VP.n23 VP.n14 161.3
R12 VP.n25 VP.n24 161.3
R13 VP.n27 VP.n26 161.3
R14 VP.n28 VP.n12 161.3
R15 VP.n30 VP.n29 161.3
R16 VP.n31 VP.n11 161.3
R17 VP.n33 VP.n32 161.3
R18 VP.n34 VP.n10 161.3
R19 VP.n64 VP.n0 161.3
R20 VP.n63 VP.n62 161.3
R21 VP.n61 VP.n1 161.3
R22 VP.n60 VP.n59 161.3
R23 VP.n58 VP.n2 161.3
R24 VP.n57 VP.n56 161.3
R25 VP.n55 VP.n54 161.3
R26 VP.n53 VP.n4 161.3
R27 VP.n52 VP.n51 161.3
R28 VP.n50 VP.n5 161.3
R29 VP.n49 VP.n48 161.3
R30 VP.n46 VP.n6 161.3
R31 VP.n45 VP.n44 161.3
R32 VP.n43 VP.n7 161.3
R33 VP.n42 VP.n41 161.3
R34 VP.n40 VP.n8 161.3
R35 VP.n39 VP.n38 161.3
R36 VP.n37 VP.n9 99.596
R37 VP.n66 VP.n65 99.596
R38 VP.n36 VP.n35 99.596
R39 VP.n41 VP.n7 56.5617
R40 VP.n59 VP.n1 56.5617
R41 VP.n29 VP.n11 56.5617
R42 VP.n37 VP.n36 54.5754
R43 VP.n17 VP.n16 52.5962
R44 VP.n52 VP.n5 40.577
R45 VP.n53 VP.n52 40.577
R46 VP.n23 VP.n22 40.577
R47 VP.n22 VP.n15 40.577
R48 VP.n40 VP.n39 24.5923
R49 VP.n41 VP.n40 24.5923
R50 VP.n45 VP.n7 24.5923
R51 VP.n46 VP.n45 24.5923
R52 VP.n48 VP.n5 24.5923
R53 VP.n54 VP.n53 24.5923
R54 VP.n58 VP.n57 24.5923
R55 VP.n59 VP.n58 24.5923
R56 VP.n63 VP.n1 24.5923
R57 VP.n64 VP.n63 24.5923
R58 VP.n33 VP.n11 24.5923
R59 VP.n34 VP.n33 24.5923
R60 VP.n24 VP.n23 24.5923
R61 VP.n28 VP.n27 24.5923
R62 VP.n29 VP.n28 24.5923
R63 VP.n18 VP.n15 24.5923
R64 VP.n48 VP.n47 20.1658
R65 VP.n54 VP.n3 20.1658
R66 VP.n24 VP.n13 20.1658
R67 VP.n18 VP.n17 20.1658
R68 VP.n39 VP.n9 11.3127
R69 VP.n65 VP.n64 11.3127
R70 VP.n35 VP.n34 11.3127
R71 VP.n19 VP.n16 6.75133
R72 VP.n47 VP.n46 4.42703
R73 VP.n57 VP.n3 4.42703
R74 VP.n27 VP.n13 4.42703
R75 VP.n36 VP.n10 0.278335
R76 VP.n38 VP.n37 0.278335
R77 VP.n66 VP.n0 0.278335
R78 VP.n20 VP.n19 0.189894
R79 VP.n21 VP.n20 0.189894
R80 VP.n21 VP.n14 0.189894
R81 VP.n25 VP.n14 0.189894
R82 VP.n26 VP.n25 0.189894
R83 VP.n26 VP.n12 0.189894
R84 VP.n30 VP.n12 0.189894
R85 VP.n31 VP.n30 0.189894
R86 VP.n32 VP.n31 0.189894
R87 VP.n32 VP.n10 0.189894
R88 VP.n38 VP.n8 0.189894
R89 VP.n42 VP.n8 0.189894
R90 VP.n43 VP.n42 0.189894
R91 VP.n44 VP.n43 0.189894
R92 VP.n44 VP.n6 0.189894
R93 VP.n49 VP.n6 0.189894
R94 VP.n50 VP.n49 0.189894
R95 VP.n51 VP.n50 0.189894
R96 VP.n51 VP.n4 0.189894
R97 VP.n55 VP.n4 0.189894
R98 VP.n56 VP.n55 0.189894
R99 VP.n56 VP.n2 0.189894
R100 VP.n60 VP.n2 0.189894
R101 VP.n61 VP.n60 0.189894
R102 VP.n62 VP.n61 0.189894
R103 VP.n62 VP.n0 0.189894
R104 VP VP.n66 0.153485
R105 VDD1 VDD1.n0 70.2959
R106 VDD1.n3 VDD1.n2 70.1822
R107 VDD1.n3 VDD1.n1 70.1822
R108 VDD1.n5 VDD1.n4 69.022
R109 VDD1.n5 VDD1.n3 50.3414
R110 VDD1.n4 VDD1.t3 1.85581
R111 VDD1.n4 VDD1.t6 1.85581
R112 VDD1.n0 VDD1.t0 1.85581
R113 VDD1.n0 VDD1.t2 1.85581
R114 VDD1.n2 VDD1.t4 1.85581
R115 VDD1.n2 VDD1.t5 1.85581
R116 VDD1.n1 VDD1.t7 1.85581
R117 VDD1.n1 VDD1.t1 1.85581
R118 VDD1 VDD1.n5 1.15783
R119 VTAIL.n786 VTAIL.n694 756.745
R120 VTAIL.n94 VTAIL.n2 756.745
R121 VTAIL.n192 VTAIL.n100 756.745
R122 VTAIL.n292 VTAIL.n200 756.745
R123 VTAIL.n688 VTAIL.n596 756.745
R124 VTAIL.n588 VTAIL.n496 756.745
R125 VTAIL.n490 VTAIL.n398 756.745
R126 VTAIL.n390 VTAIL.n298 756.745
R127 VTAIL.n727 VTAIL.n726 585
R128 VTAIL.n729 VTAIL.n728 585
R129 VTAIL.n722 VTAIL.n721 585
R130 VTAIL.n735 VTAIL.n734 585
R131 VTAIL.n737 VTAIL.n736 585
R132 VTAIL.n718 VTAIL.n717 585
R133 VTAIL.n743 VTAIL.n742 585
R134 VTAIL.n745 VTAIL.n744 585
R135 VTAIL.n714 VTAIL.n713 585
R136 VTAIL.n751 VTAIL.n750 585
R137 VTAIL.n753 VTAIL.n752 585
R138 VTAIL.n710 VTAIL.n709 585
R139 VTAIL.n759 VTAIL.n758 585
R140 VTAIL.n761 VTAIL.n760 585
R141 VTAIL.n706 VTAIL.n705 585
R142 VTAIL.n768 VTAIL.n767 585
R143 VTAIL.n769 VTAIL.n704 585
R144 VTAIL.n771 VTAIL.n770 585
R145 VTAIL.n702 VTAIL.n701 585
R146 VTAIL.n777 VTAIL.n776 585
R147 VTAIL.n779 VTAIL.n778 585
R148 VTAIL.n698 VTAIL.n697 585
R149 VTAIL.n785 VTAIL.n784 585
R150 VTAIL.n787 VTAIL.n786 585
R151 VTAIL.n35 VTAIL.n34 585
R152 VTAIL.n37 VTAIL.n36 585
R153 VTAIL.n30 VTAIL.n29 585
R154 VTAIL.n43 VTAIL.n42 585
R155 VTAIL.n45 VTAIL.n44 585
R156 VTAIL.n26 VTAIL.n25 585
R157 VTAIL.n51 VTAIL.n50 585
R158 VTAIL.n53 VTAIL.n52 585
R159 VTAIL.n22 VTAIL.n21 585
R160 VTAIL.n59 VTAIL.n58 585
R161 VTAIL.n61 VTAIL.n60 585
R162 VTAIL.n18 VTAIL.n17 585
R163 VTAIL.n67 VTAIL.n66 585
R164 VTAIL.n69 VTAIL.n68 585
R165 VTAIL.n14 VTAIL.n13 585
R166 VTAIL.n76 VTAIL.n75 585
R167 VTAIL.n77 VTAIL.n12 585
R168 VTAIL.n79 VTAIL.n78 585
R169 VTAIL.n10 VTAIL.n9 585
R170 VTAIL.n85 VTAIL.n84 585
R171 VTAIL.n87 VTAIL.n86 585
R172 VTAIL.n6 VTAIL.n5 585
R173 VTAIL.n93 VTAIL.n92 585
R174 VTAIL.n95 VTAIL.n94 585
R175 VTAIL.n133 VTAIL.n132 585
R176 VTAIL.n135 VTAIL.n134 585
R177 VTAIL.n128 VTAIL.n127 585
R178 VTAIL.n141 VTAIL.n140 585
R179 VTAIL.n143 VTAIL.n142 585
R180 VTAIL.n124 VTAIL.n123 585
R181 VTAIL.n149 VTAIL.n148 585
R182 VTAIL.n151 VTAIL.n150 585
R183 VTAIL.n120 VTAIL.n119 585
R184 VTAIL.n157 VTAIL.n156 585
R185 VTAIL.n159 VTAIL.n158 585
R186 VTAIL.n116 VTAIL.n115 585
R187 VTAIL.n165 VTAIL.n164 585
R188 VTAIL.n167 VTAIL.n166 585
R189 VTAIL.n112 VTAIL.n111 585
R190 VTAIL.n174 VTAIL.n173 585
R191 VTAIL.n175 VTAIL.n110 585
R192 VTAIL.n177 VTAIL.n176 585
R193 VTAIL.n108 VTAIL.n107 585
R194 VTAIL.n183 VTAIL.n182 585
R195 VTAIL.n185 VTAIL.n184 585
R196 VTAIL.n104 VTAIL.n103 585
R197 VTAIL.n191 VTAIL.n190 585
R198 VTAIL.n193 VTAIL.n192 585
R199 VTAIL.n233 VTAIL.n232 585
R200 VTAIL.n235 VTAIL.n234 585
R201 VTAIL.n228 VTAIL.n227 585
R202 VTAIL.n241 VTAIL.n240 585
R203 VTAIL.n243 VTAIL.n242 585
R204 VTAIL.n224 VTAIL.n223 585
R205 VTAIL.n249 VTAIL.n248 585
R206 VTAIL.n251 VTAIL.n250 585
R207 VTAIL.n220 VTAIL.n219 585
R208 VTAIL.n257 VTAIL.n256 585
R209 VTAIL.n259 VTAIL.n258 585
R210 VTAIL.n216 VTAIL.n215 585
R211 VTAIL.n265 VTAIL.n264 585
R212 VTAIL.n267 VTAIL.n266 585
R213 VTAIL.n212 VTAIL.n211 585
R214 VTAIL.n274 VTAIL.n273 585
R215 VTAIL.n275 VTAIL.n210 585
R216 VTAIL.n277 VTAIL.n276 585
R217 VTAIL.n208 VTAIL.n207 585
R218 VTAIL.n283 VTAIL.n282 585
R219 VTAIL.n285 VTAIL.n284 585
R220 VTAIL.n204 VTAIL.n203 585
R221 VTAIL.n291 VTAIL.n290 585
R222 VTAIL.n293 VTAIL.n292 585
R223 VTAIL.n689 VTAIL.n688 585
R224 VTAIL.n687 VTAIL.n686 585
R225 VTAIL.n600 VTAIL.n599 585
R226 VTAIL.n681 VTAIL.n680 585
R227 VTAIL.n679 VTAIL.n678 585
R228 VTAIL.n604 VTAIL.n603 585
R229 VTAIL.n608 VTAIL.n606 585
R230 VTAIL.n673 VTAIL.n672 585
R231 VTAIL.n671 VTAIL.n670 585
R232 VTAIL.n610 VTAIL.n609 585
R233 VTAIL.n665 VTAIL.n664 585
R234 VTAIL.n663 VTAIL.n662 585
R235 VTAIL.n614 VTAIL.n613 585
R236 VTAIL.n657 VTAIL.n656 585
R237 VTAIL.n655 VTAIL.n654 585
R238 VTAIL.n618 VTAIL.n617 585
R239 VTAIL.n649 VTAIL.n648 585
R240 VTAIL.n647 VTAIL.n646 585
R241 VTAIL.n622 VTAIL.n621 585
R242 VTAIL.n641 VTAIL.n640 585
R243 VTAIL.n639 VTAIL.n638 585
R244 VTAIL.n626 VTAIL.n625 585
R245 VTAIL.n633 VTAIL.n632 585
R246 VTAIL.n631 VTAIL.n630 585
R247 VTAIL.n589 VTAIL.n588 585
R248 VTAIL.n587 VTAIL.n586 585
R249 VTAIL.n500 VTAIL.n499 585
R250 VTAIL.n581 VTAIL.n580 585
R251 VTAIL.n579 VTAIL.n578 585
R252 VTAIL.n504 VTAIL.n503 585
R253 VTAIL.n508 VTAIL.n506 585
R254 VTAIL.n573 VTAIL.n572 585
R255 VTAIL.n571 VTAIL.n570 585
R256 VTAIL.n510 VTAIL.n509 585
R257 VTAIL.n565 VTAIL.n564 585
R258 VTAIL.n563 VTAIL.n562 585
R259 VTAIL.n514 VTAIL.n513 585
R260 VTAIL.n557 VTAIL.n556 585
R261 VTAIL.n555 VTAIL.n554 585
R262 VTAIL.n518 VTAIL.n517 585
R263 VTAIL.n549 VTAIL.n548 585
R264 VTAIL.n547 VTAIL.n546 585
R265 VTAIL.n522 VTAIL.n521 585
R266 VTAIL.n541 VTAIL.n540 585
R267 VTAIL.n539 VTAIL.n538 585
R268 VTAIL.n526 VTAIL.n525 585
R269 VTAIL.n533 VTAIL.n532 585
R270 VTAIL.n531 VTAIL.n530 585
R271 VTAIL.n491 VTAIL.n490 585
R272 VTAIL.n489 VTAIL.n488 585
R273 VTAIL.n402 VTAIL.n401 585
R274 VTAIL.n483 VTAIL.n482 585
R275 VTAIL.n481 VTAIL.n480 585
R276 VTAIL.n406 VTAIL.n405 585
R277 VTAIL.n410 VTAIL.n408 585
R278 VTAIL.n475 VTAIL.n474 585
R279 VTAIL.n473 VTAIL.n472 585
R280 VTAIL.n412 VTAIL.n411 585
R281 VTAIL.n467 VTAIL.n466 585
R282 VTAIL.n465 VTAIL.n464 585
R283 VTAIL.n416 VTAIL.n415 585
R284 VTAIL.n459 VTAIL.n458 585
R285 VTAIL.n457 VTAIL.n456 585
R286 VTAIL.n420 VTAIL.n419 585
R287 VTAIL.n451 VTAIL.n450 585
R288 VTAIL.n449 VTAIL.n448 585
R289 VTAIL.n424 VTAIL.n423 585
R290 VTAIL.n443 VTAIL.n442 585
R291 VTAIL.n441 VTAIL.n440 585
R292 VTAIL.n428 VTAIL.n427 585
R293 VTAIL.n435 VTAIL.n434 585
R294 VTAIL.n433 VTAIL.n432 585
R295 VTAIL.n391 VTAIL.n390 585
R296 VTAIL.n389 VTAIL.n388 585
R297 VTAIL.n302 VTAIL.n301 585
R298 VTAIL.n383 VTAIL.n382 585
R299 VTAIL.n381 VTAIL.n380 585
R300 VTAIL.n306 VTAIL.n305 585
R301 VTAIL.n310 VTAIL.n308 585
R302 VTAIL.n375 VTAIL.n374 585
R303 VTAIL.n373 VTAIL.n372 585
R304 VTAIL.n312 VTAIL.n311 585
R305 VTAIL.n367 VTAIL.n366 585
R306 VTAIL.n365 VTAIL.n364 585
R307 VTAIL.n316 VTAIL.n315 585
R308 VTAIL.n359 VTAIL.n358 585
R309 VTAIL.n357 VTAIL.n356 585
R310 VTAIL.n320 VTAIL.n319 585
R311 VTAIL.n351 VTAIL.n350 585
R312 VTAIL.n349 VTAIL.n348 585
R313 VTAIL.n324 VTAIL.n323 585
R314 VTAIL.n343 VTAIL.n342 585
R315 VTAIL.n341 VTAIL.n340 585
R316 VTAIL.n328 VTAIL.n327 585
R317 VTAIL.n335 VTAIL.n334 585
R318 VTAIL.n333 VTAIL.n332 585
R319 VTAIL.n725 VTAIL.t1 327.466
R320 VTAIL.n33 VTAIL.t7 327.466
R321 VTAIL.n131 VTAIL.t9 327.466
R322 VTAIL.n231 VTAIL.t11 327.466
R323 VTAIL.n629 VTAIL.t10 327.466
R324 VTAIL.n529 VTAIL.t12 327.466
R325 VTAIL.n431 VTAIL.t3 327.466
R326 VTAIL.n331 VTAIL.t4 327.466
R327 VTAIL.n728 VTAIL.n727 171.744
R328 VTAIL.n728 VTAIL.n721 171.744
R329 VTAIL.n735 VTAIL.n721 171.744
R330 VTAIL.n736 VTAIL.n735 171.744
R331 VTAIL.n736 VTAIL.n717 171.744
R332 VTAIL.n743 VTAIL.n717 171.744
R333 VTAIL.n744 VTAIL.n743 171.744
R334 VTAIL.n744 VTAIL.n713 171.744
R335 VTAIL.n751 VTAIL.n713 171.744
R336 VTAIL.n752 VTAIL.n751 171.744
R337 VTAIL.n752 VTAIL.n709 171.744
R338 VTAIL.n759 VTAIL.n709 171.744
R339 VTAIL.n760 VTAIL.n759 171.744
R340 VTAIL.n760 VTAIL.n705 171.744
R341 VTAIL.n768 VTAIL.n705 171.744
R342 VTAIL.n769 VTAIL.n768 171.744
R343 VTAIL.n770 VTAIL.n769 171.744
R344 VTAIL.n770 VTAIL.n701 171.744
R345 VTAIL.n777 VTAIL.n701 171.744
R346 VTAIL.n778 VTAIL.n777 171.744
R347 VTAIL.n778 VTAIL.n697 171.744
R348 VTAIL.n785 VTAIL.n697 171.744
R349 VTAIL.n786 VTAIL.n785 171.744
R350 VTAIL.n36 VTAIL.n35 171.744
R351 VTAIL.n36 VTAIL.n29 171.744
R352 VTAIL.n43 VTAIL.n29 171.744
R353 VTAIL.n44 VTAIL.n43 171.744
R354 VTAIL.n44 VTAIL.n25 171.744
R355 VTAIL.n51 VTAIL.n25 171.744
R356 VTAIL.n52 VTAIL.n51 171.744
R357 VTAIL.n52 VTAIL.n21 171.744
R358 VTAIL.n59 VTAIL.n21 171.744
R359 VTAIL.n60 VTAIL.n59 171.744
R360 VTAIL.n60 VTAIL.n17 171.744
R361 VTAIL.n67 VTAIL.n17 171.744
R362 VTAIL.n68 VTAIL.n67 171.744
R363 VTAIL.n68 VTAIL.n13 171.744
R364 VTAIL.n76 VTAIL.n13 171.744
R365 VTAIL.n77 VTAIL.n76 171.744
R366 VTAIL.n78 VTAIL.n77 171.744
R367 VTAIL.n78 VTAIL.n9 171.744
R368 VTAIL.n85 VTAIL.n9 171.744
R369 VTAIL.n86 VTAIL.n85 171.744
R370 VTAIL.n86 VTAIL.n5 171.744
R371 VTAIL.n93 VTAIL.n5 171.744
R372 VTAIL.n94 VTAIL.n93 171.744
R373 VTAIL.n134 VTAIL.n133 171.744
R374 VTAIL.n134 VTAIL.n127 171.744
R375 VTAIL.n141 VTAIL.n127 171.744
R376 VTAIL.n142 VTAIL.n141 171.744
R377 VTAIL.n142 VTAIL.n123 171.744
R378 VTAIL.n149 VTAIL.n123 171.744
R379 VTAIL.n150 VTAIL.n149 171.744
R380 VTAIL.n150 VTAIL.n119 171.744
R381 VTAIL.n157 VTAIL.n119 171.744
R382 VTAIL.n158 VTAIL.n157 171.744
R383 VTAIL.n158 VTAIL.n115 171.744
R384 VTAIL.n165 VTAIL.n115 171.744
R385 VTAIL.n166 VTAIL.n165 171.744
R386 VTAIL.n166 VTAIL.n111 171.744
R387 VTAIL.n174 VTAIL.n111 171.744
R388 VTAIL.n175 VTAIL.n174 171.744
R389 VTAIL.n176 VTAIL.n175 171.744
R390 VTAIL.n176 VTAIL.n107 171.744
R391 VTAIL.n183 VTAIL.n107 171.744
R392 VTAIL.n184 VTAIL.n183 171.744
R393 VTAIL.n184 VTAIL.n103 171.744
R394 VTAIL.n191 VTAIL.n103 171.744
R395 VTAIL.n192 VTAIL.n191 171.744
R396 VTAIL.n234 VTAIL.n233 171.744
R397 VTAIL.n234 VTAIL.n227 171.744
R398 VTAIL.n241 VTAIL.n227 171.744
R399 VTAIL.n242 VTAIL.n241 171.744
R400 VTAIL.n242 VTAIL.n223 171.744
R401 VTAIL.n249 VTAIL.n223 171.744
R402 VTAIL.n250 VTAIL.n249 171.744
R403 VTAIL.n250 VTAIL.n219 171.744
R404 VTAIL.n257 VTAIL.n219 171.744
R405 VTAIL.n258 VTAIL.n257 171.744
R406 VTAIL.n258 VTAIL.n215 171.744
R407 VTAIL.n265 VTAIL.n215 171.744
R408 VTAIL.n266 VTAIL.n265 171.744
R409 VTAIL.n266 VTAIL.n211 171.744
R410 VTAIL.n274 VTAIL.n211 171.744
R411 VTAIL.n275 VTAIL.n274 171.744
R412 VTAIL.n276 VTAIL.n275 171.744
R413 VTAIL.n276 VTAIL.n207 171.744
R414 VTAIL.n283 VTAIL.n207 171.744
R415 VTAIL.n284 VTAIL.n283 171.744
R416 VTAIL.n284 VTAIL.n203 171.744
R417 VTAIL.n291 VTAIL.n203 171.744
R418 VTAIL.n292 VTAIL.n291 171.744
R419 VTAIL.n688 VTAIL.n687 171.744
R420 VTAIL.n687 VTAIL.n599 171.744
R421 VTAIL.n680 VTAIL.n599 171.744
R422 VTAIL.n680 VTAIL.n679 171.744
R423 VTAIL.n679 VTAIL.n603 171.744
R424 VTAIL.n608 VTAIL.n603 171.744
R425 VTAIL.n672 VTAIL.n608 171.744
R426 VTAIL.n672 VTAIL.n671 171.744
R427 VTAIL.n671 VTAIL.n609 171.744
R428 VTAIL.n664 VTAIL.n609 171.744
R429 VTAIL.n664 VTAIL.n663 171.744
R430 VTAIL.n663 VTAIL.n613 171.744
R431 VTAIL.n656 VTAIL.n613 171.744
R432 VTAIL.n656 VTAIL.n655 171.744
R433 VTAIL.n655 VTAIL.n617 171.744
R434 VTAIL.n648 VTAIL.n617 171.744
R435 VTAIL.n648 VTAIL.n647 171.744
R436 VTAIL.n647 VTAIL.n621 171.744
R437 VTAIL.n640 VTAIL.n621 171.744
R438 VTAIL.n640 VTAIL.n639 171.744
R439 VTAIL.n639 VTAIL.n625 171.744
R440 VTAIL.n632 VTAIL.n625 171.744
R441 VTAIL.n632 VTAIL.n631 171.744
R442 VTAIL.n588 VTAIL.n587 171.744
R443 VTAIL.n587 VTAIL.n499 171.744
R444 VTAIL.n580 VTAIL.n499 171.744
R445 VTAIL.n580 VTAIL.n579 171.744
R446 VTAIL.n579 VTAIL.n503 171.744
R447 VTAIL.n508 VTAIL.n503 171.744
R448 VTAIL.n572 VTAIL.n508 171.744
R449 VTAIL.n572 VTAIL.n571 171.744
R450 VTAIL.n571 VTAIL.n509 171.744
R451 VTAIL.n564 VTAIL.n509 171.744
R452 VTAIL.n564 VTAIL.n563 171.744
R453 VTAIL.n563 VTAIL.n513 171.744
R454 VTAIL.n556 VTAIL.n513 171.744
R455 VTAIL.n556 VTAIL.n555 171.744
R456 VTAIL.n555 VTAIL.n517 171.744
R457 VTAIL.n548 VTAIL.n517 171.744
R458 VTAIL.n548 VTAIL.n547 171.744
R459 VTAIL.n547 VTAIL.n521 171.744
R460 VTAIL.n540 VTAIL.n521 171.744
R461 VTAIL.n540 VTAIL.n539 171.744
R462 VTAIL.n539 VTAIL.n525 171.744
R463 VTAIL.n532 VTAIL.n525 171.744
R464 VTAIL.n532 VTAIL.n531 171.744
R465 VTAIL.n490 VTAIL.n489 171.744
R466 VTAIL.n489 VTAIL.n401 171.744
R467 VTAIL.n482 VTAIL.n401 171.744
R468 VTAIL.n482 VTAIL.n481 171.744
R469 VTAIL.n481 VTAIL.n405 171.744
R470 VTAIL.n410 VTAIL.n405 171.744
R471 VTAIL.n474 VTAIL.n410 171.744
R472 VTAIL.n474 VTAIL.n473 171.744
R473 VTAIL.n473 VTAIL.n411 171.744
R474 VTAIL.n466 VTAIL.n411 171.744
R475 VTAIL.n466 VTAIL.n465 171.744
R476 VTAIL.n465 VTAIL.n415 171.744
R477 VTAIL.n458 VTAIL.n415 171.744
R478 VTAIL.n458 VTAIL.n457 171.744
R479 VTAIL.n457 VTAIL.n419 171.744
R480 VTAIL.n450 VTAIL.n419 171.744
R481 VTAIL.n450 VTAIL.n449 171.744
R482 VTAIL.n449 VTAIL.n423 171.744
R483 VTAIL.n442 VTAIL.n423 171.744
R484 VTAIL.n442 VTAIL.n441 171.744
R485 VTAIL.n441 VTAIL.n427 171.744
R486 VTAIL.n434 VTAIL.n427 171.744
R487 VTAIL.n434 VTAIL.n433 171.744
R488 VTAIL.n390 VTAIL.n389 171.744
R489 VTAIL.n389 VTAIL.n301 171.744
R490 VTAIL.n382 VTAIL.n301 171.744
R491 VTAIL.n382 VTAIL.n381 171.744
R492 VTAIL.n381 VTAIL.n305 171.744
R493 VTAIL.n310 VTAIL.n305 171.744
R494 VTAIL.n374 VTAIL.n310 171.744
R495 VTAIL.n374 VTAIL.n373 171.744
R496 VTAIL.n373 VTAIL.n311 171.744
R497 VTAIL.n366 VTAIL.n311 171.744
R498 VTAIL.n366 VTAIL.n365 171.744
R499 VTAIL.n365 VTAIL.n315 171.744
R500 VTAIL.n358 VTAIL.n315 171.744
R501 VTAIL.n358 VTAIL.n357 171.744
R502 VTAIL.n357 VTAIL.n319 171.744
R503 VTAIL.n350 VTAIL.n319 171.744
R504 VTAIL.n350 VTAIL.n349 171.744
R505 VTAIL.n349 VTAIL.n323 171.744
R506 VTAIL.n342 VTAIL.n323 171.744
R507 VTAIL.n342 VTAIL.n341 171.744
R508 VTAIL.n341 VTAIL.n327 171.744
R509 VTAIL.n334 VTAIL.n327 171.744
R510 VTAIL.n334 VTAIL.n333 171.744
R511 VTAIL.n727 VTAIL.t1 85.8723
R512 VTAIL.n35 VTAIL.t7 85.8723
R513 VTAIL.n133 VTAIL.t9 85.8723
R514 VTAIL.n233 VTAIL.t11 85.8723
R515 VTAIL.n631 VTAIL.t10 85.8723
R516 VTAIL.n531 VTAIL.t12 85.8723
R517 VTAIL.n433 VTAIL.t3 85.8723
R518 VTAIL.n333 VTAIL.t4 85.8723
R519 VTAIL.n595 VTAIL.n594 52.3434
R520 VTAIL.n397 VTAIL.n396 52.3434
R521 VTAIL.n1 VTAIL.n0 52.3433
R522 VTAIL.n199 VTAIL.n198 52.3433
R523 VTAIL.n791 VTAIL.n790 32.1853
R524 VTAIL.n99 VTAIL.n98 32.1853
R525 VTAIL.n197 VTAIL.n196 32.1853
R526 VTAIL.n297 VTAIL.n296 32.1853
R527 VTAIL.n693 VTAIL.n692 32.1853
R528 VTAIL.n593 VTAIL.n592 32.1853
R529 VTAIL.n495 VTAIL.n494 32.1853
R530 VTAIL.n395 VTAIL.n394 32.1853
R531 VTAIL.n791 VTAIL.n693 29.9014
R532 VTAIL.n395 VTAIL.n297 29.9014
R533 VTAIL.n726 VTAIL.n725 16.3895
R534 VTAIL.n34 VTAIL.n33 16.3895
R535 VTAIL.n132 VTAIL.n131 16.3895
R536 VTAIL.n232 VTAIL.n231 16.3895
R537 VTAIL.n630 VTAIL.n629 16.3895
R538 VTAIL.n530 VTAIL.n529 16.3895
R539 VTAIL.n432 VTAIL.n431 16.3895
R540 VTAIL.n332 VTAIL.n331 16.3895
R541 VTAIL.n771 VTAIL.n702 13.1884
R542 VTAIL.n79 VTAIL.n10 13.1884
R543 VTAIL.n177 VTAIL.n108 13.1884
R544 VTAIL.n277 VTAIL.n208 13.1884
R545 VTAIL.n606 VTAIL.n604 13.1884
R546 VTAIL.n506 VTAIL.n504 13.1884
R547 VTAIL.n408 VTAIL.n406 13.1884
R548 VTAIL.n308 VTAIL.n306 13.1884
R549 VTAIL.n729 VTAIL.n724 12.8005
R550 VTAIL.n772 VTAIL.n704 12.8005
R551 VTAIL.n776 VTAIL.n775 12.8005
R552 VTAIL.n37 VTAIL.n32 12.8005
R553 VTAIL.n80 VTAIL.n12 12.8005
R554 VTAIL.n84 VTAIL.n83 12.8005
R555 VTAIL.n135 VTAIL.n130 12.8005
R556 VTAIL.n178 VTAIL.n110 12.8005
R557 VTAIL.n182 VTAIL.n181 12.8005
R558 VTAIL.n235 VTAIL.n230 12.8005
R559 VTAIL.n278 VTAIL.n210 12.8005
R560 VTAIL.n282 VTAIL.n281 12.8005
R561 VTAIL.n678 VTAIL.n677 12.8005
R562 VTAIL.n674 VTAIL.n673 12.8005
R563 VTAIL.n633 VTAIL.n628 12.8005
R564 VTAIL.n578 VTAIL.n577 12.8005
R565 VTAIL.n574 VTAIL.n573 12.8005
R566 VTAIL.n533 VTAIL.n528 12.8005
R567 VTAIL.n480 VTAIL.n479 12.8005
R568 VTAIL.n476 VTAIL.n475 12.8005
R569 VTAIL.n435 VTAIL.n430 12.8005
R570 VTAIL.n380 VTAIL.n379 12.8005
R571 VTAIL.n376 VTAIL.n375 12.8005
R572 VTAIL.n335 VTAIL.n330 12.8005
R573 VTAIL.n730 VTAIL.n722 12.0247
R574 VTAIL.n767 VTAIL.n766 12.0247
R575 VTAIL.n779 VTAIL.n700 12.0247
R576 VTAIL.n38 VTAIL.n30 12.0247
R577 VTAIL.n75 VTAIL.n74 12.0247
R578 VTAIL.n87 VTAIL.n8 12.0247
R579 VTAIL.n136 VTAIL.n128 12.0247
R580 VTAIL.n173 VTAIL.n172 12.0247
R581 VTAIL.n185 VTAIL.n106 12.0247
R582 VTAIL.n236 VTAIL.n228 12.0247
R583 VTAIL.n273 VTAIL.n272 12.0247
R584 VTAIL.n285 VTAIL.n206 12.0247
R585 VTAIL.n681 VTAIL.n602 12.0247
R586 VTAIL.n670 VTAIL.n607 12.0247
R587 VTAIL.n634 VTAIL.n626 12.0247
R588 VTAIL.n581 VTAIL.n502 12.0247
R589 VTAIL.n570 VTAIL.n507 12.0247
R590 VTAIL.n534 VTAIL.n526 12.0247
R591 VTAIL.n483 VTAIL.n404 12.0247
R592 VTAIL.n472 VTAIL.n409 12.0247
R593 VTAIL.n436 VTAIL.n428 12.0247
R594 VTAIL.n383 VTAIL.n304 12.0247
R595 VTAIL.n372 VTAIL.n309 12.0247
R596 VTAIL.n336 VTAIL.n328 12.0247
R597 VTAIL.n734 VTAIL.n733 11.249
R598 VTAIL.n765 VTAIL.n706 11.249
R599 VTAIL.n780 VTAIL.n698 11.249
R600 VTAIL.n42 VTAIL.n41 11.249
R601 VTAIL.n73 VTAIL.n14 11.249
R602 VTAIL.n88 VTAIL.n6 11.249
R603 VTAIL.n140 VTAIL.n139 11.249
R604 VTAIL.n171 VTAIL.n112 11.249
R605 VTAIL.n186 VTAIL.n104 11.249
R606 VTAIL.n240 VTAIL.n239 11.249
R607 VTAIL.n271 VTAIL.n212 11.249
R608 VTAIL.n286 VTAIL.n204 11.249
R609 VTAIL.n682 VTAIL.n600 11.249
R610 VTAIL.n669 VTAIL.n610 11.249
R611 VTAIL.n638 VTAIL.n637 11.249
R612 VTAIL.n582 VTAIL.n500 11.249
R613 VTAIL.n569 VTAIL.n510 11.249
R614 VTAIL.n538 VTAIL.n537 11.249
R615 VTAIL.n484 VTAIL.n402 11.249
R616 VTAIL.n471 VTAIL.n412 11.249
R617 VTAIL.n440 VTAIL.n439 11.249
R618 VTAIL.n384 VTAIL.n302 11.249
R619 VTAIL.n371 VTAIL.n312 11.249
R620 VTAIL.n340 VTAIL.n339 11.249
R621 VTAIL.n737 VTAIL.n720 10.4732
R622 VTAIL.n762 VTAIL.n761 10.4732
R623 VTAIL.n784 VTAIL.n783 10.4732
R624 VTAIL.n45 VTAIL.n28 10.4732
R625 VTAIL.n70 VTAIL.n69 10.4732
R626 VTAIL.n92 VTAIL.n91 10.4732
R627 VTAIL.n143 VTAIL.n126 10.4732
R628 VTAIL.n168 VTAIL.n167 10.4732
R629 VTAIL.n190 VTAIL.n189 10.4732
R630 VTAIL.n243 VTAIL.n226 10.4732
R631 VTAIL.n268 VTAIL.n267 10.4732
R632 VTAIL.n290 VTAIL.n289 10.4732
R633 VTAIL.n686 VTAIL.n685 10.4732
R634 VTAIL.n666 VTAIL.n665 10.4732
R635 VTAIL.n641 VTAIL.n624 10.4732
R636 VTAIL.n586 VTAIL.n585 10.4732
R637 VTAIL.n566 VTAIL.n565 10.4732
R638 VTAIL.n541 VTAIL.n524 10.4732
R639 VTAIL.n488 VTAIL.n487 10.4732
R640 VTAIL.n468 VTAIL.n467 10.4732
R641 VTAIL.n443 VTAIL.n426 10.4732
R642 VTAIL.n388 VTAIL.n387 10.4732
R643 VTAIL.n368 VTAIL.n367 10.4732
R644 VTAIL.n343 VTAIL.n326 10.4732
R645 VTAIL.n738 VTAIL.n718 9.69747
R646 VTAIL.n758 VTAIL.n708 9.69747
R647 VTAIL.n787 VTAIL.n696 9.69747
R648 VTAIL.n46 VTAIL.n26 9.69747
R649 VTAIL.n66 VTAIL.n16 9.69747
R650 VTAIL.n95 VTAIL.n4 9.69747
R651 VTAIL.n144 VTAIL.n124 9.69747
R652 VTAIL.n164 VTAIL.n114 9.69747
R653 VTAIL.n193 VTAIL.n102 9.69747
R654 VTAIL.n244 VTAIL.n224 9.69747
R655 VTAIL.n264 VTAIL.n214 9.69747
R656 VTAIL.n293 VTAIL.n202 9.69747
R657 VTAIL.n689 VTAIL.n598 9.69747
R658 VTAIL.n662 VTAIL.n612 9.69747
R659 VTAIL.n642 VTAIL.n622 9.69747
R660 VTAIL.n589 VTAIL.n498 9.69747
R661 VTAIL.n562 VTAIL.n512 9.69747
R662 VTAIL.n542 VTAIL.n522 9.69747
R663 VTAIL.n491 VTAIL.n400 9.69747
R664 VTAIL.n464 VTAIL.n414 9.69747
R665 VTAIL.n444 VTAIL.n424 9.69747
R666 VTAIL.n391 VTAIL.n300 9.69747
R667 VTAIL.n364 VTAIL.n314 9.69747
R668 VTAIL.n344 VTAIL.n324 9.69747
R669 VTAIL.n790 VTAIL.n789 9.45567
R670 VTAIL.n98 VTAIL.n97 9.45567
R671 VTAIL.n196 VTAIL.n195 9.45567
R672 VTAIL.n296 VTAIL.n295 9.45567
R673 VTAIL.n692 VTAIL.n691 9.45567
R674 VTAIL.n592 VTAIL.n591 9.45567
R675 VTAIL.n494 VTAIL.n493 9.45567
R676 VTAIL.n394 VTAIL.n393 9.45567
R677 VTAIL.n789 VTAIL.n788 9.3005
R678 VTAIL.n696 VTAIL.n695 9.3005
R679 VTAIL.n783 VTAIL.n782 9.3005
R680 VTAIL.n781 VTAIL.n780 9.3005
R681 VTAIL.n700 VTAIL.n699 9.3005
R682 VTAIL.n775 VTAIL.n774 9.3005
R683 VTAIL.n747 VTAIL.n746 9.3005
R684 VTAIL.n716 VTAIL.n715 9.3005
R685 VTAIL.n741 VTAIL.n740 9.3005
R686 VTAIL.n739 VTAIL.n738 9.3005
R687 VTAIL.n720 VTAIL.n719 9.3005
R688 VTAIL.n733 VTAIL.n732 9.3005
R689 VTAIL.n731 VTAIL.n730 9.3005
R690 VTAIL.n724 VTAIL.n723 9.3005
R691 VTAIL.n749 VTAIL.n748 9.3005
R692 VTAIL.n712 VTAIL.n711 9.3005
R693 VTAIL.n755 VTAIL.n754 9.3005
R694 VTAIL.n757 VTAIL.n756 9.3005
R695 VTAIL.n708 VTAIL.n707 9.3005
R696 VTAIL.n763 VTAIL.n762 9.3005
R697 VTAIL.n765 VTAIL.n764 9.3005
R698 VTAIL.n766 VTAIL.n703 9.3005
R699 VTAIL.n773 VTAIL.n772 9.3005
R700 VTAIL.n97 VTAIL.n96 9.3005
R701 VTAIL.n4 VTAIL.n3 9.3005
R702 VTAIL.n91 VTAIL.n90 9.3005
R703 VTAIL.n89 VTAIL.n88 9.3005
R704 VTAIL.n8 VTAIL.n7 9.3005
R705 VTAIL.n83 VTAIL.n82 9.3005
R706 VTAIL.n55 VTAIL.n54 9.3005
R707 VTAIL.n24 VTAIL.n23 9.3005
R708 VTAIL.n49 VTAIL.n48 9.3005
R709 VTAIL.n47 VTAIL.n46 9.3005
R710 VTAIL.n28 VTAIL.n27 9.3005
R711 VTAIL.n41 VTAIL.n40 9.3005
R712 VTAIL.n39 VTAIL.n38 9.3005
R713 VTAIL.n32 VTAIL.n31 9.3005
R714 VTAIL.n57 VTAIL.n56 9.3005
R715 VTAIL.n20 VTAIL.n19 9.3005
R716 VTAIL.n63 VTAIL.n62 9.3005
R717 VTAIL.n65 VTAIL.n64 9.3005
R718 VTAIL.n16 VTAIL.n15 9.3005
R719 VTAIL.n71 VTAIL.n70 9.3005
R720 VTAIL.n73 VTAIL.n72 9.3005
R721 VTAIL.n74 VTAIL.n11 9.3005
R722 VTAIL.n81 VTAIL.n80 9.3005
R723 VTAIL.n195 VTAIL.n194 9.3005
R724 VTAIL.n102 VTAIL.n101 9.3005
R725 VTAIL.n189 VTAIL.n188 9.3005
R726 VTAIL.n187 VTAIL.n186 9.3005
R727 VTAIL.n106 VTAIL.n105 9.3005
R728 VTAIL.n181 VTAIL.n180 9.3005
R729 VTAIL.n153 VTAIL.n152 9.3005
R730 VTAIL.n122 VTAIL.n121 9.3005
R731 VTAIL.n147 VTAIL.n146 9.3005
R732 VTAIL.n145 VTAIL.n144 9.3005
R733 VTAIL.n126 VTAIL.n125 9.3005
R734 VTAIL.n139 VTAIL.n138 9.3005
R735 VTAIL.n137 VTAIL.n136 9.3005
R736 VTAIL.n130 VTAIL.n129 9.3005
R737 VTAIL.n155 VTAIL.n154 9.3005
R738 VTAIL.n118 VTAIL.n117 9.3005
R739 VTAIL.n161 VTAIL.n160 9.3005
R740 VTAIL.n163 VTAIL.n162 9.3005
R741 VTAIL.n114 VTAIL.n113 9.3005
R742 VTAIL.n169 VTAIL.n168 9.3005
R743 VTAIL.n171 VTAIL.n170 9.3005
R744 VTAIL.n172 VTAIL.n109 9.3005
R745 VTAIL.n179 VTAIL.n178 9.3005
R746 VTAIL.n295 VTAIL.n294 9.3005
R747 VTAIL.n202 VTAIL.n201 9.3005
R748 VTAIL.n289 VTAIL.n288 9.3005
R749 VTAIL.n287 VTAIL.n286 9.3005
R750 VTAIL.n206 VTAIL.n205 9.3005
R751 VTAIL.n281 VTAIL.n280 9.3005
R752 VTAIL.n253 VTAIL.n252 9.3005
R753 VTAIL.n222 VTAIL.n221 9.3005
R754 VTAIL.n247 VTAIL.n246 9.3005
R755 VTAIL.n245 VTAIL.n244 9.3005
R756 VTAIL.n226 VTAIL.n225 9.3005
R757 VTAIL.n239 VTAIL.n238 9.3005
R758 VTAIL.n237 VTAIL.n236 9.3005
R759 VTAIL.n230 VTAIL.n229 9.3005
R760 VTAIL.n255 VTAIL.n254 9.3005
R761 VTAIL.n218 VTAIL.n217 9.3005
R762 VTAIL.n261 VTAIL.n260 9.3005
R763 VTAIL.n263 VTAIL.n262 9.3005
R764 VTAIL.n214 VTAIL.n213 9.3005
R765 VTAIL.n269 VTAIL.n268 9.3005
R766 VTAIL.n271 VTAIL.n270 9.3005
R767 VTAIL.n272 VTAIL.n209 9.3005
R768 VTAIL.n279 VTAIL.n278 9.3005
R769 VTAIL.n616 VTAIL.n615 9.3005
R770 VTAIL.n659 VTAIL.n658 9.3005
R771 VTAIL.n661 VTAIL.n660 9.3005
R772 VTAIL.n612 VTAIL.n611 9.3005
R773 VTAIL.n667 VTAIL.n666 9.3005
R774 VTAIL.n669 VTAIL.n668 9.3005
R775 VTAIL.n607 VTAIL.n605 9.3005
R776 VTAIL.n675 VTAIL.n674 9.3005
R777 VTAIL.n691 VTAIL.n690 9.3005
R778 VTAIL.n598 VTAIL.n597 9.3005
R779 VTAIL.n685 VTAIL.n684 9.3005
R780 VTAIL.n683 VTAIL.n682 9.3005
R781 VTAIL.n602 VTAIL.n601 9.3005
R782 VTAIL.n677 VTAIL.n676 9.3005
R783 VTAIL.n653 VTAIL.n652 9.3005
R784 VTAIL.n651 VTAIL.n650 9.3005
R785 VTAIL.n620 VTAIL.n619 9.3005
R786 VTAIL.n645 VTAIL.n644 9.3005
R787 VTAIL.n643 VTAIL.n642 9.3005
R788 VTAIL.n624 VTAIL.n623 9.3005
R789 VTAIL.n637 VTAIL.n636 9.3005
R790 VTAIL.n635 VTAIL.n634 9.3005
R791 VTAIL.n628 VTAIL.n627 9.3005
R792 VTAIL.n516 VTAIL.n515 9.3005
R793 VTAIL.n559 VTAIL.n558 9.3005
R794 VTAIL.n561 VTAIL.n560 9.3005
R795 VTAIL.n512 VTAIL.n511 9.3005
R796 VTAIL.n567 VTAIL.n566 9.3005
R797 VTAIL.n569 VTAIL.n568 9.3005
R798 VTAIL.n507 VTAIL.n505 9.3005
R799 VTAIL.n575 VTAIL.n574 9.3005
R800 VTAIL.n591 VTAIL.n590 9.3005
R801 VTAIL.n498 VTAIL.n497 9.3005
R802 VTAIL.n585 VTAIL.n584 9.3005
R803 VTAIL.n583 VTAIL.n582 9.3005
R804 VTAIL.n502 VTAIL.n501 9.3005
R805 VTAIL.n577 VTAIL.n576 9.3005
R806 VTAIL.n553 VTAIL.n552 9.3005
R807 VTAIL.n551 VTAIL.n550 9.3005
R808 VTAIL.n520 VTAIL.n519 9.3005
R809 VTAIL.n545 VTAIL.n544 9.3005
R810 VTAIL.n543 VTAIL.n542 9.3005
R811 VTAIL.n524 VTAIL.n523 9.3005
R812 VTAIL.n537 VTAIL.n536 9.3005
R813 VTAIL.n535 VTAIL.n534 9.3005
R814 VTAIL.n528 VTAIL.n527 9.3005
R815 VTAIL.n418 VTAIL.n417 9.3005
R816 VTAIL.n461 VTAIL.n460 9.3005
R817 VTAIL.n463 VTAIL.n462 9.3005
R818 VTAIL.n414 VTAIL.n413 9.3005
R819 VTAIL.n469 VTAIL.n468 9.3005
R820 VTAIL.n471 VTAIL.n470 9.3005
R821 VTAIL.n409 VTAIL.n407 9.3005
R822 VTAIL.n477 VTAIL.n476 9.3005
R823 VTAIL.n493 VTAIL.n492 9.3005
R824 VTAIL.n400 VTAIL.n399 9.3005
R825 VTAIL.n487 VTAIL.n486 9.3005
R826 VTAIL.n485 VTAIL.n484 9.3005
R827 VTAIL.n404 VTAIL.n403 9.3005
R828 VTAIL.n479 VTAIL.n478 9.3005
R829 VTAIL.n455 VTAIL.n454 9.3005
R830 VTAIL.n453 VTAIL.n452 9.3005
R831 VTAIL.n422 VTAIL.n421 9.3005
R832 VTAIL.n447 VTAIL.n446 9.3005
R833 VTAIL.n445 VTAIL.n444 9.3005
R834 VTAIL.n426 VTAIL.n425 9.3005
R835 VTAIL.n439 VTAIL.n438 9.3005
R836 VTAIL.n437 VTAIL.n436 9.3005
R837 VTAIL.n430 VTAIL.n429 9.3005
R838 VTAIL.n318 VTAIL.n317 9.3005
R839 VTAIL.n361 VTAIL.n360 9.3005
R840 VTAIL.n363 VTAIL.n362 9.3005
R841 VTAIL.n314 VTAIL.n313 9.3005
R842 VTAIL.n369 VTAIL.n368 9.3005
R843 VTAIL.n371 VTAIL.n370 9.3005
R844 VTAIL.n309 VTAIL.n307 9.3005
R845 VTAIL.n377 VTAIL.n376 9.3005
R846 VTAIL.n393 VTAIL.n392 9.3005
R847 VTAIL.n300 VTAIL.n299 9.3005
R848 VTAIL.n387 VTAIL.n386 9.3005
R849 VTAIL.n385 VTAIL.n384 9.3005
R850 VTAIL.n304 VTAIL.n303 9.3005
R851 VTAIL.n379 VTAIL.n378 9.3005
R852 VTAIL.n355 VTAIL.n354 9.3005
R853 VTAIL.n353 VTAIL.n352 9.3005
R854 VTAIL.n322 VTAIL.n321 9.3005
R855 VTAIL.n347 VTAIL.n346 9.3005
R856 VTAIL.n345 VTAIL.n344 9.3005
R857 VTAIL.n326 VTAIL.n325 9.3005
R858 VTAIL.n339 VTAIL.n338 9.3005
R859 VTAIL.n337 VTAIL.n336 9.3005
R860 VTAIL.n330 VTAIL.n329 9.3005
R861 VTAIL.n742 VTAIL.n741 8.92171
R862 VTAIL.n757 VTAIL.n710 8.92171
R863 VTAIL.n788 VTAIL.n694 8.92171
R864 VTAIL.n50 VTAIL.n49 8.92171
R865 VTAIL.n65 VTAIL.n18 8.92171
R866 VTAIL.n96 VTAIL.n2 8.92171
R867 VTAIL.n148 VTAIL.n147 8.92171
R868 VTAIL.n163 VTAIL.n116 8.92171
R869 VTAIL.n194 VTAIL.n100 8.92171
R870 VTAIL.n248 VTAIL.n247 8.92171
R871 VTAIL.n263 VTAIL.n216 8.92171
R872 VTAIL.n294 VTAIL.n200 8.92171
R873 VTAIL.n690 VTAIL.n596 8.92171
R874 VTAIL.n661 VTAIL.n614 8.92171
R875 VTAIL.n646 VTAIL.n645 8.92171
R876 VTAIL.n590 VTAIL.n496 8.92171
R877 VTAIL.n561 VTAIL.n514 8.92171
R878 VTAIL.n546 VTAIL.n545 8.92171
R879 VTAIL.n492 VTAIL.n398 8.92171
R880 VTAIL.n463 VTAIL.n416 8.92171
R881 VTAIL.n448 VTAIL.n447 8.92171
R882 VTAIL.n392 VTAIL.n298 8.92171
R883 VTAIL.n363 VTAIL.n316 8.92171
R884 VTAIL.n348 VTAIL.n347 8.92171
R885 VTAIL.n745 VTAIL.n716 8.14595
R886 VTAIL.n754 VTAIL.n753 8.14595
R887 VTAIL.n53 VTAIL.n24 8.14595
R888 VTAIL.n62 VTAIL.n61 8.14595
R889 VTAIL.n151 VTAIL.n122 8.14595
R890 VTAIL.n160 VTAIL.n159 8.14595
R891 VTAIL.n251 VTAIL.n222 8.14595
R892 VTAIL.n260 VTAIL.n259 8.14595
R893 VTAIL.n658 VTAIL.n657 8.14595
R894 VTAIL.n649 VTAIL.n620 8.14595
R895 VTAIL.n558 VTAIL.n557 8.14595
R896 VTAIL.n549 VTAIL.n520 8.14595
R897 VTAIL.n460 VTAIL.n459 8.14595
R898 VTAIL.n451 VTAIL.n422 8.14595
R899 VTAIL.n360 VTAIL.n359 8.14595
R900 VTAIL.n351 VTAIL.n322 8.14595
R901 VTAIL.n746 VTAIL.n714 7.3702
R902 VTAIL.n750 VTAIL.n712 7.3702
R903 VTAIL.n54 VTAIL.n22 7.3702
R904 VTAIL.n58 VTAIL.n20 7.3702
R905 VTAIL.n152 VTAIL.n120 7.3702
R906 VTAIL.n156 VTAIL.n118 7.3702
R907 VTAIL.n252 VTAIL.n220 7.3702
R908 VTAIL.n256 VTAIL.n218 7.3702
R909 VTAIL.n654 VTAIL.n616 7.3702
R910 VTAIL.n650 VTAIL.n618 7.3702
R911 VTAIL.n554 VTAIL.n516 7.3702
R912 VTAIL.n550 VTAIL.n518 7.3702
R913 VTAIL.n456 VTAIL.n418 7.3702
R914 VTAIL.n452 VTAIL.n420 7.3702
R915 VTAIL.n356 VTAIL.n318 7.3702
R916 VTAIL.n352 VTAIL.n320 7.3702
R917 VTAIL.n749 VTAIL.n714 6.59444
R918 VTAIL.n750 VTAIL.n749 6.59444
R919 VTAIL.n57 VTAIL.n22 6.59444
R920 VTAIL.n58 VTAIL.n57 6.59444
R921 VTAIL.n155 VTAIL.n120 6.59444
R922 VTAIL.n156 VTAIL.n155 6.59444
R923 VTAIL.n255 VTAIL.n220 6.59444
R924 VTAIL.n256 VTAIL.n255 6.59444
R925 VTAIL.n654 VTAIL.n653 6.59444
R926 VTAIL.n653 VTAIL.n618 6.59444
R927 VTAIL.n554 VTAIL.n553 6.59444
R928 VTAIL.n553 VTAIL.n518 6.59444
R929 VTAIL.n456 VTAIL.n455 6.59444
R930 VTAIL.n455 VTAIL.n420 6.59444
R931 VTAIL.n356 VTAIL.n355 6.59444
R932 VTAIL.n355 VTAIL.n320 6.59444
R933 VTAIL.n746 VTAIL.n745 5.81868
R934 VTAIL.n753 VTAIL.n712 5.81868
R935 VTAIL.n54 VTAIL.n53 5.81868
R936 VTAIL.n61 VTAIL.n20 5.81868
R937 VTAIL.n152 VTAIL.n151 5.81868
R938 VTAIL.n159 VTAIL.n118 5.81868
R939 VTAIL.n252 VTAIL.n251 5.81868
R940 VTAIL.n259 VTAIL.n218 5.81868
R941 VTAIL.n657 VTAIL.n616 5.81868
R942 VTAIL.n650 VTAIL.n649 5.81868
R943 VTAIL.n557 VTAIL.n516 5.81868
R944 VTAIL.n550 VTAIL.n549 5.81868
R945 VTAIL.n459 VTAIL.n418 5.81868
R946 VTAIL.n452 VTAIL.n451 5.81868
R947 VTAIL.n359 VTAIL.n318 5.81868
R948 VTAIL.n352 VTAIL.n351 5.81868
R949 VTAIL.n742 VTAIL.n716 5.04292
R950 VTAIL.n754 VTAIL.n710 5.04292
R951 VTAIL.n790 VTAIL.n694 5.04292
R952 VTAIL.n50 VTAIL.n24 5.04292
R953 VTAIL.n62 VTAIL.n18 5.04292
R954 VTAIL.n98 VTAIL.n2 5.04292
R955 VTAIL.n148 VTAIL.n122 5.04292
R956 VTAIL.n160 VTAIL.n116 5.04292
R957 VTAIL.n196 VTAIL.n100 5.04292
R958 VTAIL.n248 VTAIL.n222 5.04292
R959 VTAIL.n260 VTAIL.n216 5.04292
R960 VTAIL.n296 VTAIL.n200 5.04292
R961 VTAIL.n692 VTAIL.n596 5.04292
R962 VTAIL.n658 VTAIL.n614 5.04292
R963 VTAIL.n646 VTAIL.n620 5.04292
R964 VTAIL.n592 VTAIL.n496 5.04292
R965 VTAIL.n558 VTAIL.n514 5.04292
R966 VTAIL.n546 VTAIL.n520 5.04292
R967 VTAIL.n494 VTAIL.n398 5.04292
R968 VTAIL.n460 VTAIL.n416 5.04292
R969 VTAIL.n448 VTAIL.n422 5.04292
R970 VTAIL.n394 VTAIL.n298 5.04292
R971 VTAIL.n360 VTAIL.n316 5.04292
R972 VTAIL.n348 VTAIL.n322 5.04292
R973 VTAIL.n741 VTAIL.n718 4.26717
R974 VTAIL.n758 VTAIL.n757 4.26717
R975 VTAIL.n788 VTAIL.n787 4.26717
R976 VTAIL.n49 VTAIL.n26 4.26717
R977 VTAIL.n66 VTAIL.n65 4.26717
R978 VTAIL.n96 VTAIL.n95 4.26717
R979 VTAIL.n147 VTAIL.n124 4.26717
R980 VTAIL.n164 VTAIL.n163 4.26717
R981 VTAIL.n194 VTAIL.n193 4.26717
R982 VTAIL.n247 VTAIL.n224 4.26717
R983 VTAIL.n264 VTAIL.n263 4.26717
R984 VTAIL.n294 VTAIL.n293 4.26717
R985 VTAIL.n690 VTAIL.n689 4.26717
R986 VTAIL.n662 VTAIL.n661 4.26717
R987 VTAIL.n645 VTAIL.n622 4.26717
R988 VTAIL.n590 VTAIL.n589 4.26717
R989 VTAIL.n562 VTAIL.n561 4.26717
R990 VTAIL.n545 VTAIL.n522 4.26717
R991 VTAIL.n492 VTAIL.n491 4.26717
R992 VTAIL.n464 VTAIL.n463 4.26717
R993 VTAIL.n447 VTAIL.n424 4.26717
R994 VTAIL.n392 VTAIL.n391 4.26717
R995 VTAIL.n364 VTAIL.n363 4.26717
R996 VTAIL.n347 VTAIL.n324 4.26717
R997 VTAIL.n725 VTAIL.n723 3.70982
R998 VTAIL.n33 VTAIL.n31 3.70982
R999 VTAIL.n131 VTAIL.n129 3.70982
R1000 VTAIL.n231 VTAIL.n229 3.70982
R1001 VTAIL.n629 VTAIL.n627 3.70982
R1002 VTAIL.n529 VTAIL.n527 3.70982
R1003 VTAIL.n431 VTAIL.n429 3.70982
R1004 VTAIL.n331 VTAIL.n329 3.70982
R1005 VTAIL.n738 VTAIL.n737 3.49141
R1006 VTAIL.n761 VTAIL.n708 3.49141
R1007 VTAIL.n784 VTAIL.n696 3.49141
R1008 VTAIL.n46 VTAIL.n45 3.49141
R1009 VTAIL.n69 VTAIL.n16 3.49141
R1010 VTAIL.n92 VTAIL.n4 3.49141
R1011 VTAIL.n144 VTAIL.n143 3.49141
R1012 VTAIL.n167 VTAIL.n114 3.49141
R1013 VTAIL.n190 VTAIL.n102 3.49141
R1014 VTAIL.n244 VTAIL.n243 3.49141
R1015 VTAIL.n267 VTAIL.n214 3.49141
R1016 VTAIL.n290 VTAIL.n202 3.49141
R1017 VTAIL.n686 VTAIL.n598 3.49141
R1018 VTAIL.n665 VTAIL.n612 3.49141
R1019 VTAIL.n642 VTAIL.n641 3.49141
R1020 VTAIL.n586 VTAIL.n498 3.49141
R1021 VTAIL.n565 VTAIL.n512 3.49141
R1022 VTAIL.n542 VTAIL.n541 3.49141
R1023 VTAIL.n488 VTAIL.n400 3.49141
R1024 VTAIL.n467 VTAIL.n414 3.49141
R1025 VTAIL.n444 VTAIL.n443 3.49141
R1026 VTAIL.n388 VTAIL.n300 3.49141
R1027 VTAIL.n367 VTAIL.n314 3.49141
R1028 VTAIL.n344 VTAIL.n343 3.49141
R1029 VTAIL.n734 VTAIL.n720 2.71565
R1030 VTAIL.n762 VTAIL.n706 2.71565
R1031 VTAIL.n783 VTAIL.n698 2.71565
R1032 VTAIL.n42 VTAIL.n28 2.71565
R1033 VTAIL.n70 VTAIL.n14 2.71565
R1034 VTAIL.n91 VTAIL.n6 2.71565
R1035 VTAIL.n140 VTAIL.n126 2.71565
R1036 VTAIL.n168 VTAIL.n112 2.71565
R1037 VTAIL.n189 VTAIL.n104 2.71565
R1038 VTAIL.n240 VTAIL.n226 2.71565
R1039 VTAIL.n268 VTAIL.n212 2.71565
R1040 VTAIL.n289 VTAIL.n204 2.71565
R1041 VTAIL.n685 VTAIL.n600 2.71565
R1042 VTAIL.n666 VTAIL.n610 2.71565
R1043 VTAIL.n638 VTAIL.n624 2.71565
R1044 VTAIL.n585 VTAIL.n500 2.71565
R1045 VTAIL.n566 VTAIL.n510 2.71565
R1046 VTAIL.n538 VTAIL.n524 2.71565
R1047 VTAIL.n487 VTAIL.n402 2.71565
R1048 VTAIL.n468 VTAIL.n412 2.71565
R1049 VTAIL.n440 VTAIL.n426 2.71565
R1050 VTAIL.n387 VTAIL.n302 2.71565
R1051 VTAIL.n368 VTAIL.n312 2.71565
R1052 VTAIL.n340 VTAIL.n326 2.71565
R1053 VTAIL.n397 VTAIL.n395 2.43153
R1054 VTAIL.n495 VTAIL.n397 2.43153
R1055 VTAIL.n595 VTAIL.n593 2.43153
R1056 VTAIL.n693 VTAIL.n595 2.43153
R1057 VTAIL.n297 VTAIL.n199 2.43153
R1058 VTAIL.n199 VTAIL.n197 2.43153
R1059 VTAIL.n99 VTAIL.n1 2.43153
R1060 VTAIL VTAIL.n791 2.37334
R1061 VTAIL.n733 VTAIL.n722 1.93989
R1062 VTAIL.n767 VTAIL.n765 1.93989
R1063 VTAIL.n780 VTAIL.n779 1.93989
R1064 VTAIL.n41 VTAIL.n30 1.93989
R1065 VTAIL.n75 VTAIL.n73 1.93989
R1066 VTAIL.n88 VTAIL.n87 1.93989
R1067 VTAIL.n139 VTAIL.n128 1.93989
R1068 VTAIL.n173 VTAIL.n171 1.93989
R1069 VTAIL.n186 VTAIL.n185 1.93989
R1070 VTAIL.n239 VTAIL.n228 1.93989
R1071 VTAIL.n273 VTAIL.n271 1.93989
R1072 VTAIL.n286 VTAIL.n285 1.93989
R1073 VTAIL.n682 VTAIL.n681 1.93989
R1074 VTAIL.n670 VTAIL.n669 1.93989
R1075 VTAIL.n637 VTAIL.n626 1.93989
R1076 VTAIL.n582 VTAIL.n581 1.93989
R1077 VTAIL.n570 VTAIL.n569 1.93989
R1078 VTAIL.n537 VTAIL.n526 1.93989
R1079 VTAIL.n484 VTAIL.n483 1.93989
R1080 VTAIL.n472 VTAIL.n471 1.93989
R1081 VTAIL.n439 VTAIL.n428 1.93989
R1082 VTAIL.n384 VTAIL.n383 1.93989
R1083 VTAIL.n372 VTAIL.n371 1.93989
R1084 VTAIL.n339 VTAIL.n328 1.93989
R1085 VTAIL.n0 VTAIL.t6 1.85581
R1086 VTAIL.n0 VTAIL.t0 1.85581
R1087 VTAIL.n198 VTAIL.t13 1.85581
R1088 VTAIL.n198 VTAIL.t8 1.85581
R1089 VTAIL.n594 VTAIL.t14 1.85581
R1090 VTAIL.n594 VTAIL.t15 1.85581
R1091 VTAIL.n396 VTAIL.t2 1.85581
R1092 VTAIL.n396 VTAIL.t5 1.85581
R1093 VTAIL.n730 VTAIL.n729 1.16414
R1094 VTAIL.n766 VTAIL.n704 1.16414
R1095 VTAIL.n776 VTAIL.n700 1.16414
R1096 VTAIL.n38 VTAIL.n37 1.16414
R1097 VTAIL.n74 VTAIL.n12 1.16414
R1098 VTAIL.n84 VTAIL.n8 1.16414
R1099 VTAIL.n136 VTAIL.n135 1.16414
R1100 VTAIL.n172 VTAIL.n110 1.16414
R1101 VTAIL.n182 VTAIL.n106 1.16414
R1102 VTAIL.n236 VTAIL.n235 1.16414
R1103 VTAIL.n272 VTAIL.n210 1.16414
R1104 VTAIL.n282 VTAIL.n206 1.16414
R1105 VTAIL.n678 VTAIL.n602 1.16414
R1106 VTAIL.n673 VTAIL.n607 1.16414
R1107 VTAIL.n634 VTAIL.n633 1.16414
R1108 VTAIL.n578 VTAIL.n502 1.16414
R1109 VTAIL.n573 VTAIL.n507 1.16414
R1110 VTAIL.n534 VTAIL.n533 1.16414
R1111 VTAIL.n480 VTAIL.n404 1.16414
R1112 VTAIL.n475 VTAIL.n409 1.16414
R1113 VTAIL.n436 VTAIL.n435 1.16414
R1114 VTAIL.n380 VTAIL.n304 1.16414
R1115 VTAIL.n375 VTAIL.n309 1.16414
R1116 VTAIL.n336 VTAIL.n335 1.16414
R1117 VTAIL.n593 VTAIL.n495 0.470328
R1118 VTAIL.n197 VTAIL.n99 0.470328
R1119 VTAIL.n726 VTAIL.n724 0.388379
R1120 VTAIL.n772 VTAIL.n771 0.388379
R1121 VTAIL.n775 VTAIL.n702 0.388379
R1122 VTAIL.n34 VTAIL.n32 0.388379
R1123 VTAIL.n80 VTAIL.n79 0.388379
R1124 VTAIL.n83 VTAIL.n10 0.388379
R1125 VTAIL.n132 VTAIL.n130 0.388379
R1126 VTAIL.n178 VTAIL.n177 0.388379
R1127 VTAIL.n181 VTAIL.n108 0.388379
R1128 VTAIL.n232 VTAIL.n230 0.388379
R1129 VTAIL.n278 VTAIL.n277 0.388379
R1130 VTAIL.n281 VTAIL.n208 0.388379
R1131 VTAIL.n677 VTAIL.n604 0.388379
R1132 VTAIL.n674 VTAIL.n606 0.388379
R1133 VTAIL.n630 VTAIL.n628 0.388379
R1134 VTAIL.n577 VTAIL.n504 0.388379
R1135 VTAIL.n574 VTAIL.n506 0.388379
R1136 VTAIL.n530 VTAIL.n528 0.388379
R1137 VTAIL.n479 VTAIL.n406 0.388379
R1138 VTAIL.n476 VTAIL.n408 0.388379
R1139 VTAIL.n432 VTAIL.n430 0.388379
R1140 VTAIL.n379 VTAIL.n306 0.388379
R1141 VTAIL.n376 VTAIL.n308 0.388379
R1142 VTAIL.n332 VTAIL.n330 0.388379
R1143 VTAIL.n731 VTAIL.n723 0.155672
R1144 VTAIL.n732 VTAIL.n731 0.155672
R1145 VTAIL.n732 VTAIL.n719 0.155672
R1146 VTAIL.n739 VTAIL.n719 0.155672
R1147 VTAIL.n740 VTAIL.n739 0.155672
R1148 VTAIL.n740 VTAIL.n715 0.155672
R1149 VTAIL.n747 VTAIL.n715 0.155672
R1150 VTAIL.n748 VTAIL.n747 0.155672
R1151 VTAIL.n748 VTAIL.n711 0.155672
R1152 VTAIL.n755 VTAIL.n711 0.155672
R1153 VTAIL.n756 VTAIL.n755 0.155672
R1154 VTAIL.n756 VTAIL.n707 0.155672
R1155 VTAIL.n763 VTAIL.n707 0.155672
R1156 VTAIL.n764 VTAIL.n763 0.155672
R1157 VTAIL.n764 VTAIL.n703 0.155672
R1158 VTAIL.n773 VTAIL.n703 0.155672
R1159 VTAIL.n774 VTAIL.n773 0.155672
R1160 VTAIL.n774 VTAIL.n699 0.155672
R1161 VTAIL.n781 VTAIL.n699 0.155672
R1162 VTAIL.n782 VTAIL.n781 0.155672
R1163 VTAIL.n782 VTAIL.n695 0.155672
R1164 VTAIL.n789 VTAIL.n695 0.155672
R1165 VTAIL.n39 VTAIL.n31 0.155672
R1166 VTAIL.n40 VTAIL.n39 0.155672
R1167 VTAIL.n40 VTAIL.n27 0.155672
R1168 VTAIL.n47 VTAIL.n27 0.155672
R1169 VTAIL.n48 VTAIL.n47 0.155672
R1170 VTAIL.n48 VTAIL.n23 0.155672
R1171 VTAIL.n55 VTAIL.n23 0.155672
R1172 VTAIL.n56 VTAIL.n55 0.155672
R1173 VTAIL.n56 VTAIL.n19 0.155672
R1174 VTAIL.n63 VTAIL.n19 0.155672
R1175 VTAIL.n64 VTAIL.n63 0.155672
R1176 VTAIL.n64 VTAIL.n15 0.155672
R1177 VTAIL.n71 VTAIL.n15 0.155672
R1178 VTAIL.n72 VTAIL.n71 0.155672
R1179 VTAIL.n72 VTAIL.n11 0.155672
R1180 VTAIL.n81 VTAIL.n11 0.155672
R1181 VTAIL.n82 VTAIL.n81 0.155672
R1182 VTAIL.n82 VTAIL.n7 0.155672
R1183 VTAIL.n89 VTAIL.n7 0.155672
R1184 VTAIL.n90 VTAIL.n89 0.155672
R1185 VTAIL.n90 VTAIL.n3 0.155672
R1186 VTAIL.n97 VTAIL.n3 0.155672
R1187 VTAIL.n137 VTAIL.n129 0.155672
R1188 VTAIL.n138 VTAIL.n137 0.155672
R1189 VTAIL.n138 VTAIL.n125 0.155672
R1190 VTAIL.n145 VTAIL.n125 0.155672
R1191 VTAIL.n146 VTAIL.n145 0.155672
R1192 VTAIL.n146 VTAIL.n121 0.155672
R1193 VTAIL.n153 VTAIL.n121 0.155672
R1194 VTAIL.n154 VTAIL.n153 0.155672
R1195 VTAIL.n154 VTAIL.n117 0.155672
R1196 VTAIL.n161 VTAIL.n117 0.155672
R1197 VTAIL.n162 VTAIL.n161 0.155672
R1198 VTAIL.n162 VTAIL.n113 0.155672
R1199 VTAIL.n169 VTAIL.n113 0.155672
R1200 VTAIL.n170 VTAIL.n169 0.155672
R1201 VTAIL.n170 VTAIL.n109 0.155672
R1202 VTAIL.n179 VTAIL.n109 0.155672
R1203 VTAIL.n180 VTAIL.n179 0.155672
R1204 VTAIL.n180 VTAIL.n105 0.155672
R1205 VTAIL.n187 VTAIL.n105 0.155672
R1206 VTAIL.n188 VTAIL.n187 0.155672
R1207 VTAIL.n188 VTAIL.n101 0.155672
R1208 VTAIL.n195 VTAIL.n101 0.155672
R1209 VTAIL.n237 VTAIL.n229 0.155672
R1210 VTAIL.n238 VTAIL.n237 0.155672
R1211 VTAIL.n238 VTAIL.n225 0.155672
R1212 VTAIL.n245 VTAIL.n225 0.155672
R1213 VTAIL.n246 VTAIL.n245 0.155672
R1214 VTAIL.n246 VTAIL.n221 0.155672
R1215 VTAIL.n253 VTAIL.n221 0.155672
R1216 VTAIL.n254 VTAIL.n253 0.155672
R1217 VTAIL.n254 VTAIL.n217 0.155672
R1218 VTAIL.n261 VTAIL.n217 0.155672
R1219 VTAIL.n262 VTAIL.n261 0.155672
R1220 VTAIL.n262 VTAIL.n213 0.155672
R1221 VTAIL.n269 VTAIL.n213 0.155672
R1222 VTAIL.n270 VTAIL.n269 0.155672
R1223 VTAIL.n270 VTAIL.n209 0.155672
R1224 VTAIL.n279 VTAIL.n209 0.155672
R1225 VTAIL.n280 VTAIL.n279 0.155672
R1226 VTAIL.n280 VTAIL.n205 0.155672
R1227 VTAIL.n287 VTAIL.n205 0.155672
R1228 VTAIL.n288 VTAIL.n287 0.155672
R1229 VTAIL.n288 VTAIL.n201 0.155672
R1230 VTAIL.n295 VTAIL.n201 0.155672
R1231 VTAIL.n691 VTAIL.n597 0.155672
R1232 VTAIL.n684 VTAIL.n597 0.155672
R1233 VTAIL.n684 VTAIL.n683 0.155672
R1234 VTAIL.n683 VTAIL.n601 0.155672
R1235 VTAIL.n676 VTAIL.n601 0.155672
R1236 VTAIL.n676 VTAIL.n675 0.155672
R1237 VTAIL.n675 VTAIL.n605 0.155672
R1238 VTAIL.n668 VTAIL.n605 0.155672
R1239 VTAIL.n668 VTAIL.n667 0.155672
R1240 VTAIL.n667 VTAIL.n611 0.155672
R1241 VTAIL.n660 VTAIL.n611 0.155672
R1242 VTAIL.n660 VTAIL.n659 0.155672
R1243 VTAIL.n659 VTAIL.n615 0.155672
R1244 VTAIL.n652 VTAIL.n615 0.155672
R1245 VTAIL.n652 VTAIL.n651 0.155672
R1246 VTAIL.n651 VTAIL.n619 0.155672
R1247 VTAIL.n644 VTAIL.n619 0.155672
R1248 VTAIL.n644 VTAIL.n643 0.155672
R1249 VTAIL.n643 VTAIL.n623 0.155672
R1250 VTAIL.n636 VTAIL.n623 0.155672
R1251 VTAIL.n636 VTAIL.n635 0.155672
R1252 VTAIL.n635 VTAIL.n627 0.155672
R1253 VTAIL.n591 VTAIL.n497 0.155672
R1254 VTAIL.n584 VTAIL.n497 0.155672
R1255 VTAIL.n584 VTAIL.n583 0.155672
R1256 VTAIL.n583 VTAIL.n501 0.155672
R1257 VTAIL.n576 VTAIL.n501 0.155672
R1258 VTAIL.n576 VTAIL.n575 0.155672
R1259 VTAIL.n575 VTAIL.n505 0.155672
R1260 VTAIL.n568 VTAIL.n505 0.155672
R1261 VTAIL.n568 VTAIL.n567 0.155672
R1262 VTAIL.n567 VTAIL.n511 0.155672
R1263 VTAIL.n560 VTAIL.n511 0.155672
R1264 VTAIL.n560 VTAIL.n559 0.155672
R1265 VTAIL.n559 VTAIL.n515 0.155672
R1266 VTAIL.n552 VTAIL.n515 0.155672
R1267 VTAIL.n552 VTAIL.n551 0.155672
R1268 VTAIL.n551 VTAIL.n519 0.155672
R1269 VTAIL.n544 VTAIL.n519 0.155672
R1270 VTAIL.n544 VTAIL.n543 0.155672
R1271 VTAIL.n543 VTAIL.n523 0.155672
R1272 VTAIL.n536 VTAIL.n523 0.155672
R1273 VTAIL.n536 VTAIL.n535 0.155672
R1274 VTAIL.n535 VTAIL.n527 0.155672
R1275 VTAIL.n493 VTAIL.n399 0.155672
R1276 VTAIL.n486 VTAIL.n399 0.155672
R1277 VTAIL.n486 VTAIL.n485 0.155672
R1278 VTAIL.n485 VTAIL.n403 0.155672
R1279 VTAIL.n478 VTAIL.n403 0.155672
R1280 VTAIL.n478 VTAIL.n477 0.155672
R1281 VTAIL.n477 VTAIL.n407 0.155672
R1282 VTAIL.n470 VTAIL.n407 0.155672
R1283 VTAIL.n470 VTAIL.n469 0.155672
R1284 VTAIL.n469 VTAIL.n413 0.155672
R1285 VTAIL.n462 VTAIL.n413 0.155672
R1286 VTAIL.n462 VTAIL.n461 0.155672
R1287 VTAIL.n461 VTAIL.n417 0.155672
R1288 VTAIL.n454 VTAIL.n417 0.155672
R1289 VTAIL.n454 VTAIL.n453 0.155672
R1290 VTAIL.n453 VTAIL.n421 0.155672
R1291 VTAIL.n446 VTAIL.n421 0.155672
R1292 VTAIL.n446 VTAIL.n445 0.155672
R1293 VTAIL.n445 VTAIL.n425 0.155672
R1294 VTAIL.n438 VTAIL.n425 0.155672
R1295 VTAIL.n438 VTAIL.n437 0.155672
R1296 VTAIL.n437 VTAIL.n429 0.155672
R1297 VTAIL.n393 VTAIL.n299 0.155672
R1298 VTAIL.n386 VTAIL.n299 0.155672
R1299 VTAIL.n386 VTAIL.n385 0.155672
R1300 VTAIL.n385 VTAIL.n303 0.155672
R1301 VTAIL.n378 VTAIL.n303 0.155672
R1302 VTAIL.n378 VTAIL.n377 0.155672
R1303 VTAIL.n377 VTAIL.n307 0.155672
R1304 VTAIL.n370 VTAIL.n307 0.155672
R1305 VTAIL.n370 VTAIL.n369 0.155672
R1306 VTAIL.n369 VTAIL.n313 0.155672
R1307 VTAIL.n362 VTAIL.n313 0.155672
R1308 VTAIL.n362 VTAIL.n361 0.155672
R1309 VTAIL.n361 VTAIL.n317 0.155672
R1310 VTAIL.n354 VTAIL.n317 0.155672
R1311 VTAIL.n354 VTAIL.n353 0.155672
R1312 VTAIL.n353 VTAIL.n321 0.155672
R1313 VTAIL.n346 VTAIL.n321 0.155672
R1314 VTAIL.n346 VTAIL.n345 0.155672
R1315 VTAIL.n345 VTAIL.n325 0.155672
R1316 VTAIL.n338 VTAIL.n325 0.155672
R1317 VTAIL.n338 VTAIL.n337 0.155672
R1318 VTAIL.n337 VTAIL.n329 0.155672
R1319 VTAIL VTAIL.n1 0.0586897
R1320 VN.n6 VN.t7 203.607
R1321 VN.n33 VN.t6 203.607
R1322 VN.n7 VN.t5 169.571
R1323 VN.n3 VN.t3 169.571
R1324 VN.n25 VN.t2 169.571
R1325 VN.n34 VN.t4 169.571
R1326 VN.n30 VN.t1 169.571
R1327 VN.n52 VN.t0 169.571
R1328 VN.n51 VN.n27 161.3
R1329 VN.n50 VN.n49 161.3
R1330 VN.n48 VN.n28 161.3
R1331 VN.n47 VN.n46 161.3
R1332 VN.n45 VN.n29 161.3
R1333 VN.n44 VN.n43 161.3
R1334 VN.n42 VN.n41 161.3
R1335 VN.n40 VN.n31 161.3
R1336 VN.n39 VN.n38 161.3
R1337 VN.n37 VN.n32 161.3
R1338 VN.n36 VN.n35 161.3
R1339 VN.n24 VN.n0 161.3
R1340 VN.n23 VN.n22 161.3
R1341 VN.n21 VN.n1 161.3
R1342 VN.n20 VN.n19 161.3
R1343 VN.n18 VN.n2 161.3
R1344 VN.n17 VN.n16 161.3
R1345 VN.n15 VN.n14 161.3
R1346 VN.n13 VN.n4 161.3
R1347 VN.n12 VN.n11 161.3
R1348 VN.n10 VN.n5 161.3
R1349 VN.n9 VN.n8 161.3
R1350 VN.n26 VN.n25 99.596
R1351 VN.n53 VN.n52 99.596
R1352 VN.n19 VN.n1 56.5617
R1353 VN.n46 VN.n28 56.5617
R1354 VN VN.n53 54.8542
R1355 VN.n7 VN.n6 52.5962
R1356 VN.n34 VN.n33 52.5962
R1357 VN.n12 VN.n5 40.577
R1358 VN.n13 VN.n12 40.577
R1359 VN.n39 VN.n32 40.577
R1360 VN.n40 VN.n39 40.577
R1361 VN.n8 VN.n5 24.5923
R1362 VN.n14 VN.n13 24.5923
R1363 VN.n18 VN.n17 24.5923
R1364 VN.n19 VN.n18 24.5923
R1365 VN.n23 VN.n1 24.5923
R1366 VN.n24 VN.n23 24.5923
R1367 VN.n35 VN.n32 24.5923
R1368 VN.n46 VN.n45 24.5923
R1369 VN.n45 VN.n44 24.5923
R1370 VN.n41 VN.n40 24.5923
R1371 VN.n51 VN.n50 24.5923
R1372 VN.n50 VN.n28 24.5923
R1373 VN.n8 VN.n7 20.1658
R1374 VN.n14 VN.n3 20.1658
R1375 VN.n35 VN.n34 20.1658
R1376 VN.n41 VN.n30 20.1658
R1377 VN.n25 VN.n24 11.3127
R1378 VN.n52 VN.n51 11.3127
R1379 VN.n36 VN.n33 6.75133
R1380 VN.n9 VN.n6 6.75133
R1381 VN.n17 VN.n3 4.42703
R1382 VN.n44 VN.n30 4.42703
R1383 VN.n53 VN.n27 0.278335
R1384 VN.n26 VN.n0 0.278335
R1385 VN.n49 VN.n27 0.189894
R1386 VN.n49 VN.n48 0.189894
R1387 VN.n48 VN.n47 0.189894
R1388 VN.n47 VN.n29 0.189894
R1389 VN.n43 VN.n29 0.189894
R1390 VN.n43 VN.n42 0.189894
R1391 VN.n42 VN.n31 0.189894
R1392 VN.n38 VN.n31 0.189894
R1393 VN.n38 VN.n37 0.189894
R1394 VN.n37 VN.n36 0.189894
R1395 VN.n10 VN.n9 0.189894
R1396 VN.n11 VN.n10 0.189894
R1397 VN.n11 VN.n4 0.189894
R1398 VN.n15 VN.n4 0.189894
R1399 VN.n16 VN.n15 0.189894
R1400 VN.n16 VN.n2 0.189894
R1401 VN.n20 VN.n2 0.189894
R1402 VN.n21 VN.n20 0.189894
R1403 VN.n22 VN.n21 0.189894
R1404 VN.n22 VN.n0 0.189894
R1405 VN VN.n26 0.153485
R1406 VDD2.n2 VDD2.n1 70.1822
R1407 VDD2.n2 VDD2.n0 70.1822
R1408 VDD2 VDD2.n5 70.1794
R1409 VDD2.n4 VDD2.n3 69.0222
R1410 VDD2.n4 VDD2.n2 49.7584
R1411 VDD2.n5 VDD2.t3 1.85581
R1412 VDD2.n5 VDD2.t1 1.85581
R1413 VDD2.n3 VDD2.t7 1.85581
R1414 VDD2.n3 VDD2.t6 1.85581
R1415 VDD2.n1 VDD2.t4 1.85581
R1416 VDD2.n1 VDD2.t5 1.85581
R1417 VDD2.n0 VDD2.t0 1.85581
R1418 VDD2.n0 VDD2.t2 1.85581
R1419 VDD2 VDD2.n4 1.27421
R1420 B.n495 B.n494 585
R1421 B.n493 B.n144 585
R1422 B.n492 B.n491 585
R1423 B.n490 B.n145 585
R1424 B.n489 B.n488 585
R1425 B.n487 B.n146 585
R1426 B.n486 B.n485 585
R1427 B.n484 B.n147 585
R1428 B.n483 B.n482 585
R1429 B.n481 B.n148 585
R1430 B.n480 B.n479 585
R1431 B.n478 B.n149 585
R1432 B.n477 B.n476 585
R1433 B.n475 B.n150 585
R1434 B.n474 B.n473 585
R1435 B.n472 B.n151 585
R1436 B.n471 B.n470 585
R1437 B.n469 B.n152 585
R1438 B.n468 B.n467 585
R1439 B.n466 B.n153 585
R1440 B.n465 B.n464 585
R1441 B.n463 B.n154 585
R1442 B.n462 B.n461 585
R1443 B.n460 B.n155 585
R1444 B.n459 B.n458 585
R1445 B.n457 B.n156 585
R1446 B.n456 B.n455 585
R1447 B.n454 B.n157 585
R1448 B.n453 B.n452 585
R1449 B.n451 B.n158 585
R1450 B.n450 B.n449 585
R1451 B.n448 B.n159 585
R1452 B.n447 B.n446 585
R1453 B.n445 B.n160 585
R1454 B.n444 B.n443 585
R1455 B.n442 B.n161 585
R1456 B.n441 B.n440 585
R1457 B.n439 B.n162 585
R1458 B.n438 B.n437 585
R1459 B.n436 B.n163 585
R1460 B.n435 B.n434 585
R1461 B.n433 B.n164 585
R1462 B.n432 B.n431 585
R1463 B.n430 B.n165 585
R1464 B.n429 B.n428 585
R1465 B.n427 B.n166 585
R1466 B.n426 B.n425 585
R1467 B.n424 B.n167 585
R1468 B.n423 B.n422 585
R1469 B.n421 B.n168 585
R1470 B.n420 B.n419 585
R1471 B.n418 B.n169 585
R1472 B.n417 B.n416 585
R1473 B.n415 B.n170 585
R1474 B.n414 B.n413 585
R1475 B.n412 B.n171 585
R1476 B.n411 B.n410 585
R1477 B.n409 B.n172 585
R1478 B.n408 B.n407 585
R1479 B.n403 B.n173 585
R1480 B.n402 B.n401 585
R1481 B.n400 B.n174 585
R1482 B.n399 B.n398 585
R1483 B.n397 B.n175 585
R1484 B.n396 B.n395 585
R1485 B.n394 B.n176 585
R1486 B.n393 B.n392 585
R1487 B.n390 B.n177 585
R1488 B.n389 B.n388 585
R1489 B.n387 B.n180 585
R1490 B.n386 B.n385 585
R1491 B.n384 B.n181 585
R1492 B.n383 B.n382 585
R1493 B.n381 B.n182 585
R1494 B.n380 B.n379 585
R1495 B.n378 B.n183 585
R1496 B.n377 B.n376 585
R1497 B.n375 B.n184 585
R1498 B.n374 B.n373 585
R1499 B.n372 B.n185 585
R1500 B.n371 B.n370 585
R1501 B.n369 B.n186 585
R1502 B.n368 B.n367 585
R1503 B.n366 B.n187 585
R1504 B.n365 B.n364 585
R1505 B.n363 B.n188 585
R1506 B.n362 B.n361 585
R1507 B.n360 B.n189 585
R1508 B.n359 B.n358 585
R1509 B.n357 B.n190 585
R1510 B.n356 B.n355 585
R1511 B.n354 B.n191 585
R1512 B.n353 B.n352 585
R1513 B.n351 B.n192 585
R1514 B.n350 B.n349 585
R1515 B.n348 B.n193 585
R1516 B.n347 B.n346 585
R1517 B.n345 B.n194 585
R1518 B.n344 B.n343 585
R1519 B.n342 B.n195 585
R1520 B.n341 B.n340 585
R1521 B.n339 B.n196 585
R1522 B.n338 B.n337 585
R1523 B.n336 B.n197 585
R1524 B.n335 B.n334 585
R1525 B.n333 B.n198 585
R1526 B.n332 B.n331 585
R1527 B.n330 B.n199 585
R1528 B.n329 B.n328 585
R1529 B.n327 B.n200 585
R1530 B.n326 B.n325 585
R1531 B.n324 B.n201 585
R1532 B.n323 B.n322 585
R1533 B.n321 B.n202 585
R1534 B.n320 B.n319 585
R1535 B.n318 B.n203 585
R1536 B.n317 B.n316 585
R1537 B.n315 B.n204 585
R1538 B.n314 B.n313 585
R1539 B.n312 B.n205 585
R1540 B.n311 B.n310 585
R1541 B.n309 B.n206 585
R1542 B.n308 B.n307 585
R1543 B.n306 B.n207 585
R1544 B.n305 B.n304 585
R1545 B.n496 B.n143 585
R1546 B.n498 B.n497 585
R1547 B.n499 B.n142 585
R1548 B.n501 B.n500 585
R1549 B.n502 B.n141 585
R1550 B.n504 B.n503 585
R1551 B.n505 B.n140 585
R1552 B.n507 B.n506 585
R1553 B.n508 B.n139 585
R1554 B.n510 B.n509 585
R1555 B.n511 B.n138 585
R1556 B.n513 B.n512 585
R1557 B.n514 B.n137 585
R1558 B.n516 B.n515 585
R1559 B.n517 B.n136 585
R1560 B.n519 B.n518 585
R1561 B.n520 B.n135 585
R1562 B.n522 B.n521 585
R1563 B.n523 B.n134 585
R1564 B.n525 B.n524 585
R1565 B.n526 B.n133 585
R1566 B.n528 B.n527 585
R1567 B.n529 B.n132 585
R1568 B.n531 B.n530 585
R1569 B.n532 B.n131 585
R1570 B.n534 B.n533 585
R1571 B.n535 B.n130 585
R1572 B.n537 B.n536 585
R1573 B.n538 B.n129 585
R1574 B.n540 B.n539 585
R1575 B.n541 B.n128 585
R1576 B.n543 B.n542 585
R1577 B.n544 B.n127 585
R1578 B.n546 B.n545 585
R1579 B.n547 B.n126 585
R1580 B.n549 B.n548 585
R1581 B.n550 B.n125 585
R1582 B.n552 B.n551 585
R1583 B.n553 B.n124 585
R1584 B.n555 B.n554 585
R1585 B.n556 B.n123 585
R1586 B.n558 B.n557 585
R1587 B.n559 B.n122 585
R1588 B.n561 B.n560 585
R1589 B.n562 B.n121 585
R1590 B.n564 B.n563 585
R1591 B.n565 B.n120 585
R1592 B.n567 B.n566 585
R1593 B.n568 B.n119 585
R1594 B.n570 B.n569 585
R1595 B.n571 B.n118 585
R1596 B.n573 B.n572 585
R1597 B.n574 B.n117 585
R1598 B.n576 B.n575 585
R1599 B.n577 B.n116 585
R1600 B.n579 B.n578 585
R1601 B.n580 B.n115 585
R1602 B.n582 B.n581 585
R1603 B.n583 B.n114 585
R1604 B.n585 B.n584 585
R1605 B.n586 B.n113 585
R1606 B.n588 B.n587 585
R1607 B.n589 B.n112 585
R1608 B.n591 B.n590 585
R1609 B.n592 B.n111 585
R1610 B.n594 B.n593 585
R1611 B.n595 B.n110 585
R1612 B.n597 B.n596 585
R1613 B.n598 B.n109 585
R1614 B.n600 B.n599 585
R1615 B.n601 B.n108 585
R1616 B.n603 B.n602 585
R1617 B.n604 B.n107 585
R1618 B.n606 B.n605 585
R1619 B.n607 B.n106 585
R1620 B.n609 B.n608 585
R1621 B.n610 B.n105 585
R1622 B.n612 B.n611 585
R1623 B.n613 B.n104 585
R1624 B.n615 B.n614 585
R1625 B.n616 B.n103 585
R1626 B.n618 B.n617 585
R1627 B.n619 B.n102 585
R1628 B.n621 B.n620 585
R1629 B.n622 B.n101 585
R1630 B.n624 B.n623 585
R1631 B.n625 B.n100 585
R1632 B.n627 B.n626 585
R1633 B.n628 B.n99 585
R1634 B.n630 B.n629 585
R1635 B.n631 B.n98 585
R1636 B.n633 B.n632 585
R1637 B.n634 B.n97 585
R1638 B.n636 B.n635 585
R1639 B.n637 B.n96 585
R1640 B.n639 B.n638 585
R1641 B.n640 B.n95 585
R1642 B.n642 B.n641 585
R1643 B.n643 B.n94 585
R1644 B.n645 B.n644 585
R1645 B.n834 B.n833 585
R1646 B.n832 B.n27 585
R1647 B.n831 B.n830 585
R1648 B.n829 B.n28 585
R1649 B.n828 B.n827 585
R1650 B.n826 B.n29 585
R1651 B.n825 B.n824 585
R1652 B.n823 B.n30 585
R1653 B.n822 B.n821 585
R1654 B.n820 B.n31 585
R1655 B.n819 B.n818 585
R1656 B.n817 B.n32 585
R1657 B.n816 B.n815 585
R1658 B.n814 B.n33 585
R1659 B.n813 B.n812 585
R1660 B.n811 B.n34 585
R1661 B.n810 B.n809 585
R1662 B.n808 B.n35 585
R1663 B.n807 B.n806 585
R1664 B.n805 B.n36 585
R1665 B.n804 B.n803 585
R1666 B.n802 B.n37 585
R1667 B.n801 B.n800 585
R1668 B.n799 B.n38 585
R1669 B.n798 B.n797 585
R1670 B.n796 B.n39 585
R1671 B.n795 B.n794 585
R1672 B.n793 B.n40 585
R1673 B.n792 B.n791 585
R1674 B.n790 B.n41 585
R1675 B.n789 B.n788 585
R1676 B.n787 B.n42 585
R1677 B.n786 B.n785 585
R1678 B.n784 B.n43 585
R1679 B.n783 B.n782 585
R1680 B.n781 B.n44 585
R1681 B.n780 B.n779 585
R1682 B.n778 B.n45 585
R1683 B.n777 B.n776 585
R1684 B.n775 B.n46 585
R1685 B.n774 B.n773 585
R1686 B.n772 B.n47 585
R1687 B.n771 B.n770 585
R1688 B.n769 B.n48 585
R1689 B.n768 B.n767 585
R1690 B.n766 B.n49 585
R1691 B.n765 B.n764 585
R1692 B.n763 B.n50 585
R1693 B.n762 B.n761 585
R1694 B.n760 B.n51 585
R1695 B.n759 B.n758 585
R1696 B.n757 B.n52 585
R1697 B.n756 B.n755 585
R1698 B.n754 B.n53 585
R1699 B.n753 B.n752 585
R1700 B.n751 B.n54 585
R1701 B.n750 B.n749 585
R1702 B.n748 B.n55 585
R1703 B.n746 B.n745 585
R1704 B.n744 B.n58 585
R1705 B.n743 B.n742 585
R1706 B.n741 B.n59 585
R1707 B.n740 B.n739 585
R1708 B.n738 B.n60 585
R1709 B.n737 B.n736 585
R1710 B.n735 B.n61 585
R1711 B.n734 B.n733 585
R1712 B.n732 B.n731 585
R1713 B.n730 B.n65 585
R1714 B.n729 B.n728 585
R1715 B.n727 B.n66 585
R1716 B.n726 B.n725 585
R1717 B.n724 B.n67 585
R1718 B.n723 B.n722 585
R1719 B.n721 B.n68 585
R1720 B.n720 B.n719 585
R1721 B.n718 B.n69 585
R1722 B.n717 B.n716 585
R1723 B.n715 B.n70 585
R1724 B.n714 B.n713 585
R1725 B.n712 B.n71 585
R1726 B.n711 B.n710 585
R1727 B.n709 B.n72 585
R1728 B.n708 B.n707 585
R1729 B.n706 B.n73 585
R1730 B.n705 B.n704 585
R1731 B.n703 B.n74 585
R1732 B.n702 B.n701 585
R1733 B.n700 B.n75 585
R1734 B.n699 B.n698 585
R1735 B.n697 B.n76 585
R1736 B.n696 B.n695 585
R1737 B.n694 B.n77 585
R1738 B.n693 B.n692 585
R1739 B.n691 B.n78 585
R1740 B.n690 B.n689 585
R1741 B.n688 B.n79 585
R1742 B.n687 B.n686 585
R1743 B.n685 B.n80 585
R1744 B.n684 B.n683 585
R1745 B.n682 B.n81 585
R1746 B.n681 B.n680 585
R1747 B.n679 B.n82 585
R1748 B.n678 B.n677 585
R1749 B.n676 B.n83 585
R1750 B.n675 B.n674 585
R1751 B.n673 B.n84 585
R1752 B.n672 B.n671 585
R1753 B.n670 B.n85 585
R1754 B.n669 B.n668 585
R1755 B.n667 B.n86 585
R1756 B.n666 B.n665 585
R1757 B.n664 B.n87 585
R1758 B.n663 B.n662 585
R1759 B.n661 B.n88 585
R1760 B.n660 B.n659 585
R1761 B.n658 B.n89 585
R1762 B.n657 B.n656 585
R1763 B.n655 B.n90 585
R1764 B.n654 B.n653 585
R1765 B.n652 B.n91 585
R1766 B.n651 B.n650 585
R1767 B.n649 B.n92 585
R1768 B.n648 B.n647 585
R1769 B.n646 B.n93 585
R1770 B.n835 B.n26 585
R1771 B.n837 B.n836 585
R1772 B.n838 B.n25 585
R1773 B.n840 B.n839 585
R1774 B.n841 B.n24 585
R1775 B.n843 B.n842 585
R1776 B.n844 B.n23 585
R1777 B.n846 B.n845 585
R1778 B.n847 B.n22 585
R1779 B.n849 B.n848 585
R1780 B.n850 B.n21 585
R1781 B.n852 B.n851 585
R1782 B.n853 B.n20 585
R1783 B.n855 B.n854 585
R1784 B.n856 B.n19 585
R1785 B.n858 B.n857 585
R1786 B.n859 B.n18 585
R1787 B.n861 B.n860 585
R1788 B.n862 B.n17 585
R1789 B.n864 B.n863 585
R1790 B.n865 B.n16 585
R1791 B.n867 B.n866 585
R1792 B.n868 B.n15 585
R1793 B.n870 B.n869 585
R1794 B.n871 B.n14 585
R1795 B.n873 B.n872 585
R1796 B.n874 B.n13 585
R1797 B.n876 B.n875 585
R1798 B.n877 B.n12 585
R1799 B.n879 B.n878 585
R1800 B.n880 B.n11 585
R1801 B.n882 B.n881 585
R1802 B.n883 B.n10 585
R1803 B.n885 B.n884 585
R1804 B.n886 B.n9 585
R1805 B.n888 B.n887 585
R1806 B.n889 B.n8 585
R1807 B.n891 B.n890 585
R1808 B.n892 B.n7 585
R1809 B.n894 B.n893 585
R1810 B.n895 B.n6 585
R1811 B.n897 B.n896 585
R1812 B.n898 B.n5 585
R1813 B.n900 B.n899 585
R1814 B.n901 B.n4 585
R1815 B.n903 B.n902 585
R1816 B.n904 B.n3 585
R1817 B.n906 B.n905 585
R1818 B.n907 B.n0 585
R1819 B.n2 B.n1 585
R1820 B.n233 B.n232 585
R1821 B.n234 B.n231 585
R1822 B.n236 B.n235 585
R1823 B.n237 B.n230 585
R1824 B.n239 B.n238 585
R1825 B.n240 B.n229 585
R1826 B.n242 B.n241 585
R1827 B.n243 B.n228 585
R1828 B.n245 B.n244 585
R1829 B.n246 B.n227 585
R1830 B.n248 B.n247 585
R1831 B.n249 B.n226 585
R1832 B.n251 B.n250 585
R1833 B.n252 B.n225 585
R1834 B.n254 B.n253 585
R1835 B.n255 B.n224 585
R1836 B.n257 B.n256 585
R1837 B.n258 B.n223 585
R1838 B.n260 B.n259 585
R1839 B.n261 B.n222 585
R1840 B.n263 B.n262 585
R1841 B.n264 B.n221 585
R1842 B.n266 B.n265 585
R1843 B.n267 B.n220 585
R1844 B.n269 B.n268 585
R1845 B.n270 B.n219 585
R1846 B.n272 B.n271 585
R1847 B.n273 B.n218 585
R1848 B.n275 B.n274 585
R1849 B.n276 B.n217 585
R1850 B.n278 B.n277 585
R1851 B.n279 B.n216 585
R1852 B.n281 B.n280 585
R1853 B.n282 B.n215 585
R1854 B.n284 B.n283 585
R1855 B.n285 B.n214 585
R1856 B.n287 B.n286 585
R1857 B.n288 B.n213 585
R1858 B.n290 B.n289 585
R1859 B.n291 B.n212 585
R1860 B.n293 B.n292 585
R1861 B.n294 B.n211 585
R1862 B.n296 B.n295 585
R1863 B.n297 B.n210 585
R1864 B.n299 B.n298 585
R1865 B.n300 B.n209 585
R1866 B.n302 B.n301 585
R1867 B.n303 B.n208 585
R1868 B.n304 B.n303 535.745
R1869 B.n494 B.n143 535.745
R1870 B.n644 B.n93 535.745
R1871 B.n835 B.n834 535.745
R1872 B.n404 B.t10 529.755
R1873 B.n62 B.t5 529.755
R1874 B.n178 B.t1 529.755
R1875 B.n56 B.t8 529.755
R1876 B.n405 B.t11 475.065
R1877 B.n63 B.t4 475.065
R1878 B.n179 B.t2 475.065
R1879 B.n57 B.t7 475.065
R1880 B.n178 B.t0 377.445
R1881 B.n404 B.t9 377.445
R1882 B.n62 B.t3 377.445
R1883 B.n56 B.t6 377.445
R1884 B.n909 B.n908 256.663
R1885 B.n908 B.n907 235.042
R1886 B.n908 B.n2 235.042
R1887 B.n304 B.n207 163.367
R1888 B.n308 B.n207 163.367
R1889 B.n309 B.n308 163.367
R1890 B.n310 B.n309 163.367
R1891 B.n310 B.n205 163.367
R1892 B.n314 B.n205 163.367
R1893 B.n315 B.n314 163.367
R1894 B.n316 B.n315 163.367
R1895 B.n316 B.n203 163.367
R1896 B.n320 B.n203 163.367
R1897 B.n321 B.n320 163.367
R1898 B.n322 B.n321 163.367
R1899 B.n322 B.n201 163.367
R1900 B.n326 B.n201 163.367
R1901 B.n327 B.n326 163.367
R1902 B.n328 B.n327 163.367
R1903 B.n328 B.n199 163.367
R1904 B.n332 B.n199 163.367
R1905 B.n333 B.n332 163.367
R1906 B.n334 B.n333 163.367
R1907 B.n334 B.n197 163.367
R1908 B.n338 B.n197 163.367
R1909 B.n339 B.n338 163.367
R1910 B.n340 B.n339 163.367
R1911 B.n340 B.n195 163.367
R1912 B.n344 B.n195 163.367
R1913 B.n345 B.n344 163.367
R1914 B.n346 B.n345 163.367
R1915 B.n346 B.n193 163.367
R1916 B.n350 B.n193 163.367
R1917 B.n351 B.n350 163.367
R1918 B.n352 B.n351 163.367
R1919 B.n352 B.n191 163.367
R1920 B.n356 B.n191 163.367
R1921 B.n357 B.n356 163.367
R1922 B.n358 B.n357 163.367
R1923 B.n358 B.n189 163.367
R1924 B.n362 B.n189 163.367
R1925 B.n363 B.n362 163.367
R1926 B.n364 B.n363 163.367
R1927 B.n364 B.n187 163.367
R1928 B.n368 B.n187 163.367
R1929 B.n369 B.n368 163.367
R1930 B.n370 B.n369 163.367
R1931 B.n370 B.n185 163.367
R1932 B.n374 B.n185 163.367
R1933 B.n375 B.n374 163.367
R1934 B.n376 B.n375 163.367
R1935 B.n376 B.n183 163.367
R1936 B.n380 B.n183 163.367
R1937 B.n381 B.n380 163.367
R1938 B.n382 B.n381 163.367
R1939 B.n382 B.n181 163.367
R1940 B.n386 B.n181 163.367
R1941 B.n387 B.n386 163.367
R1942 B.n388 B.n387 163.367
R1943 B.n388 B.n177 163.367
R1944 B.n393 B.n177 163.367
R1945 B.n394 B.n393 163.367
R1946 B.n395 B.n394 163.367
R1947 B.n395 B.n175 163.367
R1948 B.n399 B.n175 163.367
R1949 B.n400 B.n399 163.367
R1950 B.n401 B.n400 163.367
R1951 B.n401 B.n173 163.367
R1952 B.n408 B.n173 163.367
R1953 B.n409 B.n408 163.367
R1954 B.n410 B.n409 163.367
R1955 B.n410 B.n171 163.367
R1956 B.n414 B.n171 163.367
R1957 B.n415 B.n414 163.367
R1958 B.n416 B.n415 163.367
R1959 B.n416 B.n169 163.367
R1960 B.n420 B.n169 163.367
R1961 B.n421 B.n420 163.367
R1962 B.n422 B.n421 163.367
R1963 B.n422 B.n167 163.367
R1964 B.n426 B.n167 163.367
R1965 B.n427 B.n426 163.367
R1966 B.n428 B.n427 163.367
R1967 B.n428 B.n165 163.367
R1968 B.n432 B.n165 163.367
R1969 B.n433 B.n432 163.367
R1970 B.n434 B.n433 163.367
R1971 B.n434 B.n163 163.367
R1972 B.n438 B.n163 163.367
R1973 B.n439 B.n438 163.367
R1974 B.n440 B.n439 163.367
R1975 B.n440 B.n161 163.367
R1976 B.n444 B.n161 163.367
R1977 B.n445 B.n444 163.367
R1978 B.n446 B.n445 163.367
R1979 B.n446 B.n159 163.367
R1980 B.n450 B.n159 163.367
R1981 B.n451 B.n450 163.367
R1982 B.n452 B.n451 163.367
R1983 B.n452 B.n157 163.367
R1984 B.n456 B.n157 163.367
R1985 B.n457 B.n456 163.367
R1986 B.n458 B.n457 163.367
R1987 B.n458 B.n155 163.367
R1988 B.n462 B.n155 163.367
R1989 B.n463 B.n462 163.367
R1990 B.n464 B.n463 163.367
R1991 B.n464 B.n153 163.367
R1992 B.n468 B.n153 163.367
R1993 B.n469 B.n468 163.367
R1994 B.n470 B.n469 163.367
R1995 B.n470 B.n151 163.367
R1996 B.n474 B.n151 163.367
R1997 B.n475 B.n474 163.367
R1998 B.n476 B.n475 163.367
R1999 B.n476 B.n149 163.367
R2000 B.n480 B.n149 163.367
R2001 B.n481 B.n480 163.367
R2002 B.n482 B.n481 163.367
R2003 B.n482 B.n147 163.367
R2004 B.n486 B.n147 163.367
R2005 B.n487 B.n486 163.367
R2006 B.n488 B.n487 163.367
R2007 B.n488 B.n145 163.367
R2008 B.n492 B.n145 163.367
R2009 B.n493 B.n492 163.367
R2010 B.n494 B.n493 163.367
R2011 B.n644 B.n643 163.367
R2012 B.n643 B.n642 163.367
R2013 B.n642 B.n95 163.367
R2014 B.n638 B.n95 163.367
R2015 B.n638 B.n637 163.367
R2016 B.n637 B.n636 163.367
R2017 B.n636 B.n97 163.367
R2018 B.n632 B.n97 163.367
R2019 B.n632 B.n631 163.367
R2020 B.n631 B.n630 163.367
R2021 B.n630 B.n99 163.367
R2022 B.n626 B.n99 163.367
R2023 B.n626 B.n625 163.367
R2024 B.n625 B.n624 163.367
R2025 B.n624 B.n101 163.367
R2026 B.n620 B.n101 163.367
R2027 B.n620 B.n619 163.367
R2028 B.n619 B.n618 163.367
R2029 B.n618 B.n103 163.367
R2030 B.n614 B.n103 163.367
R2031 B.n614 B.n613 163.367
R2032 B.n613 B.n612 163.367
R2033 B.n612 B.n105 163.367
R2034 B.n608 B.n105 163.367
R2035 B.n608 B.n607 163.367
R2036 B.n607 B.n606 163.367
R2037 B.n606 B.n107 163.367
R2038 B.n602 B.n107 163.367
R2039 B.n602 B.n601 163.367
R2040 B.n601 B.n600 163.367
R2041 B.n600 B.n109 163.367
R2042 B.n596 B.n109 163.367
R2043 B.n596 B.n595 163.367
R2044 B.n595 B.n594 163.367
R2045 B.n594 B.n111 163.367
R2046 B.n590 B.n111 163.367
R2047 B.n590 B.n589 163.367
R2048 B.n589 B.n588 163.367
R2049 B.n588 B.n113 163.367
R2050 B.n584 B.n113 163.367
R2051 B.n584 B.n583 163.367
R2052 B.n583 B.n582 163.367
R2053 B.n582 B.n115 163.367
R2054 B.n578 B.n115 163.367
R2055 B.n578 B.n577 163.367
R2056 B.n577 B.n576 163.367
R2057 B.n576 B.n117 163.367
R2058 B.n572 B.n117 163.367
R2059 B.n572 B.n571 163.367
R2060 B.n571 B.n570 163.367
R2061 B.n570 B.n119 163.367
R2062 B.n566 B.n119 163.367
R2063 B.n566 B.n565 163.367
R2064 B.n565 B.n564 163.367
R2065 B.n564 B.n121 163.367
R2066 B.n560 B.n121 163.367
R2067 B.n560 B.n559 163.367
R2068 B.n559 B.n558 163.367
R2069 B.n558 B.n123 163.367
R2070 B.n554 B.n123 163.367
R2071 B.n554 B.n553 163.367
R2072 B.n553 B.n552 163.367
R2073 B.n552 B.n125 163.367
R2074 B.n548 B.n125 163.367
R2075 B.n548 B.n547 163.367
R2076 B.n547 B.n546 163.367
R2077 B.n546 B.n127 163.367
R2078 B.n542 B.n127 163.367
R2079 B.n542 B.n541 163.367
R2080 B.n541 B.n540 163.367
R2081 B.n540 B.n129 163.367
R2082 B.n536 B.n129 163.367
R2083 B.n536 B.n535 163.367
R2084 B.n535 B.n534 163.367
R2085 B.n534 B.n131 163.367
R2086 B.n530 B.n131 163.367
R2087 B.n530 B.n529 163.367
R2088 B.n529 B.n528 163.367
R2089 B.n528 B.n133 163.367
R2090 B.n524 B.n133 163.367
R2091 B.n524 B.n523 163.367
R2092 B.n523 B.n522 163.367
R2093 B.n522 B.n135 163.367
R2094 B.n518 B.n135 163.367
R2095 B.n518 B.n517 163.367
R2096 B.n517 B.n516 163.367
R2097 B.n516 B.n137 163.367
R2098 B.n512 B.n137 163.367
R2099 B.n512 B.n511 163.367
R2100 B.n511 B.n510 163.367
R2101 B.n510 B.n139 163.367
R2102 B.n506 B.n139 163.367
R2103 B.n506 B.n505 163.367
R2104 B.n505 B.n504 163.367
R2105 B.n504 B.n141 163.367
R2106 B.n500 B.n141 163.367
R2107 B.n500 B.n499 163.367
R2108 B.n499 B.n498 163.367
R2109 B.n498 B.n143 163.367
R2110 B.n834 B.n27 163.367
R2111 B.n830 B.n27 163.367
R2112 B.n830 B.n829 163.367
R2113 B.n829 B.n828 163.367
R2114 B.n828 B.n29 163.367
R2115 B.n824 B.n29 163.367
R2116 B.n824 B.n823 163.367
R2117 B.n823 B.n822 163.367
R2118 B.n822 B.n31 163.367
R2119 B.n818 B.n31 163.367
R2120 B.n818 B.n817 163.367
R2121 B.n817 B.n816 163.367
R2122 B.n816 B.n33 163.367
R2123 B.n812 B.n33 163.367
R2124 B.n812 B.n811 163.367
R2125 B.n811 B.n810 163.367
R2126 B.n810 B.n35 163.367
R2127 B.n806 B.n35 163.367
R2128 B.n806 B.n805 163.367
R2129 B.n805 B.n804 163.367
R2130 B.n804 B.n37 163.367
R2131 B.n800 B.n37 163.367
R2132 B.n800 B.n799 163.367
R2133 B.n799 B.n798 163.367
R2134 B.n798 B.n39 163.367
R2135 B.n794 B.n39 163.367
R2136 B.n794 B.n793 163.367
R2137 B.n793 B.n792 163.367
R2138 B.n792 B.n41 163.367
R2139 B.n788 B.n41 163.367
R2140 B.n788 B.n787 163.367
R2141 B.n787 B.n786 163.367
R2142 B.n786 B.n43 163.367
R2143 B.n782 B.n43 163.367
R2144 B.n782 B.n781 163.367
R2145 B.n781 B.n780 163.367
R2146 B.n780 B.n45 163.367
R2147 B.n776 B.n45 163.367
R2148 B.n776 B.n775 163.367
R2149 B.n775 B.n774 163.367
R2150 B.n774 B.n47 163.367
R2151 B.n770 B.n47 163.367
R2152 B.n770 B.n769 163.367
R2153 B.n769 B.n768 163.367
R2154 B.n768 B.n49 163.367
R2155 B.n764 B.n49 163.367
R2156 B.n764 B.n763 163.367
R2157 B.n763 B.n762 163.367
R2158 B.n762 B.n51 163.367
R2159 B.n758 B.n51 163.367
R2160 B.n758 B.n757 163.367
R2161 B.n757 B.n756 163.367
R2162 B.n756 B.n53 163.367
R2163 B.n752 B.n53 163.367
R2164 B.n752 B.n751 163.367
R2165 B.n751 B.n750 163.367
R2166 B.n750 B.n55 163.367
R2167 B.n745 B.n55 163.367
R2168 B.n745 B.n744 163.367
R2169 B.n744 B.n743 163.367
R2170 B.n743 B.n59 163.367
R2171 B.n739 B.n59 163.367
R2172 B.n739 B.n738 163.367
R2173 B.n738 B.n737 163.367
R2174 B.n737 B.n61 163.367
R2175 B.n733 B.n61 163.367
R2176 B.n733 B.n732 163.367
R2177 B.n732 B.n65 163.367
R2178 B.n728 B.n65 163.367
R2179 B.n728 B.n727 163.367
R2180 B.n727 B.n726 163.367
R2181 B.n726 B.n67 163.367
R2182 B.n722 B.n67 163.367
R2183 B.n722 B.n721 163.367
R2184 B.n721 B.n720 163.367
R2185 B.n720 B.n69 163.367
R2186 B.n716 B.n69 163.367
R2187 B.n716 B.n715 163.367
R2188 B.n715 B.n714 163.367
R2189 B.n714 B.n71 163.367
R2190 B.n710 B.n71 163.367
R2191 B.n710 B.n709 163.367
R2192 B.n709 B.n708 163.367
R2193 B.n708 B.n73 163.367
R2194 B.n704 B.n73 163.367
R2195 B.n704 B.n703 163.367
R2196 B.n703 B.n702 163.367
R2197 B.n702 B.n75 163.367
R2198 B.n698 B.n75 163.367
R2199 B.n698 B.n697 163.367
R2200 B.n697 B.n696 163.367
R2201 B.n696 B.n77 163.367
R2202 B.n692 B.n77 163.367
R2203 B.n692 B.n691 163.367
R2204 B.n691 B.n690 163.367
R2205 B.n690 B.n79 163.367
R2206 B.n686 B.n79 163.367
R2207 B.n686 B.n685 163.367
R2208 B.n685 B.n684 163.367
R2209 B.n684 B.n81 163.367
R2210 B.n680 B.n81 163.367
R2211 B.n680 B.n679 163.367
R2212 B.n679 B.n678 163.367
R2213 B.n678 B.n83 163.367
R2214 B.n674 B.n83 163.367
R2215 B.n674 B.n673 163.367
R2216 B.n673 B.n672 163.367
R2217 B.n672 B.n85 163.367
R2218 B.n668 B.n85 163.367
R2219 B.n668 B.n667 163.367
R2220 B.n667 B.n666 163.367
R2221 B.n666 B.n87 163.367
R2222 B.n662 B.n87 163.367
R2223 B.n662 B.n661 163.367
R2224 B.n661 B.n660 163.367
R2225 B.n660 B.n89 163.367
R2226 B.n656 B.n89 163.367
R2227 B.n656 B.n655 163.367
R2228 B.n655 B.n654 163.367
R2229 B.n654 B.n91 163.367
R2230 B.n650 B.n91 163.367
R2231 B.n650 B.n649 163.367
R2232 B.n649 B.n648 163.367
R2233 B.n648 B.n93 163.367
R2234 B.n836 B.n835 163.367
R2235 B.n836 B.n25 163.367
R2236 B.n840 B.n25 163.367
R2237 B.n841 B.n840 163.367
R2238 B.n842 B.n841 163.367
R2239 B.n842 B.n23 163.367
R2240 B.n846 B.n23 163.367
R2241 B.n847 B.n846 163.367
R2242 B.n848 B.n847 163.367
R2243 B.n848 B.n21 163.367
R2244 B.n852 B.n21 163.367
R2245 B.n853 B.n852 163.367
R2246 B.n854 B.n853 163.367
R2247 B.n854 B.n19 163.367
R2248 B.n858 B.n19 163.367
R2249 B.n859 B.n858 163.367
R2250 B.n860 B.n859 163.367
R2251 B.n860 B.n17 163.367
R2252 B.n864 B.n17 163.367
R2253 B.n865 B.n864 163.367
R2254 B.n866 B.n865 163.367
R2255 B.n866 B.n15 163.367
R2256 B.n870 B.n15 163.367
R2257 B.n871 B.n870 163.367
R2258 B.n872 B.n871 163.367
R2259 B.n872 B.n13 163.367
R2260 B.n876 B.n13 163.367
R2261 B.n877 B.n876 163.367
R2262 B.n878 B.n877 163.367
R2263 B.n878 B.n11 163.367
R2264 B.n882 B.n11 163.367
R2265 B.n883 B.n882 163.367
R2266 B.n884 B.n883 163.367
R2267 B.n884 B.n9 163.367
R2268 B.n888 B.n9 163.367
R2269 B.n889 B.n888 163.367
R2270 B.n890 B.n889 163.367
R2271 B.n890 B.n7 163.367
R2272 B.n894 B.n7 163.367
R2273 B.n895 B.n894 163.367
R2274 B.n896 B.n895 163.367
R2275 B.n896 B.n5 163.367
R2276 B.n900 B.n5 163.367
R2277 B.n901 B.n900 163.367
R2278 B.n902 B.n901 163.367
R2279 B.n902 B.n3 163.367
R2280 B.n906 B.n3 163.367
R2281 B.n907 B.n906 163.367
R2282 B.n232 B.n2 163.367
R2283 B.n232 B.n231 163.367
R2284 B.n236 B.n231 163.367
R2285 B.n237 B.n236 163.367
R2286 B.n238 B.n237 163.367
R2287 B.n238 B.n229 163.367
R2288 B.n242 B.n229 163.367
R2289 B.n243 B.n242 163.367
R2290 B.n244 B.n243 163.367
R2291 B.n244 B.n227 163.367
R2292 B.n248 B.n227 163.367
R2293 B.n249 B.n248 163.367
R2294 B.n250 B.n249 163.367
R2295 B.n250 B.n225 163.367
R2296 B.n254 B.n225 163.367
R2297 B.n255 B.n254 163.367
R2298 B.n256 B.n255 163.367
R2299 B.n256 B.n223 163.367
R2300 B.n260 B.n223 163.367
R2301 B.n261 B.n260 163.367
R2302 B.n262 B.n261 163.367
R2303 B.n262 B.n221 163.367
R2304 B.n266 B.n221 163.367
R2305 B.n267 B.n266 163.367
R2306 B.n268 B.n267 163.367
R2307 B.n268 B.n219 163.367
R2308 B.n272 B.n219 163.367
R2309 B.n273 B.n272 163.367
R2310 B.n274 B.n273 163.367
R2311 B.n274 B.n217 163.367
R2312 B.n278 B.n217 163.367
R2313 B.n279 B.n278 163.367
R2314 B.n280 B.n279 163.367
R2315 B.n280 B.n215 163.367
R2316 B.n284 B.n215 163.367
R2317 B.n285 B.n284 163.367
R2318 B.n286 B.n285 163.367
R2319 B.n286 B.n213 163.367
R2320 B.n290 B.n213 163.367
R2321 B.n291 B.n290 163.367
R2322 B.n292 B.n291 163.367
R2323 B.n292 B.n211 163.367
R2324 B.n296 B.n211 163.367
R2325 B.n297 B.n296 163.367
R2326 B.n298 B.n297 163.367
R2327 B.n298 B.n209 163.367
R2328 B.n302 B.n209 163.367
R2329 B.n303 B.n302 163.367
R2330 B.n391 B.n179 59.5399
R2331 B.n406 B.n405 59.5399
R2332 B.n64 B.n63 59.5399
R2333 B.n747 B.n57 59.5399
R2334 B.n179 B.n178 54.6914
R2335 B.n405 B.n404 54.6914
R2336 B.n63 B.n62 54.6914
R2337 B.n57 B.n56 54.6914
R2338 B.n833 B.n26 34.8103
R2339 B.n646 B.n645 34.8103
R2340 B.n305 B.n208 34.8103
R2341 B.n496 B.n495 34.8103
R2342 B B.n909 18.0485
R2343 B.n837 B.n26 10.6151
R2344 B.n838 B.n837 10.6151
R2345 B.n839 B.n838 10.6151
R2346 B.n839 B.n24 10.6151
R2347 B.n843 B.n24 10.6151
R2348 B.n844 B.n843 10.6151
R2349 B.n845 B.n844 10.6151
R2350 B.n845 B.n22 10.6151
R2351 B.n849 B.n22 10.6151
R2352 B.n850 B.n849 10.6151
R2353 B.n851 B.n850 10.6151
R2354 B.n851 B.n20 10.6151
R2355 B.n855 B.n20 10.6151
R2356 B.n856 B.n855 10.6151
R2357 B.n857 B.n856 10.6151
R2358 B.n857 B.n18 10.6151
R2359 B.n861 B.n18 10.6151
R2360 B.n862 B.n861 10.6151
R2361 B.n863 B.n862 10.6151
R2362 B.n863 B.n16 10.6151
R2363 B.n867 B.n16 10.6151
R2364 B.n868 B.n867 10.6151
R2365 B.n869 B.n868 10.6151
R2366 B.n869 B.n14 10.6151
R2367 B.n873 B.n14 10.6151
R2368 B.n874 B.n873 10.6151
R2369 B.n875 B.n874 10.6151
R2370 B.n875 B.n12 10.6151
R2371 B.n879 B.n12 10.6151
R2372 B.n880 B.n879 10.6151
R2373 B.n881 B.n880 10.6151
R2374 B.n881 B.n10 10.6151
R2375 B.n885 B.n10 10.6151
R2376 B.n886 B.n885 10.6151
R2377 B.n887 B.n886 10.6151
R2378 B.n887 B.n8 10.6151
R2379 B.n891 B.n8 10.6151
R2380 B.n892 B.n891 10.6151
R2381 B.n893 B.n892 10.6151
R2382 B.n893 B.n6 10.6151
R2383 B.n897 B.n6 10.6151
R2384 B.n898 B.n897 10.6151
R2385 B.n899 B.n898 10.6151
R2386 B.n899 B.n4 10.6151
R2387 B.n903 B.n4 10.6151
R2388 B.n904 B.n903 10.6151
R2389 B.n905 B.n904 10.6151
R2390 B.n905 B.n0 10.6151
R2391 B.n833 B.n832 10.6151
R2392 B.n832 B.n831 10.6151
R2393 B.n831 B.n28 10.6151
R2394 B.n827 B.n28 10.6151
R2395 B.n827 B.n826 10.6151
R2396 B.n826 B.n825 10.6151
R2397 B.n825 B.n30 10.6151
R2398 B.n821 B.n30 10.6151
R2399 B.n821 B.n820 10.6151
R2400 B.n820 B.n819 10.6151
R2401 B.n819 B.n32 10.6151
R2402 B.n815 B.n32 10.6151
R2403 B.n815 B.n814 10.6151
R2404 B.n814 B.n813 10.6151
R2405 B.n813 B.n34 10.6151
R2406 B.n809 B.n34 10.6151
R2407 B.n809 B.n808 10.6151
R2408 B.n808 B.n807 10.6151
R2409 B.n807 B.n36 10.6151
R2410 B.n803 B.n36 10.6151
R2411 B.n803 B.n802 10.6151
R2412 B.n802 B.n801 10.6151
R2413 B.n801 B.n38 10.6151
R2414 B.n797 B.n38 10.6151
R2415 B.n797 B.n796 10.6151
R2416 B.n796 B.n795 10.6151
R2417 B.n795 B.n40 10.6151
R2418 B.n791 B.n40 10.6151
R2419 B.n791 B.n790 10.6151
R2420 B.n790 B.n789 10.6151
R2421 B.n789 B.n42 10.6151
R2422 B.n785 B.n42 10.6151
R2423 B.n785 B.n784 10.6151
R2424 B.n784 B.n783 10.6151
R2425 B.n783 B.n44 10.6151
R2426 B.n779 B.n44 10.6151
R2427 B.n779 B.n778 10.6151
R2428 B.n778 B.n777 10.6151
R2429 B.n777 B.n46 10.6151
R2430 B.n773 B.n46 10.6151
R2431 B.n773 B.n772 10.6151
R2432 B.n772 B.n771 10.6151
R2433 B.n771 B.n48 10.6151
R2434 B.n767 B.n48 10.6151
R2435 B.n767 B.n766 10.6151
R2436 B.n766 B.n765 10.6151
R2437 B.n765 B.n50 10.6151
R2438 B.n761 B.n50 10.6151
R2439 B.n761 B.n760 10.6151
R2440 B.n760 B.n759 10.6151
R2441 B.n759 B.n52 10.6151
R2442 B.n755 B.n52 10.6151
R2443 B.n755 B.n754 10.6151
R2444 B.n754 B.n753 10.6151
R2445 B.n753 B.n54 10.6151
R2446 B.n749 B.n54 10.6151
R2447 B.n749 B.n748 10.6151
R2448 B.n746 B.n58 10.6151
R2449 B.n742 B.n58 10.6151
R2450 B.n742 B.n741 10.6151
R2451 B.n741 B.n740 10.6151
R2452 B.n740 B.n60 10.6151
R2453 B.n736 B.n60 10.6151
R2454 B.n736 B.n735 10.6151
R2455 B.n735 B.n734 10.6151
R2456 B.n731 B.n730 10.6151
R2457 B.n730 B.n729 10.6151
R2458 B.n729 B.n66 10.6151
R2459 B.n725 B.n66 10.6151
R2460 B.n725 B.n724 10.6151
R2461 B.n724 B.n723 10.6151
R2462 B.n723 B.n68 10.6151
R2463 B.n719 B.n68 10.6151
R2464 B.n719 B.n718 10.6151
R2465 B.n718 B.n717 10.6151
R2466 B.n717 B.n70 10.6151
R2467 B.n713 B.n70 10.6151
R2468 B.n713 B.n712 10.6151
R2469 B.n712 B.n711 10.6151
R2470 B.n711 B.n72 10.6151
R2471 B.n707 B.n72 10.6151
R2472 B.n707 B.n706 10.6151
R2473 B.n706 B.n705 10.6151
R2474 B.n705 B.n74 10.6151
R2475 B.n701 B.n74 10.6151
R2476 B.n701 B.n700 10.6151
R2477 B.n700 B.n699 10.6151
R2478 B.n699 B.n76 10.6151
R2479 B.n695 B.n76 10.6151
R2480 B.n695 B.n694 10.6151
R2481 B.n694 B.n693 10.6151
R2482 B.n693 B.n78 10.6151
R2483 B.n689 B.n78 10.6151
R2484 B.n689 B.n688 10.6151
R2485 B.n688 B.n687 10.6151
R2486 B.n687 B.n80 10.6151
R2487 B.n683 B.n80 10.6151
R2488 B.n683 B.n682 10.6151
R2489 B.n682 B.n681 10.6151
R2490 B.n681 B.n82 10.6151
R2491 B.n677 B.n82 10.6151
R2492 B.n677 B.n676 10.6151
R2493 B.n676 B.n675 10.6151
R2494 B.n675 B.n84 10.6151
R2495 B.n671 B.n84 10.6151
R2496 B.n671 B.n670 10.6151
R2497 B.n670 B.n669 10.6151
R2498 B.n669 B.n86 10.6151
R2499 B.n665 B.n86 10.6151
R2500 B.n665 B.n664 10.6151
R2501 B.n664 B.n663 10.6151
R2502 B.n663 B.n88 10.6151
R2503 B.n659 B.n88 10.6151
R2504 B.n659 B.n658 10.6151
R2505 B.n658 B.n657 10.6151
R2506 B.n657 B.n90 10.6151
R2507 B.n653 B.n90 10.6151
R2508 B.n653 B.n652 10.6151
R2509 B.n652 B.n651 10.6151
R2510 B.n651 B.n92 10.6151
R2511 B.n647 B.n92 10.6151
R2512 B.n647 B.n646 10.6151
R2513 B.n645 B.n94 10.6151
R2514 B.n641 B.n94 10.6151
R2515 B.n641 B.n640 10.6151
R2516 B.n640 B.n639 10.6151
R2517 B.n639 B.n96 10.6151
R2518 B.n635 B.n96 10.6151
R2519 B.n635 B.n634 10.6151
R2520 B.n634 B.n633 10.6151
R2521 B.n633 B.n98 10.6151
R2522 B.n629 B.n98 10.6151
R2523 B.n629 B.n628 10.6151
R2524 B.n628 B.n627 10.6151
R2525 B.n627 B.n100 10.6151
R2526 B.n623 B.n100 10.6151
R2527 B.n623 B.n622 10.6151
R2528 B.n622 B.n621 10.6151
R2529 B.n621 B.n102 10.6151
R2530 B.n617 B.n102 10.6151
R2531 B.n617 B.n616 10.6151
R2532 B.n616 B.n615 10.6151
R2533 B.n615 B.n104 10.6151
R2534 B.n611 B.n104 10.6151
R2535 B.n611 B.n610 10.6151
R2536 B.n610 B.n609 10.6151
R2537 B.n609 B.n106 10.6151
R2538 B.n605 B.n106 10.6151
R2539 B.n605 B.n604 10.6151
R2540 B.n604 B.n603 10.6151
R2541 B.n603 B.n108 10.6151
R2542 B.n599 B.n108 10.6151
R2543 B.n599 B.n598 10.6151
R2544 B.n598 B.n597 10.6151
R2545 B.n597 B.n110 10.6151
R2546 B.n593 B.n110 10.6151
R2547 B.n593 B.n592 10.6151
R2548 B.n592 B.n591 10.6151
R2549 B.n591 B.n112 10.6151
R2550 B.n587 B.n112 10.6151
R2551 B.n587 B.n586 10.6151
R2552 B.n586 B.n585 10.6151
R2553 B.n585 B.n114 10.6151
R2554 B.n581 B.n114 10.6151
R2555 B.n581 B.n580 10.6151
R2556 B.n580 B.n579 10.6151
R2557 B.n579 B.n116 10.6151
R2558 B.n575 B.n116 10.6151
R2559 B.n575 B.n574 10.6151
R2560 B.n574 B.n573 10.6151
R2561 B.n573 B.n118 10.6151
R2562 B.n569 B.n118 10.6151
R2563 B.n569 B.n568 10.6151
R2564 B.n568 B.n567 10.6151
R2565 B.n567 B.n120 10.6151
R2566 B.n563 B.n120 10.6151
R2567 B.n563 B.n562 10.6151
R2568 B.n562 B.n561 10.6151
R2569 B.n561 B.n122 10.6151
R2570 B.n557 B.n122 10.6151
R2571 B.n557 B.n556 10.6151
R2572 B.n556 B.n555 10.6151
R2573 B.n555 B.n124 10.6151
R2574 B.n551 B.n124 10.6151
R2575 B.n551 B.n550 10.6151
R2576 B.n550 B.n549 10.6151
R2577 B.n549 B.n126 10.6151
R2578 B.n545 B.n126 10.6151
R2579 B.n545 B.n544 10.6151
R2580 B.n544 B.n543 10.6151
R2581 B.n543 B.n128 10.6151
R2582 B.n539 B.n128 10.6151
R2583 B.n539 B.n538 10.6151
R2584 B.n538 B.n537 10.6151
R2585 B.n537 B.n130 10.6151
R2586 B.n533 B.n130 10.6151
R2587 B.n533 B.n532 10.6151
R2588 B.n532 B.n531 10.6151
R2589 B.n531 B.n132 10.6151
R2590 B.n527 B.n132 10.6151
R2591 B.n527 B.n526 10.6151
R2592 B.n526 B.n525 10.6151
R2593 B.n525 B.n134 10.6151
R2594 B.n521 B.n134 10.6151
R2595 B.n521 B.n520 10.6151
R2596 B.n520 B.n519 10.6151
R2597 B.n519 B.n136 10.6151
R2598 B.n515 B.n136 10.6151
R2599 B.n515 B.n514 10.6151
R2600 B.n514 B.n513 10.6151
R2601 B.n513 B.n138 10.6151
R2602 B.n509 B.n138 10.6151
R2603 B.n509 B.n508 10.6151
R2604 B.n508 B.n507 10.6151
R2605 B.n507 B.n140 10.6151
R2606 B.n503 B.n140 10.6151
R2607 B.n503 B.n502 10.6151
R2608 B.n502 B.n501 10.6151
R2609 B.n501 B.n142 10.6151
R2610 B.n497 B.n142 10.6151
R2611 B.n497 B.n496 10.6151
R2612 B.n233 B.n1 10.6151
R2613 B.n234 B.n233 10.6151
R2614 B.n235 B.n234 10.6151
R2615 B.n235 B.n230 10.6151
R2616 B.n239 B.n230 10.6151
R2617 B.n240 B.n239 10.6151
R2618 B.n241 B.n240 10.6151
R2619 B.n241 B.n228 10.6151
R2620 B.n245 B.n228 10.6151
R2621 B.n246 B.n245 10.6151
R2622 B.n247 B.n246 10.6151
R2623 B.n247 B.n226 10.6151
R2624 B.n251 B.n226 10.6151
R2625 B.n252 B.n251 10.6151
R2626 B.n253 B.n252 10.6151
R2627 B.n253 B.n224 10.6151
R2628 B.n257 B.n224 10.6151
R2629 B.n258 B.n257 10.6151
R2630 B.n259 B.n258 10.6151
R2631 B.n259 B.n222 10.6151
R2632 B.n263 B.n222 10.6151
R2633 B.n264 B.n263 10.6151
R2634 B.n265 B.n264 10.6151
R2635 B.n265 B.n220 10.6151
R2636 B.n269 B.n220 10.6151
R2637 B.n270 B.n269 10.6151
R2638 B.n271 B.n270 10.6151
R2639 B.n271 B.n218 10.6151
R2640 B.n275 B.n218 10.6151
R2641 B.n276 B.n275 10.6151
R2642 B.n277 B.n276 10.6151
R2643 B.n277 B.n216 10.6151
R2644 B.n281 B.n216 10.6151
R2645 B.n282 B.n281 10.6151
R2646 B.n283 B.n282 10.6151
R2647 B.n283 B.n214 10.6151
R2648 B.n287 B.n214 10.6151
R2649 B.n288 B.n287 10.6151
R2650 B.n289 B.n288 10.6151
R2651 B.n289 B.n212 10.6151
R2652 B.n293 B.n212 10.6151
R2653 B.n294 B.n293 10.6151
R2654 B.n295 B.n294 10.6151
R2655 B.n295 B.n210 10.6151
R2656 B.n299 B.n210 10.6151
R2657 B.n300 B.n299 10.6151
R2658 B.n301 B.n300 10.6151
R2659 B.n301 B.n208 10.6151
R2660 B.n306 B.n305 10.6151
R2661 B.n307 B.n306 10.6151
R2662 B.n307 B.n206 10.6151
R2663 B.n311 B.n206 10.6151
R2664 B.n312 B.n311 10.6151
R2665 B.n313 B.n312 10.6151
R2666 B.n313 B.n204 10.6151
R2667 B.n317 B.n204 10.6151
R2668 B.n318 B.n317 10.6151
R2669 B.n319 B.n318 10.6151
R2670 B.n319 B.n202 10.6151
R2671 B.n323 B.n202 10.6151
R2672 B.n324 B.n323 10.6151
R2673 B.n325 B.n324 10.6151
R2674 B.n325 B.n200 10.6151
R2675 B.n329 B.n200 10.6151
R2676 B.n330 B.n329 10.6151
R2677 B.n331 B.n330 10.6151
R2678 B.n331 B.n198 10.6151
R2679 B.n335 B.n198 10.6151
R2680 B.n336 B.n335 10.6151
R2681 B.n337 B.n336 10.6151
R2682 B.n337 B.n196 10.6151
R2683 B.n341 B.n196 10.6151
R2684 B.n342 B.n341 10.6151
R2685 B.n343 B.n342 10.6151
R2686 B.n343 B.n194 10.6151
R2687 B.n347 B.n194 10.6151
R2688 B.n348 B.n347 10.6151
R2689 B.n349 B.n348 10.6151
R2690 B.n349 B.n192 10.6151
R2691 B.n353 B.n192 10.6151
R2692 B.n354 B.n353 10.6151
R2693 B.n355 B.n354 10.6151
R2694 B.n355 B.n190 10.6151
R2695 B.n359 B.n190 10.6151
R2696 B.n360 B.n359 10.6151
R2697 B.n361 B.n360 10.6151
R2698 B.n361 B.n188 10.6151
R2699 B.n365 B.n188 10.6151
R2700 B.n366 B.n365 10.6151
R2701 B.n367 B.n366 10.6151
R2702 B.n367 B.n186 10.6151
R2703 B.n371 B.n186 10.6151
R2704 B.n372 B.n371 10.6151
R2705 B.n373 B.n372 10.6151
R2706 B.n373 B.n184 10.6151
R2707 B.n377 B.n184 10.6151
R2708 B.n378 B.n377 10.6151
R2709 B.n379 B.n378 10.6151
R2710 B.n379 B.n182 10.6151
R2711 B.n383 B.n182 10.6151
R2712 B.n384 B.n383 10.6151
R2713 B.n385 B.n384 10.6151
R2714 B.n385 B.n180 10.6151
R2715 B.n389 B.n180 10.6151
R2716 B.n390 B.n389 10.6151
R2717 B.n392 B.n176 10.6151
R2718 B.n396 B.n176 10.6151
R2719 B.n397 B.n396 10.6151
R2720 B.n398 B.n397 10.6151
R2721 B.n398 B.n174 10.6151
R2722 B.n402 B.n174 10.6151
R2723 B.n403 B.n402 10.6151
R2724 B.n407 B.n403 10.6151
R2725 B.n411 B.n172 10.6151
R2726 B.n412 B.n411 10.6151
R2727 B.n413 B.n412 10.6151
R2728 B.n413 B.n170 10.6151
R2729 B.n417 B.n170 10.6151
R2730 B.n418 B.n417 10.6151
R2731 B.n419 B.n418 10.6151
R2732 B.n419 B.n168 10.6151
R2733 B.n423 B.n168 10.6151
R2734 B.n424 B.n423 10.6151
R2735 B.n425 B.n424 10.6151
R2736 B.n425 B.n166 10.6151
R2737 B.n429 B.n166 10.6151
R2738 B.n430 B.n429 10.6151
R2739 B.n431 B.n430 10.6151
R2740 B.n431 B.n164 10.6151
R2741 B.n435 B.n164 10.6151
R2742 B.n436 B.n435 10.6151
R2743 B.n437 B.n436 10.6151
R2744 B.n437 B.n162 10.6151
R2745 B.n441 B.n162 10.6151
R2746 B.n442 B.n441 10.6151
R2747 B.n443 B.n442 10.6151
R2748 B.n443 B.n160 10.6151
R2749 B.n447 B.n160 10.6151
R2750 B.n448 B.n447 10.6151
R2751 B.n449 B.n448 10.6151
R2752 B.n449 B.n158 10.6151
R2753 B.n453 B.n158 10.6151
R2754 B.n454 B.n453 10.6151
R2755 B.n455 B.n454 10.6151
R2756 B.n455 B.n156 10.6151
R2757 B.n459 B.n156 10.6151
R2758 B.n460 B.n459 10.6151
R2759 B.n461 B.n460 10.6151
R2760 B.n461 B.n154 10.6151
R2761 B.n465 B.n154 10.6151
R2762 B.n466 B.n465 10.6151
R2763 B.n467 B.n466 10.6151
R2764 B.n467 B.n152 10.6151
R2765 B.n471 B.n152 10.6151
R2766 B.n472 B.n471 10.6151
R2767 B.n473 B.n472 10.6151
R2768 B.n473 B.n150 10.6151
R2769 B.n477 B.n150 10.6151
R2770 B.n478 B.n477 10.6151
R2771 B.n479 B.n478 10.6151
R2772 B.n479 B.n148 10.6151
R2773 B.n483 B.n148 10.6151
R2774 B.n484 B.n483 10.6151
R2775 B.n485 B.n484 10.6151
R2776 B.n485 B.n146 10.6151
R2777 B.n489 B.n146 10.6151
R2778 B.n490 B.n489 10.6151
R2779 B.n491 B.n490 10.6151
R2780 B.n491 B.n144 10.6151
R2781 B.n495 B.n144 10.6151
R2782 B.n909 B.n0 8.11757
R2783 B.n909 B.n1 8.11757
R2784 B.n747 B.n746 6.5566
R2785 B.n734 B.n64 6.5566
R2786 B.n392 B.n391 6.5566
R2787 B.n407 B.n406 6.5566
R2788 B.n748 B.n747 4.05904
R2789 B.n731 B.n64 4.05904
R2790 B.n391 B.n390 4.05904
R2791 B.n406 B.n172 4.05904
C0 VP VN 8.54424f
C1 VDD1 VP 12.7299f
C2 w_n3790_n4472# VDD2 2.17971f
C3 B VN 1.26816f
C4 VDD1 B 1.76325f
C5 VTAIL VDD2 10.015901f
C6 B VP 2.09182f
C7 VN VDD2 12.3748f
C8 VTAIL w_n3790_n4472# 5.44101f
C9 VDD1 VDD2 1.72084f
C10 w_n3790_n4472# VN 7.77422f
C11 VDD1 w_n3790_n4472# 2.06962f
C12 VP VDD2 0.5084f
C13 B VDD2 1.85581f
C14 VTAIL VN 12.5002f
C15 VTAIL VDD1 9.96227f
C16 w_n3790_n4472# VP 8.26592f
C17 w_n3790_n4472# B 11.4952f
C18 VDD1 VN 0.151964f
C19 VTAIL VP 12.514299f
C20 VTAIL B 6.7322f
C21 VDD2 VSUBS 2.001692f
C22 VDD1 VSUBS 2.62592f
C23 VTAIL VSUBS 1.569238f
C24 VN VSUBS 6.82758f
C25 VP VSUBS 3.675086f
C26 B VSUBS 5.350127f
C27 w_n3790_n4472# VSUBS 0.207343p
C28 B.n0 VSUBS 0.006069f
C29 B.n1 VSUBS 0.006069f
C30 B.n2 VSUBS 0.008976f
C31 B.n3 VSUBS 0.006878f
C32 B.n4 VSUBS 0.006878f
C33 B.n5 VSUBS 0.006878f
C34 B.n6 VSUBS 0.006878f
C35 B.n7 VSUBS 0.006878f
C36 B.n8 VSUBS 0.006878f
C37 B.n9 VSUBS 0.006878f
C38 B.n10 VSUBS 0.006878f
C39 B.n11 VSUBS 0.006878f
C40 B.n12 VSUBS 0.006878f
C41 B.n13 VSUBS 0.006878f
C42 B.n14 VSUBS 0.006878f
C43 B.n15 VSUBS 0.006878f
C44 B.n16 VSUBS 0.006878f
C45 B.n17 VSUBS 0.006878f
C46 B.n18 VSUBS 0.006878f
C47 B.n19 VSUBS 0.006878f
C48 B.n20 VSUBS 0.006878f
C49 B.n21 VSUBS 0.006878f
C50 B.n22 VSUBS 0.006878f
C51 B.n23 VSUBS 0.006878f
C52 B.n24 VSUBS 0.006878f
C53 B.n25 VSUBS 0.006878f
C54 B.n26 VSUBS 0.016466f
C55 B.n27 VSUBS 0.006878f
C56 B.n28 VSUBS 0.006878f
C57 B.n29 VSUBS 0.006878f
C58 B.n30 VSUBS 0.006878f
C59 B.n31 VSUBS 0.006878f
C60 B.n32 VSUBS 0.006878f
C61 B.n33 VSUBS 0.006878f
C62 B.n34 VSUBS 0.006878f
C63 B.n35 VSUBS 0.006878f
C64 B.n36 VSUBS 0.006878f
C65 B.n37 VSUBS 0.006878f
C66 B.n38 VSUBS 0.006878f
C67 B.n39 VSUBS 0.006878f
C68 B.n40 VSUBS 0.006878f
C69 B.n41 VSUBS 0.006878f
C70 B.n42 VSUBS 0.006878f
C71 B.n43 VSUBS 0.006878f
C72 B.n44 VSUBS 0.006878f
C73 B.n45 VSUBS 0.006878f
C74 B.n46 VSUBS 0.006878f
C75 B.n47 VSUBS 0.006878f
C76 B.n48 VSUBS 0.006878f
C77 B.n49 VSUBS 0.006878f
C78 B.n50 VSUBS 0.006878f
C79 B.n51 VSUBS 0.006878f
C80 B.n52 VSUBS 0.006878f
C81 B.n53 VSUBS 0.006878f
C82 B.n54 VSUBS 0.006878f
C83 B.n55 VSUBS 0.006878f
C84 B.t7 VSUBS 0.333608f
C85 B.t8 VSUBS 0.36531f
C86 B.t6 VSUBS 1.89889f
C87 B.n56 VSUBS 0.557418f
C88 B.n57 VSUBS 0.31688f
C89 B.n58 VSUBS 0.006878f
C90 B.n59 VSUBS 0.006878f
C91 B.n60 VSUBS 0.006878f
C92 B.n61 VSUBS 0.006878f
C93 B.t4 VSUBS 0.333612f
C94 B.t5 VSUBS 0.365313f
C95 B.t3 VSUBS 1.89889f
C96 B.n62 VSUBS 0.557415f
C97 B.n63 VSUBS 0.316876f
C98 B.n64 VSUBS 0.015937f
C99 B.n65 VSUBS 0.006878f
C100 B.n66 VSUBS 0.006878f
C101 B.n67 VSUBS 0.006878f
C102 B.n68 VSUBS 0.006878f
C103 B.n69 VSUBS 0.006878f
C104 B.n70 VSUBS 0.006878f
C105 B.n71 VSUBS 0.006878f
C106 B.n72 VSUBS 0.006878f
C107 B.n73 VSUBS 0.006878f
C108 B.n74 VSUBS 0.006878f
C109 B.n75 VSUBS 0.006878f
C110 B.n76 VSUBS 0.006878f
C111 B.n77 VSUBS 0.006878f
C112 B.n78 VSUBS 0.006878f
C113 B.n79 VSUBS 0.006878f
C114 B.n80 VSUBS 0.006878f
C115 B.n81 VSUBS 0.006878f
C116 B.n82 VSUBS 0.006878f
C117 B.n83 VSUBS 0.006878f
C118 B.n84 VSUBS 0.006878f
C119 B.n85 VSUBS 0.006878f
C120 B.n86 VSUBS 0.006878f
C121 B.n87 VSUBS 0.006878f
C122 B.n88 VSUBS 0.006878f
C123 B.n89 VSUBS 0.006878f
C124 B.n90 VSUBS 0.006878f
C125 B.n91 VSUBS 0.006878f
C126 B.n92 VSUBS 0.006878f
C127 B.n93 VSUBS 0.017117f
C128 B.n94 VSUBS 0.006878f
C129 B.n95 VSUBS 0.006878f
C130 B.n96 VSUBS 0.006878f
C131 B.n97 VSUBS 0.006878f
C132 B.n98 VSUBS 0.006878f
C133 B.n99 VSUBS 0.006878f
C134 B.n100 VSUBS 0.006878f
C135 B.n101 VSUBS 0.006878f
C136 B.n102 VSUBS 0.006878f
C137 B.n103 VSUBS 0.006878f
C138 B.n104 VSUBS 0.006878f
C139 B.n105 VSUBS 0.006878f
C140 B.n106 VSUBS 0.006878f
C141 B.n107 VSUBS 0.006878f
C142 B.n108 VSUBS 0.006878f
C143 B.n109 VSUBS 0.006878f
C144 B.n110 VSUBS 0.006878f
C145 B.n111 VSUBS 0.006878f
C146 B.n112 VSUBS 0.006878f
C147 B.n113 VSUBS 0.006878f
C148 B.n114 VSUBS 0.006878f
C149 B.n115 VSUBS 0.006878f
C150 B.n116 VSUBS 0.006878f
C151 B.n117 VSUBS 0.006878f
C152 B.n118 VSUBS 0.006878f
C153 B.n119 VSUBS 0.006878f
C154 B.n120 VSUBS 0.006878f
C155 B.n121 VSUBS 0.006878f
C156 B.n122 VSUBS 0.006878f
C157 B.n123 VSUBS 0.006878f
C158 B.n124 VSUBS 0.006878f
C159 B.n125 VSUBS 0.006878f
C160 B.n126 VSUBS 0.006878f
C161 B.n127 VSUBS 0.006878f
C162 B.n128 VSUBS 0.006878f
C163 B.n129 VSUBS 0.006878f
C164 B.n130 VSUBS 0.006878f
C165 B.n131 VSUBS 0.006878f
C166 B.n132 VSUBS 0.006878f
C167 B.n133 VSUBS 0.006878f
C168 B.n134 VSUBS 0.006878f
C169 B.n135 VSUBS 0.006878f
C170 B.n136 VSUBS 0.006878f
C171 B.n137 VSUBS 0.006878f
C172 B.n138 VSUBS 0.006878f
C173 B.n139 VSUBS 0.006878f
C174 B.n140 VSUBS 0.006878f
C175 B.n141 VSUBS 0.006878f
C176 B.n142 VSUBS 0.006878f
C177 B.n143 VSUBS 0.016466f
C178 B.n144 VSUBS 0.006878f
C179 B.n145 VSUBS 0.006878f
C180 B.n146 VSUBS 0.006878f
C181 B.n147 VSUBS 0.006878f
C182 B.n148 VSUBS 0.006878f
C183 B.n149 VSUBS 0.006878f
C184 B.n150 VSUBS 0.006878f
C185 B.n151 VSUBS 0.006878f
C186 B.n152 VSUBS 0.006878f
C187 B.n153 VSUBS 0.006878f
C188 B.n154 VSUBS 0.006878f
C189 B.n155 VSUBS 0.006878f
C190 B.n156 VSUBS 0.006878f
C191 B.n157 VSUBS 0.006878f
C192 B.n158 VSUBS 0.006878f
C193 B.n159 VSUBS 0.006878f
C194 B.n160 VSUBS 0.006878f
C195 B.n161 VSUBS 0.006878f
C196 B.n162 VSUBS 0.006878f
C197 B.n163 VSUBS 0.006878f
C198 B.n164 VSUBS 0.006878f
C199 B.n165 VSUBS 0.006878f
C200 B.n166 VSUBS 0.006878f
C201 B.n167 VSUBS 0.006878f
C202 B.n168 VSUBS 0.006878f
C203 B.n169 VSUBS 0.006878f
C204 B.n170 VSUBS 0.006878f
C205 B.n171 VSUBS 0.006878f
C206 B.n172 VSUBS 0.004754f
C207 B.n173 VSUBS 0.006878f
C208 B.n174 VSUBS 0.006878f
C209 B.n175 VSUBS 0.006878f
C210 B.n176 VSUBS 0.006878f
C211 B.n177 VSUBS 0.006878f
C212 B.t2 VSUBS 0.333608f
C213 B.t1 VSUBS 0.36531f
C214 B.t0 VSUBS 1.89889f
C215 B.n178 VSUBS 0.557418f
C216 B.n179 VSUBS 0.31688f
C217 B.n180 VSUBS 0.006878f
C218 B.n181 VSUBS 0.006878f
C219 B.n182 VSUBS 0.006878f
C220 B.n183 VSUBS 0.006878f
C221 B.n184 VSUBS 0.006878f
C222 B.n185 VSUBS 0.006878f
C223 B.n186 VSUBS 0.006878f
C224 B.n187 VSUBS 0.006878f
C225 B.n188 VSUBS 0.006878f
C226 B.n189 VSUBS 0.006878f
C227 B.n190 VSUBS 0.006878f
C228 B.n191 VSUBS 0.006878f
C229 B.n192 VSUBS 0.006878f
C230 B.n193 VSUBS 0.006878f
C231 B.n194 VSUBS 0.006878f
C232 B.n195 VSUBS 0.006878f
C233 B.n196 VSUBS 0.006878f
C234 B.n197 VSUBS 0.006878f
C235 B.n198 VSUBS 0.006878f
C236 B.n199 VSUBS 0.006878f
C237 B.n200 VSUBS 0.006878f
C238 B.n201 VSUBS 0.006878f
C239 B.n202 VSUBS 0.006878f
C240 B.n203 VSUBS 0.006878f
C241 B.n204 VSUBS 0.006878f
C242 B.n205 VSUBS 0.006878f
C243 B.n206 VSUBS 0.006878f
C244 B.n207 VSUBS 0.006878f
C245 B.n208 VSUBS 0.016466f
C246 B.n209 VSUBS 0.006878f
C247 B.n210 VSUBS 0.006878f
C248 B.n211 VSUBS 0.006878f
C249 B.n212 VSUBS 0.006878f
C250 B.n213 VSUBS 0.006878f
C251 B.n214 VSUBS 0.006878f
C252 B.n215 VSUBS 0.006878f
C253 B.n216 VSUBS 0.006878f
C254 B.n217 VSUBS 0.006878f
C255 B.n218 VSUBS 0.006878f
C256 B.n219 VSUBS 0.006878f
C257 B.n220 VSUBS 0.006878f
C258 B.n221 VSUBS 0.006878f
C259 B.n222 VSUBS 0.006878f
C260 B.n223 VSUBS 0.006878f
C261 B.n224 VSUBS 0.006878f
C262 B.n225 VSUBS 0.006878f
C263 B.n226 VSUBS 0.006878f
C264 B.n227 VSUBS 0.006878f
C265 B.n228 VSUBS 0.006878f
C266 B.n229 VSUBS 0.006878f
C267 B.n230 VSUBS 0.006878f
C268 B.n231 VSUBS 0.006878f
C269 B.n232 VSUBS 0.006878f
C270 B.n233 VSUBS 0.006878f
C271 B.n234 VSUBS 0.006878f
C272 B.n235 VSUBS 0.006878f
C273 B.n236 VSUBS 0.006878f
C274 B.n237 VSUBS 0.006878f
C275 B.n238 VSUBS 0.006878f
C276 B.n239 VSUBS 0.006878f
C277 B.n240 VSUBS 0.006878f
C278 B.n241 VSUBS 0.006878f
C279 B.n242 VSUBS 0.006878f
C280 B.n243 VSUBS 0.006878f
C281 B.n244 VSUBS 0.006878f
C282 B.n245 VSUBS 0.006878f
C283 B.n246 VSUBS 0.006878f
C284 B.n247 VSUBS 0.006878f
C285 B.n248 VSUBS 0.006878f
C286 B.n249 VSUBS 0.006878f
C287 B.n250 VSUBS 0.006878f
C288 B.n251 VSUBS 0.006878f
C289 B.n252 VSUBS 0.006878f
C290 B.n253 VSUBS 0.006878f
C291 B.n254 VSUBS 0.006878f
C292 B.n255 VSUBS 0.006878f
C293 B.n256 VSUBS 0.006878f
C294 B.n257 VSUBS 0.006878f
C295 B.n258 VSUBS 0.006878f
C296 B.n259 VSUBS 0.006878f
C297 B.n260 VSUBS 0.006878f
C298 B.n261 VSUBS 0.006878f
C299 B.n262 VSUBS 0.006878f
C300 B.n263 VSUBS 0.006878f
C301 B.n264 VSUBS 0.006878f
C302 B.n265 VSUBS 0.006878f
C303 B.n266 VSUBS 0.006878f
C304 B.n267 VSUBS 0.006878f
C305 B.n268 VSUBS 0.006878f
C306 B.n269 VSUBS 0.006878f
C307 B.n270 VSUBS 0.006878f
C308 B.n271 VSUBS 0.006878f
C309 B.n272 VSUBS 0.006878f
C310 B.n273 VSUBS 0.006878f
C311 B.n274 VSUBS 0.006878f
C312 B.n275 VSUBS 0.006878f
C313 B.n276 VSUBS 0.006878f
C314 B.n277 VSUBS 0.006878f
C315 B.n278 VSUBS 0.006878f
C316 B.n279 VSUBS 0.006878f
C317 B.n280 VSUBS 0.006878f
C318 B.n281 VSUBS 0.006878f
C319 B.n282 VSUBS 0.006878f
C320 B.n283 VSUBS 0.006878f
C321 B.n284 VSUBS 0.006878f
C322 B.n285 VSUBS 0.006878f
C323 B.n286 VSUBS 0.006878f
C324 B.n287 VSUBS 0.006878f
C325 B.n288 VSUBS 0.006878f
C326 B.n289 VSUBS 0.006878f
C327 B.n290 VSUBS 0.006878f
C328 B.n291 VSUBS 0.006878f
C329 B.n292 VSUBS 0.006878f
C330 B.n293 VSUBS 0.006878f
C331 B.n294 VSUBS 0.006878f
C332 B.n295 VSUBS 0.006878f
C333 B.n296 VSUBS 0.006878f
C334 B.n297 VSUBS 0.006878f
C335 B.n298 VSUBS 0.006878f
C336 B.n299 VSUBS 0.006878f
C337 B.n300 VSUBS 0.006878f
C338 B.n301 VSUBS 0.006878f
C339 B.n302 VSUBS 0.006878f
C340 B.n303 VSUBS 0.016466f
C341 B.n304 VSUBS 0.017117f
C342 B.n305 VSUBS 0.017117f
C343 B.n306 VSUBS 0.006878f
C344 B.n307 VSUBS 0.006878f
C345 B.n308 VSUBS 0.006878f
C346 B.n309 VSUBS 0.006878f
C347 B.n310 VSUBS 0.006878f
C348 B.n311 VSUBS 0.006878f
C349 B.n312 VSUBS 0.006878f
C350 B.n313 VSUBS 0.006878f
C351 B.n314 VSUBS 0.006878f
C352 B.n315 VSUBS 0.006878f
C353 B.n316 VSUBS 0.006878f
C354 B.n317 VSUBS 0.006878f
C355 B.n318 VSUBS 0.006878f
C356 B.n319 VSUBS 0.006878f
C357 B.n320 VSUBS 0.006878f
C358 B.n321 VSUBS 0.006878f
C359 B.n322 VSUBS 0.006878f
C360 B.n323 VSUBS 0.006878f
C361 B.n324 VSUBS 0.006878f
C362 B.n325 VSUBS 0.006878f
C363 B.n326 VSUBS 0.006878f
C364 B.n327 VSUBS 0.006878f
C365 B.n328 VSUBS 0.006878f
C366 B.n329 VSUBS 0.006878f
C367 B.n330 VSUBS 0.006878f
C368 B.n331 VSUBS 0.006878f
C369 B.n332 VSUBS 0.006878f
C370 B.n333 VSUBS 0.006878f
C371 B.n334 VSUBS 0.006878f
C372 B.n335 VSUBS 0.006878f
C373 B.n336 VSUBS 0.006878f
C374 B.n337 VSUBS 0.006878f
C375 B.n338 VSUBS 0.006878f
C376 B.n339 VSUBS 0.006878f
C377 B.n340 VSUBS 0.006878f
C378 B.n341 VSUBS 0.006878f
C379 B.n342 VSUBS 0.006878f
C380 B.n343 VSUBS 0.006878f
C381 B.n344 VSUBS 0.006878f
C382 B.n345 VSUBS 0.006878f
C383 B.n346 VSUBS 0.006878f
C384 B.n347 VSUBS 0.006878f
C385 B.n348 VSUBS 0.006878f
C386 B.n349 VSUBS 0.006878f
C387 B.n350 VSUBS 0.006878f
C388 B.n351 VSUBS 0.006878f
C389 B.n352 VSUBS 0.006878f
C390 B.n353 VSUBS 0.006878f
C391 B.n354 VSUBS 0.006878f
C392 B.n355 VSUBS 0.006878f
C393 B.n356 VSUBS 0.006878f
C394 B.n357 VSUBS 0.006878f
C395 B.n358 VSUBS 0.006878f
C396 B.n359 VSUBS 0.006878f
C397 B.n360 VSUBS 0.006878f
C398 B.n361 VSUBS 0.006878f
C399 B.n362 VSUBS 0.006878f
C400 B.n363 VSUBS 0.006878f
C401 B.n364 VSUBS 0.006878f
C402 B.n365 VSUBS 0.006878f
C403 B.n366 VSUBS 0.006878f
C404 B.n367 VSUBS 0.006878f
C405 B.n368 VSUBS 0.006878f
C406 B.n369 VSUBS 0.006878f
C407 B.n370 VSUBS 0.006878f
C408 B.n371 VSUBS 0.006878f
C409 B.n372 VSUBS 0.006878f
C410 B.n373 VSUBS 0.006878f
C411 B.n374 VSUBS 0.006878f
C412 B.n375 VSUBS 0.006878f
C413 B.n376 VSUBS 0.006878f
C414 B.n377 VSUBS 0.006878f
C415 B.n378 VSUBS 0.006878f
C416 B.n379 VSUBS 0.006878f
C417 B.n380 VSUBS 0.006878f
C418 B.n381 VSUBS 0.006878f
C419 B.n382 VSUBS 0.006878f
C420 B.n383 VSUBS 0.006878f
C421 B.n384 VSUBS 0.006878f
C422 B.n385 VSUBS 0.006878f
C423 B.n386 VSUBS 0.006878f
C424 B.n387 VSUBS 0.006878f
C425 B.n388 VSUBS 0.006878f
C426 B.n389 VSUBS 0.006878f
C427 B.n390 VSUBS 0.004754f
C428 B.n391 VSUBS 0.015937f
C429 B.n392 VSUBS 0.005563f
C430 B.n393 VSUBS 0.006878f
C431 B.n394 VSUBS 0.006878f
C432 B.n395 VSUBS 0.006878f
C433 B.n396 VSUBS 0.006878f
C434 B.n397 VSUBS 0.006878f
C435 B.n398 VSUBS 0.006878f
C436 B.n399 VSUBS 0.006878f
C437 B.n400 VSUBS 0.006878f
C438 B.n401 VSUBS 0.006878f
C439 B.n402 VSUBS 0.006878f
C440 B.n403 VSUBS 0.006878f
C441 B.t11 VSUBS 0.333612f
C442 B.t10 VSUBS 0.365313f
C443 B.t9 VSUBS 1.89889f
C444 B.n404 VSUBS 0.557415f
C445 B.n405 VSUBS 0.316876f
C446 B.n406 VSUBS 0.015937f
C447 B.n407 VSUBS 0.005563f
C448 B.n408 VSUBS 0.006878f
C449 B.n409 VSUBS 0.006878f
C450 B.n410 VSUBS 0.006878f
C451 B.n411 VSUBS 0.006878f
C452 B.n412 VSUBS 0.006878f
C453 B.n413 VSUBS 0.006878f
C454 B.n414 VSUBS 0.006878f
C455 B.n415 VSUBS 0.006878f
C456 B.n416 VSUBS 0.006878f
C457 B.n417 VSUBS 0.006878f
C458 B.n418 VSUBS 0.006878f
C459 B.n419 VSUBS 0.006878f
C460 B.n420 VSUBS 0.006878f
C461 B.n421 VSUBS 0.006878f
C462 B.n422 VSUBS 0.006878f
C463 B.n423 VSUBS 0.006878f
C464 B.n424 VSUBS 0.006878f
C465 B.n425 VSUBS 0.006878f
C466 B.n426 VSUBS 0.006878f
C467 B.n427 VSUBS 0.006878f
C468 B.n428 VSUBS 0.006878f
C469 B.n429 VSUBS 0.006878f
C470 B.n430 VSUBS 0.006878f
C471 B.n431 VSUBS 0.006878f
C472 B.n432 VSUBS 0.006878f
C473 B.n433 VSUBS 0.006878f
C474 B.n434 VSUBS 0.006878f
C475 B.n435 VSUBS 0.006878f
C476 B.n436 VSUBS 0.006878f
C477 B.n437 VSUBS 0.006878f
C478 B.n438 VSUBS 0.006878f
C479 B.n439 VSUBS 0.006878f
C480 B.n440 VSUBS 0.006878f
C481 B.n441 VSUBS 0.006878f
C482 B.n442 VSUBS 0.006878f
C483 B.n443 VSUBS 0.006878f
C484 B.n444 VSUBS 0.006878f
C485 B.n445 VSUBS 0.006878f
C486 B.n446 VSUBS 0.006878f
C487 B.n447 VSUBS 0.006878f
C488 B.n448 VSUBS 0.006878f
C489 B.n449 VSUBS 0.006878f
C490 B.n450 VSUBS 0.006878f
C491 B.n451 VSUBS 0.006878f
C492 B.n452 VSUBS 0.006878f
C493 B.n453 VSUBS 0.006878f
C494 B.n454 VSUBS 0.006878f
C495 B.n455 VSUBS 0.006878f
C496 B.n456 VSUBS 0.006878f
C497 B.n457 VSUBS 0.006878f
C498 B.n458 VSUBS 0.006878f
C499 B.n459 VSUBS 0.006878f
C500 B.n460 VSUBS 0.006878f
C501 B.n461 VSUBS 0.006878f
C502 B.n462 VSUBS 0.006878f
C503 B.n463 VSUBS 0.006878f
C504 B.n464 VSUBS 0.006878f
C505 B.n465 VSUBS 0.006878f
C506 B.n466 VSUBS 0.006878f
C507 B.n467 VSUBS 0.006878f
C508 B.n468 VSUBS 0.006878f
C509 B.n469 VSUBS 0.006878f
C510 B.n470 VSUBS 0.006878f
C511 B.n471 VSUBS 0.006878f
C512 B.n472 VSUBS 0.006878f
C513 B.n473 VSUBS 0.006878f
C514 B.n474 VSUBS 0.006878f
C515 B.n475 VSUBS 0.006878f
C516 B.n476 VSUBS 0.006878f
C517 B.n477 VSUBS 0.006878f
C518 B.n478 VSUBS 0.006878f
C519 B.n479 VSUBS 0.006878f
C520 B.n480 VSUBS 0.006878f
C521 B.n481 VSUBS 0.006878f
C522 B.n482 VSUBS 0.006878f
C523 B.n483 VSUBS 0.006878f
C524 B.n484 VSUBS 0.006878f
C525 B.n485 VSUBS 0.006878f
C526 B.n486 VSUBS 0.006878f
C527 B.n487 VSUBS 0.006878f
C528 B.n488 VSUBS 0.006878f
C529 B.n489 VSUBS 0.006878f
C530 B.n490 VSUBS 0.006878f
C531 B.n491 VSUBS 0.006878f
C532 B.n492 VSUBS 0.006878f
C533 B.n493 VSUBS 0.006878f
C534 B.n494 VSUBS 0.017117f
C535 B.n495 VSUBS 0.016355f
C536 B.n496 VSUBS 0.017229f
C537 B.n497 VSUBS 0.006878f
C538 B.n498 VSUBS 0.006878f
C539 B.n499 VSUBS 0.006878f
C540 B.n500 VSUBS 0.006878f
C541 B.n501 VSUBS 0.006878f
C542 B.n502 VSUBS 0.006878f
C543 B.n503 VSUBS 0.006878f
C544 B.n504 VSUBS 0.006878f
C545 B.n505 VSUBS 0.006878f
C546 B.n506 VSUBS 0.006878f
C547 B.n507 VSUBS 0.006878f
C548 B.n508 VSUBS 0.006878f
C549 B.n509 VSUBS 0.006878f
C550 B.n510 VSUBS 0.006878f
C551 B.n511 VSUBS 0.006878f
C552 B.n512 VSUBS 0.006878f
C553 B.n513 VSUBS 0.006878f
C554 B.n514 VSUBS 0.006878f
C555 B.n515 VSUBS 0.006878f
C556 B.n516 VSUBS 0.006878f
C557 B.n517 VSUBS 0.006878f
C558 B.n518 VSUBS 0.006878f
C559 B.n519 VSUBS 0.006878f
C560 B.n520 VSUBS 0.006878f
C561 B.n521 VSUBS 0.006878f
C562 B.n522 VSUBS 0.006878f
C563 B.n523 VSUBS 0.006878f
C564 B.n524 VSUBS 0.006878f
C565 B.n525 VSUBS 0.006878f
C566 B.n526 VSUBS 0.006878f
C567 B.n527 VSUBS 0.006878f
C568 B.n528 VSUBS 0.006878f
C569 B.n529 VSUBS 0.006878f
C570 B.n530 VSUBS 0.006878f
C571 B.n531 VSUBS 0.006878f
C572 B.n532 VSUBS 0.006878f
C573 B.n533 VSUBS 0.006878f
C574 B.n534 VSUBS 0.006878f
C575 B.n535 VSUBS 0.006878f
C576 B.n536 VSUBS 0.006878f
C577 B.n537 VSUBS 0.006878f
C578 B.n538 VSUBS 0.006878f
C579 B.n539 VSUBS 0.006878f
C580 B.n540 VSUBS 0.006878f
C581 B.n541 VSUBS 0.006878f
C582 B.n542 VSUBS 0.006878f
C583 B.n543 VSUBS 0.006878f
C584 B.n544 VSUBS 0.006878f
C585 B.n545 VSUBS 0.006878f
C586 B.n546 VSUBS 0.006878f
C587 B.n547 VSUBS 0.006878f
C588 B.n548 VSUBS 0.006878f
C589 B.n549 VSUBS 0.006878f
C590 B.n550 VSUBS 0.006878f
C591 B.n551 VSUBS 0.006878f
C592 B.n552 VSUBS 0.006878f
C593 B.n553 VSUBS 0.006878f
C594 B.n554 VSUBS 0.006878f
C595 B.n555 VSUBS 0.006878f
C596 B.n556 VSUBS 0.006878f
C597 B.n557 VSUBS 0.006878f
C598 B.n558 VSUBS 0.006878f
C599 B.n559 VSUBS 0.006878f
C600 B.n560 VSUBS 0.006878f
C601 B.n561 VSUBS 0.006878f
C602 B.n562 VSUBS 0.006878f
C603 B.n563 VSUBS 0.006878f
C604 B.n564 VSUBS 0.006878f
C605 B.n565 VSUBS 0.006878f
C606 B.n566 VSUBS 0.006878f
C607 B.n567 VSUBS 0.006878f
C608 B.n568 VSUBS 0.006878f
C609 B.n569 VSUBS 0.006878f
C610 B.n570 VSUBS 0.006878f
C611 B.n571 VSUBS 0.006878f
C612 B.n572 VSUBS 0.006878f
C613 B.n573 VSUBS 0.006878f
C614 B.n574 VSUBS 0.006878f
C615 B.n575 VSUBS 0.006878f
C616 B.n576 VSUBS 0.006878f
C617 B.n577 VSUBS 0.006878f
C618 B.n578 VSUBS 0.006878f
C619 B.n579 VSUBS 0.006878f
C620 B.n580 VSUBS 0.006878f
C621 B.n581 VSUBS 0.006878f
C622 B.n582 VSUBS 0.006878f
C623 B.n583 VSUBS 0.006878f
C624 B.n584 VSUBS 0.006878f
C625 B.n585 VSUBS 0.006878f
C626 B.n586 VSUBS 0.006878f
C627 B.n587 VSUBS 0.006878f
C628 B.n588 VSUBS 0.006878f
C629 B.n589 VSUBS 0.006878f
C630 B.n590 VSUBS 0.006878f
C631 B.n591 VSUBS 0.006878f
C632 B.n592 VSUBS 0.006878f
C633 B.n593 VSUBS 0.006878f
C634 B.n594 VSUBS 0.006878f
C635 B.n595 VSUBS 0.006878f
C636 B.n596 VSUBS 0.006878f
C637 B.n597 VSUBS 0.006878f
C638 B.n598 VSUBS 0.006878f
C639 B.n599 VSUBS 0.006878f
C640 B.n600 VSUBS 0.006878f
C641 B.n601 VSUBS 0.006878f
C642 B.n602 VSUBS 0.006878f
C643 B.n603 VSUBS 0.006878f
C644 B.n604 VSUBS 0.006878f
C645 B.n605 VSUBS 0.006878f
C646 B.n606 VSUBS 0.006878f
C647 B.n607 VSUBS 0.006878f
C648 B.n608 VSUBS 0.006878f
C649 B.n609 VSUBS 0.006878f
C650 B.n610 VSUBS 0.006878f
C651 B.n611 VSUBS 0.006878f
C652 B.n612 VSUBS 0.006878f
C653 B.n613 VSUBS 0.006878f
C654 B.n614 VSUBS 0.006878f
C655 B.n615 VSUBS 0.006878f
C656 B.n616 VSUBS 0.006878f
C657 B.n617 VSUBS 0.006878f
C658 B.n618 VSUBS 0.006878f
C659 B.n619 VSUBS 0.006878f
C660 B.n620 VSUBS 0.006878f
C661 B.n621 VSUBS 0.006878f
C662 B.n622 VSUBS 0.006878f
C663 B.n623 VSUBS 0.006878f
C664 B.n624 VSUBS 0.006878f
C665 B.n625 VSUBS 0.006878f
C666 B.n626 VSUBS 0.006878f
C667 B.n627 VSUBS 0.006878f
C668 B.n628 VSUBS 0.006878f
C669 B.n629 VSUBS 0.006878f
C670 B.n630 VSUBS 0.006878f
C671 B.n631 VSUBS 0.006878f
C672 B.n632 VSUBS 0.006878f
C673 B.n633 VSUBS 0.006878f
C674 B.n634 VSUBS 0.006878f
C675 B.n635 VSUBS 0.006878f
C676 B.n636 VSUBS 0.006878f
C677 B.n637 VSUBS 0.006878f
C678 B.n638 VSUBS 0.006878f
C679 B.n639 VSUBS 0.006878f
C680 B.n640 VSUBS 0.006878f
C681 B.n641 VSUBS 0.006878f
C682 B.n642 VSUBS 0.006878f
C683 B.n643 VSUBS 0.006878f
C684 B.n644 VSUBS 0.016466f
C685 B.n645 VSUBS 0.016466f
C686 B.n646 VSUBS 0.017117f
C687 B.n647 VSUBS 0.006878f
C688 B.n648 VSUBS 0.006878f
C689 B.n649 VSUBS 0.006878f
C690 B.n650 VSUBS 0.006878f
C691 B.n651 VSUBS 0.006878f
C692 B.n652 VSUBS 0.006878f
C693 B.n653 VSUBS 0.006878f
C694 B.n654 VSUBS 0.006878f
C695 B.n655 VSUBS 0.006878f
C696 B.n656 VSUBS 0.006878f
C697 B.n657 VSUBS 0.006878f
C698 B.n658 VSUBS 0.006878f
C699 B.n659 VSUBS 0.006878f
C700 B.n660 VSUBS 0.006878f
C701 B.n661 VSUBS 0.006878f
C702 B.n662 VSUBS 0.006878f
C703 B.n663 VSUBS 0.006878f
C704 B.n664 VSUBS 0.006878f
C705 B.n665 VSUBS 0.006878f
C706 B.n666 VSUBS 0.006878f
C707 B.n667 VSUBS 0.006878f
C708 B.n668 VSUBS 0.006878f
C709 B.n669 VSUBS 0.006878f
C710 B.n670 VSUBS 0.006878f
C711 B.n671 VSUBS 0.006878f
C712 B.n672 VSUBS 0.006878f
C713 B.n673 VSUBS 0.006878f
C714 B.n674 VSUBS 0.006878f
C715 B.n675 VSUBS 0.006878f
C716 B.n676 VSUBS 0.006878f
C717 B.n677 VSUBS 0.006878f
C718 B.n678 VSUBS 0.006878f
C719 B.n679 VSUBS 0.006878f
C720 B.n680 VSUBS 0.006878f
C721 B.n681 VSUBS 0.006878f
C722 B.n682 VSUBS 0.006878f
C723 B.n683 VSUBS 0.006878f
C724 B.n684 VSUBS 0.006878f
C725 B.n685 VSUBS 0.006878f
C726 B.n686 VSUBS 0.006878f
C727 B.n687 VSUBS 0.006878f
C728 B.n688 VSUBS 0.006878f
C729 B.n689 VSUBS 0.006878f
C730 B.n690 VSUBS 0.006878f
C731 B.n691 VSUBS 0.006878f
C732 B.n692 VSUBS 0.006878f
C733 B.n693 VSUBS 0.006878f
C734 B.n694 VSUBS 0.006878f
C735 B.n695 VSUBS 0.006878f
C736 B.n696 VSUBS 0.006878f
C737 B.n697 VSUBS 0.006878f
C738 B.n698 VSUBS 0.006878f
C739 B.n699 VSUBS 0.006878f
C740 B.n700 VSUBS 0.006878f
C741 B.n701 VSUBS 0.006878f
C742 B.n702 VSUBS 0.006878f
C743 B.n703 VSUBS 0.006878f
C744 B.n704 VSUBS 0.006878f
C745 B.n705 VSUBS 0.006878f
C746 B.n706 VSUBS 0.006878f
C747 B.n707 VSUBS 0.006878f
C748 B.n708 VSUBS 0.006878f
C749 B.n709 VSUBS 0.006878f
C750 B.n710 VSUBS 0.006878f
C751 B.n711 VSUBS 0.006878f
C752 B.n712 VSUBS 0.006878f
C753 B.n713 VSUBS 0.006878f
C754 B.n714 VSUBS 0.006878f
C755 B.n715 VSUBS 0.006878f
C756 B.n716 VSUBS 0.006878f
C757 B.n717 VSUBS 0.006878f
C758 B.n718 VSUBS 0.006878f
C759 B.n719 VSUBS 0.006878f
C760 B.n720 VSUBS 0.006878f
C761 B.n721 VSUBS 0.006878f
C762 B.n722 VSUBS 0.006878f
C763 B.n723 VSUBS 0.006878f
C764 B.n724 VSUBS 0.006878f
C765 B.n725 VSUBS 0.006878f
C766 B.n726 VSUBS 0.006878f
C767 B.n727 VSUBS 0.006878f
C768 B.n728 VSUBS 0.006878f
C769 B.n729 VSUBS 0.006878f
C770 B.n730 VSUBS 0.006878f
C771 B.n731 VSUBS 0.004754f
C772 B.n732 VSUBS 0.006878f
C773 B.n733 VSUBS 0.006878f
C774 B.n734 VSUBS 0.005563f
C775 B.n735 VSUBS 0.006878f
C776 B.n736 VSUBS 0.006878f
C777 B.n737 VSUBS 0.006878f
C778 B.n738 VSUBS 0.006878f
C779 B.n739 VSUBS 0.006878f
C780 B.n740 VSUBS 0.006878f
C781 B.n741 VSUBS 0.006878f
C782 B.n742 VSUBS 0.006878f
C783 B.n743 VSUBS 0.006878f
C784 B.n744 VSUBS 0.006878f
C785 B.n745 VSUBS 0.006878f
C786 B.n746 VSUBS 0.005563f
C787 B.n747 VSUBS 0.015937f
C788 B.n748 VSUBS 0.004754f
C789 B.n749 VSUBS 0.006878f
C790 B.n750 VSUBS 0.006878f
C791 B.n751 VSUBS 0.006878f
C792 B.n752 VSUBS 0.006878f
C793 B.n753 VSUBS 0.006878f
C794 B.n754 VSUBS 0.006878f
C795 B.n755 VSUBS 0.006878f
C796 B.n756 VSUBS 0.006878f
C797 B.n757 VSUBS 0.006878f
C798 B.n758 VSUBS 0.006878f
C799 B.n759 VSUBS 0.006878f
C800 B.n760 VSUBS 0.006878f
C801 B.n761 VSUBS 0.006878f
C802 B.n762 VSUBS 0.006878f
C803 B.n763 VSUBS 0.006878f
C804 B.n764 VSUBS 0.006878f
C805 B.n765 VSUBS 0.006878f
C806 B.n766 VSUBS 0.006878f
C807 B.n767 VSUBS 0.006878f
C808 B.n768 VSUBS 0.006878f
C809 B.n769 VSUBS 0.006878f
C810 B.n770 VSUBS 0.006878f
C811 B.n771 VSUBS 0.006878f
C812 B.n772 VSUBS 0.006878f
C813 B.n773 VSUBS 0.006878f
C814 B.n774 VSUBS 0.006878f
C815 B.n775 VSUBS 0.006878f
C816 B.n776 VSUBS 0.006878f
C817 B.n777 VSUBS 0.006878f
C818 B.n778 VSUBS 0.006878f
C819 B.n779 VSUBS 0.006878f
C820 B.n780 VSUBS 0.006878f
C821 B.n781 VSUBS 0.006878f
C822 B.n782 VSUBS 0.006878f
C823 B.n783 VSUBS 0.006878f
C824 B.n784 VSUBS 0.006878f
C825 B.n785 VSUBS 0.006878f
C826 B.n786 VSUBS 0.006878f
C827 B.n787 VSUBS 0.006878f
C828 B.n788 VSUBS 0.006878f
C829 B.n789 VSUBS 0.006878f
C830 B.n790 VSUBS 0.006878f
C831 B.n791 VSUBS 0.006878f
C832 B.n792 VSUBS 0.006878f
C833 B.n793 VSUBS 0.006878f
C834 B.n794 VSUBS 0.006878f
C835 B.n795 VSUBS 0.006878f
C836 B.n796 VSUBS 0.006878f
C837 B.n797 VSUBS 0.006878f
C838 B.n798 VSUBS 0.006878f
C839 B.n799 VSUBS 0.006878f
C840 B.n800 VSUBS 0.006878f
C841 B.n801 VSUBS 0.006878f
C842 B.n802 VSUBS 0.006878f
C843 B.n803 VSUBS 0.006878f
C844 B.n804 VSUBS 0.006878f
C845 B.n805 VSUBS 0.006878f
C846 B.n806 VSUBS 0.006878f
C847 B.n807 VSUBS 0.006878f
C848 B.n808 VSUBS 0.006878f
C849 B.n809 VSUBS 0.006878f
C850 B.n810 VSUBS 0.006878f
C851 B.n811 VSUBS 0.006878f
C852 B.n812 VSUBS 0.006878f
C853 B.n813 VSUBS 0.006878f
C854 B.n814 VSUBS 0.006878f
C855 B.n815 VSUBS 0.006878f
C856 B.n816 VSUBS 0.006878f
C857 B.n817 VSUBS 0.006878f
C858 B.n818 VSUBS 0.006878f
C859 B.n819 VSUBS 0.006878f
C860 B.n820 VSUBS 0.006878f
C861 B.n821 VSUBS 0.006878f
C862 B.n822 VSUBS 0.006878f
C863 B.n823 VSUBS 0.006878f
C864 B.n824 VSUBS 0.006878f
C865 B.n825 VSUBS 0.006878f
C866 B.n826 VSUBS 0.006878f
C867 B.n827 VSUBS 0.006878f
C868 B.n828 VSUBS 0.006878f
C869 B.n829 VSUBS 0.006878f
C870 B.n830 VSUBS 0.006878f
C871 B.n831 VSUBS 0.006878f
C872 B.n832 VSUBS 0.006878f
C873 B.n833 VSUBS 0.017117f
C874 B.n834 VSUBS 0.017117f
C875 B.n835 VSUBS 0.016466f
C876 B.n836 VSUBS 0.006878f
C877 B.n837 VSUBS 0.006878f
C878 B.n838 VSUBS 0.006878f
C879 B.n839 VSUBS 0.006878f
C880 B.n840 VSUBS 0.006878f
C881 B.n841 VSUBS 0.006878f
C882 B.n842 VSUBS 0.006878f
C883 B.n843 VSUBS 0.006878f
C884 B.n844 VSUBS 0.006878f
C885 B.n845 VSUBS 0.006878f
C886 B.n846 VSUBS 0.006878f
C887 B.n847 VSUBS 0.006878f
C888 B.n848 VSUBS 0.006878f
C889 B.n849 VSUBS 0.006878f
C890 B.n850 VSUBS 0.006878f
C891 B.n851 VSUBS 0.006878f
C892 B.n852 VSUBS 0.006878f
C893 B.n853 VSUBS 0.006878f
C894 B.n854 VSUBS 0.006878f
C895 B.n855 VSUBS 0.006878f
C896 B.n856 VSUBS 0.006878f
C897 B.n857 VSUBS 0.006878f
C898 B.n858 VSUBS 0.006878f
C899 B.n859 VSUBS 0.006878f
C900 B.n860 VSUBS 0.006878f
C901 B.n861 VSUBS 0.006878f
C902 B.n862 VSUBS 0.006878f
C903 B.n863 VSUBS 0.006878f
C904 B.n864 VSUBS 0.006878f
C905 B.n865 VSUBS 0.006878f
C906 B.n866 VSUBS 0.006878f
C907 B.n867 VSUBS 0.006878f
C908 B.n868 VSUBS 0.006878f
C909 B.n869 VSUBS 0.006878f
C910 B.n870 VSUBS 0.006878f
C911 B.n871 VSUBS 0.006878f
C912 B.n872 VSUBS 0.006878f
C913 B.n873 VSUBS 0.006878f
C914 B.n874 VSUBS 0.006878f
C915 B.n875 VSUBS 0.006878f
C916 B.n876 VSUBS 0.006878f
C917 B.n877 VSUBS 0.006878f
C918 B.n878 VSUBS 0.006878f
C919 B.n879 VSUBS 0.006878f
C920 B.n880 VSUBS 0.006878f
C921 B.n881 VSUBS 0.006878f
C922 B.n882 VSUBS 0.006878f
C923 B.n883 VSUBS 0.006878f
C924 B.n884 VSUBS 0.006878f
C925 B.n885 VSUBS 0.006878f
C926 B.n886 VSUBS 0.006878f
C927 B.n887 VSUBS 0.006878f
C928 B.n888 VSUBS 0.006878f
C929 B.n889 VSUBS 0.006878f
C930 B.n890 VSUBS 0.006878f
C931 B.n891 VSUBS 0.006878f
C932 B.n892 VSUBS 0.006878f
C933 B.n893 VSUBS 0.006878f
C934 B.n894 VSUBS 0.006878f
C935 B.n895 VSUBS 0.006878f
C936 B.n896 VSUBS 0.006878f
C937 B.n897 VSUBS 0.006878f
C938 B.n898 VSUBS 0.006878f
C939 B.n899 VSUBS 0.006878f
C940 B.n900 VSUBS 0.006878f
C941 B.n901 VSUBS 0.006878f
C942 B.n902 VSUBS 0.006878f
C943 B.n903 VSUBS 0.006878f
C944 B.n904 VSUBS 0.006878f
C945 B.n905 VSUBS 0.006878f
C946 B.n906 VSUBS 0.006878f
C947 B.n907 VSUBS 0.008976f
C948 B.n908 VSUBS 0.009562f
C949 B.n909 VSUBS 0.019015f
C950 VDD2.t0 VSUBS 0.37043f
C951 VDD2.t2 VSUBS 0.37043f
C952 VDD2.n0 VSUBS 3.08035f
C953 VDD2.t4 VSUBS 0.37043f
C954 VDD2.t5 VSUBS 0.37043f
C955 VDD2.n1 VSUBS 3.08035f
C956 VDD2.n2 VSUBS 4.41685f
C957 VDD2.t7 VSUBS 0.37043f
C958 VDD2.t6 VSUBS 0.37043f
C959 VDD2.n3 VSUBS 3.06636f
C960 VDD2.n4 VSUBS 3.87013f
C961 VDD2.t3 VSUBS 0.37043f
C962 VDD2.t1 VSUBS 0.37043f
C963 VDD2.n5 VSUBS 3.0803f
C964 VN.n0 VSUBS 0.035558f
C965 VN.t2 VSUBS 3.23484f
C966 VN.n1 VSUBS 0.033985f
C967 VN.n2 VSUBS 0.026973f
C968 VN.t3 VSUBS 3.23484f
C969 VN.n3 VSUBS 1.12388f
C970 VN.n4 VSUBS 0.026973f
C971 VN.n5 VSUBS 0.053325f
C972 VN.t7 VSUBS 3.4498f
C973 VN.n6 VSUBS 1.17303f
C974 VN.t5 VSUBS 3.23484f
C975 VN.n7 VSUBS 1.2081f
C976 VN.n8 VSUBS 0.045573f
C977 VN.n9 VSUBS 0.257716f
C978 VN.n10 VSUBS 0.026973f
C979 VN.n11 VSUBS 0.026973f
C980 VN.n12 VSUBS 0.021785f
C981 VN.n13 VSUBS 0.053325f
C982 VN.n14 VSUBS 0.045573f
C983 VN.n15 VSUBS 0.026973f
C984 VN.n16 VSUBS 0.026973f
C985 VN.n17 VSUBS 0.02977f
C986 VN.n18 VSUBS 0.050018f
C987 VN.n19 VSUBS 0.044432f
C988 VN.n20 VSUBS 0.026973f
C989 VN.n21 VSUBS 0.026973f
C990 VN.n22 VSUBS 0.026973f
C991 VN.n23 VSUBS 0.050018f
C992 VN.n24 VSUBS 0.036684f
C993 VN.n25 VSUBS 1.21172f
C994 VN.n26 VSUBS 0.04208f
C995 VN.n27 VSUBS 0.035558f
C996 VN.t0 VSUBS 3.23484f
C997 VN.n28 VSUBS 0.033985f
C998 VN.n29 VSUBS 0.026973f
C999 VN.t1 VSUBS 3.23484f
C1000 VN.n30 VSUBS 1.12388f
C1001 VN.n31 VSUBS 0.026973f
C1002 VN.n32 VSUBS 0.053325f
C1003 VN.t6 VSUBS 3.4498f
C1004 VN.n33 VSUBS 1.17303f
C1005 VN.t4 VSUBS 3.23484f
C1006 VN.n34 VSUBS 1.2081f
C1007 VN.n35 VSUBS 0.045573f
C1008 VN.n36 VSUBS 0.257716f
C1009 VN.n37 VSUBS 0.026973f
C1010 VN.n38 VSUBS 0.026973f
C1011 VN.n39 VSUBS 0.021785f
C1012 VN.n40 VSUBS 0.053325f
C1013 VN.n41 VSUBS 0.045573f
C1014 VN.n42 VSUBS 0.026973f
C1015 VN.n43 VSUBS 0.026973f
C1016 VN.n44 VSUBS 0.02977f
C1017 VN.n45 VSUBS 0.050018f
C1018 VN.n46 VSUBS 0.044432f
C1019 VN.n47 VSUBS 0.026973f
C1020 VN.n48 VSUBS 0.026973f
C1021 VN.n49 VSUBS 0.026973f
C1022 VN.n50 VSUBS 0.050018f
C1023 VN.n51 VSUBS 0.036684f
C1024 VN.n52 VSUBS 1.21172f
C1025 VN.n53 VSUBS 1.71488f
C1026 VTAIL.t6 VSUBS 0.326723f
C1027 VTAIL.t0 VSUBS 0.326723f
C1028 VTAIL.n0 VSUBS 2.55802f
C1029 VTAIL.n1 VSUBS 0.76805f
C1030 VTAIL.n2 VSUBS 0.025431f
C1031 VTAIL.n3 VSUBS 0.023599f
C1032 VTAIL.n4 VSUBS 0.012681f
C1033 VTAIL.n5 VSUBS 0.029973f
C1034 VTAIL.n6 VSUBS 0.013427f
C1035 VTAIL.n7 VSUBS 0.023599f
C1036 VTAIL.n8 VSUBS 0.012681f
C1037 VTAIL.n9 VSUBS 0.029973f
C1038 VTAIL.n10 VSUBS 0.013054f
C1039 VTAIL.n11 VSUBS 0.023599f
C1040 VTAIL.n12 VSUBS 0.013427f
C1041 VTAIL.n13 VSUBS 0.029973f
C1042 VTAIL.n14 VSUBS 0.013427f
C1043 VTAIL.n15 VSUBS 0.023599f
C1044 VTAIL.n16 VSUBS 0.012681f
C1045 VTAIL.n17 VSUBS 0.029973f
C1046 VTAIL.n18 VSUBS 0.013427f
C1047 VTAIL.n19 VSUBS 0.023599f
C1048 VTAIL.n20 VSUBS 0.012681f
C1049 VTAIL.n21 VSUBS 0.029973f
C1050 VTAIL.n22 VSUBS 0.013427f
C1051 VTAIL.n23 VSUBS 0.023599f
C1052 VTAIL.n24 VSUBS 0.012681f
C1053 VTAIL.n25 VSUBS 0.029973f
C1054 VTAIL.n26 VSUBS 0.013427f
C1055 VTAIL.n27 VSUBS 0.023599f
C1056 VTAIL.n28 VSUBS 0.012681f
C1057 VTAIL.n29 VSUBS 0.029973f
C1058 VTAIL.n30 VSUBS 0.013427f
C1059 VTAIL.n31 VSUBS 1.77681f
C1060 VTAIL.n32 VSUBS 0.012681f
C1061 VTAIL.t7 VSUBS 0.064315f
C1062 VTAIL.n33 VSUBS 0.183893f
C1063 VTAIL.n34 VSUBS 0.019068f
C1064 VTAIL.n35 VSUBS 0.02248f
C1065 VTAIL.n36 VSUBS 0.029973f
C1066 VTAIL.n37 VSUBS 0.013427f
C1067 VTAIL.n38 VSUBS 0.012681f
C1068 VTAIL.n39 VSUBS 0.023599f
C1069 VTAIL.n40 VSUBS 0.023599f
C1070 VTAIL.n41 VSUBS 0.012681f
C1071 VTAIL.n42 VSUBS 0.013427f
C1072 VTAIL.n43 VSUBS 0.029973f
C1073 VTAIL.n44 VSUBS 0.029973f
C1074 VTAIL.n45 VSUBS 0.013427f
C1075 VTAIL.n46 VSUBS 0.012681f
C1076 VTAIL.n47 VSUBS 0.023599f
C1077 VTAIL.n48 VSUBS 0.023599f
C1078 VTAIL.n49 VSUBS 0.012681f
C1079 VTAIL.n50 VSUBS 0.013427f
C1080 VTAIL.n51 VSUBS 0.029973f
C1081 VTAIL.n52 VSUBS 0.029973f
C1082 VTAIL.n53 VSUBS 0.013427f
C1083 VTAIL.n54 VSUBS 0.012681f
C1084 VTAIL.n55 VSUBS 0.023599f
C1085 VTAIL.n56 VSUBS 0.023599f
C1086 VTAIL.n57 VSUBS 0.012681f
C1087 VTAIL.n58 VSUBS 0.013427f
C1088 VTAIL.n59 VSUBS 0.029973f
C1089 VTAIL.n60 VSUBS 0.029973f
C1090 VTAIL.n61 VSUBS 0.013427f
C1091 VTAIL.n62 VSUBS 0.012681f
C1092 VTAIL.n63 VSUBS 0.023599f
C1093 VTAIL.n64 VSUBS 0.023599f
C1094 VTAIL.n65 VSUBS 0.012681f
C1095 VTAIL.n66 VSUBS 0.013427f
C1096 VTAIL.n67 VSUBS 0.029973f
C1097 VTAIL.n68 VSUBS 0.029973f
C1098 VTAIL.n69 VSUBS 0.013427f
C1099 VTAIL.n70 VSUBS 0.012681f
C1100 VTAIL.n71 VSUBS 0.023599f
C1101 VTAIL.n72 VSUBS 0.023599f
C1102 VTAIL.n73 VSUBS 0.012681f
C1103 VTAIL.n74 VSUBS 0.012681f
C1104 VTAIL.n75 VSUBS 0.013427f
C1105 VTAIL.n76 VSUBS 0.029973f
C1106 VTAIL.n77 VSUBS 0.029973f
C1107 VTAIL.n78 VSUBS 0.029973f
C1108 VTAIL.n79 VSUBS 0.013054f
C1109 VTAIL.n80 VSUBS 0.012681f
C1110 VTAIL.n81 VSUBS 0.023599f
C1111 VTAIL.n82 VSUBS 0.023599f
C1112 VTAIL.n83 VSUBS 0.012681f
C1113 VTAIL.n84 VSUBS 0.013427f
C1114 VTAIL.n85 VSUBS 0.029973f
C1115 VTAIL.n86 VSUBS 0.029973f
C1116 VTAIL.n87 VSUBS 0.013427f
C1117 VTAIL.n88 VSUBS 0.012681f
C1118 VTAIL.n89 VSUBS 0.023599f
C1119 VTAIL.n90 VSUBS 0.023599f
C1120 VTAIL.n91 VSUBS 0.012681f
C1121 VTAIL.n92 VSUBS 0.013427f
C1122 VTAIL.n93 VSUBS 0.029973f
C1123 VTAIL.n94 VSUBS 0.070863f
C1124 VTAIL.n95 VSUBS 0.013427f
C1125 VTAIL.n96 VSUBS 0.012681f
C1126 VTAIL.n97 VSUBS 0.054548f
C1127 VTAIL.n98 VSUBS 0.035561f
C1128 VTAIL.n99 VSUBS 0.240739f
C1129 VTAIL.n100 VSUBS 0.025431f
C1130 VTAIL.n101 VSUBS 0.023599f
C1131 VTAIL.n102 VSUBS 0.012681f
C1132 VTAIL.n103 VSUBS 0.029973f
C1133 VTAIL.n104 VSUBS 0.013427f
C1134 VTAIL.n105 VSUBS 0.023599f
C1135 VTAIL.n106 VSUBS 0.012681f
C1136 VTAIL.n107 VSUBS 0.029973f
C1137 VTAIL.n108 VSUBS 0.013054f
C1138 VTAIL.n109 VSUBS 0.023599f
C1139 VTAIL.n110 VSUBS 0.013427f
C1140 VTAIL.n111 VSUBS 0.029973f
C1141 VTAIL.n112 VSUBS 0.013427f
C1142 VTAIL.n113 VSUBS 0.023599f
C1143 VTAIL.n114 VSUBS 0.012681f
C1144 VTAIL.n115 VSUBS 0.029973f
C1145 VTAIL.n116 VSUBS 0.013427f
C1146 VTAIL.n117 VSUBS 0.023599f
C1147 VTAIL.n118 VSUBS 0.012681f
C1148 VTAIL.n119 VSUBS 0.029973f
C1149 VTAIL.n120 VSUBS 0.013427f
C1150 VTAIL.n121 VSUBS 0.023599f
C1151 VTAIL.n122 VSUBS 0.012681f
C1152 VTAIL.n123 VSUBS 0.029973f
C1153 VTAIL.n124 VSUBS 0.013427f
C1154 VTAIL.n125 VSUBS 0.023599f
C1155 VTAIL.n126 VSUBS 0.012681f
C1156 VTAIL.n127 VSUBS 0.029973f
C1157 VTAIL.n128 VSUBS 0.013427f
C1158 VTAIL.n129 VSUBS 1.77681f
C1159 VTAIL.n130 VSUBS 0.012681f
C1160 VTAIL.t9 VSUBS 0.064315f
C1161 VTAIL.n131 VSUBS 0.183893f
C1162 VTAIL.n132 VSUBS 0.019068f
C1163 VTAIL.n133 VSUBS 0.02248f
C1164 VTAIL.n134 VSUBS 0.029973f
C1165 VTAIL.n135 VSUBS 0.013427f
C1166 VTAIL.n136 VSUBS 0.012681f
C1167 VTAIL.n137 VSUBS 0.023599f
C1168 VTAIL.n138 VSUBS 0.023599f
C1169 VTAIL.n139 VSUBS 0.012681f
C1170 VTAIL.n140 VSUBS 0.013427f
C1171 VTAIL.n141 VSUBS 0.029973f
C1172 VTAIL.n142 VSUBS 0.029973f
C1173 VTAIL.n143 VSUBS 0.013427f
C1174 VTAIL.n144 VSUBS 0.012681f
C1175 VTAIL.n145 VSUBS 0.023599f
C1176 VTAIL.n146 VSUBS 0.023599f
C1177 VTAIL.n147 VSUBS 0.012681f
C1178 VTAIL.n148 VSUBS 0.013427f
C1179 VTAIL.n149 VSUBS 0.029973f
C1180 VTAIL.n150 VSUBS 0.029973f
C1181 VTAIL.n151 VSUBS 0.013427f
C1182 VTAIL.n152 VSUBS 0.012681f
C1183 VTAIL.n153 VSUBS 0.023599f
C1184 VTAIL.n154 VSUBS 0.023599f
C1185 VTAIL.n155 VSUBS 0.012681f
C1186 VTAIL.n156 VSUBS 0.013427f
C1187 VTAIL.n157 VSUBS 0.029973f
C1188 VTAIL.n158 VSUBS 0.029973f
C1189 VTAIL.n159 VSUBS 0.013427f
C1190 VTAIL.n160 VSUBS 0.012681f
C1191 VTAIL.n161 VSUBS 0.023599f
C1192 VTAIL.n162 VSUBS 0.023599f
C1193 VTAIL.n163 VSUBS 0.012681f
C1194 VTAIL.n164 VSUBS 0.013427f
C1195 VTAIL.n165 VSUBS 0.029973f
C1196 VTAIL.n166 VSUBS 0.029973f
C1197 VTAIL.n167 VSUBS 0.013427f
C1198 VTAIL.n168 VSUBS 0.012681f
C1199 VTAIL.n169 VSUBS 0.023599f
C1200 VTAIL.n170 VSUBS 0.023599f
C1201 VTAIL.n171 VSUBS 0.012681f
C1202 VTAIL.n172 VSUBS 0.012681f
C1203 VTAIL.n173 VSUBS 0.013427f
C1204 VTAIL.n174 VSUBS 0.029973f
C1205 VTAIL.n175 VSUBS 0.029973f
C1206 VTAIL.n176 VSUBS 0.029973f
C1207 VTAIL.n177 VSUBS 0.013054f
C1208 VTAIL.n178 VSUBS 0.012681f
C1209 VTAIL.n179 VSUBS 0.023599f
C1210 VTAIL.n180 VSUBS 0.023599f
C1211 VTAIL.n181 VSUBS 0.012681f
C1212 VTAIL.n182 VSUBS 0.013427f
C1213 VTAIL.n183 VSUBS 0.029973f
C1214 VTAIL.n184 VSUBS 0.029973f
C1215 VTAIL.n185 VSUBS 0.013427f
C1216 VTAIL.n186 VSUBS 0.012681f
C1217 VTAIL.n187 VSUBS 0.023599f
C1218 VTAIL.n188 VSUBS 0.023599f
C1219 VTAIL.n189 VSUBS 0.012681f
C1220 VTAIL.n190 VSUBS 0.013427f
C1221 VTAIL.n191 VSUBS 0.029973f
C1222 VTAIL.n192 VSUBS 0.070863f
C1223 VTAIL.n193 VSUBS 0.013427f
C1224 VTAIL.n194 VSUBS 0.012681f
C1225 VTAIL.n195 VSUBS 0.054548f
C1226 VTAIL.n196 VSUBS 0.035561f
C1227 VTAIL.n197 VSUBS 0.240739f
C1228 VTAIL.t13 VSUBS 0.326723f
C1229 VTAIL.t8 VSUBS 0.326723f
C1230 VTAIL.n198 VSUBS 2.55802f
C1231 VTAIL.n199 VSUBS 0.948484f
C1232 VTAIL.n200 VSUBS 0.025431f
C1233 VTAIL.n201 VSUBS 0.023599f
C1234 VTAIL.n202 VSUBS 0.012681f
C1235 VTAIL.n203 VSUBS 0.029973f
C1236 VTAIL.n204 VSUBS 0.013427f
C1237 VTAIL.n205 VSUBS 0.023599f
C1238 VTAIL.n206 VSUBS 0.012681f
C1239 VTAIL.n207 VSUBS 0.029973f
C1240 VTAIL.n208 VSUBS 0.013054f
C1241 VTAIL.n209 VSUBS 0.023599f
C1242 VTAIL.n210 VSUBS 0.013427f
C1243 VTAIL.n211 VSUBS 0.029973f
C1244 VTAIL.n212 VSUBS 0.013427f
C1245 VTAIL.n213 VSUBS 0.023599f
C1246 VTAIL.n214 VSUBS 0.012681f
C1247 VTAIL.n215 VSUBS 0.029973f
C1248 VTAIL.n216 VSUBS 0.013427f
C1249 VTAIL.n217 VSUBS 0.023599f
C1250 VTAIL.n218 VSUBS 0.012681f
C1251 VTAIL.n219 VSUBS 0.029973f
C1252 VTAIL.n220 VSUBS 0.013427f
C1253 VTAIL.n221 VSUBS 0.023599f
C1254 VTAIL.n222 VSUBS 0.012681f
C1255 VTAIL.n223 VSUBS 0.029973f
C1256 VTAIL.n224 VSUBS 0.013427f
C1257 VTAIL.n225 VSUBS 0.023599f
C1258 VTAIL.n226 VSUBS 0.012681f
C1259 VTAIL.n227 VSUBS 0.029973f
C1260 VTAIL.n228 VSUBS 0.013427f
C1261 VTAIL.n229 VSUBS 1.77681f
C1262 VTAIL.n230 VSUBS 0.012681f
C1263 VTAIL.t11 VSUBS 0.064315f
C1264 VTAIL.n231 VSUBS 0.183893f
C1265 VTAIL.n232 VSUBS 0.019068f
C1266 VTAIL.n233 VSUBS 0.02248f
C1267 VTAIL.n234 VSUBS 0.029973f
C1268 VTAIL.n235 VSUBS 0.013427f
C1269 VTAIL.n236 VSUBS 0.012681f
C1270 VTAIL.n237 VSUBS 0.023599f
C1271 VTAIL.n238 VSUBS 0.023599f
C1272 VTAIL.n239 VSUBS 0.012681f
C1273 VTAIL.n240 VSUBS 0.013427f
C1274 VTAIL.n241 VSUBS 0.029973f
C1275 VTAIL.n242 VSUBS 0.029973f
C1276 VTAIL.n243 VSUBS 0.013427f
C1277 VTAIL.n244 VSUBS 0.012681f
C1278 VTAIL.n245 VSUBS 0.023599f
C1279 VTAIL.n246 VSUBS 0.023599f
C1280 VTAIL.n247 VSUBS 0.012681f
C1281 VTAIL.n248 VSUBS 0.013427f
C1282 VTAIL.n249 VSUBS 0.029973f
C1283 VTAIL.n250 VSUBS 0.029973f
C1284 VTAIL.n251 VSUBS 0.013427f
C1285 VTAIL.n252 VSUBS 0.012681f
C1286 VTAIL.n253 VSUBS 0.023599f
C1287 VTAIL.n254 VSUBS 0.023599f
C1288 VTAIL.n255 VSUBS 0.012681f
C1289 VTAIL.n256 VSUBS 0.013427f
C1290 VTAIL.n257 VSUBS 0.029973f
C1291 VTAIL.n258 VSUBS 0.029973f
C1292 VTAIL.n259 VSUBS 0.013427f
C1293 VTAIL.n260 VSUBS 0.012681f
C1294 VTAIL.n261 VSUBS 0.023599f
C1295 VTAIL.n262 VSUBS 0.023599f
C1296 VTAIL.n263 VSUBS 0.012681f
C1297 VTAIL.n264 VSUBS 0.013427f
C1298 VTAIL.n265 VSUBS 0.029973f
C1299 VTAIL.n266 VSUBS 0.029973f
C1300 VTAIL.n267 VSUBS 0.013427f
C1301 VTAIL.n268 VSUBS 0.012681f
C1302 VTAIL.n269 VSUBS 0.023599f
C1303 VTAIL.n270 VSUBS 0.023599f
C1304 VTAIL.n271 VSUBS 0.012681f
C1305 VTAIL.n272 VSUBS 0.012681f
C1306 VTAIL.n273 VSUBS 0.013427f
C1307 VTAIL.n274 VSUBS 0.029973f
C1308 VTAIL.n275 VSUBS 0.029973f
C1309 VTAIL.n276 VSUBS 0.029973f
C1310 VTAIL.n277 VSUBS 0.013054f
C1311 VTAIL.n278 VSUBS 0.012681f
C1312 VTAIL.n279 VSUBS 0.023599f
C1313 VTAIL.n280 VSUBS 0.023599f
C1314 VTAIL.n281 VSUBS 0.012681f
C1315 VTAIL.n282 VSUBS 0.013427f
C1316 VTAIL.n283 VSUBS 0.029973f
C1317 VTAIL.n284 VSUBS 0.029973f
C1318 VTAIL.n285 VSUBS 0.013427f
C1319 VTAIL.n286 VSUBS 0.012681f
C1320 VTAIL.n287 VSUBS 0.023599f
C1321 VTAIL.n288 VSUBS 0.023599f
C1322 VTAIL.n289 VSUBS 0.012681f
C1323 VTAIL.n290 VSUBS 0.013427f
C1324 VTAIL.n291 VSUBS 0.029973f
C1325 VTAIL.n292 VSUBS 0.070863f
C1326 VTAIL.n293 VSUBS 0.013427f
C1327 VTAIL.n294 VSUBS 0.012681f
C1328 VTAIL.n295 VSUBS 0.054548f
C1329 VTAIL.n296 VSUBS 0.035561f
C1330 VTAIL.n297 VSUBS 1.85891f
C1331 VTAIL.n298 VSUBS 0.025431f
C1332 VTAIL.n299 VSUBS 0.023599f
C1333 VTAIL.n300 VSUBS 0.012681f
C1334 VTAIL.n301 VSUBS 0.029973f
C1335 VTAIL.n302 VSUBS 0.013427f
C1336 VTAIL.n303 VSUBS 0.023599f
C1337 VTAIL.n304 VSUBS 0.012681f
C1338 VTAIL.n305 VSUBS 0.029973f
C1339 VTAIL.n306 VSUBS 0.013054f
C1340 VTAIL.n307 VSUBS 0.023599f
C1341 VTAIL.n308 VSUBS 0.013054f
C1342 VTAIL.n309 VSUBS 0.012681f
C1343 VTAIL.n310 VSUBS 0.029973f
C1344 VTAIL.n311 VSUBS 0.029973f
C1345 VTAIL.n312 VSUBS 0.013427f
C1346 VTAIL.n313 VSUBS 0.023599f
C1347 VTAIL.n314 VSUBS 0.012681f
C1348 VTAIL.n315 VSUBS 0.029973f
C1349 VTAIL.n316 VSUBS 0.013427f
C1350 VTAIL.n317 VSUBS 0.023599f
C1351 VTAIL.n318 VSUBS 0.012681f
C1352 VTAIL.n319 VSUBS 0.029973f
C1353 VTAIL.n320 VSUBS 0.013427f
C1354 VTAIL.n321 VSUBS 0.023599f
C1355 VTAIL.n322 VSUBS 0.012681f
C1356 VTAIL.n323 VSUBS 0.029973f
C1357 VTAIL.n324 VSUBS 0.013427f
C1358 VTAIL.n325 VSUBS 0.023599f
C1359 VTAIL.n326 VSUBS 0.012681f
C1360 VTAIL.n327 VSUBS 0.029973f
C1361 VTAIL.n328 VSUBS 0.013427f
C1362 VTAIL.n329 VSUBS 1.77681f
C1363 VTAIL.n330 VSUBS 0.012681f
C1364 VTAIL.t4 VSUBS 0.064315f
C1365 VTAIL.n331 VSUBS 0.183893f
C1366 VTAIL.n332 VSUBS 0.019068f
C1367 VTAIL.n333 VSUBS 0.02248f
C1368 VTAIL.n334 VSUBS 0.029973f
C1369 VTAIL.n335 VSUBS 0.013427f
C1370 VTAIL.n336 VSUBS 0.012681f
C1371 VTAIL.n337 VSUBS 0.023599f
C1372 VTAIL.n338 VSUBS 0.023599f
C1373 VTAIL.n339 VSUBS 0.012681f
C1374 VTAIL.n340 VSUBS 0.013427f
C1375 VTAIL.n341 VSUBS 0.029973f
C1376 VTAIL.n342 VSUBS 0.029973f
C1377 VTAIL.n343 VSUBS 0.013427f
C1378 VTAIL.n344 VSUBS 0.012681f
C1379 VTAIL.n345 VSUBS 0.023599f
C1380 VTAIL.n346 VSUBS 0.023599f
C1381 VTAIL.n347 VSUBS 0.012681f
C1382 VTAIL.n348 VSUBS 0.013427f
C1383 VTAIL.n349 VSUBS 0.029973f
C1384 VTAIL.n350 VSUBS 0.029973f
C1385 VTAIL.n351 VSUBS 0.013427f
C1386 VTAIL.n352 VSUBS 0.012681f
C1387 VTAIL.n353 VSUBS 0.023599f
C1388 VTAIL.n354 VSUBS 0.023599f
C1389 VTAIL.n355 VSUBS 0.012681f
C1390 VTAIL.n356 VSUBS 0.013427f
C1391 VTAIL.n357 VSUBS 0.029973f
C1392 VTAIL.n358 VSUBS 0.029973f
C1393 VTAIL.n359 VSUBS 0.013427f
C1394 VTAIL.n360 VSUBS 0.012681f
C1395 VTAIL.n361 VSUBS 0.023599f
C1396 VTAIL.n362 VSUBS 0.023599f
C1397 VTAIL.n363 VSUBS 0.012681f
C1398 VTAIL.n364 VSUBS 0.013427f
C1399 VTAIL.n365 VSUBS 0.029973f
C1400 VTAIL.n366 VSUBS 0.029973f
C1401 VTAIL.n367 VSUBS 0.013427f
C1402 VTAIL.n368 VSUBS 0.012681f
C1403 VTAIL.n369 VSUBS 0.023599f
C1404 VTAIL.n370 VSUBS 0.023599f
C1405 VTAIL.n371 VSUBS 0.012681f
C1406 VTAIL.n372 VSUBS 0.013427f
C1407 VTAIL.n373 VSUBS 0.029973f
C1408 VTAIL.n374 VSUBS 0.029973f
C1409 VTAIL.n375 VSUBS 0.013427f
C1410 VTAIL.n376 VSUBS 0.012681f
C1411 VTAIL.n377 VSUBS 0.023599f
C1412 VTAIL.n378 VSUBS 0.023599f
C1413 VTAIL.n379 VSUBS 0.012681f
C1414 VTAIL.n380 VSUBS 0.013427f
C1415 VTAIL.n381 VSUBS 0.029973f
C1416 VTAIL.n382 VSUBS 0.029973f
C1417 VTAIL.n383 VSUBS 0.013427f
C1418 VTAIL.n384 VSUBS 0.012681f
C1419 VTAIL.n385 VSUBS 0.023599f
C1420 VTAIL.n386 VSUBS 0.023599f
C1421 VTAIL.n387 VSUBS 0.012681f
C1422 VTAIL.n388 VSUBS 0.013427f
C1423 VTAIL.n389 VSUBS 0.029973f
C1424 VTAIL.n390 VSUBS 0.070863f
C1425 VTAIL.n391 VSUBS 0.013427f
C1426 VTAIL.n392 VSUBS 0.012681f
C1427 VTAIL.n393 VSUBS 0.054548f
C1428 VTAIL.n394 VSUBS 0.035561f
C1429 VTAIL.n395 VSUBS 1.85891f
C1430 VTAIL.t2 VSUBS 0.326723f
C1431 VTAIL.t5 VSUBS 0.326723f
C1432 VTAIL.n396 VSUBS 2.55804f
C1433 VTAIL.n397 VSUBS 0.948468f
C1434 VTAIL.n398 VSUBS 0.025431f
C1435 VTAIL.n399 VSUBS 0.023599f
C1436 VTAIL.n400 VSUBS 0.012681f
C1437 VTAIL.n401 VSUBS 0.029973f
C1438 VTAIL.n402 VSUBS 0.013427f
C1439 VTAIL.n403 VSUBS 0.023599f
C1440 VTAIL.n404 VSUBS 0.012681f
C1441 VTAIL.n405 VSUBS 0.029973f
C1442 VTAIL.n406 VSUBS 0.013054f
C1443 VTAIL.n407 VSUBS 0.023599f
C1444 VTAIL.n408 VSUBS 0.013054f
C1445 VTAIL.n409 VSUBS 0.012681f
C1446 VTAIL.n410 VSUBS 0.029973f
C1447 VTAIL.n411 VSUBS 0.029973f
C1448 VTAIL.n412 VSUBS 0.013427f
C1449 VTAIL.n413 VSUBS 0.023599f
C1450 VTAIL.n414 VSUBS 0.012681f
C1451 VTAIL.n415 VSUBS 0.029973f
C1452 VTAIL.n416 VSUBS 0.013427f
C1453 VTAIL.n417 VSUBS 0.023599f
C1454 VTAIL.n418 VSUBS 0.012681f
C1455 VTAIL.n419 VSUBS 0.029973f
C1456 VTAIL.n420 VSUBS 0.013427f
C1457 VTAIL.n421 VSUBS 0.023599f
C1458 VTAIL.n422 VSUBS 0.012681f
C1459 VTAIL.n423 VSUBS 0.029973f
C1460 VTAIL.n424 VSUBS 0.013427f
C1461 VTAIL.n425 VSUBS 0.023599f
C1462 VTAIL.n426 VSUBS 0.012681f
C1463 VTAIL.n427 VSUBS 0.029973f
C1464 VTAIL.n428 VSUBS 0.013427f
C1465 VTAIL.n429 VSUBS 1.77681f
C1466 VTAIL.n430 VSUBS 0.012681f
C1467 VTAIL.t3 VSUBS 0.064315f
C1468 VTAIL.n431 VSUBS 0.183893f
C1469 VTAIL.n432 VSUBS 0.019068f
C1470 VTAIL.n433 VSUBS 0.02248f
C1471 VTAIL.n434 VSUBS 0.029973f
C1472 VTAIL.n435 VSUBS 0.013427f
C1473 VTAIL.n436 VSUBS 0.012681f
C1474 VTAIL.n437 VSUBS 0.023599f
C1475 VTAIL.n438 VSUBS 0.023599f
C1476 VTAIL.n439 VSUBS 0.012681f
C1477 VTAIL.n440 VSUBS 0.013427f
C1478 VTAIL.n441 VSUBS 0.029973f
C1479 VTAIL.n442 VSUBS 0.029973f
C1480 VTAIL.n443 VSUBS 0.013427f
C1481 VTAIL.n444 VSUBS 0.012681f
C1482 VTAIL.n445 VSUBS 0.023599f
C1483 VTAIL.n446 VSUBS 0.023599f
C1484 VTAIL.n447 VSUBS 0.012681f
C1485 VTAIL.n448 VSUBS 0.013427f
C1486 VTAIL.n449 VSUBS 0.029973f
C1487 VTAIL.n450 VSUBS 0.029973f
C1488 VTAIL.n451 VSUBS 0.013427f
C1489 VTAIL.n452 VSUBS 0.012681f
C1490 VTAIL.n453 VSUBS 0.023599f
C1491 VTAIL.n454 VSUBS 0.023599f
C1492 VTAIL.n455 VSUBS 0.012681f
C1493 VTAIL.n456 VSUBS 0.013427f
C1494 VTAIL.n457 VSUBS 0.029973f
C1495 VTAIL.n458 VSUBS 0.029973f
C1496 VTAIL.n459 VSUBS 0.013427f
C1497 VTAIL.n460 VSUBS 0.012681f
C1498 VTAIL.n461 VSUBS 0.023599f
C1499 VTAIL.n462 VSUBS 0.023599f
C1500 VTAIL.n463 VSUBS 0.012681f
C1501 VTAIL.n464 VSUBS 0.013427f
C1502 VTAIL.n465 VSUBS 0.029973f
C1503 VTAIL.n466 VSUBS 0.029973f
C1504 VTAIL.n467 VSUBS 0.013427f
C1505 VTAIL.n468 VSUBS 0.012681f
C1506 VTAIL.n469 VSUBS 0.023599f
C1507 VTAIL.n470 VSUBS 0.023599f
C1508 VTAIL.n471 VSUBS 0.012681f
C1509 VTAIL.n472 VSUBS 0.013427f
C1510 VTAIL.n473 VSUBS 0.029973f
C1511 VTAIL.n474 VSUBS 0.029973f
C1512 VTAIL.n475 VSUBS 0.013427f
C1513 VTAIL.n476 VSUBS 0.012681f
C1514 VTAIL.n477 VSUBS 0.023599f
C1515 VTAIL.n478 VSUBS 0.023599f
C1516 VTAIL.n479 VSUBS 0.012681f
C1517 VTAIL.n480 VSUBS 0.013427f
C1518 VTAIL.n481 VSUBS 0.029973f
C1519 VTAIL.n482 VSUBS 0.029973f
C1520 VTAIL.n483 VSUBS 0.013427f
C1521 VTAIL.n484 VSUBS 0.012681f
C1522 VTAIL.n485 VSUBS 0.023599f
C1523 VTAIL.n486 VSUBS 0.023599f
C1524 VTAIL.n487 VSUBS 0.012681f
C1525 VTAIL.n488 VSUBS 0.013427f
C1526 VTAIL.n489 VSUBS 0.029973f
C1527 VTAIL.n490 VSUBS 0.070863f
C1528 VTAIL.n491 VSUBS 0.013427f
C1529 VTAIL.n492 VSUBS 0.012681f
C1530 VTAIL.n493 VSUBS 0.054548f
C1531 VTAIL.n494 VSUBS 0.035561f
C1532 VTAIL.n495 VSUBS 0.240739f
C1533 VTAIL.n496 VSUBS 0.025431f
C1534 VTAIL.n497 VSUBS 0.023599f
C1535 VTAIL.n498 VSUBS 0.012681f
C1536 VTAIL.n499 VSUBS 0.029973f
C1537 VTAIL.n500 VSUBS 0.013427f
C1538 VTAIL.n501 VSUBS 0.023599f
C1539 VTAIL.n502 VSUBS 0.012681f
C1540 VTAIL.n503 VSUBS 0.029973f
C1541 VTAIL.n504 VSUBS 0.013054f
C1542 VTAIL.n505 VSUBS 0.023599f
C1543 VTAIL.n506 VSUBS 0.013054f
C1544 VTAIL.n507 VSUBS 0.012681f
C1545 VTAIL.n508 VSUBS 0.029973f
C1546 VTAIL.n509 VSUBS 0.029973f
C1547 VTAIL.n510 VSUBS 0.013427f
C1548 VTAIL.n511 VSUBS 0.023599f
C1549 VTAIL.n512 VSUBS 0.012681f
C1550 VTAIL.n513 VSUBS 0.029973f
C1551 VTAIL.n514 VSUBS 0.013427f
C1552 VTAIL.n515 VSUBS 0.023599f
C1553 VTAIL.n516 VSUBS 0.012681f
C1554 VTAIL.n517 VSUBS 0.029973f
C1555 VTAIL.n518 VSUBS 0.013427f
C1556 VTAIL.n519 VSUBS 0.023599f
C1557 VTAIL.n520 VSUBS 0.012681f
C1558 VTAIL.n521 VSUBS 0.029973f
C1559 VTAIL.n522 VSUBS 0.013427f
C1560 VTAIL.n523 VSUBS 0.023599f
C1561 VTAIL.n524 VSUBS 0.012681f
C1562 VTAIL.n525 VSUBS 0.029973f
C1563 VTAIL.n526 VSUBS 0.013427f
C1564 VTAIL.n527 VSUBS 1.77681f
C1565 VTAIL.n528 VSUBS 0.012681f
C1566 VTAIL.t12 VSUBS 0.064315f
C1567 VTAIL.n529 VSUBS 0.183893f
C1568 VTAIL.n530 VSUBS 0.019068f
C1569 VTAIL.n531 VSUBS 0.02248f
C1570 VTAIL.n532 VSUBS 0.029973f
C1571 VTAIL.n533 VSUBS 0.013427f
C1572 VTAIL.n534 VSUBS 0.012681f
C1573 VTAIL.n535 VSUBS 0.023599f
C1574 VTAIL.n536 VSUBS 0.023599f
C1575 VTAIL.n537 VSUBS 0.012681f
C1576 VTAIL.n538 VSUBS 0.013427f
C1577 VTAIL.n539 VSUBS 0.029973f
C1578 VTAIL.n540 VSUBS 0.029973f
C1579 VTAIL.n541 VSUBS 0.013427f
C1580 VTAIL.n542 VSUBS 0.012681f
C1581 VTAIL.n543 VSUBS 0.023599f
C1582 VTAIL.n544 VSUBS 0.023599f
C1583 VTAIL.n545 VSUBS 0.012681f
C1584 VTAIL.n546 VSUBS 0.013427f
C1585 VTAIL.n547 VSUBS 0.029973f
C1586 VTAIL.n548 VSUBS 0.029973f
C1587 VTAIL.n549 VSUBS 0.013427f
C1588 VTAIL.n550 VSUBS 0.012681f
C1589 VTAIL.n551 VSUBS 0.023599f
C1590 VTAIL.n552 VSUBS 0.023599f
C1591 VTAIL.n553 VSUBS 0.012681f
C1592 VTAIL.n554 VSUBS 0.013427f
C1593 VTAIL.n555 VSUBS 0.029973f
C1594 VTAIL.n556 VSUBS 0.029973f
C1595 VTAIL.n557 VSUBS 0.013427f
C1596 VTAIL.n558 VSUBS 0.012681f
C1597 VTAIL.n559 VSUBS 0.023599f
C1598 VTAIL.n560 VSUBS 0.023599f
C1599 VTAIL.n561 VSUBS 0.012681f
C1600 VTAIL.n562 VSUBS 0.013427f
C1601 VTAIL.n563 VSUBS 0.029973f
C1602 VTAIL.n564 VSUBS 0.029973f
C1603 VTAIL.n565 VSUBS 0.013427f
C1604 VTAIL.n566 VSUBS 0.012681f
C1605 VTAIL.n567 VSUBS 0.023599f
C1606 VTAIL.n568 VSUBS 0.023599f
C1607 VTAIL.n569 VSUBS 0.012681f
C1608 VTAIL.n570 VSUBS 0.013427f
C1609 VTAIL.n571 VSUBS 0.029973f
C1610 VTAIL.n572 VSUBS 0.029973f
C1611 VTAIL.n573 VSUBS 0.013427f
C1612 VTAIL.n574 VSUBS 0.012681f
C1613 VTAIL.n575 VSUBS 0.023599f
C1614 VTAIL.n576 VSUBS 0.023599f
C1615 VTAIL.n577 VSUBS 0.012681f
C1616 VTAIL.n578 VSUBS 0.013427f
C1617 VTAIL.n579 VSUBS 0.029973f
C1618 VTAIL.n580 VSUBS 0.029973f
C1619 VTAIL.n581 VSUBS 0.013427f
C1620 VTAIL.n582 VSUBS 0.012681f
C1621 VTAIL.n583 VSUBS 0.023599f
C1622 VTAIL.n584 VSUBS 0.023599f
C1623 VTAIL.n585 VSUBS 0.012681f
C1624 VTAIL.n586 VSUBS 0.013427f
C1625 VTAIL.n587 VSUBS 0.029973f
C1626 VTAIL.n588 VSUBS 0.070863f
C1627 VTAIL.n589 VSUBS 0.013427f
C1628 VTAIL.n590 VSUBS 0.012681f
C1629 VTAIL.n591 VSUBS 0.054548f
C1630 VTAIL.n592 VSUBS 0.035561f
C1631 VTAIL.n593 VSUBS 0.240739f
C1632 VTAIL.t14 VSUBS 0.326723f
C1633 VTAIL.t15 VSUBS 0.326723f
C1634 VTAIL.n594 VSUBS 2.55804f
C1635 VTAIL.n595 VSUBS 0.948468f
C1636 VTAIL.n596 VSUBS 0.025431f
C1637 VTAIL.n597 VSUBS 0.023599f
C1638 VTAIL.n598 VSUBS 0.012681f
C1639 VTAIL.n599 VSUBS 0.029973f
C1640 VTAIL.n600 VSUBS 0.013427f
C1641 VTAIL.n601 VSUBS 0.023599f
C1642 VTAIL.n602 VSUBS 0.012681f
C1643 VTAIL.n603 VSUBS 0.029973f
C1644 VTAIL.n604 VSUBS 0.013054f
C1645 VTAIL.n605 VSUBS 0.023599f
C1646 VTAIL.n606 VSUBS 0.013054f
C1647 VTAIL.n607 VSUBS 0.012681f
C1648 VTAIL.n608 VSUBS 0.029973f
C1649 VTAIL.n609 VSUBS 0.029973f
C1650 VTAIL.n610 VSUBS 0.013427f
C1651 VTAIL.n611 VSUBS 0.023599f
C1652 VTAIL.n612 VSUBS 0.012681f
C1653 VTAIL.n613 VSUBS 0.029973f
C1654 VTAIL.n614 VSUBS 0.013427f
C1655 VTAIL.n615 VSUBS 0.023599f
C1656 VTAIL.n616 VSUBS 0.012681f
C1657 VTAIL.n617 VSUBS 0.029973f
C1658 VTAIL.n618 VSUBS 0.013427f
C1659 VTAIL.n619 VSUBS 0.023599f
C1660 VTAIL.n620 VSUBS 0.012681f
C1661 VTAIL.n621 VSUBS 0.029973f
C1662 VTAIL.n622 VSUBS 0.013427f
C1663 VTAIL.n623 VSUBS 0.023599f
C1664 VTAIL.n624 VSUBS 0.012681f
C1665 VTAIL.n625 VSUBS 0.029973f
C1666 VTAIL.n626 VSUBS 0.013427f
C1667 VTAIL.n627 VSUBS 1.77681f
C1668 VTAIL.n628 VSUBS 0.012681f
C1669 VTAIL.t10 VSUBS 0.064315f
C1670 VTAIL.n629 VSUBS 0.183893f
C1671 VTAIL.n630 VSUBS 0.019068f
C1672 VTAIL.n631 VSUBS 0.02248f
C1673 VTAIL.n632 VSUBS 0.029973f
C1674 VTAIL.n633 VSUBS 0.013427f
C1675 VTAIL.n634 VSUBS 0.012681f
C1676 VTAIL.n635 VSUBS 0.023599f
C1677 VTAIL.n636 VSUBS 0.023599f
C1678 VTAIL.n637 VSUBS 0.012681f
C1679 VTAIL.n638 VSUBS 0.013427f
C1680 VTAIL.n639 VSUBS 0.029973f
C1681 VTAIL.n640 VSUBS 0.029973f
C1682 VTAIL.n641 VSUBS 0.013427f
C1683 VTAIL.n642 VSUBS 0.012681f
C1684 VTAIL.n643 VSUBS 0.023599f
C1685 VTAIL.n644 VSUBS 0.023599f
C1686 VTAIL.n645 VSUBS 0.012681f
C1687 VTAIL.n646 VSUBS 0.013427f
C1688 VTAIL.n647 VSUBS 0.029973f
C1689 VTAIL.n648 VSUBS 0.029973f
C1690 VTAIL.n649 VSUBS 0.013427f
C1691 VTAIL.n650 VSUBS 0.012681f
C1692 VTAIL.n651 VSUBS 0.023599f
C1693 VTAIL.n652 VSUBS 0.023599f
C1694 VTAIL.n653 VSUBS 0.012681f
C1695 VTAIL.n654 VSUBS 0.013427f
C1696 VTAIL.n655 VSUBS 0.029973f
C1697 VTAIL.n656 VSUBS 0.029973f
C1698 VTAIL.n657 VSUBS 0.013427f
C1699 VTAIL.n658 VSUBS 0.012681f
C1700 VTAIL.n659 VSUBS 0.023599f
C1701 VTAIL.n660 VSUBS 0.023599f
C1702 VTAIL.n661 VSUBS 0.012681f
C1703 VTAIL.n662 VSUBS 0.013427f
C1704 VTAIL.n663 VSUBS 0.029973f
C1705 VTAIL.n664 VSUBS 0.029973f
C1706 VTAIL.n665 VSUBS 0.013427f
C1707 VTAIL.n666 VSUBS 0.012681f
C1708 VTAIL.n667 VSUBS 0.023599f
C1709 VTAIL.n668 VSUBS 0.023599f
C1710 VTAIL.n669 VSUBS 0.012681f
C1711 VTAIL.n670 VSUBS 0.013427f
C1712 VTAIL.n671 VSUBS 0.029973f
C1713 VTAIL.n672 VSUBS 0.029973f
C1714 VTAIL.n673 VSUBS 0.013427f
C1715 VTAIL.n674 VSUBS 0.012681f
C1716 VTAIL.n675 VSUBS 0.023599f
C1717 VTAIL.n676 VSUBS 0.023599f
C1718 VTAIL.n677 VSUBS 0.012681f
C1719 VTAIL.n678 VSUBS 0.013427f
C1720 VTAIL.n679 VSUBS 0.029973f
C1721 VTAIL.n680 VSUBS 0.029973f
C1722 VTAIL.n681 VSUBS 0.013427f
C1723 VTAIL.n682 VSUBS 0.012681f
C1724 VTAIL.n683 VSUBS 0.023599f
C1725 VTAIL.n684 VSUBS 0.023599f
C1726 VTAIL.n685 VSUBS 0.012681f
C1727 VTAIL.n686 VSUBS 0.013427f
C1728 VTAIL.n687 VSUBS 0.029973f
C1729 VTAIL.n688 VSUBS 0.070863f
C1730 VTAIL.n689 VSUBS 0.013427f
C1731 VTAIL.n690 VSUBS 0.012681f
C1732 VTAIL.n691 VSUBS 0.054548f
C1733 VTAIL.n692 VSUBS 0.035561f
C1734 VTAIL.n693 VSUBS 1.85891f
C1735 VTAIL.n694 VSUBS 0.025431f
C1736 VTAIL.n695 VSUBS 0.023599f
C1737 VTAIL.n696 VSUBS 0.012681f
C1738 VTAIL.n697 VSUBS 0.029973f
C1739 VTAIL.n698 VSUBS 0.013427f
C1740 VTAIL.n699 VSUBS 0.023599f
C1741 VTAIL.n700 VSUBS 0.012681f
C1742 VTAIL.n701 VSUBS 0.029973f
C1743 VTAIL.n702 VSUBS 0.013054f
C1744 VTAIL.n703 VSUBS 0.023599f
C1745 VTAIL.n704 VSUBS 0.013427f
C1746 VTAIL.n705 VSUBS 0.029973f
C1747 VTAIL.n706 VSUBS 0.013427f
C1748 VTAIL.n707 VSUBS 0.023599f
C1749 VTAIL.n708 VSUBS 0.012681f
C1750 VTAIL.n709 VSUBS 0.029973f
C1751 VTAIL.n710 VSUBS 0.013427f
C1752 VTAIL.n711 VSUBS 0.023599f
C1753 VTAIL.n712 VSUBS 0.012681f
C1754 VTAIL.n713 VSUBS 0.029973f
C1755 VTAIL.n714 VSUBS 0.013427f
C1756 VTAIL.n715 VSUBS 0.023599f
C1757 VTAIL.n716 VSUBS 0.012681f
C1758 VTAIL.n717 VSUBS 0.029973f
C1759 VTAIL.n718 VSUBS 0.013427f
C1760 VTAIL.n719 VSUBS 0.023599f
C1761 VTAIL.n720 VSUBS 0.012681f
C1762 VTAIL.n721 VSUBS 0.029973f
C1763 VTAIL.n722 VSUBS 0.013427f
C1764 VTAIL.n723 VSUBS 1.77681f
C1765 VTAIL.n724 VSUBS 0.012681f
C1766 VTAIL.t1 VSUBS 0.064315f
C1767 VTAIL.n725 VSUBS 0.183893f
C1768 VTAIL.n726 VSUBS 0.019068f
C1769 VTAIL.n727 VSUBS 0.02248f
C1770 VTAIL.n728 VSUBS 0.029973f
C1771 VTAIL.n729 VSUBS 0.013427f
C1772 VTAIL.n730 VSUBS 0.012681f
C1773 VTAIL.n731 VSUBS 0.023599f
C1774 VTAIL.n732 VSUBS 0.023599f
C1775 VTAIL.n733 VSUBS 0.012681f
C1776 VTAIL.n734 VSUBS 0.013427f
C1777 VTAIL.n735 VSUBS 0.029973f
C1778 VTAIL.n736 VSUBS 0.029973f
C1779 VTAIL.n737 VSUBS 0.013427f
C1780 VTAIL.n738 VSUBS 0.012681f
C1781 VTAIL.n739 VSUBS 0.023599f
C1782 VTAIL.n740 VSUBS 0.023599f
C1783 VTAIL.n741 VSUBS 0.012681f
C1784 VTAIL.n742 VSUBS 0.013427f
C1785 VTAIL.n743 VSUBS 0.029973f
C1786 VTAIL.n744 VSUBS 0.029973f
C1787 VTAIL.n745 VSUBS 0.013427f
C1788 VTAIL.n746 VSUBS 0.012681f
C1789 VTAIL.n747 VSUBS 0.023599f
C1790 VTAIL.n748 VSUBS 0.023599f
C1791 VTAIL.n749 VSUBS 0.012681f
C1792 VTAIL.n750 VSUBS 0.013427f
C1793 VTAIL.n751 VSUBS 0.029973f
C1794 VTAIL.n752 VSUBS 0.029973f
C1795 VTAIL.n753 VSUBS 0.013427f
C1796 VTAIL.n754 VSUBS 0.012681f
C1797 VTAIL.n755 VSUBS 0.023599f
C1798 VTAIL.n756 VSUBS 0.023599f
C1799 VTAIL.n757 VSUBS 0.012681f
C1800 VTAIL.n758 VSUBS 0.013427f
C1801 VTAIL.n759 VSUBS 0.029973f
C1802 VTAIL.n760 VSUBS 0.029973f
C1803 VTAIL.n761 VSUBS 0.013427f
C1804 VTAIL.n762 VSUBS 0.012681f
C1805 VTAIL.n763 VSUBS 0.023599f
C1806 VTAIL.n764 VSUBS 0.023599f
C1807 VTAIL.n765 VSUBS 0.012681f
C1808 VTAIL.n766 VSUBS 0.012681f
C1809 VTAIL.n767 VSUBS 0.013427f
C1810 VTAIL.n768 VSUBS 0.029973f
C1811 VTAIL.n769 VSUBS 0.029973f
C1812 VTAIL.n770 VSUBS 0.029973f
C1813 VTAIL.n771 VSUBS 0.013054f
C1814 VTAIL.n772 VSUBS 0.012681f
C1815 VTAIL.n773 VSUBS 0.023599f
C1816 VTAIL.n774 VSUBS 0.023599f
C1817 VTAIL.n775 VSUBS 0.012681f
C1818 VTAIL.n776 VSUBS 0.013427f
C1819 VTAIL.n777 VSUBS 0.029973f
C1820 VTAIL.n778 VSUBS 0.029973f
C1821 VTAIL.n779 VSUBS 0.013427f
C1822 VTAIL.n780 VSUBS 0.012681f
C1823 VTAIL.n781 VSUBS 0.023599f
C1824 VTAIL.n782 VSUBS 0.023599f
C1825 VTAIL.n783 VSUBS 0.012681f
C1826 VTAIL.n784 VSUBS 0.013427f
C1827 VTAIL.n785 VSUBS 0.029973f
C1828 VTAIL.n786 VSUBS 0.070863f
C1829 VTAIL.n787 VSUBS 0.013427f
C1830 VTAIL.n788 VSUBS 0.012681f
C1831 VTAIL.n789 VSUBS 0.054548f
C1832 VTAIL.n790 VSUBS 0.035561f
C1833 VTAIL.n791 VSUBS 1.85449f
C1834 VDD1.t0 VSUBS 0.371948f
C1835 VDD1.t2 VSUBS 0.371948f
C1836 VDD1.n0 VSUBS 3.0945f
C1837 VDD1.t7 VSUBS 0.371948f
C1838 VDD1.t1 VSUBS 0.371948f
C1839 VDD1.n1 VSUBS 3.09297f
C1840 VDD1.t4 VSUBS 0.371948f
C1841 VDD1.t5 VSUBS 0.371948f
C1842 VDD1.n2 VSUBS 3.09297f
C1843 VDD1.n3 VSUBS 4.49072f
C1844 VDD1.t3 VSUBS 0.371948f
C1845 VDD1.t6 VSUBS 0.371948f
C1846 VDD1.n4 VSUBS 3.07891f
C1847 VDD1.n5 VSUBS 3.91938f
C1848 VP.n0 VSUBS 0.038096f
C1849 VP.t6 VSUBS 3.46572f
C1850 VP.n1 VSUBS 0.03641f
C1851 VP.n2 VSUBS 0.028898f
C1852 VP.t7 VSUBS 3.46572f
C1853 VP.n3 VSUBS 1.2041f
C1854 VP.n4 VSUBS 0.028898f
C1855 VP.n5 VSUBS 0.057131f
C1856 VP.n6 VSUBS 0.028898f
C1857 VP.t2 VSUBS 3.46572f
C1858 VP.n7 VSUBS 0.047604f
C1859 VP.n8 VSUBS 0.028898f
C1860 VP.t4 VSUBS 3.46572f
C1861 VP.n9 VSUBS 1.2982f
C1862 VP.n10 VSUBS 0.038096f
C1863 VP.t5 VSUBS 3.46572f
C1864 VP.n11 VSUBS 0.03641f
C1865 VP.n12 VSUBS 0.028898f
C1866 VP.t0 VSUBS 3.46572f
C1867 VP.n13 VSUBS 1.2041f
C1868 VP.n14 VSUBS 0.028898f
C1869 VP.n15 VSUBS 0.057131f
C1870 VP.t3 VSUBS 3.69603f
C1871 VP.n16 VSUBS 1.25676f
C1872 VP.t1 VSUBS 3.46572f
C1873 VP.n17 VSUBS 1.29432f
C1874 VP.n18 VSUBS 0.048826f
C1875 VP.n19 VSUBS 0.27611f
C1876 VP.n20 VSUBS 0.028898f
C1877 VP.n21 VSUBS 0.028898f
C1878 VP.n22 VSUBS 0.02334f
C1879 VP.n23 VSUBS 0.057131f
C1880 VP.n24 VSUBS 0.048826f
C1881 VP.n25 VSUBS 0.028898f
C1882 VP.n26 VSUBS 0.028898f
C1883 VP.n27 VSUBS 0.031895f
C1884 VP.n28 VSUBS 0.053588f
C1885 VP.n29 VSUBS 0.047604f
C1886 VP.n30 VSUBS 0.028898f
C1887 VP.n31 VSUBS 0.028898f
C1888 VP.n32 VSUBS 0.028898f
C1889 VP.n33 VSUBS 0.053588f
C1890 VP.n34 VSUBS 0.039302f
C1891 VP.n35 VSUBS 1.2982f
C1892 VP.n36 VSUBS 1.82196f
C1893 VP.n37 VSUBS 1.84104f
C1894 VP.n38 VSUBS 0.038096f
C1895 VP.n39 VSUBS 0.039302f
C1896 VP.n40 VSUBS 0.053588f
C1897 VP.n41 VSUBS 0.03641f
C1898 VP.n42 VSUBS 0.028898f
C1899 VP.n43 VSUBS 0.028898f
C1900 VP.n44 VSUBS 0.028898f
C1901 VP.n45 VSUBS 0.053588f
C1902 VP.n46 VSUBS 0.031895f
C1903 VP.n47 VSUBS 1.2041f
C1904 VP.n48 VSUBS 0.048826f
C1905 VP.n49 VSUBS 0.028898f
C1906 VP.n50 VSUBS 0.028898f
C1907 VP.n51 VSUBS 0.028898f
C1908 VP.n52 VSUBS 0.02334f
C1909 VP.n53 VSUBS 0.057131f
C1910 VP.n54 VSUBS 0.048826f
C1911 VP.n55 VSUBS 0.028898f
C1912 VP.n56 VSUBS 0.028898f
C1913 VP.n57 VSUBS 0.031895f
C1914 VP.n58 VSUBS 0.053588f
C1915 VP.n59 VSUBS 0.047604f
C1916 VP.n60 VSUBS 0.028898f
C1917 VP.n61 VSUBS 0.028898f
C1918 VP.n62 VSUBS 0.028898f
C1919 VP.n63 VSUBS 0.053588f
C1920 VP.n64 VSUBS 0.039302f
C1921 VP.n65 VSUBS 1.2982f
C1922 VP.n66 VSUBS 0.045084f
.ends

