* NGSPICE file created from diff_pair_sample_1580.ext - technology: sky130A

.subckt diff_pair_sample_1580 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t15 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=1.04115 ps=6.64 w=6.31 l=2.02
X1 VDD2.t9 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X2 B.t23 B.t21 B.t22 B.t15 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=0 ps=0 w=6.31 l=2.02
X3 B.t20 B.t18 B.t19 B.t11 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=0 ps=0 w=6.31 l=2.02
X4 VTAIL.t8 VN.t1 VDD2.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X5 VDD1.t8 VP.t1 VTAIL.t18 B.t5 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=2.4609 ps=13.4 w=6.31 l=2.02
X6 VDD1.t7 VP.t2 VTAIL.t17 B.t1 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X7 VDD1.t6 VP.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X8 VTAIL.t10 VP.t4 VDD1.t5 B.t8 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X9 VTAIL.t6 VN.t2 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X10 VDD2.t6 VN.t3 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=1.04115 ps=6.64 w=6.31 l=2.02
X11 VTAIL.t4 VN.t4 VDD2.t5 B.t4 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X12 VTAIL.t13 VP.t5 VDD1.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X13 VTAIL.t11 VP.t6 VDD1.t3 B.t6 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X14 VDD2.t4 VN.t5 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=2.4609 ps=13.4 w=6.31 l=2.02
X15 VTAIL.t16 VP.t7 VDD1.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X16 VDD1.t1 VP.t8 VTAIL.t19 B.t9 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=2.4609 ps=13.4 w=6.31 l=2.02
X17 B.t17 B.t14 B.t16 B.t15 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=0 ps=0 w=6.31 l=2.02
X18 VDD1.t0 VP.t9 VTAIL.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=1.04115 ps=6.64 w=6.31 l=2.02
X19 VDD2.t3 VN.t6 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=2.4609 ps=13.4 w=6.31 l=2.02
X20 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=0 ps=0 w=6.31 l=2.02
X21 VDD2.t2 VN.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.4609 pd=13.4 as=1.04115 ps=6.64 w=6.31 l=2.02
X22 VTAIL.t0 VN.t8 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
X23 VDD2.t0 VN.t9 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.04115 pd=6.64 as=1.04115 ps=6.64 w=6.31 l=2.02
R0 VP.n20 VP.n19 161.3
R1 VP.n21 VP.n16 161.3
R2 VP.n23 VP.n22 161.3
R3 VP.n24 VP.n15 161.3
R4 VP.n26 VP.n25 161.3
R5 VP.n28 VP.n14 161.3
R6 VP.n30 VP.n29 161.3
R7 VP.n31 VP.n13 161.3
R8 VP.n33 VP.n32 161.3
R9 VP.n34 VP.n12 161.3
R10 VP.n37 VP.n36 161.3
R11 VP.n38 VP.n11 161.3
R12 VP.n40 VP.n39 161.3
R13 VP.n41 VP.n10 161.3
R14 VP.n74 VP.n0 161.3
R15 VP.n73 VP.n72 161.3
R16 VP.n71 VP.n1 161.3
R17 VP.n70 VP.n69 161.3
R18 VP.n67 VP.n2 161.3
R19 VP.n66 VP.n65 161.3
R20 VP.n64 VP.n3 161.3
R21 VP.n63 VP.n62 161.3
R22 VP.n61 VP.n4 161.3
R23 VP.n59 VP.n58 161.3
R24 VP.n57 VP.n5 161.3
R25 VP.n56 VP.n55 161.3
R26 VP.n54 VP.n6 161.3
R27 VP.n53 VP.n52 161.3
R28 VP.n51 VP.n50 161.3
R29 VP.n49 VP.n8 161.3
R30 VP.n48 VP.n47 161.3
R31 VP.n46 VP.n9 161.3
R32 VP.n18 VP.t0 106.01
R33 VP.n45 VP.n44 88.7361
R34 VP.n76 VP.n75 88.7361
R35 VP.n43 VP.n42 88.7361
R36 VP.n44 VP.t9 75.2832
R37 VP.n7 VP.t6 75.2832
R38 VP.n60 VP.t2 75.2832
R39 VP.n68 VP.t5 75.2832
R40 VP.n75 VP.t1 75.2832
R41 VP.n42 VP.t8 75.2832
R42 VP.n35 VP.t7 75.2832
R43 VP.n27 VP.t3 75.2832
R44 VP.n17 VP.t4 75.2832
R45 VP.n18 VP.n17 65.1987
R46 VP.n49 VP.n48 56.5193
R47 VP.n73 VP.n1 56.5193
R48 VP.n40 VP.n11 56.5193
R49 VP.n55 VP.n5 47.7779
R50 VP.n62 VP.n3 47.7779
R51 VP.n29 VP.n13 47.7779
R52 VP.n22 VP.n15 47.7779
R53 VP.n45 VP.n43 45.7155
R54 VP.n55 VP.n54 33.2089
R55 VP.n66 VP.n3 33.2089
R56 VP.n33 VP.n13 33.2089
R57 VP.n22 VP.n21 33.2089
R58 VP.n48 VP.n9 24.4675
R59 VP.n50 VP.n49 24.4675
R60 VP.n54 VP.n53 24.4675
R61 VP.n59 VP.n5 24.4675
R62 VP.n62 VP.n61 24.4675
R63 VP.n67 VP.n66 24.4675
R64 VP.n69 VP.n1 24.4675
R65 VP.n74 VP.n73 24.4675
R66 VP.n41 VP.n40 24.4675
R67 VP.n34 VP.n33 24.4675
R68 VP.n36 VP.n11 24.4675
R69 VP.n26 VP.n15 24.4675
R70 VP.n29 VP.n28 24.4675
R71 VP.n21 VP.n20 24.4675
R72 VP.n44 VP.n9 22.0208
R73 VP.n75 VP.n74 22.0208
R74 VP.n42 VP.n41 22.0208
R75 VP.n50 VP.n7 19.5741
R76 VP.n69 VP.n68 19.5741
R77 VP.n36 VP.n35 19.5741
R78 VP.n19 VP.n18 13.0188
R79 VP.n60 VP.n59 12.234
R80 VP.n61 VP.n60 12.234
R81 VP.n27 VP.n26 12.234
R82 VP.n28 VP.n27 12.234
R83 VP.n53 VP.n7 4.8939
R84 VP.n68 VP.n67 4.8939
R85 VP.n35 VP.n34 4.8939
R86 VP.n20 VP.n17 4.8939
R87 VP.n43 VP.n10 0.278367
R88 VP.n46 VP.n45 0.278367
R89 VP.n76 VP.n0 0.278367
R90 VP.n19 VP.n16 0.189894
R91 VP.n23 VP.n16 0.189894
R92 VP.n24 VP.n23 0.189894
R93 VP.n25 VP.n24 0.189894
R94 VP.n25 VP.n14 0.189894
R95 VP.n30 VP.n14 0.189894
R96 VP.n31 VP.n30 0.189894
R97 VP.n32 VP.n31 0.189894
R98 VP.n32 VP.n12 0.189894
R99 VP.n37 VP.n12 0.189894
R100 VP.n38 VP.n37 0.189894
R101 VP.n39 VP.n38 0.189894
R102 VP.n39 VP.n10 0.189894
R103 VP.n47 VP.n46 0.189894
R104 VP.n47 VP.n8 0.189894
R105 VP.n51 VP.n8 0.189894
R106 VP.n52 VP.n51 0.189894
R107 VP.n52 VP.n6 0.189894
R108 VP.n56 VP.n6 0.189894
R109 VP.n57 VP.n56 0.189894
R110 VP.n58 VP.n57 0.189894
R111 VP.n58 VP.n4 0.189894
R112 VP.n63 VP.n4 0.189894
R113 VP.n64 VP.n63 0.189894
R114 VP.n65 VP.n64 0.189894
R115 VP.n65 VP.n2 0.189894
R116 VP.n70 VP.n2 0.189894
R117 VP.n71 VP.n70 0.189894
R118 VP.n72 VP.n71 0.189894
R119 VP.n72 VP.n0 0.189894
R120 VP VP.n76 0.153454
R121 VTAIL.n11 VTAIL.t5 52.0854
R122 VTAIL.n17 VTAIL.t9 52.0853
R123 VTAIL.n2 VTAIL.t18 52.0853
R124 VTAIL.n16 VTAIL.t19 52.0853
R125 VTAIL.n15 VTAIL.n14 48.9476
R126 VTAIL.n13 VTAIL.n12 48.9476
R127 VTAIL.n10 VTAIL.n9 48.9476
R128 VTAIL.n8 VTAIL.n7 48.9476
R129 VTAIL.n19 VTAIL.n18 48.9473
R130 VTAIL.n1 VTAIL.n0 48.9473
R131 VTAIL.n4 VTAIL.n3 48.9473
R132 VTAIL.n6 VTAIL.n5 48.9473
R133 VTAIL.n8 VTAIL.n6 21.8583
R134 VTAIL.n17 VTAIL.n16 19.8324
R135 VTAIL.n18 VTAIL.t2 3.13838
R136 VTAIL.n18 VTAIL.t4 3.13838
R137 VTAIL.n0 VTAIL.t3 3.13838
R138 VTAIL.n0 VTAIL.t8 3.13838
R139 VTAIL.n3 VTAIL.t17 3.13838
R140 VTAIL.n3 VTAIL.t13 3.13838
R141 VTAIL.n5 VTAIL.t14 3.13838
R142 VTAIL.n5 VTAIL.t11 3.13838
R143 VTAIL.n14 VTAIL.t12 3.13838
R144 VTAIL.n14 VTAIL.t16 3.13838
R145 VTAIL.n12 VTAIL.t15 3.13838
R146 VTAIL.n12 VTAIL.t10 3.13838
R147 VTAIL.n9 VTAIL.t1 3.13838
R148 VTAIL.n9 VTAIL.t0 3.13838
R149 VTAIL.n7 VTAIL.t7 3.13838
R150 VTAIL.n7 VTAIL.t6 3.13838
R151 VTAIL.n10 VTAIL.n8 2.02636
R152 VTAIL.n11 VTAIL.n10 2.02636
R153 VTAIL.n15 VTAIL.n13 2.02636
R154 VTAIL.n16 VTAIL.n15 2.02636
R155 VTAIL.n6 VTAIL.n4 2.02636
R156 VTAIL.n4 VTAIL.n2 2.02636
R157 VTAIL.n19 VTAIL.n17 2.02636
R158 VTAIL VTAIL.n1 1.57809
R159 VTAIL.n13 VTAIL.n11 1.48326
R160 VTAIL.n2 VTAIL.n1 1.48326
R161 VTAIL VTAIL.n19 0.448776
R162 VDD1.n1 VDD1.t9 70.79
R163 VDD1.n3 VDD1.t0 70.7899
R164 VDD1.n5 VDD1.n4 67.0902
R165 VDD1.n1 VDD1.n0 65.6264
R166 VDD1.n7 VDD1.n6 65.6262
R167 VDD1.n3 VDD1.n2 65.6261
R168 VDD1.n7 VDD1.n5 40.3737
R169 VDD1.n6 VDD1.t2 3.13838
R170 VDD1.n6 VDD1.t1 3.13838
R171 VDD1.n0 VDD1.t5 3.13838
R172 VDD1.n0 VDD1.t6 3.13838
R173 VDD1.n4 VDD1.t4 3.13838
R174 VDD1.n4 VDD1.t8 3.13838
R175 VDD1.n2 VDD1.t3 3.13838
R176 VDD1.n2 VDD1.t7 3.13838
R177 VDD1 VDD1.n7 1.46171
R178 VDD1 VDD1.n1 0.565155
R179 VDD1.n5 VDD1.n3 0.451619
R180 B.n704 B.n703 585
R181 B.n705 B.n704 585
R182 B.n242 B.n121 585
R183 B.n241 B.n240 585
R184 B.n239 B.n238 585
R185 B.n237 B.n236 585
R186 B.n235 B.n234 585
R187 B.n233 B.n232 585
R188 B.n231 B.n230 585
R189 B.n229 B.n228 585
R190 B.n227 B.n226 585
R191 B.n225 B.n224 585
R192 B.n223 B.n222 585
R193 B.n221 B.n220 585
R194 B.n219 B.n218 585
R195 B.n217 B.n216 585
R196 B.n215 B.n214 585
R197 B.n213 B.n212 585
R198 B.n211 B.n210 585
R199 B.n209 B.n208 585
R200 B.n207 B.n206 585
R201 B.n205 B.n204 585
R202 B.n203 B.n202 585
R203 B.n201 B.n200 585
R204 B.n199 B.n198 585
R205 B.n197 B.n196 585
R206 B.n195 B.n194 585
R207 B.n193 B.n192 585
R208 B.n191 B.n190 585
R209 B.n189 B.n188 585
R210 B.n187 B.n186 585
R211 B.n185 B.n184 585
R212 B.n183 B.n182 585
R213 B.n181 B.n180 585
R214 B.n179 B.n178 585
R215 B.n176 B.n175 585
R216 B.n174 B.n173 585
R217 B.n172 B.n171 585
R218 B.n170 B.n169 585
R219 B.n168 B.n167 585
R220 B.n166 B.n165 585
R221 B.n164 B.n163 585
R222 B.n162 B.n161 585
R223 B.n160 B.n159 585
R224 B.n158 B.n157 585
R225 B.n156 B.n155 585
R226 B.n154 B.n153 585
R227 B.n152 B.n151 585
R228 B.n150 B.n149 585
R229 B.n148 B.n147 585
R230 B.n146 B.n145 585
R231 B.n144 B.n143 585
R232 B.n142 B.n141 585
R233 B.n140 B.n139 585
R234 B.n138 B.n137 585
R235 B.n136 B.n135 585
R236 B.n134 B.n133 585
R237 B.n132 B.n131 585
R238 B.n130 B.n129 585
R239 B.n128 B.n127 585
R240 B.n702 B.n91 585
R241 B.n706 B.n91 585
R242 B.n701 B.n90 585
R243 B.n707 B.n90 585
R244 B.n700 B.n699 585
R245 B.n699 B.n86 585
R246 B.n698 B.n85 585
R247 B.n713 B.n85 585
R248 B.n697 B.n84 585
R249 B.n714 B.n84 585
R250 B.n696 B.n83 585
R251 B.n715 B.n83 585
R252 B.n695 B.n694 585
R253 B.n694 B.n82 585
R254 B.n693 B.n78 585
R255 B.n721 B.n78 585
R256 B.n692 B.n77 585
R257 B.n722 B.n77 585
R258 B.n691 B.n76 585
R259 B.n723 B.n76 585
R260 B.n690 B.n689 585
R261 B.n689 B.n72 585
R262 B.n688 B.n71 585
R263 B.n729 B.n71 585
R264 B.n687 B.n70 585
R265 B.n730 B.n70 585
R266 B.n686 B.n69 585
R267 B.n731 B.n69 585
R268 B.n685 B.n684 585
R269 B.n684 B.n65 585
R270 B.n683 B.n64 585
R271 B.n737 B.n64 585
R272 B.n682 B.n63 585
R273 B.n738 B.n63 585
R274 B.n681 B.n62 585
R275 B.n739 B.n62 585
R276 B.n680 B.n679 585
R277 B.n679 B.n58 585
R278 B.n678 B.n57 585
R279 B.n745 B.n57 585
R280 B.n677 B.n56 585
R281 B.n746 B.n56 585
R282 B.n676 B.n55 585
R283 B.n747 B.n55 585
R284 B.n675 B.n674 585
R285 B.n674 B.n51 585
R286 B.n673 B.n50 585
R287 B.n753 B.n50 585
R288 B.n672 B.n49 585
R289 B.n754 B.n49 585
R290 B.n671 B.n48 585
R291 B.n755 B.n48 585
R292 B.n670 B.n669 585
R293 B.n669 B.n44 585
R294 B.n668 B.n43 585
R295 B.n761 B.n43 585
R296 B.n667 B.n42 585
R297 B.n762 B.n42 585
R298 B.n666 B.n41 585
R299 B.n763 B.n41 585
R300 B.n665 B.n664 585
R301 B.n664 B.n40 585
R302 B.n663 B.n36 585
R303 B.n769 B.n36 585
R304 B.n662 B.n35 585
R305 B.n770 B.n35 585
R306 B.n661 B.n34 585
R307 B.n771 B.n34 585
R308 B.n660 B.n659 585
R309 B.n659 B.n30 585
R310 B.n658 B.n29 585
R311 B.n777 B.n29 585
R312 B.n657 B.n28 585
R313 B.n778 B.n28 585
R314 B.n656 B.n27 585
R315 B.n779 B.n27 585
R316 B.n655 B.n654 585
R317 B.n654 B.n23 585
R318 B.n653 B.n22 585
R319 B.n785 B.n22 585
R320 B.n652 B.n21 585
R321 B.n786 B.n21 585
R322 B.n651 B.n20 585
R323 B.n787 B.n20 585
R324 B.n650 B.n649 585
R325 B.n649 B.n16 585
R326 B.n648 B.n15 585
R327 B.n793 B.n15 585
R328 B.n647 B.n14 585
R329 B.n794 B.n14 585
R330 B.n646 B.n13 585
R331 B.n795 B.n13 585
R332 B.n645 B.n644 585
R333 B.n644 B.n12 585
R334 B.n643 B.n642 585
R335 B.n643 B.n8 585
R336 B.n641 B.n7 585
R337 B.n802 B.n7 585
R338 B.n640 B.n6 585
R339 B.n803 B.n6 585
R340 B.n639 B.n5 585
R341 B.n804 B.n5 585
R342 B.n638 B.n637 585
R343 B.n637 B.n4 585
R344 B.n636 B.n243 585
R345 B.n636 B.n635 585
R346 B.n626 B.n244 585
R347 B.n245 B.n244 585
R348 B.n628 B.n627 585
R349 B.n629 B.n628 585
R350 B.n625 B.n249 585
R351 B.n253 B.n249 585
R352 B.n624 B.n623 585
R353 B.n623 B.n622 585
R354 B.n251 B.n250 585
R355 B.n252 B.n251 585
R356 B.n615 B.n614 585
R357 B.n616 B.n615 585
R358 B.n613 B.n258 585
R359 B.n258 B.n257 585
R360 B.n612 B.n611 585
R361 B.n611 B.n610 585
R362 B.n260 B.n259 585
R363 B.n261 B.n260 585
R364 B.n603 B.n602 585
R365 B.n604 B.n603 585
R366 B.n601 B.n266 585
R367 B.n266 B.n265 585
R368 B.n600 B.n599 585
R369 B.n599 B.n598 585
R370 B.n268 B.n267 585
R371 B.n269 B.n268 585
R372 B.n591 B.n590 585
R373 B.n592 B.n591 585
R374 B.n589 B.n274 585
R375 B.n274 B.n273 585
R376 B.n588 B.n587 585
R377 B.n587 B.n586 585
R378 B.n276 B.n275 585
R379 B.n579 B.n276 585
R380 B.n578 B.n577 585
R381 B.n580 B.n578 585
R382 B.n576 B.n281 585
R383 B.n281 B.n280 585
R384 B.n575 B.n574 585
R385 B.n574 B.n573 585
R386 B.n283 B.n282 585
R387 B.n284 B.n283 585
R388 B.n566 B.n565 585
R389 B.n567 B.n566 585
R390 B.n564 B.n289 585
R391 B.n289 B.n288 585
R392 B.n563 B.n562 585
R393 B.n562 B.n561 585
R394 B.n291 B.n290 585
R395 B.n292 B.n291 585
R396 B.n554 B.n553 585
R397 B.n555 B.n554 585
R398 B.n552 B.n297 585
R399 B.n297 B.n296 585
R400 B.n551 B.n550 585
R401 B.n550 B.n549 585
R402 B.n299 B.n298 585
R403 B.n300 B.n299 585
R404 B.n542 B.n541 585
R405 B.n543 B.n542 585
R406 B.n540 B.n304 585
R407 B.n308 B.n304 585
R408 B.n539 B.n538 585
R409 B.n538 B.n537 585
R410 B.n306 B.n305 585
R411 B.n307 B.n306 585
R412 B.n530 B.n529 585
R413 B.n531 B.n530 585
R414 B.n528 B.n313 585
R415 B.n313 B.n312 585
R416 B.n527 B.n526 585
R417 B.n526 B.n525 585
R418 B.n315 B.n314 585
R419 B.n316 B.n315 585
R420 B.n518 B.n517 585
R421 B.n519 B.n518 585
R422 B.n516 B.n321 585
R423 B.n321 B.n320 585
R424 B.n515 B.n514 585
R425 B.n514 B.n513 585
R426 B.n323 B.n322 585
R427 B.n506 B.n323 585
R428 B.n505 B.n504 585
R429 B.n507 B.n505 585
R430 B.n503 B.n328 585
R431 B.n328 B.n327 585
R432 B.n502 B.n501 585
R433 B.n501 B.n500 585
R434 B.n330 B.n329 585
R435 B.n331 B.n330 585
R436 B.n493 B.n492 585
R437 B.n494 B.n493 585
R438 B.n491 B.n336 585
R439 B.n336 B.n335 585
R440 B.n485 B.n484 585
R441 B.n483 B.n367 585
R442 B.n482 B.n366 585
R443 B.n487 B.n366 585
R444 B.n481 B.n480 585
R445 B.n479 B.n478 585
R446 B.n477 B.n476 585
R447 B.n475 B.n474 585
R448 B.n473 B.n472 585
R449 B.n471 B.n470 585
R450 B.n469 B.n468 585
R451 B.n467 B.n466 585
R452 B.n465 B.n464 585
R453 B.n463 B.n462 585
R454 B.n461 B.n460 585
R455 B.n459 B.n458 585
R456 B.n457 B.n456 585
R457 B.n455 B.n454 585
R458 B.n453 B.n452 585
R459 B.n451 B.n450 585
R460 B.n449 B.n448 585
R461 B.n447 B.n446 585
R462 B.n445 B.n444 585
R463 B.n443 B.n442 585
R464 B.n441 B.n440 585
R465 B.n439 B.n438 585
R466 B.n437 B.n436 585
R467 B.n435 B.n434 585
R468 B.n433 B.n432 585
R469 B.n431 B.n430 585
R470 B.n429 B.n428 585
R471 B.n427 B.n426 585
R472 B.n425 B.n424 585
R473 B.n423 B.n422 585
R474 B.n421 B.n420 585
R475 B.n418 B.n417 585
R476 B.n416 B.n415 585
R477 B.n414 B.n413 585
R478 B.n412 B.n411 585
R479 B.n410 B.n409 585
R480 B.n408 B.n407 585
R481 B.n406 B.n405 585
R482 B.n404 B.n403 585
R483 B.n402 B.n401 585
R484 B.n400 B.n399 585
R485 B.n398 B.n397 585
R486 B.n396 B.n395 585
R487 B.n394 B.n393 585
R488 B.n392 B.n391 585
R489 B.n390 B.n389 585
R490 B.n388 B.n387 585
R491 B.n386 B.n385 585
R492 B.n384 B.n383 585
R493 B.n382 B.n381 585
R494 B.n380 B.n379 585
R495 B.n378 B.n377 585
R496 B.n376 B.n375 585
R497 B.n374 B.n373 585
R498 B.n338 B.n337 585
R499 B.n490 B.n489 585
R500 B.n334 B.n333 585
R501 B.n335 B.n334 585
R502 B.n496 B.n495 585
R503 B.n495 B.n494 585
R504 B.n497 B.n332 585
R505 B.n332 B.n331 585
R506 B.n499 B.n498 585
R507 B.n500 B.n499 585
R508 B.n326 B.n325 585
R509 B.n327 B.n326 585
R510 B.n509 B.n508 585
R511 B.n508 B.n507 585
R512 B.n510 B.n324 585
R513 B.n506 B.n324 585
R514 B.n512 B.n511 585
R515 B.n513 B.n512 585
R516 B.n319 B.n318 585
R517 B.n320 B.n319 585
R518 B.n521 B.n520 585
R519 B.n520 B.n519 585
R520 B.n522 B.n317 585
R521 B.n317 B.n316 585
R522 B.n524 B.n523 585
R523 B.n525 B.n524 585
R524 B.n311 B.n310 585
R525 B.n312 B.n311 585
R526 B.n533 B.n532 585
R527 B.n532 B.n531 585
R528 B.n534 B.n309 585
R529 B.n309 B.n307 585
R530 B.n536 B.n535 585
R531 B.n537 B.n536 585
R532 B.n303 B.n302 585
R533 B.n308 B.n303 585
R534 B.n545 B.n544 585
R535 B.n544 B.n543 585
R536 B.n546 B.n301 585
R537 B.n301 B.n300 585
R538 B.n548 B.n547 585
R539 B.n549 B.n548 585
R540 B.n295 B.n294 585
R541 B.n296 B.n295 585
R542 B.n557 B.n556 585
R543 B.n556 B.n555 585
R544 B.n558 B.n293 585
R545 B.n293 B.n292 585
R546 B.n560 B.n559 585
R547 B.n561 B.n560 585
R548 B.n287 B.n286 585
R549 B.n288 B.n287 585
R550 B.n569 B.n568 585
R551 B.n568 B.n567 585
R552 B.n570 B.n285 585
R553 B.n285 B.n284 585
R554 B.n572 B.n571 585
R555 B.n573 B.n572 585
R556 B.n279 B.n278 585
R557 B.n280 B.n279 585
R558 B.n582 B.n581 585
R559 B.n581 B.n580 585
R560 B.n583 B.n277 585
R561 B.n579 B.n277 585
R562 B.n585 B.n584 585
R563 B.n586 B.n585 585
R564 B.n272 B.n271 585
R565 B.n273 B.n272 585
R566 B.n594 B.n593 585
R567 B.n593 B.n592 585
R568 B.n595 B.n270 585
R569 B.n270 B.n269 585
R570 B.n597 B.n596 585
R571 B.n598 B.n597 585
R572 B.n264 B.n263 585
R573 B.n265 B.n264 585
R574 B.n606 B.n605 585
R575 B.n605 B.n604 585
R576 B.n607 B.n262 585
R577 B.n262 B.n261 585
R578 B.n609 B.n608 585
R579 B.n610 B.n609 585
R580 B.n256 B.n255 585
R581 B.n257 B.n256 585
R582 B.n618 B.n617 585
R583 B.n617 B.n616 585
R584 B.n619 B.n254 585
R585 B.n254 B.n252 585
R586 B.n621 B.n620 585
R587 B.n622 B.n621 585
R588 B.n248 B.n247 585
R589 B.n253 B.n248 585
R590 B.n631 B.n630 585
R591 B.n630 B.n629 585
R592 B.n632 B.n246 585
R593 B.n246 B.n245 585
R594 B.n634 B.n633 585
R595 B.n635 B.n634 585
R596 B.n3 B.n0 585
R597 B.n4 B.n3 585
R598 B.n801 B.n1 585
R599 B.n802 B.n801 585
R600 B.n800 B.n799 585
R601 B.n800 B.n8 585
R602 B.n798 B.n9 585
R603 B.n12 B.n9 585
R604 B.n797 B.n796 585
R605 B.n796 B.n795 585
R606 B.n11 B.n10 585
R607 B.n794 B.n11 585
R608 B.n792 B.n791 585
R609 B.n793 B.n792 585
R610 B.n790 B.n17 585
R611 B.n17 B.n16 585
R612 B.n789 B.n788 585
R613 B.n788 B.n787 585
R614 B.n19 B.n18 585
R615 B.n786 B.n19 585
R616 B.n784 B.n783 585
R617 B.n785 B.n784 585
R618 B.n782 B.n24 585
R619 B.n24 B.n23 585
R620 B.n781 B.n780 585
R621 B.n780 B.n779 585
R622 B.n26 B.n25 585
R623 B.n778 B.n26 585
R624 B.n776 B.n775 585
R625 B.n777 B.n776 585
R626 B.n774 B.n31 585
R627 B.n31 B.n30 585
R628 B.n773 B.n772 585
R629 B.n772 B.n771 585
R630 B.n33 B.n32 585
R631 B.n770 B.n33 585
R632 B.n768 B.n767 585
R633 B.n769 B.n768 585
R634 B.n766 B.n37 585
R635 B.n40 B.n37 585
R636 B.n765 B.n764 585
R637 B.n764 B.n763 585
R638 B.n39 B.n38 585
R639 B.n762 B.n39 585
R640 B.n760 B.n759 585
R641 B.n761 B.n760 585
R642 B.n758 B.n45 585
R643 B.n45 B.n44 585
R644 B.n757 B.n756 585
R645 B.n756 B.n755 585
R646 B.n47 B.n46 585
R647 B.n754 B.n47 585
R648 B.n752 B.n751 585
R649 B.n753 B.n752 585
R650 B.n750 B.n52 585
R651 B.n52 B.n51 585
R652 B.n749 B.n748 585
R653 B.n748 B.n747 585
R654 B.n54 B.n53 585
R655 B.n746 B.n54 585
R656 B.n744 B.n743 585
R657 B.n745 B.n744 585
R658 B.n742 B.n59 585
R659 B.n59 B.n58 585
R660 B.n741 B.n740 585
R661 B.n740 B.n739 585
R662 B.n61 B.n60 585
R663 B.n738 B.n61 585
R664 B.n736 B.n735 585
R665 B.n737 B.n736 585
R666 B.n734 B.n66 585
R667 B.n66 B.n65 585
R668 B.n733 B.n732 585
R669 B.n732 B.n731 585
R670 B.n68 B.n67 585
R671 B.n730 B.n68 585
R672 B.n728 B.n727 585
R673 B.n729 B.n728 585
R674 B.n726 B.n73 585
R675 B.n73 B.n72 585
R676 B.n725 B.n724 585
R677 B.n724 B.n723 585
R678 B.n75 B.n74 585
R679 B.n722 B.n75 585
R680 B.n720 B.n719 585
R681 B.n721 B.n720 585
R682 B.n718 B.n79 585
R683 B.n82 B.n79 585
R684 B.n717 B.n716 585
R685 B.n716 B.n715 585
R686 B.n81 B.n80 585
R687 B.n714 B.n81 585
R688 B.n712 B.n711 585
R689 B.n713 B.n712 585
R690 B.n710 B.n87 585
R691 B.n87 B.n86 585
R692 B.n709 B.n708 585
R693 B.n708 B.n707 585
R694 B.n89 B.n88 585
R695 B.n706 B.n89 585
R696 B.n805 B.n804 585
R697 B.n803 B.n2 585
R698 B.n127 B.n89 540.549
R699 B.n704 B.n91 540.549
R700 B.n489 B.n336 540.549
R701 B.n485 B.n334 540.549
R702 B.n125 B.t21 282.248
R703 B.n122 B.t14 282.248
R704 B.n371 B.t10 282.248
R705 B.n368 B.t18 282.248
R706 B.n705 B.n120 256.663
R707 B.n705 B.n119 256.663
R708 B.n705 B.n118 256.663
R709 B.n705 B.n117 256.663
R710 B.n705 B.n116 256.663
R711 B.n705 B.n115 256.663
R712 B.n705 B.n114 256.663
R713 B.n705 B.n113 256.663
R714 B.n705 B.n112 256.663
R715 B.n705 B.n111 256.663
R716 B.n705 B.n110 256.663
R717 B.n705 B.n109 256.663
R718 B.n705 B.n108 256.663
R719 B.n705 B.n107 256.663
R720 B.n705 B.n106 256.663
R721 B.n705 B.n105 256.663
R722 B.n705 B.n104 256.663
R723 B.n705 B.n103 256.663
R724 B.n705 B.n102 256.663
R725 B.n705 B.n101 256.663
R726 B.n705 B.n100 256.663
R727 B.n705 B.n99 256.663
R728 B.n705 B.n98 256.663
R729 B.n705 B.n97 256.663
R730 B.n705 B.n96 256.663
R731 B.n705 B.n95 256.663
R732 B.n705 B.n94 256.663
R733 B.n705 B.n93 256.663
R734 B.n705 B.n92 256.663
R735 B.n487 B.n486 256.663
R736 B.n487 B.n339 256.663
R737 B.n487 B.n340 256.663
R738 B.n487 B.n341 256.663
R739 B.n487 B.n342 256.663
R740 B.n487 B.n343 256.663
R741 B.n487 B.n344 256.663
R742 B.n487 B.n345 256.663
R743 B.n487 B.n346 256.663
R744 B.n487 B.n347 256.663
R745 B.n487 B.n348 256.663
R746 B.n487 B.n349 256.663
R747 B.n487 B.n350 256.663
R748 B.n487 B.n351 256.663
R749 B.n487 B.n352 256.663
R750 B.n487 B.n353 256.663
R751 B.n487 B.n354 256.663
R752 B.n487 B.n355 256.663
R753 B.n487 B.n356 256.663
R754 B.n487 B.n357 256.663
R755 B.n487 B.n358 256.663
R756 B.n487 B.n359 256.663
R757 B.n487 B.n360 256.663
R758 B.n487 B.n361 256.663
R759 B.n487 B.n362 256.663
R760 B.n487 B.n363 256.663
R761 B.n487 B.n364 256.663
R762 B.n487 B.n365 256.663
R763 B.n488 B.n487 256.663
R764 B.n807 B.n806 256.663
R765 B.n131 B.n130 163.367
R766 B.n135 B.n134 163.367
R767 B.n139 B.n138 163.367
R768 B.n143 B.n142 163.367
R769 B.n147 B.n146 163.367
R770 B.n151 B.n150 163.367
R771 B.n155 B.n154 163.367
R772 B.n159 B.n158 163.367
R773 B.n163 B.n162 163.367
R774 B.n167 B.n166 163.367
R775 B.n171 B.n170 163.367
R776 B.n175 B.n174 163.367
R777 B.n180 B.n179 163.367
R778 B.n184 B.n183 163.367
R779 B.n188 B.n187 163.367
R780 B.n192 B.n191 163.367
R781 B.n196 B.n195 163.367
R782 B.n200 B.n199 163.367
R783 B.n204 B.n203 163.367
R784 B.n208 B.n207 163.367
R785 B.n212 B.n211 163.367
R786 B.n216 B.n215 163.367
R787 B.n220 B.n219 163.367
R788 B.n224 B.n223 163.367
R789 B.n228 B.n227 163.367
R790 B.n232 B.n231 163.367
R791 B.n236 B.n235 163.367
R792 B.n240 B.n239 163.367
R793 B.n704 B.n121 163.367
R794 B.n493 B.n336 163.367
R795 B.n493 B.n330 163.367
R796 B.n501 B.n330 163.367
R797 B.n501 B.n328 163.367
R798 B.n505 B.n328 163.367
R799 B.n505 B.n323 163.367
R800 B.n514 B.n323 163.367
R801 B.n514 B.n321 163.367
R802 B.n518 B.n321 163.367
R803 B.n518 B.n315 163.367
R804 B.n526 B.n315 163.367
R805 B.n526 B.n313 163.367
R806 B.n530 B.n313 163.367
R807 B.n530 B.n306 163.367
R808 B.n538 B.n306 163.367
R809 B.n538 B.n304 163.367
R810 B.n542 B.n304 163.367
R811 B.n542 B.n299 163.367
R812 B.n550 B.n299 163.367
R813 B.n550 B.n297 163.367
R814 B.n554 B.n297 163.367
R815 B.n554 B.n291 163.367
R816 B.n562 B.n291 163.367
R817 B.n562 B.n289 163.367
R818 B.n566 B.n289 163.367
R819 B.n566 B.n283 163.367
R820 B.n574 B.n283 163.367
R821 B.n574 B.n281 163.367
R822 B.n578 B.n281 163.367
R823 B.n578 B.n276 163.367
R824 B.n587 B.n276 163.367
R825 B.n587 B.n274 163.367
R826 B.n591 B.n274 163.367
R827 B.n591 B.n268 163.367
R828 B.n599 B.n268 163.367
R829 B.n599 B.n266 163.367
R830 B.n603 B.n266 163.367
R831 B.n603 B.n260 163.367
R832 B.n611 B.n260 163.367
R833 B.n611 B.n258 163.367
R834 B.n615 B.n258 163.367
R835 B.n615 B.n251 163.367
R836 B.n623 B.n251 163.367
R837 B.n623 B.n249 163.367
R838 B.n628 B.n249 163.367
R839 B.n628 B.n244 163.367
R840 B.n636 B.n244 163.367
R841 B.n637 B.n636 163.367
R842 B.n637 B.n5 163.367
R843 B.n6 B.n5 163.367
R844 B.n7 B.n6 163.367
R845 B.n643 B.n7 163.367
R846 B.n644 B.n643 163.367
R847 B.n644 B.n13 163.367
R848 B.n14 B.n13 163.367
R849 B.n15 B.n14 163.367
R850 B.n649 B.n15 163.367
R851 B.n649 B.n20 163.367
R852 B.n21 B.n20 163.367
R853 B.n22 B.n21 163.367
R854 B.n654 B.n22 163.367
R855 B.n654 B.n27 163.367
R856 B.n28 B.n27 163.367
R857 B.n29 B.n28 163.367
R858 B.n659 B.n29 163.367
R859 B.n659 B.n34 163.367
R860 B.n35 B.n34 163.367
R861 B.n36 B.n35 163.367
R862 B.n664 B.n36 163.367
R863 B.n664 B.n41 163.367
R864 B.n42 B.n41 163.367
R865 B.n43 B.n42 163.367
R866 B.n669 B.n43 163.367
R867 B.n669 B.n48 163.367
R868 B.n49 B.n48 163.367
R869 B.n50 B.n49 163.367
R870 B.n674 B.n50 163.367
R871 B.n674 B.n55 163.367
R872 B.n56 B.n55 163.367
R873 B.n57 B.n56 163.367
R874 B.n679 B.n57 163.367
R875 B.n679 B.n62 163.367
R876 B.n63 B.n62 163.367
R877 B.n64 B.n63 163.367
R878 B.n684 B.n64 163.367
R879 B.n684 B.n69 163.367
R880 B.n70 B.n69 163.367
R881 B.n71 B.n70 163.367
R882 B.n689 B.n71 163.367
R883 B.n689 B.n76 163.367
R884 B.n77 B.n76 163.367
R885 B.n78 B.n77 163.367
R886 B.n694 B.n78 163.367
R887 B.n694 B.n83 163.367
R888 B.n84 B.n83 163.367
R889 B.n85 B.n84 163.367
R890 B.n699 B.n85 163.367
R891 B.n699 B.n90 163.367
R892 B.n91 B.n90 163.367
R893 B.n367 B.n366 163.367
R894 B.n480 B.n366 163.367
R895 B.n478 B.n477 163.367
R896 B.n474 B.n473 163.367
R897 B.n470 B.n469 163.367
R898 B.n466 B.n465 163.367
R899 B.n462 B.n461 163.367
R900 B.n458 B.n457 163.367
R901 B.n454 B.n453 163.367
R902 B.n450 B.n449 163.367
R903 B.n446 B.n445 163.367
R904 B.n442 B.n441 163.367
R905 B.n438 B.n437 163.367
R906 B.n434 B.n433 163.367
R907 B.n430 B.n429 163.367
R908 B.n426 B.n425 163.367
R909 B.n422 B.n421 163.367
R910 B.n417 B.n416 163.367
R911 B.n413 B.n412 163.367
R912 B.n409 B.n408 163.367
R913 B.n405 B.n404 163.367
R914 B.n401 B.n400 163.367
R915 B.n397 B.n396 163.367
R916 B.n393 B.n392 163.367
R917 B.n389 B.n388 163.367
R918 B.n385 B.n384 163.367
R919 B.n381 B.n380 163.367
R920 B.n377 B.n376 163.367
R921 B.n373 B.n338 163.367
R922 B.n495 B.n334 163.367
R923 B.n495 B.n332 163.367
R924 B.n499 B.n332 163.367
R925 B.n499 B.n326 163.367
R926 B.n508 B.n326 163.367
R927 B.n508 B.n324 163.367
R928 B.n512 B.n324 163.367
R929 B.n512 B.n319 163.367
R930 B.n520 B.n319 163.367
R931 B.n520 B.n317 163.367
R932 B.n524 B.n317 163.367
R933 B.n524 B.n311 163.367
R934 B.n532 B.n311 163.367
R935 B.n532 B.n309 163.367
R936 B.n536 B.n309 163.367
R937 B.n536 B.n303 163.367
R938 B.n544 B.n303 163.367
R939 B.n544 B.n301 163.367
R940 B.n548 B.n301 163.367
R941 B.n548 B.n295 163.367
R942 B.n556 B.n295 163.367
R943 B.n556 B.n293 163.367
R944 B.n560 B.n293 163.367
R945 B.n560 B.n287 163.367
R946 B.n568 B.n287 163.367
R947 B.n568 B.n285 163.367
R948 B.n572 B.n285 163.367
R949 B.n572 B.n279 163.367
R950 B.n581 B.n279 163.367
R951 B.n581 B.n277 163.367
R952 B.n585 B.n277 163.367
R953 B.n585 B.n272 163.367
R954 B.n593 B.n272 163.367
R955 B.n593 B.n270 163.367
R956 B.n597 B.n270 163.367
R957 B.n597 B.n264 163.367
R958 B.n605 B.n264 163.367
R959 B.n605 B.n262 163.367
R960 B.n609 B.n262 163.367
R961 B.n609 B.n256 163.367
R962 B.n617 B.n256 163.367
R963 B.n617 B.n254 163.367
R964 B.n621 B.n254 163.367
R965 B.n621 B.n248 163.367
R966 B.n630 B.n248 163.367
R967 B.n630 B.n246 163.367
R968 B.n634 B.n246 163.367
R969 B.n634 B.n3 163.367
R970 B.n805 B.n3 163.367
R971 B.n801 B.n2 163.367
R972 B.n801 B.n800 163.367
R973 B.n800 B.n9 163.367
R974 B.n796 B.n9 163.367
R975 B.n796 B.n11 163.367
R976 B.n792 B.n11 163.367
R977 B.n792 B.n17 163.367
R978 B.n788 B.n17 163.367
R979 B.n788 B.n19 163.367
R980 B.n784 B.n19 163.367
R981 B.n784 B.n24 163.367
R982 B.n780 B.n24 163.367
R983 B.n780 B.n26 163.367
R984 B.n776 B.n26 163.367
R985 B.n776 B.n31 163.367
R986 B.n772 B.n31 163.367
R987 B.n772 B.n33 163.367
R988 B.n768 B.n33 163.367
R989 B.n768 B.n37 163.367
R990 B.n764 B.n37 163.367
R991 B.n764 B.n39 163.367
R992 B.n760 B.n39 163.367
R993 B.n760 B.n45 163.367
R994 B.n756 B.n45 163.367
R995 B.n756 B.n47 163.367
R996 B.n752 B.n47 163.367
R997 B.n752 B.n52 163.367
R998 B.n748 B.n52 163.367
R999 B.n748 B.n54 163.367
R1000 B.n744 B.n54 163.367
R1001 B.n744 B.n59 163.367
R1002 B.n740 B.n59 163.367
R1003 B.n740 B.n61 163.367
R1004 B.n736 B.n61 163.367
R1005 B.n736 B.n66 163.367
R1006 B.n732 B.n66 163.367
R1007 B.n732 B.n68 163.367
R1008 B.n728 B.n68 163.367
R1009 B.n728 B.n73 163.367
R1010 B.n724 B.n73 163.367
R1011 B.n724 B.n75 163.367
R1012 B.n720 B.n75 163.367
R1013 B.n720 B.n79 163.367
R1014 B.n716 B.n79 163.367
R1015 B.n716 B.n81 163.367
R1016 B.n712 B.n81 163.367
R1017 B.n712 B.n87 163.367
R1018 B.n708 B.n87 163.367
R1019 B.n708 B.n89 163.367
R1020 B.n487 B.n335 122.487
R1021 B.n706 B.n705 122.487
R1022 B.n122 B.t16 118.541
R1023 B.n371 B.t13 118.541
R1024 B.n125 B.t22 118.534
R1025 B.n368 B.t20 118.534
R1026 B.n123 B.t17 72.9658
R1027 B.n372 B.t12 72.9658
R1028 B.n126 B.t23 72.9591
R1029 B.n369 B.t19 72.9591
R1030 B.n127 B.n92 71.676
R1031 B.n131 B.n93 71.676
R1032 B.n135 B.n94 71.676
R1033 B.n139 B.n95 71.676
R1034 B.n143 B.n96 71.676
R1035 B.n147 B.n97 71.676
R1036 B.n151 B.n98 71.676
R1037 B.n155 B.n99 71.676
R1038 B.n159 B.n100 71.676
R1039 B.n163 B.n101 71.676
R1040 B.n167 B.n102 71.676
R1041 B.n171 B.n103 71.676
R1042 B.n175 B.n104 71.676
R1043 B.n180 B.n105 71.676
R1044 B.n184 B.n106 71.676
R1045 B.n188 B.n107 71.676
R1046 B.n192 B.n108 71.676
R1047 B.n196 B.n109 71.676
R1048 B.n200 B.n110 71.676
R1049 B.n204 B.n111 71.676
R1050 B.n208 B.n112 71.676
R1051 B.n212 B.n113 71.676
R1052 B.n216 B.n114 71.676
R1053 B.n220 B.n115 71.676
R1054 B.n224 B.n116 71.676
R1055 B.n228 B.n117 71.676
R1056 B.n232 B.n118 71.676
R1057 B.n236 B.n119 71.676
R1058 B.n240 B.n120 71.676
R1059 B.n121 B.n120 71.676
R1060 B.n239 B.n119 71.676
R1061 B.n235 B.n118 71.676
R1062 B.n231 B.n117 71.676
R1063 B.n227 B.n116 71.676
R1064 B.n223 B.n115 71.676
R1065 B.n219 B.n114 71.676
R1066 B.n215 B.n113 71.676
R1067 B.n211 B.n112 71.676
R1068 B.n207 B.n111 71.676
R1069 B.n203 B.n110 71.676
R1070 B.n199 B.n109 71.676
R1071 B.n195 B.n108 71.676
R1072 B.n191 B.n107 71.676
R1073 B.n187 B.n106 71.676
R1074 B.n183 B.n105 71.676
R1075 B.n179 B.n104 71.676
R1076 B.n174 B.n103 71.676
R1077 B.n170 B.n102 71.676
R1078 B.n166 B.n101 71.676
R1079 B.n162 B.n100 71.676
R1080 B.n158 B.n99 71.676
R1081 B.n154 B.n98 71.676
R1082 B.n150 B.n97 71.676
R1083 B.n146 B.n96 71.676
R1084 B.n142 B.n95 71.676
R1085 B.n138 B.n94 71.676
R1086 B.n134 B.n93 71.676
R1087 B.n130 B.n92 71.676
R1088 B.n486 B.n485 71.676
R1089 B.n480 B.n339 71.676
R1090 B.n477 B.n340 71.676
R1091 B.n473 B.n341 71.676
R1092 B.n469 B.n342 71.676
R1093 B.n465 B.n343 71.676
R1094 B.n461 B.n344 71.676
R1095 B.n457 B.n345 71.676
R1096 B.n453 B.n346 71.676
R1097 B.n449 B.n347 71.676
R1098 B.n445 B.n348 71.676
R1099 B.n441 B.n349 71.676
R1100 B.n437 B.n350 71.676
R1101 B.n433 B.n351 71.676
R1102 B.n429 B.n352 71.676
R1103 B.n425 B.n353 71.676
R1104 B.n421 B.n354 71.676
R1105 B.n416 B.n355 71.676
R1106 B.n412 B.n356 71.676
R1107 B.n408 B.n357 71.676
R1108 B.n404 B.n358 71.676
R1109 B.n400 B.n359 71.676
R1110 B.n396 B.n360 71.676
R1111 B.n392 B.n361 71.676
R1112 B.n388 B.n362 71.676
R1113 B.n384 B.n363 71.676
R1114 B.n380 B.n364 71.676
R1115 B.n376 B.n365 71.676
R1116 B.n488 B.n338 71.676
R1117 B.n486 B.n367 71.676
R1118 B.n478 B.n339 71.676
R1119 B.n474 B.n340 71.676
R1120 B.n470 B.n341 71.676
R1121 B.n466 B.n342 71.676
R1122 B.n462 B.n343 71.676
R1123 B.n458 B.n344 71.676
R1124 B.n454 B.n345 71.676
R1125 B.n450 B.n346 71.676
R1126 B.n446 B.n347 71.676
R1127 B.n442 B.n348 71.676
R1128 B.n438 B.n349 71.676
R1129 B.n434 B.n350 71.676
R1130 B.n430 B.n351 71.676
R1131 B.n426 B.n352 71.676
R1132 B.n422 B.n353 71.676
R1133 B.n417 B.n354 71.676
R1134 B.n413 B.n355 71.676
R1135 B.n409 B.n356 71.676
R1136 B.n405 B.n357 71.676
R1137 B.n401 B.n358 71.676
R1138 B.n397 B.n359 71.676
R1139 B.n393 B.n360 71.676
R1140 B.n389 B.n361 71.676
R1141 B.n385 B.n362 71.676
R1142 B.n381 B.n363 71.676
R1143 B.n377 B.n364 71.676
R1144 B.n373 B.n365 71.676
R1145 B.n489 B.n488 71.676
R1146 B.n806 B.n805 71.676
R1147 B.n806 B.n2 71.676
R1148 B.n494 B.n335 64.5668
R1149 B.n494 B.n331 64.5668
R1150 B.n500 B.n331 64.5668
R1151 B.n500 B.n327 64.5668
R1152 B.n507 B.n327 64.5668
R1153 B.n507 B.n506 64.5668
R1154 B.n513 B.n320 64.5668
R1155 B.n519 B.n320 64.5668
R1156 B.n519 B.n316 64.5668
R1157 B.n525 B.n316 64.5668
R1158 B.n525 B.n312 64.5668
R1159 B.n531 B.n312 64.5668
R1160 B.n531 B.n307 64.5668
R1161 B.n537 B.n307 64.5668
R1162 B.n537 B.n308 64.5668
R1163 B.n543 B.n300 64.5668
R1164 B.n549 B.n300 64.5668
R1165 B.n549 B.n296 64.5668
R1166 B.n555 B.n296 64.5668
R1167 B.n555 B.n292 64.5668
R1168 B.n561 B.n292 64.5668
R1169 B.n567 B.n288 64.5668
R1170 B.n567 B.n284 64.5668
R1171 B.n573 B.n284 64.5668
R1172 B.n573 B.n280 64.5668
R1173 B.n580 B.n280 64.5668
R1174 B.n580 B.n579 64.5668
R1175 B.n586 B.n273 64.5668
R1176 B.n592 B.n273 64.5668
R1177 B.n592 B.n269 64.5668
R1178 B.n598 B.n269 64.5668
R1179 B.n598 B.n265 64.5668
R1180 B.n604 B.n265 64.5668
R1181 B.n610 B.n261 64.5668
R1182 B.n610 B.n257 64.5668
R1183 B.n616 B.n257 64.5668
R1184 B.n616 B.n252 64.5668
R1185 B.n622 B.n252 64.5668
R1186 B.n622 B.n253 64.5668
R1187 B.n629 B.n245 64.5668
R1188 B.n635 B.n245 64.5668
R1189 B.n635 B.n4 64.5668
R1190 B.n804 B.n4 64.5668
R1191 B.n804 B.n803 64.5668
R1192 B.n803 B.n802 64.5668
R1193 B.n802 B.n8 64.5668
R1194 B.n12 B.n8 64.5668
R1195 B.n795 B.n12 64.5668
R1196 B.n794 B.n793 64.5668
R1197 B.n793 B.n16 64.5668
R1198 B.n787 B.n16 64.5668
R1199 B.n787 B.n786 64.5668
R1200 B.n786 B.n785 64.5668
R1201 B.n785 B.n23 64.5668
R1202 B.n779 B.n778 64.5668
R1203 B.n778 B.n777 64.5668
R1204 B.n777 B.n30 64.5668
R1205 B.n771 B.n30 64.5668
R1206 B.n771 B.n770 64.5668
R1207 B.n770 B.n769 64.5668
R1208 B.n763 B.n40 64.5668
R1209 B.n763 B.n762 64.5668
R1210 B.n762 B.n761 64.5668
R1211 B.n761 B.n44 64.5668
R1212 B.n755 B.n44 64.5668
R1213 B.n755 B.n754 64.5668
R1214 B.n753 B.n51 64.5668
R1215 B.n747 B.n51 64.5668
R1216 B.n747 B.n746 64.5668
R1217 B.n746 B.n745 64.5668
R1218 B.n745 B.n58 64.5668
R1219 B.n739 B.n58 64.5668
R1220 B.n738 B.n737 64.5668
R1221 B.n737 B.n65 64.5668
R1222 B.n731 B.n65 64.5668
R1223 B.n731 B.n730 64.5668
R1224 B.n730 B.n729 64.5668
R1225 B.n729 B.n72 64.5668
R1226 B.n723 B.n72 64.5668
R1227 B.n723 B.n722 64.5668
R1228 B.n722 B.n721 64.5668
R1229 B.n715 B.n82 64.5668
R1230 B.n715 B.n714 64.5668
R1231 B.n714 B.n713 64.5668
R1232 B.n713 B.n86 64.5668
R1233 B.n707 B.n86 64.5668
R1234 B.n707 B.n706 64.5668
R1235 B.n177 B.n126 59.5399
R1236 B.n124 B.n123 59.5399
R1237 B.n419 B.n372 59.5399
R1238 B.n370 B.n369 59.5399
R1239 B.n308 B.t7 51.2737
R1240 B.t9 B.n738 51.2737
R1241 B.n561 B.t6 45.5767
R1242 B.t4 B.n753 45.5767
R1243 B.n126 B.n125 45.5763
R1244 B.n123 B.n122 45.5763
R1245 B.n372 B.n371 45.5763
R1246 B.n369 B.n368 45.5763
R1247 B.n506 B.t11 43.6777
R1248 B.n82 B.t15 43.6777
R1249 B.n579 B.t1 39.8797
R1250 B.n40 B.t2 39.8797
R1251 B.n629 B.t5 36.0816
R1252 B.n795 B.t3 36.0816
R1253 B.n484 B.n333 35.1225
R1254 B.n491 B.n490 35.1225
R1255 B.n128 B.n88 35.1225
R1256 B.n703 B.n702 35.1224
R1257 B.n604 B.t0 34.1826
R1258 B.n779 B.t8 34.1826
R1259 B.t0 B.n261 30.3846
R1260 B.t8 B.n23 30.3846
R1261 B.n253 B.t5 28.4856
R1262 B.t3 B.n794 28.4856
R1263 B.n586 B.t1 24.6876
R1264 B.n769 B.t2 24.6876
R1265 B.n513 B.t11 20.8896
R1266 B.n721 B.t15 20.8896
R1267 B.t6 B.n288 18.9906
R1268 B.n754 B.t4 18.9906
R1269 B B.n807 18.0485
R1270 B.n543 B.t7 13.2936
R1271 B.n739 B.t9 13.2936
R1272 B.n496 B.n333 10.6151
R1273 B.n497 B.n496 10.6151
R1274 B.n498 B.n497 10.6151
R1275 B.n498 B.n325 10.6151
R1276 B.n509 B.n325 10.6151
R1277 B.n510 B.n509 10.6151
R1278 B.n511 B.n510 10.6151
R1279 B.n511 B.n318 10.6151
R1280 B.n521 B.n318 10.6151
R1281 B.n522 B.n521 10.6151
R1282 B.n523 B.n522 10.6151
R1283 B.n523 B.n310 10.6151
R1284 B.n533 B.n310 10.6151
R1285 B.n534 B.n533 10.6151
R1286 B.n535 B.n534 10.6151
R1287 B.n535 B.n302 10.6151
R1288 B.n545 B.n302 10.6151
R1289 B.n546 B.n545 10.6151
R1290 B.n547 B.n546 10.6151
R1291 B.n547 B.n294 10.6151
R1292 B.n557 B.n294 10.6151
R1293 B.n558 B.n557 10.6151
R1294 B.n559 B.n558 10.6151
R1295 B.n559 B.n286 10.6151
R1296 B.n569 B.n286 10.6151
R1297 B.n570 B.n569 10.6151
R1298 B.n571 B.n570 10.6151
R1299 B.n571 B.n278 10.6151
R1300 B.n582 B.n278 10.6151
R1301 B.n583 B.n582 10.6151
R1302 B.n584 B.n583 10.6151
R1303 B.n584 B.n271 10.6151
R1304 B.n594 B.n271 10.6151
R1305 B.n595 B.n594 10.6151
R1306 B.n596 B.n595 10.6151
R1307 B.n596 B.n263 10.6151
R1308 B.n606 B.n263 10.6151
R1309 B.n607 B.n606 10.6151
R1310 B.n608 B.n607 10.6151
R1311 B.n608 B.n255 10.6151
R1312 B.n618 B.n255 10.6151
R1313 B.n619 B.n618 10.6151
R1314 B.n620 B.n619 10.6151
R1315 B.n620 B.n247 10.6151
R1316 B.n631 B.n247 10.6151
R1317 B.n632 B.n631 10.6151
R1318 B.n633 B.n632 10.6151
R1319 B.n633 B.n0 10.6151
R1320 B.n484 B.n483 10.6151
R1321 B.n483 B.n482 10.6151
R1322 B.n482 B.n481 10.6151
R1323 B.n481 B.n479 10.6151
R1324 B.n479 B.n476 10.6151
R1325 B.n476 B.n475 10.6151
R1326 B.n475 B.n472 10.6151
R1327 B.n472 B.n471 10.6151
R1328 B.n471 B.n468 10.6151
R1329 B.n468 B.n467 10.6151
R1330 B.n467 B.n464 10.6151
R1331 B.n464 B.n463 10.6151
R1332 B.n463 B.n460 10.6151
R1333 B.n460 B.n459 10.6151
R1334 B.n459 B.n456 10.6151
R1335 B.n456 B.n455 10.6151
R1336 B.n455 B.n452 10.6151
R1337 B.n452 B.n451 10.6151
R1338 B.n451 B.n448 10.6151
R1339 B.n448 B.n447 10.6151
R1340 B.n447 B.n444 10.6151
R1341 B.n444 B.n443 10.6151
R1342 B.n443 B.n440 10.6151
R1343 B.n440 B.n439 10.6151
R1344 B.n436 B.n435 10.6151
R1345 B.n435 B.n432 10.6151
R1346 B.n432 B.n431 10.6151
R1347 B.n431 B.n428 10.6151
R1348 B.n428 B.n427 10.6151
R1349 B.n427 B.n424 10.6151
R1350 B.n424 B.n423 10.6151
R1351 B.n423 B.n420 10.6151
R1352 B.n418 B.n415 10.6151
R1353 B.n415 B.n414 10.6151
R1354 B.n414 B.n411 10.6151
R1355 B.n411 B.n410 10.6151
R1356 B.n410 B.n407 10.6151
R1357 B.n407 B.n406 10.6151
R1358 B.n406 B.n403 10.6151
R1359 B.n403 B.n402 10.6151
R1360 B.n402 B.n399 10.6151
R1361 B.n399 B.n398 10.6151
R1362 B.n398 B.n395 10.6151
R1363 B.n395 B.n394 10.6151
R1364 B.n394 B.n391 10.6151
R1365 B.n391 B.n390 10.6151
R1366 B.n390 B.n387 10.6151
R1367 B.n387 B.n386 10.6151
R1368 B.n386 B.n383 10.6151
R1369 B.n383 B.n382 10.6151
R1370 B.n382 B.n379 10.6151
R1371 B.n379 B.n378 10.6151
R1372 B.n378 B.n375 10.6151
R1373 B.n375 B.n374 10.6151
R1374 B.n374 B.n337 10.6151
R1375 B.n490 B.n337 10.6151
R1376 B.n492 B.n491 10.6151
R1377 B.n492 B.n329 10.6151
R1378 B.n502 B.n329 10.6151
R1379 B.n503 B.n502 10.6151
R1380 B.n504 B.n503 10.6151
R1381 B.n504 B.n322 10.6151
R1382 B.n515 B.n322 10.6151
R1383 B.n516 B.n515 10.6151
R1384 B.n517 B.n516 10.6151
R1385 B.n517 B.n314 10.6151
R1386 B.n527 B.n314 10.6151
R1387 B.n528 B.n527 10.6151
R1388 B.n529 B.n528 10.6151
R1389 B.n529 B.n305 10.6151
R1390 B.n539 B.n305 10.6151
R1391 B.n540 B.n539 10.6151
R1392 B.n541 B.n540 10.6151
R1393 B.n541 B.n298 10.6151
R1394 B.n551 B.n298 10.6151
R1395 B.n552 B.n551 10.6151
R1396 B.n553 B.n552 10.6151
R1397 B.n553 B.n290 10.6151
R1398 B.n563 B.n290 10.6151
R1399 B.n564 B.n563 10.6151
R1400 B.n565 B.n564 10.6151
R1401 B.n565 B.n282 10.6151
R1402 B.n575 B.n282 10.6151
R1403 B.n576 B.n575 10.6151
R1404 B.n577 B.n576 10.6151
R1405 B.n577 B.n275 10.6151
R1406 B.n588 B.n275 10.6151
R1407 B.n589 B.n588 10.6151
R1408 B.n590 B.n589 10.6151
R1409 B.n590 B.n267 10.6151
R1410 B.n600 B.n267 10.6151
R1411 B.n601 B.n600 10.6151
R1412 B.n602 B.n601 10.6151
R1413 B.n602 B.n259 10.6151
R1414 B.n612 B.n259 10.6151
R1415 B.n613 B.n612 10.6151
R1416 B.n614 B.n613 10.6151
R1417 B.n614 B.n250 10.6151
R1418 B.n624 B.n250 10.6151
R1419 B.n625 B.n624 10.6151
R1420 B.n627 B.n625 10.6151
R1421 B.n627 B.n626 10.6151
R1422 B.n626 B.n243 10.6151
R1423 B.n638 B.n243 10.6151
R1424 B.n639 B.n638 10.6151
R1425 B.n640 B.n639 10.6151
R1426 B.n641 B.n640 10.6151
R1427 B.n642 B.n641 10.6151
R1428 B.n645 B.n642 10.6151
R1429 B.n646 B.n645 10.6151
R1430 B.n647 B.n646 10.6151
R1431 B.n648 B.n647 10.6151
R1432 B.n650 B.n648 10.6151
R1433 B.n651 B.n650 10.6151
R1434 B.n652 B.n651 10.6151
R1435 B.n653 B.n652 10.6151
R1436 B.n655 B.n653 10.6151
R1437 B.n656 B.n655 10.6151
R1438 B.n657 B.n656 10.6151
R1439 B.n658 B.n657 10.6151
R1440 B.n660 B.n658 10.6151
R1441 B.n661 B.n660 10.6151
R1442 B.n662 B.n661 10.6151
R1443 B.n663 B.n662 10.6151
R1444 B.n665 B.n663 10.6151
R1445 B.n666 B.n665 10.6151
R1446 B.n667 B.n666 10.6151
R1447 B.n668 B.n667 10.6151
R1448 B.n670 B.n668 10.6151
R1449 B.n671 B.n670 10.6151
R1450 B.n672 B.n671 10.6151
R1451 B.n673 B.n672 10.6151
R1452 B.n675 B.n673 10.6151
R1453 B.n676 B.n675 10.6151
R1454 B.n677 B.n676 10.6151
R1455 B.n678 B.n677 10.6151
R1456 B.n680 B.n678 10.6151
R1457 B.n681 B.n680 10.6151
R1458 B.n682 B.n681 10.6151
R1459 B.n683 B.n682 10.6151
R1460 B.n685 B.n683 10.6151
R1461 B.n686 B.n685 10.6151
R1462 B.n687 B.n686 10.6151
R1463 B.n688 B.n687 10.6151
R1464 B.n690 B.n688 10.6151
R1465 B.n691 B.n690 10.6151
R1466 B.n692 B.n691 10.6151
R1467 B.n693 B.n692 10.6151
R1468 B.n695 B.n693 10.6151
R1469 B.n696 B.n695 10.6151
R1470 B.n697 B.n696 10.6151
R1471 B.n698 B.n697 10.6151
R1472 B.n700 B.n698 10.6151
R1473 B.n701 B.n700 10.6151
R1474 B.n702 B.n701 10.6151
R1475 B.n799 B.n1 10.6151
R1476 B.n799 B.n798 10.6151
R1477 B.n798 B.n797 10.6151
R1478 B.n797 B.n10 10.6151
R1479 B.n791 B.n10 10.6151
R1480 B.n791 B.n790 10.6151
R1481 B.n790 B.n789 10.6151
R1482 B.n789 B.n18 10.6151
R1483 B.n783 B.n18 10.6151
R1484 B.n783 B.n782 10.6151
R1485 B.n782 B.n781 10.6151
R1486 B.n781 B.n25 10.6151
R1487 B.n775 B.n25 10.6151
R1488 B.n775 B.n774 10.6151
R1489 B.n774 B.n773 10.6151
R1490 B.n773 B.n32 10.6151
R1491 B.n767 B.n32 10.6151
R1492 B.n767 B.n766 10.6151
R1493 B.n766 B.n765 10.6151
R1494 B.n765 B.n38 10.6151
R1495 B.n759 B.n38 10.6151
R1496 B.n759 B.n758 10.6151
R1497 B.n758 B.n757 10.6151
R1498 B.n757 B.n46 10.6151
R1499 B.n751 B.n46 10.6151
R1500 B.n751 B.n750 10.6151
R1501 B.n750 B.n749 10.6151
R1502 B.n749 B.n53 10.6151
R1503 B.n743 B.n53 10.6151
R1504 B.n743 B.n742 10.6151
R1505 B.n742 B.n741 10.6151
R1506 B.n741 B.n60 10.6151
R1507 B.n735 B.n60 10.6151
R1508 B.n735 B.n734 10.6151
R1509 B.n734 B.n733 10.6151
R1510 B.n733 B.n67 10.6151
R1511 B.n727 B.n67 10.6151
R1512 B.n727 B.n726 10.6151
R1513 B.n726 B.n725 10.6151
R1514 B.n725 B.n74 10.6151
R1515 B.n719 B.n74 10.6151
R1516 B.n719 B.n718 10.6151
R1517 B.n718 B.n717 10.6151
R1518 B.n717 B.n80 10.6151
R1519 B.n711 B.n80 10.6151
R1520 B.n711 B.n710 10.6151
R1521 B.n710 B.n709 10.6151
R1522 B.n709 B.n88 10.6151
R1523 B.n129 B.n128 10.6151
R1524 B.n132 B.n129 10.6151
R1525 B.n133 B.n132 10.6151
R1526 B.n136 B.n133 10.6151
R1527 B.n137 B.n136 10.6151
R1528 B.n140 B.n137 10.6151
R1529 B.n141 B.n140 10.6151
R1530 B.n144 B.n141 10.6151
R1531 B.n145 B.n144 10.6151
R1532 B.n148 B.n145 10.6151
R1533 B.n149 B.n148 10.6151
R1534 B.n152 B.n149 10.6151
R1535 B.n153 B.n152 10.6151
R1536 B.n156 B.n153 10.6151
R1537 B.n157 B.n156 10.6151
R1538 B.n160 B.n157 10.6151
R1539 B.n161 B.n160 10.6151
R1540 B.n164 B.n161 10.6151
R1541 B.n165 B.n164 10.6151
R1542 B.n168 B.n165 10.6151
R1543 B.n169 B.n168 10.6151
R1544 B.n172 B.n169 10.6151
R1545 B.n173 B.n172 10.6151
R1546 B.n176 B.n173 10.6151
R1547 B.n181 B.n178 10.6151
R1548 B.n182 B.n181 10.6151
R1549 B.n185 B.n182 10.6151
R1550 B.n186 B.n185 10.6151
R1551 B.n189 B.n186 10.6151
R1552 B.n190 B.n189 10.6151
R1553 B.n193 B.n190 10.6151
R1554 B.n194 B.n193 10.6151
R1555 B.n198 B.n197 10.6151
R1556 B.n201 B.n198 10.6151
R1557 B.n202 B.n201 10.6151
R1558 B.n205 B.n202 10.6151
R1559 B.n206 B.n205 10.6151
R1560 B.n209 B.n206 10.6151
R1561 B.n210 B.n209 10.6151
R1562 B.n213 B.n210 10.6151
R1563 B.n214 B.n213 10.6151
R1564 B.n217 B.n214 10.6151
R1565 B.n218 B.n217 10.6151
R1566 B.n221 B.n218 10.6151
R1567 B.n222 B.n221 10.6151
R1568 B.n225 B.n222 10.6151
R1569 B.n226 B.n225 10.6151
R1570 B.n229 B.n226 10.6151
R1571 B.n230 B.n229 10.6151
R1572 B.n233 B.n230 10.6151
R1573 B.n234 B.n233 10.6151
R1574 B.n237 B.n234 10.6151
R1575 B.n238 B.n237 10.6151
R1576 B.n241 B.n238 10.6151
R1577 B.n242 B.n241 10.6151
R1578 B.n703 B.n242 10.6151
R1579 B.n807 B.n0 8.11757
R1580 B.n807 B.n1 8.11757
R1581 B.n436 B.n370 6.5566
R1582 B.n420 B.n419 6.5566
R1583 B.n178 B.n177 6.5566
R1584 B.n194 B.n124 6.5566
R1585 B.n439 B.n370 4.05904
R1586 B.n419 B.n418 4.05904
R1587 B.n177 B.n176 4.05904
R1588 B.n197 B.n124 4.05904
R1589 VN.n65 VN.n34 161.3
R1590 VN.n64 VN.n63 161.3
R1591 VN.n62 VN.n35 161.3
R1592 VN.n61 VN.n60 161.3
R1593 VN.n58 VN.n36 161.3
R1594 VN.n57 VN.n56 161.3
R1595 VN.n55 VN.n37 161.3
R1596 VN.n54 VN.n53 161.3
R1597 VN.n52 VN.n38 161.3
R1598 VN.n50 VN.n49 161.3
R1599 VN.n48 VN.n39 161.3
R1600 VN.n47 VN.n46 161.3
R1601 VN.n45 VN.n40 161.3
R1602 VN.n44 VN.n43 161.3
R1603 VN.n31 VN.n0 161.3
R1604 VN.n30 VN.n29 161.3
R1605 VN.n28 VN.n1 161.3
R1606 VN.n27 VN.n26 161.3
R1607 VN.n24 VN.n2 161.3
R1608 VN.n23 VN.n22 161.3
R1609 VN.n21 VN.n3 161.3
R1610 VN.n20 VN.n19 161.3
R1611 VN.n18 VN.n4 161.3
R1612 VN.n16 VN.n15 161.3
R1613 VN.n14 VN.n5 161.3
R1614 VN.n13 VN.n12 161.3
R1615 VN.n11 VN.n6 161.3
R1616 VN.n10 VN.n9 161.3
R1617 VN.n8 VN.t7 106.01
R1618 VN.n42 VN.t6 106.01
R1619 VN.n33 VN.n32 88.7361
R1620 VN.n67 VN.n66 88.7361
R1621 VN.n7 VN.t1 75.2832
R1622 VN.n17 VN.t0 75.2832
R1623 VN.n25 VN.t4 75.2832
R1624 VN.n32 VN.t5 75.2832
R1625 VN.n41 VN.t8 75.2832
R1626 VN.n51 VN.t9 75.2832
R1627 VN.n59 VN.t2 75.2832
R1628 VN.n66 VN.t3 75.2832
R1629 VN.n8 VN.n7 65.1987
R1630 VN.n42 VN.n41 65.1987
R1631 VN.n30 VN.n1 56.5193
R1632 VN.n64 VN.n35 56.5193
R1633 VN.n12 VN.n5 47.7779
R1634 VN.n19 VN.n3 47.7779
R1635 VN.n46 VN.n39 47.7779
R1636 VN.n53 VN.n37 47.7779
R1637 VN VN.n67 45.9944
R1638 VN.n12 VN.n11 33.2089
R1639 VN.n23 VN.n3 33.2089
R1640 VN.n46 VN.n45 33.2089
R1641 VN.n57 VN.n37 33.2089
R1642 VN.n11 VN.n10 24.4675
R1643 VN.n16 VN.n5 24.4675
R1644 VN.n19 VN.n18 24.4675
R1645 VN.n24 VN.n23 24.4675
R1646 VN.n26 VN.n1 24.4675
R1647 VN.n31 VN.n30 24.4675
R1648 VN.n45 VN.n44 24.4675
R1649 VN.n53 VN.n52 24.4675
R1650 VN.n50 VN.n39 24.4675
R1651 VN.n60 VN.n35 24.4675
R1652 VN.n58 VN.n57 24.4675
R1653 VN.n65 VN.n64 24.4675
R1654 VN.n32 VN.n31 22.0208
R1655 VN.n66 VN.n65 22.0208
R1656 VN.n26 VN.n25 19.5741
R1657 VN.n60 VN.n59 19.5741
R1658 VN.n43 VN.n42 13.0188
R1659 VN.n9 VN.n8 13.0188
R1660 VN.n17 VN.n16 12.234
R1661 VN.n18 VN.n17 12.234
R1662 VN.n52 VN.n51 12.234
R1663 VN.n51 VN.n50 12.234
R1664 VN.n10 VN.n7 4.8939
R1665 VN.n25 VN.n24 4.8939
R1666 VN.n44 VN.n41 4.8939
R1667 VN.n59 VN.n58 4.8939
R1668 VN.n67 VN.n34 0.278367
R1669 VN.n33 VN.n0 0.278367
R1670 VN.n63 VN.n34 0.189894
R1671 VN.n63 VN.n62 0.189894
R1672 VN.n62 VN.n61 0.189894
R1673 VN.n61 VN.n36 0.189894
R1674 VN.n56 VN.n36 0.189894
R1675 VN.n56 VN.n55 0.189894
R1676 VN.n55 VN.n54 0.189894
R1677 VN.n54 VN.n38 0.189894
R1678 VN.n49 VN.n38 0.189894
R1679 VN.n49 VN.n48 0.189894
R1680 VN.n48 VN.n47 0.189894
R1681 VN.n47 VN.n40 0.189894
R1682 VN.n43 VN.n40 0.189894
R1683 VN.n9 VN.n6 0.189894
R1684 VN.n13 VN.n6 0.189894
R1685 VN.n14 VN.n13 0.189894
R1686 VN.n15 VN.n14 0.189894
R1687 VN.n15 VN.n4 0.189894
R1688 VN.n20 VN.n4 0.189894
R1689 VN.n21 VN.n20 0.189894
R1690 VN.n22 VN.n21 0.189894
R1691 VN.n22 VN.n2 0.189894
R1692 VN.n27 VN.n2 0.189894
R1693 VN.n28 VN.n27 0.189894
R1694 VN.n29 VN.n28 0.189894
R1695 VN.n29 VN.n0 0.189894
R1696 VN VN.n33 0.153454
R1697 VDD2.n1 VDD2.t2 70.7899
R1698 VDD2.n4 VDD2.t6 68.7642
R1699 VDD2.n3 VDD2.n2 67.0902
R1700 VDD2 VDD2.n7 67.0874
R1701 VDD2.n6 VDD2.n5 65.6264
R1702 VDD2.n1 VDD2.n0 65.6261
R1703 VDD2.n4 VDD2.n3 38.7778
R1704 VDD2.n7 VDD2.t1 3.13838
R1705 VDD2.n7 VDD2.t3 3.13838
R1706 VDD2.n5 VDD2.t7 3.13838
R1707 VDD2.n5 VDD2.t0 3.13838
R1708 VDD2.n2 VDD2.t5 3.13838
R1709 VDD2.n2 VDD2.t4 3.13838
R1710 VDD2.n0 VDD2.t8 3.13838
R1711 VDD2.n0 VDD2.t9 3.13838
R1712 VDD2.n6 VDD2.n4 2.02636
R1713 VDD2 VDD2.n6 0.565155
R1714 VDD2.n3 VDD2.n1 0.451619
C0 VN VP 6.4896f
C1 VTAIL VP 6.3534f
C2 VDD1 VP 5.89231f
C3 VTAIL VN 6.33917f
C4 VDD1 VN 0.152015f
C5 VDD2 VP 0.509064f
C6 VDD1 VTAIL 7.448669f
C7 VDD2 VN 5.53797f
C8 VDD2 VTAIL 7.49665f
C9 VDD2 VDD1 1.79611f
C10 VDD2 B 5.496676f
C11 VDD1 B 5.482637f
C12 VTAIL B 5.166324f
C13 VN B 14.76934f
C14 VP B 13.310868f
C15 VDD2.t2 B 1.20531f
C16 VDD2.t8 B 0.1121f
C17 VDD2.t9 B 0.1121f
C18 VDD2.n0 B 0.940125f
C19 VDD2.n1 B 0.744386f
C20 VDD2.t5 B 0.1121f
C21 VDD2.t4 B 0.1121f
C22 VDD2.n2 B 0.949856f
C23 VDD2.n3 B 2.02878f
C24 VDD2.t6 B 1.19412f
C25 VDD2.n4 B 2.19686f
C26 VDD2.t7 B 0.1121f
C27 VDD2.t0 B 0.1121f
C28 VDD2.n5 B 0.940128f
C29 VDD2.n6 B 0.371379f
C30 VDD2.t1 B 0.1121f
C31 VDD2.t3 B 0.1121f
C32 VDD2.n7 B 0.949824f
C33 VN.n0 B 0.035754f
C34 VN.t5 B 0.917533f
C35 VN.n1 B 0.04148f
C36 VN.n2 B 0.027119f
C37 VN.t4 B 0.917533f
C38 VN.n3 B 0.023949f
C39 VN.n4 B 0.027119f
C40 VN.t0 B 0.917533f
C41 VN.n5 B 0.05103f
C42 VN.n6 B 0.027119f
C43 VN.t1 B 0.917533f
C44 VN.n7 B 0.40631f
C45 VN.t7 B 1.05775f
C46 VN.n8 B 0.414964f
C47 VN.n9 B 0.203448f
C48 VN.n10 B 0.03058f
C49 VN.n11 B 0.054746f
C50 VN.n12 B 0.023949f
C51 VN.n13 B 0.027119f
C52 VN.n14 B 0.027119f
C53 VN.n15 B 0.027119f
C54 VN.n16 B 0.038066f
C55 VN.n17 B 0.347855f
C56 VN.n18 B 0.038066f
C57 VN.n19 B 0.05103f
C58 VN.n20 B 0.027119f
C59 VN.n21 B 0.027119f
C60 VN.n22 B 0.027119f
C61 VN.n23 B 0.054746f
C62 VN.n24 B 0.03058f
C63 VN.n25 B 0.347855f
C64 VN.n26 B 0.045552f
C65 VN.n27 B 0.027119f
C66 VN.n28 B 0.027119f
C67 VN.n29 B 0.027119f
C68 VN.n30 B 0.037702f
C69 VN.n31 B 0.048047f
C70 VN.n32 B 0.43554f
C71 VN.n33 B 0.031145f
C72 VN.n34 B 0.035754f
C73 VN.t3 B 0.917533f
C74 VN.n35 B 0.04148f
C75 VN.n36 B 0.027119f
C76 VN.t2 B 0.917533f
C77 VN.n37 B 0.023949f
C78 VN.n38 B 0.027119f
C79 VN.t9 B 0.917533f
C80 VN.n39 B 0.05103f
C81 VN.n40 B 0.027119f
C82 VN.t8 B 0.917533f
C83 VN.n41 B 0.40631f
C84 VN.t6 B 1.05775f
C85 VN.n42 B 0.414964f
C86 VN.n43 B 0.203448f
C87 VN.n44 B 0.03058f
C88 VN.n45 B 0.054746f
C89 VN.n46 B 0.023949f
C90 VN.n47 B 0.027119f
C91 VN.n48 B 0.027119f
C92 VN.n49 B 0.027119f
C93 VN.n50 B 0.038066f
C94 VN.n51 B 0.347855f
C95 VN.n52 B 0.038066f
C96 VN.n53 B 0.05103f
C97 VN.n54 B 0.027119f
C98 VN.n55 B 0.027119f
C99 VN.n56 B 0.027119f
C100 VN.n57 B 0.054746f
C101 VN.n58 B 0.03058f
C102 VN.n59 B 0.347855f
C103 VN.n60 B 0.045552f
C104 VN.n61 B 0.027119f
C105 VN.n62 B 0.027119f
C106 VN.n63 B 0.027119f
C107 VN.n64 B 0.037702f
C108 VN.n65 B 0.048047f
C109 VN.n66 B 0.43554f
C110 VN.n67 B 1.32052f
C111 VDD1.t9 B 1.22531f
C112 VDD1.t5 B 0.113959f
C113 VDD1.t6 B 0.113959f
C114 VDD1.n0 B 0.955719f
C115 VDD1.n1 B 0.763909f
C116 VDD1.t0 B 1.2253f
C117 VDD1.t3 B 0.113959f
C118 VDD1.t7 B 0.113959f
C119 VDD1.n2 B 0.955715f
C120 VDD1.n3 B 0.756731f
C121 VDD1.t4 B 0.113959f
C122 VDD1.t8 B 0.113959f
C123 VDD1.n4 B 0.965608f
C124 VDD1.n5 B 2.159f
C125 VDD1.t2 B 0.113959f
C126 VDD1.t1 B 0.113959f
C127 VDD1.n6 B 0.955714f
C128 VDD1.n7 B 2.27614f
C129 VTAIL.t3 B 0.136949f
C130 VTAIL.t8 B 0.136949f
C131 VTAIL.n0 B 1.07382f
C132 VTAIL.n1 B 0.532658f
C133 VTAIL.t18 B 1.36838f
C134 VTAIL.n2 B 0.651275f
C135 VTAIL.t17 B 0.136949f
C136 VTAIL.t13 B 0.136949f
C137 VTAIL.n3 B 1.07382f
C138 VTAIL.n4 B 0.620392f
C139 VTAIL.t14 B 0.136949f
C140 VTAIL.t11 B 0.136949f
C141 VTAIL.n5 B 1.07382f
C142 VTAIL.n6 B 1.65415f
C143 VTAIL.t7 B 0.136949f
C144 VTAIL.t6 B 0.136949f
C145 VTAIL.n7 B 1.07383f
C146 VTAIL.n8 B 1.65415f
C147 VTAIL.t1 B 0.136949f
C148 VTAIL.t0 B 0.136949f
C149 VTAIL.n9 B 1.07383f
C150 VTAIL.n10 B 0.620386f
C151 VTAIL.t5 B 1.36839f
C152 VTAIL.n11 B 0.651266f
C153 VTAIL.t15 B 0.136949f
C154 VTAIL.t10 B 0.136949f
C155 VTAIL.n12 B 1.07383f
C156 VTAIL.n13 B 0.572323f
C157 VTAIL.t12 B 0.136949f
C158 VTAIL.t16 B 0.136949f
C159 VTAIL.n14 B 1.07383f
C160 VTAIL.n15 B 0.620386f
C161 VTAIL.t19 B 1.36838f
C162 VTAIL.n16 B 1.55381f
C163 VTAIL.t9 B 1.36838f
C164 VTAIL.n17 B 1.55381f
C165 VTAIL.t2 B 0.136949f
C166 VTAIL.t4 B 0.136949f
C167 VTAIL.n18 B 1.07382f
C168 VTAIL.n19 B 0.48078f
C169 VP.n0 B 0.036807f
C170 VP.t1 B 0.94457f
C171 VP.n1 B 0.042703f
C172 VP.n2 B 0.027918f
C173 VP.t5 B 0.94457f
C174 VP.n3 B 0.024654f
C175 VP.n4 B 0.027918f
C176 VP.t2 B 0.94457f
C177 VP.n5 B 0.052533f
C178 VP.n6 B 0.027918f
C179 VP.t6 B 0.94457f
C180 VP.n7 B 0.358105f
C181 VP.n8 B 0.027918f
C182 VP.n9 B 0.049463f
C183 VP.n10 B 0.036807f
C184 VP.t8 B 0.94457f
C185 VP.n11 B 0.042703f
C186 VP.n12 B 0.027918f
C187 VP.t7 B 0.94457f
C188 VP.n13 B 0.024654f
C189 VP.n14 B 0.027918f
C190 VP.t3 B 0.94457f
C191 VP.n15 B 0.052533f
C192 VP.n16 B 0.027918f
C193 VP.t4 B 0.94457f
C194 VP.n17 B 0.418282f
C195 VP.t0 B 1.08891f
C196 VP.n18 B 0.427192f
C197 VP.n19 B 0.209443f
C198 VP.n20 B 0.031481f
C199 VP.n21 B 0.05636f
C200 VP.n22 B 0.024654f
C201 VP.n23 B 0.027918f
C202 VP.n24 B 0.027918f
C203 VP.n25 B 0.027918f
C204 VP.n26 B 0.039188f
C205 VP.n27 B 0.358105f
C206 VP.n28 B 0.039188f
C207 VP.n29 B 0.052533f
C208 VP.n30 B 0.027918f
C209 VP.n31 B 0.027918f
C210 VP.n32 B 0.027918f
C211 VP.n33 B 0.05636f
C212 VP.n34 B 0.031481f
C213 VP.n35 B 0.358105f
C214 VP.n36 B 0.046894f
C215 VP.n37 B 0.027918f
C216 VP.n38 B 0.027918f
C217 VP.n39 B 0.027918f
C218 VP.n40 B 0.038813f
C219 VP.n41 B 0.049463f
C220 VP.n42 B 0.448374f
C221 VP.n43 B 1.3442f
C222 VP.t9 B 0.94457f
C223 VP.n44 B 0.448374f
C224 VP.n45 B 1.36616f
C225 VP.n46 B 0.036807f
C226 VP.n47 B 0.027918f
C227 VP.n48 B 0.038813f
C228 VP.n49 B 0.042703f
C229 VP.n50 B 0.046894f
C230 VP.n51 B 0.027918f
C231 VP.n52 B 0.027918f
C232 VP.n53 B 0.031481f
C233 VP.n54 B 0.05636f
C234 VP.n55 B 0.024654f
C235 VP.n56 B 0.027918f
C236 VP.n57 B 0.027918f
C237 VP.n58 B 0.027918f
C238 VP.n59 B 0.039188f
C239 VP.n60 B 0.358105f
C240 VP.n61 B 0.039188f
C241 VP.n62 B 0.052533f
C242 VP.n63 B 0.027918f
C243 VP.n64 B 0.027918f
C244 VP.n65 B 0.027918f
C245 VP.n66 B 0.05636f
C246 VP.n67 B 0.031481f
C247 VP.n68 B 0.358105f
C248 VP.n69 B 0.046894f
C249 VP.n70 B 0.027918f
C250 VP.n71 B 0.027918f
C251 VP.n72 B 0.027918f
C252 VP.n73 B 0.038813f
C253 VP.n74 B 0.049463f
C254 VP.n75 B 0.448374f
C255 VP.n76 B 0.032063f
.ends

