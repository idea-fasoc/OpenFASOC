* NGSPICE file created from diff_pair_sample_1301.ext - technology: sky130A

.subckt diff_pair_sample_1301 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=3.7401 ps=19.96 w=9.59 l=0.29
X1 VDD2.t8 VN.t1 VTAIL.t9 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X2 VDD1.t9 VP.t0 VTAIL.t7 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=3.7401 ps=19.96 w=9.59 l=0.29
X3 VDD2.t7 VN.t2 VTAIL.t14 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=1.58235 ps=9.92 w=9.59 l=0.29
X4 VTAIL.t12 VN.t3 VDD2.t6 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X5 VTAIL.t18 VP.t1 VDD1.t8 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X6 VTAIL.t17 VN.t4 VDD2.t5 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X7 VDD2.t4 VN.t5 VTAIL.t16 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=1.58235 ps=9.92 w=9.59 l=0.29
X8 VDD2.t3 VN.t6 VTAIL.t15 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=3.7401 ps=19.96 w=9.59 l=0.29
X9 VTAIL.t0 VP.t2 VDD1.t7 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X10 VDD1.t6 VP.t3 VTAIL.t19 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X11 VDD1.t5 VP.t4 VTAIL.t3 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=1.58235 ps=9.92 w=9.59 l=0.29
X12 VTAIL.t2 VP.t5 VDD1.t4 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X13 B.t11 B.t9 B.t10 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=0 ps=0 w=9.59 l=0.29
X14 B.t8 B.t6 B.t7 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=0 ps=0 w=9.59 l=0.29
X15 B.t5 B.t3 B.t4 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=0 ps=0 w=9.59 l=0.29
X16 VTAIL.t13 VN.t7 VDD2.t2 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X17 VDD1.t3 VP.t6 VTAIL.t6 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=3.7401 ps=19.96 w=9.59 l=0.29
X18 VDD1.t2 VP.t7 VTAIL.t4 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=1.58235 ps=9.92 w=9.59 l=0.29
X19 B.t2 B.t0 B.t1 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=3.7401 pd=19.96 as=0 ps=0 w=9.59 l=0.29
X20 VTAIL.t11 VN.t8 VDD2.t1 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X21 VDD2.t0 VN.t9 VTAIL.t8 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X22 VDD1.t1 VP.t8 VTAIL.t5 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
X23 VTAIL.t1 VP.t9 VDD1.t0 w_n1714_n2886# sky130_fd_pr__pfet_01v8 ad=1.58235 pd=9.92 as=1.58235 ps=9.92 w=9.59 l=0.29
R0 VN.n9 VN.t0 940.883
R1 VN.n3 VN.t5 940.883
R2 VN.n20 VN.t2 940.883
R3 VN.n14 VN.t6 940.883
R4 VN.n6 VN.t9 905.828
R5 VN.n8 VN.t8 905.828
R6 VN.n2 VN.t7 905.828
R7 VN.n17 VN.t1 905.828
R8 VN.n19 VN.t4 905.828
R9 VN.n13 VN.t3 905.828
R10 VN.n15 VN.n14 161.489
R11 VN.n4 VN.n3 161.489
R12 VN.n10 VN.n9 161.3
R13 VN.n21 VN.n20 161.3
R14 VN.n18 VN.n11 161.3
R15 VN.n17 VN.n16 161.3
R16 VN.n15 VN.n12 161.3
R17 VN.n7 VN.n0 161.3
R18 VN.n6 VN.n5 161.3
R19 VN.n4 VN.n1 161.3
R20 VN.n6 VN.n1 73.0308
R21 VN.n7 VN.n6 73.0308
R22 VN.n18 VN.n17 73.0308
R23 VN.n17 VN.n12 73.0308
R24 VN.n3 VN.n2 55.5035
R25 VN.n9 VN.n8 55.5035
R26 VN.n20 VN.n19 55.5035
R27 VN.n14 VN.n13 55.5035
R28 VN VN.n21 39.1463
R29 VN.n2 VN.n1 17.5278
R30 VN.n8 VN.n7 17.5278
R31 VN.n19 VN.n18 17.5278
R32 VN.n13 VN.n12 17.5278
R33 VN.n21 VN.n11 0.189894
R34 VN.n16 VN.n11 0.189894
R35 VN.n16 VN.n15 0.189894
R36 VN.n5 VN.n4 0.189894
R37 VN.n5 VN.n0 0.189894
R38 VN.n10 VN.n0 0.189894
R39 VN VN.n10 0.0516364
R40 VTAIL.n11 VTAIL.t15 64.3371
R41 VTAIL.n17 VTAIL.t10 64.3369
R42 VTAIL.n2 VTAIL.t6 64.3369
R43 VTAIL.n16 VTAIL.t7 64.3369
R44 VTAIL.n15 VTAIL.n14 60.9477
R45 VTAIL.n13 VTAIL.n12 60.9477
R46 VTAIL.n10 VTAIL.n9 60.9477
R47 VTAIL.n8 VTAIL.n7 60.9477
R48 VTAIL.n19 VTAIL.n18 60.9474
R49 VTAIL.n1 VTAIL.n0 60.9474
R50 VTAIL.n4 VTAIL.n3 60.9474
R51 VTAIL.n6 VTAIL.n5 60.9474
R52 VTAIL.n8 VTAIL.n6 21.7031
R53 VTAIL.n17 VTAIL.n16 21.1686
R54 VTAIL.n18 VTAIL.t8 3.38997
R55 VTAIL.n18 VTAIL.t11 3.38997
R56 VTAIL.n0 VTAIL.t16 3.38997
R57 VTAIL.n0 VTAIL.t13 3.38997
R58 VTAIL.n3 VTAIL.t5 3.38997
R59 VTAIL.n3 VTAIL.t1 3.38997
R60 VTAIL.n5 VTAIL.t4 3.38997
R61 VTAIL.n5 VTAIL.t0 3.38997
R62 VTAIL.n14 VTAIL.t19 3.38997
R63 VTAIL.n14 VTAIL.t18 3.38997
R64 VTAIL.n12 VTAIL.t3 3.38997
R65 VTAIL.n12 VTAIL.t2 3.38997
R66 VTAIL.n9 VTAIL.t9 3.38997
R67 VTAIL.n9 VTAIL.t12 3.38997
R68 VTAIL.n7 VTAIL.t14 3.38997
R69 VTAIL.n7 VTAIL.t17 3.38997
R70 VTAIL.n13 VTAIL.n11 0.737569
R71 VTAIL.n2 VTAIL.n1 0.737569
R72 VTAIL.n10 VTAIL.n8 0.534983
R73 VTAIL.n11 VTAIL.n10 0.534983
R74 VTAIL.n15 VTAIL.n13 0.534983
R75 VTAIL.n16 VTAIL.n15 0.534983
R76 VTAIL.n6 VTAIL.n4 0.534983
R77 VTAIL.n4 VTAIL.n2 0.534983
R78 VTAIL.n19 VTAIL.n17 0.534983
R79 VTAIL VTAIL.n1 0.459552
R80 VTAIL VTAIL.n19 0.075931
R81 VDD2.n1 VDD2.t4 81.5502
R82 VDD2.n4 VDD2.t7 81.0159
R83 VDD2.n3 VDD2.n2 77.9717
R84 VDD2 VDD2.n7 77.9689
R85 VDD2.n6 VDD2.n5 77.6265
R86 VDD2.n1 VDD2.n0 77.6262
R87 VDD2.n4 VDD2.n3 34.5213
R88 VDD2.n7 VDD2.t6 3.38997
R89 VDD2.n7 VDD2.t3 3.38997
R90 VDD2.n5 VDD2.t5 3.38997
R91 VDD2.n5 VDD2.t8 3.38997
R92 VDD2.n2 VDD2.t1 3.38997
R93 VDD2.n2 VDD2.t9 3.38997
R94 VDD2.n0 VDD2.t2 3.38997
R95 VDD2.n0 VDD2.t0 3.38997
R96 VDD2.n6 VDD2.n4 0.534983
R97 VDD2 VDD2.n6 0.19231
R98 VDD2.n3 VDD2.n1 0.0787747
R99 VP.n21 VP.t6 940.883
R100 VP.n14 VP.t7 940.883
R101 VP.n5 VP.t4 940.883
R102 VP.n11 VP.t0 940.883
R103 VP.n18 VP.t8 905.828
R104 VP.n20 VP.t9 905.828
R105 VP.n13 VP.t2 905.828
R106 VP.n8 VP.t3 905.828
R107 VP.n4 VP.t5 905.828
R108 VP.n10 VP.t1 905.828
R109 VP.n6 VP.n5 161.489
R110 VP.n22 VP.n21 161.3
R111 VP.n6 VP.n3 161.3
R112 VP.n8 VP.n7 161.3
R113 VP.n9 VP.n2 161.3
R114 VP.n12 VP.n11 161.3
R115 VP.n19 VP.n0 161.3
R116 VP.n18 VP.n17 161.3
R117 VP.n16 VP.n1 161.3
R118 VP.n15 VP.n14 161.3
R119 VP.n18 VP.n1 73.0308
R120 VP.n19 VP.n18 73.0308
R121 VP.n8 VP.n3 73.0308
R122 VP.n9 VP.n8 73.0308
R123 VP.n14 VP.n13 55.5035
R124 VP.n21 VP.n20 55.5035
R125 VP.n5 VP.n4 55.5035
R126 VP.n11 VP.n10 55.5035
R127 VP.n15 VP.n12 38.7657
R128 VP.n13 VP.n1 17.5278
R129 VP.n20 VP.n19 17.5278
R130 VP.n4 VP.n3 17.5278
R131 VP.n10 VP.n9 17.5278
R132 VP.n7 VP.n6 0.189894
R133 VP.n7 VP.n2 0.189894
R134 VP.n12 VP.n2 0.189894
R135 VP.n16 VP.n15 0.189894
R136 VP.n17 VP.n16 0.189894
R137 VP.n17 VP.n0 0.189894
R138 VP.n22 VP.n0 0.189894
R139 VP VP.n22 0.0516364
R140 VDD1.n1 VDD1.t5 81.5503
R141 VDD1.n3 VDD1.t2 81.5502
R142 VDD1.n5 VDD1.n4 77.9717
R143 VDD1.n1 VDD1.n0 77.6265
R144 VDD1.n7 VDD1.n6 77.6263
R145 VDD1.n3 VDD1.n2 77.6262
R146 VDD1.n7 VDD1.n5 35.3716
R147 VDD1.n6 VDD1.t8 3.38997
R148 VDD1.n6 VDD1.t9 3.38997
R149 VDD1.n0 VDD1.t4 3.38997
R150 VDD1.n0 VDD1.t6 3.38997
R151 VDD1.n4 VDD1.t0 3.38997
R152 VDD1.n4 VDD1.t3 3.38997
R153 VDD1.n2 VDD1.t7 3.38997
R154 VDD1.n2 VDD1.t1 3.38997
R155 VDD1 VDD1.n7 0.343172
R156 VDD1 VDD1.n1 0.19231
R157 VDD1.n5 VDD1.n3 0.0787747
R158 B.n92 B.t6 1014.61
R159 B.n100 B.t3 1014.61
R160 B.n30 B.t0 1014.61
R161 B.n36 B.t9 1014.61
R162 B.n334 B.n333 585
R163 B.n335 B.n54 585
R164 B.n337 B.n336 585
R165 B.n338 B.n53 585
R166 B.n340 B.n339 585
R167 B.n341 B.n52 585
R168 B.n343 B.n342 585
R169 B.n344 B.n51 585
R170 B.n346 B.n345 585
R171 B.n347 B.n50 585
R172 B.n349 B.n348 585
R173 B.n350 B.n49 585
R174 B.n352 B.n351 585
R175 B.n353 B.n48 585
R176 B.n355 B.n354 585
R177 B.n356 B.n47 585
R178 B.n358 B.n357 585
R179 B.n359 B.n46 585
R180 B.n361 B.n360 585
R181 B.n362 B.n45 585
R182 B.n364 B.n363 585
R183 B.n365 B.n44 585
R184 B.n367 B.n366 585
R185 B.n368 B.n43 585
R186 B.n370 B.n369 585
R187 B.n371 B.n42 585
R188 B.n373 B.n372 585
R189 B.n374 B.n41 585
R190 B.n376 B.n375 585
R191 B.n377 B.n40 585
R192 B.n379 B.n378 585
R193 B.n380 B.n39 585
R194 B.n382 B.n381 585
R195 B.n383 B.n38 585
R196 B.n385 B.n384 585
R197 B.n387 B.n35 585
R198 B.n389 B.n388 585
R199 B.n390 B.n34 585
R200 B.n392 B.n391 585
R201 B.n393 B.n33 585
R202 B.n395 B.n394 585
R203 B.n396 B.n32 585
R204 B.n398 B.n397 585
R205 B.n399 B.n29 585
R206 B.n402 B.n401 585
R207 B.n403 B.n28 585
R208 B.n405 B.n404 585
R209 B.n406 B.n27 585
R210 B.n408 B.n407 585
R211 B.n409 B.n26 585
R212 B.n411 B.n410 585
R213 B.n412 B.n25 585
R214 B.n414 B.n413 585
R215 B.n415 B.n24 585
R216 B.n417 B.n416 585
R217 B.n418 B.n23 585
R218 B.n420 B.n419 585
R219 B.n421 B.n22 585
R220 B.n423 B.n422 585
R221 B.n424 B.n21 585
R222 B.n426 B.n425 585
R223 B.n427 B.n20 585
R224 B.n429 B.n428 585
R225 B.n430 B.n19 585
R226 B.n432 B.n431 585
R227 B.n433 B.n18 585
R228 B.n435 B.n434 585
R229 B.n436 B.n17 585
R230 B.n438 B.n437 585
R231 B.n439 B.n16 585
R232 B.n441 B.n440 585
R233 B.n442 B.n15 585
R234 B.n444 B.n443 585
R235 B.n445 B.n14 585
R236 B.n447 B.n446 585
R237 B.n448 B.n13 585
R238 B.n450 B.n449 585
R239 B.n451 B.n12 585
R240 B.n453 B.n452 585
R241 B.n332 B.n55 585
R242 B.n331 B.n330 585
R243 B.n329 B.n56 585
R244 B.n328 B.n327 585
R245 B.n326 B.n57 585
R246 B.n325 B.n324 585
R247 B.n323 B.n58 585
R248 B.n322 B.n321 585
R249 B.n320 B.n59 585
R250 B.n319 B.n318 585
R251 B.n317 B.n60 585
R252 B.n316 B.n315 585
R253 B.n314 B.n61 585
R254 B.n313 B.n312 585
R255 B.n311 B.n62 585
R256 B.n310 B.n309 585
R257 B.n308 B.n63 585
R258 B.n307 B.n306 585
R259 B.n305 B.n64 585
R260 B.n304 B.n303 585
R261 B.n302 B.n65 585
R262 B.n301 B.n300 585
R263 B.n299 B.n66 585
R264 B.n298 B.n297 585
R265 B.n296 B.n67 585
R266 B.n295 B.n294 585
R267 B.n293 B.n68 585
R268 B.n292 B.n291 585
R269 B.n290 B.n69 585
R270 B.n289 B.n288 585
R271 B.n287 B.n70 585
R272 B.n286 B.n285 585
R273 B.n284 B.n71 585
R274 B.n283 B.n282 585
R275 B.n281 B.n72 585
R276 B.n280 B.n279 585
R277 B.n278 B.n73 585
R278 B.n277 B.n276 585
R279 B.n275 B.n74 585
R280 B.n155 B.n118 585
R281 B.n157 B.n156 585
R282 B.n158 B.n117 585
R283 B.n160 B.n159 585
R284 B.n161 B.n116 585
R285 B.n163 B.n162 585
R286 B.n164 B.n115 585
R287 B.n166 B.n165 585
R288 B.n167 B.n114 585
R289 B.n169 B.n168 585
R290 B.n170 B.n113 585
R291 B.n172 B.n171 585
R292 B.n173 B.n112 585
R293 B.n175 B.n174 585
R294 B.n176 B.n111 585
R295 B.n178 B.n177 585
R296 B.n179 B.n110 585
R297 B.n181 B.n180 585
R298 B.n182 B.n109 585
R299 B.n184 B.n183 585
R300 B.n185 B.n108 585
R301 B.n187 B.n186 585
R302 B.n188 B.n107 585
R303 B.n190 B.n189 585
R304 B.n191 B.n106 585
R305 B.n193 B.n192 585
R306 B.n194 B.n105 585
R307 B.n196 B.n195 585
R308 B.n197 B.n104 585
R309 B.n199 B.n198 585
R310 B.n200 B.n103 585
R311 B.n202 B.n201 585
R312 B.n203 B.n102 585
R313 B.n205 B.n204 585
R314 B.n206 B.n99 585
R315 B.n209 B.n208 585
R316 B.n210 B.n98 585
R317 B.n212 B.n211 585
R318 B.n213 B.n97 585
R319 B.n215 B.n214 585
R320 B.n216 B.n96 585
R321 B.n218 B.n217 585
R322 B.n219 B.n95 585
R323 B.n221 B.n220 585
R324 B.n223 B.n222 585
R325 B.n224 B.n91 585
R326 B.n226 B.n225 585
R327 B.n227 B.n90 585
R328 B.n229 B.n228 585
R329 B.n230 B.n89 585
R330 B.n232 B.n231 585
R331 B.n233 B.n88 585
R332 B.n235 B.n234 585
R333 B.n236 B.n87 585
R334 B.n238 B.n237 585
R335 B.n239 B.n86 585
R336 B.n241 B.n240 585
R337 B.n242 B.n85 585
R338 B.n244 B.n243 585
R339 B.n245 B.n84 585
R340 B.n247 B.n246 585
R341 B.n248 B.n83 585
R342 B.n250 B.n249 585
R343 B.n251 B.n82 585
R344 B.n253 B.n252 585
R345 B.n254 B.n81 585
R346 B.n256 B.n255 585
R347 B.n257 B.n80 585
R348 B.n259 B.n258 585
R349 B.n260 B.n79 585
R350 B.n262 B.n261 585
R351 B.n263 B.n78 585
R352 B.n265 B.n264 585
R353 B.n266 B.n77 585
R354 B.n268 B.n267 585
R355 B.n269 B.n76 585
R356 B.n271 B.n270 585
R357 B.n272 B.n75 585
R358 B.n274 B.n273 585
R359 B.n154 B.n153 585
R360 B.n152 B.n119 585
R361 B.n151 B.n150 585
R362 B.n149 B.n120 585
R363 B.n148 B.n147 585
R364 B.n146 B.n121 585
R365 B.n145 B.n144 585
R366 B.n143 B.n122 585
R367 B.n142 B.n141 585
R368 B.n140 B.n123 585
R369 B.n139 B.n138 585
R370 B.n137 B.n124 585
R371 B.n136 B.n135 585
R372 B.n134 B.n125 585
R373 B.n133 B.n132 585
R374 B.n131 B.n126 585
R375 B.n130 B.n129 585
R376 B.n128 B.n127 585
R377 B.n2 B.n0 585
R378 B.n481 B.n1 585
R379 B.n480 B.n479 585
R380 B.n478 B.n3 585
R381 B.n477 B.n476 585
R382 B.n475 B.n4 585
R383 B.n474 B.n473 585
R384 B.n472 B.n5 585
R385 B.n471 B.n470 585
R386 B.n469 B.n6 585
R387 B.n468 B.n467 585
R388 B.n466 B.n7 585
R389 B.n465 B.n464 585
R390 B.n463 B.n8 585
R391 B.n462 B.n461 585
R392 B.n460 B.n9 585
R393 B.n459 B.n458 585
R394 B.n457 B.n10 585
R395 B.n456 B.n455 585
R396 B.n454 B.n11 585
R397 B.n483 B.n482 585
R398 B.n155 B.n154 478.086
R399 B.n452 B.n11 478.086
R400 B.n275 B.n274 478.086
R401 B.n334 B.n55 478.086
R402 B.n154 B.n119 163.367
R403 B.n150 B.n119 163.367
R404 B.n150 B.n149 163.367
R405 B.n149 B.n148 163.367
R406 B.n148 B.n121 163.367
R407 B.n144 B.n121 163.367
R408 B.n144 B.n143 163.367
R409 B.n143 B.n142 163.367
R410 B.n142 B.n123 163.367
R411 B.n138 B.n123 163.367
R412 B.n138 B.n137 163.367
R413 B.n137 B.n136 163.367
R414 B.n136 B.n125 163.367
R415 B.n132 B.n125 163.367
R416 B.n132 B.n131 163.367
R417 B.n131 B.n130 163.367
R418 B.n130 B.n127 163.367
R419 B.n127 B.n2 163.367
R420 B.n482 B.n2 163.367
R421 B.n482 B.n481 163.367
R422 B.n481 B.n480 163.367
R423 B.n480 B.n3 163.367
R424 B.n476 B.n3 163.367
R425 B.n476 B.n475 163.367
R426 B.n475 B.n474 163.367
R427 B.n474 B.n5 163.367
R428 B.n470 B.n5 163.367
R429 B.n470 B.n469 163.367
R430 B.n469 B.n468 163.367
R431 B.n468 B.n7 163.367
R432 B.n464 B.n7 163.367
R433 B.n464 B.n463 163.367
R434 B.n463 B.n462 163.367
R435 B.n462 B.n9 163.367
R436 B.n458 B.n9 163.367
R437 B.n458 B.n457 163.367
R438 B.n457 B.n456 163.367
R439 B.n456 B.n11 163.367
R440 B.n156 B.n155 163.367
R441 B.n156 B.n117 163.367
R442 B.n160 B.n117 163.367
R443 B.n161 B.n160 163.367
R444 B.n162 B.n161 163.367
R445 B.n162 B.n115 163.367
R446 B.n166 B.n115 163.367
R447 B.n167 B.n166 163.367
R448 B.n168 B.n167 163.367
R449 B.n168 B.n113 163.367
R450 B.n172 B.n113 163.367
R451 B.n173 B.n172 163.367
R452 B.n174 B.n173 163.367
R453 B.n174 B.n111 163.367
R454 B.n178 B.n111 163.367
R455 B.n179 B.n178 163.367
R456 B.n180 B.n179 163.367
R457 B.n180 B.n109 163.367
R458 B.n184 B.n109 163.367
R459 B.n185 B.n184 163.367
R460 B.n186 B.n185 163.367
R461 B.n186 B.n107 163.367
R462 B.n190 B.n107 163.367
R463 B.n191 B.n190 163.367
R464 B.n192 B.n191 163.367
R465 B.n192 B.n105 163.367
R466 B.n196 B.n105 163.367
R467 B.n197 B.n196 163.367
R468 B.n198 B.n197 163.367
R469 B.n198 B.n103 163.367
R470 B.n202 B.n103 163.367
R471 B.n203 B.n202 163.367
R472 B.n204 B.n203 163.367
R473 B.n204 B.n99 163.367
R474 B.n209 B.n99 163.367
R475 B.n210 B.n209 163.367
R476 B.n211 B.n210 163.367
R477 B.n211 B.n97 163.367
R478 B.n215 B.n97 163.367
R479 B.n216 B.n215 163.367
R480 B.n217 B.n216 163.367
R481 B.n217 B.n95 163.367
R482 B.n221 B.n95 163.367
R483 B.n222 B.n221 163.367
R484 B.n222 B.n91 163.367
R485 B.n226 B.n91 163.367
R486 B.n227 B.n226 163.367
R487 B.n228 B.n227 163.367
R488 B.n228 B.n89 163.367
R489 B.n232 B.n89 163.367
R490 B.n233 B.n232 163.367
R491 B.n234 B.n233 163.367
R492 B.n234 B.n87 163.367
R493 B.n238 B.n87 163.367
R494 B.n239 B.n238 163.367
R495 B.n240 B.n239 163.367
R496 B.n240 B.n85 163.367
R497 B.n244 B.n85 163.367
R498 B.n245 B.n244 163.367
R499 B.n246 B.n245 163.367
R500 B.n246 B.n83 163.367
R501 B.n250 B.n83 163.367
R502 B.n251 B.n250 163.367
R503 B.n252 B.n251 163.367
R504 B.n252 B.n81 163.367
R505 B.n256 B.n81 163.367
R506 B.n257 B.n256 163.367
R507 B.n258 B.n257 163.367
R508 B.n258 B.n79 163.367
R509 B.n262 B.n79 163.367
R510 B.n263 B.n262 163.367
R511 B.n264 B.n263 163.367
R512 B.n264 B.n77 163.367
R513 B.n268 B.n77 163.367
R514 B.n269 B.n268 163.367
R515 B.n270 B.n269 163.367
R516 B.n270 B.n75 163.367
R517 B.n274 B.n75 163.367
R518 B.n276 B.n275 163.367
R519 B.n276 B.n73 163.367
R520 B.n280 B.n73 163.367
R521 B.n281 B.n280 163.367
R522 B.n282 B.n281 163.367
R523 B.n282 B.n71 163.367
R524 B.n286 B.n71 163.367
R525 B.n287 B.n286 163.367
R526 B.n288 B.n287 163.367
R527 B.n288 B.n69 163.367
R528 B.n292 B.n69 163.367
R529 B.n293 B.n292 163.367
R530 B.n294 B.n293 163.367
R531 B.n294 B.n67 163.367
R532 B.n298 B.n67 163.367
R533 B.n299 B.n298 163.367
R534 B.n300 B.n299 163.367
R535 B.n300 B.n65 163.367
R536 B.n304 B.n65 163.367
R537 B.n305 B.n304 163.367
R538 B.n306 B.n305 163.367
R539 B.n306 B.n63 163.367
R540 B.n310 B.n63 163.367
R541 B.n311 B.n310 163.367
R542 B.n312 B.n311 163.367
R543 B.n312 B.n61 163.367
R544 B.n316 B.n61 163.367
R545 B.n317 B.n316 163.367
R546 B.n318 B.n317 163.367
R547 B.n318 B.n59 163.367
R548 B.n322 B.n59 163.367
R549 B.n323 B.n322 163.367
R550 B.n324 B.n323 163.367
R551 B.n324 B.n57 163.367
R552 B.n328 B.n57 163.367
R553 B.n329 B.n328 163.367
R554 B.n330 B.n329 163.367
R555 B.n330 B.n55 163.367
R556 B.n452 B.n451 163.367
R557 B.n451 B.n450 163.367
R558 B.n450 B.n13 163.367
R559 B.n446 B.n13 163.367
R560 B.n446 B.n445 163.367
R561 B.n445 B.n444 163.367
R562 B.n444 B.n15 163.367
R563 B.n440 B.n15 163.367
R564 B.n440 B.n439 163.367
R565 B.n439 B.n438 163.367
R566 B.n438 B.n17 163.367
R567 B.n434 B.n17 163.367
R568 B.n434 B.n433 163.367
R569 B.n433 B.n432 163.367
R570 B.n432 B.n19 163.367
R571 B.n428 B.n19 163.367
R572 B.n428 B.n427 163.367
R573 B.n427 B.n426 163.367
R574 B.n426 B.n21 163.367
R575 B.n422 B.n21 163.367
R576 B.n422 B.n421 163.367
R577 B.n421 B.n420 163.367
R578 B.n420 B.n23 163.367
R579 B.n416 B.n23 163.367
R580 B.n416 B.n415 163.367
R581 B.n415 B.n414 163.367
R582 B.n414 B.n25 163.367
R583 B.n410 B.n25 163.367
R584 B.n410 B.n409 163.367
R585 B.n409 B.n408 163.367
R586 B.n408 B.n27 163.367
R587 B.n404 B.n27 163.367
R588 B.n404 B.n403 163.367
R589 B.n403 B.n402 163.367
R590 B.n402 B.n29 163.367
R591 B.n397 B.n29 163.367
R592 B.n397 B.n396 163.367
R593 B.n396 B.n395 163.367
R594 B.n395 B.n33 163.367
R595 B.n391 B.n33 163.367
R596 B.n391 B.n390 163.367
R597 B.n390 B.n389 163.367
R598 B.n389 B.n35 163.367
R599 B.n384 B.n35 163.367
R600 B.n384 B.n383 163.367
R601 B.n383 B.n382 163.367
R602 B.n382 B.n39 163.367
R603 B.n378 B.n39 163.367
R604 B.n378 B.n377 163.367
R605 B.n377 B.n376 163.367
R606 B.n376 B.n41 163.367
R607 B.n372 B.n41 163.367
R608 B.n372 B.n371 163.367
R609 B.n371 B.n370 163.367
R610 B.n370 B.n43 163.367
R611 B.n366 B.n43 163.367
R612 B.n366 B.n365 163.367
R613 B.n365 B.n364 163.367
R614 B.n364 B.n45 163.367
R615 B.n360 B.n45 163.367
R616 B.n360 B.n359 163.367
R617 B.n359 B.n358 163.367
R618 B.n358 B.n47 163.367
R619 B.n354 B.n47 163.367
R620 B.n354 B.n353 163.367
R621 B.n353 B.n352 163.367
R622 B.n352 B.n49 163.367
R623 B.n348 B.n49 163.367
R624 B.n348 B.n347 163.367
R625 B.n347 B.n346 163.367
R626 B.n346 B.n51 163.367
R627 B.n342 B.n51 163.367
R628 B.n342 B.n341 163.367
R629 B.n341 B.n340 163.367
R630 B.n340 B.n53 163.367
R631 B.n336 B.n53 163.367
R632 B.n336 B.n335 163.367
R633 B.n335 B.n334 163.367
R634 B.n92 B.t8 121.21
R635 B.n36 B.t10 121.21
R636 B.n100 B.t5 121.2
R637 B.n30 B.t1 121.2
R638 B.n93 B.t7 109.186
R639 B.n37 B.t11 109.186
R640 B.n101 B.t4 109.175
R641 B.n31 B.t2 109.175
R642 B.n94 B.n93 59.5399
R643 B.n207 B.n101 59.5399
R644 B.n400 B.n31 59.5399
R645 B.n386 B.n37 59.5399
R646 B.n454 B.n453 31.0639
R647 B.n333 B.n332 31.0639
R648 B.n273 B.n74 31.0639
R649 B.n153 B.n118 31.0639
R650 B B.n483 18.0485
R651 B.n93 B.n92 12.0247
R652 B.n101 B.n100 12.0247
R653 B.n31 B.n30 12.0247
R654 B.n37 B.n36 12.0247
R655 B.n453 B.n12 10.6151
R656 B.n449 B.n12 10.6151
R657 B.n449 B.n448 10.6151
R658 B.n448 B.n447 10.6151
R659 B.n447 B.n14 10.6151
R660 B.n443 B.n14 10.6151
R661 B.n443 B.n442 10.6151
R662 B.n442 B.n441 10.6151
R663 B.n441 B.n16 10.6151
R664 B.n437 B.n16 10.6151
R665 B.n437 B.n436 10.6151
R666 B.n436 B.n435 10.6151
R667 B.n435 B.n18 10.6151
R668 B.n431 B.n18 10.6151
R669 B.n431 B.n430 10.6151
R670 B.n430 B.n429 10.6151
R671 B.n429 B.n20 10.6151
R672 B.n425 B.n20 10.6151
R673 B.n425 B.n424 10.6151
R674 B.n424 B.n423 10.6151
R675 B.n423 B.n22 10.6151
R676 B.n419 B.n22 10.6151
R677 B.n419 B.n418 10.6151
R678 B.n418 B.n417 10.6151
R679 B.n417 B.n24 10.6151
R680 B.n413 B.n24 10.6151
R681 B.n413 B.n412 10.6151
R682 B.n412 B.n411 10.6151
R683 B.n411 B.n26 10.6151
R684 B.n407 B.n26 10.6151
R685 B.n407 B.n406 10.6151
R686 B.n406 B.n405 10.6151
R687 B.n405 B.n28 10.6151
R688 B.n401 B.n28 10.6151
R689 B.n399 B.n398 10.6151
R690 B.n398 B.n32 10.6151
R691 B.n394 B.n32 10.6151
R692 B.n394 B.n393 10.6151
R693 B.n393 B.n392 10.6151
R694 B.n392 B.n34 10.6151
R695 B.n388 B.n34 10.6151
R696 B.n388 B.n387 10.6151
R697 B.n385 B.n38 10.6151
R698 B.n381 B.n38 10.6151
R699 B.n381 B.n380 10.6151
R700 B.n380 B.n379 10.6151
R701 B.n379 B.n40 10.6151
R702 B.n375 B.n40 10.6151
R703 B.n375 B.n374 10.6151
R704 B.n374 B.n373 10.6151
R705 B.n373 B.n42 10.6151
R706 B.n369 B.n42 10.6151
R707 B.n369 B.n368 10.6151
R708 B.n368 B.n367 10.6151
R709 B.n367 B.n44 10.6151
R710 B.n363 B.n44 10.6151
R711 B.n363 B.n362 10.6151
R712 B.n362 B.n361 10.6151
R713 B.n361 B.n46 10.6151
R714 B.n357 B.n46 10.6151
R715 B.n357 B.n356 10.6151
R716 B.n356 B.n355 10.6151
R717 B.n355 B.n48 10.6151
R718 B.n351 B.n48 10.6151
R719 B.n351 B.n350 10.6151
R720 B.n350 B.n349 10.6151
R721 B.n349 B.n50 10.6151
R722 B.n345 B.n50 10.6151
R723 B.n345 B.n344 10.6151
R724 B.n344 B.n343 10.6151
R725 B.n343 B.n52 10.6151
R726 B.n339 B.n52 10.6151
R727 B.n339 B.n338 10.6151
R728 B.n338 B.n337 10.6151
R729 B.n337 B.n54 10.6151
R730 B.n333 B.n54 10.6151
R731 B.n277 B.n74 10.6151
R732 B.n278 B.n277 10.6151
R733 B.n279 B.n278 10.6151
R734 B.n279 B.n72 10.6151
R735 B.n283 B.n72 10.6151
R736 B.n284 B.n283 10.6151
R737 B.n285 B.n284 10.6151
R738 B.n285 B.n70 10.6151
R739 B.n289 B.n70 10.6151
R740 B.n290 B.n289 10.6151
R741 B.n291 B.n290 10.6151
R742 B.n291 B.n68 10.6151
R743 B.n295 B.n68 10.6151
R744 B.n296 B.n295 10.6151
R745 B.n297 B.n296 10.6151
R746 B.n297 B.n66 10.6151
R747 B.n301 B.n66 10.6151
R748 B.n302 B.n301 10.6151
R749 B.n303 B.n302 10.6151
R750 B.n303 B.n64 10.6151
R751 B.n307 B.n64 10.6151
R752 B.n308 B.n307 10.6151
R753 B.n309 B.n308 10.6151
R754 B.n309 B.n62 10.6151
R755 B.n313 B.n62 10.6151
R756 B.n314 B.n313 10.6151
R757 B.n315 B.n314 10.6151
R758 B.n315 B.n60 10.6151
R759 B.n319 B.n60 10.6151
R760 B.n320 B.n319 10.6151
R761 B.n321 B.n320 10.6151
R762 B.n321 B.n58 10.6151
R763 B.n325 B.n58 10.6151
R764 B.n326 B.n325 10.6151
R765 B.n327 B.n326 10.6151
R766 B.n327 B.n56 10.6151
R767 B.n331 B.n56 10.6151
R768 B.n332 B.n331 10.6151
R769 B.n157 B.n118 10.6151
R770 B.n158 B.n157 10.6151
R771 B.n159 B.n158 10.6151
R772 B.n159 B.n116 10.6151
R773 B.n163 B.n116 10.6151
R774 B.n164 B.n163 10.6151
R775 B.n165 B.n164 10.6151
R776 B.n165 B.n114 10.6151
R777 B.n169 B.n114 10.6151
R778 B.n170 B.n169 10.6151
R779 B.n171 B.n170 10.6151
R780 B.n171 B.n112 10.6151
R781 B.n175 B.n112 10.6151
R782 B.n176 B.n175 10.6151
R783 B.n177 B.n176 10.6151
R784 B.n177 B.n110 10.6151
R785 B.n181 B.n110 10.6151
R786 B.n182 B.n181 10.6151
R787 B.n183 B.n182 10.6151
R788 B.n183 B.n108 10.6151
R789 B.n187 B.n108 10.6151
R790 B.n188 B.n187 10.6151
R791 B.n189 B.n188 10.6151
R792 B.n189 B.n106 10.6151
R793 B.n193 B.n106 10.6151
R794 B.n194 B.n193 10.6151
R795 B.n195 B.n194 10.6151
R796 B.n195 B.n104 10.6151
R797 B.n199 B.n104 10.6151
R798 B.n200 B.n199 10.6151
R799 B.n201 B.n200 10.6151
R800 B.n201 B.n102 10.6151
R801 B.n205 B.n102 10.6151
R802 B.n206 B.n205 10.6151
R803 B.n208 B.n98 10.6151
R804 B.n212 B.n98 10.6151
R805 B.n213 B.n212 10.6151
R806 B.n214 B.n213 10.6151
R807 B.n214 B.n96 10.6151
R808 B.n218 B.n96 10.6151
R809 B.n219 B.n218 10.6151
R810 B.n220 B.n219 10.6151
R811 B.n224 B.n223 10.6151
R812 B.n225 B.n224 10.6151
R813 B.n225 B.n90 10.6151
R814 B.n229 B.n90 10.6151
R815 B.n230 B.n229 10.6151
R816 B.n231 B.n230 10.6151
R817 B.n231 B.n88 10.6151
R818 B.n235 B.n88 10.6151
R819 B.n236 B.n235 10.6151
R820 B.n237 B.n236 10.6151
R821 B.n237 B.n86 10.6151
R822 B.n241 B.n86 10.6151
R823 B.n242 B.n241 10.6151
R824 B.n243 B.n242 10.6151
R825 B.n243 B.n84 10.6151
R826 B.n247 B.n84 10.6151
R827 B.n248 B.n247 10.6151
R828 B.n249 B.n248 10.6151
R829 B.n249 B.n82 10.6151
R830 B.n253 B.n82 10.6151
R831 B.n254 B.n253 10.6151
R832 B.n255 B.n254 10.6151
R833 B.n255 B.n80 10.6151
R834 B.n259 B.n80 10.6151
R835 B.n260 B.n259 10.6151
R836 B.n261 B.n260 10.6151
R837 B.n261 B.n78 10.6151
R838 B.n265 B.n78 10.6151
R839 B.n266 B.n265 10.6151
R840 B.n267 B.n266 10.6151
R841 B.n267 B.n76 10.6151
R842 B.n271 B.n76 10.6151
R843 B.n272 B.n271 10.6151
R844 B.n273 B.n272 10.6151
R845 B.n153 B.n152 10.6151
R846 B.n152 B.n151 10.6151
R847 B.n151 B.n120 10.6151
R848 B.n147 B.n120 10.6151
R849 B.n147 B.n146 10.6151
R850 B.n146 B.n145 10.6151
R851 B.n145 B.n122 10.6151
R852 B.n141 B.n122 10.6151
R853 B.n141 B.n140 10.6151
R854 B.n140 B.n139 10.6151
R855 B.n139 B.n124 10.6151
R856 B.n135 B.n124 10.6151
R857 B.n135 B.n134 10.6151
R858 B.n134 B.n133 10.6151
R859 B.n133 B.n126 10.6151
R860 B.n129 B.n126 10.6151
R861 B.n129 B.n128 10.6151
R862 B.n128 B.n0 10.6151
R863 B.n479 B.n1 10.6151
R864 B.n479 B.n478 10.6151
R865 B.n478 B.n477 10.6151
R866 B.n477 B.n4 10.6151
R867 B.n473 B.n4 10.6151
R868 B.n473 B.n472 10.6151
R869 B.n472 B.n471 10.6151
R870 B.n471 B.n6 10.6151
R871 B.n467 B.n6 10.6151
R872 B.n467 B.n466 10.6151
R873 B.n466 B.n465 10.6151
R874 B.n465 B.n8 10.6151
R875 B.n461 B.n8 10.6151
R876 B.n461 B.n460 10.6151
R877 B.n460 B.n459 10.6151
R878 B.n459 B.n10 10.6151
R879 B.n455 B.n10 10.6151
R880 B.n455 B.n454 10.6151
R881 B.n400 B.n399 6.5566
R882 B.n387 B.n386 6.5566
R883 B.n208 B.n207 6.5566
R884 B.n220 B.n94 6.5566
R885 B.n401 B.n400 4.05904
R886 B.n386 B.n385 4.05904
R887 B.n207 B.n206 4.05904
R888 B.n223 B.n94 4.05904
R889 B.n483 B.n0 2.81026
R890 B.n483 B.n1 2.81026
C0 VTAIL VP 2.90379f
C1 VDD1 VTAIL 17.3716f
C2 B VDD2 1.37986f
C3 VP VDD2 0.28902f
C4 VDD1 VDD2 0.718908f
C5 B w_n1714_n2886# 6.01092f
C6 VP w_n1714_n2886# 3.13591f
C7 VDD1 w_n1714_n2886# 1.66923f
C8 VTAIL VN 2.88916f
C9 VN VDD2 3.18731f
C10 B VP 1.0138f
C11 VDD1 B 1.35125f
C12 VN w_n1714_n2886# 2.91989f
C13 VDD1 VP 3.32411f
C14 VTAIL VDD2 17.4029f
C15 VTAIL w_n1714_n2886# 2.65068f
C16 VN B 0.663284f
C17 w_n1714_n2886# VDD2 1.69286f
C18 VN VP 4.54788f
C19 VDD1 VN 0.148026f
C20 VTAIL B 2.04543f
C21 VDD2 VSUBS 1.317988f
C22 VDD1 VSUBS 0.935623f
C23 VTAIL VSUBS 0.519385f
C24 VN VSUBS 4.37931f
C25 VP VSUBS 1.218303f
C26 B VSUBS 2.291425f
C27 w_n1714_n2886# VSUBS 61.148697f
C28 B.n0 VSUBS 0.005059f
C29 B.n1 VSUBS 0.005059f
C30 B.n2 VSUBS 0.008001f
C31 B.n3 VSUBS 0.008001f
C32 B.n4 VSUBS 0.008001f
C33 B.n5 VSUBS 0.008001f
C34 B.n6 VSUBS 0.008001f
C35 B.n7 VSUBS 0.008001f
C36 B.n8 VSUBS 0.008001f
C37 B.n9 VSUBS 0.008001f
C38 B.n10 VSUBS 0.008001f
C39 B.n11 VSUBS 0.017453f
C40 B.n12 VSUBS 0.008001f
C41 B.n13 VSUBS 0.008001f
C42 B.n14 VSUBS 0.008001f
C43 B.n15 VSUBS 0.008001f
C44 B.n16 VSUBS 0.008001f
C45 B.n17 VSUBS 0.008001f
C46 B.n18 VSUBS 0.008001f
C47 B.n19 VSUBS 0.008001f
C48 B.n20 VSUBS 0.008001f
C49 B.n21 VSUBS 0.008001f
C50 B.n22 VSUBS 0.008001f
C51 B.n23 VSUBS 0.008001f
C52 B.n24 VSUBS 0.008001f
C53 B.n25 VSUBS 0.008001f
C54 B.n26 VSUBS 0.008001f
C55 B.n27 VSUBS 0.008001f
C56 B.n28 VSUBS 0.008001f
C57 B.n29 VSUBS 0.008001f
C58 B.t2 VSUBS 0.34762f
C59 B.t1 VSUBS 0.35352f
C60 B.t0 VSUBS 0.125893f
C61 B.n30 VSUBS 0.099413f
C62 B.n31 VSUBS 0.070878f
C63 B.n32 VSUBS 0.008001f
C64 B.n33 VSUBS 0.008001f
C65 B.n34 VSUBS 0.008001f
C66 B.n35 VSUBS 0.008001f
C67 B.t11 VSUBS 0.347616f
C68 B.t10 VSUBS 0.353515f
C69 B.t9 VSUBS 0.125893f
C70 B.n36 VSUBS 0.099418f
C71 B.n37 VSUBS 0.070883f
C72 B.n38 VSUBS 0.008001f
C73 B.n39 VSUBS 0.008001f
C74 B.n40 VSUBS 0.008001f
C75 B.n41 VSUBS 0.008001f
C76 B.n42 VSUBS 0.008001f
C77 B.n43 VSUBS 0.008001f
C78 B.n44 VSUBS 0.008001f
C79 B.n45 VSUBS 0.008001f
C80 B.n46 VSUBS 0.008001f
C81 B.n47 VSUBS 0.008001f
C82 B.n48 VSUBS 0.008001f
C83 B.n49 VSUBS 0.008001f
C84 B.n50 VSUBS 0.008001f
C85 B.n51 VSUBS 0.008001f
C86 B.n52 VSUBS 0.008001f
C87 B.n53 VSUBS 0.008001f
C88 B.n54 VSUBS 0.008001f
C89 B.n55 VSUBS 0.017453f
C90 B.n56 VSUBS 0.008001f
C91 B.n57 VSUBS 0.008001f
C92 B.n58 VSUBS 0.008001f
C93 B.n59 VSUBS 0.008001f
C94 B.n60 VSUBS 0.008001f
C95 B.n61 VSUBS 0.008001f
C96 B.n62 VSUBS 0.008001f
C97 B.n63 VSUBS 0.008001f
C98 B.n64 VSUBS 0.008001f
C99 B.n65 VSUBS 0.008001f
C100 B.n66 VSUBS 0.008001f
C101 B.n67 VSUBS 0.008001f
C102 B.n68 VSUBS 0.008001f
C103 B.n69 VSUBS 0.008001f
C104 B.n70 VSUBS 0.008001f
C105 B.n71 VSUBS 0.008001f
C106 B.n72 VSUBS 0.008001f
C107 B.n73 VSUBS 0.008001f
C108 B.n74 VSUBS 0.017453f
C109 B.n75 VSUBS 0.008001f
C110 B.n76 VSUBS 0.008001f
C111 B.n77 VSUBS 0.008001f
C112 B.n78 VSUBS 0.008001f
C113 B.n79 VSUBS 0.008001f
C114 B.n80 VSUBS 0.008001f
C115 B.n81 VSUBS 0.008001f
C116 B.n82 VSUBS 0.008001f
C117 B.n83 VSUBS 0.008001f
C118 B.n84 VSUBS 0.008001f
C119 B.n85 VSUBS 0.008001f
C120 B.n86 VSUBS 0.008001f
C121 B.n87 VSUBS 0.008001f
C122 B.n88 VSUBS 0.008001f
C123 B.n89 VSUBS 0.008001f
C124 B.n90 VSUBS 0.008001f
C125 B.n91 VSUBS 0.008001f
C126 B.t7 VSUBS 0.347616f
C127 B.t8 VSUBS 0.353515f
C128 B.t6 VSUBS 0.125893f
C129 B.n92 VSUBS 0.099418f
C130 B.n93 VSUBS 0.070883f
C131 B.n94 VSUBS 0.018537f
C132 B.n95 VSUBS 0.008001f
C133 B.n96 VSUBS 0.008001f
C134 B.n97 VSUBS 0.008001f
C135 B.n98 VSUBS 0.008001f
C136 B.n99 VSUBS 0.008001f
C137 B.t4 VSUBS 0.34762f
C138 B.t5 VSUBS 0.35352f
C139 B.t3 VSUBS 0.125893f
C140 B.n100 VSUBS 0.099413f
C141 B.n101 VSUBS 0.070878f
C142 B.n102 VSUBS 0.008001f
C143 B.n103 VSUBS 0.008001f
C144 B.n104 VSUBS 0.008001f
C145 B.n105 VSUBS 0.008001f
C146 B.n106 VSUBS 0.008001f
C147 B.n107 VSUBS 0.008001f
C148 B.n108 VSUBS 0.008001f
C149 B.n109 VSUBS 0.008001f
C150 B.n110 VSUBS 0.008001f
C151 B.n111 VSUBS 0.008001f
C152 B.n112 VSUBS 0.008001f
C153 B.n113 VSUBS 0.008001f
C154 B.n114 VSUBS 0.008001f
C155 B.n115 VSUBS 0.008001f
C156 B.n116 VSUBS 0.008001f
C157 B.n117 VSUBS 0.008001f
C158 B.n118 VSUBS 0.018786f
C159 B.n119 VSUBS 0.008001f
C160 B.n120 VSUBS 0.008001f
C161 B.n121 VSUBS 0.008001f
C162 B.n122 VSUBS 0.008001f
C163 B.n123 VSUBS 0.008001f
C164 B.n124 VSUBS 0.008001f
C165 B.n125 VSUBS 0.008001f
C166 B.n126 VSUBS 0.008001f
C167 B.n127 VSUBS 0.008001f
C168 B.n128 VSUBS 0.008001f
C169 B.n129 VSUBS 0.008001f
C170 B.n130 VSUBS 0.008001f
C171 B.n131 VSUBS 0.008001f
C172 B.n132 VSUBS 0.008001f
C173 B.n133 VSUBS 0.008001f
C174 B.n134 VSUBS 0.008001f
C175 B.n135 VSUBS 0.008001f
C176 B.n136 VSUBS 0.008001f
C177 B.n137 VSUBS 0.008001f
C178 B.n138 VSUBS 0.008001f
C179 B.n139 VSUBS 0.008001f
C180 B.n140 VSUBS 0.008001f
C181 B.n141 VSUBS 0.008001f
C182 B.n142 VSUBS 0.008001f
C183 B.n143 VSUBS 0.008001f
C184 B.n144 VSUBS 0.008001f
C185 B.n145 VSUBS 0.008001f
C186 B.n146 VSUBS 0.008001f
C187 B.n147 VSUBS 0.008001f
C188 B.n148 VSUBS 0.008001f
C189 B.n149 VSUBS 0.008001f
C190 B.n150 VSUBS 0.008001f
C191 B.n151 VSUBS 0.008001f
C192 B.n152 VSUBS 0.008001f
C193 B.n153 VSUBS 0.017453f
C194 B.n154 VSUBS 0.017453f
C195 B.n155 VSUBS 0.018786f
C196 B.n156 VSUBS 0.008001f
C197 B.n157 VSUBS 0.008001f
C198 B.n158 VSUBS 0.008001f
C199 B.n159 VSUBS 0.008001f
C200 B.n160 VSUBS 0.008001f
C201 B.n161 VSUBS 0.008001f
C202 B.n162 VSUBS 0.008001f
C203 B.n163 VSUBS 0.008001f
C204 B.n164 VSUBS 0.008001f
C205 B.n165 VSUBS 0.008001f
C206 B.n166 VSUBS 0.008001f
C207 B.n167 VSUBS 0.008001f
C208 B.n168 VSUBS 0.008001f
C209 B.n169 VSUBS 0.008001f
C210 B.n170 VSUBS 0.008001f
C211 B.n171 VSUBS 0.008001f
C212 B.n172 VSUBS 0.008001f
C213 B.n173 VSUBS 0.008001f
C214 B.n174 VSUBS 0.008001f
C215 B.n175 VSUBS 0.008001f
C216 B.n176 VSUBS 0.008001f
C217 B.n177 VSUBS 0.008001f
C218 B.n178 VSUBS 0.008001f
C219 B.n179 VSUBS 0.008001f
C220 B.n180 VSUBS 0.008001f
C221 B.n181 VSUBS 0.008001f
C222 B.n182 VSUBS 0.008001f
C223 B.n183 VSUBS 0.008001f
C224 B.n184 VSUBS 0.008001f
C225 B.n185 VSUBS 0.008001f
C226 B.n186 VSUBS 0.008001f
C227 B.n187 VSUBS 0.008001f
C228 B.n188 VSUBS 0.008001f
C229 B.n189 VSUBS 0.008001f
C230 B.n190 VSUBS 0.008001f
C231 B.n191 VSUBS 0.008001f
C232 B.n192 VSUBS 0.008001f
C233 B.n193 VSUBS 0.008001f
C234 B.n194 VSUBS 0.008001f
C235 B.n195 VSUBS 0.008001f
C236 B.n196 VSUBS 0.008001f
C237 B.n197 VSUBS 0.008001f
C238 B.n198 VSUBS 0.008001f
C239 B.n199 VSUBS 0.008001f
C240 B.n200 VSUBS 0.008001f
C241 B.n201 VSUBS 0.008001f
C242 B.n202 VSUBS 0.008001f
C243 B.n203 VSUBS 0.008001f
C244 B.n204 VSUBS 0.008001f
C245 B.n205 VSUBS 0.008001f
C246 B.n206 VSUBS 0.00553f
C247 B.n207 VSUBS 0.018537f
C248 B.n208 VSUBS 0.006471f
C249 B.n209 VSUBS 0.008001f
C250 B.n210 VSUBS 0.008001f
C251 B.n211 VSUBS 0.008001f
C252 B.n212 VSUBS 0.008001f
C253 B.n213 VSUBS 0.008001f
C254 B.n214 VSUBS 0.008001f
C255 B.n215 VSUBS 0.008001f
C256 B.n216 VSUBS 0.008001f
C257 B.n217 VSUBS 0.008001f
C258 B.n218 VSUBS 0.008001f
C259 B.n219 VSUBS 0.008001f
C260 B.n220 VSUBS 0.006471f
C261 B.n221 VSUBS 0.008001f
C262 B.n222 VSUBS 0.008001f
C263 B.n223 VSUBS 0.00553f
C264 B.n224 VSUBS 0.008001f
C265 B.n225 VSUBS 0.008001f
C266 B.n226 VSUBS 0.008001f
C267 B.n227 VSUBS 0.008001f
C268 B.n228 VSUBS 0.008001f
C269 B.n229 VSUBS 0.008001f
C270 B.n230 VSUBS 0.008001f
C271 B.n231 VSUBS 0.008001f
C272 B.n232 VSUBS 0.008001f
C273 B.n233 VSUBS 0.008001f
C274 B.n234 VSUBS 0.008001f
C275 B.n235 VSUBS 0.008001f
C276 B.n236 VSUBS 0.008001f
C277 B.n237 VSUBS 0.008001f
C278 B.n238 VSUBS 0.008001f
C279 B.n239 VSUBS 0.008001f
C280 B.n240 VSUBS 0.008001f
C281 B.n241 VSUBS 0.008001f
C282 B.n242 VSUBS 0.008001f
C283 B.n243 VSUBS 0.008001f
C284 B.n244 VSUBS 0.008001f
C285 B.n245 VSUBS 0.008001f
C286 B.n246 VSUBS 0.008001f
C287 B.n247 VSUBS 0.008001f
C288 B.n248 VSUBS 0.008001f
C289 B.n249 VSUBS 0.008001f
C290 B.n250 VSUBS 0.008001f
C291 B.n251 VSUBS 0.008001f
C292 B.n252 VSUBS 0.008001f
C293 B.n253 VSUBS 0.008001f
C294 B.n254 VSUBS 0.008001f
C295 B.n255 VSUBS 0.008001f
C296 B.n256 VSUBS 0.008001f
C297 B.n257 VSUBS 0.008001f
C298 B.n258 VSUBS 0.008001f
C299 B.n259 VSUBS 0.008001f
C300 B.n260 VSUBS 0.008001f
C301 B.n261 VSUBS 0.008001f
C302 B.n262 VSUBS 0.008001f
C303 B.n263 VSUBS 0.008001f
C304 B.n264 VSUBS 0.008001f
C305 B.n265 VSUBS 0.008001f
C306 B.n266 VSUBS 0.008001f
C307 B.n267 VSUBS 0.008001f
C308 B.n268 VSUBS 0.008001f
C309 B.n269 VSUBS 0.008001f
C310 B.n270 VSUBS 0.008001f
C311 B.n271 VSUBS 0.008001f
C312 B.n272 VSUBS 0.008001f
C313 B.n273 VSUBS 0.018786f
C314 B.n274 VSUBS 0.018786f
C315 B.n275 VSUBS 0.017453f
C316 B.n276 VSUBS 0.008001f
C317 B.n277 VSUBS 0.008001f
C318 B.n278 VSUBS 0.008001f
C319 B.n279 VSUBS 0.008001f
C320 B.n280 VSUBS 0.008001f
C321 B.n281 VSUBS 0.008001f
C322 B.n282 VSUBS 0.008001f
C323 B.n283 VSUBS 0.008001f
C324 B.n284 VSUBS 0.008001f
C325 B.n285 VSUBS 0.008001f
C326 B.n286 VSUBS 0.008001f
C327 B.n287 VSUBS 0.008001f
C328 B.n288 VSUBS 0.008001f
C329 B.n289 VSUBS 0.008001f
C330 B.n290 VSUBS 0.008001f
C331 B.n291 VSUBS 0.008001f
C332 B.n292 VSUBS 0.008001f
C333 B.n293 VSUBS 0.008001f
C334 B.n294 VSUBS 0.008001f
C335 B.n295 VSUBS 0.008001f
C336 B.n296 VSUBS 0.008001f
C337 B.n297 VSUBS 0.008001f
C338 B.n298 VSUBS 0.008001f
C339 B.n299 VSUBS 0.008001f
C340 B.n300 VSUBS 0.008001f
C341 B.n301 VSUBS 0.008001f
C342 B.n302 VSUBS 0.008001f
C343 B.n303 VSUBS 0.008001f
C344 B.n304 VSUBS 0.008001f
C345 B.n305 VSUBS 0.008001f
C346 B.n306 VSUBS 0.008001f
C347 B.n307 VSUBS 0.008001f
C348 B.n308 VSUBS 0.008001f
C349 B.n309 VSUBS 0.008001f
C350 B.n310 VSUBS 0.008001f
C351 B.n311 VSUBS 0.008001f
C352 B.n312 VSUBS 0.008001f
C353 B.n313 VSUBS 0.008001f
C354 B.n314 VSUBS 0.008001f
C355 B.n315 VSUBS 0.008001f
C356 B.n316 VSUBS 0.008001f
C357 B.n317 VSUBS 0.008001f
C358 B.n318 VSUBS 0.008001f
C359 B.n319 VSUBS 0.008001f
C360 B.n320 VSUBS 0.008001f
C361 B.n321 VSUBS 0.008001f
C362 B.n322 VSUBS 0.008001f
C363 B.n323 VSUBS 0.008001f
C364 B.n324 VSUBS 0.008001f
C365 B.n325 VSUBS 0.008001f
C366 B.n326 VSUBS 0.008001f
C367 B.n327 VSUBS 0.008001f
C368 B.n328 VSUBS 0.008001f
C369 B.n329 VSUBS 0.008001f
C370 B.n330 VSUBS 0.008001f
C371 B.n331 VSUBS 0.008001f
C372 B.n332 VSUBS 0.018446f
C373 B.n333 VSUBS 0.017792f
C374 B.n334 VSUBS 0.018786f
C375 B.n335 VSUBS 0.008001f
C376 B.n336 VSUBS 0.008001f
C377 B.n337 VSUBS 0.008001f
C378 B.n338 VSUBS 0.008001f
C379 B.n339 VSUBS 0.008001f
C380 B.n340 VSUBS 0.008001f
C381 B.n341 VSUBS 0.008001f
C382 B.n342 VSUBS 0.008001f
C383 B.n343 VSUBS 0.008001f
C384 B.n344 VSUBS 0.008001f
C385 B.n345 VSUBS 0.008001f
C386 B.n346 VSUBS 0.008001f
C387 B.n347 VSUBS 0.008001f
C388 B.n348 VSUBS 0.008001f
C389 B.n349 VSUBS 0.008001f
C390 B.n350 VSUBS 0.008001f
C391 B.n351 VSUBS 0.008001f
C392 B.n352 VSUBS 0.008001f
C393 B.n353 VSUBS 0.008001f
C394 B.n354 VSUBS 0.008001f
C395 B.n355 VSUBS 0.008001f
C396 B.n356 VSUBS 0.008001f
C397 B.n357 VSUBS 0.008001f
C398 B.n358 VSUBS 0.008001f
C399 B.n359 VSUBS 0.008001f
C400 B.n360 VSUBS 0.008001f
C401 B.n361 VSUBS 0.008001f
C402 B.n362 VSUBS 0.008001f
C403 B.n363 VSUBS 0.008001f
C404 B.n364 VSUBS 0.008001f
C405 B.n365 VSUBS 0.008001f
C406 B.n366 VSUBS 0.008001f
C407 B.n367 VSUBS 0.008001f
C408 B.n368 VSUBS 0.008001f
C409 B.n369 VSUBS 0.008001f
C410 B.n370 VSUBS 0.008001f
C411 B.n371 VSUBS 0.008001f
C412 B.n372 VSUBS 0.008001f
C413 B.n373 VSUBS 0.008001f
C414 B.n374 VSUBS 0.008001f
C415 B.n375 VSUBS 0.008001f
C416 B.n376 VSUBS 0.008001f
C417 B.n377 VSUBS 0.008001f
C418 B.n378 VSUBS 0.008001f
C419 B.n379 VSUBS 0.008001f
C420 B.n380 VSUBS 0.008001f
C421 B.n381 VSUBS 0.008001f
C422 B.n382 VSUBS 0.008001f
C423 B.n383 VSUBS 0.008001f
C424 B.n384 VSUBS 0.008001f
C425 B.n385 VSUBS 0.00553f
C426 B.n386 VSUBS 0.018537f
C427 B.n387 VSUBS 0.006471f
C428 B.n388 VSUBS 0.008001f
C429 B.n389 VSUBS 0.008001f
C430 B.n390 VSUBS 0.008001f
C431 B.n391 VSUBS 0.008001f
C432 B.n392 VSUBS 0.008001f
C433 B.n393 VSUBS 0.008001f
C434 B.n394 VSUBS 0.008001f
C435 B.n395 VSUBS 0.008001f
C436 B.n396 VSUBS 0.008001f
C437 B.n397 VSUBS 0.008001f
C438 B.n398 VSUBS 0.008001f
C439 B.n399 VSUBS 0.006471f
C440 B.n400 VSUBS 0.018537f
C441 B.n401 VSUBS 0.00553f
C442 B.n402 VSUBS 0.008001f
C443 B.n403 VSUBS 0.008001f
C444 B.n404 VSUBS 0.008001f
C445 B.n405 VSUBS 0.008001f
C446 B.n406 VSUBS 0.008001f
C447 B.n407 VSUBS 0.008001f
C448 B.n408 VSUBS 0.008001f
C449 B.n409 VSUBS 0.008001f
C450 B.n410 VSUBS 0.008001f
C451 B.n411 VSUBS 0.008001f
C452 B.n412 VSUBS 0.008001f
C453 B.n413 VSUBS 0.008001f
C454 B.n414 VSUBS 0.008001f
C455 B.n415 VSUBS 0.008001f
C456 B.n416 VSUBS 0.008001f
C457 B.n417 VSUBS 0.008001f
C458 B.n418 VSUBS 0.008001f
C459 B.n419 VSUBS 0.008001f
C460 B.n420 VSUBS 0.008001f
C461 B.n421 VSUBS 0.008001f
C462 B.n422 VSUBS 0.008001f
C463 B.n423 VSUBS 0.008001f
C464 B.n424 VSUBS 0.008001f
C465 B.n425 VSUBS 0.008001f
C466 B.n426 VSUBS 0.008001f
C467 B.n427 VSUBS 0.008001f
C468 B.n428 VSUBS 0.008001f
C469 B.n429 VSUBS 0.008001f
C470 B.n430 VSUBS 0.008001f
C471 B.n431 VSUBS 0.008001f
C472 B.n432 VSUBS 0.008001f
C473 B.n433 VSUBS 0.008001f
C474 B.n434 VSUBS 0.008001f
C475 B.n435 VSUBS 0.008001f
C476 B.n436 VSUBS 0.008001f
C477 B.n437 VSUBS 0.008001f
C478 B.n438 VSUBS 0.008001f
C479 B.n439 VSUBS 0.008001f
C480 B.n440 VSUBS 0.008001f
C481 B.n441 VSUBS 0.008001f
C482 B.n442 VSUBS 0.008001f
C483 B.n443 VSUBS 0.008001f
C484 B.n444 VSUBS 0.008001f
C485 B.n445 VSUBS 0.008001f
C486 B.n446 VSUBS 0.008001f
C487 B.n447 VSUBS 0.008001f
C488 B.n448 VSUBS 0.008001f
C489 B.n449 VSUBS 0.008001f
C490 B.n450 VSUBS 0.008001f
C491 B.n451 VSUBS 0.008001f
C492 B.n452 VSUBS 0.018786f
C493 B.n453 VSUBS 0.018786f
C494 B.n454 VSUBS 0.017453f
C495 B.n455 VSUBS 0.008001f
C496 B.n456 VSUBS 0.008001f
C497 B.n457 VSUBS 0.008001f
C498 B.n458 VSUBS 0.008001f
C499 B.n459 VSUBS 0.008001f
C500 B.n460 VSUBS 0.008001f
C501 B.n461 VSUBS 0.008001f
C502 B.n462 VSUBS 0.008001f
C503 B.n463 VSUBS 0.008001f
C504 B.n464 VSUBS 0.008001f
C505 B.n465 VSUBS 0.008001f
C506 B.n466 VSUBS 0.008001f
C507 B.n467 VSUBS 0.008001f
C508 B.n468 VSUBS 0.008001f
C509 B.n469 VSUBS 0.008001f
C510 B.n470 VSUBS 0.008001f
C511 B.n471 VSUBS 0.008001f
C512 B.n472 VSUBS 0.008001f
C513 B.n473 VSUBS 0.008001f
C514 B.n474 VSUBS 0.008001f
C515 B.n475 VSUBS 0.008001f
C516 B.n476 VSUBS 0.008001f
C517 B.n477 VSUBS 0.008001f
C518 B.n478 VSUBS 0.008001f
C519 B.n479 VSUBS 0.008001f
C520 B.n480 VSUBS 0.008001f
C521 B.n481 VSUBS 0.008001f
C522 B.n482 VSUBS 0.008001f
C523 B.n483 VSUBS 0.018116f
C524 VDD1.t5 VSUBS 2.24102f
C525 VDD1.t4 VSUBS 0.227575f
C526 VDD1.t6 VSUBS 0.227575f
C527 VDD1.n0 VSUBS 1.70356f
C528 VDD1.n1 VSUBS 1.29381f
C529 VDD1.t2 VSUBS 2.24101f
C530 VDD1.t7 VSUBS 0.227575f
C531 VDD1.t1 VSUBS 0.227575f
C532 VDD1.n2 VSUBS 1.70355f
C533 VDD1.n3 VSUBS 1.29173f
C534 VDD1.t0 VSUBS 0.227575f
C535 VDD1.t3 VSUBS 0.227575f
C536 VDD1.n4 VSUBS 1.70638f
C537 VDD1.n5 VSUBS 2.21628f
C538 VDD1.t8 VSUBS 0.227575f
C539 VDD1.t9 VSUBS 0.227575f
C540 VDD1.n6 VSUBS 1.70355f
C541 VDD1.n7 VSUBS 2.72679f
C542 VP.n0 VSUBS 0.070198f
C543 VP.t9 VSUBS 0.553012f
C544 VP.t8 VSUBS 0.553012f
C545 VP.n1 VSUBS 0.02848f
C546 VP.n2 VSUBS 0.070198f
C547 VP.t1 VSUBS 0.553012f
C548 VP.t3 VSUBS 0.553012f
C549 VP.n3 VSUBS 0.02848f
C550 VP.t4 VSUBS 0.56159f
C551 VP.t5 VSUBS 0.553012f
C552 VP.n4 VSUBS 0.228925f
C553 VP.n5 VSUBS 0.250222f
C554 VP.n6 VSUBS 0.151985f
C555 VP.n7 VSUBS 0.070198f
C556 VP.n8 VSUBS 0.252211f
C557 VP.n9 VSUBS 0.02848f
C558 VP.n10 VSUBS 0.228925f
C559 VP.t0 VSUBS 0.56159f
C560 VP.n11 VSUBS 0.250126f
C561 VP.n12 VSUBS 2.52549f
C562 VP.t7 VSUBS 0.56159f
C563 VP.t2 VSUBS 0.553012f
C564 VP.n13 VSUBS 0.228925f
C565 VP.n14 VSUBS 0.250126f
C566 VP.n15 VSUBS 2.59058f
C567 VP.n16 VSUBS 0.070198f
C568 VP.n17 VSUBS 0.070198f
C569 VP.n18 VSUBS 0.252211f
C570 VP.n19 VSUBS 0.02848f
C571 VP.n20 VSUBS 0.228925f
C572 VP.t6 VSUBS 0.56159f
C573 VP.n21 VSUBS 0.250126f
C574 VP.n22 VSUBS 0.054401f
C575 VDD2.t4 VSUBS 2.2422f
C576 VDD2.t2 VSUBS 0.227695f
C577 VDD2.t0 VSUBS 0.227695f
C578 VDD2.n0 VSUBS 1.70446f
C579 VDD2.n1 VSUBS 1.29242f
C580 VDD2.t1 VSUBS 0.227695f
C581 VDD2.t9 VSUBS 0.227695f
C582 VDD2.n2 VSUBS 1.70728f
C583 VDD2.n3 VSUBS 2.13682f
C584 VDD2.t7 VSUBS 2.23769f
C585 VDD2.n4 VSUBS 2.75248f
C586 VDD2.t5 VSUBS 0.227695f
C587 VDD2.t8 VSUBS 0.227695f
C588 VDD2.n5 VSUBS 1.70446f
C589 VDD2.n6 VSUBS 0.608863f
C590 VDD2.t6 VSUBS 0.227695f
C591 VDD2.t3 VSUBS 0.227695f
C592 VDD2.n7 VSUBS 1.70725f
C593 VTAIL.t16 VSUBS 0.265765f
C594 VTAIL.t13 VSUBS 0.265765f
C595 VTAIL.n0 VSUBS 1.81924f
C596 VTAIL.n1 VSUBS 0.886286f
C597 VTAIL.t6 VSUBS 2.42402f
C598 VTAIL.n2 VSUBS 1.01484f
C599 VTAIL.t5 VSUBS 0.265765f
C600 VTAIL.t1 VSUBS 0.265765f
C601 VTAIL.n3 VSUBS 1.81924f
C602 VTAIL.n4 VSUBS 0.871918f
C603 VTAIL.t4 VSUBS 0.265765f
C604 VTAIL.t0 VSUBS 0.265765f
C605 VTAIL.n5 VSUBS 1.81924f
C606 VTAIL.n6 VSUBS 2.34289f
C607 VTAIL.t14 VSUBS 0.265765f
C608 VTAIL.t17 VSUBS 0.265765f
C609 VTAIL.n7 VSUBS 1.81924f
C610 VTAIL.n8 VSUBS 2.34288f
C611 VTAIL.t9 VSUBS 0.265765f
C612 VTAIL.t12 VSUBS 0.265765f
C613 VTAIL.n9 VSUBS 1.81924f
C614 VTAIL.n10 VSUBS 0.87191f
C615 VTAIL.t15 VSUBS 2.42403f
C616 VTAIL.n11 VSUBS 1.01483f
C617 VTAIL.t3 VSUBS 0.265765f
C618 VTAIL.t2 VSUBS 0.265765f
C619 VTAIL.n12 VSUBS 1.81924f
C620 VTAIL.n13 VSUBS 0.894803f
C621 VTAIL.t19 VSUBS 0.265765f
C622 VTAIL.t18 VSUBS 0.265765f
C623 VTAIL.n14 VSUBS 1.81924f
C624 VTAIL.n15 VSUBS 0.87191f
C625 VTAIL.t7 VSUBS 2.42402f
C626 VTAIL.n16 VSUBS 2.40253f
C627 VTAIL.t10 VSUBS 2.42402f
C628 VTAIL.n17 VSUBS 2.40253f
C629 VTAIL.t8 VSUBS 0.265765f
C630 VTAIL.t11 VSUBS 0.265765f
C631 VTAIL.n18 VSUBS 1.81924f
C632 VTAIL.n19 VSUBS 0.820045f
C633 VN.n0 VSUBS 0.068184f
C634 VN.t8 VSUBS 0.53715f
C635 VN.t9 VSUBS 0.53715f
C636 VN.n1 VSUBS 0.027664f
C637 VN.t5 VSUBS 0.545481f
C638 VN.t7 VSUBS 0.53715f
C639 VN.n2 VSUBS 0.222358f
C640 VN.n3 VSUBS 0.243045f
C641 VN.n4 VSUBS 0.147625f
C642 VN.n5 VSUBS 0.068184f
C643 VN.n6 VSUBS 0.244977f
C644 VN.n7 VSUBS 0.027664f
C645 VN.n8 VSUBS 0.222358f
C646 VN.t0 VSUBS 0.545481f
C647 VN.n9 VSUBS 0.242951f
C648 VN.n10 VSUBS 0.05284f
C649 VN.n11 VSUBS 0.068184f
C650 VN.t2 VSUBS 0.545481f
C651 VN.t4 VSUBS 0.53715f
C652 VN.t1 VSUBS 0.53715f
C653 VN.n12 VSUBS 0.027664f
C654 VN.t3 VSUBS 0.53715f
C655 VN.n13 VSUBS 0.222358f
C656 VN.t6 VSUBS 0.545481f
C657 VN.n14 VSUBS 0.243045f
C658 VN.n15 VSUBS 0.147625f
C659 VN.n16 VSUBS 0.068184f
C660 VN.n17 VSUBS 0.244977f
C661 VN.n18 VSUBS 0.027664f
C662 VN.n19 VSUBS 0.222358f
C663 VN.n20 VSUBS 0.242951f
C664 VN.n21 VSUBS 2.49804f
.ends

