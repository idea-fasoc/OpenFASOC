* NGSPICE file created from diff_pair_sample_1038.ext - technology: sky130A

.subckt diff_pair_sample_1038 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t3 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=1.35465 ps=8.54 w=8.21 l=1.25
X1 VTAIL.t0 VN.t0 VDD2.t3 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=1.35465 ps=8.54 w=8.21 l=1.25
X2 VDD2.t2 VN.t1 VTAIL.t3 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=1.35465 pd=8.54 as=3.2019 ps=17.2 w=8.21 l=1.25
X3 VTAIL.t2 VN.t2 VDD2.t1 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=1.35465 ps=8.54 w=8.21 l=1.25
X4 VDD1.t1 VP.t1 VTAIL.t6 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=1.35465 pd=8.54 as=3.2019 ps=17.2 w=8.21 l=1.25
X5 VDD2.t0 VN.t3 VTAIL.t1 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=1.35465 pd=8.54 as=3.2019 ps=17.2 w=8.21 l=1.25
X6 B.t11 B.t9 B.t10 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=0 ps=0 w=8.21 l=1.25
X7 VTAIL.t5 VP.t2 VDD1.t0 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=1.35465 ps=8.54 w=8.21 l=1.25
X8 VDD1.t2 VP.t3 VTAIL.t4 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=1.35465 pd=8.54 as=3.2019 ps=17.2 w=8.21 l=1.25
X9 B.t8 B.t6 B.t7 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=0 ps=0 w=8.21 l=1.25
X10 B.t5 B.t3 B.t4 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=0 ps=0 w=8.21 l=1.25
X11 B.t2 B.t0 B.t1 w_n1918_n2610# sky130_fd_pr__pfet_01v8 ad=3.2019 pd=17.2 as=0 ps=0 w=8.21 l=1.25
R0 VP.n2 VP.t2 195.058
R1 VP.n2 VP.t3 194.835
R2 VP.n4 VP.n3 171.577
R3 VP.n10 VP.n9 171.577
R4 VP.n8 VP.n0 161.3
R5 VP.n7 VP.n6 161.3
R6 VP.n5 VP.n1 161.3
R7 VP.n3 VP.t0 158.29
R8 VP.n9 VP.t1 158.29
R9 VP.n4 VP.n2 57.4434
R10 VP.n7 VP.n1 40.4934
R11 VP.n8 VP.n7 40.4934
R12 VP.n3 VP.n1 14.1914
R13 VP.n9 VP.n8 14.1914
R14 VP.n5 VP.n4 0.189894
R15 VP.n6 VP.n5 0.189894
R16 VP.n6 VP.n0 0.189894
R17 VP.n10 VP.n0 0.189894
R18 VP VP.n10 0.0516364
R19 VDD1 VDD1.n1 117.657
R20 VDD1 VDD1.n0 82.3126
R21 VDD1.n0 VDD1.t0 3.9597
R22 VDD1.n0 VDD1.t2 3.9597
R23 VDD1.n1 VDD1.t3 3.9597
R24 VDD1.n1 VDD1.t1 3.9597
R25 VTAIL.n5 VTAIL.t5 69.5349
R26 VTAIL.n4 VTAIL.t1 69.5349
R27 VTAIL.n3 VTAIL.t2 69.5349
R28 VTAIL.n7 VTAIL.t3 69.5348
R29 VTAIL.n0 VTAIL.t0 69.5348
R30 VTAIL.n1 VTAIL.t6 69.5348
R31 VTAIL.n2 VTAIL.t7 69.5348
R32 VTAIL.n6 VTAIL.t4 69.5348
R33 VTAIL.n7 VTAIL.n6 20.8065
R34 VTAIL.n3 VTAIL.n2 20.8065
R35 VTAIL.n4 VTAIL.n3 1.36257
R36 VTAIL.n6 VTAIL.n5 1.36257
R37 VTAIL.n2 VTAIL.n1 1.36257
R38 VTAIL VTAIL.n0 0.739724
R39 VTAIL VTAIL.n7 0.623345
R40 VTAIL.n5 VTAIL.n4 0.470328
R41 VTAIL.n1 VTAIL.n0 0.470328
R42 VN.n0 VN.t0 195.058
R43 VN.n1 VN.t3 195.058
R44 VN.n0 VN.t1 194.835
R45 VN.n1 VN.t2 194.835
R46 VN VN.n1 57.8241
R47 VN VN.n0 18.2521
R48 VDD2.n2 VDD2.n0 117.132
R49 VDD2.n2 VDD2.n1 82.2544
R50 VDD2.n1 VDD2.t1 3.9597
R51 VDD2.n1 VDD2.t0 3.9597
R52 VDD2.n0 VDD2.t3 3.9597
R53 VDD2.n0 VDD2.t2 3.9597
R54 VDD2 VDD2.n2 0.0586897
R55 B.n334 B.n53 585
R56 B.n336 B.n335 585
R57 B.n337 B.n52 585
R58 B.n339 B.n338 585
R59 B.n340 B.n51 585
R60 B.n342 B.n341 585
R61 B.n343 B.n50 585
R62 B.n345 B.n344 585
R63 B.n346 B.n49 585
R64 B.n348 B.n347 585
R65 B.n349 B.n48 585
R66 B.n351 B.n350 585
R67 B.n352 B.n47 585
R68 B.n354 B.n353 585
R69 B.n355 B.n46 585
R70 B.n357 B.n356 585
R71 B.n358 B.n45 585
R72 B.n360 B.n359 585
R73 B.n361 B.n44 585
R74 B.n363 B.n362 585
R75 B.n364 B.n43 585
R76 B.n366 B.n365 585
R77 B.n367 B.n42 585
R78 B.n369 B.n368 585
R79 B.n370 B.n41 585
R80 B.n372 B.n371 585
R81 B.n373 B.n40 585
R82 B.n375 B.n374 585
R83 B.n376 B.n39 585
R84 B.n378 B.n377 585
R85 B.n379 B.n36 585
R86 B.n382 B.n381 585
R87 B.n383 B.n35 585
R88 B.n385 B.n384 585
R89 B.n386 B.n34 585
R90 B.n388 B.n387 585
R91 B.n389 B.n33 585
R92 B.n391 B.n390 585
R93 B.n392 B.n29 585
R94 B.n394 B.n393 585
R95 B.n395 B.n28 585
R96 B.n397 B.n396 585
R97 B.n398 B.n27 585
R98 B.n400 B.n399 585
R99 B.n401 B.n26 585
R100 B.n403 B.n402 585
R101 B.n404 B.n25 585
R102 B.n406 B.n405 585
R103 B.n407 B.n24 585
R104 B.n409 B.n408 585
R105 B.n410 B.n23 585
R106 B.n412 B.n411 585
R107 B.n413 B.n22 585
R108 B.n415 B.n414 585
R109 B.n416 B.n21 585
R110 B.n418 B.n417 585
R111 B.n419 B.n20 585
R112 B.n421 B.n420 585
R113 B.n422 B.n19 585
R114 B.n424 B.n423 585
R115 B.n425 B.n18 585
R116 B.n427 B.n426 585
R117 B.n428 B.n17 585
R118 B.n430 B.n429 585
R119 B.n431 B.n16 585
R120 B.n433 B.n432 585
R121 B.n434 B.n15 585
R122 B.n436 B.n435 585
R123 B.n437 B.n14 585
R124 B.n439 B.n438 585
R125 B.n440 B.n13 585
R126 B.n333 B.n332 585
R127 B.n331 B.n54 585
R128 B.n330 B.n329 585
R129 B.n328 B.n55 585
R130 B.n327 B.n326 585
R131 B.n325 B.n56 585
R132 B.n324 B.n323 585
R133 B.n322 B.n57 585
R134 B.n321 B.n320 585
R135 B.n319 B.n58 585
R136 B.n318 B.n317 585
R137 B.n316 B.n59 585
R138 B.n315 B.n314 585
R139 B.n313 B.n60 585
R140 B.n312 B.n311 585
R141 B.n310 B.n61 585
R142 B.n309 B.n308 585
R143 B.n307 B.n62 585
R144 B.n306 B.n305 585
R145 B.n304 B.n63 585
R146 B.n303 B.n302 585
R147 B.n301 B.n64 585
R148 B.n300 B.n299 585
R149 B.n298 B.n65 585
R150 B.n297 B.n296 585
R151 B.n295 B.n66 585
R152 B.n294 B.n293 585
R153 B.n292 B.n67 585
R154 B.n291 B.n290 585
R155 B.n289 B.n68 585
R156 B.n288 B.n287 585
R157 B.n286 B.n69 585
R158 B.n285 B.n284 585
R159 B.n283 B.n70 585
R160 B.n282 B.n281 585
R161 B.n280 B.n71 585
R162 B.n279 B.n278 585
R163 B.n277 B.n72 585
R164 B.n276 B.n275 585
R165 B.n274 B.n73 585
R166 B.n273 B.n272 585
R167 B.n271 B.n74 585
R168 B.n270 B.n269 585
R169 B.n268 B.n75 585
R170 B.n267 B.n266 585
R171 B.n156 B.n113 585
R172 B.n158 B.n157 585
R173 B.n159 B.n112 585
R174 B.n161 B.n160 585
R175 B.n162 B.n111 585
R176 B.n164 B.n163 585
R177 B.n165 B.n110 585
R178 B.n167 B.n166 585
R179 B.n168 B.n109 585
R180 B.n170 B.n169 585
R181 B.n171 B.n108 585
R182 B.n173 B.n172 585
R183 B.n174 B.n107 585
R184 B.n176 B.n175 585
R185 B.n177 B.n106 585
R186 B.n179 B.n178 585
R187 B.n180 B.n105 585
R188 B.n182 B.n181 585
R189 B.n183 B.n104 585
R190 B.n185 B.n184 585
R191 B.n186 B.n103 585
R192 B.n188 B.n187 585
R193 B.n189 B.n102 585
R194 B.n191 B.n190 585
R195 B.n192 B.n101 585
R196 B.n194 B.n193 585
R197 B.n195 B.n100 585
R198 B.n197 B.n196 585
R199 B.n198 B.n99 585
R200 B.n200 B.n199 585
R201 B.n201 B.n96 585
R202 B.n204 B.n203 585
R203 B.n205 B.n95 585
R204 B.n207 B.n206 585
R205 B.n208 B.n94 585
R206 B.n210 B.n209 585
R207 B.n211 B.n93 585
R208 B.n213 B.n212 585
R209 B.n214 B.n92 585
R210 B.n219 B.n218 585
R211 B.n220 B.n91 585
R212 B.n222 B.n221 585
R213 B.n223 B.n90 585
R214 B.n225 B.n224 585
R215 B.n226 B.n89 585
R216 B.n228 B.n227 585
R217 B.n229 B.n88 585
R218 B.n231 B.n230 585
R219 B.n232 B.n87 585
R220 B.n234 B.n233 585
R221 B.n235 B.n86 585
R222 B.n237 B.n236 585
R223 B.n238 B.n85 585
R224 B.n240 B.n239 585
R225 B.n241 B.n84 585
R226 B.n243 B.n242 585
R227 B.n244 B.n83 585
R228 B.n246 B.n245 585
R229 B.n247 B.n82 585
R230 B.n249 B.n248 585
R231 B.n250 B.n81 585
R232 B.n252 B.n251 585
R233 B.n253 B.n80 585
R234 B.n255 B.n254 585
R235 B.n256 B.n79 585
R236 B.n258 B.n257 585
R237 B.n259 B.n78 585
R238 B.n261 B.n260 585
R239 B.n262 B.n77 585
R240 B.n264 B.n263 585
R241 B.n265 B.n76 585
R242 B.n155 B.n154 585
R243 B.n153 B.n114 585
R244 B.n152 B.n151 585
R245 B.n150 B.n115 585
R246 B.n149 B.n148 585
R247 B.n147 B.n116 585
R248 B.n146 B.n145 585
R249 B.n144 B.n117 585
R250 B.n143 B.n142 585
R251 B.n141 B.n118 585
R252 B.n140 B.n139 585
R253 B.n138 B.n119 585
R254 B.n137 B.n136 585
R255 B.n135 B.n120 585
R256 B.n134 B.n133 585
R257 B.n132 B.n121 585
R258 B.n131 B.n130 585
R259 B.n129 B.n122 585
R260 B.n128 B.n127 585
R261 B.n126 B.n123 585
R262 B.n125 B.n124 585
R263 B.n2 B.n0 585
R264 B.n473 B.n1 585
R265 B.n472 B.n471 585
R266 B.n470 B.n3 585
R267 B.n469 B.n468 585
R268 B.n467 B.n4 585
R269 B.n466 B.n465 585
R270 B.n464 B.n5 585
R271 B.n463 B.n462 585
R272 B.n461 B.n6 585
R273 B.n460 B.n459 585
R274 B.n458 B.n7 585
R275 B.n457 B.n456 585
R276 B.n455 B.n8 585
R277 B.n454 B.n453 585
R278 B.n452 B.n9 585
R279 B.n451 B.n450 585
R280 B.n449 B.n10 585
R281 B.n448 B.n447 585
R282 B.n446 B.n11 585
R283 B.n445 B.n444 585
R284 B.n443 B.n12 585
R285 B.n442 B.n441 585
R286 B.n475 B.n474 585
R287 B.n156 B.n155 468.476
R288 B.n442 B.n13 468.476
R289 B.n267 B.n76 468.476
R290 B.n334 B.n333 468.476
R291 B.n215 B.t9 362.659
R292 B.n97 B.t3 362.659
R293 B.n30 B.t0 362.659
R294 B.n37 B.t6 362.659
R295 B.n155 B.n114 163.367
R296 B.n151 B.n114 163.367
R297 B.n151 B.n150 163.367
R298 B.n150 B.n149 163.367
R299 B.n149 B.n116 163.367
R300 B.n145 B.n116 163.367
R301 B.n145 B.n144 163.367
R302 B.n144 B.n143 163.367
R303 B.n143 B.n118 163.367
R304 B.n139 B.n118 163.367
R305 B.n139 B.n138 163.367
R306 B.n138 B.n137 163.367
R307 B.n137 B.n120 163.367
R308 B.n133 B.n120 163.367
R309 B.n133 B.n132 163.367
R310 B.n132 B.n131 163.367
R311 B.n131 B.n122 163.367
R312 B.n127 B.n122 163.367
R313 B.n127 B.n126 163.367
R314 B.n126 B.n125 163.367
R315 B.n125 B.n2 163.367
R316 B.n474 B.n2 163.367
R317 B.n474 B.n473 163.367
R318 B.n473 B.n472 163.367
R319 B.n472 B.n3 163.367
R320 B.n468 B.n3 163.367
R321 B.n468 B.n467 163.367
R322 B.n467 B.n466 163.367
R323 B.n466 B.n5 163.367
R324 B.n462 B.n5 163.367
R325 B.n462 B.n461 163.367
R326 B.n461 B.n460 163.367
R327 B.n460 B.n7 163.367
R328 B.n456 B.n7 163.367
R329 B.n456 B.n455 163.367
R330 B.n455 B.n454 163.367
R331 B.n454 B.n9 163.367
R332 B.n450 B.n9 163.367
R333 B.n450 B.n449 163.367
R334 B.n449 B.n448 163.367
R335 B.n448 B.n11 163.367
R336 B.n444 B.n11 163.367
R337 B.n444 B.n443 163.367
R338 B.n443 B.n442 163.367
R339 B.n157 B.n156 163.367
R340 B.n157 B.n112 163.367
R341 B.n161 B.n112 163.367
R342 B.n162 B.n161 163.367
R343 B.n163 B.n162 163.367
R344 B.n163 B.n110 163.367
R345 B.n167 B.n110 163.367
R346 B.n168 B.n167 163.367
R347 B.n169 B.n168 163.367
R348 B.n169 B.n108 163.367
R349 B.n173 B.n108 163.367
R350 B.n174 B.n173 163.367
R351 B.n175 B.n174 163.367
R352 B.n175 B.n106 163.367
R353 B.n179 B.n106 163.367
R354 B.n180 B.n179 163.367
R355 B.n181 B.n180 163.367
R356 B.n181 B.n104 163.367
R357 B.n185 B.n104 163.367
R358 B.n186 B.n185 163.367
R359 B.n187 B.n186 163.367
R360 B.n187 B.n102 163.367
R361 B.n191 B.n102 163.367
R362 B.n192 B.n191 163.367
R363 B.n193 B.n192 163.367
R364 B.n193 B.n100 163.367
R365 B.n197 B.n100 163.367
R366 B.n198 B.n197 163.367
R367 B.n199 B.n198 163.367
R368 B.n199 B.n96 163.367
R369 B.n204 B.n96 163.367
R370 B.n205 B.n204 163.367
R371 B.n206 B.n205 163.367
R372 B.n206 B.n94 163.367
R373 B.n210 B.n94 163.367
R374 B.n211 B.n210 163.367
R375 B.n212 B.n211 163.367
R376 B.n212 B.n92 163.367
R377 B.n219 B.n92 163.367
R378 B.n220 B.n219 163.367
R379 B.n221 B.n220 163.367
R380 B.n221 B.n90 163.367
R381 B.n225 B.n90 163.367
R382 B.n226 B.n225 163.367
R383 B.n227 B.n226 163.367
R384 B.n227 B.n88 163.367
R385 B.n231 B.n88 163.367
R386 B.n232 B.n231 163.367
R387 B.n233 B.n232 163.367
R388 B.n233 B.n86 163.367
R389 B.n237 B.n86 163.367
R390 B.n238 B.n237 163.367
R391 B.n239 B.n238 163.367
R392 B.n239 B.n84 163.367
R393 B.n243 B.n84 163.367
R394 B.n244 B.n243 163.367
R395 B.n245 B.n244 163.367
R396 B.n245 B.n82 163.367
R397 B.n249 B.n82 163.367
R398 B.n250 B.n249 163.367
R399 B.n251 B.n250 163.367
R400 B.n251 B.n80 163.367
R401 B.n255 B.n80 163.367
R402 B.n256 B.n255 163.367
R403 B.n257 B.n256 163.367
R404 B.n257 B.n78 163.367
R405 B.n261 B.n78 163.367
R406 B.n262 B.n261 163.367
R407 B.n263 B.n262 163.367
R408 B.n263 B.n76 163.367
R409 B.n268 B.n267 163.367
R410 B.n269 B.n268 163.367
R411 B.n269 B.n74 163.367
R412 B.n273 B.n74 163.367
R413 B.n274 B.n273 163.367
R414 B.n275 B.n274 163.367
R415 B.n275 B.n72 163.367
R416 B.n279 B.n72 163.367
R417 B.n280 B.n279 163.367
R418 B.n281 B.n280 163.367
R419 B.n281 B.n70 163.367
R420 B.n285 B.n70 163.367
R421 B.n286 B.n285 163.367
R422 B.n287 B.n286 163.367
R423 B.n287 B.n68 163.367
R424 B.n291 B.n68 163.367
R425 B.n292 B.n291 163.367
R426 B.n293 B.n292 163.367
R427 B.n293 B.n66 163.367
R428 B.n297 B.n66 163.367
R429 B.n298 B.n297 163.367
R430 B.n299 B.n298 163.367
R431 B.n299 B.n64 163.367
R432 B.n303 B.n64 163.367
R433 B.n304 B.n303 163.367
R434 B.n305 B.n304 163.367
R435 B.n305 B.n62 163.367
R436 B.n309 B.n62 163.367
R437 B.n310 B.n309 163.367
R438 B.n311 B.n310 163.367
R439 B.n311 B.n60 163.367
R440 B.n315 B.n60 163.367
R441 B.n316 B.n315 163.367
R442 B.n317 B.n316 163.367
R443 B.n317 B.n58 163.367
R444 B.n321 B.n58 163.367
R445 B.n322 B.n321 163.367
R446 B.n323 B.n322 163.367
R447 B.n323 B.n56 163.367
R448 B.n327 B.n56 163.367
R449 B.n328 B.n327 163.367
R450 B.n329 B.n328 163.367
R451 B.n329 B.n54 163.367
R452 B.n333 B.n54 163.367
R453 B.n438 B.n13 163.367
R454 B.n438 B.n437 163.367
R455 B.n437 B.n436 163.367
R456 B.n436 B.n15 163.367
R457 B.n432 B.n15 163.367
R458 B.n432 B.n431 163.367
R459 B.n431 B.n430 163.367
R460 B.n430 B.n17 163.367
R461 B.n426 B.n17 163.367
R462 B.n426 B.n425 163.367
R463 B.n425 B.n424 163.367
R464 B.n424 B.n19 163.367
R465 B.n420 B.n19 163.367
R466 B.n420 B.n419 163.367
R467 B.n419 B.n418 163.367
R468 B.n418 B.n21 163.367
R469 B.n414 B.n21 163.367
R470 B.n414 B.n413 163.367
R471 B.n413 B.n412 163.367
R472 B.n412 B.n23 163.367
R473 B.n408 B.n23 163.367
R474 B.n408 B.n407 163.367
R475 B.n407 B.n406 163.367
R476 B.n406 B.n25 163.367
R477 B.n402 B.n25 163.367
R478 B.n402 B.n401 163.367
R479 B.n401 B.n400 163.367
R480 B.n400 B.n27 163.367
R481 B.n396 B.n27 163.367
R482 B.n396 B.n395 163.367
R483 B.n395 B.n394 163.367
R484 B.n394 B.n29 163.367
R485 B.n390 B.n29 163.367
R486 B.n390 B.n389 163.367
R487 B.n389 B.n388 163.367
R488 B.n388 B.n34 163.367
R489 B.n384 B.n34 163.367
R490 B.n384 B.n383 163.367
R491 B.n383 B.n382 163.367
R492 B.n382 B.n36 163.367
R493 B.n377 B.n36 163.367
R494 B.n377 B.n376 163.367
R495 B.n376 B.n375 163.367
R496 B.n375 B.n40 163.367
R497 B.n371 B.n40 163.367
R498 B.n371 B.n370 163.367
R499 B.n370 B.n369 163.367
R500 B.n369 B.n42 163.367
R501 B.n365 B.n42 163.367
R502 B.n365 B.n364 163.367
R503 B.n364 B.n363 163.367
R504 B.n363 B.n44 163.367
R505 B.n359 B.n44 163.367
R506 B.n359 B.n358 163.367
R507 B.n358 B.n357 163.367
R508 B.n357 B.n46 163.367
R509 B.n353 B.n46 163.367
R510 B.n353 B.n352 163.367
R511 B.n352 B.n351 163.367
R512 B.n351 B.n48 163.367
R513 B.n347 B.n48 163.367
R514 B.n347 B.n346 163.367
R515 B.n346 B.n345 163.367
R516 B.n345 B.n50 163.367
R517 B.n341 B.n50 163.367
R518 B.n341 B.n340 163.367
R519 B.n340 B.n339 163.367
R520 B.n339 B.n52 163.367
R521 B.n335 B.n52 163.367
R522 B.n335 B.n334 163.367
R523 B.n215 B.t11 140.133
R524 B.n37 B.t7 140.133
R525 B.n97 B.t5 140.124
R526 B.n30 B.t1 140.124
R527 B.n216 B.t10 109.49
R528 B.n38 B.t8 109.49
R529 B.n98 B.t4 109.481
R530 B.n31 B.t2 109.481
R531 B.n217 B.n216 59.5399
R532 B.n202 B.n98 59.5399
R533 B.n32 B.n31 59.5399
R534 B.n380 B.n38 59.5399
R535 B.n216 B.n215 30.6429
R536 B.n98 B.n97 30.6429
R537 B.n31 B.n30 30.6429
R538 B.n38 B.n37 30.6429
R539 B.n332 B.n53 30.4395
R540 B.n441 B.n440 30.4395
R541 B.n266 B.n265 30.4395
R542 B.n154 B.n113 30.4395
R543 B B.n475 18.0485
R544 B.n440 B.n439 10.6151
R545 B.n439 B.n14 10.6151
R546 B.n435 B.n14 10.6151
R547 B.n435 B.n434 10.6151
R548 B.n434 B.n433 10.6151
R549 B.n433 B.n16 10.6151
R550 B.n429 B.n16 10.6151
R551 B.n429 B.n428 10.6151
R552 B.n428 B.n427 10.6151
R553 B.n427 B.n18 10.6151
R554 B.n423 B.n18 10.6151
R555 B.n423 B.n422 10.6151
R556 B.n422 B.n421 10.6151
R557 B.n421 B.n20 10.6151
R558 B.n417 B.n20 10.6151
R559 B.n417 B.n416 10.6151
R560 B.n416 B.n415 10.6151
R561 B.n415 B.n22 10.6151
R562 B.n411 B.n22 10.6151
R563 B.n411 B.n410 10.6151
R564 B.n410 B.n409 10.6151
R565 B.n409 B.n24 10.6151
R566 B.n405 B.n24 10.6151
R567 B.n405 B.n404 10.6151
R568 B.n404 B.n403 10.6151
R569 B.n403 B.n26 10.6151
R570 B.n399 B.n26 10.6151
R571 B.n399 B.n398 10.6151
R572 B.n398 B.n397 10.6151
R573 B.n397 B.n28 10.6151
R574 B.n393 B.n392 10.6151
R575 B.n392 B.n391 10.6151
R576 B.n391 B.n33 10.6151
R577 B.n387 B.n33 10.6151
R578 B.n387 B.n386 10.6151
R579 B.n386 B.n385 10.6151
R580 B.n385 B.n35 10.6151
R581 B.n381 B.n35 10.6151
R582 B.n379 B.n378 10.6151
R583 B.n378 B.n39 10.6151
R584 B.n374 B.n39 10.6151
R585 B.n374 B.n373 10.6151
R586 B.n373 B.n372 10.6151
R587 B.n372 B.n41 10.6151
R588 B.n368 B.n41 10.6151
R589 B.n368 B.n367 10.6151
R590 B.n367 B.n366 10.6151
R591 B.n366 B.n43 10.6151
R592 B.n362 B.n43 10.6151
R593 B.n362 B.n361 10.6151
R594 B.n361 B.n360 10.6151
R595 B.n360 B.n45 10.6151
R596 B.n356 B.n45 10.6151
R597 B.n356 B.n355 10.6151
R598 B.n355 B.n354 10.6151
R599 B.n354 B.n47 10.6151
R600 B.n350 B.n47 10.6151
R601 B.n350 B.n349 10.6151
R602 B.n349 B.n348 10.6151
R603 B.n348 B.n49 10.6151
R604 B.n344 B.n49 10.6151
R605 B.n344 B.n343 10.6151
R606 B.n343 B.n342 10.6151
R607 B.n342 B.n51 10.6151
R608 B.n338 B.n51 10.6151
R609 B.n338 B.n337 10.6151
R610 B.n337 B.n336 10.6151
R611 B.n336 B.n53 10.6151
R612 B.n266 B.n75 10.6151
R613 B.n270 B.n75 10.6151
R614 B.n271 B.n270 10.6151
R615 B.n272 B.n271 10.6151
R616 B.n272 B.n73 10.6151
R617 B.n276 B.n73 10.6151
R618 B.n277 B.n276 10.6151
R619 B.n278 B.n277 10.6151
R620 B.n278 B.n71 10.6151
R621 B.n282 B.n71 10.6151
R622 B.n283 B.n282 10.6151
R623 B.n284 B.n283 10.6151
R624 B.n284 B.n69 10.6151
R625 B.n288 B.n69 10.6151
R626 B.n289 B.n288 10.6151
R627 B.n290 B.n289 10.6151
R628 B.n290 B.n67 10.6151
R629 B.n294 B.n67 10.6151
R630 B.n295 B.n294 10.6151
R631 B.n296 B.n295 10.6151
R632 B.n296 B.n65 10.6151
R633 B.n300 B.n65 10.6151
R634 B.n301 B.n300 10.6151
R635 B.n302 B.n301 10.6151
R636 B.n302 B.n63 10.6151
R637 B.n306 B.n63 10.6151
R638 B.n307 B.n306 10.6151
R639 B.n308 B.n307 10.6151
R640 B.n308 B.n61 10.6151
R641 B.n312 B.n61 10.6151
R642 B.n313 B.n312 10.6151
R643 B.n314 B.n313 10.6151
R644 B.n314 B.n59 10.6151
R645 B.n318 B.n59 10.6151
R646 B.n319 B.n318 10.6151
R647 B.n320 B.n319 10.6151
R648 B.n320 B.n57 10.6151
R649 B.n324 B.n57 10.6151
R650 B.n325 B.n324 10.6151
R651 B.n326 B.n325 10.6151
R652 B.n326 B.n55 10.6151
R653 B.n330 B.n55 10.6151
R654 B.n331 B.n330 10.6151
R655 B.n332 B.n331 10.6151
R656 B.n158 B.n113 10.6151
R657 B.n159 B.n158 10.6151
R658 B.n160 B.n159 10.6151
R659 B.n160 B.n111 10.6151
R660 B.n164 B.n111 10.6151
R661 B.n165 B.n164 10.6151
R662 B.n166 B.n165 10.6151
R663 B.n166 B.n109 10.6151
R664 B.n170 B.n109 10.6151
R665 B.n171 B.n170 10.6151
R666 B.n172 B.n171 10.6151
R667 B.n172 B.n107 10.6151
R668 B.n176 B.n107 10.6151
R669 B.n177 B.n176 10.6151
R670 B.n178 B.n177 10.6151
R671 B.n178 B.n105 10.6151
R672 B.n182 B.n105 10.6151
R673 B.n183 B.n182 10.6151
R674 B.n184 B.n183 10.6151
R675 B.n184 B.n103 10.6151
R676 B.n188 B.n103 10.6151
R677 B.n189 B.n188 10.6151
R678 B.n190 B.n189 10.6151
R679 B.n190 B.n101 10.6151
R680 B.n194 B.n101 10.6151
R681 B.n195 B.n194 10.6151
R682 B.n196 B.n195 10.6151
R683 B.n196 B.n99 10.6151
R684 B.n200 B.n99 10.6151
R685 B.n201 B.n200 10.6151
R686 B.n203 B.n95 10.6151
R687 B.n207 B.n95 10.6151
R688 B.n208 B.n207 10.6151
R689 B.n209 B.n208 10.6151
R690 B.n209 B.n93 10.6151
R691 B.n213 B.n93 10.6151
R692 B.n214 B.n213 10.6151
R693 B.n218 B.n214 10.6151
R694 B.n222 B.n91 10.6151
R695 B.n223 B.n222 10.6151
R696 B.n224 B.n223 10.6151
R697 B.n224 B.n89 10.6151
R698 B.n228 B.n89 10.6151
R699 B.n229 B.n228 10.6151
R700 B.n230 B.n229 10.6151
R701 B.n230 B.n87 10.6151
R702 B.n234 B.n87 10.6151
R703 B.n235 B.n234 10.6151
R704 B.n236 B.n235 10.6151
R705 B.n236 B.n85 10.6151
R706 B.n240 B.n85 10.6151
R707 B.n241 B.n240 10.6151
R708 B.n242 B.n241 10.6151
R709 B.n242 B.n83 10.6151
R710 B.n246 B.n83 10.6151
R711 B.n247 B.n246 10.6151
R712 B.n248 B.n247 10.6151
R713 B.n248 B.n81 10.6151
R714 B.n252 B.n81 10.6151
R715 B.n253 B.n252 10.6151
R716 B.n254 B.n253 10.6151
R717 B.n254 B.n79 10.6151
R718 B.n258 B.n79 10.6151
R719 B.n259 B.n258 10.6151
R720 B.n260 B.n259 10.6151
R721 B.n260 B.n77 10.6151
R722 B.n264 B.n77 10.6151
R723 B.n265 B.n264 10.6151
R724 B.n154 B.n153 10.6151
R725 B.n153 B.n152 10.6151
R726 B.n152 B.n115 10.6151
R727 B.n148 B.n115 10.6151
R728 B.n148 B.n147 10.6151
R729 B.n147 B.n146 10.6151
R730 B.n146 B.n117 10.6151
R731 B.n142 B.n117 10.6151
R732 B.n142 B.n141 10.6151
R733 B.n141 B.n140 10.6151
R734 B.n140 B.n119 10.6151
R735 B.n136 B.n119 10.6151
R736 B.n136 B.n135 10.6151
R737 B.n135 B.n134 10.6151
R738 B.n134 B.n121 10.6151
R739 B.n130 B.n121 10.6151
R740 B.n130 B.n129 10.6151
R741 B.n129 B.n128 10.6151
R742 B.n128 B.n123 10.6151
R743 B.n124 B.n123 10.6151
R744 B.n124 B.n0 10.6151
R745 B.n471 B.n1 10.6151
R746 B.n471 B.n470 10.6151
R747 B.n470 B.n469 10.6151
R748 B.n469 B.n4 10.6151
R749 B.n465 B.n4 10.6151
R750 B.n465 B.n464 10.6151
R751 B.n464 B.n463 10.6151
R752 B.n463 B.n6 10.6151
R753 B.n459 B.n6 10.6151
R754 B.n459 B.n458 10.6151
R755 B.n458 B.n457 10.6151
R756 B.n457 B.n8 10.6151
R757 B.n453 B.n8 10.6151
R758 B.n453 B.n452 10.6151
R759 B.n452 B.n451 10.6151
R760 B.n451 B.n10 10.6151
R761 B.n447 B.n10 10.6151
R762 B.n447 B.n446 10.6151
R763 B.n446 B.n445 10.6151
R764 B.n445 B.n12 10.6151
R765 B.n441 B.n12 10.6151
R766 B.n393 B.n32 6.5566
R767 B.n381 B.n380 6.5566
R768 B.n203 B.n202 6.5566
R769 B.n218 B.n217 6.5566
R770 B.n32 B.n28 4.05904
R771 B.n380 B.n379 4.05904
R772 B.n202 B.n201 4.05904
R773 B.n217 B.n91 4.05904
R774 B.n475 B.n0 2.81026
R775 B.n475 B.n1 2.81026
C0 VDD1 w_n1918_n2610# 1.07919f
C1 VP VN 4.51714f
C2 VDD2 VN 2.80529f
C3 VTAIL B 3.10774f
C4 VDD2 VP 0.308216f
C5 VTAIL w_n1918_n2610# 3.12642f
C6 VDD1 VN 0.147593f
C7 w_n1918_n2610# B 6.52154f
C8 VDD1 VP 2.96552f
C9 VDD1 VDD2 0.696497f
C10 VTAIL VN 2.65813f
C11 VTAIL VP 2.67224f
C12 VTAIL VDD2 4.52107f
C13 VN B 0.807767f
C14 VN w_n1918_n2610# 2.93281f
C15 VP B 1.20498f
C16 VDD2 B 0.951739f
C17 VTAIL VDD1 4.47591f
C18 VP w_n1918_n2610# 3.17597f
C19 VDD2 w_n1918_n2610# 1.10535f
C20 VDD1 B 0.921589f
C21 VDD2 VSUBS 0.654185f
C22 VDD1 VSUBS 4.517119f
C23 VTAIL VSUBS 0.811427f
C24 VN VSUBS 5.019741f
C25 VP VSUBS 1.429025f
C26 B VSUBS 2.78205f
C27 w_n1918_n2610# VSUBS 62.074104f
C28 B.n0 VSUBS 0.005241f
C29 B.n1 VSUBS 0.005241f
C30 B.n2 VSUBS 0.008289f
C31 B.n3 VSUBS 0.008289f
C32 B.n4 VSUBS 0.008289f
C33 B.n5 VSUBS 0.008289f
C34 B.n6 VSUBS 0.008289f
C35 B.n7 VSUBS 0.008289f
C36 B.n8 VSUBS 0.008289f
C37 B.n9 VSUBS 0.008289f
C38 B.n10 VSUBS 0.008289f
C39 B.n11 VSUBS 0.008289f
C40 B.n12 VSUBS 0.008289f
C41 B.n13 VSUBS 0.019284f
C42 B.n14 VSUBS 0.008289f
C43 B.n15 VSUBS 0.008289f
C44 B.n16 VSUBS 0.008289f
C45 B.n17 VSUBS 0.008289f
C46 B.n18 VSUBS 0.008289f
C47 B.n19 VSUBS 0.008289f
C48 B.n20 VSUBS 0.008289f
C49 B.n21 VSUBS 0.008289f
C50 B.n22 VSUBS 0.008289f
C51 B.n23 VSUBS 0.008289f
C52 B.n24 VSUBS 0.008289f
C53 B.n25 VSUBS 0.008289f
C54 B.n26 VSUBS 0.008289f
C55 B.n27 VSUBS 0.008289f
C56 B.n28 VSUBS 0.005729f
C57 B.n29 VSUBS 0.008289f
C58 B.t2 VSUBS 0.301285f
C59 B.t1 VSUBS 0.315738f
C60 B.t0 VSUBS 0.538083f
C61 B.n30 VSUBS 0.145747f
C62 B.n31 VSUBS 0.077914f
C63 B.n32 VSUBS 0.019204f
C64 B.n33 VSUBS 0.008289f
C65 B.n34 VSUBS 0.008289f
C66 B.n35 VSUBS 0.008289f
C67 B.n36 VSUBS 0.008289f
C68 B.t8 VSUBS 0.301282f
C69 B.t7 VSUBS 0.315735f
C70 B.t6 VSUBS 0.538083f
C71 B.n37 VSUBS 0.14575f
C72 B.n38 VSUBS 0.077917f
C73 B.n39 VSUBS 0.008289f
C74 B.n40 VSUBS 0.008289f
C75 B.n41 VSUBS 0.008289f
C76 B.n42 VSUBS 0.008289f
C77 B.n43 VSUBS 0.008289f
C78 B.n44 VSUBS 0.008289f
C79 B.n45 VSUBS 0.008289f
C80 B.n46 VSUBS 0.008289f
C81 B.n47 VSUBS 0.008289f
C82 B.n48 VSUBS 0.008289f
C83 B.n49 VSUBS 0.008289f
C84 B.n50 VSUBS 0.008289f
C85 B.n51 VSUBS 0.008289f
C86 B.n52 VSUBS 0.008289f
C87 B.n53 VSUBS 0.018233f
C88 B.n54 VSUBS 0.008289f
C89 B.n55 VSUBS 0.008289f
C90 B.n56 VSUBS 0.008289f
C91 B.n57 VSUBS 0.008289f
C92 B.n58 VSUBS 0.008289f
C93 B.n59 VSUBS 0.008289f
C94 B.n60 VSUBS 0.008289f
C95 B.n61 VSUBS 0.008289f
C96 B.n62 VSUBS 0.008289f
C97 B.n63 VSUBS 0.008289f
C98 B.n64 VSUBS 0.008289f
C99 B.n65 VSUBS 0.008289f
C100 B.n66 VSUBS 0.008289f
C101 B.n67 VSUBS 0.008289f
C102 B.n68 VSUBS 0.008289f
C103 B.n69 VSUBS 0.008289f
C104 B.n70 VSUBS 0.008289f
C105 B.n71 VSUBS 0.008289f
C106 B.n72 VSUBS 0.008289f
C107 B.n73 VSUBS 0.008289f
C108 B.n74 VSUBS 0.008289f
C109 B.n75 VSUBS 0.008289f
C110 B.n76 VSUBS 0.019284f
C111 B.n77 VSUBS 0.008289f
C112 B.n78 VSUBS 0.008289f
C113 B.n79 VSUBS 0.008289f
C114 B.n80 VSUBS 0.008289f
C115 B.n81 VSUBS 0.008289f
C116 B.n82 VSUBS 0.008289f
C117 B.n83 VSUBS 0.008289f
C118 B.n84 VSUBS 0.008289f
C119 B.n85 VSUBS 0.008289f
C120 B.n86 VSUBS 0.008289f
C121 B.n87 VSUBS 0.008289f
C122 B.n88 VSUBS 0.008289f
C123 B.n89 VSUBS 0.008289f
C124 B.n90 VSUBS 0.008289f
C125 B.n91 VSUBS 0.005729f
C126 B.n92 VSUBS 0.008289f
C127 B.n93 VSUBS 0.008289f
C128 B.n94 VSUBS 0.008289f
C129 B.n95 VSUBS 0.008289f
C130 B.n96 VSUBS 0.008289f
C131 B.t4 VSUBS 0.301285f
C132 B.t5 VSUBS 0.315738f
C133 B.t3 VSUBS 0.538083f
C134 B.n97 VSUBS 0.145747f
C135 B.n98 VSUBS 0.077914f
C136 B.n99 VSUBS 0.008289f
C137 B.n100 VSUBS 0.008289f
C138 B.n101 VSUBS 0.008289f
C139 B.n102 VSUBS 0.008289f
C140 B.n103 VSUBS 0.008289f
C141 B.n104 VSUBS 0.008289f
C142 B.n105 VSUBS 0.008289f
C143 B.n106 VSUBS 0.008289f
C144 B.n107 VSUBS 0.008289f
C145 B.n108 VSUBS 0.008289f
C146 B.n109 VSUBS 0.008289f
C147 B.n110 VSUBS 0.008289f
C148 B.n111 VSUBS 0.008289f
C149 B.n112 VSUBS 0.008289f
C150 B.n113 VSUBS 0.019284f
C151 B.n114 VSUBS 0.008289f
C152 B.n115 VSUBS 0.008289f
C153 B.n116 VSUBS 0.008289f
C154 B.n117 VSUBS 0.008289f
C155 B.n118 VSUBS 0.008289f
C156 B.n119 VSUBS 0.008289f
C157 B.n120 VSUBS 0.008289f
C158 B.n121 VSUBS 0.008289f
C159 B.n122 VSUBS 0.008289f
C160 B.n123 VSUBS 0.008289f
C161 B.n124 VSUBS 0.008289f
C162 B.n125 VSUBS 0.008289f
C163 B.n126 VSUBS 0.008289f
C164 B.n127 VSUBS 0.008289f
C165 B.n128 VSUBS 0.008289f
C166 B.n129 VSUBS 0.008289f
C167 B.n130 VSUBS 0.008289f
C168 B.n131 VSUBS 0.008289f
C169 B.n132 VSUBS 0.008289f
C170 B.n133 VSUBS 0.008289f
C171 B.n134 VSUBS 0.008289f
C172 B.n135 VSUBS 0.008289f
C173 B.n136 VSUBS 0.008289f
C174 B.n137 VSUBS 0.008289f
C175 B.n138 VSUBS 0.008289f
C176 B.n139 VSUBS 0.008289f
C177 B.n140 VSUBS 0.008289f
C178 B.n141 VSUBS 0.008289f
C179 B.n142 VSUBS 0.008289f
C180 B.n143 VSUBS 0.008289f
C181 B.n144 VSUBS 0.008289f
C182 B.n145 VSUBS 0.008289f
C183 B.n146 VSUBS 0.008289f
C184 B.n147 VSUBS 0.008289f
C185 B.n148 VSUBS 0.008289f
C186 B.n149 VSUBS 0.008289f
C187 B.n150 VSUBS 0.008289f
C188 B.n151 VSUBS 0.008289f
C189 B.n152 VSUBS 0.008289f
C190 B.n153 VSUBS 0.008289f
C191 B.n154 VSUBS 0.017772f
C192 B.n155 VSUBS 0.017772f
C193 B.n156 VSUBS 0.019284f
C194 B.n157 VSUBS 0.008289f
C195 B.n158 VSUBS 0.008289f
C196 B.n159 VSUBS 0.008289f
C197 B.n160 VSUBS 0.008289f
C198 B.n161 VSUBS 0.008289f
C199 B.n162 VSUBS 0.008289f
C200 B.n163 VSUBS 0.008289f
C201 B.n164 VSUBS 0.008289f
C202 B.n165 VSUBS 0.008289f
C203 B.n166 VSUBS 0.008289f
C204 B.n167 VSUBS 0.008289f
C205 B.n168 VSUBS 0.008289f
C206 B.n169 VSUBS 0.008289f
C207 B.n170 VSUBS 0.008289f
C208 B.n171 VSUBS 0.008289f
C209 B.n172 VSUBS 0.008289f
C210 B.n173 VSUBS 0.008289f
C211 B.n174 VSUBS 0.008289f
C212 B.n175 VSUBS 0.008289f
C213 B.n176 VSUBS 0.008289f
C214 B.n177 VSUBS 0.008289f
C215 B.n178 VSUBS 0.008289f
C216 B.n179 VSUBS 0.008289f
C217 B.n180 VSUBS 0.008289f
C218 B.n181 VSUBS 0.008289f
C219 B.n182 VSUBS 0.008289f
C220 B.n183 VSUBS 0.008289f
C221 B.n184 VSUBS 0.008289f
C222 B.n185 VSUBS 0.008289f
C223 B.n186 VSUBS 0.008289f
C224 B.n187 VSUBS 0.008289f
C225 B.n188 VSUBS 0.008289f
C226 B.n189 VSUBS 0.008289f
C227 B.n190 VSUBS 0.008289f
C228 B.n191 VSUBS 0.008289f
C229 B.n192 VSUBS 0.008289f
C230 B.n193 VSUBS 0.008289f
C231 B.n194 VSUBS 0.008289f
C232 B.n195 VSUBS 0.008289f
C233 B.n196 VSUBS 0.008289f
C234 B.n197 VSUBS 0.008289f
C235 B.n198 VSUBS 0.008289f
C236 B.n199 VSUBS 0.008289f
C237 B.n200 VSUBS 0.008289f
C238 B.n201 VSUBS 0.005729f
C239 B.n202 VSUBS 0.019204f
C240 B.n203 VSUBS 0.006704f
C241 B.n204 VSUBS 0.008289f
C242 B.n205 VSUBS 0.008289f
C243 B.n206 VSUBS 0.008289f
C244 B.n207 VSUBS 0.008289f
C245 B.n208 VSUBS 0.008289f
C246 B.n209 VSUBS 0.008289f
C247 B.n210 VSUBS 0.008289f
C248 B.n211 VSUBS 0.008289f
C249 B.n212 VSUBS 0.008289f
C250 B.n213 VSUBS 0.008289f
C251 B.n214 VSUBS 0.008289f
C252 B.t10 VSUBS 0.301282f
C253 B.t11 VSUBS 0.315735f
C254 B.t9 VSUBS 0.538083f
C255 B.n215 VSUBS 0.14575f
C256 B.n216 VSUBS 0.077917f
C257 B.n217 VSUBS 0.019204f
C258 B.n218 VSUBS 0.006704f
C259 B.n219 VSUBS 0.008289f
C260 B.n220 VSUBS 0.008289f
C261 B.n221 VSUBS 0.008289f
C262 B.n222 VSUBS 0.008289f
C263 B.n223 VSUBS 0.008289f
C264 B.n224 VSUBS 0.008289f
C265 B.n225 VSUBS 0.008289f
C266 B.n226 VSUBS 0.008289f
C267 B.n227 VSUBS 0.008289f
C268 B.n228 VSUBS 0.008289f
C269 B.n229 VSUBS 0.008289f
C270 B.n230 VSUBS 0.008289f
C271 B.n231 VSUBS 0.008289f
C272 B.n232 VSUBS 0.008289f
C273 B.n233 VSUBS 0.008289f
C274 B.n234 VSUBS 0.008289f
C275 B.n235 VSUBS 0.008289f
C276 B.n236 VSUBS 0.008289f
C277 B.n237 VSUBS 0.008289f
C278 B.n238 VSUBS 0.008289f
C279 B.n239 VSUBS 0.008289f
C280 B.n240 VSUBS 0.008289f
C281 B.n241 VSUBS 0.008289f
C282 B.n242 VSUBS 0.008289f
C283 B.n243 VSUBS 0.008289f
C284 B.n244 VSUBS 0.008289f
C285 B.n245 VSUBS 0.008289f
C286 B.n246 VSUBS 0.008289f
C287 B.n247 VSUBS 0.008289f
C288 B.n248 VSUBS 0.008289f
C289 B.n249 VSUBS 0.008289f
C290 B.n250 VSUBS 0.008289f
C291 B.n251 VSUBS 0.008289f
C292 B.n252 VSUBS 0.008289f
C293 B.n253 VSUBS 0.008289f
C294 B.n254 VSUBS 0.008289f
C295 B.n255 VSUBS 0.008289f
C296 B.n256 VSUBS 0.008289f
C297 B.n257 VSUBS 0.008289f
C298 B.n258 VSUBS 0.008289f
C299 B.n259 VSUBS 0.008289f
C300 B.n260 VSUBS 0.008289f
C301 B.n261 VSUBS 0.008289f
C302 B.n262 VSUBS 0.008289f
C303 B.n263 VSUBS 0.008289f
C304 B.n264 VSUBS 0.008289f
C305 B.n265 VSUBS 0.019284f
C306 B.n266 VSUBS 0.017772f
C307 B.n267 VSUBS 0.017772f
C308 B.n268 VSUBS 0.008289f
C309 B.n269 VSUBS 0.008289f
C310 B.n270 VSUBS 0.008289f
C311 B.n271 VSUBS 0.008289f
C312 B.n272 VSUBS 0.008289f
C313 B.n273 VSUBS 0.008289f
C314 B.n274 VSUBS 0.008289f
C315 B.n275 VSUBS 0.008289f
C316 B.n276 VSUBS 0.008289f
C317 B.n277 VSUBS 0.008289f
C318 B.n278 VSUBS 0.008289f
C319 B.n279 VSUBS 0.008289f
C320 B.n280 VSUBS 0.008289f
C321 B.n281 VSUBS 0.008289f
C322 B.n282 VSUBS 0.008289f
C323 B.n283 VSUBS 0.008289f
C324 B.n284 VSUBS 0.008289f
C325 B.n285 VSUBS 0.008289f
C326 B.n286 VSUBS 0.008289f
C327 B.n287 VSUBS 0.008289f
C328 B.n288 VSUBS 0.008289f
C329 B.n289 VSUBS 0.008289f
C330 B.n290 VSUBS 0.008289f
C331 B.n291 VSUBS 0.008289f
C332 B.n292 VSUBS 0.008289f
C333 B.n293 VSUBS 0.008289f
C334 B.n294 VSUBS 0.008289f
C335 B.n295 VSUBS 0.008289f
C336 B.n296 VSUBS 0.008289f
C337 B.n297 VSUBS 0.008289f
C338 B.n298 VSUBS 0.008289f
C339 B.n299 VSUBS 0.008289f
C340 B.n300 VSUBS 0.008289f
C341 B.n301 VSUBS 0.008289f
C342 B.n302 VSUBS 0.008289f
C343 B.n303 VSUBS 0.008289f
C344 B.n304 VSUBS 0.008289f
C345 B.n305 VSUBS 0.008289f
C346 B.n306 VSUBS 0.008289f
C347 B.n307 VSUBS 0.008289f
C348 B.n308 VSUBS 0.008289f
C349 B.n309 VSUBS 0.008289f
C350 B.n310 VSUBS 0.008289f
C351 B.n311 VSUBS 0.008289f
C352 B.n312 VSUBS 0.008289f
C353 B.n313 VSUBS 0.008289f
C354 B.n314 VSUBS 0.008289f
C355 B.n315 VSUBS 0.008289f
C356 B.n316 VSUBS 0.008289f
C357 B.n317 VSUBS 0.008289f
C358 B.n318 VSUBS 0.008289f
C359 B.n319 VSUBS 0.008289f
C360 B.n320 VSUBS 0.008289f
C361 B.n321 VSUBS 0.008289f
C362 B.n322 VSUBS 0.008289f
C363 B.n323 VSUBS 0.008289f
C364 B.n324 VSUBS 0.008289f
C365 B.n325 VSUBS 0.008289f
C366 B.n326 VSUBS 0.008289f
C367 B.n327 VSUBS 0.008289f
C368 B.n328 VSUBS 0.008289f
C369 B.n329 VSUBS 0.008289f
C370 B.n330 VSUBS 0.008289f
C371 B.n331 VSUBS 0.008289f
C372 B.n332 VSUBS 0.018823f
C373 B.n333 VSUBS 0.017772f
C374 B.n334 VSUBS 0.019284f
C375 B.n335 VSUBS 0.008289f
C376 B.n336 VSUBS 0.008289f
C377 B.n337 VSUBS 0.008289f
C378 B.n338 VSUBS 0.008289f
C379 B.n339 VSUBS 0.008289f
C380 B.n340 VSUBS 0.008289f
C381 B.n341 VSUBS 0.008289f
C382 B.n342 VSUBS 0.008289f
C383 B.n343 VSUBS 0.008289f
C384 B.n344 VSUBS 0.008289f
C385 B.n345 VSUBS 0.008289f
C386 B.n346 VSUBS 0.008289f
C387 B.n347 VSUBS 0.008289f
C388 B.n348 VSUBS 0.008289f
C389 B.n349 VSUBS 0.008289f
C390 B.n350 VSUBS 0.008289f
C391 B.n351 VSUBS 0.008289f
C392 B.n352 VSUBS 0.008289f
C393 B.n353 VSUBS 0.008289f
C394 B.n354 VSUBS 0.008289f
C395 B.n355 VSUBS 0.008289f
C396 B.n356 VSUBS 0.008289f
C397 B.n357 VSUBS 0.008289f
C398 B.n358 VSUBS 0.008289f
C399 B.n359 VSUBS 0.008289f
C400 B.n360 VSUBS 0.008289f
C401 B.n361 VSUBS 0.008289f
C402 B.n362 VSUBS 0.008289f
C403 B.n363 VSUBS 0.008289f
C404 B.n364 VSUBS 0.008289f
C405 B.n365 VSUBS 0.008289f
C406 B.n366 VSUBS 0.008289f
C407 B.n367 VSUBS 0.008289f
C408 B.n368 VSUBS 0.008289f
C409 B.n369 VSUBS 0.008289f
C410 B.n370 VSUBS 0.008289f
C411 B.n371 VSUBS 0.008289f
C412 B.n372 VSUBS 0.008289f
C413 B.n373 VSUBS 0.008289f
C414 B.n374 VSUBS 0.008289f
C415 B.n375 VSUBS 0.008289f
C416 B.n376 VSUBS 0.008289f
C417 B.n377 VSUBS 0.008289f
C418 B.n378 VSUBS 0.008289f
C419 B.n379 VSUBS 0.005729f
C420 B.n380 VSUBS 0.019204f
C421 B.n381 VSUBS 0.006704f
C422 B.n382 VSUBS 0.008289f
C423 B.n383 VSUBS 0.008289f
C424 B.n384 VSUBS 0.008289f
C425 B.n385 VSUBS 0.008289f
C426 B.n386 VSUBS 0.008289f
C427 B.n387 VSUBS 0.008289f
C428 B.n388 VSUBS 0.008289f
C429 B.n389 VSUBS 0.008289f
C430 B.n390 VSUBS 0.008289f
C431 B.n391 VSUBS 0.008289f
C432 B.n392 VSUBS 0.008289f
C433 B.n393 VSUBS 0.006704f
C434 B.n394 VSUBS 0.008289f
C435 B.n395 VSUBS 0.008289f
C436 B.n396 VSUBS 0.008289f
C437 B.n397 VSUBS 0.008289f
C438 B.n398 VSUBS 0.008289f
C439 B.n399 VSUBS 0.008289f
C440 B.n400 VSUBS 0.008289f
C441 B.n401 VSUBS 0.008289f
C442 B.n402 VSUBS 0.008289f
C443 B.n403 VSUBS 0.008289f
C444 B.n404 VSUBS 0.008289f
C445 B.n405 VSUBS 0.008289f
C446 B.n406 VSUBS 0.008289f
C447 B.n407 VSUBS 0.008289f
C448 B.n408 VSUBS 0.008289f
C449 B.n409 VSUBS 0.008289f
C450 B.n410 VSUBS 0.008289f
C451 B.n411 VSUBS 0.008289f
C452 B.n412 VSUBS 0.008289f
C453 B.n413 VSUBS 0.008289f
C454 B.n414 VSUBS 0.008289f
C455 B.n415 VSUBS 0.008289f
C456 B.n416 VSUBS 0.008289f
C457 B.n417 VSUBS 0.008289f
C458 B.n418 VSUBS 0.008289f
C459 B.n419 VSUBS 0.008289f
C460 B.n420 VSUBS 0.008289f
C461 B.n421 VSUBS 0.008289f
C462 B.n422 VSUBS 0.008289f
C463 B.n423 VSUBS 0.008289f
C464 B.n424 VSUBS 0.008289f
C465 B.n425 VSUBS 0.008289f
C466 B.n426 VSUBS 0.008289f
C467 B.n427 VSUBS 0.008289f
C468 B.n428 VSUBS 0.008289f
C469 B.n429 VSUBS 0.008289f
C470 B.n430 VSUBS 0.008289f
C471 B.n431 VSUBS 0.008289f
C472 B.n432 VSUBS 0.008289f
C473 B.n433 VSUBS 0.008289f
C474 B.n434 VSUBS 0.008289f
C475 B.n435 VSUBS 0.008289f
C476 B.n436 VSUBS 0.008289f
C477 B.n437 VSUBS 0.008289f
C478 B.n438 VSUBS 0.008289f
C479 B.n439 VSUBS 0.008289f
C480 B.n440 VSUBS 0.019284f
C481 B.n441 VSUBS 0.017772f
C482 B.n442 VSUBS 0.017772f
C483 B.n443 VSUBS 0.008289f
C484 B.n444 VSUBS 0.008289f
C485 B.n445 VSUBS 0.008289f
C486 B.n446 VSUBS 0.008289f
C487 B.n447 VSUBS 0.008289f
C488 B.n448 VSUBS 0.008289f
C489 B.n449 VSUBS 0.008289f
C490 B.n450 VSUBS 0.008289f
C491 B.n451 VSUBS 0.008289f
C492 B.n452 VSUBS 0.008289f
C493 B.n453 VSUBS 0.008289f
C494 B.n454 VSUBS 0.008289f
C495 B.n455 VSUBS 0.008289f
C496 B.n456 VSUBS 0.008289f
C497 B.n457 VSUBS 0.008289f
C498 B.n458 VSUBS 0.008289f
C499 B.n459 VSUBS 0.008289f
C500 B.n460 VSUBS 0.008289f
C501 B.n461 VSUBS 0.008289f
C502 B.n462 VSUBS 0.008289f
C503 B.n463 VSUBS 0.008289f
C504 B.n464 VSUBS 0.008289f
C505 B.n465 VSUBS 0.008289f
C506 B.n466 VSUBS 0.008289f
C507 B.n467 VSUBS 0.008289f
C508 B.n468 VSUBS 0.008289f
C509 B.n469 VSUBS 0.008289f
C510 B.n470 VSUBS 0.008289f
C511 B.n471 VSUBS 0.008289f
C512 B.n472 VSUBS 0.008289f
C513 B.n473 VSUBS 0.008289f
C514 B.n474 VSUBS 0.008289f
C515 B.n475 VSUBS 0.018769f
C516 VDD2.t3 VSUBS 0.174302f
C517 VDD2.t2 VSUBS 0.174302f
C518 VDD2.n0 VSUBS 1.73631f
C519 VDD2.t1 VSUBS 0.174302f
C520 VDD2.t0 VSUBS 0.174302f
C521 VDD2.n1 VSUBS 1.26663f
C522 VDD2.n2 VSUBS 3.47616f
C523 VN.t0 VSUBS 1.54334f
C524 VN.t1 VSUBS 1.54249f
C525 VN.n0 VSUBS 1.20289f
C526 VN.t3 VSUBS 1.54334f
C527 VN.t2 VSUBS 1.54249f
C528 VN.n1 VSUBS 2.66609f
C529 VTAIL.t0 VSUBS 1.39377f
C530 VTAIL.n0 VSUBS 0.656284f
C531 VTAIL.t6 VSUBS 1.39377f
C532 VTAIL.n1 VSUBS 0.70497f
C533 VTAIL.t7 VSUBS 1.39377f
C534 VTAIL.n2 VSUBS 1.65748f
C535 VTAIL.t2 VSUBS 1.39378f
C536 VTAIL.n3 VSUBS 1.65747f
C537 VTAIL.t1 VSUBS 1.39378f
C538 VTAIL.n4 VSUBS 0.70496f
C539 VTAIL.t5 VSUBS 1.39378f
C540 VTAIL.n5 VSUBS 0.70496f
C541 VTAIL.t4 VSUBS 1.39377f
C542 VTAIL.n6 VSUBS 1.65748f
C543 VTAIL.t3 VSUBS 1.39377f
C544 VTAIL.n7 VSUBS 1.5997f
C545 VDD1.t0 VSUBS 0.176676f
C546 VDD1.t2 VSUBS 0.176676f
C547 VDD1.n0 VSUBS 1.28431f
C548 VDD1.t3 VSUBS 0.176676f
C549 VDD1.t1 VSUBS 0.176676f
C550 VDD1.n1 VSUBS 1.78162f
C551 VP.n0 VSUBS 0.053384f
C552 VP.t1 VSUBS 1.47301f
C553 VP.n1 VSUBS 0.08547f
C554 VP.t2 VSUBS 1.61214f
C555 VP.t3 VSUBS 1.61125f
C556 VP.n2 VSUBS 2.75623f
C557 VP.t0 VSUBS 1.47301f
C558 VP.n3 VSUBS 0.658135f
C559 VP.n4 VSUBS 2.71338f
C560 VP.n5 VSUBS 0.053384f
C561 VP.n6 VSUBS 0.053384f
C562 VP.n7 VSUBS 0.043156f
C563 VP.n8 VSUBS 0.08547f
C564 VP.n9 VSUBS 0.658135f
C565 VP.n10 VSUBS 0.047565f
.ends

