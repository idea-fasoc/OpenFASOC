* NGSPICE file created from diff_pair_sample_1295.ext - technology: sky130A

.subckt diff_pair_sample_1295 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=0 ps=0 w=17.08 l=3.67
X1 VTAIL.t14 VN.t0 VDD2.t7 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X2 VTAIL.t2 VP.t0 VDD1.t7 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X3 VTAIL.t13 VN.t1 VDD2.t3 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=2.8182 ps=17.41 w=17.08 l=3.67
X4 VTAIL.t12 VN.t2 VDD2.t0 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=2.8182 ps=17.41 w=17.08 l=3.67
X5 VTAIL.t5 VP.t1 VDD1.t6 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=2.8182 ps=17.41 w=17.08 l=3.67
X6 B.t8 B.t6 B.t7 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=0 ps=0 w=17.08 l=3.67
X7 VDD2.t1 VN.t3 VTAIL.t11 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X8 VDD1.t5 VP.t2 VTAIL.t6 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=6.6612 ps=34.94 w=17.08 l=3.67
X9 VDD2.t2 VN.t4 VTAIL.t10 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=6.6612 ps=34.94 w=17.08 l=3.67
X10 VDD1.t4 VP.t3 VTAIL.t4 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=6.6612 ps=34.94 w=17.08 l=3.67
X11 VTAIL.t9 VN.t5 VDD2.t4 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X12 VDD1.t3 VP.t4 VTAIL.t15 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X13 VTAIL.t3 VP.t5 VDD1.t2 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X14 VDD2.t6 VN.t6 VTAIL.t8 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X15 VDD2.t5 VN.t7 VTAIL.t7 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=6.6612 ps=34.94 w=17.08 l=3.67
X16 VDD1.t1 VP.t6 VTAIL.t0 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=2.8182 pd=17.41 as=2.8182 ps=17.41 w=17.08 l=3.67
X17 B.t5 B.t3 B.t4 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=0 ps=0 w=17.08 l=3.67
X18 VTAIL.t1 VP.t7 VDD1.t0 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=2.8182 ps=17.41 w=17.08 l=3.67
X19 B.t2 B.t0 B.t1 w_n4970_n4384# sky130_fd_pr__pfet_01v8 ad=6.6612 pd=34.94 as=0 ps=0 w=17.08 l=3.67
R0 B.n756 B.n101 585
R1 B.n758 B.n757 585
R2 B.n759 B.n100 585
R3 B.n761 B.n760 585
R4 B.n762 B.n99 585
R5 B.n764 B.n763 585
R6 B.n765 B.n98 585
R7 B.n767 B.n766 585
R8 B.n768 B.n97 585
R9 B.n770 B.n769 585
R10 B.n771 B.n96 585
R11 B.n773 B.n772 585
R12 B.n774 B.n95 585
R13 B.n776 B.n775 585
R14 B.n777 B.n94 585
R15 B.n779 B.n778 585
R16 B.n780 B.n93 585
R17 B.n782 B.n781 585
R18 B.n783 B.n92 585
R19 B.n785 B.n784 585
R20 B.n786 B.n91 585
R21 B.n788 B.n787 585
R22 B.n789 B.n90 585
R23 B.n791 B.n790 585
R24 B.n792 B.n89 585
R25 B.n794 B.n793 585
R26 B.n795 B.n88 585
R27 B.n797 B.n796 585
R28 B.n798 B.n87 585
R29 B.n800 B.n799 585
R30 B.n801 B.n86 585
R31 B.n803 B.n802 585
R32 B.n804 B.n85 585
R33 B.n806 B.n805 585
R34 B.n807 B.n84 585
R35 B.n809 B.n808 585
R36 B.n810 B.n83 585
R37 B.n812 B.n811 585
R38 B.n813 B.n82 585
R39 B.n815 B.n814 585
R40 B.n816 B.n81 585
R41 B.n818 B.n817 585
R42 B.n819 B.n80 585
R43 B.n821 B.n820 585
R44 B.n822 B.n79 585
R45 B.n824 B.n823 585
R46 B.n825 B.n78 585
R47 B.n827 B.n826 585
R48 B.n828 B.n77 585
R49 B.n830 B.n829 585
R50 B.n831 B.n76 585
R51 B.n833 B.n832 585
R52 B.n834 B.n75 585
R53 B.n836 B.n835 585
R54 B.n837 B.n74 585
R55 B.n839 B.n838 585
R56 B.n840 B.n71 585
R57 B.n843 B.n842 585
R58 B.n844 B.n70 585
R59 B.n846 B.n845 585
R60 B.n847 B.n69 585
R61 B.n849 B.n848 585
R62 B.n850 B.n68 585
R63 B.n852 B.n851 585
R64 B.n853 B.n67 585
R65 B.n855 B.n854 585
R66 B.n857 B.n856 585
R67 B.n858 B.n63 585
R68 B.n860 B.n859 585
R69 B.n861 B.n62 585
R70 B.n863 B.n862 585
R71 B.n864 B.n61 585
R72 B.n866 B.n865 585
R73 B.n867 B.n60 585
R74 B.n869 B.n868 585
R75 B.n870 B.n59 585
R76 B.n872 B.n871 585
R77 B.n873 B.n58 585
R78 B.n875 B.n874 585
R79 B.n876 B.n57 585
R80 B.n878 B.n877 585
R81 B.n879 B.n56 585
R82 B.n881 B.n880 585
R83 B.n882 B.n55 585
R84 B.n884 B.n883 585
R85 B.n885 B.n54 585
R86 B.n887 B.n886 585
R87 B.n888 B.n53 585
R88 B.n890 B.n889 585
R89 B.n891 B.n52 585
R90 B.n893 B.n892 585
R91 B.n894 B.n51 585
R92 B.n896 B.n895 585
R93 B.n897 B.n50 585
R94 B.n899 B.n898 585
R95 B.n900 B.n49 585
R96 B.n902 B.n901 585
R97 B.n903 B.n48 585
R98 B.n905 B.n904 585
R99 B.n906 B.n47 585
R100 B.n908 B.n907 585
R101 B.n909 B.n46 585
R102 B.n911 B.n910 585
R103 B.n912 B.n45 585
R104 B.n914 B.n913 585
R105 B.n915 B.n44 585
R106 B.n917 B.n916 585
R107 B.n918 B.n43 585
R108 B.n920 B.n919 585
R109 B.n921 B.n42 585
R110 B.n923 B.n922 585
R111 B.n924 B.n41 585
R112 B.n926 B.n925 585
R113 B.n927 B.n40 585
R114 B.n929 B.n928 585
R115 B.n930 B.n39 585
R116 B.n932 B.n931 585
R117 B.n933 B.n38 585
R118 B.n935 B.n934 585
R119 B.n936 B.n37 585
R120 B.n938 B.n937 585
R121 B.n939 B.n36 585
R122 B.n941 B.n940 585
R123 B.n755 B.n754 585
R124 B.n753 B.n102 585
R125 B.n752 B.n751 585
R126 B.n750 B.n103 585
R127 B.n749 B.n748 585
R128 B.n747 B.n104 585
R129 B.n746 B.n745 585
R130 B.n744 B.n105 585
R131 B.n743 B.n742 585
R132 B.n741 B.n106 585
R133 B.n740 B.n739 585
R134 B.n738 B.n107 585
R135 B.n737 B.n736 585
R136 B.n735 B.n108 585
R137 B.n734 B.n733 585
R138 B.n732 B.n109 585
R139 B.n731 B.n730 585
R140 B.n729 B.n110 585
R141 B.n728 B.n727 585
R142 B.n726 B.n111 585
R143 B.n725 B.n724 585
R144 B.n723 B.n112 585
R145 B.n722 B.n721 585
R146 B.n720 B.n113 585
R147 B.n719 B.n718 585
R148 B.n717 B.n114 585
R149 B.n716 B.n715 585
R150 B.n714 B.n115 585
R151 B.n713 B.n712 585
R152 B.n711 B.n116 585
R153 B.n710 B.n709 585
R154 B.n708 B.n117 585
R155 B.n707 B.n706 585
R156 B.n705 B.n118 585
R157 B.n704 B.n703 585
R158 B.n702 B.n119 585
R159 B.n701 B.n700 585
R160 B.n699 B.n120 585
R161 B.n698 B.n697 585
R162 B.n696 B.n121 585
R163 B.n695 B.n694 585
R164 B.n693 B.n122 585
R165 B.n692 B.n691 585
R166 B.n690 B.n123 585
R167 B.n689 B.n688 585
R168 B.n687 B.n124 585
R169 B.n686 B.n685 585
R170 B.n684 B.n125 585
R171 B.n683 B.n682 585
R172 B.n681 B.n126 585
R173 B.n680 B.n679 585
R174 B.n678 B.n127 585
R175 B.n677 B.n676 585
R176 B.n675 B.n128 585
R177 B.n674 B.n673 585
R178 B.n672 B.n129 585
R179 B.n671 B.n670 585
R180 B.n669 B.n130 585
R181 B.n668 B.n667 585
R182 B.n666 B.n131 585
R183 B.n665 B.n664 585
R184 B.n663 B.n132 585
R185 B.n662 B.n661 585
R186 B.n660 B.n133 585
R187 B.n659 B.n658 585
R188 B.n657 B.n134 585
R189 B.n656 B.n655 585
R190 B.n654 B.n135 585
R191 B.n653 B.n652 585
R192 B.n651 B.n136 585
R193 B.n650 B.n649 585
R194 B.n648 B.n137 585
R195 B.n647 B.n646 585
R196 B.n645 B.n138 585
R197 B.n644 B.n643 585
R198 B.n642 B.n139 585
R199 B.n641 B.n640 585
R200 B.n639 B.n140 585
R201 B.n638 B.n637 585
R202 B.n636 B.n141 585
R203 B.n635 B.n634 585
R204 B.n633 B.n142 585
R205 B.n632 B.n631 585
R206 B.n630 B.n143 585
R207 B.n629 B.n628 585
R208 B.n627 B.n144 585
R209 B.n626 B.n625 585
R210 B.n624 B.n145 585
R211 B.n623 B.n622 585
R212 B.n621 B.n146 585
R213 B.n620 B.n619 585
R214 B.n618 B.n147 585
R215 B.n617 B.n616 585
R216 B.n615 B.n148 585
R217 B.n614 B.n613 585
R218 B.n612 B.n149 585
R219 B.n611 B.n610 585
R220 B.n609 B.n150 585
R221 B.n608 B.n607 585
R222 B.n606 B.n151 585
R223 B.n605 B.n604 585
R224 B.n603 B.n152 585
R225 B.n602 B.n601 585
R226 B.n600 B.n153 585
R227 B.n599 B.n598 585
R228 B.n597 B.n154 585
R229 B.n596 B.n595 585
R230 B.n594 B.n155 585
R231 B.n593 B.n592 585
R232 B.n591 B.n156 585
R233 B.n590 B.n589 585
R234 B.n588 B.n157 585
R235 B.n587 B.n586 585
R236 B.n585 B.n158 585
R237 B.n584 B.n583 585
R238 B.n582 B.n159 585
R239 B.n581 B.n580 585
R240 B.n579 B.n160 585
R241 B.n578 B.n577 585
R242 B.n576 B.n161 585
R243 B.n575 B.n574 585
R244 B.n573 B.n162 585
R245 B.n572 B.n571 585
R246 B.n570 B.n163 585
R247 B.n569 B.n568 585
R248 B.n567 B.n164 585
R249 B.n566 B.n565 585
R250 B.n564 B.n165 585
R251 B.n563 B.n562 585
R252 B.n561 B.n166 585
R253 B.n560 B.n559 585
R254 B.n558 B.n167 585
R255 B.n557 B.n556 585
R256 B.n555 B.n168 585
R257 B.n554 B.n553 585
R258 B.n368 B.n367 585
R259 B.n369 B.n234 585
R260 B.n371 B.n370 585
R261 B.n372 B.n233 585
R262 B.n374 B.n373 585
R263 B.n375 B.n232 585
R264 B.n377 B.n376 585
R265 B.n378 B.n231 585
R266 B.n380 B.n379 585
R267 B.n381 B.n230 585
R268 B.n383 B.n382 585
R269 B.n384 B.n229 585
R270 B.n386 B.n385 585
R271 B.n387 B.n228 585
R272 B.n389 B.n388 585
R273 B.n390 B.n227 585
R274 B.n392 B.n391 585
R275 B.n393 B.n226 585
R276 B.n395 B.n394 585
R277 B.n396 B.n225 585
R278 B.n398 B.n397 585
R279 B.n399 B.n224 585
R280 B.n401 B.n400 585
R281 B.n402 B.n223 585
R282 B.n404 B.n403 585
R283 B.n405 B.n222 585
R284 B.n407 B.n406 585
R285 B.n408 B.n221 585
R286 B.n410 B.n409 585
R287 B.n411 B.n220 585
R288 B.n413 B.n412 585
R289 B.n414 B.n219 585
R290 B.n416 B.n415 585
R291 B.n417 B.n218 585
R292 B.n419 B.n418 585
R293 B.n420 B.n217 585
R294 B.n422 B.n421 585
R295 B.n423 B.n216 585
R296 B.n425 B.n424 585
R297 B.n426 B.n215 585
R298 B.n428 B.n427 585
R299 B.n429 B.n214 585
R300 B.n431 B.n430 585
R301 B.n432 B.n213 585
R302 B.n434 B.n433 585
R303 B.n435 B.n212 585
R304 B.n437 B.n436 585
R305 B.n438 B.n211 585
R306 B.n440 B.n439 585
R307 B.n441 B.n210 585
R308 B.n443 B.n442 585
R309 B.n444 B.n209 585
R310 B.n446 B.n445 585
R311 B.n447 B.n208 585
R312 B.n449 B.n448 585
R313 B.n450 B.n207 585
R314 B.n452 B.n451 585
R315 B.n454 B.n453 585
R316 B.n455 B.n203 585
R317 B.n457 B.n456 585
R318 B.n458 B.n202 585
R319 B.n460 B.n459 585
R320 B.n461 B.n201 585
R321 B.n463 B.n462 585
R322 B.n464 B.n200 585
R323 B.n466 B.n465 585
R324 B.n468 B.n197 585
R325 B.n470 B.n469 585
R326 B.n471 B.n196 585
R327 B.n473 B.n472 585
R328 B.n474 B.n195 585
R329 B.n476 B.n475 585
R330 B.n477 B.n194 585
R331 B.n479 B.n478 585
R332 B.n480 B.n193 585
R333 B.n482 B.n481 585
R334 B.n483 B.n192 585
R335 B.n485 B.n484 585
R336 B.n486 B.n191 585
R337 B.n488 B.n487 585
R338 B.n489 B.n190 585
R339 B.n491 B.n490 585
R340 B.n492 B.n189 585
R341 B.n494 B.n493 585
R342 B.n495 B.n188 585
R343 B.n497 B.n496 585
R344 B.n498 B.n187 585
R345 B.n500 B.n499 585
R346 B.n501 B.n186 585
R347 B.n503 B.n502 585
R348 B.n504 B.n185 585
R349 B.n506 B.n505 585
R350 B.n507 B.n184 585
R351 B.n509 B.n508 585
R352 B.n510 B.n183 585
R353 B.n512 B.n511 585
R354 B.n513 B.n182 585
R355 B.n515 B.n514 585
R356 B.n516 B.n181 585
R357 B.n518 B.n517 585
R358 B.n519 B.n180 585
R359 B.n521 B.n520 585
R360 B.n522 B.n179 585
R361 B.n524 B.n523 585
R362 B.n525 B.n178 585
R363 B.n527 B.n526 585
R364 B.n528 B.n177 585
R365 B.n530 B.n529 585
R366 B.n531 B.n176 585
R367 B.n533 B.n532 585
R368 B.n534 B.n175 585
R369 B.n536 B.n535 585
R370 B.n537 B.n174 585
R371 B.n539 B.n538 585
R372 B.n540 B.n173 585
R373 B.n542 B.n541 585
R374 B.n543 B.n172 585
R375 B.n545 B.n544 585
R376 B.n546 B.n171 585
R377 B.n548 B.n547 585
R378 B.n549 B.n170 585
R379 B.n551 B.n550 585
R380 B.n552 B.n169 585
R381 B.n366 B.n235 585
R382 B.n365 B.n364 585
R383 B.n363 B.n236 585
R384 B.n362 B.n361 585
R385 B.n360 B.n237 585
R386 B.n359 B.n358 585
R387 B.n357 B.n238 585
R388 B.n356 B.n355 585
R389 B.n354 B.n239 585
R390 B.n353 B.n352 585
R391 B.n351 B.n240 585
R392 B.n350 B.n349 585
R393 B.n348 B.n241 585
R394 B.n347 B.n346 585
R395 B.n345 B.n242 585
R396 B.n344 B.n343 585
R397 B.n342 B.n243 585
R398 B.n341 B.n340 585
R399 B.n339 B.n244 585
R400 B.n338 B.n337 585
R401 B.n336 B.n245 585
R402 B.n335 B.n334 585
R403 B.n333 B.n246 585
R404 B.n332 B.n331 585
R405 B.n330 B.n247 585
R406 B.n329 B.n328 585
R407 B.n327 B.n248 585
R408 B.n326 B.n325 585
R409 B.n324 B.n249 585
R410 B.n323 B.n322 585
R411 B.n321 B.n250 585
R412 B.n320 B.n319 585
R413 B.n318 B.n251 585
R414 B.n317 B.n316 585
R415 B.n315 B.n252 585
R416 B.n314 B.n313 585
R417 B.n312 B.n253 585
R418 B.n311 B.n310 585
R419 B.n309 B.n254 585
R420 B.n308 B.n307 585
R421 B.n306 B.n255 585
R422 B.n305 B.n304 585
R423 B.n303 B.n256 585
R424 B.n302 B.n301 585
R425 B.n300 B.n257 585
R426 B.n299 B.n298 585
R427 B.n297 B.n258 585
R428 B.n296 B.n295 585
R429 B.n294 B.n259 585
R430 B.n293 B.n292 585
R431 B.n291 B.n260 585
R432 B.n290 B.n289 585
R433 B.n288 B.n261 585
R434 B.n287 B.n286 585
R435 B.n285 B.n262 585
R436 B.n284 B.n283 585
R437 B.n282 B.n263 585
R438 B.n281 B.n280 585
R439 B.n279 B.n264 585
R440 B.n278 B.n277 585
R441 B.n276 B.n265 585
R442 B.n275 B.n274 585
R443 B.n273 B.n266 585
R444 B.n272 B.n271 585
R445 B.n270 B.n267 585
R446 B.n269 B.n268 585
R447 B.n2 B.n0 585
R448 B.n1041 B.n1 585
R449 B.n1040 B.n1039 585
R450 B.n1038 B.n3 585
R451 B.n1037 B.n1036 585
R452 B.n1035 B.n4 585
R453 B.n1034 B.n1033 585
R454 B.n1032 B.n5 585
R455 B.n1031 B.n1030 585
R456 B.n1029 B.n6 585
R457 B.n1028 B.n1027 585
R458 B.n1026 B.n7 585
R459 B.n1025 B.n1024 585
R460 B.n1023 B.n8 585
R461 B.n1022 B.n1021 585
R462 B.n1020 B.n9 585
R463 B.n1019 B.n1018 585
R464 B.n1017 B.n10 585
R465 B.n1016 B.n1015 585
R466 B.n1014 B.n11 585
R467 B.n1013 B.n1012 585
R468 B.n1011 B.n12 585
R469 B.n1010 B.n1009 585
R470 B.n1008 B.n13 585
R471 B.n1007 B.n1006 585
R472 B.n1005 B.n14 585
R473 B.n1004 B.n1003 585
R474 B.n1002 B.n15 585
R475 B.n1001 B.n1000 585
R476 B.n999 B.n16 585
R477 B.n998 B.n997 585
R478 B.n996 B.n17 585
R479 B.n995 B.n994 585
R480 B.n993 B.n18 585
R481 B.n992 B.n991 585
R482 B.n990 B.n19 585
R483 B.n989 B.n988 585
R484 B.n987 B.n20 585
R485 B.n986 B.n985 585
R486 B.n984 B.n21 585
R487 B.n983 B.n982 585
R488 B.n981 B.n22 585
R489 B.n980 B.n979 585
R490 B.n978 B.n23 585
R491 B.n977 B.n976 585
R492 B.n975 B.n24 585
R493 B.n974 B.n973 585
R494 B.n972 B.n25 585
R495 B.n971 B.n970 585
R496 B.n969 B.n26 585
R497 B.n968 B.n967 585
R498 B.n966 B.n27 585
R499 B.n965 B.n964 585
R500 B.n963 B.n28 585
R501 B.n962 B.n961 585
R502 B.n960 B.n29 585
R503 B.n959 B.n958 585
R504 B.n957 B.n30 585
R505 B.n956 B.n955 585
R506 B.n954 B.n31 585
R507 B.n953 B.n952 585
R508 B.n951 B.n32 585
R509 B.n950 B.n949 585
R510 B.n948 B.n33 585
R511 B.n947 B.n946 585
R512 B.n945 B.n34 585
R513 B.n944 B.n943 585
R514 B.n942 B.n35 585
R515 B.n1043 B.n1042 585
R516 B.n368 B.n235 463.671
R517 B.n940 B.n35 463.671
R518 B.n554 B.n169 463.671
R519 B.n754 B.n101 463.671
R520 B.n198 B.t9 321.401
R521 B.n204 B.t0 321.401
R522 B.n64 B.t6 321.401
R523 B.n72 B.t3 321.401
R524 B.n198 B.t11 185.428
R525 B.n72 B.t4 185.428
R526 B.n204 B.t2 185.405
R527 B.n64 B.t7 185.405
R528 B.n364 B.n235 163.367
R529 B.n364 B.n363 163.367
R530 B.n363 B.n362 163.367
R531 B.n362 B.n237 163.367
R532 B.n358 B.n237 163.367
R533 B.n358 B.n357 163.367
R534 B.n357 B.n356 163.367
R535 B.n356 B.n239 163.367
R536 B.n352 B.n239 163.367
R537 B.n352 B.n351 163.367
R538 B.n351 B.n350 163.367
R539 B.n350 B.n241 163.367
R540 B.n346 B.n241 163.367
R541 B.n346 B.n345 163.367
R542 B.n345 B.n344 163.367
R543 B.n344 B.n243 163.367
R544 B.n340 B.n243 163.367
R545 B.n340 B.n339 163.367
R546 B.n339 B.n338 163.367
R547 B.n338 B.n245 163.367
R548 B.n334 B.n245 163.367
R549 B.n334 B.n333 163.367
R550 B.n333 B.n332 163.367
R551 B.n332 B.n247 163.367
R552 B.n328 B.n247 163.367
R553 B.n328 B.n327 163.367
R554 B.n327 B.n326 163.367
R555 B.n326 B.n249 163.367
R556 B.n322 B.n249 163.367
R557 B.n322 B.n321 163.367
R558 B.n321 B.n320 163.367
R559 B.n320 B.n251 163.367
R560 B.n316 B.n251 163.367
R561 B.n316 B.n315 163.367
R562 B.n315 B.n314 163.367
R563 B.n314 B.n253 163.367
R564 B.n310 B.n253 163.367
R565 B.n310 B.n309 163.367
R566 B.n309 B.n308 163.367
R567 B.n308 B.n255 163.367
R568 B.n304 B.n255 163.367
R569 B.n304 B.n303 163.367
R570 B.n303 B.n302 163.367
R571 B.n302 B.n257 163.367
R572 B.n298 B.n257 163.367
R573 B.n298 B.n297 163.367
R574 B.n297 B.n296 163.367
R575 B.n296 B.n259 163.367
R576 B.n292 B.n259 163.367
R577 B.n292 B.n291 163.367
R578 B.n291 B.n290 163.367
R579 B.n290 B.n261 163.367
R580 B.n286 B.n261 163.367
R581 B.n286 B.n285 163.367
R582 B.n285 B.n284 163.367
R583 B.n284 B.n263 163.367
R584 B.n280 B.n263 163.367
R585 B.n280 B.n279 163.367
R586 B.n279 B.n278 163.367
R587 B.n278 B.n265 163.367
R588 B.n274 B.n265 163.367
R589 B.n274 B.n273 163.367
R590 B.n273 B.n272 163.367
R591 B.n272 B.n267 163.367
R592 B.n268 B.n267 163.367
R593 B.n268 B.n2 163.367
R594 B.n1042 B.n2 163.367
R595 B.n1042 B.n1041 163.367
R596 B.n1041 B.n1040 163.367
R597 B.n1040 B.n3 163.367
R598 B.n1036 B.n3 163.367
R599 B.n1036 B.n1035 163.367
R600 B.n1035 B.n1034 163.367
R601 B.n1034 B.n5 163.367
R602 B.n1030 B.n5 163.367
R603 B.n1030 B.n1029 163.367
R604 B.n1029 B.n1028 163.367
R605 B.n1028 B.n7 163.367
R606 B.n1024 B.n7 163.367
R607 B.n1024 B.n1023 163.367
R608 B.n1023 B.n1022 163.367
R609 B.n1022 B.n9 163.367
R610 B.n1018 B.n9 163.367
R611 B.n1018 B.n1017 163.367
R612 B.n1017 B.n1016 163.367
R613 B.n1016 B.n11 163.367
R614 B.n1012 B.n11 163.367
R615 B.n1012 B.n1011 163.367
R616 B.n1011 B.n1010 163.367
R617 B.n1010 B.n13 163.367
R618 B.n1006 B.n13 163.367
R619 B.n1006 B.n1005 163.367
R620 B.n1005 B.n1004 163.367
R621 B.n1004 B.n15 163.367
R622 B.n1000 B.n15 163.367
R623 B.n1000 B.n999 163.367
R624 B.n999 B.n998 163.367
R625 B.n998 B.n17 163.367
R626 B.n994 B.n17 163.367
R627 B.n994 B.n993 163.367
R628 B.n993 B.n992 163.367
R629 B.n992 B.n19 163.367
R630 B.n988 B.n19 163.367
R631 B.n988 B.n987 163.367
R632 B.n987 B.n986 163.367
R633 B.n986 B.n21 163.367
R634 B.n982 B.n21 163.367
R635 B.n982 B.n981 163.367
R636 B.n981 B.n980 163.367
R637 B.n980 B.n23 163.367
R638 B.n976 B.n23 163.367
R639 B.n976 B.n975 163.367
R640 B.n975 B.n974 163.367
R641 B.n974 B.n25 163.367
R642 B.n970 B.n25 163.367
R643 B.n970 B.n969 163.367
R644 B.n969 B.n968 163.367
R645 B.n968 B.n27 163.367
R646 B.n964 B.n27 163.367
R647 B.n964 B.n963 163.367
R648 B.n963 B.n962 163.367
R649 B.n962 B.n29 163.367
R650 B.n958 B.n29 163.367
R651 B.n958 B.n957 163.367
R652 B.n957 B.n956 163.367
R653 B.n956 B.n31 163.367
R654 B.n952 B.n31 163.367
R655 B.n952 B.n951 163.367
R656 B.n951 B.n950 163.367
R657 B.n950 B.n33 163.367
R658 B.n946 B.n33 163.367
R659 B.n946 B.n945 163.367
R660 B.n945 B.n944 163.367
R661 B.n944 B.n35 163.367
R662 B.n369 B.n368 163.367
R663 B.n370 B.n369 163.367
R664 B.n370 B.n233 163.367
R665 B.n374 B.n233 163.367
R666 B.n375 B.n374 163.367
R667 B.n376 B.n375 163.367
R668 B.n376 B.n231 163.367
R669 B.n380 B.n231 163.367
R670 B.n381 B.n380 163.367
R671 B.n382 B.n381 163.367
R672 B.n382 B.n229 163.367
R673 B.n386 B.n229 163.367
R674 B.n387 B.n386 163.367
R675 B.n388 B.n387 163.367
R676 B.n388 B.n227 163.367
R677 B.n392 B.n227 163.367
R678 B.n393 B.n392 163.367
R679 B.n394 B.n393 163.367
R680 B.n394 B.n225 163.367
R681 B.n398 B.n225 163.367
R682 B.n399 B.n398 163.367
R683 B.n400 B.n399 163.367
R684 B.n400 B.n223 163.367
R685 B.n404 B.n223 163.367
R686 B.n405 B.n404 163.367
R687 B.n406 B.n405 163.367
R688 B.n406 B.n221 163.367
R689 B.n410 B.n221 163.367
R690 B.n411 B.n410 163.367
R691 B.n412 B.n411 163.367
R692 B.n412 B.n219 163.367
R693 B.n416 B.n219 163.367
R694 B.n417 B.n416 163.367
R695 B.n418 B.n417 163.367
R696 B.n418 B.n217 163.367
R697 B.n422 B.n217 163.367
R698 B.n423 B.n422 163.367
R699 B.n424 B.n423 163.367
R700 B.n424 B.n215 163.367
R701 B.n428 B.n215 163.367
R702 B.n429 B.n428 163.367
R703 B.n430 B.n429 163.367
R704 B.n430 B.n213 163.367
R705 B.n434 B.n213 163.367
R706 B.n435 B.n434 163.367
R707 B.n436 B.n435 163.367
R708 B.n436 B.n211 163.367
R709 B.n440 B.n211 163.367
R710 B.n441 B.n440 163.367
R711 B.n442 B.n441 163.367
R712 B.n442 B.n209 163.367
R713 B.n446 B.n209 163.367
R714 B.n447 B.n446 163.367
R715 B.n448 B.n447 163.367
R716 B.n448 B.n207 163.367
R717 B.n452 B.n207 163.367
R718 B.n453 B.n452 163.367
R719 B.n453 B.n203 163.367
R720 B.n457 B.n203 163.367
R721 B.n458 B.n457 163.367
R722 B.n459 B.n458 163.367
R723 B.n459 B.n201 163.367
R724 B.n463 B.n201 163.367
R725 B.n464 B.n463 163.367
R726 B.n465 B.n464 163.367
R727 B.n465 B.n197 163.367
R728 B.n470 B.n197 163.367
R729 B.n471 B.n470 163.367
R730 B.n472 B.n471 163.367
R731 B.n472 B.n195 163.367
R732 B.n476 B.n195 163.367
R733 B.n477 B.n476 163.367
R734 B.n478 B.n477 163.367
R735 B.n478 B.n193 163.367
R736 B.n482 B.n193 163.367
R737 B.n483 B.n482 163.367
R738 B.n484 B.n483 163.367
R739 B.n484 B.n191 163.367
R740 B.n488 B.n191 163.367
R741 B.n489 B.n488 163.367
R742 B.n490 B.n489 163.367
R743 B.n490 B.n189 163.367
R744 B.n494 B.n189 163.367
R745 B.n495 B.n494 163.367
R746 B.n496 B.n495 163.367
R747 B.n496 B.n187 163.367
R748 B.n500 B.n187 163.367
R749 B.n501 B.n500 163.367
R750 B.n502 B.n501 163.367
R751 B.n502 B.n185 163.367
R752 B.n506 B.n185 163.367
R753 B.n507 B.n506 163.367
R754 B.n508 B.n507 163.367
R755 B.n508 B.n183 163.367
R756 B.n512 B.n183 163.367
R757 B.n513 B.n512 163.367
R758 B.n514 B.n513 163.367
R759 B.n514 B.n181 163.367
R760 B.n518 B.n181 163.367
R761 B.n519 B.n518 163.367
R762 B.n520 B.n519 163.367
R763 B.n520 B.n179 163.367
R764 B.n524 B.n179 163.367
R765 B.n525 B.n524 163.367
R766 B.n526 B.n525 163.367
R767 B.n526 B.n177 163.367
R768 B.n530 B.n177 163.367
R769 B.n531 B.n530 163.367
R770 B.n532 B.n531 163.367
R771 B.n532 B.n175 163.367
R772 B.n536 B.n175 163.367
R773 B.n537 B.n536 163.367
R774 B.n538 B.n537 163.367
R775 B.n538 B.n173 163.367
R776 B.n542 B.n173 163.367
R777 B.n543 B.n542 163.367
R778 B.n544 B.n543 163.367
R779 B.n544 B.n171 163.367
R780 B.n548 B.n171 163.367
R781 B.n549 B.n548 163.367
R782 B.n550 B.n549 163.367
R783 B.n550 B.n169 163.367
R784 B.n555 B.n554 163.367
R785 B.n556 B.n555 163.367
R786 B.n556 B.n167 163.367
R787 B.n560 B.n167 163.367
R788 B.n561 B.n560 163.367
R789 B.n562 B.n561 163.367
R790 B.n562 B.n165 163.367
R791 B.n566 B.n165 163.367
R792 B.n567 B.n566 163.367
R793 B.n568 B.n567 163.367
R794 B.n568 B.n163 163.367
R795 B.n572 B.n163 163.367
R796 B.n573 B.n572 163.367
R797 B.n574 B.n573 163.367
R798 B.n574 B.n161 163.367
R799 B.n578 B.n161 163.367
R800 B.n579 B.n578 163.367
R801 B.n580 B.n579 163.367
R802 B.n580 B.n159 163.367
R803 B.n584 B.n159 163.367
R804 B.n585 B.n584 163.367
R805 B.n586 B.n585 163.367
R806 B.n586 B.n157 163.367
R807 B.n590 B.n157 163.367
R808 B.n591 B.n590 163.367
R809 B.n592 B.n591 163.367
R810 B.n592 B.n155 163.367
R811 B.n596 B.n155 163.367
R812 B.n597 B.n596 163.367
R813 B.n598 B.n597 163.367
R814 B.n598 B.n153 163.367
R815 B.n602 B.n153 163.367
R816 B.n603 B.n602 163.367
R817 B.n604 B.n603 163.367
R818 B.n604 B.n151 163.367
R819 B.n608 B.n151 163.367
R820 B.n609 B.n608 163.367
R821 B.n610 B.n609 163.367
R822 B.n610 B.n149 163.367
R823 B.n614 B.n149 163.367
R824 B.n615 B.n614 163.367
R825 B.n616 B.n615 163.367
R826 B.n616 B.n147 163.367
R827 B.n620 B.n147 163.367
R828 B.n621 B.n620 163.367
R829 B.n622 B.n621 163.367
R830 B.n622 B.n145 163.367
R831 B.n626 B.n145 163.367
R832 B.n627 B.n626 163.367
R833 B.n628 B.n627 163.367
R834 B.n628 B.n143 163.367
R835 B.n632 B.n143 163.367
R836 B.n633 B.n632 163.367
R837 B.n634 B.n633 163.367
R838 B.n634 B.n141 163.367
R839 B.n638 B.n141 163.367
R840 B.n639 B.n638 163.367
R841 B.n640 B.n639 163.367
R842 B.n640 B.n139 163.367
R843 B.n644 B.n139 163.367
R844 B.n645 B.n644 163.367
R845 B.n646 B.n645 163.367
R846 B.n646 B.n137 163.367
R847 B.n650 B.n137 163.367
R848 B.n651 B.n650 163.367
R849 B.n652 B.n651 163.367
R850 B.n652 B.n135 163.367
R851 B.n656 B.n135 163.367
R852 B.n657 B.n656 163.367
R853 B.n658 B.n657 163.367
R854 B.n658 B.n133 163.367
R855 B.n662 B.n133 163.367
R856 B.n663 B.n662 163.367
R857 B.n664 B.n663 163.367
R858 B.n664 B.n131 163.367
R859 B.n668 B.n131 163.367
R860 B.n669 B.n668 163.367
R861 B.n670 B.n669 163.367
R862 B.n670 B.n129 163.367
R863 B.n674 B.n129 163.367
R864 B.n675 B.n674 163.367
R865 B.n676 B.n675 163.367
R866 B.n676 B.n127 163.367
R867 B.n680 B.n127 163.367
R868 B.n681 B.n680 163.367
R869 B.n682 B.n681 163.367
R870 B.n682 B.n125 163.367
R871 B.n686 B.n125 163.367
R872 B.n687 B.n686 163.367
R873 B.n688 B.n687 163.367
R874 B.n688 B.n123 163.367
R875 B.n692 B.n123 163.367
R876 B.n693 B.n692 163.367
R877 B.n694 B.n693 163.367
R878 B.n694 B.n121 163.367
R879 B.n698 B.n121 163.367
R880 B.n699 B.n698 163.367
R881 B.n700 B.n699 163.367
R882 B.n700 B.n119 163.367
R883 B.n704 B.n119 163.367
R884 B.n705 B.n704 163.367
R885 B.n706 B.n705 163.367
R886 B.n706 B.n117 163.367
R887 B.n710 B.n117 163.367
R888 B.n711 B.n710 163.367
R889 B.n712 B.n711 163.367
R890 B.n712 B.n115 163.367
R891 B.n716 B.n115 163.367
R892 B.n717 B.n716 163.367
R893 B.n718 B.n717 163.367
R894 B.n718 B.n113 163.367
R895 B.n722 B.n113 163.367
R896 B.n723 B.n722 163.367
R897 B.n724 B.n723 163.367
R898 B.n724 B.n111 163.367
R899 B.n728 B.n111 163.367
R900 B.n729 B.n728 163.367
R901 B.n730 B.n729 163.367
R902 B.n730 B.n109 163.367
R903 B.n734 B.n109 163.367
R904 B.n735 B.n734 163.367
R905 B.n736 B.n735 163.367
R906 B.n736 B.n107 163.367
R907 B.n740 B.n107 163.367
R908 B.n741 B.n740 163.367
R909 B.n742 B.n741 163.367
R910 B.n742 B.n105 163.367
R911 B.n746 B.n105 163.367
R912 B.n747 B.n746 163.367
R913 B.n748 B.n747 163.367
R914 B.n748 B.n103 163.367
R915 B.n752 B.n103 163.367
R916 B.n753 B.n752 163.367
R917 B.n754 B.n753 163.367
R918 B.n940 B.n939 163.367
R919 B.n939 B.n938 163.367
R920 B.n938 B.n37 163.367
R921 B.n934 B.n37 163.367
R922 B.n934 B.n933 163.367
R923 B.n933 B.n932 163.367
R924 B.n932 B.n39 163.367
R925 B.n928 B.n39 163.367
R926 B.n928 B.n927 163.367
R927 B.n927 B.n926 163.367
R928 B.n926 B.n41 163.367
R929 B.n922 B.n41 163.367
R930 B.n922 B.n921 163.367
R931 B.n921 B.n920 163.367
R932 B.n920 B.n43 163.367
R933 B.n916 B.n43 163.367
R934 B.n916 B.n915 163.367
R935 B.n915 B.n914 163.367
R936 B.n914 B.n45 163.367
R937 B.n910 B.n45 163.367
R938 B.n910 B.n909 163.367
R939 B.n909 B.n908 163.367
R940 B.n908 B.n47 163.367
R941 B.n904 B.n47 163.367
R942 B.n904 B.n903 163.367
R943 B.n903 B.n902 163.367
R944 B.n902 B.n49 163.367
R945 B.n898 B.n49 163.367
R946 B.n898 B.n897 163.367
R947 B.n897 B.n896 163.367
R948 B.n896 B.n51 163.367
R949 B.n892 B.n51 163.367
R950 B.n892 B.n891 163.367
R951 B.n891 B.n890 163.367
R952 B.n890 B.n53 163.367
R953 B.n886 B.n53 163.367
R954 B.n886 B.n885 163.367
R955 B.n885 B.n884 163.367
R956 B.n884 B.n55 163.367
R957 B.n880 B.n55 163.367
R958 B.n880 B.n879 163.367
R959 B.n879 B.n878 163.367
R960 B.n878 B.n57 163.367
R961 B.n874 B.n57 163.367
R962 B.n874 B.n873 163.367
R963 B.n873 B.n872 163.367
R964 B.n872 B.n59 163.367
R965 B.n868 B.n59 163.367
R966 B.n868 B.n867 163.367
R967 B.n867 B.n866 163.367
R968 B.n866 B.n61 163.367
R969 B.n862 B.n61 163.367
R970 B.n862 B.n861 163.367
R971 B.n861 B.n860 163.367
R972 B.n860 B.n63 163.367
R973 B.n856 B.n63 163.367
R974 B.n856 B.n855 163.367
R975 B.n855 B.n67 163.367
R976 B.n851 B.n67 163.367
R977 B.n851 B.n850 163.367
R978 B.n850 B.n849 163.367
R979 B.n849 B.n69 163.367
R980 B.n845 B.n69 163.367
R981 B.n845 B.n844 163.367
R982 B.n844 B.n843 163.367
R983 B.n843 B.n71 163.367
R984 B.n838 B.n71 163.367
R985 B.n838 B.n837 163.367
R986 B.n837 B.n836 163.367
R987 B.n836 B.n75 163.367
R988 B.n832 B.n75 163.367
R989 B.n832 B.n831 163.367
R990 B.n831 B.n830 163.367
R991 B.n830 B.n77 163.367
R992 B.n826 B.n77 163.367
R993 B.n826 B.n825 163.367
R994 B.n825 B.n824 163.367
R995 B.n824 B.n79 163.367
R996 B.n820 B.n79 163.367
R997 B.n820 B.n819 163.367
R998 B.n819 B.n818 163.367
R999 B.n818 B.n81 163.367
R1000 B.n814 B.n81 163.367
R1001 B.n814 B.n813 163.367
R1002 B.n813 B.n812 163.367
R1003 B.n812 B.n83 163.367
R1004 B.n808 B.n83 163.367
R1005 B.n808 B.n807 163.367
R1006 B.n807 B.n806 163.367
R1007 B.n806 B.n85 163.367
R1008 B.n802 B.n85 163.367
R1009 B.n802 B.n801 163.367
R1010 B.n801 B.n800 163.367
R1011 B.n800 B.n87 163.367
R1012 B.n796 B.n87 163.367
R1013 B.n796 B.n795 163.367
R1014 B.n795 B.n794 163.367
R1015 B.n794 B.n89 163.367
R1016 B.n790 B.n89 163.367
R1017 B.n790 B.n789 163.367
R1018 B.n789 B.n788 163.367
R1019 B.n788 B.n91 163.367
R1020 B.n784 B.n91 163.367
R1021 B.n784 B.n783 163.367
R1022 B.n783 B.n782 163.367
R1023 B.n782 B.n93 163.367
R1024 B.n778 B.n93 163.367
R1025 B.n778 B.n777 163.367
R1026 B.n777 B.n776 163.367
R1027 B.n776 B.n95 163.367
R1028 B.n772 B.n95 163.367
R1029 B.n772 B.n771 163.367
R1030 B.n771 B.n770 163.367
R1031 B.n770 B.n97 163.367
R1032 B.n766 B.n97 163.367
R1033 B.n766 B.n765 163.367
R1034 B.n765 B.n764 163.367
R1035 B.n764 B.n99 163.367
R1036 B.n760 B.n99 163.367
R1037 B.n760 B.n759 163.367
R1038 B.n759 B.n758 163.367
R1039 B.n758 B.n101 163.367
R1040 B.n199 B.t10 107.852
R1041 B.n73 B.t5 107.852
R1042 B.n205 B.t1 107.829
R1043 B.n65 B.t8 107.829
R1044 B.n199 B.n198 77.5763
R1045 B.n205 B.n204 77.5763
R1046 B.n65 B.n64 77.5763
R1047 B.n73 B.n72 77.5763
R1048 B.n467 B.n199 59.5399
R1049 B.n206 B.n205 59.5399
R1050 B.n66 B.n65 59.5399
R1051 B.n841 B.n73 59.5399
R1052 B.n942 B.n941 30.1273
R1053 B.n756 B.n755 30.1273
R1054 B.n553 B.n552 30.1273
R1055 B.n367 B.n366 30.1273
R1056 B B.n1043 18.0485
R1057 B.n941 B.n36 10.6151
R1058 B.n937 B.n36 10.6151
R1059 B.n937 B.n936 10.6151
R1060 B.n936 B.n935 10.6151
R1061 B.n935 B.n38 10.6151
R1062 B.n931 B.n38 10.6151
R1063 B.n931 B.n930 10.6151
R1064 B.n930 B.n929 10.6151
R1065 B.n929 B.n40 10.6151
R1066 B.n925 B.n40 10.6151
R1067 B.n925 B.n924 10.6151
R1068 B.n924 B.n923 10.6151
R1069 B.n923 B.n42 10.6151
R1070 B.n919 B.n42 10.6151
R1071 B.n919 B.n918 10.6151
R1072 B.n918 B.n917 10.6151
R1073 B.n917 B.n44 10.6151
R1074 B.n913 B.n44 10.6151
R1075 B.n913 B.n912 10.6151
R1076 B.n912 B.n911 10.6151
R1077 B.n911 B.n46 10.6151
R1078 B.n907 B.n46 10.6151
R1079 B.n907 B.n906 10.6151
R1080 B.n906 B.n905 10.6151
R1081 B.n905 B.n48 10.6151
R1082 B.n901 B.n48 10.6151
R1083 B.n901 B.n900 10.6151
R1084 B.n900 B.n899 10.6151
R1085 B.n899 B.n50 10.6151
R1086 B.n895 B.n50 10.6151
R1087 B.n895 B.n894 10.6151
R1088 B.n894 B.n893 10.6151
R1089 B.n893 B.n52 10.6151
R1090 B.n889 B.n52 10.6151
R1091 B.n889 B.n888 10.6151
R1092 B.n888 B.n887 10.6151
R1093 B.n887 B.n54 10.6151
R1094 B.n883 B.n54 10.6151
R1095 B.n883 B.n882 10.6151
R1096 B.n882 B.n881 10.6151
R1097 B.n881 B.n56 10.6151
R1098 B.n877 B.n56 10.6151
R1099 B.n877 B.n876 10.6151
R1100 B.n876 B.n875 10.6151
R1101 B.n875 B.n58 10.6151
R1102 B.n871 B.n58 10.6151
R1103 B.n871 B.n870 10.6151
R1104 B.n870 B.n869 10.6151
R1105 B.n869 B.n60 10.6151
R1106 B.n865 B.n60 10.6151
R1107 B.n865 B.n864 10.6151
R1108 B.n864 B.n863 10.6151
R1109 B.n863 B.n62 10.6151
R1110 B.n859 B.n62 10.6151
R1111 B.n859 B.n858 10.6151
R1112 B.n858 B.n857 10.6151
R1113 B.n854 B.n853 10.6151
R1114 B.n853 B.n852 10.6151
R1115 B.n852 B.n68 10.6151
R1116 B.n848 B.n68 10.6151
R1117 B.n848 B.n847 10.6151
R1118 B.n847 B.n846 10.6151
R1119 B.n846 B.n70 10.6151
R1120 B.n842 B.n70 10.6151
R1121 B.n840 B.n839 10.6151
R1122 B.n839 B.n74 10.6151
R1123 B.n835 B.n74 10.6151
R1124 B.n835 B.n834 10.6151
R1125 B.n834 B.n833 10.6151
R1126 B.n833 B.n76 10.6151
R1127 B.n829 B.n76 10.6151
R1128 B.n829 B.n828 10.6151
R1129 B.n828 B.n827 10.6151
R1130 B.n827 B.n78 10.6151
R1131 B.n823 B.n78 10.6151
R1132 B.n823 B.n822 10.6151
R1133 B.n822 B.n821 10.6151
R1134 B.n821 B.n80 10.6151
R1135 B.n817 B.n80 10.6151
R1136 B.n817 B.n816 10.6151
R1137 B.n816 B.n815 10.6151
R1138 B.n815 B.n82 10.6151
R1139 B.n811 B.n82 10.6151
R1140 B.n811 B.n810 10.6151
R1141 B.n810 B.n809 10.6151
R1142 B.n809 B.n84 10.6151
R1143 B.n805 B.n84 10.6151
R1144 B.n805 B.n804 10.6151
R1145 B.n804 B.n803 10.6151
R1146 B.n803 B.n86 10.6151
R1147 B.n799 B.n86 10.6151
R1148 B.n799 B.n798 10.6151
R1149 B.n798 B.n797 10.6151
R1150 B.n797 B.n88 10.6151
R1151 B.n793 B.n88 10.6151
R1152 B.n793 B.n792 10.6151
R1153 B.n792 B.n791 10.6151
R1154 B.n791 B.n90 10.6151
R1155 B.n787 B.n90 10.6151
R1156 B.n787 B.n786 10.6151
R1157 B.n786 B.n785 10.6151
R1158 B.n785 B.n92 10.6151
R1159 B.n781 B.n92 10.6151
R1160 B.n781 B.n780 10.6151
R1161 B.n780 B.n779 10.6151
R1162 B.n779 B.n94 10.6151
R1163 B.n775 B.n94 10.6151
R1164 B.n775 B.n774 10.6151
R1165 B.n774 B.n773 10.6151
R1166 B.n773 B.n96 10.6151
R1167 B.n769 B.n96 10.6151
R1168 B.n769 B.n768 10.6151
R1169 B.n768 B.n767 10.6151
R1170 B.n767 B.n98 10.6151
R1171 B.n763 B.n98 10.6151
R1172 B.n763 B.n762 10.6151
R1173 B.n762 B.n761 10.6151
R1174 B.n761 B.n100 10.6151
R1175 B.n757 B.n100 10.6151
R1176 B.n757 B.n756 10.6151
R1177 B.n553 B.n168 10.6151
R1178 B.n557 B.n168 10.6151
R1179 B.n558 B.n557 10.6151
R1180 B.n559 B.n558 10.6151
R1181 B.n559 B.n166 10.6151
R1182 B.n563 B.n166 10.6151
R1183 B.n564 B.n563 10.6151
R1184 B.n565 B.n564 10.6151
R1185 B.n565 B.n164 10.6151
R1186 B.n569 B.n164 10.6151
R1187 B.n570 B.n569 10.6151
R1188 B.n571 B.n570 10.6151
R1189 B.n571 B.n162 10.6151
R1190 B.n575 B.n162 10.6151
R1191 B.n576 B.n575 10.6151
R1192 B.n577 B.n576 10.6151
R1193 B.n577 B.n160 10.6151
R1194 B.n581 B.n160 10.6151
R1195 B.n582 B.n581 10.6151
R1196 B.n583 B.n582 10.6151
R1197 B.n583 B.n158 10.6151
R1198 B.n587 B.n158 10.6151
R1199 B.n588 B.n587 10.6151
R1200 B.n589 B.n588 10.6151
R1201 B.n589 B.n156 10.6151
R1202 B.n593 B.n156 10.6151
R1203 B.n594 B.n593 10.6151
R1204 B.n595 B.n594 10.6151
R1205 B.n595 B.n154 10.6151
R1206 B.n599 B.n154 10.6151
R1207 B.n600 B.n599 10.6151
R1208 B.n601 B.n600 10.6151
R1209 B.n601 B.n152 10.6151
R1210 B.n605 B.n152 10.6151
R1211 B.n606 B.n605 10.6151
R1212 B.n607 B.n606 10.6151
R1213 B.n607 B.n150 10.6151
R1214 B.n611 B.n150 10.6151
R1215 B.n612 B.n611 10.6151
R1216 B.n613 B.n612 10.6151
R1217 B.n613 B.n148 10.6151
R1218 B.n617 B.n148 10.6151
R1219 B.n618 B.n617 10.6151
R1220 B.n619 B.n618 10.6151
R1221 B.n619 B.n146 10.6151
R1222 B.n623 B.n146 10.6151
R1223 B.n624 B.n623 10.6151
R1224 B.n625 B.n624 10.6151
R1225 B.n625 B.n144 10.6151
R1226 B.n629 B.n144 10.6151
R1227 B.n630 B.n629 10.6151
R1228 B.n631 B.n630 10.6151
R1229 B.n631 B.n142 10.6151
R1230 B.n635 B.n142 10.6151
R1231 B.n636 B.n635 10.6151
R1232 B.n637 B.n636 10.6151
R1233 B.n637 B.n140 10.6151
R1234 B.n641 B.n140 10.6151
R1235 B.n642 B.n641 10.6151
R1236 B.n643 B.n642 10.6151
R1237 B.n643 B.n138 10.6151
R1238 B.n647 B.n138 10.6151
R1239 B.n648 B.n647 10.6151
R1240 B.n649 B.n648 10.6151
R1241 B.n649 B.n136 10.6151
R1242 B.n653 B.n136 10.6151
R1243 B.n654 B.n653 10.6151
R1244 B.n655 B.n654 10.6151
R1245 B.n655 B.n134 10.6151
R1246 B.n659 B.n134 10.6151
R1247 B.n660 B.n659 10.6151
R1248 B.n661 B.n660 10.6151
R1249 B.n661 B.n132 10.6151
R1250 B.n665 B.n132 10.6151
R1251 B.n666 B.n665 10.6151
R1252 B.n667 B.n666 10.6151
R1253 B.n667 B.n130 10.6151
R1254 B.n671 B.n130 10.6151
R1255 B.n672 B.n671 10.6151
R1256 B.n673 B.n672 10.6151
R1257 B.n673 B.n128 10.6151
R1258 B.n677 B.n128 10.6151
R1259 B.n678 B.n677 10.6151
R1260 B.n679 B.n678 10.6151
R1261 B.n679 B.n126 10.6151
R1262 B.n683 B.n126 10.6151
R1263 B.n684 B.n683 10.6151
R1264 B.n685 B.n684 10.6151
R1265 B.n685 B.n124 10.6151
R1266 B.n689 B.n124 10.6151
R1267 B.n690 B.n689 10.6151
R1268 B.n691 B.n690 10.6151
R1269 B.n691 B.n122 10.6151
R1270 B.n695 B.n122 10.6151
R1271 B.n696 B.n695 10.6151
R1272 B.n697 B.n696 10.6151
R1273 B.n697 B.n120 10.6151
R1274 B.n701 B.n120 10.6151
R1275 B.n702 B.n701 10.6151
R1276 B.n703 B.n702 10.6151
R1277 B.n703 B.n118 10.6151
R1278 B.n707 B.n118 10.6151
R1279 B.n708 B.n707 10.6151
R1280 B.n709 B.n708 10.6151
R1281 B.n709 B.n116 10.6151
R1282 B.n713 B.n116 10.6151
R1283 B.n714 B.n713 10.6151
R1284 B.n715 B.n714 10.6151
R1285 B.n715 B.n114 10.6151
R1286 B.n719 B.n114 10.6151
R1287 B.n720 B.n719 10.6151
R1288 B.n721 B.n720 10.6151
R1289 B.n721 B.n112 10.6151
R1290 B.n725 B.n112 10.6151
R1291 B.n726 B.n725 10.6151
R1292 B.n727 B.n726 10.6151
R1293 B.n727 B.n110 10.6151
R1294 B.n731 B.n110 10.6151
R1295 B.n732 B.n731 10.6151
R1296 B.n733 B.n732 10.6151
R1297 B.n733 B.n108 10.6151
R1298 B.n737 B.n108 10.6151
R1299 B.n738 B.n737 10.6151
R1300 B.n739 B.n738 10.6151
R1301 B.n739 B.n106 10.6151
R1302 B.n743 B.n106 10.6151
R1303 B.n744 B.n743 10.6151
R1304 B.n745 B.n744 10.6151
R1305 B.n745 B.n104 10.6151
R1306 B.n749 B.n104 10.6151
R1307 B.n750 B.n749 10.6151
R1308 B.n751 B.n750 10.6151
R1309 B.n751 B.n102 10.6151
R1310 B.n755 B.n102 10.6151
R1311 B.n367 B.n234 10.6151
R1312 B.n371 B.n234 10.6151
R1313 B.n372 B.n371 10.6151
R1314 B.n373 B.n372 10.6151
R1315 B.n373 B.n232 10.6151
R1316 B.n377 B.n232 10.6151
R1317 B.n378 B.n377 10.6151
R1318 B.n379 B.n378 10.6151
R1319 B.n379 B.n230 10.6151
R1320 B.n383 B.n230 10.6151
R1321 B.n384 B.n383 10.6151
R1322 B.n385 B.n384 10.6151
R1323 B.n385 B.n228 10.6151
R1324 B.n389 B.n228 10.6151
R1325 B.n390 B.n389 10.6151
R1326 B.n391 B.n390 10.6151
R1327 B.n391 B.n226 10.6151
R1328 B.n395 B.n226 10.6151
R1329 B.n396 B.n395 10.6151
R1330 B.n397 B.n396 10.6151
R1331 B.n397 B.n224 10.6151
R1332 B.n401 B.n224 10.6151
R1333 B.n402 B.n401 10.6151
R1334 B.n403 B.n402 10.6151
R1335 B.n403 B.n222 10.6151
R1336 B.n407 B.n222 10.6151
R1337 B.n408 B.n407 10.6151
R1338 B.n409 B.n408 10.6151
R1339 B.n409 B.n220 10.6151
R1340 B.n413 B.n220 10.6151
R1341 B.n414 B.n413 10.6151
R1342 B.n415 B.n414 10.6151
R1343 B.n415 B.n218 10.6151
R1344 B.n419 B.n218 10.6151
R1345 B.n420 B.n419 10.6151
R1346 B.n421 B.n420 10.6151
R1347 B.n421 B.n216 10.6151
R1348 B.n425 B.n216 10.6151
R1349 B.n426 B.n425 10.6151
R1350 B.n427 B.n426 10.6151
R1351 B.n427 B.n214 10.6151
R1352 B.n431 B.n214 10.6151
R1353 B.n432 B.n431 10.6151
R1354 B.n433 B.n432 10.6151
R1355 B.n433 B.n212 10.6151
R1356 B.n437 B.n212 10.6151
R1357 B.n438 B.n437 10.6151
R1358 B.n439 B.n438 10.6151
R1359 B.n439 B.n210 10.6151
R1360 B.n443 B.n210 10.6151
R1361 B.n444 B.n443 10.6151
R1362 B.n445 B.n444 10.6151
R1363 B.n445 B.n208 10.6151
R1364 B.n449 B.n208 10.6151
R1365 B.n450 B.n449 10.6151
R1366 B.n451 B.n450 10.6151
R1367 B.n455 B.n454 10.6151
R1368 B.n456 B.n455 10.6151
R1369 B.n456 B.n202 10.6151
R1370 B.n460 B.n202 10.6151
R1371 B.n461 B.n460 10.6151
R1372 B.n462 B.n461 10.6151
R1373 B.n462 B.n200 10.6151
R1374 B.n466 B.n200 10.6151
R1375 B.n469 B.n468 10.6151
R1376 B.n469 B.n196 10.6151
R1377 B.n473 B.n196 10.6151
R1378 B.n474 B.n473 10.6151
R1379 B.n475 B.n474 10.6151
R1380 B.n475 B.n194 10.6151
R1381 B.n479 B.n194 10.6151
R1382 B.n480 B.n479 10.6151
R1383 B.n481 B.n480 10.6151
R1384 B.n481 B.n192 10.6151
R1385 B.n485 B.n192 10.6151
R1386 B.n486 B.n485 10.6151
R1387 B.n487 B.n486 10.6151
R1388 B.n487 B.n190 10.6151
R1389 B.n491 B.n190 10.6151
R1390 B.n492 B.n491 10.6151
R1391 B.n493 B.n492 10.6151
R1392 B.n493 B.n188 10.6151
R1393 B.n497 B.n188 10.6151
R1394 B.n498 B.n497 10.6151
R1395 B.n499 B.n498 10.6151
R1396 B.n499 B.n186 10.6151
R1397 B.n503 B.n186 10.6151
R1398 B.n504 B.n503 10.6151
R1399 B.n505 B.n504 10.6151
R1400 B.n505 B.n184 10.6151
R1401 B.n509 B.n184 10.6151
R1402 B.n510 B.n509 10.6151
R1403 B.n511 B.n510 10.6151
R1404 B.n511 B.n182 10.6151
R1405 B.n515 B.n182 10.6151
R1406 B.n516 B.n515 10.6151
R1407 B.n517 B.n516 10.6151
R1408 B.n517 B.n180 10.6151
R1409 B.n521 B.n180 10.6151
R1410 B.n522 B.n521 10.6151
R1411 B.n523 B.n522 10.6151
R1412 B.n523 B.n178 10.6151
R1413 B.n527 B.n178 10.6151
R1414 B.n528 B.n527 10.6151
R1415 B.n529 B.n528 10.6151
R1416 B.n529 B.n176 10.6151
R1417 B.n533 B.n176 10.6151
R1418 B.n534 B.n533 10.6151
R1419 B.n535 B.n534 10.6151
R1420 B.n535 B.n174 10.6151
R1421 B.n539 B.n174 10.6151
R1422 B.n540 B.n539 10.6151
R1423 B.n541 B.n540 10.6151
R1424 B.n541 B.n172 10.6151
R1425 B.n545 B.n172 10.6151
R1426 B.n546 B.n545 10.6151
R1427 B.n547 B.n546 10.6151
R1428 B.n547 B.n170 10.6151
R1429 B.n551 B.n170 10.6151
R1430 B.n552 B.n551 10.6151
R1431 B.n366 B.n365 10.6151
R1432 B.n365 B.n236 10.6151
R1433 B.n361 B.n236 10.6151
R1434 B.n361 B.n360 10.6151
R1435 B.n360 B.n359 10.6151
R1436 B.n359 B.n238 10.6151
R1437 B.n355 B.n238 10.6151
R1438 B.n355 B.n354 10.6151
R1439 B.n354 B.n353 10.6151
R1440 B.n353 B.n240 10.6151
R1441 B.n349 B.n240 10.6151
R1442 B.n349 B.n348 10.6151
R1443 B.n348 B.n347 10.6151
R1444 B.n347 B.n242 10.6151
R1445 B.n343 B.n242 10.6151
R1446 B.n343 B.n342 10.6151
R1447 B.n342 B.n341 10.6151
R1448 B.n341 B.n244 10.6151
R1449 B.n337 B.n244 10.6151
R1450 B.n337 B.n336 10.6151
R1451 B.n336 B.n335 10.6151
R1452 B.n335 B.n246 10.6151
R1453 B.n331 B.n246 10.6151
R1454 B.n331 B.n330 10.6151
R1455 B.n330 B.n329 10.6151
R1456 B.n329 B.n248 10.6151
R1457 B.n325 B.n248 10.6151
R1458 B.n325 B.n324 10.6151
R1459 B.n324 B.n323 10.6151
R1460 B.n323 B.n250 10.6151
R1461 B.n319 B.n250 10.6151
R1462 B.n319 B.n318 10.6151
R1463 B.n318 B.n317 10.6151
R1464 B.n317 B.n252 10.6151
R1465 B.n313 B.n252 10.6151
R1466 B.n313 B.n312 10.6151
R1467 B.n312 B.n311 10.6151
R1468 B.n311 B.n254 10.6151
R1469 B.n307 B.n254 10.6151
R1470 B.n307 B.n306 10.6151
R1471 B.n306 B.n305 10.6151
R1472 B.n305 B.n256 10.6151
R1473 B.n301 B.n256 10.6151
R1474 B.n301 B.n300 10.6151
R1475 B.n300 B.n299 10.6151
R1476 B.n299 B.n258 10.6151
R1477 B.n295 B.n258 10.6151
R1478 B.n295 B.n294 10.6151
R1479 B.n294 B.n293 10.6151
R1480 B.n293 B.n260 10.6151
R1481 B.n289 B.n260 10.6151
R1482 B.n289 B.n288 10.6151
R1483 B.n288 B.n287 10.6151
R1484 B.n287 B.n262 10.6151
R1485 B.n283 B.n262 10.6151
R1486 B.n283 B.n282 10.6151
R1487 B.n282 B.n281 10.6151
R1488 B.n281 B.n264 10.6151
R1489 B.n277 B.n264 10.6151
R1490 B.n277 B.n276 10.6151
R1491 B.n276 B.n275 10.6151
R1492 B.n275 B.n266 10.6151
R1493 B.n271 B.n266 10.6151
R1494 B.n271 B.n270 10.6151
R1495 B.n270 B.n269 10.6151
R1496 B.n269 B.n0 10.6151
R1497 B.n1039 B.n1 10.6151
R1498 B.n1039 B.n1038 10.6151
R1499 B.n1038 B.n1037 10.6151
R1500 B.n1037 B.n4 10.6151
R1501 B.n1033 B.n4 10.6151
R1502 B.n1033 B.n1032 10.6151
R1503 B.n1032 B.n1031 10.6151
R1504 B.n1031 B.n6 10.6151
R1505 B.n1027 B.n6 10.6151
R1506 B.n1027 B.n1026 10.6151
R1507 B.n1026 B.n1025 10.6151
R1508 B.n1025 B.n8 10.6151
R1509 B.n1021 B.n8 10.6151
R1510 B.n1021 B.n1020 10.6151
R1511 B.n1020 B.n1019 10.6151
R1512 B.n1019 B.n10 10.6151
R1513 B.n1015 B.n10 10.6151
R1514 B.n1015 B.n1014 10.6151
R1515 B.n1014 B.n1013 10.6151
R1516 B.n1013 B.n12 10.6151
R1517 B.n1009 B.n12 10.6151
R1518 B.n1009 B.n1008 10.6151
R1519 B.n1008 B.n1007 10.6151
R1520 B.n1007 B.n14 10.6151
R1521 B.n1003 B.n14 10.6151
R1522 B.n1003 B.n1002 10.6151
R1523 B.n1002 B.n1001 10.6151
R1524 B.n1001 B.n16 10.6151
R1525 B.n997 B.n16 10.6151
R1526 B.n997 B.n996 10.6151
R1527 B.n996 B.n995 10.6151
R1528 B.n995 B.n18 10.6151
R1529 B.n991 B.n18 10.6151
R1530 B.n991 B.n990 10.6151
R1531 B.n990 B.n989 10.6151
R1532 B.n989 B.n20 10.6151
R1533 B.n985 B.n20 10.6151
R1534 B.n985 B.n984 10.6151
R1535 B.n984 B.n983 10.6151
R1536 B.n983 B.n22 10.6151
R1537 B.n979 B.n22 10.6151
R1538 B.n979 B.n978 10.6151
R1539 B.n978 B.n977 10.6151
R1540 B.n977 B.n24 10.6151
R1541 B.n973 B.n24 10.6151
R1542 B.n973 B.n972 10.6151
R1543 B.n972 B.n971 10.6151
R1544 B.n971 B.n26 10.6151
R1545 B.n967 B.n26 10.6151
R1546 B.n967 B.n966 10.6151
R1547 B.n966 B.n965 10.6151
R1548 B.n965 B.n28 10.6151
R1549 B.n961 B.n28 10.6151
R1550 B.n961 B.n960 10.6151
R1551 B.n960 B.n959 10.6151
R1552 B.n959 B.n30 10.6151
R1553 B.n955 B.n30 10.6151
R1554 B.n955 B.n954 10.6151
R1555 B.n954 B.n953 10.6151
R1556 B.n953 B.n32 10.6151
R1557 B.n949 B.n32 10.6151
R1558 B.n949 B.n948 10.6151
R1559 B.n948 B.n947 10.6151
R1560 B.n947 B.n34 10.6151
R1561 B.n943 B.n34 10.6151
R1562 B.n943 B.n942 10.6151
R1563 B.n854 B.n66 6.5566
R1564 B.n842 B.n841 6.5566
R1565 B.n454 B.n206 6.5566
R1566 B.n467 B.n466 6.5566
R1567 B.n857 B.n66 4.05904
R1568 B.n841 B.n840 4.05904
R1569 B.n451 B.n206 4.05904
R1570 B.n468 B.n467 4.05904
R1571 B.n1043 B.n0 2.81026
R1572 B.n1043 B.n1 2.81026
R1573 VN.n65 VN.n34 161.3
R1574 VN.n64 VN.n63 161.3
R1575 VN.n62 VN.n35 161.3
R1576 VN.n61 VN.n60 161.3
R1577 VN.n59 VN.n36 161.3
R1578 VN.n58 VN.n57 161.3
R1579 VN.n56 VN.n37 161.3
R1580 VN.n55 VN.n54 161.3
R1581 VN.n53 VN.n38 161.3
R1582 VN.n52 VN.n51 161.3
R1583 VN.n50 VN.n39 161.3
R1584 VN.n49 VN.n48 161.3
R1585 VN.n47 VN.n40 161.3
R1586 VN.n46 VN.n45 161.3
R1587 VN.n44 VN.n41 161.3
R1588 VN.n31 VN.n0 161.3
R1589 VN.n30 VN.n29 161.3
R1590 VN.n28 VN.n1 161.3
R1591 VN.n27 VN.n26 161.3
R1592 VN.n25 VN.n2 161.3
R1593 VN.n24 VN.n23 161.3
R1594 VN.n22 VN.n3 161.3
R1595 VN.n21 VN.n20 161.3
R1596 VN.n19 VN.n4 161.3
R1597 VN.n18 VN.n17 161.3
R1598 VN.n16 VN.n5 161.3
R1599 VN.n15 VN.n14 161.3
R1600 VN.n13 VN.n6 161.3
R1601 VN.n12 VN.n11 161.3
R1602 VN.n10 VN.n7 161.3
R1603 VN.n9 VN.t2 144.345
R1604 VN.n43 VN.t4 144.345
R1605 VN.n32 VN.t7 112.16
R1606 VN.n20 VN.t5 112.16
R1607 VN.n8 VN.t3 112.16
R1608 VN.n66 VN.t1 112.16
R1609 VN.n54 VN.t6 112.16
R1610 VN.n42 VN.t0 112.16
R1611 VN VN.n67 60.0195
R1612 VN.n33 VN.n32 57.7881
R1613 VN.n67 VN.n66 57.7881
R1614 VN.n9 VN.n8 50.586
R1615 VN.n43 VN.n42 50.586
R1616 VN.n14 VN.n13 40.577
R1617 VN.n14 VN.n5 40.577
R1618 VN.n26 VN.n25 40.577
R1619 VN.n26 VN.n1 40.577
R1620 VN.n48 VN.n47 40.577
R1621 VN.n48 VN.n39 40.577
R1622 VN.n60 VN.n59 40.577
R1623 VN.n60 VN.n35 40.577
R1624 VN.n8 VN.n7 24.5923
R1625 VN.n12 VN.n7 24.5923
R1626 VN.n13 VN.n12 24.5923
R1627 VN.n18 VN.n5 24.5923
R1628 VN.n19 VN.n18 24.5923
R1629 VN.n20 VN.n19 24.5923
R1630 VN.n20 VN.n3 24.5923
R1631 VN.n24 VN.n3 24.5923
R1632 VN.n25 VN.n24 24.5923
R1633 VN.n30 VN.n1 24.5923
R1634 VN.n31 VN.n30 24.5923
R1635 VN.n32 VN.n31 24.5923
R1636 VN.n47 VN.n46 24.5923
R1637 VN.n46 VN.n41 24.5923
R1638 VN.n42 VN.n41 24.5923
R1639 VN.n59 VN.n58 24.5923
R1640 VN.n58 VN.n37 24.5923
R1641 VN.n54 VN.n37 24.5923
R1642 VN.n54 VN.n53 24.5923
R1643 VN.n53 VN.n52 24.5923
R1644 VN.n52 VN.n39 24.5923
R1645 VN.n66 VN.n65 24.5923
R1646 VN.n65 VN.n64 24.5923
R1647 VN.n64 VN.n35 24.5923
R1648 VN.n44 VN.n43 2.51557
R1649 VN.n10 VN.n9 2.51557
R1650 VN.n67 VN.n34 0.417304
R1651 VN.n33 VN.n0 0.417304
R1652 VN VN.n33 0.394524
R1653 VN.n63 VN.n34 0.189894
R1654 VN.n63 VN.n62 0.189894
R1655 VN.n62 VN.n61 0.189894
R1656 VN.n61 VN.n36 0.189894
R1657 VN.n57 VN.n36 0.189894
R1658 VN.n57 VN.n56 0.189894
R1659 VN.n56 VN.n55 0.189894
R1660 VN.n55 VN.n38 0.189894
R1661 VN.n51 VN.n38 0.189894
R1662 VN.n51 VN.n50 0.189894
R1663 VN.n50 VN.n49 0.189894
R1664 VN.n49 VN.n40 0.189894
R1665 VN.n45 VN.n40 0.189894
R1666 VN.n45 VN.n44 0.189894
R1667 VN.n11 VN.n10 0.189894
R1668 VN.n11 VN.n6 0.189894
R1669 VN.n15 VN.n6 0.189894
R1670 VN.n16 VN.n15 0.189894
R1671 VN.n17 VN.n16 0.189894
R1672 VN.n17 VN.n4 0.189894
R1673 VN.n21 VN.n4 0.189894
R1674 VN.n22 VN.n21 0.189894
R1675 VN.n23 VN.n22 0.189894
R1676 VN.n23 VN.n2 0.189894
R1677 VN.n27 VN.n2 0.189894
R1678 VN.n28 VN.n27 0.189894
R1679 VN.n29 VN.n28 0.189894
R1680 VN.n29 VN.n0 0.189894
R1681 VDD2.n2 VDD2.n1 69.3192
R1682 VDD2.n2 VDD2.n0 69.3192
R1683 VDD2 VDD2.n5 69.3164
R1684 VDD2.n4 VDD2.n3 67.6507
R1685 VDD2.n4 VDD2.n2 53.9567
R1686 VDD2.n5 VDD2.t7 1.9036
R1687 VDD2.n5 VDD2.t2 1.9036
R1688 VDD2.n3 VDD2.t3 1.9036
R1689 VDD2.n3 VDD2.t6 1.9036
R1690 VDD2.n1 VDD2.t4 1.9036
R1691 VDD2.n1 VDD2.t5 1.9036
R1692 VDD2.n0 VDD2.t0 1.9036
R1693 VDD2.n0 VDD2.t1 1.9036
R1694 VDD2 VDD2.n4 1.78283
R1695 VTAIL.n11 VTAIL.t5 52.8749
R1696 VTAIL.n10 VTAIL.t10 52.8749
R1697 VTAIL.n7 VTAIL.t13 52.8749
R1698 VTAIL.n15 VTAIL.t7 52.8748
R1699 VTAIL.n2 VTAIL.t12 52.8748
R1700 VTAIL.n3 VTAIL.t4 52.8748
R1701 VTAIL.n6 VTAIL.t1 52.8748
R1702 VTAIL.n14 VTAIL.t6 52.8748
R1703 VTAIL.n13 VTAIL.n12 50.9719
R1704 VTAIL.n9 VTAIL.n8 50.9719
R1705 VTAIL.n1 VTAIL.n0 50.9716
R1706 VTAIL.n5 VTAIL.n4 50.9716
R1707 VTAIL.n15 VTAIL.n14 30.5393
R1708 VTAIL.n7 VTAIL.n6 30.5393
R1709 VTAIL.n9 VTAIL.n7 3.44878
R1710 VTAIL.n10 VTAIL.n9 3.44878
R1711 VTAIL.n13 VTAIL.n11 3.44878
R1712 VTAIL.n14 VTAIL.n13 3.44878
R1713 VTAIL.n6 VTAIL.n5 3.44878
R1714 VTAIL.n5 VTAIL.n3 3.44878
R1715 VTAIL.n2 VTAIL.n1 3.44878
R1716 VTAIL VTAIL.n15 3.39059
R1717 VTAIL.n0 VTAIL.t11 1.9036
R1718 VTAIL.n0 VTAIL.t9 1.9036
R1719 VTAIL.n4 VTAIL.t0 1.9036
R1720 VTAIL.n4 VTAIL.t3 1.9036
R1721 VTAIL.n12 VTAIL.t15 1.9036
R1722 VTAIL.n12 VTAIL.t2 1.9036
R1723 VTAIL.n8 VTAIL.t8 1.9036
R1724 VTAIL.n8 VTAIL.t14 1.9036
R1725 VTAIL.n11 VTAIL.n10 0.470328
R1726 VTAIL.n3 VTAIL.n2 0.470328
R1727 VTAIL VTAIL.n1 0.0586897
R1728 VP.n22 VP.n19 161.3
R1729 VP.n24 VP.n23 161.3
R1730 VP.n25 VP.n18 161.3
R1731 VP.n27 VP.n26 161.3
R1732 VP.n28 VP.n17 161.3
R1733 VP.n30 VP.n29 161.3
R1734 VP.n31 VP.n16 161.3
R1735 VP.n33 VP.n32 161.3
R1736 VP.n34 VP.n15 161.3
R1737 VP.n36 VP.n35 161.3
R1738 VP.n37 VP.n14 161.3
R1739 VP.n39 VP.n38 161.3
R1740 VP.n40 VP.n13 161.3
R1741 VP.n42 VP.n41 161.3
R1742 VP.n43 VP.n12 161.3
R1743 VP.n81 VP.n0 161.3
R1744 VP.n80 VP.n79 161.3
R1745 VP.n78 VP.n1 161.3
R1746 VP.n77 VP.n76 161.3
R1747 VP.n75 VP.n2 161.3
R1748 VP.n74 VP.n73 161.3
R1749 VP.n72 VP.n3 161.3
R1750 VP.n71 VP.n70 161.3
R1751 VP.n69 VP.n4 161.3
R1752 VP.n68 VP.n67 161.3
R1753 VP.n66 VP.n5 161.3
R1754 VP.n65 VP.n64 161.3
R1755 VP.n63 VP.n6 161.3
R1756 VP.n62 VP.n61 161.3
R1757 VP.n60 VP.n7 161.3
R1758 VP.n59 VP.n58 161.3
R1759 VP.n57 VP.n8 161.3
R1760 VP.n56 VP.n55 161.3
R1761 VP.n54 VP.n9 161.3
R1762 VP.n53 VP.n52 161.3
R1763 VP.n51 VP.n10 161.3
R1764 VP.n50 VP.n49 161.3
R1765 VP.n48 VP.n11 161.3
R1766 VP.n21 VP.t1 144.345
R1767 VP.n82 VP.t3 112.16
R1768 VP.n70 VP.t5 112.16
R1769 VP.n58 VP.t6 112.16
R1770 VP.n46 VP.t7 112.16
R1771 VP.n20 VP.t4 112.16
R1772 VP.n32 VP.t0 112.16
R1773 VP.n44 VP.t2 112.16
R1774 VP.n47 VP.n45 59.9817
R1775 VP.n47 VP.n46 57.7881
R1776 VP.n83 VP.n82 57.7881
R1777 VP.n45 VP.n44 57.7881
R1778 VP.n21 VP.n20 50.586
R1779 VP.n52 VP.n51 40.577
R1780 VP.n52 VP.n9 40.577
R1781 VP.n64 VP.n63 40.577
R1782 VP.n64 VP.n5 40.577
R1783 VP.n76 VP.n75 40.577
R1784 VP.n76 VP.n1 40.577
R1785 VP.n38 VP.n13 40.577
R1786 VP.n38 VP.n37 40.577
R1787 VP.n26 VP.n17 40.577
R1788 VP.n26 VP.n25 40.577
R1789 VP.n46 VP.n11 24.5923
R1790 VP.n50 VP.n11 24.5923
R1791 VP.n51 VP.n50 24.5923
R1792 VP.n56 VP.n9 24.5923
R1793 VP.n57 VP.n56 24.5923
R1794 VP.n58 VP.n57 24.5923
R1795 VP.n58 VP.n7 24.5923
R1796 VP.n62 VP.n7 24.5923
R1797 VP.n63 VP.n62 24.5923
R1798 VP.n68 VP.n5 24.5923
R1799 VP.n69 VP.n68 24.5923
R1800 VP.n70 VP.n69 24.5923
R1801 VP.n70 VP.n3 24.5923
R1802 VP.n74 VP.n3 24.5923
R1803 VP.n75 VP.n74 24.5923
R1804 VP.n80 VP.n1 24.5923
R1805 VP.n81 VP.n80 24.5923
R1806 VP.n82 VP.n81 24.5923
R1807 VP.n42 VP.n13 24.5923
R1808 VP.n43 VP.n42 24.5923
R1809 VP.n44 VP.n43 24.5923
R1810 VP.n30 VP.n17 24.5923
R1811 VP.n31 VP.n30 24.5923
R1812 VP.n32 VP.n31 24.5923
R1813 VP.n32 VP.n15 24.5923
R1814 VP.n36 VP.n15 24.5923
R1815 VP.n37 VP.n36 24.5923
R1816 VP.n20 VP.n19 24.5923
R1817 VP.n24 VP.n19 24.5923
R1818 VP.n25 VP.n24 24.5923
R1819 VP.n22 VP.n21 2.51554
R1820 VP.n45 VP.n12 0.417304
R1821 VP.n48 VP.n47 0.417304
R1822 VP.n83 VP.n0 0.417304
R1823 VP VP.n83 0.394524
R1824 VP.n23 VP.n22 0.189894
R1825 VP.n23 VP.n18 0.189894
R1826 VP.n27 VP.n18 0.189894
R1827 VP.n28 VP.n27 0.189894
R1828 VP.n29 VP.n28 0.189894
R1829 VP.n29 VP.n16 0.189894
R1830 VP.n33 VP.n16 0.189894
R1831 VP.n34 VP.n33 0.189894
R1832 VP.n35 VP.n34 0.189894
R1833 VP.n35 VP.n14 0.189894
R1834 VP.n39 VP.n14 0.189894
R1835 VP.n40 VP.n39 0.189894
R1836 VP.n41 VP.n40 0.189894
R1837 VP.n41 VP.n12 0.189894
R1838 VP.n49 VP.n48 0.189894
R1839 VP.n49 VP.n10 0.189894
R1840 VP.n53 VP.n10 0.189894
R1841 VP.n54 VP.n53 0.189894
R1842 VP.n55 VP.n54 0.189894
R1843 VP.n55 VP.n8 0.189894
R1844 VP.n59 VP.n8 0.189894
R1845 VP.n60 VP.n59 0.189894
R1846 VP.n61 VP.n60 0.189894
R1847 VP.n61 VP.n6 0.189894
R1848 VP.n65 VP.n6 0.189894
R1849 VP.n66 VP.n65 0.189894
R1850 VP.n67 VP.n66 0.189894
R1851 VP.n67 VP.n4 0.189894
R1852 VP.n71 VP.n4 0.189894
R1853 VP.n72 VP.n71 0.189894
R1854 VP.n73 VP.n72 0.189894
R1855 VP.n73 VP.n2 0.189894
R1856 VP.n77 VP.n2 0.189894
R1857 VP.n78 VP.n77 0.189894
R1858 VP.n79 VP.n78 0.189894
R1859 VP.n79 VP.n0 0.189894
R1860 VDD1 VDD1.n0 69.433
R1861 VDD1.n3 VDD1.n2 69.3192
R1862 VDD1.n3 VDD1.n1 69.3192
R1863 VDD1.n5 VDD1.n4 67.6505
R1864 VDD1.n5 VDD1.n3 54.5397
R1865 VDD1.n4 VDD1.t7 1.9036
R1866 VDD1.n4 VDD1.t5 1.9036
R1867 VDD1.n0 VDD1.t6 1.9036
R1868 VDD1.n0 VDD1.t3 1.9036
R1869 VDD1.n2 VDD1.t2 1.9036
R1870 VDD1.n2 VDD1.t4 1.9036
R1871 VDD1.n1 VDD1.t0 1.9036
R1872 VDD1.n1 VDD1.t1 1.9036
R1873 VDD1 VDD1.n5 1.66645
C0 VTAIL VN 13.4313f
C1 VDD1 VTAIL 9.95803f
C2 VDD2 B 2.24271f
C3 w_n4970_n4384# VTAIL 5.40421f
C4 VP B 2.63118f
C5 VDD2 VP 0.633406f
C6 VDD1 VN 0.153539f
C7 w_n4970_n4384# VN 10.5135f
C8 VDD1 w_n4970_n4384# 2.42705f
C9 VTAIL B 7.17688f
C10 VTAIL VDD2 10.019599f
C11 VTAIL VP 13.4454f
C12 VN B 1.5386f
C13 VN VDD2 12.924f
C14 VN VP 9.909491f
C15 VDD1 B 2.11302f
C16 VDD1 VDD2 2.32923f
C17 w_n4970_n4384# B 13.1774f
C18 w_n4970_n4384# VDD2 2.58664f
C19 VDD1 VP 13.402f
C20 w_n4970_n4384# VP 11.161799f
C21 VDD2 VSUBS 2.54299f
C22 VDD1 VSUBS 3.37638f
C23 VTAIL VSUBS 1.751912f
C24 VN VSUBS 8.34799f
C25 VP VSUBS 4.882145f
C26 B VSUBS 6.625776f
C27 w_n4970_n4384# VSUBS 0.26665p
C28 VDD1.t6 VSUBS 0.425882f
C29 VDD1.t3 VSUBS 0.425882f
C30 VDD1.n0 VSUBS 3.53531f
C31 VDD1.t0 VSUBS 0.425882f
C32 VDD1.t1 VSUBS 0.425882f
C33 VDD1.n1 VSUBS 3.53317f
C34 VDD1.t2 VSUBS 0.425882f
C35 VDD1.t4 VSUBS 0.425882f
C36 VDD1.n2 VSUBS 3.53317f
C37 VDD1.n3 VSUBS 6.11114f
C38 VDD1.t7 VSUBS 0.425882f
C39 VDD1.t5 VSUBS 0.425882f
C40 VDD1.n4 VSUBS 3.50521f
C41 VDD1.n5 VSUBS 5.08252f
C42 VP.n0 VSUBS 0.044011f
C43 VP.t3 VSUBS 4.0312f
C44 VP.n1 VSUBS 0.046271f
C45 VP.n2 VSUBS 0.023404f
C46 VP.n3 VSUBS 0.043401f
C47 VP.n4 VSUBS 0.023404f
C48 VP.t5 VSUBS 4.0312f
C49 VP.n5 VSUBS 0.046271f
C50 VP.n6 VSUBS 0.023404f
C51 VP.n7 VSUBS 0.043401f
C52 VP.n8 VSUBS 0.023404f
C53 VP.t6 VSUBS 4.0312f
C54 VP.n9 VSUBS 0.046271f
C55 VP.n10 VSUBS 0.023404f
C56 VP.n11 VSUBS 0.043401f
C57 VP.n12 VSUBS 0.044011f
C58 VP.t2 VSUBS 4.0312f
C59 VP.n13 VSUBS 0.046271f
C60 VP.n14 VSUBS 0.023404f
C61 VP.n15 VSUBS 0.043401f
C62 VP.n16 VSUBS 0.023404f
C63 VP.t0 VSUBS 4.0312f
C64 VP.n17 VSUBS 0.046271f
C65 VP.n18 VSUBS 0.023404f
C66 VP.n19 VSUBS 0.043401f
C67 VP.t1 VSUBS 4.38208f
C68 VP.t4 VSUBS 4.0312f
C69 VP.n20 VSUBS 1.48682f
C70 VP.n21 VSUBS 1.42135f
C71 VP.n22 VSUBS 0.297954f
C72 VP.n23 VSUBS 0.023404f
C73 VP.n24 VSUBS 0.043401f
C74 VP.n25 VSUBS 0.046271f
C75 VP.n26 VSUBS 0.018903f
C76 VP.n27 VSUBS 0.023404f
C77 VP.n28 VSUBS 0.023404f
C78 VP.n29 VSUBS 0.023404f
C79 VP.n30 VSUBS 0.043401f
C80 VP.n31 VSUBS 0.043401f
C81 VP.n32 VSUBS 1.41388f
C82 VP.n33 VSUBS 0.023404f
C83 VP.n34 VSUBS 0.023404f
C84 VP.n35 VSUBS 0.023404f
C85 VP.n36 VSUBS 0.043401f
C86 VP.n37 VSUBS 0.046271f
C87 VP.n38 VSUBS 0.018903f
C88 VP.n39 VSUBS 0.023404f
C89 VP.n40 VSUBS 0.023404f
C90 VP.n41 VSUBS 0.023404f
C91 VP.n42 VSUBS 0.043401f
C92 VP.n43 VSUBS 0.043401f
C93 VP.n44 VSUBS 1.49493f
C94 VP.n45 VSUBS 1.73398f
C95 VP.t7 VSUBS 4.0312f
C96 VP.n46 VSUBS 1.49493f
C97 VP.n47 VSUBS 1.74805f
C98 VP.n48 VSUBS 0.044011f
C99 VP.n49 VSUBS 0.023404f
C100 VP.n50 VSUBS 0.043401f
C101 VP.n51 VSUBS 0.046271f
C102 VP.n52 VSUBS 0.018903f
C103 VP.n53 VSUBS 0.023404f
C104 VP.n54 VSUBS 0.023404f
C105 VP.n55 VSUBS 0.023404f
C106 VP.n56 VSUBS 0.043401f
C107 VP.n57 VSUBS 0.043401f
C108 VP.n58 VSUBS 1.41388f
C109 VP.n59 VSUBS 0.023404f
C110 VP.n60 VSUBS 0.023404f
C111 VP.n61 VSUBS 0.023404f
C112 VP.n62 VSUBS 0.043401f
C113 VP.n63 VSUBS 0.046271f
C114 VP.n64 VSUBS 0.018903f
C115 VP.n65 VSUBS 0.023404f
C116 VP.n66 VSUBS 0.023404f
C117 VP.n67 VSUBS 0.023404f
C118 VP.n68 VSUBS 0.043401f
C119 VP.n69 VSUBS 0.043401f
C120 VP.n70 VSUBS 1.41388f
C121 VP.n71 VSUBS 0.023404f
C122 VP.n72 VSUBS 0.023404f
C123 VP.n73 VSUBS 0.023404f
C124 VP.n74 VSUBS 0.043401f
C125 VP.n75 VSUBS 0.046271f
C126 VP.n76 VSUBS 0.018903f
C127 VP.n77 VSUBS 0.023404f
C128 VP.n78 VSUBS 0.023404f
C129 VP.n79 VSUBS 0.023404f
C130 VP.n80 VSUBS 0.043401f
C131 VP.n81 VSUBS 0.043401f
C132 VP.n82 VSUBS 1.49493f
C133 VP.n83 VSUBS 0.065799f
C134 VTAIL.t11 VSUBS 0.329902f
C135 VTAIL.t9 VSUBS 0.329902f
C136 VTAIL.n0 VSUBS 2.55776f
C137 VTAIL.n1 VSUBS 0.886454f
C138 VTAIL.t12 VSUBS 3.34491f
C139 VTAIL.n2 VSUBS 1.03146f
C140 VTAIL.t4 VSUBS 3.34491f
C141 VTAIL.n3 VSUBS 1.03146f
C142 VTAIL.t0 VSUBS 0.329902f
C143 VTAIL.t3 VSUBS 0.329902f
C144 VTAIL.n4 VSUBS 2.55776f
C145 VTAIL.n5 VSUBS 1.15345f
C146 VTAIL.t1 VSUBS 3.34491f
C147 VTAIL.n6 VSUBS 2.75771f
C148 VTAIL.t13 VSUBS 3.34494f
C149 VTAIL.n7 VSUBS 2.75769f
C150 VTAIL.t8 VSUBS 0.329902f
C151 VTAIL.t14 VSUBS 0.329902f
C152 VTAIL.n8 VSUBS 2.55776f
C153 VTAIL.n9 VSUBS 1.15345f
C154 VTAIL.t10 VSUBS 3.34494f
C155 VTAIL.n10 VSUBS 1.03143f
C156 VTAIL.t5 VSUBS 3.34494f
C157 VTAIL.n11 VSUBS 1.03143f
C158 VTAIL.t15 VSUBS 0.329902f
C159 VTAIL.t2 VSUBS 0.329902f
C160 VTAIL.n12 VSUBS 2.55776f
C161 VTAIL.n13 VSUBS 1.15345f
C162 VTAIL.t6 VSUBS 3.34491f
C163 VTAIL.n14 VSUBS 2.75771f
C164 VTAIL.t7 VSUBS 3.34491f
C165 VTAIL.n15 VSUBS 2.75313f
C166 VDD2.t0 VSUBS 0.424701f
C167 VDD2.t1 VSUBS 0.424701f
C168 VDD2.n0 VSUBS 3.52337f
C169 VDD2.t4 VSUBS 0.424701f
C170 VDD2.t5 VSUBS 0.424701f
C171 VDD2.n1 VSUBS 3.52337f
C172 VDD2.n2 VSUBS 6.02957f
C173 VDD2.t3 VSUBS 0.424701f
C174 VDD2.t6 VSUBS 0.424701f
C175 VDD2.n3 VSUBS 3.4955f
C176 VDD2.n4 VSUBS 5.0286f
C177 VDD2.t7 VSUBS 0.424701f
C178 VDD2.t2 VSUBS 0.424701f
C179 VDD2.n5 VSUBS 3.52329f
C180 VN.n0 VSUBS 0.040673f
C181 VN.t7 VSUBS 3.72543f
C182 VN.n1 VSUBS 0.042762f
C183 VN.n2 VSUBS 0.021629f
C184 VN.n3 VSUBS 0.04011f
C185 VN.n4 VSUBS 0.021629f
C186 VN.t5 VSUBS 3.72543f
C187 VN.n5 VSUBS 0.042762f
C188 VN.n6 VSUBS 0.021629f
C189 VN.n7 VSUBS 0.04011f
C190 VN.t2 VSUBS 4.04971f
C191 VN.t3 VSUBS 3.72543f
C192 VN.n8 VSUBS 1.37404f
C193 VN.n9 VSUBS 1.31354f
C194 VN.n10 VSUBS 0.275354f
C195 VN.n11 VSUBS 0.021629f
C196 VN.n12 VSUBS 0.04011f
C197 VN.n13 VSUBS 0.042762f
C198 VN.n14 VSUBS 0.017469f
C199 VN.n15 VSUBS 0.021629f
C200 VN.n16 VSUBS 0.021629f
C201 VN.n17 VSUBS 0.021629f
C202 VN.n18 VSUBS 0.04011f
C203 VN.n19 VSUBS 0.04011f
C204 VN.n20 VSUBS 1.30664f
C205 VN.n21 VSUBS 0.021629f
C206 VN.n22 VSUBS 0.021629f
C207 VN.n23 VSUBS 0.021629f
C208 VN.n24 VSUBS 0.04011f
C209 VN.n25 VSUBS 0.042762f
C210 VN.n26 VSUBS 0.017469f
C211 VN.n27 VSUBS 0.021629f
C212 VN.n28 VSUBS 0.021629f
C213 VN.n29 VSUBS 0.021629f
C214 VN.n30 VSUBS 0.04011f
C215 VN.n31 VSUBS 0.04011f
C216 VN.n32 VSUBS 1.38154f
C217 VN.n33 VSUBS 0.060808f
C218 VN.n34 VSUBS 0.040673f
C219 VN.t1 VSUBS 3.72543f
C220 VN.n35 VSUBS 0.042762f
C221 VN.n36 VSUBS 0.021629f
C222 VN.n37 VSUBS 0.04011f
C223 VN.n38 VSUBS 0.021629f
C224 VN.t6 VSUBS 3.72543f
C225 VN.n39 VSUBS 0.042762f
C226 VN.n40 VSUBS 0.021629f
C227 VN.n41 VSUBS 0.04011f
C228 VN.t4 VSUBS 4.04971f
C229 VN.t0 VSUBS 3.72543f
C230 VN.n42 VSUBS 1.37404f
C231 VN.n43 VSUBS 1.31354f
C232 VN.n44 VSUBS 0.275354f
C233 VN.n45 VSUBS 0.021629f
C234 VN.n46 VSUBS 0.04011f
C235 VN.n47 VSUBS 0.042762f
C236 VN.n48 VSUBS 0.017469f
C237 VN.n49 VSUBS 0.021629f
C238 VN.n50 VSUBS 0.021629f
C239 VN.n51 VSUBS 0.021629f
C240 VN.n52 VSUBS 0.04011f
C241 VN.n53 VSUBS 0.04011f
C242 VN.n54 VSUBS 1.30664f
C243 VN.n55 VSUBS 0.021629f
C244 VN.n56 VSUBS 0.021629f
C245 VN.n57 VSUBS 0.021629f
C246 VN.n58 VSUBS 0.04011f
C247 VN.n59 VSUBS 0.042762f
C248 VN.n60 VSUBS 0.017469f
C249 VN.n61 VSUBS 0.021629f
C250 VN.n62 VSUBS 0.021629f
C251 VN.n63 VSUBS 0.021629f
C252 VN.n64 VSUBS 0.04011f
C253 VN.n65 VSUBS 0.04011f
C254 VN.n66 VSUBS 1.38154f
C255 VN.n67 VSUBS 1.6074f
C256 B.n0 VSUBS 0.004769f
C257 B.n1 VSUBS 0.004769f
C258 B.n2 VSUBS 0.007542f
C259 B.n3 VSUBS 0.007542f
C260 B.n4 VSUBS 0.007542f
C261 B.n5 VSUBS 0.007542f
C262 B.n6 VSUBS 0.007542f
C263 B.n7 VSUBS 0.007542f
C264 B.n8 VSUBS 0.007542f
C265 B.n9 VSUBS 0.007542f
C266 B.n10 VSUBS 0.007542f
C267 B.n11 VSUBS 0.007542f
C268 B.n12 VSUBS 0.007542f
C269 B.n13 VSUBS 0.007542f
C270 B.n14 VSUBS 0.007542f
C271 B.n15 VSUBS 0.007542f
C272 B.n16 VSUBS 0.007542f
C273 B.n17 VSUBS 0.007542f
C274 B.n18 VSUBS 0.007542f
C275 B.n19 VSUBS 0.007542f
C276 B.n20 VSUBS 0.007542f
C277 B.n21 VSUBS 0.007542f
C278 B.n22 VSUBS 0.007542f
C279 B.n23 VSUBS 0.007542f
C280 B.n24 VSUBS 0.007542f
C281 B.n25 VSUBS 0.007542f
C282 B.n26 VSUBS 0.007542f
C283 B.n27 VSUBS 0.007542f
C284 B.n28 VSUBS 0.007542f
C285 B.n29 VSUBS 0.007542f
C286 B.n30 VSUBS 0.007542f
C287 B.n31 VSUBS 0.007542f
C288 B.n32 VSUBS 0.007542f
C289 B.n33 VSUBS 0.007542f
C290 B.n34 VSUBS 0.007542f
C291 B.n35 VSUBS 0.016218f
C292 B.n36 VSUBS 0.007542f
C293 B.n37 VSUBS 0.007542f
C294 B.n38 VSUBS 0.007542f
C295 B.n39 VSUBS 0.007542f
C296 B.n40 VSUBS 0.007542f
C297 B.n41 VSUBS 0.007542f
C298 B.n42 VSUBS 0.007542f
C299 B.n43 VSUBS 0.007542f
C300 B.n44 VSUBS 0.007542f
C301 B.n45 VSUBS 0.007542f
C302 B.n46 VSUBS 0.007542f
C303 B.n47 VSUBS 0.007542f
C304 B.n48 VSUBS 0.007542f
C305 B.n49 VSUBS 0.007542f
C306 B.n50 VSUBS 0.007542f
C307 B.n51 VSUBS 0.007542f
C308 B.n52 VSUBS 0.007542f
C309 B.n53 VSUBS 0.007542f
C310 B.n54 VSUBS 0.007542f
C311 B.n55 VSUBS 0.007542f
C312 B.n56 VSUBS 0.007542f
C313 B.n57 VSUBS 0.007542f
C314 B.n58 VSUBS 0.007542f
C315 B.n59 VSUBS 0.007542f
C316 B.n60 VSUBS 0.007542f
C317 B.n61 VSUBS 0.007542f
C318 B.n62 VSUBS 0.007542f
C319 B.n63 VSUBS 0.007542f
C320 B.t8 VSUBS 0.618937f
C321 B.t7 VSUBS 0.648936f
C322 B.t6 VSUBS 3.08048f
C323 B.n64 VSUBS 0.394358f
C324 B.n65 VSUBS 0.082455f
C325 B.n66 VSUBS 0.017475f
C326 B.n67 VSUBS 0.007542f
C327 B.n68 VSUBS 0.007542f
C328 B.n69 VSUBS 0.007542f
C329 B.n70 VSUBS 0.007542f
C330 B.n71 VSUBS 0.007542f
C331 B.t5 VSUBS 0.618915f
C332 B.t4 VSUBS 0.64892f
C333 B.t3 VSUBS 3.08048f
C334 B.n72 VSUBS 0.394375f
C335 B.n73 VSUBS 0.082477f
C336 B.n74 VSUBS 0.007542f
C337 B.n75 VSUBS 0.007542f
C338 B.n76 VSUBS 0.007542f
C339 B.n77 VSUBS 0.007542f
C340 B.n78 VSUBS 0.007542f
C341 B.n79 VSUBS 0.007542f
C342 B.n80 VSUBS 0.007542f
C343 B.n81 VSUBS 0.007542f
C344 B.n82 VSUBS 0.007542f
C345 B.n83 VSUBS 0.007542f
C346 B.n84 VSUBS 0.007542f
C347 B.n85 VSUBS 0.007542f
C348 B.n86 VSUBS 0.007542f
C349 B.n87 VSUBS 0.007542f
C350 B.n88 VSUBS 0.007542f
C351 B.n89 VSUBS 0.007542f
C352 B.n90 VSUBS 0.007542f
C353 B.n91 VSUBS 0.007542f
C354 B.n92 VSUBS 0.007542f
C355 B.n93 VSUBS 0.007542f
C356 B.n94 VSUBS 0.007542f
C357 B.n95 VSUBS 0.007542f
C358 B.n96 VSUBS 0.007542f
C359 B.n97 VSUBS 0.007542f
C360 B.n98 VSUBS 0.007542f
C361 B.n99 VSUBS 0.007542f
C362 B.n100 VSUBS 0.007542f
C363 B.n101 VSUBS 0.017279f
C364 B.n102 VSUBS 0.007542f
C365 B.n103 VSUBS 0.007542f
C366 B.n104 VSUBS 0.007542f
C367 B.n105 VSUBS 0.007542f
C368 B.n106 VSUBS 0.007542f
C369 B.n107 VSUBS 0.007542f
C370 B.n108 VSUBS 0.007542f
C371 B.n109 VSUBS 0.007542f
C372 B.n110 VSUBS 0.007542f
C373 B.n111 VSUBS 0.007542f
C374 B.n112 VSUBS 0.007542f
C375 B.n113 VSUBS 0.007542f
C376 B.n114 VSUBS 0.007542f
C377 B.n115 VSUBS 0.007542f
C378 B.n116 VSUBS 0.007542f
C379 B.n117 VSUBS 0.007542f
C380 B.n118 VSUBS 0.007542f
C381 B.n119 VSUBS 0.007542f
C382 B.n120 VSUBS 0.007542f
C383 B.n121 VSUBS 0.007542f
C384 B.n122 VSUBS 0.007542f
C385 B.n123 VSUBS 0.007542f
C386 B.n124 VSUBS 0.007542f
C387 B.n125 VSUBS 0.007542f
C388 B.n126 VSUBS 0.007542f
C389 B.n127 VSUBS 0.007542f
C390 B.n128 VSUBS 0.007542f
C391 B.n129 VSUBS 0.007542f
C392 B.n130 VSUBS 0.007542f
C393 B.n131 VSUBS 0.007542f
C394 B.n132 VSUBS 0.007542f
C395 B.n133 VSUBS 0.007542f
C396 B.n134 VSUBS 0.007542f
C397 B.n135 VSUBS 0.007542f
C398 B.n136 VSUBS 0.007542f
C399 B.n137 VSUBS 0.007542f
C400 B.n138 VSUBS 0.007542f
C401 B.n139 VSUBS 0.007542f
C402 B.n140 VSUBS 0.007542f
C403 B.n141 VSUBS 0.007542f
C404 B.n142 VSUBS 0.007542f
C405 B.n143 VSUBS 0.007542f
C406 B.n144 VSUBS 0.007542f
C407 B.n145 VSUBS 0.007542f
C408 B.n146 VSUBS 0.007542f
C409 B.n147 VSUBS 0.007542f
C410 B.n148 VSUBS 0.007542f
C411 B.n149 VSUBS 0.007542f
C412 B.n150 VSUBS 0.007542f
C413 B.n151 VSUBS 0.007542f
C414 B.n152 VSUBS 0.007542f
C415 B.n153 VSUBS 0.007542f
C416 B.n154 VSUBS 0.007542f
C417 B.n155 VSUBS 0.007542f
C418 B.n156 VSUBS 0.007542f
C419 B.n157 VSUBS 0.007542f
C420 B.n158 VSUBS 0.007542f
C421 B.n159 VSUBS 0.007542f
C422 B.n160 VSUBS 0.007542f
C423 B.n161 VSUBS 0.007542f
C424 B.n162 VSUBS 0.007542f
C425 B.n163 VSUBS 0.007542f
C426 B.n164 VSUBS 0.007542f
C427 B.n165 VSUBS 0.007542f
C428 B.n166 VSUBS 0.007542f
C429 B.n167 VSUBS 0.007542f
C430 B.n168 VSUBS 0.007542f
C431 B.n169 VSUBS 0.017279f
C432 B.n170 VSUBS 0.007542f
C433 B.n171 VSUBS 0.007542f
C434 B.n172 VSUBS 0.007542f
C435 B.n173 VSUBS 0.007542f
C436 B.n174 VSUBS 0.007542f
C437 B.n175 VSUBS 0.007542f
C438 B.n176 VSUBS 0.007542f
C439 B.n177 VSUBS 0.007542f
C440 B.n178 VSUBS 0.007542f
C441 B.n179 VSUBS 0.007542f
C442 B.n180 VSUBS 0.007542f
C443 B.n181 VSUBS 0.007542f
C444 B.n182 VSUBS 0.007542f
C445 B.n183 VSUBS 0.007542f
C446 B.n184 VSUBS 0.007542f
C447 B.n185 VSUBS 0.007542f
C448 B.n186 VSUBS 0.007542f
C449 B.n187 VSUBS 0.007542f
C450 B.n188 VSUBS 0.007542f
C451 B.n189 VSUBS 0.007542f
C452 B.n190 VSUBS 0.007542f
C453 B.n191 VSUBS 0.007542f
C454 B.n192 VSUBS 0.007542f
C455 B.n193 VSUBS 0.007542f
C456 B.n194 VSUBS 0.007542f
C457 B.n195 VSUBS 0.007542f
C458 B.n196 VSUBS 0.007542f
C459 B.n197 VSUBS 0.007542f
C460 B.t10 VSUBS 0.618915f
C461 B.t11 VSUBS 0.64892f
C462 B.t9 VSUBS 3.08048f
C463 B.n198 VSUBS 0.394375f
C464 B.n199 VSUBS 0.082477f
C465 B.n200 VSUBS 0.007542f
C466 B.n201 VSUBS 0.007542f
C467 B.n202 VSUBS 0.007542f
C468 B.n203 VSUBS 0.007542f
C469 B.t1 VSUBS 0.618937f
C470 B.t2 VSUBS 0.648936f
C471 B.t0 VSUBS 3.08048f
C472 B.n204 VSUBS 0.394358f
C473 B.n205 VSUBS 0.082455f
C474 B.n206 VSUBS 0.017475f
C475 B.n207 VSUBS 0.007542f
C476 B.n208 VSUBS 0.007542f
C477 B.n209 VSUBS 0.007542f
C478 B.n210 VSUBS 0.007542f
C479 B.n211 VSUBS 0.007542f
C480 B.n212 VSUBS 0.007542f
C481 B.n213 VSUBS 0.007542f
C482 B.n214 VSUBS 0.007542f
C483 B.n215 VSUBS 0.007542f
C484 B.n216 VSUBS 0.007542f
C485 B.n217 VSUBS 0.007542f
C486 B.n218 VSUBS 0.007542f
C487 B.n219 VSUBS 0.007542f
C488 B.n220 VSUBS 0.007542f
C489 B.n221 VSUBS 0.007542f
C490 B.n222 VSUBS 0.007542f
C491 B.n223 VSUBS 0.007542f
C492 B.n224 VSUBS 0.007542f
C493 B.n225 VSUBS 0.007542f
C494 B.n226 VSUBS 0.007542f
C495 B.n227 VSUBS 0.007542f
C496 B.n228 VSUBS 0.007542f
C497 B.n229 VSUBS 0.007542f
C498 B.n230 VSUBS 0.007542f
C499 B.n231 VSUBS 0.007542f
C500 B.n232 VSUBS 0.007542f
C501 B.n233 VSUBS 0.007542f
C502 B.n234 VSUBS 0.007542f
C503 B.n235 VSUBS 0.016218f
C504 B.n236 VSUBS 0.007542f
C505 B.n237 VSUBS 0.007542f
C506 B.n238 VSUBS 0.007542f
C507 B.n239 VSUBS 0.007542f
C508 B.n240 VSUBS 0.007542f
C509 B.n241 VSUBS 0.007542f
C510 B.n242 VSUBS 0.007542f
C511 B.n243 VSUBS 0.007542f
C512 B.n244 VSUBS 0.007542f
C513 B.n245 VSUBS 0.007542f
C514 B.n246 VSUBS 0.007542f
C515 B.n247 VSUBS 0.007542f
C516 B.n248 VSUBS 0.007542f
C517 B.n249 VSUBS 0.007542f
C518 B.n250 VSUBS 0.007542f
C519 B.n251 VSUBS 0.007542f
C520 B.n252 VSUBS 0.007542f
C521 B.n253 VSUBS 0.007542f
C522 B.n254 VSUBS 0.007542f
C523 B.n255 VSUBS 0.007542f
C524 B.n256 VSUBS 0.007542f
C525 B.n257 VSUBS 0.007542f
C526 B.n258 VSUBS 0.007542f
C527 B.n259 VSUBS 0.007542f
C528 B.n260 VSUBS 0.007542f
C529 B.n261 VSUBS 0.007542f
C530 B.n262 VSUBS 0.007542f
C531 B.n263 VSUBS 0.007542f
C532 B.n264 VSUBS 0.007542f
C533 B.n265 VSUBS 0.007542f
C534 B.n266 VSUBS 0.007542f
C535 B.n267 VSUBS 0.007542f
C536 B.n268 VSUBS 0.007542f
C537 B.n269 VSUBS 0.007542f
C538 B.n270 VSUBS 0.007542f
C539 B.n271 VSUBS 0.007542f
C540 B.n272 VSUBS 0.007542f
C541 B.n273 VSUBS 0.007542f
C542 B.n274 VSUBS 0.007542f
C543 B.n275 VSUBS 0.007542f
C544 B.n276 VSUBS 0.007542f
C545 B.n277 VSUBS 0.007542f
C546 B.n278 VSUBS 0.007542f
C547 B.n279 VSUBS 0.007542f
C548 B.n280 VSUBS 0.007542f
C549 B.n281 VSUBS 0.007542f
C550 B.n282 VSUBS 0.007542f
C551 B.n283 VSUBS 0.007542f
C552 B.n284 VSUBS 0.007542f
C553 B.n285 VSUBS 0.007542f
C554 B.n286 VSUBS 0.007542f
C555 B.n287 VSUBS 0.007542f
C556 B.n288 VSUBS 0.007542f
C557 B.n289 VSUBS 0.007542f
C558 B.n290 VSUBS 0.007542f
C559 B.n291 VSUBS 0.007542f
C560 B.n292 VSUBS 0.007542f
C561 B.n293 VSUBS 0.007542f
C562 B.n294 VSUBS 0.007542f
C563 B.n295 VSUBS 0.007542f
C564 B.n296 VSUBS 0.007542f
C565 B.n297 VSUBS 0.007542f
C566 B.n298 VSUBS 0.007542f
C567 B.n299 VSUBS 0.007542f
C568 B.n300 VSUBS 0.007542f
C569 B.n301 VSUBS 0.007542f
C570 B.n302 VSUBS 0.007542f
C571 B.n303 VSUBS 0.007542f
C572 B.n304 VSUBS 0.007542f
C573 B.n305 VSUBS 0.007542f
C574 B.n306 VSUBS 0.007542f
C575 B.n307 VSUBS 0.007542f
C576 B.n308 VSUBS 0.007542f
C577 B.n309 VSUBS 0.007542f
C578 B.n310 VSUBS 0.007542f
C579 B.n311 VSUBS 0.007542f
C580 B.n312 VSUBS 0.007542f
C581 B.n313 VSUBS 0.007542f
C582 B.n314 VSUBS 0.007542f
C583 B.n315 VSUBS 0.007542f
C584 B.n316 VSUBS 0.007542f
C585 B.n317 VSUBS 0.007542f
C586 B.n318 VSUBS 0.007542f
C587 B.n319 VSUBS 0.007542f
C588 B.n320 VSUBS 0.007542f
C589 B.n321 VSUBS 0.007542f
C590 B.n322 VSUBS 0.007542f
C591 B.n323 VSUBS 0.007542f
C592 B.n324 VSUBS 0.007542f
C593 B.n325 VSUBS 0.007542f
C594 B.n326 VSUBS 0.007542f
C595 B.n327 VSUBS 0.007542f
C596 B.n328 VSUBS 0.007542f
C597 B.n329 VSUBS 0.007542f
C598 B.n330 VSUBS 0.007542f
C599 B.n331 VSUBS 0.007542f
C600 B.n332 VSUBS 0.007542f
C601 B.n333 VSUBS 0.007542f
C602 B.n334 VSUBS 0.007542f
C603 B.n335 VSUBS 0.007542f
C604 B.n336 VSUBS 0.007542f
C605 B.n337 VSUBS 0.007542f
C606 B.n338 VSUBS 0.007542f
C607 B.n339 VSUBS 0.007542f
C608 B.n340 VSUBS 0.007542f
C609 B.n341 VSUBS 0.007542f
C610 B.n342 VSUBS 0.007542f
C611 B.n343 VSUBS 0.007542f
C612 B.n344 VSUBS 0.007542f
C613 B.n345 VSUBS 0.007542f
C614 B.n346 VSUBS 0.007542f
C615 B.n347 VSUBS 0.007542f
C616 B.n348 VSUBS 0.007542f
C617 B.n349 VSUBS 0.007542f
C618 B.n350 VSUBS 0.007542f
C619 B.n351 VSUBS 0.007542f
C620 B.n352 VSUBS 0.007542f
C621 B.n353 VSUBS 0.007542f
C622 B.n354 VSUBS 0.007542f
C623 B.n355 VSUBS 0.007542f
C624 B.n356 VSUBS 0.007542f
C625 B.n357 VSUBS 0.007542f
C626 B.n358 VSUBS 0.007542f
C627 B.n359 VSUBS 0.007542f
C628 B.n360 VSUBS 0.007542f
C629 B.n361 VSUBS 0.007542f
C630 B.n362 VSUBS 0.007542f
C631 B.n363 VSUBS 0.007542f
C632 B.n364 VSUBS 0.007542f
C633 B.n365 VSUBS 0.007542f
C634 B.n366 VSUBS 0.016218f
C635 B.n367 VSUBS 0.017279f
C636 B.n368 VSUBS 0.017279f
C637 B.n369 VSUBS 0.007542f
C638 B.n370 VSUBS 0.007542f
C639 B.n371 VSUBS 0.007542f
C640 B.n372 VSUBS 0.007542f
C641 B.n373 VSUBS 0.007542f
C642 B.n374 VSUBS 0.007542f
C643 B.n375 VSUBS 0.007542f
C644 B.n376 VSUBS 0.007542f
C645 B.n377 VSUBS 0.007542f
C646 B.n378 VSUBS 0.007542f
C647 B.n379 VSUBS 0.007542f
C648 B.n380 VSUBS 0.007542f
C649 B.n381 VSUBS 0.007542f
C650 B.n382 VSUBS 0.007542f
C651 B.n383 VSUBS 0.007542f
C652 B.n384 VSUBS 0.007542f
C653 B.n385 VSUBS 0.007542f
C654 B.n386 VSUBS 0.007542f
C655 B.n387 VSUBS 0.007542f
C656 B.n388 VSUBS 0.007542f
C657 B.n389 VSUBS 0.007542f
C658 B.n390 VSUBS 0.007542f
C659 B.n391 VSUBS 0.007542f
C660 B.n392 VSUBS 0.007542f
C661 B.n393 VSUBS 0.007542f
C662 B.n394 VSUBS 0.007542f
C663 B.n395 VSUBS 0.007542f
C664 B.n396 VSUBS 0.007542f
C665 B.n397 VSUBS 0.007542f
C666 B.n398 VSUBS 0.007542f
C667 B.n399 VSUBS 0.007542f
C668 B.n400 VSUBS 0.007542f
C669 B.n401 VSUBS 0.007542f
C670 B.n402 VSUBS 0.007542f
C671 B.n403 VSUBS 0.007542f
C672 B.n404 VSUBS 0.007542f
C673 B.n405 VSUBS 0.007542f
C674 B.n406 VSUBS 0.007542f
C675 B.n407 VSUBS 0.007542f
C676 B.n408 VSUBS 0.007542f
C677 B.n409 VSUBS 0.007542f
C678 B.n410 VSUBS 0.007542f
C679 B.n411 VSUBS 0.007542f
C680 B.n412 VSUBS 0.007542f
C681 B.n413 VSUBS 0.007542f
C682 B.n414 VSUBS 0.007542f
C683 B.n415 VSUBS 0.007542f
C684 B.n416 VSUBS 0.007542f
C685 B.n417 VSUBS 0.007542f
C686 B.n418 VSUBS 0.007542f
C687 B.n419 VSUBS 0.007542f
C688 B.n420 VSUBS 0.007542f
C689 B.n421 VSUBS 0.007542f
C690 B.n422 VSUBS 0.007542f
C691 B.n423 VSUBS 0.007542f
C692 B.n424 VSUBS 0.007542f
C693 B.n425 VSUBS 0.007542f
C694 B.n426 VSUBS 0.007542f
C695 B.n427 VSUBS 0.007542f
C696 B.n428 VSUBS 0.007542f
C697 B.n429 VSUBS 0.007542f
C698 B.n430 VSUBS 0.007542f
C699 B.n431 VSUBS 0.007542f
C700 B.n432 VSUBS 0.007542f
C701 B.n433 VSUBS 0.007542f
C702 B.n434 VSUBS 0.007542f
C703 B.n435 VSUBS 0.007542f
C704 B.n436 VSUBS 0.007542f
C705 B.n437 VSUBS 0.007542f
C706 B.n438 VSUBS 0.007542f
C707 B.n439 VSUBS 0.007542f
C708 B.n440 VSUBS 0.007542f
C709 B.n441 VSUBS 0.007542f
C710 B.n442 VSUBS 0.007542f
C711 B.n443 VSUBS 0.007542f
C712 B.n444 VSUBS 0.007542f
C713 B.n445 VSUBS 0.007542f
C714 B.n446 VSUBS 0.007542f
C715 B.n447 VSUBS 0.007542f
C716 B.n448 VSUBS 0.007542f
C717 B.n449 VSUBS 0.007542f
C718 B.n450 VSUBS 0.007542f
C719 B.n451 VSUBS 0.005213f
C720 B.n452 VSUBS 0.007542f
C721 B.n453 VSUBS 0.007542f
C722 B.n454 VSUBS 0.0061f
C723 B.n455 VSUBS 0.007542f
C724 B.n456 VSUBS 0.007542f
C725 B.n457 VSUBS 0.007542f
C726 B.n458 VSUBS 0.007542f
C727 B.n459 VSUBS 0.007542f
C728 B.n460 VSUBS 0.007542f
C729 B.n461 VSUBS 0.007542f
C730 B.n462 VSUBS 0.007542f
C731 B.n463 VSUBS 0.007542f
C732 B.n464 VSUBS 0.007542f
C733 B.n465 VSUBS 0.007542f
C734 B.n466 VSUBS 0.0061f
C735 B.n467 VSUBS 0.017475f
C736 B.n468 VSUBS 0.005213f
C737 B.n469 VSUBS 0.007542f
C738 B.n470 VSUBS 0.007542f
C739 B.n471 VSUBS 0.007542f
C740 B.n472 VSUBS 0.007542f
C741 B.n473 VSUBS 0.007542f
C742 B.n474 VSUBS 0.007542f
C743 B.n475 VSUBS 0.007542f
C744 B.n476 VSUBS 0.007542f
C745 B.n477 VSUBS 0.007542f
C746 B.n478 VSUBS 0.007542f
C747 B.n479 VSUBS 0.007542f
C748 B.n480 VSUBS 0.007542f
C749 B.n481 VSUBS 0.007542f
C750 B.n482 VSUBS 0.007542f
C751 B.n483 VSUBS 0.007542f
C752 B.n484 VSUBS 0.007542f
C753 B.n485 VSUBS 0.007542f
C754 B.n486 VSUBS 0.007542f
C755 B.n487 VSUBS 0.007542f
C756 B.n488 VSUBS 0.007542f
C757 B.n489 VSUBS 0.007542f
C758 B.n490 VSUBS 0.007542f
C759 B.n491 VSUBS 0.007542f
C760 B.n492 VSUBS 0.007542f
C761 B.n493 VSUBS 0.007542f
C762 B.n494 VSUBS 0.007542f
C763 B.n495 VSUBS 0.007542f
C764 B.n496 VSUBS 0.007542f
C765 B.n497 VSUBS 0.007542f
C766 B.n498 VSUBS 0.007542f
C767 B.n499 VSUBS 0.007542f
C768 B.n500 VSUBS 0.007542f
C769 B.n501 VSUBS 0.007542f
C770 B.n502 VSUBS 0.007542f
C771 B.n503 VSUBS 0.007542f
C772 B.n504 VSUBS 0.007542f
C773 B.n505 VSUBS 0.007542f
C774 B.n506 VSUBS 0.007542f
C775 B.n507 VSUBS 0.007542f
C776 B.n508 VSUBS 0.007542f
C777 B.n509 VSUBS 0.007542f
C778 B.n510 VSUBS 0.007542f
C779 B.n511 VSUBS 0.007542f
C780 B.n512 VSUBS 0.007542f
C781 B.n513 VSUBS 0.007542f
C782 B.n514 VSUBS 0.007542f
C783 B.n515 VSUBS 0.007542f
C784 B.n516 VSUBS 0.007542f
C785 B.n517 VSUBS 0.007542f
C786 B.n518 VSUBS 0.007542f
C787 B.n519 VSUBS 0.007542f
C788 B.n520 VSUBS 0.007542f
C789 B.n521 VSUBS 0.007542f
C790 B.n522 VSUBS 0.007542f
C791 B.n523 VSUBS 0.007542f
C792 B.n524 VSUBS 0.007542f
C793 B.n525 VSUBS 0.007542f
C794 B.n526 VSUBS 0.007542f
C795 B.n527 VSUBS 0.007542f
C796 B.n528 VSUBS 0.007542f
C797 B.n529 VSUBS 0.007542f
C798 B.n530 VSUBS 0.007542f
C799 B.n531 VSUBS 0.007542f
C800 B.n532 VSUBS 0.007542f
C801 B.n533 VSUBS 0.007542f
C802 B.n534 VSUBS 0.007542f
C803 B.n535 VSUBS 0.007542f
C804 B.n536 VSUBS 0.007542f
C805 B.n537 VSUBS 0.007542f
C806 B.n538 VSUBS 0.007542f
C807 B.n539 VSUBS 0.007542f
C808 B.n540 VSUBS 0.007542f
C809 B.n541 VSUBS 0.007542f
C810 B.n542 VSUBS 0.007542f
C811 B.n543 VSUBS 0.007542f
C812 B.n544 VSUBS 0.007542f
C813 B.n545 VSUBS 0.007542f
C814 B.n546 VSUBS 0.007542f
C815 B.n547 VSUBS 0.007542f
C816 B.n548 VSUBS 0.007542f
C817 B.n549 VSUBS 0.007542f
C818 B.n550 VSUBS 0.007542f
C819 B.n551 VSUBS 0.007542f
C820 B.n552 VSUBS 0.017279f
C821 B.n553 VSUBS 0.016218f
C822 B.n554 VSUBS 0.016218f
C823 B.n555 VSUBS 0.007542f
C824 B.n556 VSUBS 0.007542f
C825 B.n557 VSUBS 0.007542f
C826 B.n558 VSUBS 0.007542f
C827 B.n559 VSUBS 0.007542f
C828 B.n560 VSUBS 0.007542f
C829 B.n561 VSUBS 0.007542f
C830 B.n562 VSUBS 0.007542f
C831 B.n563 VSUBS 0.007542f
C832 B.n564 VSUBS 0.007542f
C833 B.n565 VSUBS 0.007542f
C834 B.n566 VSUBS 0.007542f
C835 B.n567 VSUBS 0.007542f
C836 B.n568 VSUBS 0.007542f
C837 B.n569 VSUBS 0.007542f
C838 B.n570 VSUBS 0.007542f
C839 B.n571 VSUBS 0.007542f
C840 B.n572 VSUBS 0.007542f
C841 B.n573 VSUBS 0.007542f
C842 B.n574 VSUBS 0.007542f
C843 B.n575 VSUBS 0.007542f
C844 B.n576 VSUBS 0.007542f
C845 B.n577 VSUBS 0.007542f
C846 B.n578 VSUBS 0.007542f
C847 B.n579 VSUBS 0.007542f
C848 B.n580 VSUBS 0.007542f
C849 B.n581 VSUBS 0.007542f
C850 B.n582 VSUBS 0.007542f
C851 B.n583 VSUBS 0.007542f
C852 B.n584 VSUBS 0.007542f
C853 B.n585 VSUBS 0.007542f
C854 B.n586 VSUBS 0.007542f
C855 B.n587 VSUBS 0.007542f
C856 B.n588 VSUBS 0.007542f
C857 B.n589 VSUBS 0.007542f
C858 B.n590 VSUBS 0.007542f
C859 B.n591 VSUBS 0.007542f
C860 B.n592 VSUBS 0.007542f
C861 B.n593 VSUBS 0.007542f
C862 B.n594 VSUBS 0.007542f
C863 B.n595 VSUBS 0.007542f
C864 B.n596 VSUBS 0.007542f
C865 B.n597 VSUBS 0.007542f
C866 B.n598 VSUBS 0.007542f
C867 B.n599 VSUBS 0.007542f
C868 B.n600 VSUBS 0.007542f
C869 B.n601 VSUBS 0.007542f
C870 B.n602 VSUBS 0.007542f
C871 B.n603 VSUBS 0.007542f
C872 B.n604 VSUBS 0.007542f
C873 B.n605 VSUBS 0.007542f
C874 B.n606 VSUBS 0.007542f
C875 B.n607 VSUBS 0.007542f
C876 B.n608 VSUBS 0.007542f
C877 B.n609 VSUBS 0.007542f
C878 B.n610 VSUBS 0.007542f
C879 B.n611 VSUBS 0.007542f
C880 B.n612 VSUBS 0.007542f
C881 B.n613 VSUBS 0.007542f
C882 B.n614 VSUBS 0.007542f
C883 B.n615 VSUBS 0.007542f
C884 B.n616 VSUBS 0.007542f
C885 B.n617 VSUBS 0.007542f
C886 B.n618 VSUBS 0.007542f
C887 B.n619 VSUBS 0.007542f
C888 B.n620 VSUBS 0.007542f
C889 B.n621 VSUBS 0.007542f
C890 B.n622 VSUBS 0.007542f
C891 B.n623 VSUBS 0.007542f
C892 B.n624 VSUBS 0.007542f
C893 B.n625 VSUBS 0.007542f
C894 B.n626 VSUBS 0.007542f
C895 B.n627 VSUBS 0.007542f
C896 B.n628 VSUBS 0.007542f
C897 B.n629 VSUBS 0.007542f
C898 B.n630 VSUBS 0.007542f
C899 B.n631 VSUBS 0.007542f
C900 B.n632 VSUBS 0.007542f
C901 B.n633 VSUBS 0.007542f
C902 B.n634 VSUBS 0.007542f
C903 B.n635 VSUBS 0.007542f
C904 B.n636 VSUBS 0.007542f
C905 B.n637 VSUBS 0.007542f
C906 B.n638 VSUBS 0.007542f
C907 B.n639 VSUBS 0.007542f
C908 B.n640 VSUBS 0.007542f
C909 B.n641 VSUBS 0.007542f
C910 B.n642 VSUBS 0.007542f
C911 B.n643 VSUBS 0.007542f
C912 B.n644 VSUBS 0.007542f
C913 B.n645 VSUBS 0.007542f
C914 B.n646 VSUBS 0.007542f
C915 B.n647 VSUBS 0.007542f
C916 B.n648 VSUBS 0.007542f
C917 B.n649 VSUBS 0.007542f
C918 B.n650 VSUBS 0.007542f
C919 B.n651 VSUBS 0.007542f
C920 B.n652 VSUBS 0.007542f
C921 B.n653 VSUBS 0.007542f
C922 B.n654 VSUBS 0.007542f
C923 B.n655 VSUBS 0.007542f
C924 B.n656 VSUBS 0.007542f
C925 B.n657 VSUBS 0.007542f
C926 B.n658 VSUBS 0.007542f
C927 B.n659 VSUBS 0.007542f
C928 B.n660 VSUBS 0.007542f
C929 B.n661 VSUBS 0.007542f
C930 B.n662 VSUBS 0.007542f
C931 B.n663 VSUBS 0.007542f
C932 B.n664 VSUBS 0.007542f
C933 B.n665 VSUBS 0.007542f
C934 B.n666 VSUBS 0.007542f
C935 B.n667 VSUBS 0.007542f
C936 B.n668 VSUBS 0.007542f
C937 B.n669 VSUBS 0.007542f
C938 B.n670 VSUBS 0.007542f
C939 B.n671 VSUBS 0.007542f
C940 B.n672 VSUBS 0.007542f
C941 B.n673 VSUBS 0.007542f
C942 B.n674 VSUBS 0.007542f
C943 B.n675 VSUBS 0.007542f
C944 B.n676 VSUBS 0.007542f
C945 B.n677 VSUBS 0.007542f
C946 B.n678 VSUBS 0.007542f
C947 B.n679 VSUBS 0.007542f
C948 B.n680 VSUBS 0.007542f
C949 B.n681 VSUBS 0.007542f
C950 B.n682 VSUBS 0.007542f
C951 B.n683 VSUBS 0.007542f
C952 B.n684 VSUBS 0.007542f
C953 B.n685 VSUBS 0.007542f
C954 B.n686 VSUBS 0.007542f
C955 B.n687 VSUBS 0.007542f
C956 B.n688 VSUBS 0.007542f
C957 B.n689 VSUBS 0.007542f
C958 B.n690 VSUBS 0.007542f
C959 B.n691 VSUBS 0.007542f
C960 B.n692 VSUBS 0.007542f
C961 B.n693 VSUBS 0.007542f
C962 B.n694 VSUBS 0.007542f
C963 B.n695 VSUBS 0.007542f
C964 B.n696 VSUBS 0.007542f
C965 B.n697 VSUBS 0.007542f
C966 B.n698 VSUBS 0.007542f
C967 B.n699 VSUBS 0.007542f
C968 B.n700 VSUBS 0.007542f
C969 B.n701 VSUBS 0.007542f
C970 B.n702 VSUBS 0.007542f
C971 B.n703 VSUBS 0.007542f
C972 B.n704 VSUBS 0.007542f
C973 B.n705 VSUBS 0.007542f
C974 B.n706 VSUBS 0.007542f
C975 B.n707 VSUBS 0.007542f
C976 B.n708 VSUBS 0.007542f
C977 B.n709 VSUBS 0.007542f
C978 B.n710 VSUBS 0.007542f
C979 B.n711 VSUBS 0.007542f
C980 B.n712 VSUBS 0.007542f
C981 B.n713 VSUBS 0.007542f
C982 B.n714 VSUBS 0.007542f
C983 B.n715 VSUBS 0.007542f
C984 B.n716 VSUBS 0.007542f
C985 B.n717 VSUBS 0.007542f
C986 B.n718 VSUBS 0.007542f
C987 B.n719 VSUBS 0.007542f
C988 B.n720 VSUBS 0.007542f
C989 B.n721 VSUBS 0.007542f
C990 B.n722 VSUBS 0.007542f
C991 B.n723 VSUBS 0.007542f
C992 B.n724 VSUBS 0.007542f
C993 B.n725 VSUBS 0.007542f
C994 B.n726 VSUBS 0.007542f
C995 B.n727 VSUBS 0.007542f
C996 B.n728 VSUBS 0.007542f
C997 B.n729 VSUBS 0.007542f
C998 B.n730 VSUBS 0.007542f
C999 B.n731 VSUBS 0.007542f
C1000 B.n732 VSUBS 0.007542f
C1001 B.n733 VSUBS 0.007542f
C1002 B.n734 VSUBS 0.007542f
C1003 B.n735 VSUBS 0.007542f
C1004 B.n736 VSUBS 0.007542f
C1005 B.n737 VSUBS 0.007542f
C1006 B.n738 VSUBS 0.007542f
C1007 B.n739 VSUBS 0.007542f
C1008 B.n740 VSUBS 0.007542f
C1009 B.n741 VSUBS 0.007542f
C1010 B.n742 VSUBS 0.007542f
C1011 B.n743 VSUBS 0.007542f
C1012 B.n744 VSUBS 0.007542f
C1013 B.n745 VSUBS 0.007542f
C1014 B.n746 VSUBS 0.007542f
C1015 B.n747 VSUBS 0.007542f
C1016 B.n748 VSUBS 0.007542f
C1017 B.n749 VSUBS 0.007542f
C1018 B.n750 VSUBS 0.007542f
C1019 B.n751 VSUBS 0.007542f
C1020 B.n752 VSUBS 0.007542f
C1021 B.n753 VSUBS 0.007542f
C1022 B.n754 VSUBS 0.016218f
C1023 B.n755 VSUBS 0.017184f
C1024 B.n756 VSUBS 0.016313f
C1025 B.n757 VSUBS 0.007542f
C1026 B.n758 VSUBS 0.007542f
C1027 B.n759 VSUBS 0.007542f
C1028 B.n760 VSUBS 0.007542f
C1029 B.n761 VSUBS 0.007542f
C1030 B.n762 VSUBS 0.007542f
C1031 B.n763 VSUBS 0.007542f
C1032 B.n764 VSUBS 0.007542f
C1033 B.n765 VSUBS 0.007542f
C1034 B.n766 VSUBS 0.007542f
C1035 B.n767 VSUBS 0.007542f
C1036 B.n768 VSUBS 0.007542f
C1037 B.n769 VSUBS 0.007542f
C1038 B.n770 VSUBS 0.007542f
C1039 B.n771 VSUBS 0.007542f
C1040 B.n772 VSUBS 0.007542f
C1041 B.n773 VSUBS 0.007542f
C1042 B.n774 VSUBS 0.007542f
C1043 B.n775 VSUBS 0.007542f
C1044 B.n776 VSUBS 0.007542f
C1045 B.n777 VSUBS 0.007542f
C1046 B.n778 VSUBS 0.007542f
C1047 B.n779 VSUBS 0.007542f
C1048 B.n780 VSUBS 0.007542f
C1049 B.n781 VSUBS 0.007542f
C1050 B.n782 VSUBS 0.007542f
C1051 B.n783 VSUBS 0.007542f
C1052 B.n784 VSUBS 0.007542f
C1053 B.n785 VSUBS 0.007542f
C1054 B.n786 VSUBS 0.007542f
C1055 B.n787 VSUBS 0.007542f
C1056 B.n788 VSUBS 0.007542f
C1057 B.n789 VSUBS 0.007542f
C1058 B.n790 VSUBS 0.007542f
C1059 B.n791 VSUBS 0.007542f
C1060 B.n792 VSUBS 0.007542f
C1061 B.n793 VSUBS 0.007542f
C1062 B.n794 VSUBS 0.007542f
C1063 B.n795 VSUBS 0.007542f
C1064 B.n796 VSUBS 0.007542f
C1065 B.n797 VSUBS 0.007542f
C1066 B.n798 VSUBS 0.007542f
C1067 B.n799 VSUBS 0.007542f
C1068 B.n800 VSUBS 0.007542f
C1069 B.n801 VSUBS 0.007542f
C1070 B.n802 VSUBS 0.007542f
C1071 B.n803 VSUBS 0.007542f
C1072 B.n804 VSUBS 0.007542f
C1073 B.n805 VSUBS 0.007542f
C1074 B.n806 VSUBS 0.007542f
C1075 B.n807 VSUBS 0.007542f
C1076 B.n808 VSUBS 0.007542f
C1077 B.n809 VSUBS 0.007542f
C1078 B.n810 VSUBS 0.007542f
C1079 B.n811 VSUBS 0.007542f
C1080 B.n812 VSUBS 0.007542f
C1081 B.n813 VSUBS 0.007542f
C1082 B.n814 VSUBS 0.007542f
C1083 B.n815 VSUBS 0.007542f
C1084 B.n816 VSUBS 0.007542f
C1085 B.n817 VSUBS 0.007542f
C1086 B.n818 VSUBS 0.007542f
C1087 B.n819 VSUBS 0.007542f
C1088 B.n820 VSUBS 0.007542f
C1089 B.n821 VSUBS 0.007542f
C1090 B.n822 VSUBS 0.007542f
C1091 B.n823 VSUBS 0.007542f
C1092 B.n824 VSUBS 0.007542f
C1093 B.n825 VSUBS 0.007542f
C1094 B.n826 VSUBS 0.007542f
C1095 B.n827 VSUBS 0.007542f
C1096 B.n828 VSUBS 0.007542f
C1097 B.n829 VSUBS 0.007542f
C1098 B.n830 VSUBS 0.007542f
C1099 B.n831 VSUBS 0.007542f
C1100 B.n832 VSUBS 0.007542f
C1101 B.n833 VSUBS 0.007542f
C1102 B.n834 VSUBS 0.007542f
C1103 B.n835 VSUBS 0.007542f
C1104 B.n836 VSUBS 0.007542f
C1105 B.n837 VSUBS 0.007542f
C1106 B.n838 VSUBS 0.007542f
C1107 B.n839 VSUBS 0.007542f
C1108 B.n840 VSUBS 0.005213f
C1109 B.n841 VSUBS 0.017475f
C1110 B.n842 VSUBS 0.0061f
C1111 B.n843 VSUBS 0.007542f
C1112 B.n844 VSUBS 0.007542f
C1113 B.n845 VSUBS 0.007542f
C1114 B.n846 VSUBS 0.007542f
C1115 B.n847 VSUBS 0.007542f
C1116 B.n848 VSUBS 0.007542f
C1117 B.n849 VSUBS 0.007542f
C1118 B.n850 VSUBS 0.007542f
C1119 B.n851 VSUBS 0.007542f
C1120 B.n852 VSUBS 0.007542f
C1121 B.n853 VSUBS 0.007542f
C1122 B.n854 VSUBS 0.0061f
C1123 B.n855 VSUBS 0.007542f
C1124 B.n856 VSUBS 0.007542f
C1125 B.n857 VSUBS 0.005213f
C1126 B.n858 VSUBS 0.007542f
C1127 B.n859 VSUBS 0.007542f
C1128 B.n860 VSUBS 0.007542f
C1129 B.n861 VSUBS 0.007542f
C1130 B.n862 VSUBS 0.007542f
C1131 B.n863 VSUBS 0.007542f
C1132 B.n864 VSUBS 0.007542f
C1133 B.n865 VSUBS 0.007542f
C1134 B.n866 VSUBS 0.007542f
C1135 B.n867 VSUBS 0.007542f
C1136 B.n868 VSUBS 0.007542f
C1137 B.n869 VSUBS 0.007542f
C1138 B.n870 VSUBS 0.007542f
C1139 B.n871 VSUBS 0.007542f
C1140 B.n872 VSUBS 0.007542f
C1141 B.n873 VSUBS 0.007542f
C1142 B.n874 VSUBS 0.007542f
C1143 B.n875 VSUBS 0.007542f
C1144 B.n876 VSUBS 0.007542f
C1145 B.n877 VSUBS 0.007542f
C1146 B.n878 VSUBS 0.007542f
C1147 B.n879 VSUBS 0.007542f
C1148 B.n880 VSUBS 0.007542f
C1149 B.n881 VSUBS 0.007542f
C1150 B.n882 VSUBS 0.007542f
C1151 B.n883 VSUBS 0.007542f
C1152 B.n884 VSUBS 0.007542f
C1153 B.n885 VSUBS 0.007542f
C1154 B.n886 VSUBS 0.007542f
C1155 B.n887 VSUBS 0.007542f
C1156 B.n888 VSUBS 0.007542f
C1157 B.n889 VSUBS 0.007542f
C1158 B.n890 VSUBS 0.007542f
C1159 B.n891 VSUBS 0.007542f
C1160 B.n892 VSUBS 0.007542f
C1161 B.n893 VSUBS 0.007542f
C1162 B.n894 VSUBS 0.007542f
C1163 B.n895 VSUBS 0.007542f
C1164 B.n896 VSUBS 0.007542f
C1165 B.n897 VSUBS 0.007542f
C1166 B.n898 VSUBS 0.007542f
C1167 B.n899 VSUBS 0.007542f
C1168 B.n900 VSUBS 0.007542f
C1169 B.n901 VSUBS 0.007542f
C1170 B.n902 VSUBS 0.007542f
C1171 B.n903 VSUBS 0.007542f
C1172 B.n904 VSUBS 0.007542f
C1173 B.n905 VSUBS 0.007542f
C1174 B.n906 VSUBS 0.007542f
C1175 B.n907 VSUBS 0.007542f
C1176 B.n908 VSUBS 0.007542f
C1177 B.n909 VSUBS 0.007542f
C1178 B.n910 VSUBS 0.007542f
C1179 B.n911 VSUBS 0.007542f
C1180 B.n912 VSUBS 0.007542f
C1181 B.n913 VSUBS 0.007542f
C1182 B.n914 VSUBS 0.007542f
C1183 B.n915 VSUBS 0.007542f
C1184 B.n916 VSUBS 0.007542f
C1185 B.n917 VSUBS 0.007542f
C1186 B.n918 VSUBS 0.007542f
C1187 B.n919 VSUBS 0.007542f
C1188 B.n920 VSUBS 0.007542f
C1189 B.n921 VSUBS 0.007542f
C1190 B.n922 VSUBS 0.007542f
C1191 B.n923 VSUBS 0.007542f
C1192 B.n924 VSUBS 0.007542f
C1193 B.n925 VSUBS 0.007542f
C1194 B.n926 VSUBS 0.007542f
C1195 B.n927 VSUBS 0.007542f
C1196 B.n928 VSUBS 0.007542f
C1197 B.n929 VSUBS 0.007542f
C1198 B.n930 VSUBS 0.007542f
C1199 B.n931 VSUBS 0.007542f
C1200 B.n932 VSUBS 0.007542f
C1201 B.n933 VSUBS 0.007542f
C1202 B.n934 VSUBS 0.007542f
C1203 B.n935 VSUBS 0.007542f
C1204 B.n936 VSUBS 0.007542f
C1205 B.n937 VSUBS 0.007542f
C1206 B.n938 VSUBS 0.007542f
C1207 B.n939 VSUBS 0.007542f
C1208 B.n940 VSUBS 0.017279f
C1209 B.n941 VSUBS 0.017279f
C1210 B.n942 VSUBS 0.016218f
C1211 B.n943 VSUBS 0.007542f
C1212 B.n944 VSUBS 0.007542f
C1213 B.n945 VSUBS 0.007542f
C1214 B.n946 VSUBS 0.007542f
C1215 B.n947 VSUBS 0.007542f
C1216 B.n948 VSUBS 0.007542f
C1217 B.n949 VSUBS 0.007542f
C1218 B.n950 VSUBS 0.007542f
C1219 B.n951 VSUBS 0.007542f
C1220 B.n952 VSUBS 0.007542f
C1221 B.n953 VSUBS 0.007542f
C1222 B.n954 VSUBS 0.007542f
C1223 B.n955 VSUBS 0.007542f
C1224 B.n956 VSUBS 0.007542f
C1225 B.n957 VSUBS 0.007542f
C1226 B.n958 VSUBS 0.007542f
C1227 B.n959 VSUBS 0.007542f
C1228 B.n960 VSUBS 0.007542f
C1229 B.n961 VSUBS 0.007542f
C1230 B.n962 VSUBS 0.007542f
C1231 B.n963 VSUBS 0.007542f
C1232 B.n964 VSUBS 0.007542f
C1233 B.n965 VSUBS 0.007542f
C1234 B.n966 VSUBS 0.007542f
C1235 B.n967 VSUBS 0.007542f
C1236 B.n968 VSUBS 0.007542f
C1237 B.n969 VSUBS 0.007542f
C1238 B.n970 VSUBS 0.007542f
C1239 B.n971 VSUBS 0.007542f
C1240 B.n972 VSUBS 0.007542f
C1241 B.n973 VSUBS 0.007542f
C1242 B.n974 VSUBS 0.007542f
C1243 B.n975 VSUBS 0.007542f
C1244 B.n976 VSUBS 0.007542f
C1245 B.n977 VSUBS 0.007542f
C1246 B.n978 VSUBS 0.007542f
C1247 B.n979 VSUBS 0.007542f
C1248 B.n980 VSUBS 0.007542f
C1249 B.n981 VSUBS 0.007542f
C1250 B.n982 VSUBS 0.007542f
C1251 B.n983 VSUBS 0.007542f
C1252 B.n984 VSUBS 0.007542f
C1253 B.n985 VSUBS 0.007542f
C1254 B.n986 VSUBS 0.007542f
C1255 B.n987 VSUBS 0.007542f
C1256 B.n988 VSUBS 0.007542f
C1257 B.n989 VSUBS 0.007542f
C1258 B.n990 VSUBS 0.007542f
C1259 B.n991 VSUBS 0.007542f
C1260 B.n992 VSUBS 0.007542f
C1261 B.n993 VSUBS 0.007542f
C1262 B.n994 VSUBS 0.007542f
C1263 B.n995 VSUBS 0.007542f
C1264 B.n996 VSUBS 0.007542f
C1265 B.n997 VSUBS 0.007542f
C1266 B.n998 VSUBS 0.007542f
C1267 B.n999 VSUBS 0.007542f
C1268 B.n1000 VSUBS 0.007542f
C1269 B.n1001 VSUBS 0.007542f
C1270 B.n1002 VSUBS 0.007542f
C1271 B.n1003 VSUBS 0.007542f
C1272 B.n1004 VSUBS 0.007542f
C1273 B.n1005 VSUBS 0.007542f
C1274 B.n1006 VSUBS 0.007542f
C1275 B.n1007 VSUBS 0.007542f
C1276 B.n1008 VSUBS 0.007542f
C1277 B.n1009 VSUBS 0.007542f
C1278 B.n1010 VSUBS 0.007542f
C1279 B.n1011 VSUBS 0.007542f
C1280 B.n1012 VSUBS 0.007542f
C1281 B.n1013 VSUBS 0.007542f
C1282 B.n1014 VSUBS 0.007542f
C1283 B.n1015 VSUBS 0.007542f
C1284 B.n1016 VSUBS 0.007542f
C1285 B.n1017 VSUBS 0.007542f
C1286 B.n1018 VSUBS 0.007542f
C1287 B.n1019 VSUBS 0.007542f
C1288 B.n1020 VSUBS 0.007542f
C1289 B.n1021 VSUBS 0.007542f
C1290 B.n1022 VSUBS 0.007542f
C1291 B.n1023 VSUBS 0.007542f
C1292 B.n1024 VSUBS 0.007542f
C1293 B.n1025 VSUBS 0.007542f
C1294 B.n1026 VSUBS 0.007542f
C1295 B.n1027 VSUBS 0.007542f
C1296 B.n1028 VSUBS 0.007542f
C1297 B.n1029 VSUBS 0.007542f
C1298 B.n1030 VSUBS 0.007542f
C1299 B.n1031 VSUBS 0.007542f
C1300 B.n1032 VSUBS 0.007542f
C1301 B.n1033 VSUBS 0.007542f
C1302 B.n1034 VSUBS 0.007542f
C1303 B.n1035 VSUBS 0.007542f
C1304 B.n1036 VSUBS 0.007542f
C1305 B.n1037 VSUBS 0.007542f
C1306 B.n1038 VSUBS 0.007542f
C1307 B.n1039 VSUBS 0.007542f
C1308 B.n1040 VSUBS 0.007542f
C1309 B.n1041 VSUBS 0.007542f
C1310 B.n1042 VSUBS 0.007542f
C1311 B.n1043 VSUBS 0.017079f
.ends

