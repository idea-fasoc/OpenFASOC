* NGSPICE file created from diff_pair_sample_0751.ext - technology: sky130A

.subckt diff_pair_sample_0751 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 B.t23 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X1 VTAIL.t17 VN.t0 VDD2.t9 B.t23 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X2 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=3.26
X3 VTAIL.t19 VN.t1 VDD2.t8 B.t20 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X4 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=3.26
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=3.26
X6 VDD2.t7 VN.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=3.26
X7 VDD1.t6 VP.t1 VTAIL.t14 B.t0 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=3.26
X8 VDD1.t5 VP.t2 VTAIL.t13 B.t4 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X9 VDD1.t4 VP.t3 VTAIL.t12 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=3.26
X10 VDD2.t6 VN.t3 VTAIL.t16 B.t22 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=3.26
X11 VTAIL.t18 VN.t4 VDD2.t5 B.t21 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X12 VDD2.t4 VN.t5 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=3.26
X13 VDD1.t1 VP.t4 VTAIL.t11 B.t22 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=7.7805 ps=40.68 w=19.95 l=3.26
X14 VTAIL.t5 VN.t6 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X15 VDD2.t2 VN.t7 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=3.26
X16 VDD2.t1 VN.t8 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X17 VTAIL.t10 VP.t5 VDD1.t0 B.t21 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X18 VDD1.t9 VP.t6 VTAIL.t9 B.t1 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=3.29175 ps=20.28 w=19.95 l=3.26
X19 VTAIL.t8 VP.t7 VDD1.t8 B.t5 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X20 VDD2.t0 VN.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X21 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=7.7805 pd=40.68 as=0 ps=0 w=19.95 l=3.26
X22 VDD1.t3 VP.t8 VTAIL.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
X23 VTAIL.t6 VP.t9 VDD1.t2 B.t20 sky130_fd_pr__nfet_01v8 ad=3.29175 pd=20.28 as=3.29175 ps=20.28 w=19.95 l=3.26
R0 VP.n30 VP.t6 179.388
R1 VP.n32 VP.n31 161.3
R2 VP.n33 VP.n28 161.3
R3 VP.n35 VP.n34 161.3
R4 VP.n36 VP.n27 161.3
R5 VP.n38 VP.n37 161.3
R6 VP.n39 VP.n26 161.3
R7 VP.n41 VP.n40 161.3
R8 VP.n42 VP.n25 161.3
R9 VP.n44 VP.n43 161.3
R10 VP.n45 VP.n24 161.3
R11 VP.n47 VP.n46 161.3
R12 VP.n48 VP.n23 161.3
R13 VP.n50 VP.n49 161.3
R14 VP.n51 VP.n22 161.3
R15 VP.n53 VP.n52 161.3
R16 VP.n55 VP.n54 161.3
R17 VP.n56 VP.n20 161.3
R18 VP.n58 VP.n57 161.3
R19 VP.n59 VP.n19 161.3
R20 VP.n61 VP.n60 161.3
R21 VP.n62 VP.n18 161.3
R22 VP.n64 VP.n63 161.3
R23 VP.n111 VP.n110 161.3
R24 VP.n109 VP.n1 161.3
R25 VP.n108 VP.n107 161.3
R26 VP.n106 VP.n2 161.3
R27 VP.n105 VP.n104 161.3
R28 VP.n103 VP.n3 161.3
R29 VP.n102 VP.n101 161.3
R30 VP.n100 VP.n99 161.3
R31 VP.n98 VP.n5 161.3
R32 VP.n97 VP.n96 161.3
R33 VP.n95 VP.n6 161.3
R34 VP.n94 VP.n93 161.3
R35 VP.n92 VP.n7 161.3
R36 VP.n91 VP.n90 161.3
R37 VP.n89 VP.n8 161.3
R38 VP.n88 VP.n87 161.3
R39 VP.n86 VP.n9 161.3
R40 VP.n85 VP.n84 161.3
R41 VP.n83 VP.n10 161.3
R42 VP.n82 VP.n81 161.3
R43 VP.n80 VP.n11 161.3
R44 VP.n79 VP.n78 161.3
R45 VP.n77 VP.n76 161.3
R46 VP.n75 VP.n13 161.3
R47 VP.n74 VP.n73 161.3
R48 VP.n72 VP.n14 161.3
R49 VP.n71 VP.n70 161.3
R50 VP.n69 VP.n15 161.3
R51 VP.n68 VP.n67 161.3
R52 VP.n8 VP.t2 147.483
R53 VP.n16 VP.t3 147.483
R54 VP.n12 VP.t5 147.483
R55 VP.n4 VP.t7 147.483
R56 VP.n0 VP.t1 147.483
R57 VP.n25 VP.t8 147.483
R58 VP.n17 VP.t4 147.483
R59 VP.n21 VP.t9 147.483
R60 VP.n29 VP.t0 147.483
R61 VP.n66 VP.n16 81.2593
R62 VP.n112 VP.n0 81.2593
R63 VP.n65 VP.n17 81.2593
R64 VP.n30 VP.n29 70.1236
R65 VP.n66 VP.n65 62.738
R66 VP.n85 VP.n10 56.5193
R67 VP.n93 VP.n6 56.5193
R68 VP.n46 VP.n23 56.5193
R69 VP.n38 VP.n27 56.5193
R70 VP.n74 VP.n14 51.663
R71 VP.n104 VP.n2 51.663
R72 VP.n57 VP.n19 51.663
R73 VP.n70 VP.n14 29.3238
R74 VP.n108 VP.n2 29.3238
R75 VP.n61 VP.n19 29.3238
R76 VP.n69 VP.n68 24.4675
R77 VP.n70 VP.n69 24.4675
R78 VP.n75 VP.n74 24.4675
R79 VP.n76 VP.n75 24.4675
R80 VP.n80 VP.n79 24.4675
R81 VP.n81 VP.n80 24.4675
R82 VP.n81 VP.n10 24.4675
R83 VP.n86 VP.n85 24.4675
R84 VP.n87 VP.n86 24.4675
R85 VP.n87 VP.n8 24.4675
R86 VP.n91 VP.n8 24.4675
R87 VP.n92 VP.n91 24.4675
R88 VP.n93 VP.n92 24.4675
R89 VP.n97 VP.n6 24.4675
R90 VP.n98 VP.n97 24.4675
R91 VP.n99 VP.n98 24.4675
R92 VP.n103 VP.n102 24.4675
R93 VP.n104 VP.n103 24.4675
R94 VP.n109 VP.n108 24.4675
R95 VP.n110 VP.n109 24.4675
R96 VP.n62 VP.n61 24.4675
R97 VP.n63 VP.n62 24.4675
R98 VP.n50 VP.n23 24.4675
R99 VP.n51 VP.n50 24.4675
R100 VP.n52 VP.n51 24.4675
R101 VP.n56 VP.n55 24.4675
R102 VP.n57 VP.n56 24.4675
R103 VP.n39 VP.n38 24.4675
R104 VP.n40 VP.n39 24.4675
R105 VP.n40 VP.n25 24.4675
R106 VP.n44 VP.n25 24.4675
R107 VP.n45 VP.n44 24.4675
R108 VP.n46 VP.n45 24.4675
R109 VP.n33 VP.n32 24.4675
R110 VP.n34 VP.n33 24.4675
R111 VP.n34 VP.n27 24.4675
R112 VP.n76 VP.n12 20.0634
R113 VP.n102 VP.n4 20.0634
R114 VP.n55 VP.n21 20.0634
R115 VP.n68 VP.n16 8.80862
R116 VP.n110 VP.n0 8.80862
R117 VP.n63 VP.n17 8.80862
R118 VP.n31 VP.n30 4.46391
R119 VP.n79 VP.n12 4.40456
R120 VP.n99 VP.n4 4.40456
R121 VP.n52 VP.n21 4.40456
R122 VP.n32 VP.n29 4.40456
R123 VP.n65 VP.n64 0.354971
R124 VP.n67 VP.n66 0.354971
R125 VP.n112 VP.n111 0.354971
R126 VP VP.n112 0.26696
R127 VP.n31 VP.n28 0.189894
R128 VP.n35 VP.n28 0.189894
R129 VP.n36 VP.n35 0.189894
R130 VP.n37 VP.n36 0.189894
R131 VP.n37 VP.n26 0.189894
R132 VP.n41 VP.n26 0.189894
R133 VP.n42 VP.n41 0.189894
R134 VP.n43 VP.n42 0.189894
R135 VP.n43 VP.n24 0.189894
R136 VP.n47 VP.n24 0.189894
R137 VP.n48 VP.n47 0.189894
R138 VP.n49 VP.n48 0.189894
R139 VP.n49 VP.n22 0.189894
R140 VP.n53 VP.n22 0.189894
R141 VP.n54 VP.n53 0.189894
R142 VP.n54 VP.n20 0.189894
R143 VP.n58 VP.n20 0.189894
R144 VP.n59 VP.n58 0.189894
R145 VP.n60 VP.n59 0.189894
R146 VP.n60 VP.n18 0.189894
R147 VP.n64 VP.n18 0.189894
R148 VP.n67 VP.n15 0.189894
R149 VP.n71 VP.n15 0.189894
R150 VP.n72 VP.n71 0.189894
R151 VP.n73 VP.n72 0.189894
R152 VP.n73 VP.n13 0.189894
R153 VP.n77 VP.n13 0.189894
R154 VP.n78 VP.n77 0.189894
R155 VP.n78 VP.n11 0.189894
R156 VP.n82 VP.n11 0.189894
R157 VP.n83 VP.n82 0.189894
R158 VP.n84 VP.n83 0.189894
R159 VP.n84 VP.n9 0.189894
R160 VP.n88 VP.n9 0.189894
R161 VP.n89 VP.n88 0.189894
R162 VP.n90 VP.n89 0.189894
R163 VP.n90 VP.n7 0.189894
R164 VP.n94 VP.n7 0.189894
R165 VP.n95 VP.n94 0.189894
R166 VP.n96 VP.n95 0.189894
R167 VP.n96 VP.n5 0.189894
R168 VP.n100 VP.n5 0.189894
R169 VP.n101 VP.n100 0.189894
R170 VP.n101 VP.n3 0.189894
R171 VP.n105 VP.n3 0.189894
R172 VP.n106 VP.n105 0.189894
R173 VP.n107 VP.n106 0.189894
R174 VP.n107 VP.n1 0.189894
R175 VP.n111 VP.n1 0.189894
R176 VDD1.n1 VDD1.t9 62.936
R177 VDD1.n3 VDD1.t4 62.9359
R178 VDD1.n5 VDD1.n4 61.1145
R179 VDD1.n7 VDD1.n6 58.8488
R180 VDD1.n1 VDD1.n0 58.8488
R181 VDD1.n3 VDD1.n2 58.8487
R182 VDD1.n7 VDD1.n5 57.7444
R183 VDD1 VDD1.n7 2.26343
R184 VDD1.n6 VDD1.t2 0.992981
R185 VDD1.n6 VDD1.t1 0.992981
R186 VDD1.n0 VDD1.t7 0.992981
R187 VDD1.n0 VDD1.t3 0.992981
R188 VDD1.n4 VDD1.t8 0.992981
R189 VDD1.n4 VDD1.t6 0.992981
R190 VDD1.n2 VDD1.t0 0.992981
R191 VDD1.n2 VDD1.t5 0.992981
R192 VDD1 VDD1.n1 0.832397
R193 VDD1.n5 VDD1.n3 0.718861
R194 VTAIL.n16 VTAIL.t11 43.1624
R195 VTAIL.n11 VTAIL.t0 43.1624
R196 VTAIL.n17 VTAIL.t16 43.1623
R197 VTAIL.n2 VTAIL.t14 43.1623
R198 VTAIL.n15 VTAIL.n14 42.17
R199 VTAIL.n13 VTAIL.n12 42.17
R200 VTAIL.n10 VTAIL.n9 42.17
R201 VTAIL.n8 VTAIL.n7 42.17
R202 VTAIL.n19 VTAIL.n18 42.1699
R203 VTAIL.n1 VTAIL.n0 42.1699
R204 VTAIL.n4 VTAIL.n3 42.1699
R205 VTAIL.n6 VTAIL.n5 42.1699
R206 VTAIL.n8 VTAIL.n6 35.7548
R207 VTAIL.n17 VTAIL.n16 32.66
R208 VTAIL.n10 VTAIL.n8 3.09533
R209 VTAIL.n11 VTAIL.n10 3.09533
R210 VTAIL.n15 VTAIL.n13 3.09533
R211 VTAIL.n16 VTAIL.n15 3.09533
R212 VTAIL.n6 VTAIL.n4 3.09533
R213 VTAIL.n4 VTAIL.n2 3.09533
R214 VTAIL.n19 VTAIL.n17 3.09533
R215 VTAIL VTAIL.n1 2.37981
R216 VTAIL.n13 VTAIL.n11 2.01774
R217 VTAIL.n2 VTAIL.n1 2.01774
R218 VTAIL.n18 VTAIL.t3 0.992981
R219 VTAIL.n18 VTAIL.t19 0.992981
R220 VTAIL.n0 VTAIL.t1 0.992981
R221 VTAIL.n0 VTAIL.t17 0.992981
R222 VTAIL.n3 VTAIL.t13 0.992981
R223 VTAIL.n3 VTAIL.t8 0.992981
R224 VTAIL.n5 VTAIL.t12 0.992981
R225 VTAIL.n5 VTAIL.t10 0.992981
R226 VTAIL.n14 VTAIL.t7 0.992981
R227 VTAIL.n14 VTAIL.t6 0.992981
R228 VTAIL.n12 VTAIL.t9 0.992981
R229 VTAIL.n12 VTAIL.t15 0.992981
R230 VTAIL.n9 VTAIL.t4 0.992981
R231 VTAIL.n9 VTAIL.t5 0.992981
R232 VTAIL.n7 VTAIL.t2 0.992981
R233 VTAIL.n7 VTAIL.t18 0.992981
R234 VTAIL VTAIL.n19 0.716017
R235 B.n1281 B.n1280 585
R236 B.n480 B.n200 585
R237 B.n479 B.n478 585
R238 B.n477 B.n476 585
R239 B.n475 B.n474 585
R240 B.n473 B.n472 585
R241 B.n471 B.n470 585
R242 B.n469 B.n468 585
R243 B.n467 B.n466 585
R244 B.n465 B.n464 585
R245 B.n463 B.n462 585
R246 B.n461 B.n460 585
R247 B.n459 B.n458 585
R248 B.n457 B.n456 585
R249 B.n455 B.n454 585
R250 B.n453 B.n452 585
R251 B.n451 B.n450 585
R252 B.n449 B.n448 585
R253 B.n447 B.n446 585
R254 B.n445 B.n444 585
R255 B.n443 B.n442 585
R256 B.n441 B.n440 585
R257 B.n439 B.n438 585
R258 B.n437 B.n436 585
R259 B.n435 B.n434 585
R260 B.n433 B.n432 585
R261 B.n431 B.n430 585
R262 B.n429 B.n428 585
R263 B.n427 B.n426 585
R264 B.n425 B.n424 585
R265 B.n423 B.n422 585
R266 B.n421 B.n420 585
R267 B.n419 B.n418 585
R268 B.n417 B.n416 585
R269 B.n415 B.n414 585
R270 B.n413 B.n412 585
R271 B.n411 B.n410 585
R272 B.n409 B.n408 585
R273 B.n407 B.n406 585
R274 B.n405 B.n404 585
R275 B.n403 B.n402 585
R276 B.n401 B.n400 585
R277 B.n399 B.n398 585
R278 B.n397 B.n396 585
R279 B.n395 B.n394 585
R280 B.n393 B.n392 585
R281 B.n391 B.n390 585
R282 B.n389 B.n388 585
R283 B.n387 B.n386 585
R284 B.n385 B.n384 585
R285 B.n383 B.n382 585
R286 B.n381 B.n380 585
R287 B.n379 B.n378 585
R288 B.n377 B.n376 585
R289 B.n375 B.n374 585
R290 B.n373 B.n372 585
R291 B.n371 B.n370 585
R292 B.n369 B.n368 585
R293 B.n367 B.n366 585
R294 B.n365 B.n364 585
R295 B.n363 B.n362 585
R296 B.n361 B.n360 585
R297 B.n359 B.n358 585
R298 B.n357 B.n356 585
R299 B.n355 B.n354 585
R300 B.n352 B.n351 585
R301 B.n350 B.n349 585
R302 B.n348 B.n347 585
R303 B.n346 B.n345 585
R304 B.n344 B.n343 585
R305 B.n342 B.n341 585
R306 B.n340 B.n339 585
R307 B.n338 B.n337 585
R308 B.n336 B.n335 585
R309 B.n334 B.n333 585
R310 B.n331 B.n330 585
R311 B.n329 B.n328 585
R312 B.n327 B.n326 585
R313 B.n325 B.n324 585
R314 B.n323 B.n322 585
R315 B.n321 B.n320 585
R316 B.n319 B.n318 585
R317 B.n317 B.n316 585
R318 B.n315 B.n314 585
R319 B.n313 B.n312 585
R320 B.n311 B.n310 585
R321 B.n309 B.n308 585
R322 B.n307 B.n306 585
R323 B.n305 B.n304 585
R324 B.n303 B.n302 585
R325 B.n301 B.n300 585
R326 B.n299 B.n298 585
R327 B.n297 B.n296 585
R328 B.n295 B.n294 585
R329 B.n293 B.n292 585
R330 B.n291 B.n290 585
R331 B.n289 B.n288 585
R332 B.n287 B.n286 585
R333 B.n285 B.n284 585
R334 B.n283 B.n282 585
R335 B.n281 B.n280 585
R336 B.n279 B.n278 585
R337 B.n277 B.n276 585
R338 B.n275 B.n274 585
R339 B.n273 B.n272 585
R340 B.n271 B.n270 585
R341 B.n269 B.n268 585
R342 B.n267 B.n266 585
R343 B.n265 B.n264 585
R344 B.n263 B.n262 585
R345 B.n261 B.n260 585
R346 B.n259 B.n258 585
R347 B.n257 B.n256 585
R348 B.n255 B.n254 585
R349 B.n253 B.n252 585
R350 B.n251 B.n250 585
R351 B.n249 B.n248 585
R352 B.n247 B.n246 585
R353 B.n245 B.n244 585
R354 B.n243 B.n242 585
R355 B.n241 B.n240 585
R356 B.n239 B.n238 585
R357 B.n237 B.n236 585
R358 B.n235 B.n234 585
R359 B.n233 B.n232 585
R360 B.n231 B.n230 585
R361 B.n229 B.n228 585
R362 B.n227 B.n226 585
R363 B.n225 B.n224 585
R364 B.n223 B.n222 585
R365 B.n221 B.n220 585
R366 B.n219 B.n218 585
R367 B.n217 B.n216 585
R368 B.n215 B.n214 585
R369 B.n213 B.n212 585
R370 B.n211 B.n210 585
R371 B.n209 B.n208 585
R372 B.n207 B.n206 585
R373 B.n131 B.n130 585
R374 B.n1286 B.n1285 585
R375 B.n1279 B.n201 585
R376 B.n201 B.n128 585
R377 B.n1278 B.n127 585
R378 B.n1290 B.n127 585
R379 B.n1277 B.n126 585
R380 B.n1291 B.n126 585
R381 B.n1276 B.n125 585
R382 B.n1292 B.n125 585
R383 B.n1275 B.n1274 585
R384 B.n1274 B.n121 585
R385 B.n1273 B.n120 585
R386 B.n1298 B.n120 585
R387 B.n1272 B.n119 585
R388 B.n1299 B.n119 585
R389 B.n1271 B.n118 585
R390 B.n1300 B.n118 585
R391 B.n1270 B.n1269 585
R392 B.n1269 B.n117 585
R393 B.n1268 B.n113 585
R394 B.n1306 B.n113 585
R395 B.n1267 B.n112 585
R396 B.n1307 B.n112 585
R397 B.n1266 B.n111 585
R398 B.n1308 B.n111 585
R399 B.n1265 B.n1264 585
R400 B.n1264 B.n107 585
R401 B.n1263 B.n106 585
R402 B.n1314 B.n106 585
R403 B.n1262 B.n105 585
R404 B.n1315 B.n105 585
R405 B.n1261 B.n104 585
R406 B.n1316 B.n104 585
R407 B.n1260 B.n1259 585
R408 B.n1259 B.n100 585
R409 B.n1258 B.n99 585
R410 B.n1322 B.n99 585
R411 B.n1257 B.n98 585
R412 B.n1323 B.n98 585
R413 B.n1256 B.n97 585
R414 B.n1324 B.n97 585
R415 B.n1255 B.n1254 585
R416 B.n1254 B.n93 585
R417 B.n1253 B.n92 585
R418 B.n1330 B.n92 585
R419 B.n1252 B.n91 585
R420 B.n1331 B.n91 585
R421 B.n1251 B.n90 585
R422 B.n1332 B.n90 585
R423 B.n1250 B.n1249 585
R424 B.n1249 B.n86 585
R425 B.n1248 B.n85 585
R426 B.n1338 B.n85 585
R427 B.n1247 B.n84 585
R428 B.n1339 B.n84 585
R429 B.n1246 B.n83 585
R430 B.n1340 B.n83 585
R431 B.n1245 B.n1244 585
R432 B.n1244 B.n79 585
R433 B.n1243 B.n78 585
R434 B.n1346 B.n78 585
R435 B.n1242 B.n77 585
R436 B.n1347 B.n77 585
R437 B.n1241 B.n76 585
R438 B.n1348 B.n76 585
R439 B.n1240 B.n1239 585
R440 B.n1239 B.n75 585
R441 B.n1238 B.n71 585
R442 B.n1354 B.n71 585
R443 B.n1237 B.n70 585
R444 B.n1355 B.n70 585
R445 B.n1236 B.n69 585
R446 B.n1356 B.n69 585
R447 B.n1235 B.n1234 585
R448 B.n1234 B.n65 585
R449 B.n1233 B.n64 585
R450 B.n1362 B.n64 585
R451 B.n1232 B.n63 585
R452 B.n1363 B.n63 585
R453 B.n1231 B.n62 585
R454 B.n1364 B.n62 585
R455 B.n1230 B.n1229 585
R456 B.n1229 B.n58 585
R457 B.n1228 B.n57 585
R458 B.n1370 B.n57 585
R459 B.n1227 B.n56 585
R460 B.n1371 B.n56 585
R461 B.n1226 B.n55 585
R462 B.n1372 B.n55 585
R463 B.n1225 B.n1224 585
R464 B.n1224 B.n51 585
R465 B.n1223 B.n50 585
R466 B.n1378 B.n50 585
R467 B.n1222 B.n49 585
R468 B.n1379 B.n49 585
R469 B.n1221 B.n48 585
R470 B.n1380 B.n48 585
R471 B.n1220 B.n1219 585
R472 B.n1219 B.n44 585
R473 B.n1218 B.n43 585
R474 B.n1386 B.n43 585
R475 B.n1217 B.n42 585
R476 B.n1387 B.n42 585
R477 B.n1216 B.n41 585
R478 B.n1388 B.n41 585
R479 B.n1215 B.n1214 585
R480 B.n1214 B.n37 585
R481 B.n1213 B.n36 585
R482 B.n1394 B.n36 585
R483 B.n1212 B.n35 585
R484 B.n1395 B.n35 585
R485 B.n1211 B.n34 585
R486 B.n1396 B.n34 585
R487 B.n1210 B.n1209 585
R488 B.n1209 B.n30 585
R489 B.n1208 B.n29 585
R490 B.n1402 B.n29 585
R491 B.n1207 B.n28 585
R492 B.n1403 B.n28 585
R493 B.n1206 B.n27 585
R494 B.n1404 B.n27 585
R495 B.n1205 B.n1204 585
R496 B.n1204 B.n23 585
R497 B.n1203 B.n22 585
R498 B.n1410 B.n22 585
R499 B.n1202 B.n21 585
R500 B.n1411 B.n21 585
R501 B.n1201 B.n20 585
R502 B.n1412 B.n20 585
R503 B.n1200 B.n1199 585
R504 B.n1199 B.n19 585
R505 B.n1198 B.n15 585
R506 B.n1418 B.n15 585
R507 B.n1197 B.n14 585
R508 B.n1419 B.n14 585
R509 B.n1196 B.n13 585
R510 B.n1420 B.n13 585
R511 B.n1195 B.n1194 585
R512 B.n1194 B.n12 585
R513 B.n1193 B.n1192 585
R514 B.n1193 B.n8 585
R515 B.n1191 B.n7 585
R516 B.n1427 B.n7 585
R517 B.n1190 B.n6 585
R518 B.n1428 B.n6 585
R519 B.n1189 B.n5 585
R520 B.n1429 B.n5 585
R521 B.n1188 B.n1187 585
R522 B.n1187 B.n4 585
R523 B.n1186 B.n481 585
R524 B.n1186 B.n1185 585
R525 B.n1176 B.n482 585
R526 B.n483 B.n482 585
R527 B.n1178 B.n1177 585
R528 B.n1179 B.n1178 585
R529 B.n1175 B.n488 585
R530 B.n488 B.n487 585
R531 B.n1174 B.n1173 585
R532 B.n1173 B.n1172 585
R533 B.n490 B.n489 585
R534 B.n1165 B.n490 585
R535 B.n1164 B.n1163 585
R536 B.n1166 B.n1164 585
R537 B.n1162 B.n495 585
R538 B.n495 B.n494 585
R539 B.n1161 B.n1160 585
R540 B.n1160 B.n1159 585
R541 B.n497 B.n496 585
R542 B.n498 B.n497 585
R543 B.n1152 B.n1151 585
R544 B.n1153 B.n1152 585
R545 B.n1150 B.n503 585
R546 B.n503 B.n502 585
R547 B.n1149 B.n1148 585
R548 B.n1148 B.n1147 585
R549 B.n505 B.n504 585
R550 B.n506 B.n505 585
R551 B.n1140 B.n1139 585
R552 B.n1141 B.n1140 585
R553 B.n1138 B.n510 585
R554 B.n514 B.n510 585
R555 B.n1137 B.n1136 585
R556 B.n1136 B.n1135 585
R557 B.n512 B.n511 585
R558 B.n513 B.n512 585
R559 B.n1128 B.n1127 585
R560 B.n1129 B.n1128 585
R561 B.n1126 B.n519 585
R562 B.n519 B.n518 585
R563 B.n1125 B.n1124 585
R564 B.n1124 B.n1123 585
R565 B.n521 B.n520 585
R566 B.n522 B.n521 585
R567 B.n1116 B.n1115 585
R568 B.n1117 B.n1116 585
R569 B.n1114 B.n527 585
R570 B.n527 B.n526 585
R571 B.n1113 B.n1112 585
R572 B.n1112 B.n1111 585
R573 B.n529 B.n528 585
R574 B.n530 B.n529 585
R575 B.n1104 B.n1103 585
R576 B.n1105 B.n1104 585
R577 B.n1102 B.n535 585
R578 B.n535 B.n534 585
R579 B.n1101 B.n1100 585
R580 B.n1100 B.n1099 585
R581 B.n537 B.n536 585
R582 B.n538 B.n537 585
R583 B.n1092 B.n1091 585
R584 B.n1093 B.n1092 585
R585 B.n1090 B.n543 585
R586 B.n543 B.n542 585
R587 B.n1089 B.n1088 585
R588 B.n1088 B.n1087 585
R589 B.n545 B.n544 585
R590 B.n546 B.n545 585
R591 B.n1080 B.n1079 585
R592 B.n1081 B.n1080 585
R593 B.n1078 B.n551 585
R594 B.n551 B.n550 585
R595 B.n1077 B.n1076 585
R596 B.n1076 B.n1075 585
R597 B.n553 B.n552 585
R598 B.n1068 B.n553 585
R599 B.n1067 B.n1066 585
R600 B.n1069 B.n1067 585
R601 B.n1065 B.n558 585
R602 B.n558 B.n557 585
R603 B.n1064 B.n1063 585
R604 B.n1063 B.n1062 585
R605 B.n560 B.n559 585
R606 B.n561 B.n560 585
R607 B.n1055 B.n1054 585
R608 B.n1056 B.n1055 585
R609 B.n1053 B.n566 585
R610 B.n566 B.n565 585
R611 B.n1052 B.n1051 585
R612 B.n1051 B.n1050 585
R613 B.n568 B.n567 585
R614 B.n569 B.n568 585
R615 B.n1043 B.n1042 585
R616 B.n1044 B.n1043 585
R617 B.n1041 B.n573 585
R618 B.n577 B.n573 585
R619 B.n1040 B.n1039 585
R620 B.n1039 B.n1038 585
R621 B.n575 B.n574 585
R622 B.n576 B.n575 585
R623 B.n1031 B.n1030 585
R624 B.n1032 B.n1031 585
R625 B.n1029 B.n582 585
R626 B.n582 B.n581 585
R627 B.n1028 B.n1027 585
R628 B.n1027 B.n1026 585
R629 B.n584 B.n583 585
R630 B.n585 B.n584 585
R631 B.n1019 B.n1018 585
R632 B.n1020 B.n1019 585
R633 B.n1017 B.n590 585
R634 B.n590 B.n589 585
R635 B.n1016 B.n1015 585
R636 B.n1015 B.n1014 585
R637 B.n592 B.n591 585
R638 B.n593 B.n592 585
R639 B.n1007 B.n1006 585
R640 B.n1008 B.n1007 585
R641 B.n1005 B.n598 585
R642 B.n598 B.n597 585
R643 B.n1004 B.n1003 585
R644 B.n1003 B.n1002 585
R645 B.n600 B.n599 585
R646 B.n995 B.n600 585
R647 B.n994 B.n993 585
R648 B.n996 B.n994 585
R649 B.n992 B.n605 585
R650 B.n605 B.n604 585
R651 B.n991 B.n990 585
R652 B.n990 B.n989 585
R653 B.n607 B.n606 585
R654 B.n608 B.n607 585
R655 B.n982 B.n981 585
R656 B.n983 B.n982 585
R657 B.n980 B.n613 585
R658 B.n613 B.n612 585
R659 B.n979 B.n978 585
R660 B.n978 B.n977 585
R661 B.n615 B.n614 585
R662 B.n616 B.n615 585
R663 B.n973 B.n972 585
R664 B.n619 B.n618 585
R665 B.n969 B.n968 585
R666 B.n970 B.n969 585
R667 B.n967 B.n689 585
R668 B.n966 B.n965 585
R669 B.n964 B.n963 585
R670 B.n962 B.n961 585
R671 B.n960 B.n959 585
R672 B.n958 B.n957 585
R673 B.n956 B.n955 585
R674 B.n954 B.n953 585
R675 B.n952 B.n951 585
R676 B.n950 B.n949 585
R677 B.n948 B.n947 585
R678 B.n946 B.n945 585
R679 B.n944 B.n943 585
R680 B.n942 B.n941 585
R681 B.n940 B.n939 585
R682 B.n938 B.n937 585
R683 B.n936 B.n935 585
R684 B.n934 B.n933 585
R685 B.n932 B.n931 585
R686 B.n930 B.n929 585
R687 B.n928 B.n927 585
R688 B.n926 B.n925 585
R689 B.n924 B.n923 585
R690 B.n922 B.n921 585
R691 B.n920 B.n919 585
R692 B.n918 B.n917 585
R693 B.n916 B.n915 585
R694 B.n914 B.n913 585
R695 B.n912 B.n911 585
R696 B.n910 B.n909 585
R697 B.n908 B.n907 585
R698 B.n906 B.n905 585
R699 B.n904 B.n903 585
R700 B.n902 B.n901 585
R701 B.n900 B.n899 585
R702 B.n898 B.n897 585
R703 B.n896 B.n895 585
R704 B.n894 B.n893 585
R705 B.n892 B.n891 585
R706 B.n890 B.n889 585
R707 B.n888 B.n887 585
R708 B.n886 B.n885 585
R709 B.n884 B.n883 585
R710 B.n882 B.n881 585
R711 B.n880 B.n879 585
R712 B.n878 B.n877 585
R713 B.n876 B.n875 585
R714 B.n874 B.n873 585
R715 B.n872 B.n871 585
R716 B.n870 B.n869 585
R717 B.n868 B.n867 585
R718 B.n866 B.n865 585
R719 B.n864 B.n863 585
R720 B.n862 B.n861 585
R721 B.n860 B.n859 585
R722 B.n858 B.n857 585
R723 B.n856 B.n855 585
R724 B.n854 B.n853 585
R725 B.n852 B.n851 585
R726 B.n850 B.n849 585
R727 B.n848 B.n847 585
R728 B.n846 B.n845 585
R729 B.n844 B.n843 585
R730 B.n842 B.n841 585
R731 B.n840 B.n839 585
R732 B.n838 B.n837 585
R733 B.n836 B.n835 585
R734 B.n834 B.n833 585
R735 B.n832 B.n831 585
R736 B.n830 B.n829 585
R737 B.n828 B.n827 585
R738 B.n826 B.n825 585
R739 B.n824 B.n823 585
R740 B.n822 B.n821 585
R741 B.n820 B.n819 585
R742 B.n818 B.n817 585
R743 B.n816 B.n815 585
R744 B.n814 B.n813 585
R745 B.n812 B.n811 585
R746 B.n810 B.n809 585
R747 B.n808 B.n807 585
R748 B.n806 B.n805 585
R749 B.n804 B.n803 585
R750 B.n802 B.n801 585
R751 B.n800 B.n799 585
R752 B.n798 B.n797 585
R753 B.n796 B.n795 585
R754 B.n794 B.n793 585
R755 B.n792 B.n791 585
R756 B.n790 B.n789 585
R757 B.n788 B.n787 585
R758 B.n786 B.n785 585
R759 B.n784 B.n783 585
R760 B.n782 B.n781 585
R761 B.n780 B.n779 585
R762 B.n778 B.n777 585
R763 B.n776 B.n775 585
R764 B.n774 B.n773 585
R765 B.n772 B.n771 585
R766 B.n770 B.n769 585
R767 B.n768 B.n767 585
R768 B.n766 B.n765 585
R769 B.n764 B.n763 585
R770 B.n762 B.n761 585
R771 B.n760 B.n759 585
R772 B.n758 B.n757 585
R773 B.n756 B.n755 585
R774 B.n754 B.n753 585
R775 B.n752 B.n751 585
R776 B.n750 B.n749 585
R777 B.n748 B.n747 585
R778 B.n746 B.n745 585
R779 B.n744 B.n743 585
R780 B.n742 B.n741 585
R781 B.n740 B.n739 585
R782 B.n738 B.n737 585
R783 B.n736 B.n735 585
R784 B.n734 B.n733 585
R785 B.n732 B.n731 585
R786 B.n730 B.n729 585
R787 B.n728 B.n727 585
R788 B.n726 B.n725 585
R789 B.n724 B.n723 585
R790 B.n722 B.n721 585
R791 B.n720 B.n719 585
R792 B.n718 B.n717 585
R793 B.n716 B.n715 585
R794 B.n714 B.n713 585
R795 B.n712 B.n711 585
R796 B.n710 B.n709 585
R797 B.n708 B.n707 585
R798 B.n706 B.n705 585
R799 B.n704 B.n703 585
R800 B.n702 B.n701 585
R801 B.n700 B.n699 585
R802 B.n698 B.n697 585
R803 B.n696 B.n688 585
R804 B.n970 B.n688 585
R805 B.n974 B.n617 585
R806 B.n617 B.n616 585
R807 B.n976 B.n975 585
R808 B.n977 B.n976 585
R809 B.n611 B.n610 585
R810 B.n612 B.n611 585
R811 B.n985 B.n984 585
R812 B.n984 B.n983 585
R813 B.n986 B.n609 585
R814 B.n609 B.n608 585
R815 B.n988 B.n987 585
R816 B.n989 B.n988 585
R817 B.n603 B.n602 585
R818 B.n604 B.n603 585
R819 B.n998 B.n997 585
R820 B.n997 B.n996 585
R821 B.n999 B.n601 585
R822 B.n995 B.n601 585
R823 B.n1001 B.n1000 585
R824 B.n1002 B.n1001 585
R825 B.n596 B.n595 585
R826 B.n597 B.n596 585
R827 B.n1010 B.n1009 585
R828 B.n1009 B.n1008 585
R829 B.n1011 B.n594 585
R830 B.n594 B.n593 585
R831 B.n1013 B.n1012 585
R832 B.n1014 B.n1013 585
R833 B.n588 B.n587 585
R834 B.n589 B.n588 585
R835 B.n1022 B.n1021 585
R836 B.n1021 B.n1020 585
R837 B.n1023 B.n586 585
R838 B.n586 B.n585 585
R839 B.n1025 B.n1024 585
R840 B.n1026 B.n1025 585
R841 B.n580 B.n579 585
R842 B.n581 B.n580 585
R843 B.n1034 B.n1033 585
R844 B.n1033 B.n1032 585
R845 B.n1035 B.n578 585
R846 B.n578 B.n576 585
R847 B.n1037 B.n1036 585
R848 B.n1038 B.n1037 585
R849 B.n572 B.n571 585
R850 B.n577 B.n572 585
R851 B.n1046 B.n1045 585
R852 B.n1045 B.n1044 585
R853 B.n1047 B.n570 585
R854 B.n570 B.n569 585
R855 B.n1049 B.n1048 585
R856 B.n1050 B.n1049 585
R857 B.n564 B.n563 585
R858 B.n565 B.n564 585
R859 B.n1058 B.n1057 585
R860 B.n1057 B.n1056 585
R861 B.n1059 B.n562 585
R862 B.n562 B.n561 585
R863 B.n1061 B.n1060 585
R864 B.n1062 B.n1061 585
R865 B.n556 B.n555 585
R866 B.n557 B.n556 585
R867 B.n1071 B.n1070 585
R868 B.n1070 B.n1069 585
R869 B.n1072 B.n554 585
R870 B.n1068 B.n554 585
R871 B.n1074 B.n1073 585
R872 B.n1075 B.n1074 585
R873 B.n549 B.n548 585
R874 B.n550 B.n549 585
R875 B.n1083 B.n1082 585
R876 B.n1082 B.n1081 585
R877 B.n1084 B.n547 585
R878 B.n547 B.n546 585
R879 B.n1086 B.n1085 585
R880 B.n1087 B.n1086 585
R881 B.n541 B.n540 585
R882 B.n542 B.n541 585
R883 B.n1095 B.n1094 585
R884 B.n1094 B.n1093 585
R885 B.n1096 B.n539 585
R886 B.n539 B.n538 585
R887 B.n1098 B.n1097 585
R888 B.n1099 B.n1098 585
R889 B.n533 B.n532 585
R890 B.n534 B.n533 585
R891 B.n1107 B.n1106 585
R892 B.n1106 B.n1105 585
R893 B.n1108 B.n531 585
R894 B.n531 B.n530 585
R895 B.n1110 B.n1109 585
R896 B.n1111 B.n1110 585
R897 B.n525 B.n524 585
R898 B.n526 B.n525 585
R899 B.n1119 B.n1118 585
R900 B.n1118 B.n1117 585
R901 B.n1120 B.n523 585
R902 B.n523 B.n522 585
R903 B.n1122 B.n1121 585
R904 B.n1123 B.n1122 585
R905 B.n517 B.n516 585
R906 B.n518 B.n517 585
R907 B.n1131 B.n1130 585
R908 B.n1130 B.n1129 585
R909 B.n1132 B.n515 585
R910 B.n515 B.n513 585
R911 B.n1134 B.n1133 585
R912 B.n1135 B.n1134 585
R913 B.n509 B.n508 585
R914 B.n514 B.n509 585
R915 B.n1143 B.n1142 585
R916 B.n1142 B.n1141 585
R917 B.n1144 B.n507 585
R918 B.n507 B.n506 585
R919 B.n1146 B.n1145 585
R920 B.n1147 B.n1146 585
R921 B.n501 B.n500 585
R922 B.n502 B.n501 585
R923 B.n1155 B.n1154 585
R924 B.n1154 B.n1153 585
R925 B.n1156 B.n499 585
R926 B.n499 B.n498 585
R927 B.n1158 B.n1157 585
R928 B.n1159 B.n1158 585
R929 B.n493 B.n492 585
R930 B.n494 B.n493 585
R931 B.n1168 B.n1167 585
R932 B.n1167 B.n1166 585
R933 B.n1169 B.n491 585
R934 B.n1165 B.n491 585
R935 B.n1171 B.n1170 585
R936 B.n1172 B.n1171 585
R937 B.n486 B.n485 585
R938 B.n487 B.n486 585
R939 B.n1181 B.n1180 585
R940 B.n1180 B.n1179 585
R941 B.n1182 B.n484 585
R942 B.n484 B.n483 585
R943 B.n1184 B.n1183 585
R944 B.n1185 B.n1184 585
R945 B.n3 B.n0 585
R946 B.n4 B.n3 585
R947 B.n1426 B.n1 585
R948 B.n1427 B.n1426 585
R949 B.n1425 B.n1424 585
R950 B.n1425 B.n8 585
R951 B.n1423 B.n9 585
R952 B.n12 B.n9 585
R953 B.n1422 B.n1421 585
R954 B.n1421 B.n1420 585
R955 B.n11 B.n10 585
R956 B.n1419 B.n11 585
R957 B.n1417 B.n1416 585
R958 B.n1418 B.n1417 585
R959 B.n1415 B.n16 585
R960 B.n19 B.n16 585
R961 B.n1414 B.n1413 585
R962 B.n1413 B.n1412 585
R963 B.n18 B.n17 585
R964 B.n1411 B.n18 585
R965 B.n1409 B.n1408 585
R966 B.n1410 B.n1409 585
R967 B.n1407 B.n24 585
R968 B.n24 B.n23 585
R969 B.n1406 B.n1405 585
R970 B.n1405 B.n1404 585
R971 B.n26 B.n25 585
R972 B.n1403 B.n26 585
R973 B.n1401 B.n1400 585
R974 B.n1402 B.n1401 585
R975 B.n1399 B.n31 585
R976 B.n31 B.n30 585
R977 B.n1398 B.n1397 585
R978 B.n1397 B.n1396 585
R979 B.n33 B.n32 585
R980 B.n1395 B.n33 585
R981 B.n1393 B.n1392 585
R982 B.n1394 B.n1393 585
R983 B.n1391 B.n38 585
R984 B.n38 B.n37 585
R985 B.n1390 B.n1389 585
R986 B.n1389 B.n1388 585
R987 B.n40 B.n39 585
R988 B.n1387 B.n40 585
R989 B.n1385 B.n1384 585
R990 B.n1386 B.n1385 585
R991 B.n1383 B.n45 585
R992 B.n45 B.n44 585
R993 B.n1382 B.n1381 585
R994 B.n1381 B.n1380 585
R995 B.n47 B.n46 585
R996 B.n1379 B.n47 585
R997 B.n1377 B.n1376 585
R998 B.n1378 B.n1377 585
R999 B.n1375 B.n52 585
R1000 B.n52 B.n51 585
R1001 B.n1374 B.n1373 585
R1002 B.n1373 B.n1372 585
R1003 B.n54 B.n53 585
R1004 B.n1371 B.n54 585
R1005 B.n1369 B.n1368 585
R1006 B.n1370 B.n1369 585
R1007 B.n1367 B.n59 585
R1008 B.n59 B.n58 585
R1009 B.n1366 B.n1365 585
R1010 B.n1365 B.n1364 585
R1011 B.n61 B.n60 585
R1012 B.n1363 B.n61 585
R1013 B.n1361 B.n1360 585
R1014 B.n1362 B.n1361 585
R1015 B.n1359 B.n66 585
R1016 B.n66 B.n65 585
R1017 B.n1358 B.n1357 585
R1018 B.n1357 B.n1356 585
R1019 B.n68 B.n67 585
R1020 B.n1355 B.n68 585
R1021 B.n1353 B.n1352 585
R1022 B.n1354 B.n1353 585
R1023 B.n1351 B.n72 585
R1024 B.n75 B.n72 585
R1025 B.n1350 B.n1349 585
R1026 B.n1349 B.n1348 585
R1027 B.n74 B.n73 585
R1028 B.n1347 B.n74 585
R1029 B.n1345 B.n1344 585
R1030 B.n1346 B.n1345 585
R1031 B.n1343 B.n80 585
R1032 B.n80 B.n79 585
R1033 B.n1342 B.n1341 585
R1034 B.n1341 B.n1340 585
R1035 B.n82 B.n81 585
R1036 B.n1339 B.n82 585
R1037 B.n1337 B.n1336 585
R1038 B.n1338 B.n1337 585
R1039 B.n1335 B.n87 585
R1040 B.n87 B.n86 585
R1041 B.n1334 B.n1333 585
R1042 B.n1333 B.n1332 585
R1043 B.n89 B.n88 585
R1044 B.n1331 B.n89 585
R1045 B.n1329 B.n1328 585
R1046 B.n1330 B.n1329 585
R1047 B.n1327 B.n94 585
R1048 B.n94 B.n93 585
R1049 B.n1326 B.n1325 585
R1050 B.n1325 B.n1324 585
R1051 B.n96 B.n95 585
R1052 B.n1323 B.n96 585
R1053 B.n1321 B.n1320 585
R1054 B.n1322 B.n1321 585
R1055 B.n1319 B.n101 585
R1056 B.n101 B.n100 585
R1057 B.n1318 B.n1317 585
R1058 B.n1317 B.n1316 585
R1059 B.n103 B.n102 585
R1060 B.n1315 B.n103 585
R1061 B.n1313 B.n1312 585
R1062 B.n1314 B.n1313 585
R1063 B.n1311 B.n108 585
R1064 B.n108 B.n107 585
R1065 B.n1310 B.n1309 585
R1066 B.n1309 B.n1308 585
R1067 B.n110 B.n109 585
R1068 B.n1307 B.n110 585
R1069 B.n1305 B.n1304 585
R1070 B.n1306 B.n1305 585
R1071 B.n1303 B.n114 585
R1072 B.n117 B.n114 585
R1073 B.n1302 B.n1301 585
R1074 B.n1301 B.n1300 585
R1075 B.n116 B.n115 585
R1076 B.n1299 B.n116 585
R1077 B.n1297 B.n1296 585
R1078 B.n1298 B.n1297 585
R1079 B.n1295 B.n122 585
R1080 B.n122 B.n121 585
R1081 B.n1294 B.n1293 585
R1082 B.n1293 B.n1292 585
R1083 B.n124 B.n123 585
R1084 B.n1291 B.n124 585
R1085 B.n1289 B.n1288 585
R1086 B.n1290 B.n1289 585
R1087 B.n1287 B.n129 585
R1088 B.n129 B.n128 585
R1089 B.n1430 B.n1429 585
R1090 B.n1428 B.n2 585
R1091 B.n1285 B.n129 458.866
R1092 B.n1281 B.n201 458.866
R1093 B.n688 B.n615 458.866
R1094 B.n972 B.n617 458.866
R1095 B.n204 B.t10 356.348
R1096 B.n202 B.t17 356.348
R1097 B.n693 B.t6 356.348
R1098 B.n690 B.t14 356.348
R1099 B.n1283 B.n1282 256.663
R1100 B.n1283 B.n199 256.663
R1101 B.n1283 B.n198 256.663
R1102 B.n1283 B.n197 256.663
R1103 B.n1283 B.n196 256.663
R1104 B.n1283 B.n195 256.663
R1105 B.n1283 B.n194 256.663
R1106 B.n1283 B.n193 256.663
R1107 B.n1283 B.n192 256.663
R1108 B.n1283 B.n191 256.663
R1109 B.n1283 B.n190 256.663
R1110 B.n1283 B.n189 256.663
R1111 B.n1283 B.n188 256.663
R1112 B.n1283 B.n187 256.663
R1113 B.n1283 B.n186 256.663
R1114 B.n1283 B.n185 256.663
R1115 B.n1283 B.n184 256.663
R1116 B.n1283 B.n183 256.663
R1117 B.n1283 B.n182 256.663
R1118 B.n1283 B.n181 256.663
R1119 B.n1283 B.n180 256.663
R1120 B.n1283 B.n179 256.663
R1121 B.n1283 B.n178 256.663
R1122 B.n1283 B.n177 256.663
R1123 B.n1283 B.n176 256.663
R1124 B.n1283 B.n175 256.663
R1125 B.n1283 B.n174 256.663
R1126 B.n1283 B.n173 256.663
R1127 B.n1283 B.n172 256.663
R1128 B.n1283 B.n171 256.663
R1129 B.n1283 B.n170 256.663
R1130 B.n1283 B.n169 256.663
R1131 B.n1283 B.n168 256.663
R1132 B.n1283 B.n167 256.663
R1133 B.n1283 B.n166 256.663
R1134 B.n1283 B.n165 256.663
R1135 B.n1283 B.n164 256.663
R1136 B.n1283 B.n163 256.663
R1137 B.n1283 B.n162 256.663
R1138 B.n1283 B.n161 256.663
R1139 B.n1283 B.n160 256.663
R1140 B.n1283 B.n159 256.663
R1141 B.n1283 B.n158 256.663
R1142 B.n1283 B.n157 256.663
R1143 B.n1283 B.n156 256.663
R1144 B.n1283 B.n155 256.663
R1145 B.n1283 B.n154 256.663
R1146 B.n1283 B.n153 256.663
R1147 B.n1283 B.n152 256.663
R1148 B.n1283 B.n151 256.663
R1149 B.n1283 B.n150 256.663
R1150 B.n1283 B.n149 256.663
R1151 B.n1283 B.n148 256.663
R1152 B.n1283 B.n147 256.663
R1153 B.n1283 B.n146 256.663
R1154 B.n1283 B.n145 256.663
R1155 B.n1283 B.n144 256.663
R1156 B.n1283 B.n143 256.663
R1157 B.n1283 B.n142 256.663
R1158 B.n1283 B.n141 256.663
R1159 B.n1283 B.n140 256.663
R1160 B.n1283 B.n139 256.663
R1161 B.n1283 B.n138 256.663
R1162 B.n1283 B.n137 256.663
R1163 B.n1283 B.n136 256.663
R1164 B.n1283 B.n135 256.663
R1165 B.n1283 B.n134 256.663
R1166 B.n1283 B.n133 256.663
R1167 B.n1283 B.n132 256.663
R1168 B.n1284 B.n1283 256.663
R1169 B.n971 B.n970 256.663
R1170 B.n970 B.n620 256.663
R1171 B.n970 B.n621 256.663
R1172 B.n970 B.n622 256.663
R1173 B.n970 B.n623 256.663
R1174 B.n970 B.n624 256.663
R1175 B.n970 B.n625 256.663
R1176 B.n970 B.n626 256.663
R1177 B.n970 B.n627 256.663
R1178 B.n970 B.n628 256.663
R1179 B.n970 B.n629 256.663
R1180 B.n970 B.n630 256.663
R1181 B.n970 B.n631 256.663
R1182 B.n970 B.n632 256.663
R1183 B.n970 B.n633 256.663
R1184 B.n970 B.n634 256.663
R1185 B.n970 B.n635 256.663
R1186 B.n970 B.n636 256.663
R1187 B.n970 B.n637 256.663
R1188 B.n970 B.n638 256.663
R1189 B.n970 B.n639 256.663
R1190 B.n970 B.n640 256.663
R1191 B.n970 B.n641 256.663
R1192 B.n970 B.n642 256.663
R1193 B.n970 B.n643 256.663
R1194 B.n970 B.n644 256.663
R1195 B.n970 B.n645 256.663
R1196 B.n970 B.n646 256.663
R1197 B.n970 B.n647 256.663
R1198 B.n970 B.n648 256.663
R1199 B.n970 B.n649 256.663
R1200 B.n970 B.n650 256.663
R1201 B.n970 B.n651 256.663
R1202 B.n970 B.n652 256.663
R1203 B.n970 B.n653 256.663
R1204 B.n970 B.n654 256.663
R1205 B.n970 B.n655 256.663
R1206 B.n970 B.n656 256.663
R1207 B.n970 B.n657 256.663
R1208 B.n970 B.n658 256.663
R1209 B.n970 B.n659 256.663
R1210 B.n970 B.n660 256.663
R1211 B.n970 B.n661 256.663
R1212 B.n970 B.n662 256.663
R1213 B.n970 B.n663 256.663
R1214 B.n970 B.n664 256.663
R1215 B.n970 B.n665 256.663
R1216 B.n970 B.n666 256.663
R1217 B.n970 B.n667 256.663
R1218 B.n970 B.n668 256.663
R1219 B.n970 B.n669 256.663
R1220 B.n970 B.n670 256.663
R1221 B.n970 B.n671 256.663
R1222 B.n970 B.n672 256.663
R1223 B.n970 B.n673 256.663
R1224 B.n970 B.n674 256.663
R1225 B.n970 B.n675 256.663
R1226 B.n970 B.n676 256.663
R1227 B.n970 B.n677 256.663
R1228 B.n970 B.n678 256.663
R1229 B.n970 B.n679 256.663
R1230 B.n970 B.n680 256.663
R1231 B.n970 B.n681 256.663
R1232 B.n970 B.n682 256.663
R1233 B.n970 B.n683 256.663
R1234 B.n970 B.n684 256.663
R1235 B.n970 B.n685 256.663
R1236 B.n970 B.n686 256.663
R1237 B.n970 B.n687 256.663
R1238 B.n1432 B.n1431 256.663
R1239 B.n206 B.n131 163.367
R1240 B.n210 B.n209 163.367
R1241 B.n214 B.n213 163.367
R1242 B.n218 B.n217 163.367
R1243 B.n222 B.n221 163.367
R1244 B.n226 B.n225 163.367
R1245 B.n230 B.n229 163.367
R1246 B.n234 B.n233 163.367
R1247 B.n238 B.n237 163.367
R1248 B.n242 B.n241 163.367
R1249 B.n246 B.n245 163.367
R1250 B.n250 B.n249 163.367
R1251 B.n254 B.n253 163.367
R1252 B.n258 B.n257 163.367
R1253 B.n262 B.n261 163.367
R1254 B.n266 B.n265 163.367
R1255 B.n270 B.n269 163.367
R1256 B.n274 B.n273 163.367
R1257 B.n278 B.n277 163.367
R1258 B.n282 B.n281 163.367
R1259 B.n286 B.n285 163.367
R1260 B.n290 B.n289 163.367
R1261 B.n294 B.n293 163.367
R1262 B.n298 B.n297 163.367
R1263 B.n302 B.n301 163.367
R1264 B.n306 B.n305 163.367
R1265 B.n310 B.n309 163.367
R1266 B.n314 B.n313 163.367
R1267 B.n318 B.n317 163.367
R1268 B.n322 B.n321 163.367
R1269 B.n326 B.n325 163.367
R1270 B.n330 B.n329 163.367
R1271 B.n335 B.n334 163.367
R1272 B.n339 B.n338 163.367
R1273 B.n343 B.n342 163.367
R1274 B.n347 B.n346 163.367
R1275 B.n351 B.n350 163.367
R1276 B.n356 B.n355 163.367
R1277 B.n360 B.n359 163.367
R1278 B.n364 B.n363 163.367
R1279 B.n368 B.n367 163.367
R1280 B.n372 B.n371 163.367
R1281 B.n376 B.n375 163.367
R1282 B.n380 B.n379 163.367
R1283 B.n384 B.n383 163.367
R1284 B.n388 B.n387 163.367
R1285 B.n392 B.n391 163.367
R1286 B.n396 B.n395 163.367
R1287 B.n400 B.n399 163.367
R1288 B.n404 B.n403 163.367
R1289 B.n408 B.n407 163.367
R1290 B.n412 B.n411 163.367
R1291 B.n416 B.n415 163.367
R1292 B.n420 B.n419 163.367
R1293 B.n424 B.n423 163.367
R1294 B.n428 B.n427 163.367
R1295 B.n432 B.n431 163.367
R1296 B.n436 B.n435 163.367
R1297 B.n440 B.n439 163.367
R1298 B.n444 B.n443 163.367
R1299 B.n448 B.n447 163.367
R1300 B.n452 B.n451 163.367
R1301 B.n456 B.n455 163.367
R1302 B.n460 B.n459 163.367
R1303 B.n464 B.n463 163.367
R1304 B.n468 B.n467 163.367
R1305 B.n472 B.n471 163.367
R1306 B.n476 B.n475 163.367
R1307 B.n478 B.n200 163.367
R1308 B.n978 B.n615 163.367
R1309 B.n978 B.n613 163.367
R1310 B.n982 B.n613 163.367
R1311 B.n982 B.n607 163.367
R1312 B.n990 B.n607 163.367
R1313 B.n990 B.n605 163.367
R1314 B.n994 B.n605 163.367
R1315 B.n994 B.n600 163.367
R1316 B.n1003 B.n600 163.367
R1317 B.n1003 B.n598 163.367
R1318 B.n1007 B.n598 163.367
R1319 B.n1007 B.n592 163.367
R1320 B.n1015 B.n592 163.367
R1321 B.n1015 B.n590 163.367
R1322 B.n1019 B.n590 163.367
R1323 B.n1019 B.n584 163.367
R1324 B.n1027 B.n584 163.367
R1325 B.n1027 B.n582 163.367
R1326 B.n1031 B.n582 163.367
R1327 B.n1031 B.n575 163.367
R1328 B.n1039 B.n575 163.367
R1329 B.n1039 B.n573 163.367
R1330 B.n1043 B.n573 163.367
R1331 B.n1043 B.n568 163.367
R1332 B.n1051 B.n568 163.367
R1333 B.n1051 B.n566 163.367
R1334 B.n1055 B.n566 163.367
R1335 B.n1055 B.n560 163.367
R1336 B.n1063 B.n560 163.367
R1337 B.n1063 B.n558 163.367
R1338 B.n1067 B.n558 163.367
R1339 B.n1067 B.n553 163.367
R1340 B.n1076 B.n553 163.367
R1341 B.n1076 B.n551 163.367
R1342 B.n1080 B.n551 163.367
R1343 B.n1080 B.n545 163.367
R1344 B.n1088 B.n545 163.367
R1345 B.n1088 B.n543 163.367
R1346 B.n1092 B.n543 163.367
R1347 B.n1092 B.n537 163.367
R1348 B.n1100 B.n537 163.367
R1349 B.n1100 B.n535 163.367
R1350 B.n1104 B.n535 163.367
R1351 B.n1104 B.n529 163.367
R1352 B.n1112 B.n529 163.367
R1353 B.n1112 B.n527 163.367
R1354 B.n1116 B.n527 163.367
R1355 B.n1116 B.n521 163.367
R1356 B.n1124 B.n521 163.367
R1357 B.n1124 B.n519 163.367
R1358 B.n1128 B.n519 163.367
R1359 B.n1128 B.n512 163.367
R1360 B.n1136 B.n512 163.367
R1361 B.n1136 B.n510 163.367
R1362 B.n1140 B.n510 163.367
R1363 B.n1140 B.n505 163.367
R1364 B.n1148 B.n505 163.367
R1365 B.n1148 B.n503 163.367
R1366 B.n1152 B.n503 163.367
R1367 B.n1152 B.n497 163.367
R1368 B.n1160 B.n497 163.367
R1369 B.n1160 B.n495 163.367
R1370 B.n1164 B.n495 163.367
R1371 B.n1164 B.n490 163.367
R1372 B.n1173 B.n490 163.367
R1373 B.n1173 B.n488 163.367
R1374 B.n1178 B.n488 163.367
R1375 B.n1178 B.n482 163.367
R1376 B.n1186 B.n482 163.367
R1377 B.n1187 B.n1186 163.367
R1378 B.n1187 B.n5 163.367
R1379 B.n6 B.n5 163.367
R1380 B.n7 B.n6 163.367
R1381 B.n1193 B.n7 163.367
R1382 B.n1194 B.n1193 163.367
R1383 B.n1194 B.n13 163.367
R1384 B.n14 B.n13 163.367
R1385 B.n15 B.n14 163.367
R1386 B.n1199 B.n15 163.367
R1387 B.n1199 B.n20 163.367
R1388 B.n21 B.n20 163.367
R1389 B.n22 B.n21 163.367
R1390 B.n1204 B.n22 163.367
R1391 B.n1204 B.n27 163.367
R1392 B.n28 B.n27 163.367
R1393 B.n29 B.n28 163.367
R1394 B.n1209 B.n29 163.367
R1395 B.n1209 B.n34 163.367
R1396 B.n35 B.n34 163.367
R1397 B.n36 B.n35 163.367
R1398 B.n1214 B.n36 163.367
R1399 B.n1214 B.n41 163.367
R1400 B.n42 B.n41 163.367
R1401 B.n43 B.n42 163.367
R1402 B.n1219 B.n43 163.367
R1403 B.n1219 B.n48 163.367
R1404 B.n49 B.n48 163.367
R1405 B.n50 B.n49 163.367
R1406 B.n1224 B.n50 163.367
R1407 B.n1224 B.n55 163.367
R1408 B.n56 B.n55 163.367
R1409 B.n57 B.n56 163.367
R1410 B.n1229 B.n57 163.367
R1411 B.n1229 B.n62 163.367
R1412 B.n63 B.n62 163.367
R1413 B.n64 B.n63 163.367
R1414 B.n1234 B.n64 163.367
R1415 B.n1234 B.n69 163.367
R1416 B.n70 B.n69 163.367
R1417 B.n71 B.n70 163.367
R1418 B.n1239 B.n71 163.367
R1419 B.n1239 B.n76 163.367
R1420 B.n77 B.n76 163.367
R1421 B.n78 B.n77 163.367
R1422 B.n1244 B.n78 163.367
R1423 B.n1244 B.n83 163.367
R1424 B.n84 B.n83 163.367
R1425 B.n85 B.n84 163.367
R1426 B.n1249 B.n85 163.367
R1427 B.n1249 B.n90 163.367
R1428 B.n91 B.n90 163.367
R1429 B.n92 B.n91 163.367
R1430 B.n1254 B.n92 163.367
R1431 B.n1254 B.n97 163.367
R1432 B.n98 B.n97 163.367
R1433 B.n99 B.n98 163.367
R1434 B.n1259 B.n99 163.367
R1435 B.n1259 B.n104 163.367
R1436 B.n105 B.n104 163.367
R1437 B.n106 B.n105 163.367
R1438 B.n1264 B.n106 163.367
R1439 B.n1264 B.n111 163.367
R1440 B.n112 B.n111 163.367
R1441 B.n113 B.n112 163.367
R1442 B.n1269 B.n113 163.367
R1443 B.n1269 B.n118 163.367
R1444 B.n119 B.n118 163.367
R1445 B.n120 B.n119 163.367
R1446 B.n1274 B.n120 163.367
R1447 B.n1274 B.n125 163.367
R1448 B.n126 B.n125 163.367
R1449 B.n127 B.n126 163.367
R1450 B.n201 B.n127 163.367
R1451 B.n969 B.n619 163.367
R1452 B.n969 B.n689 163.367
R1453 B.n965 B.n964 163.367
R1454 B.n961 B.n960 163.367
R1455 B.n957 B.n956 163.367
R1456 B.n953 B.n952 163.367
R1457 B.n949 B.n948 163.367
R1458 B.n945 B.n944 163.367
R1459 B.n941 B.n940 163.367
R1460 B.n937 B.n936 163.367
R1461 B.n933 B.n932 163.367
R1462 B.n929 B.n928 163.367
R1463 B.n925 B.n924 163.367
R1464 B.n921 B.n920 163.367
R1465 B.n917 B.n916 163.367
R1466 B.n913 B.n912 163.367
R1467 B.n909 B.n908 163.367
R1468 B.n905 B.n904 163.367
R1469 B.n901 B.n900 163.367
R1470 B.n897 B.n896 163.367
R1471 B.n893 B.n892 163.367
R1472 B.n889 B.n888 163.367
R1473 B.n885 B.n884 163.367
R1474 B.n881 B.n880 163.367
R1475 B.n877 B.n876 163.367
R1476 B.n873 B.n872 163.367
R1477 B.n869 B.n868 163.367
R1478 B.n865 B.n864 163.367
R1479 B.n861 B.n860 163.367
R1480 B.n857 B.n856 163.367
R1481 B.n853 B.n852 163.367
R1482 B.n849 B.n848 163.367
R1483 B.n845 B.n844 163.367
R1484 B.n841 B.n840 163.367
R1485 B.n837 B.n836 163.367
R1486 B.n833 B.n832 163.367
R1487 B.n829 B.n828 163.367
R1488 B.n825 B.n824 163.367
R1489 B.n821 B.n820 163.367
R1490 B.n817 B.n816 163.367
R1491 B.n813 B.n812 163.367
R1492 B.n809 B.n808 163.367
R1493 B.n805 B.n804 163.367
R1494 B.n801 B.n800 163.367
R1495 B.n797 B.n796 163.367
R1496 B.n793 B.n792 163.367
R1497 B.n789 B.n788 163.367
R1498 B.n785 B.n784 163.367
R1499 B.n781 B.n780 163.367
R1500 B.n777 B.n776 163.367
R1501 B.n773 B.n772 163.367
R1502 B.n769 B.n768 163.367
R1503 B.n765 B.n764 163.367
R1504 B.n761 B.n760 163.367
R1505 B.n757 B.n756 163.367
R1506 B.n753 B.n752 163.367
R1507 B.n749 B.n748 163.367
R1508 B.n745 B.n744 163.367
R1509 B.n741 B.n740 163.367
R1510 B.n737 B.n736 163.367
R1511 B.n733 B.n732 163.367
R1512 B.n729 B.n728 163.367
R1513 B.n725 B.n724 163.367
R1514 B.n721 B.n720 163.367
R1515 B.n717 B.n716 163.367
R1516 B.n713 B.n712 163.367
R1517 B.n709 B.n708 163.367
R1518 B.n705 B.n704 163.367
R1519 B.n701 B.n700 163.367
R1520 B.n697 B.n688 163.367
R1521 B.n976 B.n617 163.367
R1522 B.n976 B.n611 163.367
R1523 B.n984 B.n611 163.367
R1524 B.n984 B.n609 163.367
R1525 B.n988 B.n609 163.367
R1526 B.n988 B.n603 163.367
R1527 B.n997 B.n603 163.367
R1528 B.n997 B.n601 163.367
R1529 B.n1001 B.n601 163.367
R1530 B.n1001 B.n596 163.367
R1531 B.n1009 B.n596 163.367
R1532 B.n1009 B.n594 163.367
R1533 B.n1013 B.n594 163.367
R1534 B.n1013 B.n588 163.367
R1535 B.n1021 B.n588 163.367
R1536 B.n1021 B.n586 163.367
R1537 B.n1025 B.n586 163.367
R1538 B.n1025 B.n580 163.367
R1539 B.n1033 B.n580 163.367
R1540 B.n1033 B.n578 163.367
R1541 B.n1037 B.n578 163.367
R1542 B.n1037 B.n572 163.367
R1543 B.n1045 B.n572 163.367
R1544 B.n1045 B.n570 163.367
R1545 B.n1049 B.n570 163.367
R1546 B.n1049 B.n564 163.367
R1547 B.n1057 B.n564 163.367
R1548 B.n1057 B.n562 163.367
R1549 B.n1061 B.n562 163.367
R1550 B.n1061 B.n556 163.367
R1551 B.n1070 B.n556 163.367
R1552 B.n1070 B.n554 163.367
R1553 B.n1074 B.n554 163.367
R1554 B.n1074 B.n549 163.367
R1555 B.n1082 B.n549 163.367
R1556 B.n1082 B.n547 163.367
R1557 B.n1086 B.n547 163.367
R1558 B.n1086 B.n541 163.367
R1559 B.n1094 B.n541 163.367
R1560 B.n1094 B.n539 163.367
R1561 B.n1098 B.n539 163.367
R1562 B.n1098 B.n533 163.367
R1563 B.n1106 B.n533 163.367
R1564 B.n1106 B.n531 163.367
R1565 B.n1110 B.n531 163.367
R1566 B.n1110 B.n525 163.367
R1567 B.n1118 B.n525 163.367
R1568 B.n1118 B.n523 163.367
R1569 B.n1122 B.n523 163.367
R1570 B.n1122 B.n517 163.367
R1571 B.n1130 B.n517 163.367
R1572 B.n1130 B.n515 163.367
R1573 B.n1134 B.n515 163.367
R1574 B.n1134 B.n509 163.367
R1575 B.n1142 B.n509 163.367
R1576 B.n1142 B.n507 163.367
R1577 B.n1146 B.n507 163.367
R1578 B.n1146 B.n501 163.367
R1579 B.n1154 B.n501 163.367
R1580 B.n1154 B.n499 163.367
R1581 B.n1158 B.n499 163.367
R1582 B.n1158 B.n493 163.367
R1583 B.n1167 B.n493 163.367
R1584 B.n1167 B.n491 163.367
R1585 B.n1171 B.n491 163.367
R1586 B.n1171 B.n486 163.367
R1587 B.n1180 B.n486 163.367
R1588 B.n1180 B.n484 163.367
R1589 B.n1184 B.n484 163.367
R1590 B.n1184 B.n3 163.367
R1591 B.n1430 B.n3 163.367
R1592 B.n1426 B.n2 163.367
R1593 B.n1426 B.n1425 163.367
R1594 B.n1425 B.n9 163.367
R1595 B.n1421 B.n9 163.367
R1596 B.n1421 B.n11 163.367
R1597 B.n1417 B.n11 163.367
R1598 B.n1417 B.n16 163.367
R1599 B.n1413 B.n16 163.367
R1600 B.n1413 B.n18 163.367
R1601 B.n1409 B.n18 163.367
R1602 B.n1409 B.n24 163.367
R1603 B.n1405 B.n24 163.367
R1604 B.n1405 B.n26 163.367
R1605 B.n1401 B.n26 163.367
R1606 B.n1401 B.n31 163.367
R1607 B.n1397 B.n31 163.367
R1608 B.n1397 B.n33 163.367
R1609 B.n1393 B.n33 163.367
R1610 B.n1393 B.n38 163.367
R1611 B.n1389 B.n38 163.367
R1612 B.n1389 B.n40 163.367
R1613 B.n1385 B.n40 163.367
R1614 B.n1385 B.n45 163.367
R1615 B.n1381 B.n45 163.367
R1616 B.n1381 B.n47 163.367
R1617 B.n1377 B.n47 163.367
R1618 B.n1377 B.n52 163.367
R1619 B.n1373 B.n52 163.367
R1620 B.n1373 B.n54 163.367
R1621 B.n1369 B.n54 163.367
R1622 B.n1369 B.n59 163.367
R1623 B.n1365 B.n59 163.367
R1624 B.n1365 B.n61 163.367
R1625 B.n1361 B.n61 163.367
R1626 B.n1361 B.n66 163.367
R1627 B.n1357 B.n66 163.367
R1628 B.n1357 B.n68 163.367
R1629 B.n1353 B.n68 163.367
R1630 B.n1353 B.n72 163.367
R1631 B.n1349 B.n72 163.367
R1632 B.n1349 B.n74 163.367
R1633 B.n1345 B.n74 163.367
R1634 B.n1345 B.n80 163.367
R1635 B.n1341 B.n80 163.367
R1636 B.n1341 B.n82 163.367
R1637 B.n1337 B.n82 163.367
R1638 B.n1337 B.n87 163.367
R1639 B.n1333 B.n87 163.367
R1640 B.n1333 B.n89 163.367
R1641 B.n1329 B.n89 163.367
R1642 B.n1329 B.n94 163.367
R1643 B.n1325 B.n94 163.367
R1644 B.n1325 B.n96 163.367
R1645 B.n1321 B.n96 163.367
R1646 B.n1321 B.n101 163.367
R1647 B.n1317 B.n101 163.367
R1648 B.n1317 B.n103 163.367
R1649 B.n1313 B.n103 163.367
R1650 B.n1313 B.n108 163.367
R1651 B.n1309 B.n108 163.367
R1652 B.n1309 B.n110 163.367
R1653 B.n1305 B.n110 163.367
R1654 B.n1305 B.n114 163.367
R1655 B.n1301 B.n114 163.367
R1656 B.n1301 B.n116 163.367
R1657 B.n1297 B.n116 163.367
R1658 B.n1297 B.n122 163.367
R1659 B.n1293 B.n122 163.367
R1660 B.n1293 B.n124 163.367
R1661 B.n1289 B.n124 163.367
R1662 B.n1289 B.n129 163.367
R1663 B.n202 B.t18 141.228
R1664 B.n693 B.t9 141.228
R1665 B.n204 B.t12 141.202
R1666 B.n690 B.t16 141.202
R1667 B.n1285 B.n1284 71.676
R1668 B.n206 B.n132 71.676
R1669 B.n210 B.n133 71.676
R1670 B.n214 B.n134 71.676
R1671 B.n218 B.n135 71.676
R1672 B.n222 B.n136 71.676
R1673 B.n226 B.n137 71.676
R1674 B.n230 B.n138 71.676
R1675 B.n234 B.n139 71.676
R1676 B.n238 B.n140 71.676
R1677 B.n242 B.n141 71.676
R1678 B.n246 B.n142 71.676
R1679 B.n250 B.n143 71.676
R1680 B.n254 B.n144 71.676
R1681 B.n258 B.n145 71.676
R1682 B.n262 B.n146 71.676
R1683 B.n266 B.n147 71.676
R1684 B.n270 B.n148 71.676
R1685 B.n274 B.n149 71.676
R1686 B.n278 B.n150 71.676
R1687 B.n282 B.n151 71.676
R1688 B.n286 B.n152 71.676
R1689 B.n290 B.n153 71.676
R1690 B.n294 B.n154 71.676
R1691 B.n298 B.n155 71.676
R1692 B.n302 B.n156 71.676
R1693 B.n306 B.n157 71.676
R1694 B.n310 B.n158 71.676
R1695 B.n314 B.n159 71.676
R1696 B.n318 B.n160 71.676
R1697 B.n322 B.n161 71.676
R1698 B.n326 B.n162 71.676
R1699 B.n330 B.n163 71.676
R1700 B.n335 B.n164 71.676
R1701 B.n339 B.n165 71.676
R1702 B.n343 B.n166 71.676
R1703 B.n347 B.n167 71.676
R1704 B.n351 B.n168 71.676
R1705 B.n356 B.n169 71.676
R1706 B.n360 B.n170 71.676
R1707 B.n364 B.n171 71.676
R1708 B.n368 B.n172 71.676
R1709 B.n372 B.n173 71.676
R1710 B.n376 B.n174 71.676
R1711 B.n380 B.n175 71.676
R1712 B.n384 B.n176 71.676
R1713 B.n388 B.n177 71.676
R1714 B.n392 B.n178 71.676
R1715 B.n396 B.n179 71.676
R1716 B.n400 B.n180 71.676
R1717 B.n404 B.n181 71.676
R1718 B.n408 B.n182 71.676
R1719 B.n412 B.n183 71.676
R1720 B.n416 B.n184 71.676
R1721 B.n420 B.n185 71.676
R1722 B.n424 B.n186 71.676
R1723 B.n428 B.n187 71.676
R1724 B.n432 B.n188 71.676
R1725 B.n436 B.n189 71.676
R1726 B.n440 B.n190 71.676
R1727 B.n444 B.n191 71.676
R1728 B.n448 B.n192 71.676
R1729 B.n452 B.n193 71.676
R1730 B.n456 B.n194 71.676
R1731 B.n460 B.n195 71.676
R1732 B.n464 B.n196 71.676
R1733 B.n468 B.n197 71.676
R1734 B.n472 B.n198 71.676
R1735 B.n476 B.n199 71.676
R1736 B.n1282 B.n200 71.676
R1737 B.n1282 B.n1281 71.676
R1738 B.n478 B.n199 71.676
R1739 B.n475 B.n198 71.676
R1740 B.n471 B.n197 71.676
R1741 B.n467 B.n196 71.676
R1742 B.n463 B.n195 71.676
R1743 B.n459 B.n194 71.676
R1744 B.n455 B.n193 71.676
R1745 B.n451 B.n192 71.676
R1746 B.n447 B.n191 71.676
R1747 B.n443 B.n190 71.676
R1748 B.n439 B.n189 71.676
R1749 B.n435 B.n188 71.676
R1750 B.n431 B.n187 71.676
R1751 B.n427 B.n186 71.676
R1752 B.n423 B.n185 71.676
R1753 B.n419 B.n184 71.676
R1754 B.n415 B.n183 71.676
R1755 B.n411 B.n182 71.676
R1756 B.n407 B.n181 71.676
R1757 B.n403 B.n180 71.676
R1758 B.n399 B.n179 71.676
R1759 B.n395 B.n178 71.676
R1760 B.n391 B.n177 71.676
R1761 B.n387 B.n176 71.676
R1762 B.n383 B.n175 71.676
R1763 B.n379 B.n174 71.676
R1764 B.n375 B.n173 71.676
R1765 B.n371 B.n172 71.676
R1766 B.n367 B.n171 71.676
R1767 B.n363 B.n170 71.676
R1768 B.n359 B.n169 71.676
R1769 B.n355 B.n168 71.676
R1770 B.n350 B.n167 71.676
R1771 B.n346 B.n166 71.676
R1772 B.n342 B.n165 71.676
R1773 B.n338 B.n164 71.676
R1774 B.n334 B.n163 71.676
R1775 B.n329 B.n162 71.676
R1776 B.n325 B.n161 71.676
R1777 B.n321 B.n160 71.676
R1778 B.n317 B.n159 71.676
R1779 B.n313 B.n158 71.676
R1780 B.n309 B.n157 71.676
R1781 B.n305 B.n156 71.676
R1782 B.n301 B.n155 71.676
R1783 B.n297 B.n154 71.676
R1784 B.n293 B.n153 71.676
R1785 B.n289 B.n152 71.676
R1786 B.n285 B.n151 71.676
R1787 B.n281 B.n150 71.676
R1788 B.n277 B.n149 71.676
R1789 B.n273 B.n148 71.676
R1790 B.n269 B.n147 71.676
R1791 B.n265 B.n146 71.676
R1792 B.n261 B.n145 71.676
R1793 B.n257 B.n144 71.676
R1794 B.n253 B.n143 71.676
R1795 B.n249 B.n142 71.676
R1796 B.n245 B.n141 71.676
R1797 B.n241 B.n140 71.676
R1798 B.n237 B.n139 71.676
R1799 B.n233 B.n138 71.676
R1800 B.n229 B.n137 71.676
R1801 B.n225 B.n136 71.676
R1802 B.n221 B.n135 71.676
R1803 B.n217 B.n134 71.676
R1804 B.n213 B.n133 71.676
R1805 B.n209 B.n132 71.676
R1806 B.n1284 B.n131 71.676
R1807 B.n972 B.n971 71.676
R1808 B.n689 B.n620 71.676
R1809 B.n964 B.n621 71.676
R1810 B.n960 B.n622 71.676
R1811 B.n956 B.n623 71.676
R1812 B.n952 B.n624 71.676
R1813 B.n948 B.n625 71.676
R1814 B.n944 B.n626 71.676
R1815 B.n940 B.n627 71.676
R1816 B.n936 B.n628 71.676
R1817 B.n932 B.n629 71.676
R1818 B.n928 B.n630 71.676
R1819 B.n924 B.n631 71.676
R1820 B.n920 B.n632 71.676
R1821 B.n916 B.n633 71.676
R1822 B.n912 B.n634 71.676
R1823 B.n908 B.n635 71.676
R1824 B.n904 B.n636 71.676
R1825 B.n900 B.n637 71.676
R1826 B.n896 B.n638 71.676
R1827 B.n892 B.n639 71.676
R1828 B.n888 B.n640 71.676
R1829 B.n884 B.n641 71.676
R1830 B.n880 B.n642 71.676
R1831 B.n876 B.n643 71.676
R1832 B.n872 B.n644 71.676
R1833 B.n868 B.n645 71.676
R1834 B.n864 B.n646 71.676
R1835 B.n860 B.n647 71.676
R1836 B.n856 B.n648 71.676
R1837 B.n852 B.n649 71.676
R1838 B.n848 B.n650 71.676
R1839 B.n844 B.n651 71.676
R1840 B.n840 B.n652 71.676
R1841 B.n836 B.n653 71.676
R1842 B.n832 B.n654 71.676
R1843 B.n828 B.n655 71.676
R1844 B.n824 B.n656 71.676
R1845 B.n820 B.n657 71.676
R1846 B.n816 B.n658 71.676
R1847 B.n812 B.n659 71.676
R1848 B.n808 B.n660 71.676
R1849 B.n804 B.n661 71.676
R1850 B.n800 B.n662 71.676
R1851 B.n796 B.n663 71.676
R1852 B.n792 B.n664 71.676
R1853 B.n788 B.n665 71.676
R1854 B.n784 B.n666 71.676
R1855 B.n780 B.n667 71.676
R1856 B.n776 B.n668 71.676
R1857 B.n772 B.n669 71.676
R1858 B.n768 B.n670 71.676
R1859 B.n764 B.n671 71.676
R1860 B.n760 B.n672 71.676
R1861 B.n756 B.n673 71.676
R1862 B.n752 B.n674 71.676
R1863 B.n748 B.n675 71.676
R1864 B.n744 B.n676 71.676
R1865 B.n740 B.n677 71.676
R1866 B.n736 B.n678 71.676
R1867 B.n732 B.n679 71.676
R1868 B.n728 B.n680 71.676
R1869 B.n724 B.n681 71.676
R1870 B.n720 B.n682 71.676
R1871 B.n716 B.n683 71.676
R1872 B.n712 B.n684 71.676
R1873 B.n708 B.n685 71.676
R1874 B.n704 B.n686 71.676
R1875 B.n700 B.n687 71.676
R1876 B.n971 B.n619 71.676
R1877 B.n965 B.n620 71.676
R1878 B.n961 B.n621 71.676
R1879 B.n957 B.n622 71.676
R1880 B.n953 B.n623 71.676
R1881 B.n949 B.n624 71.676
R1882 B.n945 B.n625 71.676
R1883 B.n941 B.n626 71.676
R1884 B.n937 B.n627 71.676
R1885 B.n933 B.n628 71.676
R1886 B.n929 B.n629 71.676
R1887 B.n925 B.n630 71.676
R1888 B.n921 B.n631 71.676
R1889 B.n917 B.n632 71.676
R1890 B.n913 B.n633 71.676
R1891 B.n909 B.n634 71.676
R1892 B.n905 B.n635 71.676
R1893 B.n901 B.n636 71.676
R1894 B.n897 B.n637 71.676
R1895 B.n893 B.n638 71.676
R1896 B.n889 B.n639 71.676
R1897 B.n885 B.n640 71.676
R1898 B.n881 B.n641 71.676
R1899 B.n877 B.n642 71.676
R1900 B.n873 B.n643 71.676
R1901 B.n869 B.n644 71.676
R1902 B.n865 B.n645 71.676
R1903 B.n861 B.n646 71.676
R1904 B.n857 B.n647 71.676
R1905 B.n853 B.n648 71.676
R1906 B.n849 B.n649 71.676
R1907 B.n845 B.n650 71.676
R1908 B.n841 B.n651 71.676
R1909 B.n837 B.n652 71.676
R1910 B.n833 B.n653 71.676
R1911 B.n829 B.n654 71.676
R1912 B.n825 B.n655 71.676
R1913 B.n821 B.n656 71.676
R1914 B.n817 B.n657 71.676
R1915 B.n813 B.n658 71.676
R1916 B.n809 B.n659 71.676
R1917 B.n805 B.n660 71.676
R1918 B.n801 B.n661 71.676
R1919 B.n797 B.n662 71.676
R1920 B.n793 B.n663 71.676
R1921 B.n789 B.n664 71.676
R1922 B.n785 B.n665 71.676
R1923 B.n781 B.n666 71.676
R1924 B.n777 B.n667 71.676
R1925 B.n773 B.n668 71.676
R1926 B.n769 B.n669 71.676
R1927 B.n765 B.n670 71.676
R1928 B.n761 B.n671 71.676
R1929 B.n757 B.n672 71.676
R1930 B.n753 B.n673 71.676
R1931 B.n749 B.n674 71.676
R1932 B.n745 B.n675 71.676
R1933 B.n741 B.n676 71.676
R1934 B.n737 B.n677 71.676
R1935 B.n733 B.n678 71.676
R1936 B.n729 B.n679 71.676
R1937 B.n725 B.n680 71.676
R1938 B.n721 B.n681 71.676
R1939 B.n717 B.n682 71.676
R1940 B.n713 B.n683 71.676
R1941 B.n709 B.n684 71.676
R1942 B.n705 B.n685 71.676
R1943 B.n701 B.n686 71.676
R1944 B.n697 B.n687 71.676
R1945 B.n1431 B.n1430 71.676
R1946 B.n1431 B.n2 71.676
R1947 B.n203 B.t19 71.6045
R1948 B.n694 B.t8 71.6045
R1949 B.n205 B.t13 71.5777
R1950 B.n691 B.t15 71.5777
R1951 B.n205 B.n204 69.6247
R1952 B.n203 B.n202 69.6247
R1953 B.n694 B.n693 69.6247
R1954 B.n691 B.n690 69.6247
R1955 B.n332 B.n205 59.5399
R1956 B.n353 B.n203 59.5399
R1957 B.n695 B.n694 59.5399
R1958 B.n692 B.n691 59.5399
R1959 B.n970 B.n616 52.7656
R1960 B.n1283 B.n128 52.7656
R1961 B.n1280 B.n1279 29.8151
R1962 B.n974 B.n973 29.8151
R1963 B.n696 B.n614 29.8151
R1964 B.n1287 B.n1286 29.8151
R1965 B.n977 B.n616 29.6536
R1966 B.n977 B.n612 29.6536
R1967 B.n983 B.n612 29.6536
R1968 B.n983 B.n608 29.6536
R1969 B.n989 B.n608 29.6536
R1970 B.n989 B.n604 29.6536
R1971 B.n996 B.n604 29.6536
R1972 B.n996 B.n995 29.6536
R1973 B.n1002 B.n597 29.6536
R1974 B.n1008 B.n597 29.6536
R1975 B.n1008 B.n593 29.6536
R1976 B.n1014 B.n593 29.6536
R1977 B.n1014 B.n589 29.6536
R1978 B.n1020 B.n589 29.6536
R1979 B.n1020 B.n585 29.6536
R1980 B.n1026 B.n585 29.6536
R1981 B.n1026 B.n581 29.6536
R1982 B.n1032 B.n581 29.6536
R1983 B.n1032 B.n576 29.6536
R1984 B.n1038 B.n576 29.6536
R1985 B.n1038 B.n577 29.6536
R1986 B.n1044 B.n569 29.6536
R1987 B.n1050 B.n569 29.6536
R1988 B.n1050 B.n565 29.6536
R1989 B.n1056 B.n565 29.6536
R1990 B.n1056 B.n561 29.6536
R1991 B.n1062 B.n561 29.6536
R1992 B.n1062 B.n557 29.6536
R1993 B.n1069 B.n557 29.6536
R1994 B.n1069 B.n1068 29.6536
R1995 B.n1075 B.n550 29.6536
R1996 B.n1081 B.n550 29.6536
R1997 B.n1081 B.n546 29.6536
R1998 B.n1087 B.n546 29.6536
R1999 B.n1087 B.n542 29.6536
R2000 B.n1093 B.n542 29.6536
R2001 B.n1093 B.n538 29.6536
R2002 B.n1099 B.n538 29.6536
R2003 B.n1099 B.n534 29.6536
R2004 B.n1105 B.n534 29.6536
R2005 B.n1111 B.n530 29.6536
R2006 B.n1111 B.n526 29.6536
R2007 B.n1117 B.n526 29.6536
R2008 B.n1117 B.n522 29.6536
R2009 B.n1123 B.n522 29.6536
R2010 B.n1123 B.n518 29.6536
R2011 B.n1129 B.n518 29.6536
R2012 B.n1129 B.n513 29.6536
R2013 B.n1135 B.n513 29.6536
R2014 B.n1135 B.n514 29.6536
R2015 B.n1141 B.n506 29.6536
R2016 B.n1147 B.n506 29.6536
R2017 B.n1147 B.n502 29.6536
R2018 B.n1153 B.n502 29.6536
R2019 B.n1153 B.n498 29.6536
R2020 B.n1159 B.n498 29.6536
R2021 B.n1159 B.n494 29.6536
R2022 B.n1166 B.n494 29.6536
R2023 B.n1166 B.n1165 29.6536
R2024 B.n1172 B.n487 29.6536
R2025 B.n1179 B.n487 29.6536
R2026 B.n1179 B.n483 29.6536
R2027 B.n1185 B.n483 29.6536
R2028 B.n1185 B.n4 29.6536
R2029 B.n1429 B.n4 29.6536
R2030 B.n1429 B.n1428 29.6536
R2031 B.n1428 B.n1427 29.6536
R2032 B.n1427 B.n8 29.6536
R2033 B.n12 B.n8 29.6536
R2034 B.n1420 B.n12 29.6536
R2035 B.n1420 B.n1419 29.6536
R2036 B.n1419 B.n1418 29.6536
R2037 B.n1412 B.n19 29.6536
R2038 B.n1412 B.n1411 29.6536
R2039 B.n1411 B.n1410 29.6536
R2040 B.n1410 B.n23 29.6536
R2041 B.n1404 B.n23 29.6536
R2042 B.n1404 B.n1403 29.6536
R2043 B.n1403 B.n1402 29.6536
R2044 B.n1402 B.n30 29.6536
R2045 B.n1396 B.n30 29.6536
R2046 B.n1395 B.n1394 29.6536
R2047 B.n1394 B.n37 29.6536
R2048 B.n1388 B.n37 29.6536
R2049 B.n1388 B.n1387 29.6536
R2050 B.n1387 B.n1386 29.6536
R2051 B.n1386 B.n44 29.6536
R2052 B.n1380 B.n44 29.6536
R2053 B.n1380 B.n1379 29.6536
R2054 B.n1379 B.n1378 29.6536
R2055 B.n1378 B.n51 29.6536
R2056 B.n1372 B.n1371 29.6536
R2057 B.n1371 B.n1370 29.6536
R2058 B.n1370 B.n58 29.6536
R2059 B.n1364 B.n58 29.6536
R2060 B.n1364 B.n1363 29.6536
R2061 B.n1363 B.n1362 29.6536
R2062 B.n1362 B.n65 29.6536
R2063 B.n1356 B.n65 29.6536
R2064 B.n1356 B.n1355 29.6536
R2065 B.n1355 B.n1354 29.6536
R2066 B.n1348 B.n75 29.6536
R2067 B.n1348 B.n1347 29.6536
R2068 B.n1347 B.n1346 29.6536
R2069 B.n1346 B.n79 29.6536
R2070 B.n1340 B.n79 29.6536
R2071 B.n1340 B.n1339 29.6536
R2072 B.n1339 B.n1338 29.6536
R2073 B.n1338 B.n86 29.6536
R2074 B.n1332 B.n86 29.6536
R2075 B.n1331 B.n1330 29.6536
R2076 B.n1330 B.n93 29.6536
R2077 B.n1324 B.n93 29.6536
R2078 B.n1324 B.n1323 29.6536
R2079 B.n1323 B.n1322 29.6536
R2080 B.n1322 B.n100 29.6536
R2081 B.n1316 B.n100 29.6536
R2082 B.n1316 B.n1315 29.6536
R2083 B.n1315 B.n1314 29.6536
R2084 B.n1314 B.n107 29.6536
R2085 B.n1308 B.n107 29.6536
R2086 B.n1308 B.n1307 29.6536
R2087 B.n1307 B.n1306 29.6536
R2088 B.n1300 B.n117 29.6536
R2089 B.n1300 B.n1299 29.6536
R2090 B.n1299 B.n1298 29.6536
R2091 B.n1298 B.n121 29.6536
R2092 B.n1292 B.n121 29.6536
R2093 B.n1292 B.n1291 29.6536
R2094 B.n1291 B.n1290 29.6536
R2095 B.n1290 B.n128 29.6536
R2096 B.n1068 B.t21 27.9093
R2097 B.n1141 B.t5 27.9093
R2098 B.n1396 B.t23 27.9093
R2099 B.n75 B.t20 27.9093
R2100 B.n995 B.t7 18.3157
R2101 B.n1044 B.t2 18.3157
R2102 B.n1165 B.t0 18.3157
R2103 B.n19 B.t1 18.3157
R2104 B.n1332 B.t22 18.3157
R2105 B.n117 B.t11 18.3157
R2106 B B.n1432 18.0485
R2107 B.n1105 B.t4 14.8271
R2108 B.t4 B.n530 14.8271
R2109 B.t3 B.n51 14.8271
R2110 B.n1372 B.t3 14.8271
R2111 B.n1002 B.t7 11.3385
R2112 B.n577 B.t2 11.3385
R2113 B.n1172 B.t0 11.3385
R2114 B.n1418 B.t1 11.3385
R2115 B.t22 B.n1331 11.3385
R2116 B.n1306 B.t11 11.3385
R2117 B.n975 B.n974 10.6151
R2118 B.n975 B.n610 10.6151
R2119 B.n985 B.n610 10.6151
R2120 B.n986 B.n985 10.6151
R2121 B.n987 B.n986 10.6151
R2122 B.n987 B.n602 10.6151
R2123 B.n998 B.n602 10.6151
R2124 B.n999 B.n998 10.6151
R2125 B.n1000 B.n999 10.6151
R2126 B.n1000 B.n595 10.6151
R2127 B.n1010 B.n595 10.6151
R2128 B.n1011 B.n1010 10.6151
R2129 B.n1012 B.n1011 10.6151
R2130 B.n1012 B.n587 10.6151
R2131 B.n1022 B.n587 10.6151
R2132 B.n1023 B.n1022 10.6151
R2133 B.n1024 B.n1023 10.6151
R2134 B.n1024 B.n579 10.6151
R2135 B.n1034 B.n579 10.6151
R2136 B.n1035 B.n1034 10.6151
R2137 B.n1036 B.n1035 10.6151
R2138 B.n1036 B.n571 10.6151
R2139 B.n1046 B.n571 10.6151
R2140 B.n1047 B.n1046 10.6151
R2141 B.n1048 B.n1047 10.6151
R2142 B.n1048 B.n563 10.6151
R2143 B.n1058 B.n563 10.6151
R2144 B.n1059 B.n1058 10.6151
R2145 B.n1060 B.n1059 10.6151
R2146 B.n1060 B.n555 10.6151
R2147 B.n1071 B.n555 10.6151
R2148 B.n1072 B.n1071 10.6151
R2149 B.n1073 B.n1072 10.6151
R2150 B.n1073 B.n548 10.6151
R2151 B.n1083 B.n548 10.6151
R2152 B.n1084 B.n1083 10.6151
R2153 B.n1085 B.n1084 10.6151
R2154 B.n1085 B.n540 10.6151
R2155 B.n1095 B.n540 10.6151
R2156 B.n1096 B.n1095 10.6151
R2157 B.n1097 B.n1096 10.6151
R2158 B.n1097 B.n532 10.6151
R2159 B.n1107 B.n532 10.6151
R2160 B.n1108 B.n1107 10.6151
R2161 B.n1109 B.n1108 10.6151
R2162 B.n1109 B.n524 10.6151
R2163 B.n1119 B.n524 10.6151
R2164 B.n1120 B.n1119 10.6151
R2165 B.n1121 B.n1120 10.6151
R2166 B.n1121 B.n516 10.6151
R2167 B.n1131 B.n516 10.6151
R2168 B.n1132 B.n1131 10.6151
R2169 B.n1133 B.n1132 10.6151
R2170 B.n1133 B.n508 10.6151
R2171 B.n1143 B.n508 10.6151
R2172 B.n1144 B.n1143 10.6151
R2173 B.n1145 B.n1144 10.6151
R2174 B.n1145 B.n500 10.6151
R2175 B.n1155 B.n500 10.6151
R2176 B.n1156 B.n1155 10.6151
R2177 B.n1157 B.n1156 10.6151
R2178 B.n1157 B.n492 10.6151
R2179 B.n1168 B.n492 10.6151
R2180 B.n1169 B.n1168 10.6151
R2181 B.n1170 B.n1169 10.6151
R2182 B.n1170 B.n485 10.6151
R2183 B.n1181 B.n485 10.6151
R2184 B.n1182 B.n1181 10.6151
R2185 B.n1183 B.n1182 10.6151
R2186 B.n1183 B.n0 10.6151
R2187 B.n973 B.n618 10.6151
R2188 B.n968 B.n618 10.6151
R2189 B.n968 B.n967 10.6151
R2190 B.n967 B.n966 10.6151
R2191 B.n966 B.n963 10.6151
R2192 B.n963 B.n962 10.6151
R2193 B.n962 B.n959 10.6151
R2194 B.n959 B.n958 10.6151
R2195 B.n958 B.n955 10.6151
R2196 B.n955 B.n954 10.6151
R2197 B.n954 B.n951 10.6151
R2198 B.n951 B.n950 10.6151
R2199 B.n950 B.n947 10.6151
R2200 B.n947 B.n946 10.6151
R2201 B.n946 B.n943 10.6151
R2202 B.n943 B.n942 10.6151
R2203 B.n942 B.n939 10.6151
R2204 B.n939 B.n938 10.6151
R2205 B.n938 B.n935 10.6151
R2206 B.n935 B.n934 10.6151
R2207 B.n934 B.n931 10.6151
R2208 B.n931 B.n930 10.6151
R2209 B.n930 B.n927 10.6151
R2210 B.n927 B.n926 10.6151
R2211 B.n926 B.n923 10.6151
R2212 B.n923 B.n922 10.6151
R2213 B.n922 B.n919 10.6151
R2214 B.n919 B.n918 10.6151
R2215 B.n918 B.n915 10.6151
R2216 B.n915 B.n914 10.6151
R2217 B.n914 B.n911 10.6151
R2218 B.n911 B.n910 10.6151
R2219 B.n910 B.n907 10.6151
R2220 B.n907 B.n906 10.6151
R2221 B.n906 B.n903 10.6151
R2222 B.n903 B.n902 10.6151
R2223 B.n902 B.n899 10.6151
R2224 B.n899 B.n898 10.6151
R2225 B.n898 B.n895 10.6151
R2226 B.n895 B.n894 10.6151
R2227 B.n894 B.n891 10.6151
R2228 B.n891 B.n890 10.6151
R2229 B.n890 B.n887 10.6151
R2230 B.n887 B.n886 10.6151
R2231 B.n886 B.n883 10.6151
R2232 B.n883 B.n882 10.6151
R2233 B.n882 B.n879 10.6151
R2234 B.n879 B.n878 10.6151
R2235 B.n878 B.n875 10.6151
R2236 B.n875 B.n874 10.6151
R2237 B.n874 B.n871 10.6151
R2238 B.n871 B.n870 10.6151
R2239 B.n870 B.n867 10.6151
R2240 B.n867 B.n866 10.6151
R2241 B.n866 B.n863 10.6151
R2242 B.n863 B.n862 10.6151
R2243 B.n862 B.n859 10.6151
R2244 B.n859 B.n858 10.6151
R2245 B.n858 B.n855 10.6151
R2246 B.n855 B.n854 10.6151
R2247 B.n854 B.n851 10.6151
R2248 B.n851 B.n850 10.6151
R2249 B.n850 B.n847 10.6151
R2250 B.n847 B.n846 10.6151
R2251 B.n843 B.n842 10.6151
R2252 B.n842 B.n839 10.6151
R2253 B.n839 B.n838 10.6151
R2254 B.n838 B.n835 10.6151
R2255 B.n835 B.n834 10.6151
R2256 B.n834 B.n831 10.6151
R2257 B.n831 B.n830 10.6151
R2258 B.n830 B.n827 10.6151
R2259 B.n827 B.n826 10.6151
R2260 B.n823 B.n822 10.6151
R2261 B.n822 B.n819 10.6151
R2262 B.n819 B.n818 10.6151
R2263 B.n818 B.n815 10.6151
R2264 B.n815 B.n814 10.6151
R2265 B.n814 B.n811 10.6151
R2266 B.n811 B.n810 10.6151
R2267 B.n810 B.n807 10.6151
R2268 B.n807 B.n806 10.6151
R2269 B.n806 B.n803 10.6151
R2270 B.n803 B.n802 10.6151
R2271 B.n802 B.n799 10.6151
R2272 B.n799 B.n798 10.6151
R2273 B.n798 B.n795 10.6151
R2274 B.n795 B.n794 10.6151
R2275 B.n794 B.n791 10.6151
R2276 B.n791 B.n790 10.6151
R2277 B.n790 B.n787 10.6151
R2278 B.n787 B.n786 10.6151
R2279 B.n786 B.n783 10.6151
R2280 B.n783 B.n782 10.6151
R2281 B.n782 B.n779 10.6151
R2282 B.n779 B.n778 10.6151
R2283 B.n778 B.n775 10.6151
R2284 B.n775 B.n774 10.6151
R2285 B.n774 B.n771 10.6151
R2286 B.n771 B.n770 10.6151
R2287 B.n770 B.n767 10.6151
R2288 B.n767 B.n766 10.6151
R2289 B.n766 B.n763 10.6151
R2290 B.n763 B.n762 10.6151
R2291 B.n762 B.n759 10.6151
R2292 B.n759 B.n758 10.6151
R2293 B.n758 B.n755 10.6151
R2294 B.n755 B.n754 10.6151
R2295 B.n754 B.n751 10.6151
R2296 B.n751 B.n750 10.6151
R2297 B.n750 B.n747 10.6151
R2298 B.n747 B.n746 10.6151
R2299 B.n746 B.n743 10.6151
R2300 B.n743 B.n742 10.6151
R2301 B.n742 B.n739 10.6151
R2302 B.n739 B.n738 10.6151
R2303 B.n738 B.n735 10.6151
R2304 B.n735 B.n734 10.6151
R2305 B.n734 B.n731 10.6151
R2306 B.n731 B.n730 10.6151
R2307 B.n730 B.n727 10.6151
R2308 B.n727 B.n726 10.6151
R2309 B.n726 B.n723 10.6151
R2310 B.n723 B.n722 10.6151
R2311 B.n722 B.n719 10.6151
R2312 B.n719 B.n718 10.6151
R2313 B.n718 B.n715 10.6151
R2314 B.n715 B.n714 10.6151
R2315 B.n714 B.n711 10.6151
R2316 B.n711 B.n710 10.6151
R2317 B.n710 B.n707 10.6151
R2318 B.n707 B.n706 10.6151
R2319 B.n706 B.n703 10.6151
R2320 B.n703 B.n702 10.6151
R2321 B.n702 B.n699 10.6151
R2322 B.n699 B.n698 10.6151
R2323 B.n698 B.n696 10.6151
R2324 B.n979 B.n614 10.6151
R2325 B.n980 B.n979 10.6151
R2326 B.n981 B.n980 10.6151
R2327 B.n981 B.n606 10.6151
R2328 B.n991 B.n606 10.6151
R2329 B.n992 B.n991 10.6151
R2330 B.n993 B.n992 10.6151
R2331 B.n993 B.n599 10.6151
R2332 B.n1004 B.n599 10.6151
R2333 B.n1005 B.n1004 10.6151
R2334 B.n1006 B.n1005 10.6151
R2335 B.n1006 B.n591 10.6151
R2336 B.n1016 B.n591 10.6151
R2337 B.n1017 B.n1016 10.6151
R2338 B.n1018 B.n1017 10.6151
R2339 B.n1018 B.n583 10.6151
R2340 B.n1028 B.n583 10.6151
R2341 B.n1029 B.n1028 10.6151
R2342 B.n1030 B.n1029 10.6151
R2343 B.n1030 B.n574 10.6151
R2344 B.n1040 B.n574 10.6151
R2345 B.n1041 B.n1040 10.6151
R2346 B.n1042 B.n1041 10.6151
R2347 B.n1042 B.n567 10.6151
R2348 B.n1052 B.n567 10.6151
R2349 B.n1053 B.n1052 10.6151
R2350 B.n1054 B.n1053 10.6151
R2351 B.n1054 B.n559 10.6151
R2352 B.n1064 B.n559 10.6151
R2353 B.n1065 B.n1064 10.6151
R2354 B.n1066 B.n1065 10.6151
R2355 B.n1066 B.n552 10.6151
R2356 B.n1077 B.n552 10.6151
R2357 B.n1078 B.n1077 10.6151
R2358 B.n1079 B.n1078 10.6151
R2359 B.n1079 B.n544 10.6151
R2360 B.n1089 B.n544 10.6151
R2361 B.n1090 B.n1089 10.6151
R2362 B.n1091 B.n1090 10.6151
R2363 B.n1091 B.n536 10.6151
R2364 B.n1101 B.n536 10.6151
R2365 B.n1102 B.n1101 10.6151
R2366 B.n1103 B.n1102 10.6151
R2367 B.n1103 B.n528 10.6151
R2368 B.n1113 B.n528 10.6151
R2369 B.n1114 B.n1113 10.6151
R2370 B.n1115 B.n1114 10.6151
R2371 B.n1115 B.n520 10.6151
R2372 B.n1125 B.n520 10.6151
R2373 B.n1126 B.n1125 10.6151
R2374 B.n1127 B.n1126 10.6151
R2375 B.n1127 B.n511 10.6151
R2376 B.n1137 B.n511 10.6151
R2377 B.n1138 B.n1137 10.6151
R2378 B.n1139 B.n1138 10.6151
R2379 B.n1139 B.n504 10.6151
R2380 B.n1149 B.n504 10.6151
R2381 B.n1150 B.n1149 10.6151
R2382 B.n1151 B.n1150 10.6151
R2383 B.n1151 B.n496 10.6151
R2384 B.n1161 B.n496 10.6151
R2385 B.n1162 B.n1161 10.6151
R2386 B.n1163 B.n1162 10.6151
R2387 B.n1163 B.n489 10.6151
R2388 B.n1174 B.n489 10.6151
R2389 B.n1175 B.n1174 10.6151
R2390 B.n1177 B.n1175 10.6151
R2391 B.n1177 B.n1176 10.6151
R2392 B.n1176 B.n481 10.6151
R2393 B.n1188 B.n481 10.6151
R2394 B.n1189 B.n1188 10.6151
R2395 B.n1190 B.n1189 10.6151
R2396 B.n1191 B.n1190 10.6151
R2397 B.n1192 B.n1191 10.6151
R2398 B.n1195 B.n1192 10.6151
R2399 B.n1196 B.n1195 10.6151
R2400 B.n1197 B.n1196 10.6151
R2401 B.n1198 B.n1197 10.6151
R2402 B.n1200 B.n1198 10.6151
R2403 B.n1201 B.n1200 10.6151
R2404 B.n1202 B.n1201 10.6151
R2405 B.n1203 B.n1202 10.6151
R2406 B.n1205 B.n1203 10.6151
R2407 B.n1206 B.n1205 10.6151
R2408 B.n1207 B.n1206 10.6151
R2409 B.n1208 B.n1207 10.6151
R2410 B.n1210 B.n1208 10.6151
R2411 B.n1211 B.n1210 10.6151
R2412 B.n1212 B.n1211 10.6151
R2413 B.n1213 B.n1212 10.6151
R2414 B.n1215 B.n1213 10.6151
R2415 B.n1216 B.n1215 10.6151
R2416 B.n1217 B.n1216 10.6151
R2417 B.n1218 B.n1217 10.6151
R2418 B.n1220 B.n1218 10.6151
R2419 B.n1221 B.n1220 10.6151
R2420 B.n1222 B.n1221 10.6151
R2421 B.n1223 B.n1222 10.6151
R2422 B.n1225 B.n1223 10.6151
R2423 B.n1226 B.n1225 10.6151
R2424 B.n1227 B.n1226 10.6151
R2425 B.n1228 B.n1227 10.6151
R2426 B.n1230 B.n1228 10.6151
R2427 B.n1231 B.n1230 10.6151
R2428 B.n1232 B.n1231 10.6151
R2429 B.n1233 B.n1232 10.6151
R2430 B.n1235 B.n1233 10.6151
R2431 B.n1236 B.n1235 10.6151
R2432 B.n1237 B.n1236 10.6151
R2433 B.n1238 B.n1237 10.6151
R2434 B.n1240 B.n1238 10.6151
R2435 B.n1241 B.n1240 10.6151
R2436 B.n1242 B.n1241 10.6151
R2437 B.n1243 B.n1242 10.6151
R2438 B.n1245 B.n1243 10.6151
R2439 B.n1246 B.n1245 10.6151
R2440 B.n1247 B.n1246 10.6151
R2441 B.n1248 B.n1247 10.6151
R2442 B.n1250 B.n1248 10.6151
R2443 B.n1251 B.n1250 10.6151
R2444 B.n1252 B.n1251 10.6151
R2445 B.n1253 B.n1252 10.6151
R2446 B.n1255 B.n1253 10.6151
R2447 B.n1256 B.n1255 10.6151
R2448 B.n1257 B.n1256 10.6151
R2449 B.n1258 B.n1257 10.6151
R2450 B.n1260 B.n1258 10.6151
R2451 B.n1261 B.n1260 10.6151
R2452 B.n1262 B.n1261 10.6151
R2453 B.n1263 B.n1262 10.6151
R2454 B.n1265 B.n1263 10.6151
R2455 B.n1266 B.n1265 10.6151
R2456 B.n1267 B.n1266 10.6151
R2457 B.n1268 B.n1267 10.6151
R2458 B.n1270 B.n1268 10.6151
R2459 B.n1271 B.n1270 10.6151
R2460 B.n1272 B.n1271 10.6151
R2461 B.n1273 B.n1272 10.6151
R2462 B.n1275 B.n1273 10.6151
R2463 B.n1276 B.n1275 10.6151
R2464 B.n1277 B.n1276 10.6151
R2465 B.n1278 B.n1277 10.6151
R2466 B.n1279 B.n1278 10.6151
R2467 B.n1424 B.n1 10.6151
R2468 B.n1424 B.n1423 10.6151
R2469 B.n1423 B.n1422 10.6151
R2470 B.n1422 B.n10 10.6151
R2471 B.n1416 B.n10 10.6151
R2472 B.n1416 B.n1415 10.6151
R2473 B.n1415 B.n1414 10.6151
R2474 B.n1414 B.n17 10.6151
R2475 B.n1408 B.n17 10.6151
R2476 B.n1408 B.n1407 10.6151
R2477 B.n1407 B.n1406 10.6151
R2478 B.n1406 B.n25 10.6151
R2479 B.n1400 B.n25 10.6151
R2480 B.n1400 B.n1399 10.6151
R2481 B.n1399 B.n1398 10.6151
R2482 B.n1398 B.n32 10.6151
R2483 B.n1392 B.n32 10.6151
R2484 B.n1392 B.n1391 10.6151
R2485 B.n1391 B.n1390 10.6151
R2486 B.n1390 B.n39 10.6151
R2487 B.n1384 B.n39 10.6151
R2488 B.n1384 B.n1383 10.6151
R2489 B.n1383 B.n1382 10.6151
R2490 B.n1382 B.n46 10.6151
R2491 B.n1376 B.n46 10.6151
R2492 B.n1376 B.n1375 10.6151
R2493 B.n1375 B.n1374 10.6151
R2494 B.n1374 B.n53 10.6151
R2495 B.n1368 B.n53 10.6151
R2496 B.n1368 B.n1367 10.6151
R2497 B.n1367 B.n1366 10.6151
R2498 B.n1366 B.n60 10.6151
R2499 B.n1360 B.n60 10.6151
R2500 B.n1360 B.n1359 10.6151
R2501 B.n1359 B.n1358 10.6151
R2502 B.n1358 B.n67 10.6151
R2503 B.n1352 B.n67 10.6151
R2504 B.n1352 B.n1351 10.6151
R2505 B.n1351 B.n1350 10.6151
R2506 B.n1350 B.n73 10.6151
R2507 B.n1344 B.n73 10.6151
R2508 B.n1344 B.n1343 10.6151
R2509 B.n1343 B.n1342 10.6151
R2510 B.n1342 B.n81 10.6151
R2511 B.n1336 B.n81 10.6151
R2512 B.n1336 B.n1335 10.6151
R2513 B.n1335 B.n1334 10.6151
R2514 B.n1334 B.n88 10.6151
R2515 B.n1328 B.n88 10.6151
R2516 B.n1328 B.n1327 10.6151
R2517 B.n1327 B.n1326 10.6151
R2518 B.n1326 B.n95 10.6151
R2519 B.n1320 B.n95 10.6151
R2520 B.n1320 B.n1319 10.6151
R2521 B.n1319 B.n1318 10.6151
R2522 B.n1318 B.n102 10.6151
R2523 B.n1312 B.n102 10.6151
R2524 B.n1312 B.n1311 10.6151
R2525 B.n1311 B.n1310 10.6151
R2526 B.n1310 B.n109 10.6151
R2527 B.n1304 B.n109 10.6151
R2528 B.n1304 B.n1303 10.6151
R2529 B.n1303 B.n1302 10.6151
R2530 B.n1302 B.n115 10.6151
R2531 B.n1296 B.n115 10.6151
R2532 B.n1296 B.n1295 10.6151
R2533 B.n1295 B.n1294 10.6151
R2534 B.n1294 B.n123 10.6151
R2535 B.n1288 B.n123 10.6151
R2536 B.n1288 B.n1287 10.6151
R2537 B.n1286 B.n130 10.6151
R2538 B.n207 B.n130 10.6151
R2539 B.n208 B.n207 10.6151
R2540 B.n211 B.n208 10.6151
R2541 B.n212 B.n211 10.6151
R2542 B.n215 B.n212 10.6151
R2543 B.n216 B.n215 10.6151
R2544 B.n219 B.n216 10.6151
R2545 B.n220 B.n219 10.6151
R2546 B.n223 B.n220 10.6151
R2547 B.n224 B.n223 10.6151
R2548 B.n227 B.n224 10.6151
R2549 B.n228 B.n227 10.6151
R2550 B.n231 B.n228 10.6151
R2551 B.n232 B.n231 10.6151
R2552 B.n235 B.n232 10.6151
R2553 B.n236 B.n235 10.6151
R2554 B.n239 B.n236 10.6151
R2555 B.n240 B.n239 10.6151
R2556 B.n243 B.n240 10.6151
R2557 B.n244 B.n243 10.6151
R2558 B.n247 B.n244 10.6151
R2559 B.n248 B.n247 10.6151
R2560 B.n251 B.n248 10.6151
R2561 B.n252 B.n251 10.6151
R2562 B.n255 B.n252 10.6151
R2563 B.n256 B.n255 10.6151
R2564 B.n259 B.n256 10.6151
R2565 B.n260 B.n259 10.6151
R2566 B.n263 B.n260 10.6151
R2567 B.n264 B.n263 10.6151
R2568 B.n267 B.n264 10.6151
R2569 B.n268 B.n267 10.6151
R2570 B.n271 B.n268 10.6151
R2571 B.n272 B.n271 10.6151
R2572 B.n275 B.n272 10.6151
R2573 B.n276 B.n275 10.6151
R2574 B.n279 B.n276 10.6151
R2575 B.n280 B.n279 10.6151
R2576 B.n283 B.n280 10.6151
R2577 B.n284 B.n283 10.6151
R2578 B.n287 B.n284 10.6151
R2579 B.n288 B.n287 10.6151
R2580 B.n291 B.n288 10.6151
R2581 B.n292 B.n291 10.6151
R2582 B.n295 B.n292 10.6151
R2583 B.n296 B.n295 10.6151
R2584 B.n299 B.n296 10.6151
R2585 B.n300 B.n299 10.6151
R2586 B.n303 B.n300 10.6151
R2587 B.n304 B.n303 10.6151
R2588 B.n307 B.n304 10.6151
R2589 B.n308 B.n307 10.6151
R2590 B.n311 B.n308 10.6151
R2591 B.n312 B.n311 10.6151
R2592 B.n315 B.n312 10.6151
R2593 B.n316 B.n315 10.6151
R2594 B.n319 B.n316 10.6151
R2595 B.n320 B.n319 10.6151
R2596 B.n323 B.n320 10.6151
R2597 B.n324 B.n323 10.6151
R2598 B.n327 B.n324 10.6151
R2599 B.n328 B.n327 10.6151
R2600 B.n331 B.n328 10.6151
R2601 B.n336 B.n333 10.6151
R2602 B.n337 B.n336 10.6151
R2603 B.n340 B.n337 10.6151
R2604 B.n341 B.n340 10.6151
R2605 B.n344 B.n341 10.6151
R2606 B.n345 B.n344 10.6151
R2607 B.n348 B.n345 10.6151
R2608 B.n349 B.n348 10.6151
R2609 B.n352 B.n349 10.6151
R2610 B.n357 B.n354 10.6151
R2611 B.n358 B.n357 10.6151
R2612 B.n361 B.n358 10.6151
R2613 B.n362 B.n361 10.6151
R2614 B.n365 B.n362 10.6151
R2615 B.n366 B.n365 10.6151
R2616 B.n369 B.n366 10.6151
R2617 B.n370 B.n369 10.6151
R2618 B.n373 B.n370 10.6151
R2619 B.n374 B.n373 10.6151
R2620 B.n377 B.n374 10.6151
R2621 B.n378 B.n377 10.6151
R2622 B.n381 B.n378 10.6151
R2623 B.n382 B.n381 10.6151
R2624 B.n385 B.n382 10.6151
R2625 B.n386 B.n385 10.6151
R2626 B.n389 B.n386 10.6151
R2627 B.n390 B.n389 10.6151
R2628 B.n393 B.n390 10.6151
R2629 B.n394 B.n393 10.6151
R2630 B.n397 B.n394 10.6151
R2631 B.n398 B.n397 10.6151
R2632 B.n401 B.n398 10.6151
R2633 B.n402 B.n401 10.6151
R2634 B.n405 B.n402 10.6151
R2635 B.n406 B.n405 10.6151
R2636 B.n409 B.n406 10.6151
R2637 B.n410 B.n409 10.6151
R2638 B.n413 B.n410 10.6151
R2639 B.n414 B.n413 10.6151
R2640 B.n417 B.n414 10.6151
R2641 B.n418 B.n417 10.6151
R2642 B.n421 B.n418 10.6151
R2643 B.n422 B.n421 10.6151
R2644 B.n425 B.n422 10.6151
R2645 B.n426 B.n425 10.6151
R2646 B.n429 B.n426 10.6151
R2647 B.n430 B.n429 10.6151
R2648 B.n433 B.n430 10.6151
R2649 B.n434 B.n433 10.6151
R2650 B.n437 B.n434 10.6151
R2651 B.n438 B.n437 10.6151
R2652 B.n441 B.n438 10.6151
R2653 B.n442 B.n441 10.6151
R2654 B.n445 B.n442 10.6151
R2655 B.n446 B.n445 10.6151
R2656 B.n449 B.n446 10.6151
R2657 B.n450 B.n449 10.6151
R2658 B.n453 B.n450 10.6151
R2659 B.n454 B.n453 10.6151
R2660 B.n457 B.n454 10.6151
R2661 B.n458 B.n457 10.6151
R2662 B.n461 B.n458 10.6151
R2663 B.n462 B.n461 10.6151
R2664 B.n465 B.n462 10.6151
R2665 B.n466 B.n465 10.6151
R2666 B.n469 B.n466 10.6151
R2667 B.n470 B.n469 10.6151
R2668 B.n473 B.n470 10.6151
R2669 B.n474 B.n473 10.6151
R2670 B.n477 B.n474 10.6151
R2671 B.n479 B.n477 10.6151
R2672 B.n480 B.n479 10.6151
R2673 B.n1280 B.n480 10.6151
R2674 B.n846 B.n692 9.36635
R2675 B.n823 B.n695 9.36635
R2676 B.n332 B.n331 9.36635
R2677 B.n354 B.n353 9.36635
R2678 B.n1432 B.n0 8.11757
R2679 B.n1432 B.n1 8.11757
R2680 B.n1075 B.t21 1.7448
R2681 B.n514 B.t5 1.7448
R2682 B.t23 B.n1395 1.7448
R2683 B.n1354 B.t20 1.7448
R2684 B.n843 B.n692 1.24928
R2685 B.n826 B.n695 1.24928
R2686 B.n333 B.n332 1.24928
R2687 B.n353 B.n352 1.24928
R2688 VN.n62 VN.t5 179.389
R2689 VN.n13 VN.t2 179.389
R2690 VN.n96 VN.n95 161.3
R2691 VN.n94 VN.n50 161.3
R2692 VN.n93 VN.n92 161.3
R2693 VN.n91 VN.n51 161.3
R2694 VN.n90 VN.n89 161.3
R2695 VN.n88 VN.n52 161.3
R2696 VN.n87 VN.n86 161.3
R2697 VN.n85 VN.n84 161.3
R2698 VN.n83 VN.n54 161.3
R2699 VN.n82 VN.n81 161.3
R2700 VN.n80 VN.n55 161.3
R2701 VN.n79 VN.n78 161.3
R2702 VN.n77 VN.n56 161.3
R2703 VN.n76 VN.n75 161.3
R2704 VN.n74 VN.n57 161.3
R2705 VN.n73 VN.n72 161.3
R2706 VN.n71 VN.n58 161.3
R2707 VN.n70 VN.n69 161.3
R2708 VN.n68 VN.n59 161.3
R2709 VN.n67 VN.n66 161.3
R2710 VN.n65 VN.n60 161.3
R2711 VN.n64 VN.n63 161.3
R2712 VN.n47 VN.n46 161.3
R2713 VN.n45 VN.n1 161.3
R2714 VN.n44 VN.n43 161.3
R2715 VN.n42 VN.n2 161.3
R2716 VN.n41 VN.n40 161.3
R2717 VN.n39 VN.n3 161.3
R2718 VN.n38 VN.n37 161.3
R2719 VN.n36 VN.n35 161.3
R2720 VN.n34 VN.n5 161.3
R2721 VN.n33 VN.n32 161.3
R2722 VN.n31 VN.n6 161.3
R2723 VN.n30 VN.n29 161.3
R2724 VN.n28 VN.n7 161.3
R2725 VN.n27 VN.n26 161.3
R2726 VN.n25 VN.n8 161.3
R2727 VN.n24 VN.n23 161.3
R2728 VN.n22 VN.n9 161.3
R2729 VN.n21 VN.n20 161.3
R2730 VN.n19 VN.n10 161.3
R2731 VN.n18 VN.n17 161.3
R2732 VN.n16 VN.n11 161.3
R2733 VN.n15 VN.n14 161.3
R2734 VN.n8 VN.t8 147.483
R2735 VN.n12 VN.t0 147.483
R2736 VN.n4 VN.t1 147.483
R2737 VN.n0 VN.t3 147.483
R2738 VN.n57 VN.t9 147.483
R2739 VN.n61 VN.t6 147.483
R2740 VN.n53 VN.t4 147.483
R2741 VN.n49 VN.t7 147.483
R2742 VN.n48 VN.n0 81.2593
R2743 VN.n97 VN.n49 81.2593
R2744 VN.n13 VN.n12 70.1236
R2745 VN.n62 VN.n61 70.1236
R2746 VN VN.n97 62.9033
R2747 VN.n21 VN.n10 56.5193
R2748 VN.n29 VN.n6 56.5193
R2749 VN.n70 VN.n59 56.5193
R2750 VN.n78 VN.n55 56.5193
R2751 VN.n40 VN.n2 51.663
R2752 VN.n89 VN.n51 51.663
R2753 VN.n44 VN.n2 29.3238
R2754 VN.n93 VN.n51 29.3238
R2755 VN.n16 VN.n15 24.4675
R2756 VN.n17 VN.n16 24.4675
R2757 VN.n17 VN.n10 24.4675
R2758 VN.n22 VN.n21 24.4675
R2759 VN.n23 VN.n22 24.4675
R2760 VN.n23 VN.n8 24.4675
R2761 VN.n27 VN.n8 24.4675
R2762 VN.n28 VN.n27 24.4675
R2763 VN.n29 VN.n28 24.4675
R2764 VN.n33 VN.n6 24.4675
R2765 VN.n34 VN.n33 24.4675
R2766 VN.n35 VN.n34 24.4675
R2767 VN.n39 VN.n38 24.4675
R2768 VN.n40 VN.n39 24.4675
R2769 VN.n45 VN.n44 24.4675
R2770 VN.n46 VN.n45 24.4675
R2771 VN.n66 VN.n59 24.4675
R2772 VN.n66 VN.n65 24.4675
R2773 VN.n65 VN.n64 24.4675
R2774 VN.n78 VN.n77 24.4675
R2775 VN.n77 VN.n76 24.4675
R2776 VN.n76 VN.n57 24.4675
R2777 VN.n72 VN.n57 24.4675
R2778 VN.n72 VN.n71 24.4675
R2779 VN.n71 VN.n70 24.4675
R2780 VN.n89 VN.n88 24.4675
R2781 VN.n88 VN.n87 24.4675
R2782 VN.n84 VN.n83 24.4675
R2783 VN.n83 VN.n82 24.4675
R2784 VN.n82 VN.n55 24.4675
R2785 VN.n95 VN.n94 24.4675
R2786 VN.n94 VN.n93 24.4675
R2787 VN.n38 VN.n4 20.0634
R2788 VN.n87 VN.n53 20.0634
R2789 VN.n46 VN.n0 8.80862
R2790 VN.n95 VN.n49 8.80862
R2791 VN.n63 VN.n62 4.46393
R2792 VN.n14 VN.n13 4.46393
R2793 VN.n15 VN.n12 4.40456
R2794 VN.n35 VN.n4 4.40456
R2795 VN.n64 VN.n61 4.40456
R2796 VN.n84 VN.n53 4.40456
R2797 VN.n97 VN.n96 0.354971
R2798 VN.n48 VN.n47 0.354971
R2799 VN VN.n48 0.26696
R2800 VN.n96 VN.n50 0.189894
R2801 VN.n92 VN.n50 0.189894
R2802 VN.n92 VN.n91 0.189894
R2803 VN.n91 VN.n90 0.189894
R2804 VN.n90 VN.n52 0.189894
R2805 VN.n86 VN.n52 0.189894
R2806 VN.n86 VN.n85 0.189894
R2807 VN.n85 VN.n54 0.189894
R2808 VN.n81 VN.n54 0.189894
R2809 VN.n81 VN.n80 0.189894
R2810 VN.n80 VN.n79 0.189894
R2811 VN.n79 VN.n56 0.189894
R2812 VN.n75 VN.n56 0.189894
R2813 VN.n75 VN.n74 0.189894
R2814 VN.n74 VN.n73 0.189894
R2815 VN.n73 VN.n58 0.189894
R2816 VN.n69 VN.n58 0.189894
R2817 VN.n69 VN.n68 0.189894
R2818 VN.n68 VN.n67 0.189894
R2819 VN.n67 VN.n60 0.189894
R2820 VN.n63 VN.n60 0.189894
R2821 VN.n14 VN.n11 0.189894
R2822 VN.n18 VN.n11 0.189894
R2823 VN.n19 VN.n18 0.189894
R2824 VN.n20 VN.n19 0.189894
R2825 VN.n20 VN.n9 0.189894
R2826 VN.n24 VN.n9 0.189894
R2827 VN.n25 VN.n24 0.189894
R2828 VN.n26 VN.n25 0.189894
R2829 VN.n26 VN.n7 0.189894
R2830 VN.n30 VN.n7 0.189894
R2831 VN.n31 VN.n30 0.189894
R2832 VN.n32 VN.n31 0.189894
R2833 VN.n32 VN.n5 0.189894
R2834 VN.n36 VN.n5 0.189894
R2835 VN.n37 VN.n36 0.189894
R2836 VN.n37 VN.n3 0.189894
R2837 VN.n41 VN.n3 0.189894
R2838 VN.n42 VN.n41 0.189894
R2839 VN.n43 VN.n42 0.189894
R2840 VN.n43 VN.n1 0.189894
R2841 VN.n47 VN.n1 0.189894
R2842 VDD2.n1 VDD2.t7 62.9359
R2843 VDD2.n3 VDD2.n2 61.1145
R2844 VDD2 VDD2.n7 61.1117
R2845 VDD2.n4 VDD2.t2 59.8412
R2846 VDD2.n6 VDD2.n5 58.8488
R2847 VDD2.n1 VDD2.n0 58.8487
R2848 VDD2.n4 VDD2.n3 55.614
R2849 VDD2.n6 VDD2.n4 3.09533
R2850 VDD2.n7 VDD2.t3 0.992981
R2851 VDD2.n7 VDD2.t4 0.992981
R2852 VDD2.n5 VDD2.t5 0.992981
R2853 VDD2.n5 VDD2.t0 0.992981
R2854 VDD2.n2 VDD2.t8 0.992981
R2855 VDD2.n2 VDD2.t6 0.992981
R2856 VDD2.n0 VDD2.t9 0.992981
R2857 VDD2.n0 VDD2.t1 0.992981
R2858 VDD2 VDD2.n6 0.832397
R2859 VDD2.n3 VDD2.n1 0.718861
C0 VTAIL VDD1 13.9488f
C1 VN VTAIL 18.675901f
C2 VTAIL VDD2 14.0033f
C3 VTAIL VP 18.6903f
C4 VN VDD1 0.154942f
C5 VDD1 VDD2 2.60553f
C6 VN VDD2 18.1191f
C7 VP VDD1 18.6275f
C8 VN VP 10.849299f
C9 VP VDD2 0.668387f
C10 VDD2 B 9.360055f
C11 VDD1 B 9.350011f
C12 VTAIL B 11.932043f
C13 VN B 21.927628f
C14 VP B 20.405878f
C15 VDD2.t7 B 4.33939f
C16 VDD2.t9 B 0.36923f
C17 VDD2.t1 B 0.36923f
C18 VDD2.n0 B 3.37395f
C19 VDD2.n1 B 0.970912f
C20 VDD2.t8 B 0.36923f
C21 VDD2.t6 B 0.36923f
C22 VDD2.n2 B 3.39668f
C23 VDD2.n3 B 3.51829f
C24 VDD2.t2 B 4.3144f
C25 VDD2.n4 B 3.74313f
C26 VDD2.t5 B 0.36923f
C27 VDD2.t0 B 0.36923f
C28 VDD2.n5 B 3.37394f
C29 VDD2.n6 B 0.495267f
C30 VDD2.t3 B 0.36923f
C31 VDD2.t4 B 0.36923f
C32 VDD2.n7 B 3.39663f
C33 VN.t3 B 3.10925f
C34 VN.n0 B 1.13154f
C35 VN.n1 B 0.017349f
C36 VN.n2 B 0.017215f
C37 VN.n3 B 0.017349f
C38 VN.t1 B 3.10925f
C39 VN.n4 B 1.06999f
C40 VN.n5 B 0.017349f
C41 VN.n6 B 0.023152f
C42 VN.n7 B 0.017349f
C43 VN.t8 B 3.10925f
C44 VN.n8 B 1.08636f
C45 VN.n9 B 0.017349f
C46 VN.n10 B 0.023152f
C47 VN.n11 B 0.017349f
C48 VN.t0 B 3.10925f
C49 VN.n12 B 1.12321f
C50 VN.t2 B 3.32086f
C51 VN.n13 B 1.08724f
C52 VN.n14 B 0.204364f
C53 VN.n15 B 0.019244f
C54 VN.n16 B 0.032334f
C55 VN.n17 B 0.032334f
C56 VN.n18 B 0.017349f
C57 VN.n19 B 0.017349f
C58 VN.n20 B 0.017349f
C59 VN.n21 B 0.027503f
C60 VN.n22 B 0.032334f
C61 VN.n23 B 0.032334f
C62 VN.n24 B 0.017349f
C63 VN.n25 B 0.017349f
C64 VN.n26 B 0.017349f
C65 VN.n27 B 0.032334f
C66 VN.n28 B 0.032334f
C67 VN.n29 B 0.027503f
C68 VN.n30 B 0.017349f
C69 VN.n31 B 0.017349f
C70 VN.n32 B 0.017349f
C71 VN.n33 B 0.032334f
C72 VN.n34 B 0.032334f
C73 VN.n35 B 0.019244f
C74 VN.n36 B 0.017349f
C75 VN.n37 B 0.017349f
C76 VN.n38 B 0.029461f
C77 VN.n39 B 0.032334f
C78 VN.n40 B 0.031326f
C79 VN.n41 B 0.017349f
C80 VN.n42 B 0.017349f
C81 VN.n43 B 0.017349f
C82 VN.n44 B 0.034449f
C83 VN.n45 B 0.032334f
C84 VN.n46 B 0.022117f
C85 VN.n47 B 0.028001f
C86 VN.n48 B 0.045278f
C87 VN.t7 B 3.10925f
C88 VN.n49 B 1.13154f
C89 VN.n50 B 0.017349f
C90 VN.n51 B 0.017215f
C91 VN.n52 B 0.017349f
C92 VN.t4 B 3.10925f
C93 VN.n53 B 1.06999f
C94 VN.n54 B 0.017349f
C95 VN.n55 B 0.023152f
C96 VN.n56 B 0.017349f
C97 VN.t9 B 3.10925f
C98 VN.n57 B 1.08636f
C99 VN.n58 B 0.017349f
C100 VN.n59 B 0.023152f
C101 VN.n60 B 0.017349f
C102 VN.t6 B 3.10925f
C103 VN.n61 B 1.12321f
C104 VN.t5 B 3.32086f
C105 VN.n62 B 1.08724f
C106 VN.n63 B 0.204364f
C107 VN.n64 B 0.019244f
C108 VN.n65 B 0.032334f
C109 VN.n66 B 0.032334f
C110 VN.n67 B 0.017349f
C111 VN.n68 B 0.017349f
C112 VN.n69 B 0.017349f
C113 VN.n70 B 0.027503f
C114 VN.n71 B 0.032334f
C115 VN.n72 B 0.032334f
C116 VN.n73 B 0.017349f
C117 VN.n74 B 0.017349f
C118 VN.n75 B 0.017349f
C119 VN.n76 B 0.032334f
C120 VN.n77 B 0.032334f
C121 VN.n78 B 0.027503f
C122 VN.n79 B 0.017349f
C123 VN.n80 B 0.017349f
C124 VN.n81 B 0.017349f
C125 VN.n82 B 0.032334f
C126 VN.n83 B 0.032334f
C127 VN.n84 B 0.019244f
C128 VN.n85 B 0.017349f
C129 VN.n86 B 0.017349f
C130 VN.n87 B 0.029461f
C131 VN.n88 B 0.032334f
C132 VN.n89 B 0.031326f
C133 VN.n90 B 0.017349f
C134 VN.n91 B 0.017349f
C135 VN.n92 B 0.017349f
C136 VN.n93 B 0.034449f
C137 VN.n94 B 0.032334f
C138 VN.n95 B 0.022117f
C139 VN.n96 B 0.028001f
C140 VN.n97 B 1.3562f
C141 VTAIL.t1 B 0.373003f
C142 VTAIL.t17 B 0.373003f
C143 VTAIL.n0 B 3.33073f
C144 VTAIL.n1 B 0.581684f
C145 VTAIL.t14 B 4.25658f
C146 VTAIL.n2 B 0.727658f
C147 VTAIL.t13 B 0.373003f
C148 VTAIL.t8 B 0.373003f
C149 VTAIL.n3 B 3.33073f
C150 VTAIL.n4 B 0.718387f
C151 VTAIL.t12 B 0.373003f
C152 VTAIL.t10 B 0.373003f
C153 VTAIL.n5 B 3.33073f
C154 VTAIL.n6 B 2.58689f
C155 VTAIL.t2 B 0.373003f
C156 VTAIL.t18 B 0.373003f
C157 VTAIL.n7 B 3.33072f
C158 VTAIL.n8 B 2.58689f
C159 VTAIL.t4 B 0.373003f
C160 VTAIL.t5 B 0.373003f
C161 VTAIL.n9 B 3.33072f
C162 VTAIL.n10 B 0.718394f
C163 VTAIL.t0 B 4.25661f
C164 VTAIL.n11 B 0.727634f
C165 VTAIL.t9 B 0.373003f
C166 VTAIL.t15 B 0.373003f
C167 VTAIL.n12 B 3.33072f
C168 VTAIL.n13 B 0.636241f
C169 VTAIL.t7 B 0.373003f
C170 VTAIL.t6 B 0.373003f
C171 VTAIL.n14 B 3.33072f
C172 VTAIL.n15 B 0.718394f
C173 VTAIL.t11 B 4.2566f
C174 VTAIL.n16 B 2.44235f
C175 VTAIL.t16 B 4.25658f
C176 VTAIL.n17 B 2.44237f
C177 VTAIL.t3 B 0.373003f
C178 VTAIL.t19 B 0.373003f
C179 VTAIL.n18 B 3.33073f
C180 VTAIL.n19 B 0.536993f
C181 VDD1.t9 B 4.37851f
C182 VDD1.t7 B 0.372557f
C183 VDD1.t3 B 0.372557f
C184 VDD1.n0 B 3.40435f
C185 VDD1.n1 B 0.987534f
C186 VDD1.t4 B 4.3785f
C187 VDD1.t0 B 0.372557f
C188 VDD1.t5 B 0.372557f
C189 VDD1.n2 B 3.40435f
C190 VDD1.n3 B 0.979662f
C191 VDD1.t8 B 0.372557f
C192 VDD1.t6 B 0.372557f
C193 VDD1.n4 B 3.42729f
C194 VDD1.n5 B 3.69004f
C195 VDD1.t2 B 0.372557f
C196 VDD1.t1 B 0.372557f
C197 VDD1.n6 B 3.40435f
C198 VDD1.n7 B 3.82929f
C199 VP.t1 B 3.14352f
C200 VP.n0 B 1.14401f
C201 VP.n1 B 0.01754f
C202 VP.n2 B 0.017405f
C203 VP.n3 B 0.01754f
C204 VP.t7 B 3.14352f
C205 VP.n4 B 1.08178f
C206 VP.n5 B 0.01754f
C207 VP.n6 B 0.023408f
C208 VP.n7 B 0.01754f
C209 VP.t2 B 3.14352f
C210 VP.n8 B 1.09834f
C211 VP.n9 B 0.01754f
C212 VP.n10 B 0.023408f
C213 VP.n11 B 0.01754f
C214 VP.t5 B 3.14352f
C215 VP.n12 B 1.08178f
C216 VP.n13 B 0.01754f
C217 VP.n14 B 0.017405f
C218 VP.n15 B 0.01754f
C219 VP.t3 B 3.14352f
C220 VP.n16 B 1.14401f
C221 VP.t4 B 3.14352f
C222 VP.n17 B 1.14401f
C223 VP.n18 B 0.01754f
C224 VP.n19 B 0.017405f
C225 VP.n20 B 0.01754f
C226 VP.t9 B 3.14352f
C227 VP.n21 B 1.08178f
C228 VP.n22 B 0.01754f
C229 VP.n23 B 0.023408f
C230 VP.n24 B 0.01754f
C231 VP.t8 B 3.14352f
C232 VP.n25 B 1.09834f
C233 VP.n26 B 0.01754f
C234 VP.n27 B 0.023408f
C235 VP.n28 B 0.01754f
C236 VP.t0 B 3.14352f
C237 VP.n29 B 1.13559f
C238 VP.t6 B 3.35746f
C239 VP.n30 B 1.09923f
C240 VP.n31 B 0.206617f
C241 VP.n32 B 0.019456f
C242 VP.n33 B 0.03269f
C243 VP.n34 B 0.03269f
C244 VP.n35 B 0.01754f
C245 VP.n36 B 0.01754f
C246 VP.n37 B 0.01754f
C247 VP.n38 B 0.027806f
C248 VP.n39 B 0.03269f
C249 VP.n40 B 0.03269f
C250 VP.n41 B 0.01754f
C251 VP.n42 B 0.01754f
C252 VP.n43 B 0.01754f
C253 VP.n44 B 0.03269f
C254 VP.n45 B 0.03269f
C255 VP.n46 B 0.027806f
C256 VP.n47 B 0.01754f
C257 VP.n48 B 0.01754f
C258 VP.n49 B 0.01754f
C259 VP.n50 B 0.03269f
C260 VP.n51 B 0.03269f
C261 VP.n52 B 0.019456f
C262 VP.n53 B 0.01754f
C263 VP.n54 B 0.01754f
C264 VP.n55 B 0.029785f
C265 VP.n56 B 0.03269f
C266 VP.n57 B 0.031671f
C267 VP.n58 B 0.01754f
C268 VP.n59 B 0.01754f
C269 VP.n60 B 0.01754f
C270 VP.n61 B 0.034829f
C271 VP.n62 B 0.03269f
C272 VP.n63 B 0.022361f
C273 VP.n64 B 0.028309f
C274 VP.n65 B 1.36446f
C275 VP.n66 B 1.37451f
C276 VP.n67 B 0.028309f
C277 VP.n68 B 0.022361f
C278 VP.n69 B 0.03269f
C279 VP.n70 B 0.034829f
C280 VP.n71 B 0.01754f
C281 VP.n72 B 0.01754f
C282 VP.n73 B 0.01754f
C283 VP.n74 B 0.031671f
C284 VP.n75 B 0.03269f
C285 VP.n76 B 0.029785f
C286 VP.n77 B 0.01754f
C287 VP.n78 B 0.01754f
C288 VP.n79 B 0.019456f
C289 VP.n80 B 0.03269f
C290 VP.n81 B 0.03269f
C291 VP.n82 B 0.01754f
C292 VP.n83 B 0.01754f
C293 VP.n84 B 0.01754f
C294 VP.n85 B 0.027806f
C295 VP.n86 B 0.03269f
C296 VP.n87 B 0.03269f
C297 VP.n88 B 0.01754f
C298 VP.n89 B 0.01754f
C299 VP.n90 B 0.01754f
C300 VP.n91 B 0.03269f
C301 VP.n92 B 0.03269f
C302 VP.n93 B 0.027806f
C303 VP.n94 B 0.01754f
C304 VP.n95 B 0.01754f
C305 VP.n96 B 0.01754f
C306 VP.n97 B 0.03269f
C307 VP.n98 B 0.03269f
C308 VP.n99 B 0.019456f
C309 VP.n100 B 0.01754f
C310 VP.n101 B 0.01754f
C311 VP.n102 B 0.029785f
C312 VP.n103 B 0.03269f
C313 VP.n104 B 0.031671f
C314 VP.n105 B 0.01754f
C315 VP.n106 B 0.01754f
C316 VP.n107 B 0.01754f
C317 VP.n108 B 0.034829f
C318 VP.n109 B 0.03269f
C319 VP.n110 B 0.022361f
C320 VP.n111 B 0.028309f
C321 VP.n112 B 0.045777f
.ends

