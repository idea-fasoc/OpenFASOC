* NGSPICE file created from diff_pair_sample_1692.ext - technology: sky130A

.subckt diff_pair_sample_1692 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=0.38
X1 VTAIL.t7 VP.t0 VDD1.t0 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=0.38
X2 VDD1.t1 VP.t1 VTAIL.t6 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=0.38
X3 VDD1.t3 VP.t2 VTAIL.t5 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=0.38
X4 VTAIL.t4 VP.t3 VDD1.t2 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=0.38
X5 VTAIL.t2 VN.t0 VDD2.t3 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=0.38
X6 B.t8 B.t6 B.t7 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=0.38
X7 VDD2.t2 VN.t1 VTAIL.t3 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=0.38
X8 B.t5 B.t3 B.t4 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=0.38
X9 VDD2.t1 VN.t2 VTAIL.t0 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.24255 pd=1.8 as=0.5733 ps=3.72 w=1.47 l=0.38
X10 VTAIL.t1 VN.t3 VDD2.t0 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0.24255 ps=1.8 w=1.47 l=0.38
X11 B.t2 B.t0 B.t1 w_n1396_n1266# sky130_fd_pr__pfet_01v8 ad=0.5733 pd=3.72 as=0 ps=0 w=1.47 l=0.38
R0 B.n138 B.n137 585
R1 B.n136 B.n45 585
R2 B.n135 B.n134 585
R3 B.n133 B.n46 585
R4 B.n132 B.n131 585
R5 B.n130 B.n47 585
R6 B.n129 B.n128 585
R7 B.n127 B.n48 585
R8 B.n126 B.n125 585
R9 B.n124 B.n49 585
R10 B.n123 B.n122 585
R11 B.n120 B.n50 585
R12 B.n119 B.n118 585
R13 B.n117 B.n53 585
R14 B.n116 B.n115 585
R15 B.n114 B.n54 585
R16 B.n113 B.n112 585
R17 B.n111 B.n55 585
R18 B.n110 B.n109 585
R19 B.n108 B.n56 585
R20 B.n106 B.n105 585
R21 B.n104 B.n59 585
R22 B.n103 B.n102 585
R23 B.n101 B.n60 585
R24 B.n100 B.n99 585
R25 B.n98 B.n61 585
R26 B.n97 B.n96 585
R27 B.n95 B.n62 585
R28 B.n94 B.n93 585
R29 B.n92 B.n63 585
R30 B.n91 B.n90 585
R31 B.n139 B.n44 585
R32 B.n141 B.n140 585
R33 B.n142 B.n43 585
R34 B.n144 B.n143 585
R35 B.n145 B.n42 585
R36 B.n147 B.n146 585
R37 B.n148 B.n41 585
R38 B.n150 B.n149 585
R39 B.n151 B.n40 585
R40 B.n153 B.n152 585
R41 B.n154 B.n39 585
R42 B.n156 B.n155 585
R43 B.n157 B.n38 585
R44 B.n159 B.n158 585
R45 B.n160 B.n37 585
R46 B.n162 B.n161 585
R47 B.n163 B.n36 585
R48 B.n165 B.n164 585
R49 B.n166 B.n35 585
R50 B.n168 B.n167 585
R51 B.n169 B.n34 585
R52 B.n171 B.n170 585
R53 B.n172 B.n33 585
R54 B.n174 B.n173 585
R55 B.n175 B.n32 585
R56 B.n177 B.n176 585
R57 B.n178 B.n31 585
R58 B.n180 B.n179 585
R59 B.n181 B.n30 585
R60 B.n183 B.n182 585
R61 B.n230 B.n9 585
R62 B.n229 B.n228 585
R63 B.n227 B.n10 585
R64 B.n226 B.n225 585
R65 B.n224 B.n11 585
R66 B.n223 B.n222 585
R67 B.n221 B.n12 585
R68 B.n220 B.n219 585
R69 B.n218 B.n13 585
R70 B.n217 B.n216 585
R71 B.n215 B.n14 585
R72 B.n214 B.n213 585
R73 B.n212 B.n15 585
R74 B.n211 B.n210 585
R75 B.n209 B.n19 585
R76 B.n208 B.n207 585
R77 B.n206 B.n20 585
R78 B.n205 B.n204 585
R79 B.n203 B.n21 585
R80 B.n202 B.n201 585
R81 B.n199 B.n22 585
R82 B.n198 B.n197 585
R83 B.n196 B.n25 585
R84 B.n195 B.n194 585
R85 B.n193 B.n26 585
R86 B.n192 B.n191 585
R87 B.n190 B.n27 585
R88 B.n189 B.n188 585
R89 B.n187 B.n28 585
R90 B.n186 B.n185 585
R91 B.n184 B.n29 585
R92 B.n232 B.n231 585
R93 B.n233 B.n8 585
R94 B.n235 B.n234 585
R95 B.n236 B.n7 585
R96 B.n238 B.n237 585
R97 B.n239 B.n6 585
R98 B.n241 B.n240 585
R99 B.n242 B.n5 585
R100 B.n244 B.n243 585
R101 B.n245 B.n4 585
R102 B.n247 B.n246 585
R103 B.n248 B.n3 585
R104 B.n250 B.n249 585
R105 B.n251 B.n0 585
R106 B.n2 B.n1 585
R107 B.n71 B.n70 585
R108 B.n73 B.n72 585
R109 B.n74 B.n69 585
R110 B.n76 B.n75 585
R111 B.n77 B.n68 585
R112 B.n79 B.n78 585
R113 B.n80 B.n67 585
R114 B.n82 B.n81 585
R115 B.n83 B.n66 585
R116 B.n85 B.n84 585
R117 B.n86 B.n65 585
R118 B.n88 B.n87 585
R119 B.n89 B.n64 585
R120 B.n91 B.n64 478.086
R121 B.n137 B.n44 478.086
R122 B.n184 B.n183 478.086
R123 B.n232 B.n9 478.086
R124 B.n57 B.t9 303.442
R125 B.n51 B.t0 303.442
R126 B.n23 B.t6 303.442
R127 B.n16 B.t3 303.442
R128 B.n51 B.t1 263.077
R129 B.n23 B.t8 263.077
R130 B.n57 B.t10 263.077
R131 B.n16 B.t5 263.077
R132 B.n253 B.n252 256.663
R133 B.n52 B.t2 249.309
R134 B.n24 B.t7 249.309
R135 B.n58 B.t11 249.308
R136 B.n17 B.t4 249.308
R137 B.n252 B.n251 235.042
R138 B.n252 B.n2 235.042
R139 B.n92 B.n91 163.367
R140 B.n93 B.n92 163.367
R141 B.n93 B.n62 163.367
R142 B.n97 B.n62 163.367
R143 B.n98 B.n97 163.367
R144 B.n99 B.n98 163.367
R145 B.n99 B.n60 163.367
R146 B.n103 B.n60 163.367
R147 B.n104 B.n103 163.367
R148 B.n105 B.n104 163.367
R149 B.n105 B.n56 163.367
R150 B.n110 B.n56 163.367
R151 B.n111 B.n110 163.367
R152 B.n112 B.n111 163.367
R153 B.n112 B.n54 163.367
R154 B.n116 B.n54 163.367
R155 B.n117 B.n116 163.367
R156 B.n118 B.n117 163.367
R157 B.n118 B.n50 163.367
R158 B.n123 B.n50 163.367
R159 B.n124 B.n123 163.367
R160 B.n125 B.n124 163.367
R161 B.n125 B.n48 163.367
R162 B.n129 B.n48 163.367
R163 B.n130 B.n129 163.367
R164 B.n131 B.n130 163.367
R165 B.n131 B.n46 163.367
R166 B.n135 B.n46 163.367
R167 B.n136 B.n135 163.367
R168 B.n137 B.n136 163.367
R169 B.n183 B.n30 163.367
R170 B.n179 B.n30 163.367
R171 B.n179 B.n178 163.367
R172 B.n178 B.n177 163.367
R173 B.n177 B.n32 163.367
R174 B.n173 B.n32 163.367
R175 B.n173 B.n172 163.367
R176 B.n172 B.n171 163.367
R177 B.n171 B.n34 163.367
R178 B.n167 B.n34 163.367
R179 B.n167 B.n166 163.367
R180 B.n166 B.n165 163.367
R181 B.n165 B.n36 163.367
R182 B.n161 B.n36 163.367
R183 B.n161 B.n160 163.367
R184 B.n160 B.n159 163.367
R185 B.n159 B.n38 163.367
R186 B.n155 B.n38 163.367
R187 B.n155 B.n154 163.367
R188 B.n154 B.n153 163.367
R189 B.n153 B.n40 163.367
R190 B.n149 B.n40 163.367
R191 B.n149 B.n148 163.367
R192 B.n148 B.n147 163.367
R193 B.n147 B.n42 163.367
R194 B.n143 B.n42 163.367
R195 B.n143 B.n142 163.367
R196 B.n142 B.n141 163.367
R197 B.n141 B.n44 163.367
R198 B.n228 B.n9 163.367
R199 B.n228 B.n227 163.367
R200 B.n227 B.n226 163.367
R201 B.n226 B.n11 163.367
R202 B.n222 B.n11 163.367
R203 B.n222 B.n221 163.367
R204 B.n221 B.n220 163.367
R205 B.n220 B.n13 163.367
R206 B.n216 B.n13 163.367
R207 B.n216 B.n215 163.367
R208 B.n215 B.n214 163.367
R209 B.n214 B.n15 163.367
R210 B.n210 B.n15 163.367
R211 B.n210 B.n209 163.367
R212 B.n209 B.n208 163.367
R213 B.n208 B.n20 163.367
R214 B.n204 B.n20 163.367
R215 B.n204 B.n203 163.367
R216 B.n203 B.n202 163.367
R217 B.n202 B.n22 163.367
R218 B.n197 B.n22 163.367
R219 B.n197 B.n196 163.367
R220 B.n196 B.n195 163.367
R221 B.n195 B.n26 163.367
R222 B.n191 B.n26 163.367
R223 B.n191 B.n190 163.367
R224 B.n190 B.n189 163.367
R225 B.n189 B.n28 163.367
R226 B.n185 B.n28 163.367
R227 B.n185 B.n184 163.367
R228 B.n233 B.n232 163.367
R229 B.n234 B.n233 163.367
R230 B.n234 B.n7 163.367
R231 B.n238 B.n7 163.367
R232 B.n239 B.n238 163.367
R233 B.n240 B.n239 163.367
R234 B.n240 B.n5 163.367
R235 B.n244 B.n5 163.367
R236 B.n245 B.n244 163.367
R237 B.n246 B.n245 163.367
R238 B.n246 B.n3 163.367
R239 B.n250 B.n3 163.367
R240 B.n251 B.n250 163.367
R241 B.n70 B.n2 163.367
R242 B.n73 B.n70 163.367
R243 B.n74 B.n73 163.367
R244 B.n75 B.n74 163.367
R245 B.n75 B.n68 163.367
R246 B.n79 B.n68 163.367
R247 B.n80 B.n79 163.367
R248 B.n81 B.n80 163.367
R249 B.n81 B.n66 163.367
R250 B.n85 B.n66 163.367
R251 B.n86 B.n85 163.367
R252 B.n87 B.n86 163.367
R253 B.n87 B.n64 163.367
R254 B.n107 B.n58 59.5399
R255 B.n121 B.n52 59.5399
R256 B.n200 B.n24 59.5399
R257 B.n18 B.n17 59.5399
R258 B.n231 B.n230 31.0639
R259 B.n182 B.n29 31.0639
R260 B.n139 B.n138 31.0639
R261 B.n90 B.n89 31.0639
R262 B B.n253 18.0485
R263 B.n58 B.n57 13.7702
R264 B.n52 B.n51 13.7702
R265 B.n24 B.n23 13.7702
R266 B.n17 B.n16 13.7702
R267 B.n231 B.n8 10.6151
R268 B.n235 B.n8 10.6151
R269 B.n236 B.n235 10.6151
R270 B.n237 B.n236 10.6151
R271 B.n237 B.n6 10.6151
R272 B.n241 B.n6 10.6151
R273 B.n242 B.n241 10.6151
R274 B.n243 B.n242 10.6151
R275 B.n243 B.n4 10.6151
R276 B.n247 B.n4 10.6151
R277 B.n248 B.n247 10.6151
R278 B.n249 B.n248 10.6151
R279 B.n249 B.n0 10.6151
R280 B.n230 B.n229 10.6151
R281 B.n229 B.n10 10.6151
R282 B.n225 B.n10 10.6151
R283 B.n225 B.n224 10.6151
R284 B.n224 B.n223 10.6151
R285 B.n223 B.n12 10.6151
R286 B.n219 B.n12 10.6151
R287 B.n219 B.n218 10.6151
R288 B.n218 B.n217 10.6151
R289 B.n217 B.n14 10.6151
R290 B.n213 B.n212 10.6151
R291 B.n212 B.n211 10.6151
R292 B.n211 B.n19 10.6151
R293 B.n207 B.n19 10.6151
R294 B.n207 B.n206 10.6151
R295 B.n206 B.n205 10.6151
R296 B.n205 B.n21 10.6151
R297 B.n201 B.n21 10.6151
R298 B.n199 B.n198 10.6151
R299 B.n198 B.n25 10.6151
R300 B.n194 B.n25 10.6151
R301 B.n194 B.n193 10.6151
R302 B.n193 B.n192 10.6151
R303 B.n192 B.n27 10.6151
R304 B.n188 B.n27 10.6151
R305 B.n188 B.n187 10.6151
R306 B.n187 B.n186 10.6151
R307 B.n186 B.n29 10.6151
R308 B.n182 B.n181 10.6151
R309 B.n181 B.n180 10.6151
R310 B.n180 B.n31 10.6151
R311 B.n176 B.n31 10.6151
R312 B.n176 B.n175 10.6151
R313 B.n175 B.n174 10.6151
R314 B.n174 B.n33 10.6151
R315 B.n170 B.n33 10.6151
R316 B.n170 B.n169 10.6151
R317 B.n169 B.n168 10.6151
R318 B.n168 B.n35 10.6151
R319 B.n164 B.n35 10.6151
R320 B.n164 B.n163 10.6151
R321 B.n163 B.n162 10.6151
R322 B.n162 B.n37 10.6151
R323 B.n158 B.n37 10.6151
R324 B.n158 B.n157 10.6151
R325 B.n157 B.n156 10.6151
R326 B.n156 B.n39 10.6151
R327 B.n152 B.n39 10.6151
R328 B.n152 B.n151 10.6151
R329 B.n151 B.n150 10.6151
R330 B.n150 B.n41 10.6151
R331 B.n146 B.n41 10.6151
R332 B.n146 B.n145 10.6151
R333 B.n145 B.n144 10.6151
R334 B.n144 B.n43 10.6151
R335 B.n140 B.n43 10.6151
R336 B.n140 B.n139 10.6151
R337 B.n71 B.n1 10.6151
R338 B.n72 B.n71 10.6151
R339 B.n72 B.n69 10.6151
R340 B.n76 B.n69 10.6151
R341 B.n77 B.n76 10.6151
R342 B.n78 B.n77 10.6151
R343 B.n78 B.n67 10.6151
R344 B.n82 B.n67 10.6151
R345 B.n83 B.n82 10.6151
R346 B.n84 B.n83 10.6151
R347 B.n84 B.n65 10.6151
R348 B.n88 B.n65 10.6151
R349 B.n89 B.n88 10.6151
R350 B.n90 B.n63 10.6151
R351 B.n94 B.n63 10.6151
R352 B.n95 B.n94 10.6151
R353 B.n96 B.n95 10.6151
R354 B.n96 B.n61 10.6151
R355 B.n100 B.n61 10.6151
R356 B.n101 B.n100 10.6151
R357 B.n102 B.n101 10.6151
R358 B.n102 B.n59 10.6151
R359 B.n106 B.n59 10.6151
R360 B.n109 B.n108 10.6151
R361 B.n109 B.n55 10.6151
R362 B.n113 B.n55 10.6151
R363 B.n114 B.n113 10.6151
R364 B.n115 B.n114 10.6151
R365 B.n115 B.n53 10.6151
R366 B.n119 B.n53 10.6151
R367 B.n120 B.n119 10.6151
R368 B.n122 B.n49 10.6151
R369 B.n126 B.n49 10.6151
R370 B.n127 B.n126 10.6151
R371 B.n128 B.n127 10.6151
R372 B.n128 B.n47 10.6151
R373 B.n132 B.n47 10.6151
R374 B.n133 B.n132 10.6151
R375 B.n134 B.n133 10.6151
R376 B.n134 B.n45 10.6151
R377 B.n138 B.n45 10.6151
R378 B.n253 B.n0 8.11757
R379 B.n253 B.n1 8.11757
R380 B.n213 B.n18 7.18099
R381 B.n201 B.n200 7.18099
R382 B.n108 B.n107 7.18099
R383 B.n121 B.n120 7.18099
R384 B.n18 B.n14 3.43465
R385 B.n200 B.n199 3.43465
R386 B.n107 B.n106 3.43465
R387 B.n122 B.n121 3.43465
R388 VP.n1 VP.t2 221.339
R389 VP.n1 VP.t3 221.339
R390 VP.n0 VP.t1 221.339
R391 VP.n0 VP.t0 221.339
R392 VP.n2 VP.n0 192.915
R393 VP.n2 VP.n1 161.3
R394 VP VP.n2 0.0516364
R395 VDD1 VDD1.n1 277.731
R396 VDD1 VDD1.n0 250.429
R397 VDD1.n0 VDD1.t0 22.1127
R398 VDD1.n0 VDD1.t1 22.1127
R399 VDD1.n1 VDD1.t2 22.1127
R400 VDD1.n1 VDD1.t3 22.1127
R401 VTAIL.n5 VTAIL.t7 255.804
R402 VTAIL.n4 VTAIL.t0 255.804
R403 VTAIL.n3 VTAIL.t1 255.804
R404 VTAIL.n7 VTAIL.t3 255.804
R405 VTAIL.n0 VTAIL.t2 255.804
R406 VTAIL.n1 VTAIL.t5 255.804
R407 VTAIL.n2 VTAIL.t4 255.804
R408 VTAIL.n6 VTAIL.t6 255.804
R409 VTAIL.n7 VTAIL.n6 14.2634
R410 VTAIL.n3 VTAIL.n2 14.2634
R411 VTAIL.n4 VTAIL.n3 0.612569
R412 VTAIL.n6 VTAIL.n5 0.612569
R413 VTAIL.n2 VTAIL.n1 0.612569
R414 VTAIL.n5 VTAIL.n4 0.470328
R415 VTAIL.n1 VTAIL.n0 0.470328
R416 VTAIL VTAIL.n0 0.364724
R417 VTAIL VTAIL.n7 0.248345
R418 VN.n0 VN.t1 221.339
R419 VN.n0 VN.t0 221.339
R420 VN.n1 VN.t2 221.339
R421 VN.n1 VN.t3 221.339
R422 VN VN.n1 193.294
R423 VN VN.n0 161.351
R424 VDD2.n2 VDD2.n0 277.205
R425 VDD2.n2 VDD2.n1 250.37
R426 VDD2.n1 VDD2.t0 22.1127
R427 VDD2.n1 VDD2.t1 22.1127
R428 VDD2.n0 VDD2.t3 22.1127
R429 VDD2.n0 VDD2.t2 22.1127
R430 VDD2 VDD2.n2 0.0586897
C0 VTAIL VDD1 2.19817f
C1 VDD2 VN 0.534123f
C2 w_n1396_n1266# VP 1.86825f
C3 B VP 0.817443f
C4 VN VTAIL 0.588957f
C5 VDD2 w_n1396_n1266# 0.705478f
C6 VDD2 B 0.601045f
C7 VTAIL w_n1396_n1266# 1.37948f
C8 VTAIL B 0.838318f
C9 VN VDD1 0.154488f
C10 VDD2 VP 0.261318f
C11 w_n1396_n1266# VDD1 0.697998f
C12 VDD1 B 0.583796f
C13 VTAIL VP 0.603064f
C14 VN w_n1396_n1266# 1.70064f
C15 VDD2 VTAIL 2.23749f
C16 VN B 0.540267f
C17 VDD1 VP 0.640019f
C18 w_n1396_n1266# B 3.54282f
C19 VDD2 VDD1 0.495772f
C20 VN VP 2.64102f
C21 VDD2 VSUBS 0.361172f
C22 VDD1 VSUBS 2.315188f
C23 VTAIL VSUBS 0.259774f
C24 VN VSUBS 3.09805f
C25 VP VSUBS 0.662095f
C26 B VSUBS 1.396699f
C27 w_n1396_n1266# VSUBS 22.6655f
C28 VDD2.t3 VSUBS 0.025649f
C29 VDD2.t2 VSUBS 0.025649f
C30 VDD2.n0 VSUBS 0.169465f
C31 VDD2.t0 VSUBS 0.025649f
C32 VDD2.t1 VSUBS 0.025649f
C33 VDD2.n1 VSUBS 0.097841f
C34 VDD2.n2 VSUBS 1.7818f
C35 VN.t0 VSUBS 0.077836f
C36 VN.t1 VSUBS 0.077836f
C37 VN.n0 VSUBS 0.111546f
C38 VN.t3 VSUBS 0.077836f
C39 VN.t2 VSUBS 0.077836f
C40 VN.n1 VSUBS 0.278465f
C41 VTAIL.t2 VSUBS 0.126922f
C42 VTAIL.n0 VSUBS 0.228711f
C43 VTAIL.t5 VSUBS 0.126922f
C44 VTAIL.n1 VSUBS 0.244408f
C45 VTAIL.t4 VSUBS 0.126922f
C46 VTAIL.n2 VSUBS 0.601749f
C47 VTAIL.t1 VSUBS 0.126922f
C48 VTAIL.n3 VSUBS 0.601749f
C49 VTAIL.t0 VSUBS 0.126922f
C50 VTAIL.n4 VSUBS 0.244408f
C51 VTAIL.t7 VSUBS 0.126922f
C52 VTAIL.n5 VSUBS 0.244408f
C53 VTAIL.t6 VSUBS 0.126922f
C54 VTAIL.n6 VSUBS 0.601749f
C55 VTAIL.t3 VSUBS 0.126922f
C56 VTAIL.n7 VSUBS 0.578682f
C57 VDD1.t0 VSUBS 0.024732f
C58 VDD1.t1 VSUBS 0.024732f
C59 VDD1.n0 VSUBS 0.094402f
C60 VDD1.t2 VSUBS 0.024732f
C61 VDD1.t3 VSUBS 0.024732f
C62 VDD1.n1 VSUBS 0.168983f
C63 VP.t0 VSUBS 0.079554f
C64 VP.t1 VSUBS 0.079554f
C65 VP.n0 VSUBS 0.278429f
C66 VP.t3 VSUBS 0.079554f
C67 VP.t2 VSUBS 0.079554f
C68 VP.n1 VSUBS 0.113992f
C69 VP.n2 VSUBS 1.86534f
C70 B.n0 VSUBS 0.008269f
C71 B.n1 VSUBS 0.008269f
C72 B.n2 VSUBS 0.012229f
C73 B.n3 VSUBS 0.009371f
C74 B.n4 VSUBS 0.009371f
C75 B.n5 VSUBS 0.009371f
C76 B.n6 VSUBS 0.009371f
C77 B.n7 VSUBS 0.009371f
C78 B.n8 VSUBS 0.009371f
C79 B.n9 VSUBS 0.021664f
C80 B.n10 VSUBS 0.009371f
C81 B.n11 VSUBS 0.009371f
C82 B.n12 VSUBS 0.009371f
C83 B.n13 VSUBS 0.009371f
C84 B.n14 VSUBS 0.006202f
C85 B.n15 VSUBS 0.009371f
C86 B.t4 VSUBS 0.039867f
C87 B.t5 VSUBS 0.042192f
C88 B.t3 VSUBS 0.036183f
C89 B.n16 VSUBS 0.058668f
C90 B.n17 VSUBS 0.057797f
C91 B.n18 VSUBS 0.021713f
C92 B.n19 VSUBS 0.009371f
C93 B.n20 VSUBS 0.009371f
C94 B.n21 VSUBS 0.009371f
C95 B.n22 VSUBS 0.009371f
C96 B.t7 VSUBS 0.039867f
C97 B.t8 VSUBS 0.042192f
C98 B.t6 VSUBS 0.036183f
C99 B.n23 VSUBS 0.058668f
C100 B.n24 VSUBS 0.057797f
C101 B.n25 VSUBS 0.009371f
C102 B.n26 VSUBS 0.009371f
C103 B.n27 VSUBS 0.009371f
C104 B.n28 VSUBS 0.009371f
C105 B.n29 VSUBS 0.021664f
C106 B.n30 VSUBS 0.009371f
C107 B.n31 VSUBS 0.009371f
C108 B.n32 VSUBS 0.009371f
C109 B.n33 VSUBS 0.009371f
C110 B.n34 VSUBS 0.009371f
C111 B.n35 VSUBS 0.009371f
C112 B.n36 VSUBS 0.009371f
C113 B.n37 VSUBS 0.009371f
C114 B.n38 VSUBS 0.009371f
C115 B.n39 VSUBS 0.009371f
C116 B.n40 VSUBS 0.009371f
C117 B.n41 VSUBS 0.009371f
C118 B.n42 VSUBS 0.009371f
C119 B.n43 VSUBS 0.009371f
C120 B.n44 VSUBS 0.020783f
C121 B.n45 VSUBS 0.009371f
C122 B.n46 VSUBS 0.009371f
C123 B.n47 VSUBS 0.009371f
C124 B.n48 VSUBS 0.009371f
C125 B.n49 VSUBS 0.009371f
C126 B.n50 VSUBS 0.009371f
C127 B.t2 VSUBS 0.039867f
C128 B.t1 VSUBS 0.042192f
C129 B.t0 VSUBS 0.036183f
C130 B.n51 VSUBS 0.058668f
C131 B.n52 VSUBS 0.057797f
C132 B.n53 VSUBS 0.009371f
C133 B.n54 VSUBS 0.009371f
C134 B.n55 VSUBS 0.009371f
C135 B.n56 VSUBS 0.009371f
C136 B.t11 VSUBS 0.039867f
C137 B.t10 VSUBS 0.042192f
C138 B.t9 VSUBS 0.036183f
C139 B.n57 VSUBS 0.058668f
C140 B.n58 VSUBS 0.057797f
C141 B.n59 VSUBS 0.009371f
C142 B.n60 VSUBS 0.009371f
C143 B.n61 VSUBS 0.009371f
C144 B.n62 VSUBS 0.009371f
C145 B.n63 VSUBS 0.009371f
C146 B.n64 VSUBS 0.020783f
C147 B.n65 VSUBS 0.009371f
C148 B.n66 VSUBS 0.009371f
C149 B.n67 VSUBS 0.009371f
C150 B.n68 VSUBS 0.009371f
C151 B.n69 VSUBS 0.009371f
C152 B.n70 VSUBS 0.009371f
C153 B.n71 VSUBS 0.009371f
C154 B.n72 VSUBS 0.009371f
C155 B.n73 VSUBS 0.009371f
C156 B.n74 VSUBS 0.009371f
C157 B.n75 VSUBS 0.009371f
C158 B.n76 VSUBS 0.009371f
C159 B.n77 VSUBS 0.009371f
C160 B.n78 VSUBS 0.009371f
C161 B.n79 VSUBS 0.009371f
C162 B.n80 VSUBS 0.009371f
C163 B.n81 VSUBS 0.009371f
C164 B.n82 VSUBS 0.009371f
C165 B.n83 VSUBS 0.009371f
C166 B.n84 VSUBS 0.009371f
C167 B.n85 VSUBS 0.009371f
C168 B.n86 VSUBS 0.009371f
C169 B.n87 VSUBS 0.009371f
C170 B.n88 VSUBS 0.009371f
C171 B.n89 VSUBS 0.020783f
C172 B.n90 VSUBS 0.021664f
C173 B.n91 VSUBS 0.021664f
C174 B.n92 VSUBS 0.009371f
C175 B.n93 VSUBS 0.009371f
C176 B.n94 VSUBS 0.009371f
C177 B.n95 VSUBS 0.009371f
C178 B.n96 VSUBS 0.009371f
C179 B.n97 VSUBS 0.009371f
C180 B.n98 VSUBS 0.009371f
C181 B.n99 VSUBS 0.009371f
C182 B.n100 VSUBS 0.009371f
C183 B.n101 VSUBS 0.009371f
C184 B.n102 VSUBS 0.009371f
C185 B.n103 VSUBS 0.009371f
C186 B.n104 VSUBS 0.009371f
C187 B.n105 VSUBS 0.009371f
C188 B.n106 VSUBS 0.006202f
C189 B.n107 VSUBS 0.021713f
C190 B.n108 VSUBS 0.007855f
C191 B.n109 VSUBS 0.009371f
C192 B.n110 VSUBS 0.009371f
C193 B.n111 VSUBS 0.009371f
C194 B.n112 VSUBS 0.009371f
C195 B.n113 VSUBS 0.009371f
C196 B.n114 VSUBS 0.009371f
C197 B.n115 VSUBS 0.009371f
C198 B.n116 VSUBS 0.009371f
C199 B.n117 VSUBS 0.009371f
C200 B.n118 VSUBS 0.009371f
C201 B.n119 VSUBS 0.009371f
C202 B.n120 VSUBS 0.007855f
C203 B.n121 VSUBS 0.021713f
C204 B.n122 VSUBS 0.006202f
C205 B.n123 VSUBS 0.009371f
C206 B.n124 VSUBS 0.009371f
C207 B.n125 VSUBS 0.009371f
C208 B.n126 VSUBS 0.009371f
C209 B.n127 VSUBS 0.009371f
C210 B.n128 VSUBS 0.009371f
C211 B.n129 VSUBS 0.009371f
C212 B.n130 VSUBS 0.009371f
C213 B.n131 VSUBS 0.009371f
C214 B.n132 VSUBS 0.009371f
C215 B.n133 VSUBS 0.009371f
C216 B.n134 VSUBS 0.009371f
C217 B.n135 VSUBS 0.009371f
C218 B.n136 VSUBS 0.009371f
C219 B.n137 VSUBS 0.021664f
C220 B.n138 VSUBS 0.020499f
C221 B.n139 VSUBS 0.021948f
C222 B.n140 VSUBS 0.009371f
C223 B.n141 VSUBS 0.009371f
C224 B.n142 VSUBS 0.009371f
C225 B.n143 VSUBS 0.009371f
C226 B.n144 VSUBS 0.009371f
C227 B.n145 VSUBS 0.009371f
C228 B.n146 VSUBS 0.009371f
C229 B.n147 VSUBS 0.009371f
C230 B.n148 VSUBS 0.009371f
C231 B.n149 VSUBS 0.009371f
C232 B.n150 VSUBS 0.009371f
C233 B.n151 VSUBS 0.009371f
C234 B.n152 VSUBS 0.009371f
C235 B.n153 VSUBS 0.009371f
C236 B.n154 VSUBS 0.009371f
C237 B.n155 VSUBS 0.009371f
C238 B.n156 VSUBS 0.009371f
C239 B.n157 VSUBS 0.009371f
C240 B.n158 VSUBS 0.009371f
C241 B.n159 VSUBS 0.009371f
C242 B.n160 VSUBS 0.009371f
C243 B.n161 VSUBS 0.009371f
C244 B.n162 VSUBS 0.009371f
C245 B.n163 VSUBS 0.009371f
C246 B.n164 VSUBS 0.009371f
C247 B.n165 VSUBS 0.009371f
C248 B.n166 VSUBS 0.009371f
C249 B.n167 VSUBS 0.009371f
C250 B.n168 VSUBS 0.009371f
C251 B.n169 VSUBS 0.009371f
C252 B.n170 VSUBS 0.009371f
C253 B.n171 VSUBS 0.009371f
C254 B.n172 VSUBS 0.009371f
C255 B.n173 VSUBS 0.009371f
C256 B.n174 VSUBS 0.009371f
C257 B.n175 VSUBS 0.009371f
C258 B.n176 VSUBS 0.009371f
C259 B.n177 VSUBS 0.009371f
C260 B.n178 VSUBS 0.009371f
C261 B.n179 VSUBS 0.009371f
C262 B.n180 VSUBS 0.009371f
C263 B.n181 VSUBS 0.009371f
C264 B.n182 VSUBS 0.020783f
C265 B.n183 VSUBS 0.020783f
C266 B.n184 VSUBS 0.021664f
C267 B.n185 VSUBS 0.009371f
C268 B.n186 VSUBS 0.009371f
C269 B.n187 VSUBS 0.009371f
C270 B.n188 VSUBS 0.009371f
C271 B.n189 VSUBS 0.009371f
C272 B.n190 VSUBS 0.009371f
C273 B.n191 VSUBS 0.009371f
C274 B.n192 VSUBS 0.009371f
C275 B.n193 VSUBS 0.009371f
C276 B.n194 VSUBS 0.009371f
C277 B.n195 VSUBS 0.009371f
C278 B.n196 VSUBS 0.009371f
C279 B.n197 VSUBS 0.009371f
C280 B.n198 VSUBS 0.009371f
C281 B.n199 VSUBS 0.006202f
C282 B.n200 VSUBS 0.021713f
C283 B.n201 VSUBS 0.007855f
C284 B.n202 VSUBS 0.009371f
C285 B.n203 VSUBS 0.009371f
C286 B.n204 VSUBS 0.009371f
C287 B.n205 VSUBS 0.009371f
C288 B.n206 VSUBS 0.009371f
C289 B.n207 VSUBS 0.009371f
C290 B.n208 VSUBS 0.009371f
C291 B.n209 VSUBS 0.009371f
C292 B.n210 VSUBS 0.009371f
C293 B.n211 VSUBS 0.009371f
C294 B.n212 VSUBS 0.009371f
C295 B.n213 VSUBS 0.007855f
C296 B.n214 VSUBS 0.009371f
C297 B.n215 VSUBS 0.009371f
C298 B.n216 VSUBS 0.009371f
C299 B.n217 VSUBS 0.009371f
C300 B.n218 VSUBS 0.009371f
C301 B.n219 VSUBS 0.009371f
C302 B.n220 VSUBS 0.009371f
C303 B.n221 VSUBS 0.009371f
C304 B.n222 VSUBS 0.009371f
C305 B.n223 VSUBS 0.009371f
C306 B.n224 VSUBS 0.009371f
C307 B.n225 VSUBS 0.009371f
C308 B.n226 VSUBS 0.009371f
C309 B.n227 VSUBS 0.009371f
C310 B.n228 VSUBS 0.009371f
C311 B.n229 VSUBS 0.009371f
C312 B.n230 VSUBS 0.021664f
C313 B.n231 VSUBS 0.020783f
C314 B.n232 VSUBS 0.020783f
C315 B.n233 VSUBS 0.009371f
C316 B.n234 VSUBS 0.009371f
C317 B.n235 VSUBS 0.009371f
C318 B.n236 VSUBS 0.009371f
C319 B.n237 VSUBS 0.009371f
C320 B.n238 VSUBS 0.009371f
C321 B.n239 VSUBS 0.009371f
C322 B.n240 VSUBS 0.009371f
C323 B.n241 VSUBS 0.009371f
C324 B.n242 VSUBS 0.009371f
C325 B.n243 VSUBS 0.009371f
C326 B.n244 VSUBS 0.009371f
C327 B.n245 VSUBS 0.009371f
C328 B.n246 VSUBS 0.009371f
C329 B.n247 VSUBS 0.009371f
C330 B.n248 VSUBS 0.009371f
C331 B.n249 VSUBS 0.009371f
C332 B.n250 VSUBS 0.009371f
C333 B.n251 VSUBS 0.012229f
C334 B.n252 VSUBS 0.013027f
C335 B.n253 VSUBS 0.025906f
.ends

