* NGSPICE file created from diff_pair_sample_0231.ext - technology: sky130A

.subckt diff_pair_sample_0231 VTAIL VN VP B VDD2 VDD1
X0 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=0 ps=0 w=9.31 l=1.3
X1 VTAIL.t19 VP.t0 VDD1.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X2 VTAIL.t3 VN.t0 VDD2.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X3 VDD2.t8 VN.t1 VTAIL.t6 B.t4 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=1.53615 ps=9.64 w=9.31 l=1.3
X4 VTAIL.t18 VP.t1 VDD1.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X5 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=0 ps=0 w=9.31 l=1.3
X6 VDD1.t2 VP.t2 VTAIL.t17 B.t2 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=3.6309 ps=19.4 w=9.31 l=1.3
X7 VTAIL.t7 VN.t2 VDD2.t7 B.t6 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X8 VDD1.t9 VP.t3 VTAIL.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=3.6309 ps=19.4 w=9.31 l=1.3
X9 VTAIL.t15 VP.t4 VDD1.t5 B.t6 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X10 VDD2.t6 VN.t3 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=1.53615 ps=9.64 w=9.31 l=1.3
X11 VDD1.t1 VP.t5 VTAIL.t14 B.t4 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=1.53615 ps=9.64 w=9.31 l=1.3
X12 VDD2.t5 VN.t4 VTAIL.t4 B.t2 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=3.6309 ps=19.4 w=9.31 l=1.3
X13 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=0 ps=0 w=9.31 l=1.3
X14 VDD1.t6 VP.t6 VTAIL.t13 B.t8 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=1.53615 ps=9.64 w=9.31 l=1.3
X15 VTAIL.t2 VN.t5 VDD2.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X16 VTAIL.t12 VP.t7 VDD1.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X17 VDD1.t8 VP.t8 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X18 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6309 pd=19.4 as=0 ps=0 w=9.31 l=1.3
X19 VTAIL.t1 VN.t6 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X20 VDD2.t2 VN.t7 VTAIL.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=3.6309 ps=19.4 w=9.31 l=1.3
X21 VDD2.t1 VN.t8 VTAIL.t5 B.t9 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X22 VDD2.t0 VN.t9 VTAIL.t9 B.t3 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
X23 VDD1.t0 VP.t9 VTAIL.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=1.53615 pd=9.64 as=1.53615 ps=9.64 w=9.31 l=1.3
R0 B.n694 B.n693 585
R1 B.n695 B.n694 585
R2 B.n265 B.n108 585
R3 B.n264 B.n263 585
R4 B.n262 B.n261 585
R5 B.n260 B.n259 585
R6 B.n258 B.n257 585
R7 B.n256 B.n255 585
R8 B.n254 B.n253 585
R9 B.n252 B.n251 585
R10 B.n250 B.n249 585
R11 B.n248 B.n247 585
R12 B.n246 B.n245 585
R13 B.n244 B.n243 585
R14 B.n242 B.n241 585
R15 B.n240 B.n239 585
R16 B.n238 B.n237 585
R17 B.n236 B.n235 585
R18 B.n234 B.n233 585
R19 B.n232 B.n231 585
R20 B.n230 B.n229 585
R21 B.n228 B.n227 585
R22 B.n226 B.n225 585
R23 B.n224 B.n223 585
R24 B.n222 B.n221 585
R25 B.n220 B.n219 585
R26 B.n218 B.n217 585
R27 B.n216 B.n215 585
R28 B.n214 B.n213 585
R29 B.n212 B.n211 585
R30 B.n210 B.n209 585
R31 B.n208 B.n207 585
R32 B.n206 B.n205 585
R33 B.n204 B.n203 585
R34 B.n202 B.n201 585
R35 B.n199 B.n198 585
R36 B.n197 B.n196 585
R37 B.n195 B.n194 585
R38 B.n193 B.n192 585
R39 B.n191 B.n190 585
R40 B.n189 B.n188 585
R41 B.n187 B.n186 585
R42 B.n185 B.n184 585
R43 B.n183 B.n182 585
R44 B.n181 B.n180 585
R45 B.n179 B.n178 585
R46 B.n177 B.n176 585
R47 B.n175 B.n174 585
R48 B.n173 B.n172 585
R49 B.n171 B.n170 585
R50 B.n169 B.n168 585
R51 B.n167 B.n166 585
R52 B.n165 B.n164 585
R53 B.n163 B.n162 585
R54 B.n161 B.n160 585
R55 B.n159 B.n158 585
R56 B.n157 B.n156 585
R57 B.n155 B.n154 585
R58 B.n153 B.n152 585
R59 B.n151 B.n150 585
R60 B.n149 B.n148 585
R61 B.n147 B.n146 585
R62 B.n145 B.n144 585
R63 B.n143 B.n142 585
R64 B.n141 B.n140 585
R65 B.n139 B.n138 585
R66 B.n137 B.n136 585
R67 B.n135 B.n134 585
R68 B.n133 B.n132 585
R69 B.n131 B.n130 585
R70 B.n129 B.n128 585
R71 B.n127 B.n126 585
R72 B.n125 B.n124 585
R73 B.n123 B.n122 585
R74 B.n121 B.n120 585
R75 B.n119 B.n118 585
R76 B.n117 B.n116 585
R77 B.n115 B.n114 585
R78 B.n692 B.n69 585
R79 B.n696 B.n69 585
R80 B.n691 B.n68 585
R81 B.n697 B.n68 585
R82 B.n690 B.n689 585
R83 B.n689 B.n64 585
R84 B.n688 B.n63 585
R85 B.n703 B.n63 585
R86 B.n687 B.n62 585
R87 B.n704 B.n62 585
R88 B.n686 B.n61 585
R89 B.n705 B.n61 585
R90 B.n685 B.n684 585
R91 B.n684 B.n57 585
R92 B.n683 B.n56 585
R93 B.n711 B.n56 585
R94 B.n682 B.n55 585
R95 B.n712 B.n55 585
R96 B.n681 B.n54 585
R97 B.n713 B.n54 585
R98 B.n680 B.n679 585
R99 B.n679 B.n50 585
R100 B.n678 B.n49 585
R101 B.n719 B.n49 585
R102 B.n677 B.n48 585
R103 B.n720 B.n48 585
R104 B.n676 B.n47 585
R105 B.n721 B.n47 585
R106 B.n675 B.n674 585
R107 B.n674 B.n43 585
R108 B.n673 B.n42 585
R109 B.n727 B.n42 585
R110 B.n672 B.n41 585
R111 B.n728 B.n41 585
R112 B.n671 B.n40 585
R113 B.n729 B.n40 585
R114 B.n670 B.n669 585
R115 B.n669 B.n39 585
R116 B.n668 B.n35 585
R117 B.n735 B.n35 585
R118 B.n667 B.n34 585
R119 B.n736 B.n34 585
R120 B.n666 B.n33 585
R121 B.n737 B.n33 585
R122 B.n665 B.n664 585
R123 B.n664 B.n29 585
R124 B.n663 B.n28 585
R125 B.n743 B.n28 585
R126 B.n662 B.n27 585
R127 B.n744 B.n27 585
R128 B.n661 B.n26 585
R129 B.n745 B.n26 585
R130 B.n660 B.n659 585
R131 B.n659 B.n22 585
R132 B.n658 B.n21 585
R133 B.n751 B.n21 585
R134 B.n657 B.n20 585
R135 B.n752 B.n20 585
R136 B.n656 B.n19 585
R137 B.n753 B.n19 585
R138 B.n655 B.n654 585
R139 B.n654 B.n15 585
R140 B.n653 B.n14 585
R141 B.n759 B.n14 585
R142 B.n652 B.n13 585
R143 B.n760 B.n13 585
R144 B.n651 B.n12 585
R145 B.t4 B.n12 585
R146 B.n650 B.n649 585
R147 B.n649 B.n8 585
R148 B.n648 B.n7 585
R149 B.n766 B.n7 585
R150 B.n647 B.n6 585
R151 B.n767 B.n6 585
R152 B.n646 B.n5 585
R153 B.n768 B.n5 585
R154 B.n645 B.n644 585
R155 B.n644 B.n4 585
R156 B.n643 B.n266 585
R157 B.n643 B.n642 585
R158 B.n634 B.n267 585
R159 B.n268 B.n267 585
R160 B.n636 B.n635 585
R161 B.t2 B.n636 585
R162 B.n633 B.n273 585
R163 B.n273 B.n272 585
R164 B.n632 B.n631 585
R165 B.n631 B.n630 585
R166 B.n275 B.n274 585
R167 B.n276 B.n275 585
R168 B.n623 B.n622 585
R169 B.n624 B.n623 585
R170 B.n621 B.n280 585
R171 B.n284 B.n280 585
R172 B.n620 B.n619 585
R173 B.n619 B.n618 585
R174 B.n282 B.n281 585
R175 B.n283 B.n282 585
R176 B.n611 B.n610 585
R177 B.n612 B.n611 585
R178 B.n609 B.n289 585
R179 B.n289 B.n288 585
R180 B.n608 B.n607 585
R181 B.n607 B.n606 585
R182 B.n291 B.n290 585
R183 B.n292 B.n291 585
R184 B.n599 B.n598 585
R185 B.n600 B.n599 585
R186 B.n597 B.n297 585
R187 B.n297 B.n296 585
R188 B.n596 B.n595 585
R189 B.n595 B.n594 585
R190 B.n299 B.n298 585
R191 B.n587 B.n299 585
R192 B.n586 B.n585 585
R193 B.n588 B.n586 585
R194 B.n584 B.n304 585
R195 B.n304 B.n303 585
R196 B.n583 B.n582 585
R197 B.n582 B.n581 585
R198 B.n306 B.n305 585
R199 B.n307 B.n306 585
R200 B.n574 B.n573 585
R201 B.n575 B.n574 585
R202 B.n572 B.n312 585
R203 B.n312 B.n311 585
R204 B.n571 B.n570 585
R205 B.n570 B.n569 585
R206 B.n314 B.n313 585
R207 B.n315 B.n314 585
R208 B.n562 B.n561 585
R209 B.n563 B.n562 585
R210 B.n560 B.n320 585
R211 B.n320 B.n319 585
R212 B.n559 B.n558 585
R213 B.n558 B.n557 585
R214 B.n322 B.n321 585
R215 B.n323 B.n322 585
R216 B.n550 B.n549 585
R217 B.n551 B.n550 585
R218 B.n548 B.n328 585
R219 B.n328 B.n327 585
R220 B.n547 B.n546 585
R221 B.n546 B.n545 585
R222 B.n330 B.n329 585
R223 B.n331 B.n330 585
R224 B.n538 B.n537 585
R225 B.n539 B.n538 585
R226 B.n536 B.n336 585
R227 B.n336 B.n335 585
R228 B.n530 B.n529 585
R229 B.n528 B.n376 585
R230 B.n527 B.n375 585
R231 B.n532 B.n375 585
R232 B.n526 B.n525 585
R233 B.n524 B.n523 585
R234 B.n522 B.n521 585
R235 B.n520 B.n519 585
R236 B.n518 B.n517 585
R237 B.n516 B.n515 585
R238 B.n514 B.n513 585
R239 B.n512 B.n511 585
R240 B.n510 B.n509 585
R241 B.n508 B.n507 585
R242 B.n506 B.n505 585
R243 B.n504 B.n503 585
R244 B.n502 B.n501 585
R245 B.n500 B.n499 585
R246 B.n498 B.n497 585
R247 B.n496 B.n495 585
R248 B.n494 B.n493 585
R249 B.n492 B.n491 585
R250 B.n490 B.n489 585
R251 B.n488 B.n487 585
R252 B.n486 B.n485 585
R253 B.n484 B.n483 585
R254 B.n482 B.n481 585
R255 B.n480 B.n479 585
R256 B.n478 B.n477 585
R257 B.n476 B.n475 585
R258 B.n474 B.n473 585
R259 B.n472 B.n471 585
R260 B.n470 B.n469 585
R261 B.n468 B.n467 585
R262 B.n466 B.n465 585
R263 B.n463 B.n462 585
R264 B.n461 B.n460 585
R265 B.n459 B.n458 585
R266 B.n457 B.n456 585
R267 B.n455 B.n454 585
R268 B.n453 B.n452 585
R269 B.n451 B.n450 585
R270 B.n449 B.n448 585
R271 B.n447 B.n446 585
R272 B.n445 B.n444 585
R273 B.n443 B.n442 585
R274 B.n441 B.n440 585
R275 B.n439 B.n438 585
R276 B.n437 B.n436 585
R277 B.n435 B.n434 585
R278 B.n433 B.n432 585
R279 B.n431 B.n430 585
R280 B.n429 B.n428 585
R281 B.n427 B.n426 585
R282 B.n425 B.n424 585
R283 B.n423 B.n422 585
R284 B.n421 B.n420 585
R285 B.n419 B.n418 585
R286 B.n417 B.n416 585
R287 B.n415 B.n414 585
R288 B.n413 B.n412 585
R289 B.n411 B.n410 585
R290 B.n409 B.n408 585
R291 B.n407 B.n406 585
R292 B.n405 B.n404 585
R293 B.n403 B.n402 585
R294 B.n401 B.n400 585
R295 B.n399 B.n398 585
R296 B.n397 B.n396 585
R297 B.n395 B.n394 585
R298 B.n393 B.n392 585
R299 B.n391 B.n390 585
R300 B.n389 B.n388 585
R301 B.n387 B.n386 585
R302 B.n385 B.n384 585
R303 B.n383 B.n382 585
R304 B.n338 B.n337 585
R305 B.n535 B.n534 585
R306 B.n334 B.n333 585
R307 B.n335 B.n334 585
R308 B.n541 B.n540 585
R309 B.n540 B.n539 585
R310 B.n542 B.n332 585
R311 B.n332 B.n331 585
R312 B.n544 B.n543 585
R313 B.n545 B.n544 585
R314 B.n326 B.n325 585
R315 B.n327 B.n326 585
R316 B.n553 B.n552 585
R317 B.n552 B.n551 585
R318 B.n554 B.n324 585
R319 B.n324 B.n323 585
R320 B.n556 B.n555 585
R321 B.n557 B.n556 585
R322 B.n318 B.n317 585
R323 B.n319 B.n318 585
R324 B.n565 B.n564 585
R325 B.n564 B.n563 585
R326 B.n566 B.n316 585
R327 B.n316 B.n315 585
R328 B.n568 B.n567 585
R329 B.n569 B.n568 585
R330 B.n310 B.n309 585
R331 B.n311 B.n310 585
R332 B.n577 B.n576 585
R333 B.n576 B.n575 585
R334 B.n578 B.n308 585
R335 B.n308 B.n307 585
R336 B.n580 B.n579 585
R337 B.n581 B.n580 585
R338 B.n302 B.n301 585
R339 B.n303 B.n302 585
R340 B.n590 B.n589 585
R341 B.n589 B.n588 585
R342 B.n591 B.n300 585
R343 B.n587 B.n300 585
R344 B.n593 B.n592 585
R345 B.n594 B.n593 585
R346 B.n295 B.n294 585
R347 B.n296 B.n295 585
R348 B.n602 B.n601 585
R349 B.n601 B.n600 585
R350 B.n603 B.n293 585
R351 B.n293 B.n292 585
R352 B.n605 B.n604 585
R353 B.n606 B.n605 585
R354 B.n287 B.n286 585
R355 B.n288 B.n287 585
R356 B.n614 B.n613 585
R357 B.n613 B.n612 585
R358 B.n615 B.n285 585
R359 B.n285 B.n283 585
R360 B.n617 B.n616 585
R361 B.n618 B.n617 585
R362 B.n279 B.n278 585
R363 B.n284 B.n279 585
R364 B.n626 B.n625 585
R365 B.n625 B.n624 585
R366 B.n627 B.n277 585
R367 B.n277 B.n276 585
R368 B.n629 B.n628 585
R369 B.n630 B.n629 585
R370 B.n271 B.n270 585
R371 B.n272 B.n271 585
R372 B.n638 B.n637 585
R373 B.n637 B.t2 585
R374 B.n639 B.n269 585
R375 B.n269 B.n268 585
R376 B.n641 B.n640 585
R377 B.n642 B.n641 585
R378 B.n2 B.n0 585
R379 B.n4 B.n2 585
R380 B.n3 B.n1 585
R381 B.n767 B.n3 585
R382 B.n765 B.n764 585
R383 B.n766 B.n765 585
R384 B.n763 B.n9 585
R385 B.n9 B.n8 585
R386 B.n762 B.n761 585
R387 B.n761 B.t4 585
R388 B.n11 B.n10 585
R389 B.n760 B.n11 585
R390 B.n758 B.n757 585
R391 B.n759 B.n758 585
R392 B.n756 B.n16 585
R393 B.n16 B.n15 585
R394 B.n755 B.n754 585
R395 B.n754 B.n753 585
R396 B.n18 B.n17 585
R397 B.n752 B.n18 585
R398 B.n750 B.n749 585
R399 B.n751 B.n750 585
R400 B.n748 B.n23 585
R401 B.n23 B.n22 585
R402 B.n747 B.n746 585
R403 B.n746 B.n745 585
R404 B.n25 B.n24 585
R405 B.n744 B.n25 585
R406 B.n742 B.n741 585
R407 B.n743 B.n742 585
R408 B.n740 B.n30 585
R409 B.n30 B.n29 585
R410 B.n739 B.n738 585
R411 B.n738 B.n737 585
R412 B.n32 B.n31 585
R413 B.n736 B.n32 585
R414 B.n734 B.n733 585
R415 B.n735 B.n734 585
R416 B.n732 B.n36 585
R417 B.n39 B.n36 585
R418 B.n731 B.n730 585
R419 B.n730 B.n729 585
R420 B.n38 B.n37 585
R421 B.n728 B.n38 585
R422 B.n726 B.n725 585
R423 B.n727 B.n726 585
R424 B.n724 B.n44 585
R425 B.n44 B.n43 585
R426 B.n723 B.n722 585
R427 B.n722 B.n721 585
R428 B.n46 B.n45 585
R429 B.n720 B.n46 585
R430 B.n718 B.n717 585
R431 B.n719 B.n718 585
R432 B.n716 B.n51 585
R433 B.n51 B.n50 585
R434 B.n715 B.n714 585
R435 B.n714 B.n713 585
R436 B.n53 B.n52 585
R437 B.n712 B.n53 585
R438 B.n710 B.n709 585
R439 B.n711 B.n710 585
R440 B.n708 B.n58 585
R441 B.n58 B.n57 585
R442 B.n707 B.n706 585
R443 B.n706 B.n705 585
R444 B.n60 B.n59 585
R445 B.n704 B.n60 585
R446 B.n702 B.n701 585
R447 B.n703 B.n702 585
R448 B.n700 B.n65 585
R449 B.n65 B.n64 585
R450 B.n699 B.n698 585
R451 B.n698 B.n697 585
R452 B.n67 B.n66 585
R453 B.n696 B.n67 585
R454 B.n770 B.n769 585
R455 B.n769 B.n768 585
R456 B.n530 B.n334 478.086
R457 B.n114 B.n67 478.086
R458 B.n534 B.n336 478.086
R459 B.n694 B.n69 478.086
R460 B.n379 B.t10 377.202
R461 B.n377 B.t14 377.202
R462 B.n111 B.t17 377.202
R463 B.n109 B.t21 377.202
R464 B.n379 B.t13 267.353
R465 B.n109 B.t22 267.353
R466 B.n377 B.t16 267.353
R467 B.n111 B.t19 267.353
R468 B.n695 B.n107 256.663
R469 B.n695 B.n106 256.663
R470 B.n695 B.n105 256.663
R471 B.n695 B.n104 256.663
R472 B.n695 B.n103 256.663
R473 B.n695 B.n102 256.663
R474 B.n695 B.n101 256.663
R475 B.n695 B.n100 256.663
R476 B.n695 B.n99 256.663
R477 B.n695 B.n98 256.663
R478 B.n695 B.n97 256.663
R479 B.n695 B.n96 256.663
R480 B.n695 B.n95 256.663
R481 B.n695 B.n94 256.663
R482 B.n695 B.n93 256.663
R483 B.n695 B.n92 256.663
R484 B.n695 B.n91 256.663
R485 B.n695 B.n90 256.663
R486 B.n695 B.n89 256.663
R487 B.n695 B.n88 256.663
R488 B.n695 B.n87 256.663
R489 B.n695 B.n86 256.663
R490 B.n695 B.n85 256.663
R491 B.n695 B.n84 256.663
R492 B.n695 B.n83 256.663
R493 B.n695 B.n82 256.663
R494 B.n695 B.n81 256.663
R495 B.n695 B.n80 256.663
R496 B.n695 B.n79 256.663
R497 B.n695 B.n78 256.663
R498 B.n695 B.n77 256.663
R499 B.n695 B.n76 256.663
R500 B.n695 B.n75 256.663
R501 B.n695 B.n74 256.663
R502 B.n695 B.n73 256.663
R503 B.n695 B.n72 256.663
R504 B.n695 B.n71 256.663
R505 B.n695 B.n70 256.663
R506 B.n532 B.n531 256.663
R507 B.n532 B.n339 256.663
R508 B.n532 B.n340 256.663
R509 B.n532 B.n341 256.663
R510 B.n532 B.n342 256.663
R511 B.n532 B.n343 256.663
R512 B.n532 B.n344 256.663
R513 B.n532 B.n345 256.663
R514 B.n532 B.n346 256.663
R515 B.n532 B.n347 256.663
R516 B.n532 B.n348 256.663
R517 B.n532 B.n349 256.663
R518 B.n532 B.n350 256.663
R519 B.n532 B.n351 256.663
R520 B.n532 B.n352 256.663
R521 B.n532 B.n353 256.663
R522 B.n532 B.n354 256.663
R523 B.n532 B.n355 256.663
R524 B.n532 B.n356 256.663
R525 B.n532 B.n357 256.663
R526 B.n532 B.n358 256.663
R527 B.n532 B.n359 256.663
R528 B.n532 B.n360 256.663
R529 B.n532 B.n361 256.663
R530 B.n532 B.n362 256.663
R531 B.n532 B.n363 256.663
R532 B.n532 B.n364 256.663
R533 B.n532 B.n365 256.663
R534 B.n532 B.n366 256.663
R535 B.n532 B.n367 256.663
R536 B.n532 B.n368 256.663
R537 B.n532 B.n369 256.663
R538 B.n532 B.n370 256.663
R539 B.n532 B.n371 256.663
R540 B.n532 B.n372 256.663
R541 B.n532 B.n373 256.663
R542 B.n532 B.n374 256.663
R543 B.n533 B.n532 256.663
R544 B.n380 B.t12 235.742
R545 B.n110 B.t23 235.742
R546 B.n378 B.t15 235.742
R547 B.n112 B.t20 235.742
R548 B.n540 B.n334 163.367
R549 B.n540 B.n332 163.367
R550 B.n544 B.n332 163.367
R551 B.n544 B.n326 163.367
R552 B.n552 B.n326 163.367
R553 B.n552 B.n324 163.367
R554 B.n556 B.n324 163.367
R555 B.n556 B.n318 163.367
R556 B.n564 B.n318 163.367
R557 B.n564 B.n316 163.367
R558 B.n568 B.n316 163.367
R559 B.n568 B.n310 163.367
R560 B.n576 B.n310 163.367
R561 B.n576 B.n308 163.367
R562 B.n580 B.n308 163.367
R563 B.n580 B.n302 163.367
R564 B.n589 B.n302 163.367
R565 B.n589 B.n300 163.367
R566 B.n593 B.n300 163.367
R567 B.n593 B.n295 163.367
R568 B.n601 B.n295 163.367
R569 B.n601 B.n293 163.367
R570 B.n605 B.n293 163.367
R571 B.n605 B.n287 163.367
R572 B.n613 B.n287 163.367
R573 B.n613 B.n285 163.367
R574 B.n617 B.n285 163.367
R575 B.n617 B.n279 163.367
R576 B.n625 B.n279 163.367
R577 B.n625 B.n277 163.367
R578 B.n629 B.n277 163.367
R579 B.n629 B.n271 163.367
R580 B.n637 B.n271 163.367
R581 B.n637 B.n269 163.367
R582 B.n641 B.n269 163.367
R583 B.n641 B.n2 163.367
R584 B.n769 B.n2 163.367
R585 B.n769 B.n3 163.367
R586 B.n765 B.n3 163.367
R587 B.n765 B.n9 163.367
R588 B.n761 B.n9 163.367
R589 B.n761 B.n11 163.367
R590 B.n758 B.n11 163.367
R591 B.n758 B.n16 163.367
R592 B.n754 B.n16 163.367
R593 B.n754 B.n18 163.367
R594 B.n750 B.n18 163.367
R595 B.n750 B.n23 163.367
R596 B.n746 B.n23 163.367
R597 B.n746 B.n25 163.367
R598 B.n742 B.n25 163.367
R599 B.n742 B.n30 163.367
R600 B.n738 B.n30 163.367
R601 B.n738 B.n32 163.367
R602 B.n734 B.n32 163.367
R603 B.n734 B.n36 163.367
R604 B.n730 B.n36 163.367
R605 B.n730 B.n38 163.367
R606 B.n726 B.n38 163.367
R607 B.n726 B.n44 163.367
R608 B.n722 B.n44 163.367
R609 B.n722 B.n46 163.367
R610 B.n718 B.n46 163.367
R611 B.n718 B.n51 163.367
R612 B.n714 B.n51 163.367
R613 B.n714 B.n53 163.367
R614 B.n710 B.n53 163.367
R615 B.n710 B.n58 163.367
R616 B.n706 B.n58 163.367
R617 B.n706 B.n60 163.367
R618 B.n702 B.n60 163.367
R619 B.n702 B.n65 163.367
R620 B.n698 B.n65 163.367
R621 B.n698 B.n67 163.367
R622 B.n376 B.n375 163.367
R623 B.n525 B.n375 163.367
R624 B.n523 B.n522 163.367
R625 B.n519 B.n518 163.367
R626 B.n515 B.n514 163.367
R627 B.n511 B.n510 163.367
R628 B.n507 B.n506 163.367
R629 B.n503 B.n502 163.367
R630 B.n499 B.n498 163.367
R631 B.n495 B.n494 163.367
R632 B.n491 B.n490 163.367
R633 B.n487 B.n486 163.367
R634 B.n483 B.n482 163.367
R635 B.n479 B.n478 163.367
R636 B.n475 B.n474 163.367
R637 B.n471 B.n470 163.367
R638 B.n467 B.n466 163.367
R639 B.n462 B.n461 163.367
R640 B.n458 B.n457 163.367
R641 B.n454 B.n453 163.367
R642 B.n450 B.n449 163.367
R643 B.n446 B.n445 163.367
R644 B.n442 B.n441 163.367
R645 B.n438 B.n437 163.367
R646 B.n434 B.n433 163.367
R647 B.n430 B.n429 163.367
R648 B.n426 B.n425 163.367
R649 B.n422 B.n421 163.367
R650 B.n418 B.n417 163.367
R651 B.n414 B.n413 163.367
R652 B.n410 B.n409 163.367
R653 B.n406 B.n405 163.367
R654 B.n402 B.n401 163.367
R655 B.n398 B.n397 163.367
R656 B.n394 B.n393 163.367
R657 B.n390 B.n389 163.367
R658 B.n386 B.n385 163.367
R659 B.n382 B.n338 163.367
R660 B.n538 B.n336 163.367
R661 B.n538 B.n330 163.367
R662 B.n546 B.n330 163.367
R663 B.n546 B.n328 163.367
R664 B.n550 B.n328 163.367
R665 B.n550 B.n322 163.367
R666 B.n558 B.n322 163.367
R667 B.n558 B.n320 163.367
R668 B.n562 B.n320 163.367
R669 B.n562 B.n314 163.367
R670 B.n570 B.n314 163.367
R671 B.n570 B.n312 163.367
R672 B.n574 B.n312 163.367
R673 B.n574 B.n306 163.367
R674 B.n582 B.n306 163.367
R675 B.n582 B.n304 163.367
R676 B.n586 B.n304 163.367
R677 B.n586 B.n299 163.367
R678 B.n595 B.n299 163.367
R679 B.n595 B.n297 163.367
R680 B.n599 B.n297 163.367
R681 B.n599 B.n291 163.367
R682 B.n607 B.n291 163.367
R683 B.n607 B.n289 163.367
R684 B.n611 B.n289 163.367
R685 B.n611 B.n282 163.367
R686 B.n619 B.n282 163.367
R687 B.n619 B.n280 163.367
R688 B.n623 B.n280 163.367
R689 B.n623 B.n275 163.367
R690 B.n631 B.n275 163.367
R691 B.n631 B.n273 163.367
R692 B.n636 B.n273 163.367
R693 B.n636 B.n267 163.367
R694 B.n643 B.n267 163.367
R695 B.n644 B.n643 163.367
R696 B.n644 B.n5 163.367
R697 B.n6 B.n5 163.367
R698 B.n7 B.n6 163.367
R699 B.n649 B.n7 163.367
R700 B.n649 B.n12 163.367
R701 B.n13 B.n12 163.367
R702 B.n14 B.n13 163.367
R703 B.n654 B.n14 163.367
R704 B.n654 B.n19 163.367
R705 B.n20 B.n19 163.367
R706 B.n21 B.n20 163.367
R707 B.n659 B.n21 163.367
R708 B.n659 B.n26 163.367
R709 B.n27 B.n26 163.367
R710 B.n28 B.n27 163.367
R711 B.n664 B.n28 163.367
R712 B.n664 B.n33 163.367
R713 B.n34 B.n33 163.367
R714 B.n35 B.n34 163.367
R715 B.n669 B.n35 163.367
R716 B.n669 B.n40 163.367
R717 B.n41 B.n40 163.367
R718 B.n42 B.n41 163.367
R719 B.n674 B.n42 163.367
R720 B.n674 B.n47 163.367
R721 B.n48 B.n47 163.367
R722 B.n49 B.n48 163.367
R723 B.n679 B.n49 163.367
R724 B.n679 B.n54 163.367
R725 B.n55 B.n54 163.367
R726 B.n56 B.n55 163.367
R727 B.n684 B.n56 163.367
R728 B.n684 B.n61 163.367
R729 B.n62 B.n61 163.367
R730 B.n63 B.n62 163.367
R731 B.n689 B.n63 163.367
R732 B.n689 B.n68 163.367
R733 B.n69 B.n68 163.367
R734 B.n118 B.n117 163.367
R735 B.n122 B.n121 163.367
R736 B.n126 B.n125 163.367
R737 B.n130 B.n129 163.367
R738 B.n134 B.n133 163.367
R739 B.n138 B.n137 163.367
R740 B.n142 B.n141 163.367
R741 B.n146 B.n145 163.367
R742 B.n150 B.n149 163.367
R743 B.n154 B.n153 163.367
R744 B.n158 B.n157 163.367
R745 B.n162 B.n161 163.367
R746 B.n166 B.n165 163.367
R747 B.n170 B.n169 163.367
R748 B.n174 B.n173 163.367
R749 B.n178 B.n177 163.367
R750 B.n182 B.n181 163.367
R751 B.n186 B.n185 163.367
R752 B.n190 B.n189 163.367
R753 B.n194 B.n193 163.367
R754 B.n198 B.n197 163.367
R755 B.n203 B.n202 163.367
R756 B.n207 B.n206 163.367
R757 B.n211 B.n210 163.367
R758 B.n215 B.n214 163.367
R759 B.n219 B.n218 163.367
R760 B.n223 B.n222 163.367
R761 B.n227 B.n226 163.367
R762 B.n231 B.n230 163.367
R763 B.n235 B.n234 163.367
R764 B.n239 B.n238 163.367
R765 B.n243 B.n242 163.367
R766 B.n247 B.n246 163.367
R767 B.n251 B.n250 163.367
R768 B.n255 B.n254 163.367
R769 B.n259 B.n258 163.367
R770 B.n263 B.n262 163.367
R771 B.n694 B.n108 163.367
R772 B.n532 B.n335 86.7334
R773 B.n696 B.n695 86.7334
R774 B.n531 B.n530 71.676
R775 B.n525 B.n339 71.676
R776 B.n522 B.n340 71.676
R777 B.n518 B.n341 71.676
R778 B.n514 B.n342 71.676
R779 B.n510 B.n343 71.676
R780 B.n506 B.n344 71.676
R781 B.n502 B.n345 71.676
R782 B.n498 B.n346 71.676
R783 B.n494 B.n347 71.676
R784 B.n490 B.n348 71.676
R785 B.n486 B.n349 71.676
R786 B.n482 B.n350 71.676
R787 B.n478 B.n351 71.676
R788 B.n474 B.n352 71.676
R789 B.n470 B.n353 71.676
R790 B.n466 B.n354 71.676
R791 B.n461 B.n355 71.676
R792 B.n457 B.n356 71.676
R793 B.n453 B.n357 71.676
R794 B.n449 B.n358 71.676
R795 B.n445 B.n359 71.676
R796 B.n441 B.n360 71.676
R797 B.n437 B.n361 71.676
R798 B.n433 B.n362 71.676
R799 B.n429 B.n363 71.676
R800 B.n425 B.n364 71.676
R801 B.n421 B.n365 71.676
R802 B.n417 B.n366 71.676
R803 B.n413 B.n367 71.676
R804 B.n409 B.n368 71.676
R805 B.n405 B.n369 71.676
R806 B.n401 B.n370 71.676
R807 B.n397 B.n371 71.676
R808 B.n393 B.n372 71.676
R809 B.n389 B.n373 71.676
R810 B.n385 B.n374 71.676
R811 B.n533 B.n338 71.676
R812 B.n114 B.n70 71.676
R813 B.n118 B.n71 71.676
R814 B.n122 B.n72 71.676
R815 B.n126 B.n73 71.676
R816 B.n130 B.n74 71.676
R817 B.n134 B.n75 71.676
R818 B.n138 B.n76 71.676
R819 B.n142 B.n77 71.676
R820 B.n146 B.n78 71.676
R821 B.n150 B.n79 71.676
R822 B.n154 B.n80 71.676
R823 B.n158 B.n81 71.676
R824 B.n162 B.n82 71.676
R825 B.n166 B.n83 71.676
R826 B.n170 B.n84 71.676
R827 B.n174 B.n85 71.676
R828 B.n178 B.n86 71.676
R829 B.n182 B.n87 71.676
R830 B.n186 B.n88 71.676
R831 B.n190 B.n89 71.676
R832 B.n194 B.n90 71.676
R833 B.n198 B.n91 71.676
R834 B.n203 B.n92 71.676
R835 B.n207 B.n93 71.676
R836 B.n211 B.n94 71.676
R837 B.n215 B.n95 71.676
R838 B.n219 B.n96 71.676
R839 B.n223 B.n97 71.676
R840 B.n227 B.n98 71.676
R841 B.n231 B.n99 71.676
R842 B.n235 B.n100 71.676
R843 B.n239 B.n101 71.676
R844 B.n243 B.n102 71.676
R845 B.n247 B.n103 71.676
R846 B.n251 B.n104 71.676
R847 B.n255 B.n105 71.676
R848 B.n259 B.n106 71.676
R849 B.n263 B.n107 71.676
R850 B.n108 B.n107 71.676
R851 B.n262 B.n106 71.676
R852 B.n258 B.n105 71.676
R853 B.n254 B.n104 71.676
R854 B.n250 B.n103 71.676
R855 B.n246 B.n102 71.676
R856 B.n242 B.n101 71.676
R857 B.n238 B.n100 71.676
R858 B.n234 B.n99 71.676
R859 B.n230 B.n98 71.676
R860 B.n226 B.n97 71.676
R861 B.n222 B.n96 71.676
R862 B.n218 B.n95 71.676
R863 B.n214 B.n94 71.676
R864 B.n210 B.n93 71.676
R865 B.n206 B.n92 71.676
R866 B.n202 B.n91 71.676
R867 B.n197 B.n90 71.676
R868 B.n193 B.n89 71.676
R869 B.n189 B.n88 71.676
R870 B.n185 B.n87 71.676
R871 B.n181 B.n86 71.676
R872 B.n177 B.n85 71.676
R873 B.n173 B.n84 71.676
R874 B.n169 B.n83 71.676
R875 B.n165 B.n82 71.676
R876 B.n161 B.n81 71.676
R877 B.n157 B.n80 71.676
R878 B.n153 B.n79 71.676
R879 B.n149 B.n78 71.676
R880 B.n145 B.n77 71.676
R881 B.n141 B.n76 71.676
R882 B.n137 B.n75 71.676
R883 B.n133 B.n74 71.676
R884 B.n129 B.n73 71.676
R885 B.n125 B.n72 71.676
R886 B.n121 B.n71 71.676
R887 B.n117 B.n70 71.676
R888 B.n531 B.n376 71.676
R889 B.n523 B.n339 71.676
R890 B.n519 B.n340 71.676
R891 B.n515 B.n341 71.676
R892 B.n511 B.n342 71.676
R893 B.n507 B.n343 71.676
R894 B.n503 B.n344 71.676
R895 B.n499 B.n345 71.676
R896 B.n495 B.n346 71.676
R897 B.n491 B.n347 71.676
R898 B.n487 B.n348 71.676
R899 B.n483 B.n349 71.676
R900 B.n479 B.n350 71.676
R901 B.n475 B.n351 71.676
R902 B.n471 B.n352 71.676
R903 B.n467 B.n353 71.676
R904 B.n462 B.n354 71.676
R905 B.n458 B.n355 71.676
R906 B.n454 B.n356 71.676
R907 B.n450 B.n357 71.676
R908 B.n446 B.n358 71.676
R909 B.n442 B.n359 71.676
R910 B.n438 B.n360 71.676
R911 B.n434 B.n361 71.676
R912 B.n430 B.n362 71.676
R913 B.n426 B.n363 71.676
R914 B.n422 B.n364 71.676
R915 B.n418 B.n365 71.676
R916 B.n414 B.n366 71.676
R917 B.n410 B.n367 71.676
R918 B.n406 B.n368 71.676
R919 B.n402 B.n369 71.676
R920 B.n398 B.n370 71.676
R921 B.n394 B.n371 71.676
R922 B.n390 B.n372 71.676
R923 B.n386 B.n373 71.676
R924 B.n382 B.n374 71.676
R925 B.n534 B.n533 71.676
R926 B.n381 B.n380 59.5399
R927 B.n464 B.n378 59.5399
R928 B.n113 B.n112 59.5399
R929 B.n200 B.n110 59.5399
R930 B.n539 B.n335 51.2861
R931 B.n539 B.n331 51.2861
R932 B.n545 B.n331 51.2861
R933 B.n545 B.n327 51.2861
R934 B.n551 B.n327 51.2861
R935 B.n557 B.n323 51.2861
R936 B.n557 B.n319 51.2861
R937 B.n563 B.n319 51.2861
R938 B.n563 B.n315 51.2861
R939 B.n569 B.n315 51.2861
R940 B.n569 B.n311 51.2861
R941 B.n575 B.n311 51.2861
R942 B.n581 B.n307 51.2861
R943 B.n581 B.n303 51.2861
R944 B.n588 B.n303 51.2861
R945 B.n588 B.n587 51.2861
R946 B.n594 B.n296 51.2861
R947 B.n600 B.n296 51.2861
R948 B.n600 B.n292 51.2861
R949 B.n606 B.n292 51.2861
R950 B.n612 B.n288 51.2861
R951 B.n612 B.n283 51.2861
R952 B.n618 B.n283 51.2861
R953 B.n618 B.n284 51.2861
R954 B.n624 B.n276 51.2861
R955 B.n630 B.n276 51.2861
R956 B.n630 B.n272 51.2861
R957 B.t2 B.n272 51.2861
R958 B.t2 B.n268 51.2861
R959 B.n642 B.n268 51.2861
R960 B.n642 B.n4 51.2861
R961 B.n768 B.n4 51.2861
R962 B.n768 B.n767 51.2861
R963 B.n767 B.n766 51.2861
R964 B.n766 B.n8 51.2861
R965 B.t4 B.n8 51.2861
R966 B.t4 B.n760 51.2861
R967 B.n760 B.n759 51.2861
R968 B.n759 B.n15 51.2861
R969 B.n753 B.n15 51.2861
R970 B.n752 B.n751 51.2861
R971 B.n751 B.n22 51.2861
R972 B.n745 B.n22 51.2861
R973 B.n745 B.n744 51.2861
R974 B.n743 B.n29 51.2861
R975 B.n737 B.n29 51.2861
R976 B.n737 B.n736 51.2861
R977 B.n736 B.n735 51.2861
R978 B.n729 B.n39 51.2861
R979 B.n729 B.n728 51.2861
R980 B.n728 B.n727 51.2861
R981 B.n727 B.n43 51.2861
R982 B.n721 B.n720 51.2861
R983 B.n720 B.n719 51.2861
R984 B.n719 B.n50 51.2861
R985 B.n713 B.n50 51.2861
R986 B.n713 B.n712 51.2861
R987 B.n712 B.n711 51.2861
R988 B.n711 B.n57 51.2861
R989 B.n705 B.n704 51.2861
R990 B.n704 B.n703 51.2861
R991 B.n703 B.n64 51.2861
R992 B.n697 B.n64 51.2861
R993 B.n697 B.n696 51.2861
R994 B.n551 B.t11 42.2357
R995 B.n575 B.t8 42.2357
R996 B.n721 B.t5 42.2357
R997 B.n705 B.t18 42.2357
R998 B.n624 B.t7 40.7273
R999 B.n753 B.t1 40.7273
R1000 B.n587 B.t0 31.6769
R1001 B.n39 B.t6 31.6769
R1002 B.n380 B.n379 31.6126
R1003 B.n378 B.n377 31.6126
R1004 B.n112 B.n111 31.6126
R1005 B.n110 B.n109 31.6126
R1006 B.n115 B.n66 31.0639
R1007 B.n693 B.n692 31.0639
R1008 B.n536 B.n535 31.0639
R1009 B.n529 B.n333 31.0639
R1010 B.t9 B.n288 30.1685
R1011 B.n744 B.t3 30.1685
R1012 B.n606 B.t9 21.1181
R1013 B.t3 B.n743 21.1181
R1014 B.n594 B.t0 19.6097
R1015 B.n735 B.t6 19.6097
R1016 B B.n770 18.0485
R1017 B.n116 B.n115 10.6151
R1018 B.n119 B.n116 10.6151
R1019 B.n120 B.n119 10.6151
R1020 B.n123 B.n120 10.6151
R1021 B.n124 B.n123 10.6151
R1022 B.n127 B.n124 10.6151
R1023 B.n128 B.n127 10.6151
R1024 B.n131 B.n128 10.6151
R1025 B.n132 B.n131 10.6151
R1026 B.n135 B.n132 10.6151
R1027 B.n136 B.n135 10.6151
R1028 B.n139 B.n136 10.6151
R1029 B.n140 B.n139 10.6151
R1030 B.n143 B.n140 10.6151
R1031 B.n144 B.n143 10.6151
R1032 B.n147 B.n144 10.6151
R1033 B.n148 B.n147 10.6151
R1034 B.n151 B.n148 10.6151
R1035 B.n152 B.n151 10.6151
R1036 B.n155 B.n152 10.6151
R1037 B.n156 B.n155 10.6151
R1038 B.n159 B.n156 10.6151
R1039 B.n160 B.n159 10.6151
R1040 B.n163 B.n160 10.6151
R1041 B.n164 B.n163 10.6151
R1042 B.n167 B.n164 10.6151
R1043 B.n168 B.n167 10.6151
R1044 B.n171 B.n168 10.6151
R1045 B.n172 B.n171 10.6151
R1046 B.n175 B.n172 10.6151
R1047 B.n176 B.n175 10.6151
R1048 B.n179 B.n176 10.6151
R1049 B.n180 B.n179 10.6151
R1050 B.n184 B.n183 10.6151
R1051 B.n187 B.n184 10.6151
R1052 B.n188 B.n187 10.6151
R1053 B.n191 B.n188 10.6151
R1054 B.n192 B.n191 10.6151
R1055 B.n195 B.n192 10.6151
R1056 B.n196 B.n195 10.6151
R1057 B.n199 B.n196 10.6151
R1058 B.n204 B.n201 10.6151
R1059 B.n205 B.n204 10.6151
R1060 B.n208 B.n205 10.6151
R1061 B.n209 B.n208 10.6151
R1062 B.n212 B.n209 10.6151
R1063 B.n213 B.n212 10.6151
R1064 B.n216 B.n213 10.6151
R1065 B.n217 B.n216 10.6151
R1066 B.n220 B.n217 10.6151
R1067 B.n221 B.n220 10.6151
R1068 B.n224 B.n221 10.6151
R1069 B.n225 B.n224 10.6151
R1070 B.n228 B.n225 10.6151
R1071 B.n229 B.n228 10.6151
R1072 B.n232 B.n229 10.6151
R1073 B.n233 B.n232 10.6151
R1074 B.n236 B.n233 10.6151
R1075 B.n237 B.n236 10.6151
R1076 B.n240 B.n237 10.6151
R1077 B.n241 B.n240 10.6151
R1078 B.n244 B.n241 10.6151
R1079 B.n245 B.n244 10.6151
R1080 B.n248 B.n245 10.6151
R1081 B.n249 B.n248 10.6151
R1082 B.n252 B.n249 10.6151
R1083 B.n253 B.n252 10.6151
R1084 B.n256 B.n253 10.6151
R1085 B.n257 B.n256 10.6151
R1086 B.n260 B.n257 10.6151
R1087 B.n261 B.n260 10.6151
R1088 B.n264 B.n261 10.6151
R1089 B.n265 B.n264 10.6151
R1090 B.n693 B.n265 10.6151
R1091 B.n537 B.n536 10.6151
R1092 B.n537 B.n329 10.6151
R1093 B.n547 B.n329 10.6151
R1094 B.n548 B.n547 10.6151
R1095 B.n549 B.n548 10.6151
R1096 B.n549 B.n321 10.6151
R1097 B.n559 B.n321 10.6151
R1098 B.n560 B.n559 10.6151
R1099 B.n561 B.n560 10.6151
R1100 B.n561 B.n313 10.6151
R1101 B.n571 B.n313 10.6151
R1102 B.n572 B.n571 10.6151
R1103 B.n573 B.n572 10.6151
R1104 B.n573 B.n305 10.6151
R1105 B.n583 B.n305 10.6151
R1106 B.n584 B.n583 10.6151
R1107 B.n585 B.n584 10.6151
R1108 B.n585 B.n298 10.6151
R1109 B.n596 B.n298 10.6151
R1110 B.n597 B.n596 10.6151
R1111 B.n598 B.n597 10.6151
R1112 B.n598 B.n290 10.6151
R1113 B.n608 B.n290 10.6151
R1114 B.n609 B.n608 10.6151
R1115 B.n610 B.n609 10.6151
R1116 B.n610 B.n281 10.6151
R1117 B.n620 B.n281 10.6151
R1118 B.n621 B.n620 10.6151
R1119 B.n622 B.n621 10.6151
R1120 B.n622 B.n274 10.6151
R1121 B.n632 B.n274 10.6151
R1122 B.n633 B.n632 10.6151
R1123 B.n635 B.n633 10.6151
R1124 B.n635 B.n634 10.6151
R1125 B.n634 B.n266 10.6151
R1126 B.n645 B.n266 10.6151
R1127 B.n646 B.n645 10.6151
R1128 B.n647 B.n646 10.6151
R1129 B.n648 B.n647 10.6151
R1130 B.n650 B.n648 10.6151
R1131 B.n651 B.n650 10.6151
R1132 B.n652 B.n651 10.6151
R1133 B.n653 B.n652 10.6151
R1134 B.n655 B.n653 10.6151
R1135 B.n656 B.n655 10.6151
R1136 B.n657 B.n656 10.6151
R1137 B.n658 B.n657 10.6151
R1138 B.n660 B.n658 10.6151
R1139 B.n661 B.n660 10.6151
R1140 B.n662 B.n661 10.6151
R1141 B.n663 B.n662 10.6151
R1142 B.n665 B.n663 10.6151
R1143 B.n666 B.n665 10.6151
R1144 B.n667 B.n666 10.6151
R1145 B.n668 B.n667 10.6151
R1146 B.n670 B.n668 10.6151
R1147 B.n671 B.n670 10.6151
R1148 B.n672 B.n671 10.6151
R1149 B.n673 B.n672 10.6151
R1150 B.n675 B.n673 10.6151
R1151 B.n676 B.n675 10.6151
R1152 B.n677 B.n676 10.6151
R1153 B.n678 B.n677 10.6151
R1154 B.n680 B.n678 10.6151
R1155 B.n681 B.n680 10.6151
R1156 B.n682 B.n681 10.6151
R1157 B.n683 B.n682 10.6151
R1158 B.n685 B.n683 10.6151
R1159 B.n686 B.n685 10.6151
R1160 B.n687 B.n686 10.6151
R1161 B.n688 B.n687 10.6151
R1162 B.n690 B.n688 10.6151
R1163 B.n691 B.n690 10.6151
R1164 B.n692 B.n691 10.6151
R1165 B.n529 B.n528 10.6151
R1166 B.n528 B.n527 10.6151
R1167 B.n527 B.n526 10.6151
R1168 B.n526 B.n524 10.6151
R1169 B.n524 B.n521 10.6151
R1170 B.n521 B.n520 10.6151
R1171 B.n520 B.n517 10.6151
R1172 B.n517 B.n516 10.6151
R1173 B.n516 B.n513 10.6151
R1174 B.n513 B.n512 10.6151
R1175 B.n512 B.n509 10.6151
R1176 B.n509 B.n508 10.6151
R1177 B.n508 B.n505 10.6151
R1178 B.n505 B.n504 10.6151
R1179 B.n504 B.n501 10.6151
R1180 B.n501 B.n500 10.6151
R1181 B.n500 B.n497 10.6151
R1182 B.n497 B.n496 10.6151
R1183 B.n496 B.n493 10.6151
R1184 B.n493 B.n492 10.6151
R1185 B.n492 B.n489 10.6151
R1186 B.n489 B.n488 10.6151
R1187 B.n488 B.n485 10.6151
R1188 B.n485 B.n484 10.6151
R1189 B.n484 B.n481 10.6151
R1190 B.n481 B.n480 10.6151
R1191 B.n480 B.n477 10.6151
R1192 B.n477 B.n476 10.6151
R1193 B.n476 B.n473 10.6151
R1194 B.n473 B.n472 10.6151
R1195 B.n472 B.n469 10.6151
R1196 B.n469 B.n468 10.6151
R1197 B.n468 B.n465 10.6151
R1198 B.n463 B.n460 10.6151
R1199 B.n460 B.n459 10.6151
R1200 B.n459 B.n456 10.6151
R1201 B.n456 B.n455 10.6151
R1202 B.n455 B.n452 10.6151
R1203 B.n452 B.n451 10.6151
R1204 B.n451 B.n448 10.6151
R1205 B.n448 B.n447 10.6151
R1206 B.n444 B.n443 10.6151
R1207 B.n443 B.n440 10.6151
R1208 B.n440 B.n439 10.6151
R1209 B.n439 B.n436 10.6151
R1210 B.n436 B.n435 10.6151
R1211 B.n435 B.n432 10.6151
R1212 B.n432 B.n431 10.6151
R1213 B.n431 B.n428 10.6151
R1214 B.n428 B.n427 10.6151
R1215 B.n427 B.n424 10.6151
R1216 B.n424 B.n423 10.6151
R1217 B.n423 B.n420 10.6151
R1218 B.n420 B.n419 10.6151
R1219 B.n419 B.n416 10.6151
R1220 B.n416 B.n415 10.6151
R1221 B.n415 B.n412 10.6151
R1222 B.n412 B.n411 10.6151
R1223 B.n411 B.n408 10.6151
R1224 B.n408 B.n407 10.6151
R1225 B.n407 B.n404 10.6151
R1226 B.n404 B.n403 10.6151
R1227 B.n403 B.n400 10.6151
R1228 B.n400 B.n399 10.6151
R1229 B.n399 B.n396 10.6151
R1230 B.n396 B.n395 10.6151
R1231 B.n395 B.n392 10.6151
R1232 B.n392 B.n391 10.6151
R1233 B.n391 B.n388 10.6151
R1234 B.n388 B.n387 10.6151
R1235 B.n387 B.n384 10.6151
R1236 B.n384 B.n383 10.6151
R1237 B.n383 B.n337 10.6151
R1238 B.n535 B.n337 10.6151
R1239 B.n541 B.n333 10.6151
R1240 B.n542 B.n541 10.6151
R1241 B.n543 B.n542 10.6151
R1242 B.n543 B.n325 10.6151
R1243 B.n553 B.n325 10.6151
R1244 B.n554 B.n553 10.6151
R1245 B.n555 B.n554 10.6151
R1246 B.n555 B.n317 10.6151
R1247 B.n565 B.n317 10.6151
R1248 B.n566 B.n565 10.6151
R1249 B.n567 B.n566 10.6151
R1250 B.n567 B.n309 10.6151
R1251 B.n577 B.n309 10.6151
R1252 B.n578 B.n577 10.6151
R1253 B.n579 B.n578 10.6151
R1254 B.n579 B.n301 10.6151
R1255 B.n590 B.n301 10.6151
R1256 B.n591 B.n590 10.6151
R1257 B.n592 B.n591 10.6151
R1258 B.n592 B.n294 10.6151
R1259 B.n602 B.n294 10.6151
R1260 B.n603 B.n602 10.6151
R1261 B.n604 B.n603 10.6151
R1262 B.n604 B.n286 10.6151
R1263 B.n614 B.n286 10.6151
R1264 B.n615 B.n614 10.6151
R1265 B.n616 B.n615 10.6151
R1266 B.n616 B.n278 10.6151
R1267 B.n626 B.n278 10.6151
R1268 B.n627 B.n626 10.6151
R1269 B.n628 B.n627 10.6151
R1270 B.n628 B.n270 10.6151
R1271 B.n638 B.n270 10.6151
R1272 B.n639 B.n638 10.6151
R1273 B.n640 B.n639 10.6151
R1274 B.n640 B.n0 10.6151
R1275 B.n764 B.n1 10.6151
R1276 B.n764 B.n763 10.6151
R1277 B.n763 B.n762 10.6151
R1278 B.n762 B.n10 10.6151
R1279 B.n757 B.n10 10.6151
R1280 B.n757 B.n756 10.6151
R1281 B.n756 B.n755 10.6151
R1282 B.n755 B.n17 10.6151
R1283 B.n749 B.n17 10.6151
R1284 B.n749 B.n748 10.6151
R1285 B.n748 B.n747 10.6151
R1286 B.n747 B.n24 10.6151
R1287 B.n741 B.n24 10.6151
R1288 B.n741 B.n740 10.6151
R1289 B.n740 B.n739 10.6151
R1290 B.n739 B.n31 10.6151
R1291 B.n733 B.n31 10.6151
R1292 B.n733 B.n732 10.6151
R1293 B.n732 B.n731 10.6151
R1294 B.n731 B.n37 10.6151
R1295 B.n725 B.n37 10.6151
R1296 B.n725 B.n724 10.6151
R1297 B.n724 B.n723 10.6151
R1298 B.n723 B.n45 10.6151
R1299 B.n717 B.n45 10.6151
R1300 B.n717 B.n716 10.6151
R1301 B.n716 B.n715 10.6151
R1302 B.n715 B.n52 10.6151
R1303 B.n709 B.n52 10.6151
R1304 B.n709 B.n708 10.6151
R1305 B.n708 B.n707 10.6151
R1306 B.n707 B.n59 10.6151
R1307 B.n701 B.n59 10.6151
R1308 B.n701 B.n700 10.6151
R1309 B.n700 B.n699 10.6151
R1310 B.n699 B.n66 10.6151
R1311 B.n284 B.t7 10.5593
R1312 B.t1 B.n752 10.5593
R1313 B.t11 B.n323 9.05089
R1314 B.t8 B.n307 9.05089
R1315 B.t5 B.n43 9.05089
R1316 B.t18 B.n57 9.05089
R1317 B.n183 B.n113 6.5566
R1318 B.n200 B.n199 6.5566
R1319 B.n464 B.n463 6.5566
R1320 B.n447 B.n381 6.5566
R1321 B.n180 B.n113 4.05904
R1322 B.n201 B.n200 4.05904
R1323 B.n465 B.n464 4.05904
R1324 B.n444 B.n381 4.05904
R1325 B.n770 B.n0 2.81026
R1326 B.n770 B.n1 2.81026
R1327 VP.n14 VP.t5 202.195
R1328 VP.n33 VP.n7 173.044
R1329 VP.n56 VP.n55 173.044
R1330 VP.n32 VP.n31 173.044
R1331 VP.n3 VP.t9 172.594
R1332 VP.n7 VP.t6 172.594
R1333 VP.n5 VP.t1 172.594
R1334 VP.n48 VP.t7 172.594
R1335 VP.n55 VP.t2 172.594
R1336 VP.n11 VP.t8 172.594
R1337 VP.n31 VP.t3 172.594
R1338 VP.n24 VP.t4 172.594
R1339 VP.n13 VP.t0 172.594
R1340 VP.n16 VP.n15 161.3
R1341 VP.n17 VP.n12 161.3
R1342 VP.n19 VP.n18 161.3
R1343 VP.n20 VP.n11 161.3
R1344 VP.n22 VP.n21 161.3
R1345 VP.n23 VP.n10 161.3
R1346 VP.n26 VP.n25 161.3
R1347 VP.n27 VP.n9 161.3
R1348 VP.n29 VP.n28 161.3
R1349 VP.n30 VP.n8 161.3
R1350 VP.n54 VP.n0 161.3
R1351 VP.n53 VP.n52 161.3
R1352 VP.n51 VP.n1 161.3
R1353 VP.n50 VP.n49 161.3
R1354 VP.n47 VP.n2 161.3
R1355 VP.n46 VP.n45 161.3
R1356 VP.n44 VP.n3 161.3
R1357 VP.n43 VP.n42 161.3
R1358 VP.n41 VP.n4 161.3
R1359 VP.n40 VP.n39 161.3
R1360 VP.n38 VP.n37 161.3
R1361 VP.n36 VP.n6 161.3
R1362 VP.n35 VP.n34 161.3
R1363 VP.n14 VP.n13 58.4685
R1364 VP.n42 VP.n41 56.5193
R1365 VP.n47 VP.n46 56.5193
R1366 VP.n23 VP.n22 56.5193
R1367 VP.n18 VP.n17 56.5193
R1368 VP.n37 VP.n36 45.8354
R1369 VP.n53 VP.n1 45.8354
R1370 VP.n29 VP.n9 45.8354
R1371 VP.n33 VP.n32 43.9285
R1372 VP.n36 VP.n35 35.1514
R1373 VP.n54 VP.n53 35.1514
R1374 VP.n30 VP.n29 35.1514
R1375 VP.n15 VP.n14 27.0985
R1376 VP.n41 VP.n40 24.4675
R1377 VP.n42 VP.n3 24.4675
R1378 VP.n46 VP.n3 24.4675
R1379 VP.n49 VP.n47 24.4675
R1380 VP.n25 VP.n23 24.4675
R1381 VP.n18 VP.n11 24.4675
R1382 VP.n22 VP.n11 24.4675
R1383 VP.n17 VP.n16 24.4675
R1384 VP.n37 VP.n5 18.1061
R1385 VP.n48 VP.n1 18.1061
R1386 VP.n24 VP.n9 18.1061
R1387 VP.n35 VP.n7 12.7233
R1388 VP.n55 VP.n54 12.7233
R1389 VP.n31 VP.n30 12.7233
R1390 VP.n40 VP.n5 6.36192
R1391 VP.n49 VP.n48 6.36192
R1392 VP.n25 VP.n24 6.36192
R1393 VP.n16 VP.n13 6.36192
R1394 VP.n15 VP.n12 0.189894
R1395 VP.n19 VP.n12 0.189894
R1396 VP.n20 VP.n19 0.189894
R1397 VP.n21 VP.n20 0.189894
R1398 VP.n21 VP.n10 0.189894
R1399 VP.n26 VP.n10 0.189894
R1400 VP.n27 VP.n26 0.189894
R1401 VP.n28 VP.n27 0.189894
R1402 VP.n28 VP.n8 0.189894
R1403 VP.n32 VP.n8 0.189894
R1404 VP.n34 VP.n33 0.189894
R1405 VP.n34 VP.n6 0.189894
R1406 VP.n38 VP.n6 0.189894
R1407 VP.n39 VP.n38 0.189894
R1408 VP.n39 VP.n4 0.189894
R1409 VP.n43 VP.n4 0.189894
R1410 VP.n44 VP.n43 0.189894
R1411 VP.n45 VP.n44 0.189894
R1412 VP.n45 VP.n2 0.189894
R1413 VP.n50 VP.n2 0.189894
R1414 VP.n51 VP.n50 0.189894
R1415 VP.n52 VP.n51 0.189894
R1416 VP.n52 VP.n0 0.189894
R1417 VP.n56 VP.n0 0.189894
R1418 VP VP.n56 0.0516364
R1419 VDD1.n44 VDD1.n0 289.615
R1420 VDD1.n95 VDD1.n51 289.615
R1421 VDD1.n45 VDD1.n44 185
R1422 VDD1.n43 VDD1.n42 185
R1423 VDD1.n4 VDD1.n3 185
R1424 VDD1.n8 VDD1.n6 185
R1425 VDD1.n37 VDD1.n36 185
R1426 VDD1.n35 VDD1.n34 185
R1427 VDD1.n10 VDD1.n9 185
R1428 VDD1.n29 VDD1.n28 185
R1429 VDD1.n27 VDD1.n26 185
R1430 VDD1.n14 VDD1.n13 185
R1431 VDD1.n21 VDD1.n20 185
R1432 VDD1.n19 VDD1.n18 185
R1433 VDD1.n68 VDD1.n67 185
R1434 VDD1.n70 VDD1.n69 185
R1435 VDD1.n63 VDD1.n62 185
R1436 VDD1.n76 VDD1.n75 185
R1437 VDD1.n78 VDD1.n77 185
R1438 VDD1.n59 VDD1.n58 185
R1439 VDD1.n85 VDD1.n84 185
R1440 VDD1.n86 VDD1.n57 185
R1441 VDD1.n88 VDD1.n87 185
R1442 VDD1.n55 VDD1.n54 185
R1443 VDD1.n94 VDD1.n93 185
R1444 VDD1.n96 VDD1.n95 185
R1445 VDD1.n17 VDD1.t1 149.524
R1446 VDD1.n66 VDD1.t6 149.524
R1447 VDD1.n44 VDD1.n43 104.615
R1448 VDD1.n43 VDD1.n3 104.615
R1449 VDD1.n8 VDD1.n3 104.615
R1450 VDD1.n36 VDD1.n8 104.615
R1451 VDD1.n36 VDD1.n35 104.615
R1452 VDD1.n35 VDD1.n9 104.615
R1453 VDD1.n28 VDD1.n9 104.615
R1454 VDD1.n28 VDD1.n27 104.615
R1455 VDD1.n27 VDD1.n13 104.615
R1456 VDD1.n20 VDD1.n13 104.615
R1457 VDD1.n20 VDD1.n19 104.615
R1458 VDD1.n69 VDD1.n68 104.615
R1459 VDD1.n69 VDD1.n62 104.615
R1460 VDD1.n76 VDD1.n62 104.615
R1461 VDD1.n77 VDD1.n76 104.615
R1462 VDD1.n77 VDD1.n58 104.615
R1463 VDD1.n85 VDD1.n58 104.615
R1464 VDD1.n86 VDD1.n85 104.615
R1465 VDD1.n87 VDD1.n86 104.615
R1466 VDD1.n87 VDD1.n54 104.615
R1467 VDD1.n94 VDD1.n54 104.615
R1468 VDD1.n95 VDD1.n94 104.615
R1469 VDD1.n103 VDD1.n102 65.358
R1470 VDD1.n50 VDD1.n49 64.3596
R1471 VDD1.n105 VDD1.n104 64.3594
R1472 VDD1.n101 VDD1.n100 64.3594
R1473 VDD1.n19 VDD1.t1 52.3082
R1474 VDD1.n68 VDD1.t6 52.3082
R1475 VDD1.n50 VDD1.n48 51.6269
R1476 VDD1.n101 VDD1.n99 51.6269
R1477 VDD1.n105 VDD1.n103 39.7013
R1478 VDD1.n6 VDD1.n4 13.1884
R1479 VDD1.n88 VDD1.n55 13.1884
R1480 VDD1.n42 VDD1.n41 12.8005
R1481 VDD1.n38 VDD1.n37 12.8005
R1482 VDD1.n89 VDD1.n57 12.8005
R1483 VDD1.n93 VDD1.n92 12.8005
R1484 VDD1.n45 VDD1.n2 12.0247
R1485 VDD1.n34 VDD1.n7 12.0247
R1486 VDD1.n84 VDD1.n83 12.0247
R1487 VDD1.n96 VDD1.n53 12.0247
R1488 VDD1.n46 VDD1.n0 11.249
R1489 VDD1.n33 VDD1.n10 11.249
R1490 VDD1.n82 VDD1.n59 11.249
R1491 VDD1.n97 VDD1.n51 11.249
R1492 VDD1.n30 VDD1.n29 10.4732
R1493 VDD1.n79 VDD1.n78 10.4732
R1494 VDD1.n18 VDD1.n17 10.2747
R1495 VDD1.n67 VDD1.n66 10.2747
R1496 VDD1.n26 VDD1.n12 9.69747
R1497 VDD1.n75 VDD1.n61 9.69747
R1498 VDD1.n48 VDD1.n47 9.45567
R1499 VDD1.n99 VDD1.n98 9.45567
R1500 VDD1.n16 VDD1.n15 9.3005
R1501 VDD1.n23 VDD1.n22 9.3005
R1502 VDD1.n25 VDD1.n24 9.3005
R1503 VDD1.n12 VDD1.n11 9.3005
R1504 VDD1.n31 VDD1.n30 9.3005
R1505 VDD1.n33 VDD1.n32 9.3005
R1506 VDD1.n7 VDD1.n5 9.3005
R1507 VDD1.n39 VDD1.n38 9.3005
R1508 VDD1.n47 VDD1.n46 9.3005
R1509 VDD1.n2 VDD1.n1 9.3005
R1510 VDD1.n41 VDD1.n40 9.3005
R1511 VDD1.n98 VDD1.n97 9.3005
R1512 VDD1.n53 VDD1.n52 9.3005
R1513 VDD1.n92 VDD1.n91 9.3005
R1514 VDD1.n65 VDD1.n64 9.3005
R1515 VDD1.n72 VDD1.n71 9.3005
R1516 VDD1.n74 VDD1.n73 9.3005
R1517 VDD1.n61 VDD1.n60 9.3005
R1518 VDD1.n80 VDD1.n79 9.3005
R1519 VDD1.n82 VDD1.n81 9.3005
R1520 VDD1.n83 VDD1.n56 9.3005
R1521 VDD1.n90 VDD1.n89 9.3005
R1522 VDD1.n25 VDD1.n14 8.92171
R1523 VDD1.n74 VDD1.n63 8.92171
R1524 VDD1.n22 VDD1.n21 8.14595
R1525 VDD1.n71 VDD1.n70 8.14595
R1526 VDD1.n18 VDD1.n16 7.3702
R1527 VDD1.n67 VDD1.n65 7.3702
R1528 VDD1.n21 VDD1.n16 5.81868
R1529 VDD1.n70 VDD1.n65 5.81868
R1530 VDD1.n22 VDD1.n14 5.04292
R1531 VDD1.n71 VDD1.n63 5.04292
R1532 VDD1.n26 VDD1.n25 4.26717
R1533 VDD1.n75 VDD1.n74 4.26717
R1534 VDD1.n29 VDD1.n12 3.49141
R1535 VDD1.n78 VDD1.n61 3.49141
R1536 VDD1.n17 VDD1.n15 2.84303
R1537 VDD1.n66 VDD1.n64 2.84303
R1538 VDD1.n48 VDD1.n0 2.71565
R1539 VDD1.n30 VDD1.n10 2.71565
R1540 VDD1.n79 VDD1.n59 2.71565
R1541 VDD1.n99 VDD1.n51 2.71565
R1542 VDD1.n104 VDD1.t5 2.12725
R1543 VDD1.n104 VDD1.t9 2.12725
R1544 VDD1.n49 VDD1.t4 2.12725
R1545 VDD1.n49 VDD1.t8 2.12725
R1546 VDD1.n102 VDD1.t7 2.12725
R1547 VDD1.n102 VDD1.t2 2.12725
R1548 VDD1.n100 VDD1.t3 2.12725
R1549 VDD1.n100 VDD1.t0 2.12725
R1550 VDD1.n46 VDD1.n45 1.93989
R1551 VDD1.n34 VDD1.n33 1.93989
R1552 VDD1.n84 VDD1.n82 1.93989
R1553 VDD1.n97 VDD1.n96 1.93989
R1554 VDD1.n42 VDD1.n2 1.16414
R1555 VDD1.n37 VDD1.n7 1.16414
R1556 VDD1.n83 VDD1.n57 1.16414
R1557 VDD1.n93 VDD1.n53 1.16414
R1558 VDD1 VDD1.n105 0.99619
R1559 VDD1 VDD1.n50 0.409983
R1560 VDD1.n41 VDD1.n4 0.388379
R1561 VDD1.n38 VDD1.n6 0.388379
R1562 VDD1.n89 VDD1.n88 0.388379
R1563 VDD1.n92 VDD1.n55 0.388379
R1564 VDD1.n103 VDD1.n101 0.296447
R1565 VDD1.n47 VDD1.n1 0.155672
R1566 VDD1.n40 VDD1.n1 0.155672
R1567 VDD1.n40 VDD1.n39 0.155672
R1568 VDD1.n39 VDD1.n5 0.155672
R1569 VDD1.n32 VDD1.n5 0.155672
R1570 VDD1.n32 VDD1.n31 0.155672
R1571 VDD1.n31 VDD1.n11 0.155672
R1572 VDD1.n24 VDD1.n11 0.155672
R1573 VDD1.n24 VDD1.n23 0.155672
R1574 VDD1.n23 VDD1.n15 0.155672
R1575 VDD1.n72 VDD1.n64 0.155672
R1576 VDD1.n73 VDD1.n72 0.155672
R1577 VDD1.n73 VDD1.n60 0.155672
R1578 VDD1.n80 VDD1.n60 0.155672
R1579 VDD1.n81 VDD1.n80 0.155672
R1580 VDD1.n81 VDD1.n56 0.155672
R1581 VDD1.n90 VDD1.n56 0.155672
R1582 VDD1.n91 VDD1.n90 0.155672
R1583 VDD1.n91 VDD1.n52 0.155672
R1584 VDD1.n98 VDD1.n52 0.155672
R1585 VTAIL.n208 VTAIL.n164 289.615
R1586 VTAIL.n46 VTAIL.n2 289.615
R1587 VTAIL.n158 VTAIL.n114 289.615
R1588 VTAIL.n104 VTAIL.n60 289.615
R1589 VTAIL.n181 VTAIL.n180 185
R1590 VTAIL.n183 VTAIL.n182 185
R1591 VTAIL.n176 VTAIL.n175 185
R1592 VTAIL.n189 VTAIL.n188 185
R1593 VTAIL.n191 VTAIL.n190 185
R1594 VTAIL.n172 VTAIL.n171 185
R1595 VTAIL.n198 VTAIL.n197 185
R1596 VTAIL.n199 VTAIL.n170 185
R1597 VTAIL.n201 VTAIL.n200 185
R1598 VTAIL.n168 VTAIL.n167 185
R1599 VTAIL.n207 VTAIL.n206 185
R1600 VTAIL.n209 VTAIL.n208 185
R1601 VTAIL.n19 VTAIL.n18 185
R1602 VTAIL.n21 VTAIL.n20 185
R1603 VTAIL.n14 VTAIL.n13 185
R1604 VTAIL.n27 VTAIL.n26 185
R1605 VTAIL.n29 VTAIL.n28 185
R1606 VTAIL.n10 VTAIL.n9 185
R1607 VTAIL.n36 VTAIL.n35 185
R1608 VTAIL.n37 VTAIL.n8 185
R1609 VTAIL.n39 VTAIL.n38 185
R1610 VTAIL.n6 VTAIL.n5 185
R1611 VTAIL.n45 VTAIL.n44 185
R1612 VTAIL.n47 VTAIL.n46 185
R1613 VTAIL.n159 VTAIL.n158 185
R1614 VTAIL.n157 VTAIL.n156 185
R1615 VTAIL.n118 VTAIL.n117 185
R1616 VTAIL.n122 VTAIL.n120 185
R1617 VTAIL.n151 VTAIL.n150 185
R1618 VTAIL.n149 VTAIL.n148 185
R1619 VTAIL.n124 VTAIL.n123 185
R1620 VTAIL.n143 VTAIL.n142 185
R1621 VTAIL.n141 VTAIL.n140 185
R1622 VTAIL.n128 VTAIL.n127 185
R1623 VTAIL.n135 VTAIL.n134 185
R1624 VTAIL.n133 VTAIL.n132 185
R1625 VTAIL.n105 VTAIL.n104 185
R1626 VTAIL.n103 VTAIL.n102 185
R1627 VTAIL.n64 VTAIL.n63 185
R1628 VTAIL.n68 VTAIL.n66 185
R1629 VTAIL.n97 VTAIL.n96 185
R1630 VTAIL.n95 VTAIL.n94 185
R1631 VTAIL.n70 VTAIL.n69 185
R1632 VTAIL.n89 VTAIL.n88 185
R1633 VTAIL.n87 VTAIL.n86 185
R1634 VTAIL.n74 VTAIL.n73 185
R1635 VTAIL.n81 VTAIL.n80 185
R1636 VTAIL.n79 VTAIL.n78 185
R1637 VTAIL.n179 VTAIL.t0 149.524
R1638 VTAIL.n17 VTAIL.t17 149.524
R1639 VTAIL.n131 VTAIL.t16 149.524
R1640 VTAIL.n77 VTAIL.t4 149.524
R1641 VTAIL.n182 VTAIL.n181 104.615
R1642 VTAIL.n182 VTAIL.n175 104.615
R1643 VTAIL.n189 VTAIL.n175 104.615
R1644 VTAIL.n190 VTAIL.n189 104.615
R1645 VTAIL.n190 VTAIL.n171 104.615
R1646 VTAIL.n198 VTAIL.n171 104.615
R1647 VTAIL.n199 VTAIL.n198 104.615
R1648 VTAIL.n200 VTAIL.n199 104.615
R1649 VTAIL.n200 VTAIL.n167 104.615
R1650 VTAIL.n207 VTAIL.n167 104.615
R1651 VTAIL.n208 VTAIL.n207 104.615
R1652 VTAIL.n20 VTAIL.n19 104.615
R1653 VTAIL.n20 VTAIL.n13 104.615
R1654 VTAIL.n27 VTAIL.n13 104.615
R1655 VTAIL.n28 VTAIL.n27 104.615
R1656 VTAIL.n28 VTAIL.n9 104.615
R1657 VTAIL.n36 VTAIL.n9 104.615
R1658 VTAIL.n37 VTAIL.n36 104.615
R1659 VTAIL.n38 VTAIL.n37 104.615
R1660 VTAIL.n38 VTAIL.n5 104.615
R1661 VTAIL.n45 VTAIL.n5 104.615
R1662 VTAIL.n46 VTAIL.n45 104.615
R1663 VTAIL.n158 VTAIL.n157 104.615
R1664 VTAIL.n157 VTAIL.n117 104.615
R1665 VTAIL.n122 VTAIL.n117 104.615
R1666 VTAIL.n150 VTAIL.n122 104.615
R1667 VTAIL.n150 VTAIL.n149 104.615
R1668 VTAIL.n149 VTAIL.n123 104.615
R1669 VTAIL.n142 VTAIL.n123 104.615
R1670 VTAIL.n142 VTAIL.n141 104.615
R1671 VTAIL.n141 VTAIL.n127 104.615
R1672 VTAIL.n134 VTAIL.n127 104.615
R1673 VTAIL.n134 VTAIL.n133 104.615
R1674 VTAIL.n104 VTAIL.n103 104.615
R1675 VTAIL.n103 VTAIL.n63 104.615
R1676 VTAIL.n68 VTAIL.n63 104.615
R1677 VTAIL.n96 VTAIL.n68 104.615
R1678 VTAIL.n96 VTAIL.n95 104.615
R1679 VTAIL.n95 VTAIL.n69 104.615
R1680 VTAIL.n88 VTAIL.n69 104.615
R1681 VTAIL.n88 VTAIL.n87 104.615
R1682 VTAIL.n87 VTAIL.n73 104.615
R1683 VTAIL.n80 VTAIL.n73 104.615
R1684 VTAIL.n80 VTAIL.n79 104.615
R1685 VTAIL.n181 VTAIL.t0 52.3082
R1686 VTAIL.n19 VTAIL.t17 52.3082
R1687 VTAIL.n133 VTAIL.t16 52.3082
R1688 VTAIL.n79 VTAIL.t4 52.3082
R1689 VTAIL.n113 VTAIL.n112 47.6808
R1690 VTAIL.n111 VTAIL.n110 47.6808
R1691 VTAIL.n59 VTAIL.n58 47.6808
R1692 VTAIL.n57 VTAIL.n56 47.6808
R1693 VTAIL.n215 VTAIL.n214 47.6807
R1694 VTAIL.n1 VTAIL.n0 47.6807
R1695 VTAIL.n53 VTAIL.n52 47.6807
R1696 VTAIL.n55 VTAIL.n54 47.6807
R1697 VTAIL.n213 VTAIL.n212 33.5429
R1698 VTAIL.n51 VTAIL.n50 33.5429
R1699 VTAIL.n163 VTAIL.n162 33.5429
R1700 VTAIL.n109 VTAIL.n108 33.5429
R1701 VTAIL.n57 VTAIL.n55 23.2031
R1702 VTAIL.n213 VTAIL.n163 21.7979
R1703 VTAIL.n201 VTAIL.n168 13.1884
R1704 VTAIL.n39 VTAIL.n6 13.1884
R1705 VTAIL.n120 VTAIL.n118 13.1884
R1706 VTAIL.n66 VTAIL.n64 13.1884
R1707 VTAIL.n202 VTAIL.n170 12.8005
R1708 VTAIL.n206 VTAIL.n205 12.8005
R1709 VTAIL.n40 VTAIL.n8 12.8005
R1710 VTAIL.n44 VTAIL.n43 12.8005
R1711 VTAIL.n156 VTAIL.n155 12.8005
R1712 VTAIL.n152 VTAIL.n151 12.8005
R1713 VTAIL.n102 VTAIL.n101 12.8005
R1714 VTAIL.n98 VTAIL.n97 12.8005
R1715 VTAIL.n197 VTAIL.n196 12.0247
R1716 VTAIL.n209 VTAIL.n166 12.0247
R1717 VTAIL.n35 VTAIL.n34 12.0247
R1718 VTAIL.n47 VTAIL.n4 12.0247
R1719 VTAIL.n159 VTAIL.n116 12.0247
R1720 VTAIL.n148 VTAIL.n121 12.0247
R1721 VTAIL.n105 VTAIL.n62 12.0247
R1722 VTAIL.n94 VTAIL.n67 12.0247
R1723 VTAIL.n195 VTAIL.n172 11.249
R1724 VTAIL.n210 VTAIL.n164 11.249
R1725 VTAIL.n33 VTAIL.n10 11.249
R1726 VTAIL.n48 VTAIL.n2 11.249
R1727 VTAIL.n160 VTAIL.n114 11.249
R1728 VTAIL.n147 VTAIL.n124 11.249
R1729 VTAIL.n106 VTAIL.n60 11.249
R1730 VTAIL.n93 VTAIL.n70 11.249
R1731 VTAIL.n192 VTAIL.n191 10.4732
R1732 VTAIL.n30 VTAIL.n29 10.4732
R1733 VTAIL.n144 VTAIL.n143 10.4732
R1734 VTAIL.n90 VTAIL.n89 10.4732
R1735 VTAIL.n180 VTAIL.n179 10.2747
R1736 VTAIL.n18 VTAIL.n17 10.2747
R1737 VTAIL.n132 VTAIL.n131 10.2747
R1738 VTAIL.n78 VTAIL.n77 10.2747
R1739 VTAIL.n188 VTAIL.n174 9.69747
R1740 VTAIL.n26 VTAIL.n12 9.69747
R1741 VTAIL.n140 VTAIL.n126 9.69747
R1742 VTAIL.n86 VTAIL.n72 9.69747
R1743 VTAIL.n212 VTAIL.n211 9.45567
R1744 VTAIL.n50 VTAIL.n49 9.45567
R1745 VTAIL.n162 VTAIL.n161 9.45567
R1746 VTAIL.n108 VTAIL.n107 9.45567
R1747 VTAIL.n211 VTAIL.n210 9.3005
R1748 VTAIL.n166 VTAIL.n165 9.3005
R1749 VTAIL.n205 VTAIL.n204 9.3005
R1750 VTAIL.n178 VTAIL.n177 9.3005
R1751 VTAIL.n185 VTAIL.n184 9.3005
R1752 VTAIL.n187 VTAIL.n186 9.3005
R1753 VTAIL.n174 VTAIL.n173 9.3005
R1754 VTAIL.n193 VTAIL.n192 9.3005
R1755 VTAIL.n195 VTAIL.n194 9.3005
R1756 VTAIL.n196 VTAIL.n169 9.3005
R1757 VTAIL.n203 VTAIL.n202 9.3005
R1758 VTAIL.n49 VTAIL.n48 9.3005
R1759 VTAIL.n4 VTAIL.n3 9.3005
R1760 VTAIL.n43 VTAIL.n42 9.3005
R1761 VTAIL.n16 VTAIL.n15 9.3005
R1762 VTAIL.n23 VTAIL.n22 9.3005
R1763 VTAIL.n25 VTAIL.n24 9.3005
R1764 VTAIL.n12 VTAIL.n11 9.3005
R1765 VTAIL.n31 VTAIL.n30 9.3005
R1766 VTAIL.n33 VTAIL.n32 9.3005
R1767 VTAIL.n34 VTAIL.n7 9.3005
R1768 VTAIL.n41 VTAIL.n40 9.3005
R1769 VTAIL.n130 VTAIL.n129 9.3005
R1770 VTAIL.n137 VTAIL.n136 9.3005
R1771 VTAIL.n139 VTAIL.n138 9.3005
R1772 VTAIL.n126 VTAIL.n125 9.3005
R1773 VTAIL.n145 VTAIL.n144 9.3005
R1774 VTAIL.n147 VTAIL.n146 9.3005
R1775 VTAIL.n121 VTAIL.n119 9.3005
R1776 VTAIL.n153 VTAIL.n152 9.3005
R1777 VTAIL.n161 VTAIL.n160 9.3005
R1778 VTAIL.n116 VTAIL.n115 9.3005
R1779 VTAIL.n155 VTAIL.n154 9.3005
R1780 VTAIL.n76 VTAIL.n75 9.3005
R1781 VTAIL.n83 VTAIL.n82 9.3005
R1782 VTAIL.n85 VTAIL.n84 9.3005
R1783 VTAIL.n72 VTAIL.n71 9.3005
R1784 VTAIL.n91 VTAIL.n90 9.3005
R1785 VTAIL.n93 VTAIL.n92 9.3005
R1786 VTAIL.n67 VTAIL.n65 9.3005
R1787 VTAIL.n99 VTAIL.n98 9.3005
R1788 VTAIL.n107 VTAIL.n106 9.3005
R1789 VTAIL.n62 VTAIL.n61 9.3005
R1790 VTAIL.n101 VTAIL.n100 9.3005
R1791 VTAIL.n187 VTAIL.n176 8.92171
R1792 VTAIL.n25 VTAIL.n14 8.92171
R1793 VTAIL.n139 VTAIL.n128 8.92171
R1794 VTAIL.n85 VTAIL.n74 8.92171
R1795 VTAIL.n184 VTAIL.n183 8.14595
R1796 VTAIL.n22 VTAIL.n21 8.14595
R1797 VTAIL.n136 VTAIL.n135 8.14595
R1798 VTAIL.n82 VTAIL.n81 8.14595
R1799 VTAIL.n180 VTAIL.n178 7.3702
R1800 VTAIL.n18 VTAIL.n16 7.3702
R1801 VTAIL.n132 VTAIL.n130 7.3702
R1802 VTAIL.n78 VTAIL.n76 7.3702
R1803 VTAIL.n183 VTAIL.n178 5.81868
R1804 VTAIL.n21 VTAIL.n16 5.81868
R1805 VTAIL.n135 VTAIL.n130 5.81868
R1806 VTAIL.n81 VTAIL.n76 5.81868
R1807 VTAIL.n184 VTAIL.n176 5.04292
R1808 VTAIL.n22 VTAIL.n14 5.04292
R1809 VTAIL.n136 VTAIL.n128 5.04292
R1810 VTAIL.n82 VTAIL.n74 5.04292
R1811 VTAIL.n188 VTAIL.n187 4.26717
R1812 VTAIL.n26 VTAIL.n25 4.26717
R1813 VTAIL.n140 VTAIL.n139 4.26717
R1814 VTAIL.n86 VTAIL.n85 4.26717
R1815 VTAIL.n191 VTAIL.n174 3.49141
R1816 VTAIL.n29 VTAIL.n12 3.49141
R1817 VTAIL.n143 VTAIL.n126 3.49141
R1818 VTAIL.n89 VTAIL.n72 3.49141
R1819 VTAIL.n179 VTAIL.n177 2.84303
R1820 VTAIL.n17 VTAIL.n15 2.84303
R1821 VTAIL.n131 VTAIL.n129 2.84303
R1822 VTAIL.n77 VTAIL.n75 2.84303
R1823 VTAIL.n192 VTAIL.n172 2.71565
R1824 VTAIL.n212 VTAIL.n164 2.71565
R1825 VTAIL.n30 VTAIL.n10 2.71565
R1826 VTAIL.n50 VTAIL.n2 2.71565
R1827 VTAIL.n162 VTAIL.n114 2.71565
R1828 VTAIL.n144 VTAIL.n124 2.71565
R1829 VTAIL.n108 VTAIL.n60 2.71565
R1830 VTAIL.n90 VTAIL.n70 2.71565
R1831 VTAIL.n214 VTAIL.t9 2.12725
R1832 VTAIL.n214 VTAIL.t7 2.12725
R1833 VTAIL.n0 VTAIL.t6 2.12725
R1834 VTAIL.n0 VTAIL.t2 2.12725
R1835 VTAIL.n52 VTAIL.t10 2.12725
R1836 VTAIL.n52 VTAIL.t12 2.12725
R1837 VTAIL.n54 VTAIL.t13 2.12725
R1838 VTAIL.n54 VTAIL.t18 2.12725
R1839 VTAIL.n112 VTAIL.t11 2.12725
R1840 VTAIL.n112 VTAIL.t15 2.12725
R1841 VTAIL.n110 VTAIL.t14 2.12725
R1842 VTAIL.n110 VTAIL.t19 2.12725
R1843 VTAIL.n58 VTAIL.t5 2.12725
R1844 VTAIL.n58 VTAIL.t3 2.12725
R1845 VTAIL.n56 VTAIL.t8 2.12725
R1846 VTAIL.n56 VTAIL.t1 2.12725
R1847 VTAIL.n197 VTAIL.n195 1.93989
R1848 VTAIL.n210 VTAIL.n209 1.93989
R1849 VTAIL.n35 VTAIL.n33 1.93989
R1850 VTAIL.n48 VTAIL.n47 1.93989
R1851 VTAIL.n160 VTAIL.n159 1.93989
R1852 VTAIL.n148 VTAIL.n147 1.93989
R1853 VTAIL.n106 VTAIL.n105 1.93989
R1854 VTAIL.n94 VTAIL.n93 1.93989
R1855 VTAIL.n59 VTAIL.n57 1.40567
R1856 VTAIL.n109 VTAIL.n59 1.40567
R1857 VTAIL.n113 VTAIL.n111 1.40567
R1858 VTAIL.n163 VTAIL.n113 1.40567
R1859 VTAIL.n55 VTAIL.n53 1.40567
R1860 VTAIL.n53 VTAIL.n51 1.40567
R1861 VTAIL.n215 VTAIL.n213 1.40567
R1862 VTAIL.n111 VTAIL.n109 1.17291
R1863 VTAIL.n51 VTAIL.n1 1.17291
R1864 VTAIL.n196 VTAIL.n170 1.16414
R1865 VTAIL.n206 VTAIL.n166 1.16414
R1866 VTAIL.n34 VTAIL.n8 1.16414
R1867 VTAIL.n44 VTAIL.n4 1.16414
R1868 VTAIL.n156 VTAIL.n116 1.16414
R1869 VTAIL.n151 VTAIL.n121 1.16414
R1870 VTAIL.n102 VTAIL.n62 1.16414
R1871 VTAIL.n97 VTAIL.n67 1.16414
R1872 VTAIL VTAIL.n1 1.11257
R1873 VTAIL.n202 VTAIL.n201 0.388379
R1874 VTAIL.n205 VTAIL.n168 0.388379
R1875 VTAIL.n40 VTAIL.n39 0.388379
R1876 VTAIL.n43 VTAIL.n6 0.388379
R1877 VTAIL.n155 VTAIL.n118 0.388379
R1878 VTAIL.n152 VTAIL.n120 0.388379
R1879 VTAIL.n101 VTAIL.n64 0.388379
R1880 VTAIL.n98 VTAIL.n66 0.388379
R1881 VTAIL VTAIL.n215 0.293603
R1882 VTAIL.n185 VTAIL.n177 0.155672
R1883 VTAIL.n186 VTAIL.n185 0.155672
R1884 VTAIL.n186 VTAIL.n173 0.155672
R1885 VTAIL.n193 VTAIL.n173 0.155672
R1886 VTAIL.n194 VTAIL.n193 0.155672
R1887 VTAIL.n194 VTAIL.n169 0.155672
R1888 VTAIL.n203 VTAIL.n169 0.155672
R1889 VTAIL.n204 VTAIL.n203 0.155672
R1890 VTAIL.n204 VTAIL.n165 0.155672
R1891 VTAIL.n211 VTAIL.n165 0.155672
R1892 VTAIL.n23 VTAIL.n15 0.155672
R1893 VTAIL.n24 VTAIL.n23 0.155672
R1894 VTAIL.n24 VTAIL.n11 0.155672
R1895 VTAIL.n31 VTAIL.n11 0.155672
R1896 VTAIL.n32 VTAIL.n31 0.155672
R1897 VTAIL.n32 VTAIL.n7 0.155672
R1898 VTAIL.n41 VTAIL.n7 0.155672
R1899 VTAIL.n42 VTAIL.n41 0.155672
R1900 VTAIL.n42 VTAIL.n3 0.155672
R1901 VTAIL.n49 VTAIL.n3 0.155672
R1902 VTAIL.n161 VTAIL.n115 0.155672
R1903 VTAIL.n154 VTAIL.n115 0.155672
R1904 VTAIL.n154 VTAIL.n153 0.155672
R1905 VTAIL.n153 VTAIL.n119 0.155672
R1906 VTAIL.n146 VTAIL.n119 0.155672
R1907 VTAIL.n146 VTAIL.n145 0.155672
R1908 VTAIL.n145 VTAIL.n125 0.155672
R1909 VTAIL.n138 VTAIL.n125 0.155672
R1910 VTAIL.n138 VTAIL.n137 0.155672
R1911 VTAIL.n137 VTAIL.n129 0.155672
R1912 VTAIL.n107 VTAIL.n61 0.155672
R1913 VTAIL.n100 VTAIL.n61 0.155672
R1914 VTAIL.n100 VTAIL.n99 0.155672
R1915 VTAIL.n99 VTAIL.n65 0.155672
R1916 VTAIL.n92 VTAIL.n65 0.155672
R1917 VTAIL.n92 VTAIL.n91 0.155672
R1918 VTAIL.n91 VTAIL.n71 0.155672
R1919 VTAIL.n84 VTAIL.n71 0.155672
R1920 VTAIL.n84 VTAIL.n83 0.155672
R1921 VTAIL.n83 VTAIL.n75 0.155672
R1922 VN.n6 VN.t1 202.195
R1923 VN.n32 VN.t4 202.195
R1924 VN.n24 VN.n23 173.044
R1925 VN.n49 VN.n48 173.044
R1926 VN.n3 VN.t9 172.594
R1927 VN.n5 VN.t5 172.594
R1928 VN.n16 VN.t2 172.594
R1929 VN.n23 VN.t7 172.594
R1930 VN.n29 VN.t8 172.594
R1931 VN.n31 VN.t0 172.594
R1932 VN.n28 VN.t6 172.594
R1933 VN.n48 VN.t3 172.594
R1934 VN.n47 VN.n25 161.3
R1935 VN.n46 VN.n45 161.3
R1936 VN.n44 VN.n26 161.3
R1937 VN.n43 VN.n42 161.3
R1938 VN.n41 VN.n27 161.3
R1939 VN.n40 VN.n39 161.3
R1940 VN.n38 VN.n29 161.3
R1941 VN.n37 VN.n36 161.3
R1942 VN.n35 VN.n30 161.3
R1943 VN.n34 VN.n33 161.3
R1944 VN.n22 VN.n0 161.3
R1945 VN.n21 VN.n20 161.3
R1946 VN.n19 VN.n1 161.3
R1947 VN.n18 VN.n17 161.3
R1948 VN.n15 VN.n2 161.3
R1949 VN.n14 VN.n13 161.3
R1950 VN.n12 VN.n3 161.3
R1951 VN.n11 VN.n10 161.3
R1952 VN.n9 VN.n4 161.3
R1953 VN.n8 VN.n7 161.3
R1954 VN.n6 VN.n5 58.4685
R1955 VN.n32 VN.n31 58.4685
R1956 VN.n10 VN.n9 56.5193
R1957 VN.n15 VN.n14 56.5193
R1958 VN.n36 VN.n35 56.5193
R1959 VN.n41 VN.n40 56.5193
R1960 VN.n21 VN.n1 45.8354
R1961 VN.n46 VN.n26 45.8354
R1962 VN VN.n49 44.3092
R1963 VN.n22 VN.n21 35.1514
R1964 VN.n47 VN.n46 35.1514
R1965 VN.n33 VN.n32 27.0985
R1966 VN.n7 VN.n6 27.0985
R1967 VN.n9 VN.n8 24.4675
R1968 VN.n10 VN.n3 24.4675
R1969 VN.n14 VN.n3 24.4675
R1970 VN.n17 VN.n15 24.4675
R1971 VN.n35 VN.n34 24.4675
R1972 VN.n40 VN.n29 24.4675
R1973 VN.n36 VN.n29 24.4675
R1974 VN.n42 VN.n41 24.4675
R1975 VN.n16 VN.n1 18.1061
R1976 VN.n28 VN.n26 18.1061
R1977 VN.n23 VN.n22 12.7233
R1978 VN.n48 VN.n47 12.7233
R1979 VN.n8 VN.n5 6.36192
R1980 VN.n17 VN.n16 6.36192
R1981 VN.n34 VN.n31 6.36192
R1982 VN.n42 VN.n28 6.36192
R1983 VN.n49 VN.n25 0.189894
R1984 VN.n45 VN.n25 0.189894
R1985 VN.n45 VN.n44 0.189894
R1986 VN.n44 VN.n43 0.189894
R1987 VN.n43 VN.n27 0.189894
R1988 VN.n39 VN.n27 0.189894
R1989 VN.n39 VN.n38 0.189894
R1990 VN.n38 VN.n37 0.189894
R1991 VN.n37 VN.n30 0.189894
R1992 VN.n33 VN.n30 0.189894
R1993 VN.n7 VN.n4 0.189894
R1994 VN.n11 VN.n4 0.189894
R1995 VN.n12 VN.n11 0.189894
R1996 VN.n13 VN.n12 0.189894
R1997 VN.n13 VN.n2 0.189894
R1998 VN.n18 VN.n2 0.189894
R1999 VN.n19 VN.n18 0.189894
R2000 VN.n20 VN.n19 0.189894
R2001 VN.n20 VN.n0 0.189894
R2002 VN.n24 VN.n0 0.189894
R2003 VN VN.n24 0.0516364
R2004 VDD2.n97 VDD2.n53 289.615
R2005 VDD2.n44 VDD2.n0 289.615
R2006 VDD2.n98 VDD2.n97 185
R2007 VDD2.n96 VDD2.n95 185
R2008 VDD2.n57 VDD2.n56 185
R2009 VDD2.n61 VDD2.n59 185
R2010 VDD2.n90 VDD2.n89 185
R2011 VDD2.n88 VDD2.n87 185
R2012 VDD2.n63 VDD2.n62 185
R2013 VDD2.n82 VDD2.n81 185
R2014 VDD2.n80 VDD2.n79 185
R2015 VDD2.n67 VDD2.n66 185
R2016 VDD2.n74 VDD2.n73 185
R2017 VDD2.n72 VDD2.n71 185
R2018 VDD2.n17 VDD2.n16 185
R2019 VDD2.n19 VDD2.n18 185
R2020 VDD2.n12 VDD2.n11 185
R2021 VDD2.n25 VDD2.n24 185
R2022 VDD2.n27 VDD2.n26 185
R2023 VDD2.n8 VDD2.n7 185
R2024 VDD2.n34 VDD2.n33 185
R2025 VDD2.n35 VDD2.n6 185
R2026 VDD2.n37 VDD2.n36 185
R2027 VDD2.n4 VDD2.n3 185
R2028 VDD2.n43 VDD2.n42 185
R2029 VDD2.n45 VDD2.n44 185
R2030 VDD2.n70 VDD2.t6 149.524
R2031 VDD2.n15 VDD2.t8 149.524
R2032 VDD2.n97 VDD2.n96 104.615
R2033 VDD2.n96 VDD2.n56 104.615
R2034 VDD2.n61 VDD2.n56 104.615
R2035 VDD2.n89 VDD2.n61 104.615
R2036 VDD2.n89 VDD2.n88 104.615
R2037 VDD2.n88 VDD2.n62 104.615
R2038 VDD2.n81 VDD2.n62 104.615
R2039 VDD2.n81 VDD2.n80 104.615
R2040 VDD2.n80 VDD2.n66 104.615
R2041 VDD2.n73 VDD2.n66 104.615
R2042 VDD2.n73 VDD2.n72 104.615
R2043 VDD2.n18 VDD2.n17 104.615
R2044 VDD2.n18 VDD2.n11 104.615
R2045 VDD2.n25 VDD2.n11 104.615
R2046 VDD2.n26 VDD2.n25 104.615
R2047 VDD2.n26 VDD2.n7 104.615
R2048 VDD2.n34 VDD2.n7 104.615
R2049 VDD2.n35 VDD2.n34 104.615
R2050 VDD2.n36 VDD2.n35 104.615
R2051 VDD2.n36 VDD2.n3 104.615
R2052 VDD2.n43 VDD2.n3 104.615
R2053 VDD2.n44 VDD2.n43 104.615
R2054 VDD2.n52 VDD2.n51 65.358
R2055 VDD2 VDD2.n105 65.3551
R2056 VDD2.n104 VDD2.n103 64.3596
R2057 VDD2.n50 VDD2.n49 64.3594
R2058 VDD2.n72 VDD2.t6 52.3082
R2059 VDD2.n17 VDD2.t8 52.3082
R2060 VDD2.n50 VDD2.n48 51.6269
R2061 VDD2.n102 VDD2.n101 50.2217
R2062 VDD2.n102 VDD2.n52 38.4157
R2063 VDD2.n59 VDD2.n57 13.1884
R2064 VDD2.n37 VDD2.n4 13.1884
R2065 VDD2.n95 VDD2.n94 12.8005
R2066 VDD2.n91 VDD2.n90 12.8005
R2067 VDD2.n38 VDD2.n6 12.8005
R2068 VDD2.n42 VDD2.n41 12.8005
R2069 VDD2.n98 VDD2.n55 12.0247
R2070 VDD2.n87 VDD2.n60 12.0247
R2071 VDD2.n33 VDD2.n32 12.0247
R2072 VDD2.n45 VDD2.n2 12.0247
R2073 VDD2.n99 VDD2.n53 11.249
R2074 VDD2.n86 VDD2.n63 11.249
R2075 VDD2.n31 VDD2.n8 11.249
R2076 VDD2.n46 VDD2.n0 11.249
R2077 VDD2.n83 VDD2.n82 10.4732
R2078 VDD2.n28 VDD2.n27 10.4732
R2079 VDD2.n71 VDD2.n70 10.2747
R2080 VDD2.n16 VDD2.n15 10.2747
R2081 VDD2.n79 VDD2.n65 9.69747
R2082 VDD2.n24 VDD2.n10 9.69747
R2083 VDD2.n101 VDD2.n100 9.45567
R2084 VDD2.n48 VDD2.n47 9.45567
R2085 VDD2.n69 VDD2.n68 9.3005
R2086 VDD2.n76 VDD2.n75 9.3005
R2087 VDD2.n78 VDD2.n77 9.3005
R2088 VDD2.n65 VDD2.n64 9.3005
R2089 VDD2.n84 VDD2.n83 9.3005
R2090 VDD2.n86 VDD2.n85 9.3005
R2091 VDD2.n60 VDD2.n58 9.3005
R2092 VDD2.n92 VDD2.n91 9.3005
R2093 VDD2.n100 VDD2.n99 9.3005
R2094 VDD2.n55 VDD2.n54 9.3005
R2095 VDD2.n94 VDD2.n93 9.3005
R2096 VDD2.n47 VDD2.n46 9.3005
R2097 VDD2.n2 VDD2.n1 9.3005
R2098 VDD2.n41 VDD2.n40 9.3005
R2099 VDD2.n14 VDD2.n13 9.3005
R2100 VDD2.n21 VDD2.n20 9.3005
R2101 VDD2.n23 VDD2.n22 9.3005
R2102 VDD2.n10 VDD2.n9 9.3005
R2103 VDD2.n29 VDD2.n28 9.3005
R2104 VDD2.n31 VDD2.n30 9.3005
R2105 VDD2.n32 VDD2.n5 9.3005
R2106 VDD2.n39 VDD2.n38 9.3005
R2107 VDD2.n78 VDD2.n67 8.92171
R2108 VDD2.n23 VDD2.n12 8.92171
R2109 VDD2.n75 VDD2.n74 8.14595
R2110 VDD2.n20 VDD2.n19 8.14595
R2111 VDD2.n71 VDD2.n69 7.3702
R2112 VDD2.n16 VDD2.n14 7.3702
R2113 VDD2.n74 VDD2.n69 5.81868
R2114 VDD2.n19 VDD2.n14 5.81868
R2115 VDD2.n75 VDD2.n67 5.04292
R2116 VDD2.n20 VDD2.n12 5.04292
R2117 VDD2.n79 VDD2.n78 4.26717
R2118 VDD2.n24 VDD2.n23 4.26717
R2119 VDD2.n82 VDD2.n65 3.49141
R2120 VDD2.n27 VDD2.n10 3.49141
R2121 VDD2.n70 VDD2.n68 2.84303
R2122 VDD2.n15 VDD2.n13 2.84303
R2123 VDD2.n101 VDD2.n53 2.71565
R2124 VDD2.n83 VDD2.n63 2.71565
R2125 VDD2.n28 VDD2.n8 2.71565
R2126 VDD2.n48 VDD2.n0 2.71565
R2127 VDD2.n105 VDD2.t9 2.12725
R2128 VDD2.n105 VDD2.t5 2.12725
R2129 VDD2.n103 VDD2.t3 2.12725
R2130 VDD2.n103 VDD2.t1 2.12725
R2131 VDD2.n51 VDD2.t7 2.12725
R2132 VDD2.n51 VDD2.t2 2.12725
R2133 VDD2.n49 VDD2.t4 2.12725
R2134 VDD2.n49 VDD2.t0 2.12725
R2135 VDD2.n99 VDD2.n98 1.93989
R2136 VDD2.n87 VDD2.n86 1.93989
R2137 VDD2.n33 VDD2.n31 1.93989
R2138 VDD2.n46 VDD2.n45 1.93989
R2139 VDD2.n104 VDD2.n102 1.40567
R2140 VDD2.n95 VDD2.n55 1.16414
R2141 VDD2.n90 VDD2.n60 1.16414
R2142 VDD2.n32 VDD2.n6 1.16414
R2143 VDD2.n42 VDD2.n2 1.16414
R2144 VDD2 VDD2.n104 0.409983
R2145 VDD2.n94 VDD2.n57 0.388379
R2146 VDD2.n91 VDD2.n59 0.388379
R2147 VDD2.n38 VDD2.n37 0.388379
R2148 VDD2.n41 VDD2.n4 0.388379
R2149 VDD2.n52 VDD2.n50 0.296447
R2150 VDD2.n100 VDD2.n54 0.155672
R2151 VDD2.n93 VDD2.n54 0.155672
R2152 VDD2.n93 VDD2.n92 0.155672
R2153 VDD2.n92 VDD2.n58 0.155672
R2154 VDD2.n85 VDD2.n58 0.155672
R2155 VDD2.n85 VDD2.n84 0.155672
R2156 VDD2.n84 VDD2.n64 0.155672
R2157 VDD2.n77 VDD2.n64 0.155672
R2158 VDD2.n77 VDD2.n76 0.155672
R2159 VDD2.n76 VDD2.n68 0.155672
R2160 VDD2.n21 VDD2.n13 0.155672
R2161 VDD2.n22 VDD2.n21 0.155672
R2162 VDD2.n22 VDD2.n9 0.155672
R2163 VDD2.n29 VDD2.n9 0.155672
R2164 VDD2.n30 VDD2.n29 0.155672
R2165 VDD2.n30 VDD2.n5 0.155672
R2166 VDD2.n39 VDD2.n5 0.155672
R2167 VDD2.n40 VDD2.n39 0.155672
R2168 VDD2.n40 VDD2.n1 0.155672
R2169 VDD2.n47 VDD2.n1 0.155672
C0 VDD2 VP 0.41751f
C1 VN VTAIL 7.15237f
C2 VDD2 VDD1 1.34319f
C3 VP VTAIL 7.16675f
C4 VN VP 5.98487f
C5 VDD1 VTAIL 9.50906f
C6 VN VDD1 0.150322f
C7 VDD2 VTAIL 9.55023f
C8 VDD1 VP 7.207221f
C9 VDD2 VN 6.943491f
C10 VDD2 B 5.193217f
C11 VDD1 B 5.157248f
C12 VTAIL B 6.103149f
C13 VN B 11.828039f
C14 VP B 10.209024f
C15 VDD2.n0 B 0.030685f
C16 VDD2.n1 B 0.022816f
C17 VDD2.n2 B 0.012261f
C18 VDD2.n3 B 0.028979f
C19 VDD2.n4 B 0.012621f
C20 VDD2.n5 B 0.022816f
C21 VDD2.n6 B 0.012982f
C22 VDD2.n7 B 0.028979f
C23 VDD2.n8 B 0.012982f
C24 VDD2.n9 B 0.022816f
C25 VDD2.n10 B 0.012261f
C26 VDD2.n11 B 0.028979f
C27 VDD2.n12 B 0.012982f
C28 VDD2.n13 B 0.878042f
C29 VDD2.n14 B 0.012261f
C30 VDD2.t8 B 0.048617f
C31 VDD2.n15 B 0.140946f
C32 VDD2.n16 B 0.020486f
C33 VDD2.n17 B 0.021735f
C34 VDD2.n18 B 0.028979f
C35 VDD2.n19 B 0.012982f
C36 VDD2.n20 B 0.012261f
C37 VDD2.n21 B 0.022816f
C38 VDD2.n22 B 0.022816f
C39 VDD2.n23 B 0.012261f
C40 VDD2.n24 B 0.012982f
C41 VDD2.n25 B 0.028979f
C42 VDD2.n26 B 0.028979f
C43 VDD2.n27 B 0.012982f
C44 VDD2.n28 B 0.012261f
C45 VDD2.n29 B 0.022816f
C46 VDD2.n30 B 0.022816f
C47 VDD2.n31 B 0.012261f
C48 VDD2.n32 B 0.012261f
C49 VDD2.n33 B 0.012982f
C50 VDD2.n34 B 0.028979f
C51 VDD2.n35 B 0.028979f
C52 VDD2.n36 B 0.028979f
C53 VDD2.n37 B 0.012621f
C54 VDD2.n38 B 0.012261f
C55 VDD2.n39 B 0.022816f
C56 VDD2.n40 B 0.022816f
C57 VDD2.n41 B 0.012261f
C58 VDD2.n42 B 0.012982f
C59 VDD2.n43 B 0.028979f
C60 VDD2.n44 B 0.060285f
C61 VDD2.n45 B 0.012982f
C62 VDD2.n46 B 0.012261f
C63 VDD2.n47 B 0.054921f
C64 VDD2.n48 B 0.053325f
C65 VDD2.t4 B 0.167861f
C66 VDD2.t0 B 0.167861f
C67 VDD2.n49 B 1.47136f
C68 VDD2.n50 B 0.455223f
C69 VDD2.t7 B 0.167861f
C70 VDD2.t2 B 0.167861f
C71 VDD2.n51 B 1.47701f
C72 VDD2.n52 B 1.87552f
C73 VDD2.n53 B 0.030685f
C74 VDD2.n54 B 0.022816f
C75 VDD2.n55 B 0.012261f
C76 VDD2.n56 B 0.028979f
C77 VDD2.n57 B 0.012621f
C78 VDD2.n58 B 0.022816f
C79 VDD2.n59 B 0.012621f
C80 VDD2.n60 B 0.012261f
C81 VDD2.n61 B 0.028979f
C82 VDD2.n62 B 0.028979f
C83 VDD2.n63 B 0.012982f
C84 VDD2.n64 B 0.022816f
C85 VDD2.n65 B 0.012261f
C86 VDD2.n66 B 0.028979f
C87 VDD2.n67 B 0.012982f
C88 VDD2.n68 B 0.878042f
C89 VDD2.n69 B 0.012261f
C90 VDD2.t6 B 0.048617f
C91 VDD2.n70 B 0.140946f
C92 VDD2.n71 B 0.020486f
C93 VDD2.n72 B 0.021735f
C94 VDD2.n73 B 0.028979f
C95 VDD2.n74 B 0.012982f
C96 VDD2.n75 B 0.012261f
C97 VDD2.n76 B 0.022816f
C98 VDD2.n77 B 0.022816f
C99 VDD2.n78 B 0.012261f
C100 VDD2.n79 B 0.012982f
C101 VDD2.n80 B 0.028979f
C102 VDD2.n81 B 0.028979f
C103 VDD2.n82 B 0.012982f
C104 VDD2.n83 B 0.012261f
C105 VDD2.n84 B 0.022816f
C106 VDD2.n85 B 0.022816f
C107 VDD2.n86 B 0.012261f
C108 VDD2.n87 B 0.012982f
C109 VDD2.n88 B 0.028979f
C110 VDD2.n89 B 0.028979f
C111 VDD2.n90 B 0.012982f
C112 VDD2.n91 B 0.012261f
C113 VDD2.n92 B 0.022816f
C114 VDD2.n93 B 0.022816f
C115 VDD2.n94 B 0.012261f
C116 VDD2.n95 B 0.012982f
C117 VDD2.n96 B 0.028979f
C118 VDD2.n97 B 0.060285f
C119 VDD2.n98 B 0.012982f
C120 VDD2.n99 B 0.012261f
C121 VDD2.n100 B 0.054921f
C122 VDD2.n101 B 0.049284f
C123 VDD2.n102 B 1.98682f
C124 VDD2.t3 B 0.167861f
C125 VDD2.t1 B 0.167861f
C126 VDD2.n103 B 1.47136f
C127 VDD2.n104 B 0.317327f
C128 VDD2.t9 B 0.167861f
C129 VDD2.t5 B 0.167861f
C130 VDD2.n105 B 1.47699f
C131 VN.n0 B 0.032876f
C132 VN.t7 B 1.07516f
C133 VN.n1 B 0.055099f
C134 VN.n2 B 0.032876f
C135 VN.t9 B 1.07516f
C136 VN.n3 B 0.432967f
C137 VN.n4 B 0.032876f
C138 VN.t5 B 1.07516f
C139 VN.n5 B 0.448231f
C140 VN.t1 B 1.14936f
C141 VN.n6 B 0.478503f
C142 VN.n7 B 0.173603f
C143 VN.n8 B 0.038887f
C144 VN.n9 B 0.042041f
C145 VN.n10 B 0.05395f
C146 VN.n11 B 0.032876f
C147 VN.n12 B 0.032876f
C148 VN.n13 B 0.032876f
C149 VN.n14 B 0.05395f
C150 VN.n15 B 0.042041f
C151 VN.t2 B 1.07516f
C152 VN.n16 B 0.401946f
C153 VN.n17 B 0.038887f
C154 VN.n18 B 0.032876f
C155 VN.n19 B 0.032876f
C156 VN.n20 B 0.032876f
C157 VN.n21 B 0.027878f
C158 VN.n22 B 0.051901f
C159 VN.n23 B 0.462443f
C160 VN.n24 B 0.029882f
C161 VN.n25 B 0.032876f
C162 VN.t3 B 1.07516f
C163 VN.n26 B 0.055099f
C164 VN.n27 B 0.032876f
C165 VN.t6 B 1.07516f
C166 VN.n28 B 0.401946f
C167 VN.t8 B 1.07516f
C168 VN.n29 B 0.432967f
C169 VN.n30 B 0.032876f
C170 VN.t0 B 1.07516f
C171 VN.n31 B 0.448231f
C172 VN.t4 B 1.14936f
C173 VN.n32 B 0.478503f
C174 VN.n33 B 0.173603f
C175 VN.n34 B 0.038887f
C176 VN.n35 B 0.042041f
C177 VN.n36 B 0.05395f
C178 VN.n37 B 0.032876f
C179 VN.n38 B 0.032876f
C180 VN.n39 B 0.032876f
C181 VN.n40 B 0.05395f
C182 VN.n41 B 0.042041f
C183 VN.n42 B 0.038887f
C184 VN.n43 B 0.032876f
C185 VN.n44 B 0.032876f
C186 VN.n45 B 0.032876f
C187 VN.n46 B 0.027878f
C188 VN.n47 B 0.051901f
C189 VN.n48 B 0.462443f
C190 VN.n49 B 1.48675f
C191 VTAIL.t6 B 0.186045f
C192 VTAIL.t2 B 0.186045f
C193 VTAIL.n0 B 1.56113f
C194 VTAIL.n1 B 0.425245f
C195 VTAIL.n2 B 0.034009f
C196 VTAIL.n3 B 0.025288f
C197 VTAIL.n4 B 0.013589f
C198 VTAIL.n5 B 0.032119f
C199 VTAIL.n6 B 0.013988f
C200 VTAIL.n7 B 0.025288f
C201 VTAIL.n8 B 0.014388f
C202 VTAIL.n9 B 0.032119f
C203 VTAIL.n10 B 0.014388f
C204 VTAIL.n11 B 0.025288f
C205 VTAIL.n12 B 0.013589f
C206 VTAIL.n13 B 0.032119f
C207 VTAIL.n14 B 0.014388f
C208 VTAIL.n15 B 0.973161f
C209 VTAIL.n16 B 0.013589f
C210 VTAIL.t17 B 0.053884f
C211 VTAIL.n17 B 0.156215f
C212 VTAIL.n18 B 0.022705f
C213 VTAIL.n19 B 0.024089f
C214 VTAIL.n20 B 0.032119f
C215 VTAIL.n21 B 0.014388f
C216 VTAIL.n22 B 0.013589f
C217 VTAIL.n23 B 0.025288f
C218 VTAIL.n24 B 0.025288f
C219 VTAIL.n25 B 0.013589f
C220 VTAIL.n26 B 0.014388f
C221 VTAIL.n27 B 0.032119f
C222 VTAIL.n28 B 0.032119f
C223 VTAIL.n29 B 0.014388f
C224 VTAIL.n30 B 0.013589f
C225 VTAIL.n31 B 0.025288f
C226 VTAIL.n32 B 0.025288f
C227 VTAIL.n33 B 0.013589f
C228 VTAIL.n34 B 0.013589f
C229 VTAIL.n35 B 0.014388f
C230 VTAIL.n36 B 0.032119f
C231 VTAIL.n37 B 0.032119f
C232 VTAIL.n38 B 0.032119f
C233 VTAIL.n39 B 0.013988f
C234 VTAIL.n40 B 0.013589f
C235 VTAIL.n41 B 0.025288f
C236 VTAIL.n42 B 0.025288f
C237 VTAIL.n43 B 0.013589f
C238 VTAIL.n44 B 0.014388f
C239 VTAIL.n45 B 0.032119f
C240 VTAIL.n46 B 0.066816f
C241 VTAIL.n47 B 0.014388f
C242 VTAIL.n48 B 0.013589f
C243 VTAIL.n49 B 0.06087f
C244 VTAIL.n50 B 0.03718f
C245 VTAIL.n51 B 0.232995f
C246 VTAIL.t10 B 0.186045f
C247 VTAIL.t12 B 0.186045f
C248 VTAIL.n52 B 1.56113f
C249 VTAIL.n53 B 0.468094f
C250 VTAIL.t13 B 0.186045f
C251 VTAIL.t18 B 0.186045f
C252 VTAIL.n54 B 1.56113f
C253 VTAIL.n55 B 1.58008f
C254 VTAIL.t8 B 0.186045f
C255 VTAIL.t1 B 0.186045f
C256 VTAIL.n56 B 1.56113f
C257 VTAIL.n57 B 1.58007f
C258 VTAIL.t5 B 0.186045f
C259 VTAIL.t3 B 0.186045f
C260 VTAIL.n58 B 1.56113f
C261 VTAIL.n59 B 0.468084f
C262 VTAIL.n60 B 0.034009f
C263 VTAIL.n61 B 0.025288f
C264 VTAIL.n62 B 0.013589f
C265 VTAIL.n63 B 0.032119f
C266 VTAIL.n64 B 0.013988f
C267 VTAIL.n65 B 0.025288f
C268 VTAIL.n66 B 0.013988f
C269 VTAIL.n67 B 0.013589f
C270 VTAIL.n68 B 0.032119f
C271 VTAIL.n69 B 0.032119f
C272 VTAIL.n70 B 0.014388f
C273 VTAIL.n71 B 0.025288f
C274 VTAIL.n72 B 0.013589f
C275 VTAIL.n73 B 0.032119f
C276 VTAIL.n74 B 0.014388f
C277 VTAIL.n75 B 0.973161f
C278 VTAIL.n76 B 0.013589f
C279 VTAIL.t4 B 0.053884f
C280 VTAIL.n77 B 0.156215f
C281 VTAIL.n78 B 0.022705f
C282 VTAIL.n79 B 0.024089f
C283 VTAIL.n80 B 0.032119f
C284 VTAIL.n81 B 0.014388f
C285 VTAIL.n82 B 0.013589f
C286 VTAIL.n83 B 0.025288f
C287 VTAIL.n84 B 0.025288f
C288 VTAIL.n85 B 0.013589f
C289 VTAIL.n86 B 0.014388f
C290 VTAIL.n87 B 0.032119f
C291 VTAIL.n88 B 0.032119f
C292 VTAIL.n89 B 0.014388f
C293 VTAIL.n90 B 0.013589f
C294 VTAIL.n91 B 0.025288f
C295 VTAIL.n92 B 0.025288f
C296 VTAIL.n93 B 0.013589f
C297 VTAIL.n94 B 0.014388f
C298 VTAIL.n95 B 0.032119f
C299 VTAIL.n96 B 0.032119f
C300 VTAIL.n97 B 0.014388f
C301 VTAIL.n98 B 0.013589f
C302 VTAIL.n99 B 0.025288f
C303 VTAIL.n100 B 0.025288f
C304 VTAIL.n101 B 0.013589f
C305 VTAIL.n102 B 0.014388f
C306 VTAIL.n103 B 0.032119f
C307 VTAIL.n104 B 0.066816f
C308 VTAIL.n105 B 0.014388f
C309 VTAIL.n106 B 0.013589f
C310 VTAIL.n107 B 0.06087f
C311 VTAIL.n108 B 0.03718f
C312 VTAIL.n109 B 0.232995f
C313 VTAIL.t14 B 0.186045f
C314 VTAIL.t19 B 0.186045f
C315 VTAIL.n110 B 1.56113f
C316 VTAIL.n111 B 0.449118f
C317 VTAIL.t11 B 0.186045f
C318 VTAIL.t15 B 0.186045f
C319 VTAIL.n112 B 1.56113f
C320 VTAIL.n113 B 0.468084f
C321 VTAIL.n114 B 0.034009f
C322 VTAIL.n115 B 0.025288f
C323 VTAIL.n116 B 0.013589f
C324 VTAIL.n117 B 0.032119f
C325 VTAIL.n118 B 0.013988f
C326 VTAIL.n119 B 0.025288f
C327 VTAIL.n120 B 0.013988f
C328 VTAIL.n121 B 0.013589f
C329 VTAIL.n122 B 0.032119f
C330 VTAIL.n123 B 0.032119f
C331 VTAIL.n124 B 0.014388f
C332 VTAIL.n125 B 0.025288f
C333 VTAIL.n126 B 0.013589f
C334 VTAIL.n127 B 0.032119f
C335 VTAIL.n128 B 0.014388f
C336 VTAIL.n129 B 0.973161f
C337 VTAIL.n130 B 0.013589f
C338 VTAIL.t16 B 0.053884f
C339 VTAIL.n131 B 0.156215f
C340 VTAIL.n132 B 0.022705f
C341 VTAIL.n133 B 0.024089f
C342 VTAIL.n134 B 0.032119f
C343 VTAIL.n135 B 0.014388f
C344 VTAIL.n136 B 0.013589f
C345 VTAIL.n137 B 0.025288f
C346 VTAIL.n138 B 0.025288f
C347 VTAIL.n139 B 0.013589f
C348 VTAIL.n140 B 0.014388f
C349 VTAIL.n141 B 0.032119f
C350 VTAIL.n142 B 0.032119f
C351 VTAIL.n143 B 0.014388f
C352 VTAIL.n144 B 0.013589f
C353 VTAIL.n145 B 0.025288f
C354 VTAIL.n146 B 0.025288f
C355 VTAIL.n147 B 0.013589f
C356 VTAIL.n148 B 0.014388f
C357 VTAIL.n149 B 0.032119f
C358 VTAIL.n150 B 0.032119f
C359 VTAIL.n151 B 0.014388f
C360 VTAIL.n152 B 0.013589f
C361 VTAIL.n153 B 0.025288f
C362 VTAIL.n154 B 0.025288f
C363 VTAIL.n155 B 0.013589f
C364 VTAIL.n156 B 0.014388f
C365 VTAIL.n157 B 0.032119f
C366 VTAIL.n158 B 0.066816f
C367 VTAIL.n159 B 0.014388f
C368 VTAIL.n160 B 0.013589f
C369 VTAIL.n161 B 0.06087f
C370 VTAIL.n162 B 0.03718f
C371 VTAIL.n163 B 1.24945f
C372 VTAIL.n164 B 0.034009f
C373 VTAIL.n165 B 0.025288f
C374 VTAIL.n166 B 0.013589f
C375 VTAIL.n167 B 0.032119f
C376 VTAIL.n168 B 0.013988f
C377 VTAIL.n169 B 0.025288f
C378 VTAIL.n170 B 0.014388f
C379 VTAIL.n171 B 0.032119f
C380 VTAIL.n172 B 0.014388f
C381 VTAIL.n173 B 0.025288f
C382 VTAIL.n174 B 0.013589f
C383 VTAIL.n175 B 0.032119f
C384 VTAIL.n176 B 0.014388f
C385 VTAIL.n177 B 0.973161f
C386 VTAIL.n178 B 0.013589f
C387 VTAIL.t0 B 0.053884f
C388 VTAIL.n179 B 0.156215f
C389 VTAIL.n180 B 0.022705f
C390 VTAIL.n181 B 0.024089f
C391 VTAIL.n182 B 0.032119f
C392 VTAIL.n183 B 0.014388f
C393 VTAIL.n184 B 0.013589f
C394 VTAIL.n185 B 0.025288f
C395 VTAIL.n186 B 0.025288f
C396 VTAIL.n187 B 0.013589f
C397 VTAIL.n188 B 0.014388f
C398 VTAIL.n189 B 0.032119f
C399 VTAIL.n190 B 0.032119f
C400 VTAIL.n191 B 0.014388f
C401 VTAIL.n192 B 0.013589f
C402 VTAIL.n193 B 0.025288f
C403 VTAIL.n194 B 0.025288f
C404 VTAIL.n195 B 0.013589f
C405 VTAIL.n196 B 0.013589f
C406 VTAIL.n197 B 0.014388f
C407 VTAIL.n198 B 0.032119f
C408 VTAIL.n199 B 0.032119f
C409 VTAIL.n200 B 0.032119f
C410 VTAIL.n201 B 0.013988f
C411 VTAIL.n202 B 0.013589f
C412 VTAIL.n203 B 0.025288f
C413 VTAIL.n204 B 0.025288f
C414 VTAIL.n205 B 0.013589f
C415 VTAIL.n206 B 0.014388f
C416 VTAIL.n207 B 0.032119f
C417 VTAIL.n208 B 0.066816f
C418 VTAIL.n209 B 0.014388f
C419 VTAIL.n210 B 0.013589f
C420 VTAIL.n211 B 0.06087f
C421 VTAIL.n212 B 0.03718f
C422 VTAIL.n213 B 1.24945f
C423 VTAIL.t9 B 0.186045f
C424 VTAIL.t7 B 0.186045f
C425 VTAIL.n214 B 1.56113f
C426 VTAIL.n215 B 0.377478f
C427 VDD1.n0 B 0.030899f
C428 VDD1.n1 B 0.022976f
C429 VDD1.n2 B 0.012346f
C430 VDD1.n3 B 0.029182f
C431 VDD1.n4 B 0.012709f
C432 VDD1.n5 B 0.022976f
C433 VDD1.n6 B 0.012709f
C434 VDD1.n7 B 0.012346f
C435 VDD1.n8 B 0.029182f
C436 VDD1.n9 B 0.029182f
C437 VDD1.n10 B 0.013072f
C438 VDD1.n11 B 0.022976f
C439 VDD1.n12 B 0.012346f
C440 VDD1.n13 B 0.029182f
C441 VDD1.n14 B 0.013072f
C442 VDD1.n15 B 0.88417f
C443 VDD1.n16 B 0.012346f
C444 VDD1.t1 B 0.048957f
C445 VDD1.n17 B 0.14193f
C446 VDD1.n18 B 0.020629f
C447 VDD1.n19 B 0.021886f
C448 VDD1.n20 B 0.029182f
C449 VDD1.n21 B 0.013072f
C450 VDD1.n22 B 0.012346f
C451 VDD1.n23 B 0.022976f
C452 VDD1.n24 B 0.022976f
C453 VDD1.n25 B 0.012346f
C454 VDD1.n26 B 0.013072f
C455 VDD1.n27 B 0.029182f
C456 VDD1.n28 B 0.029182f
C457 VDD1.n29 B 0.013072f
C458 VDD1.n30 B 0.012346f
C459 VDD1.n31 B 0.022976f
C460 VDD1.n32 B 0.022976f
C461 VDD1.n33 B 0.012346f
C462 VDD1.n34 B 0.013072f
C463 VDD1.n35 B 0.029182f
C464 VDD1.n36 B 0.029182f
C465 VDD1.n37 B 0.013072f
C466 VDD1.n38 B 0.012346f
C467 VDD1.n39 B 0.022976f
C468 VDD1.n40 B 0.022976f
C469 VDD1.n41 B 0.012346f
C470 VDD1.n42 B 0.013072f
C471 VDD1.n43 B 0.029182f
C472 VDD1.n44 B 0.060706f
C473 VDD1.n45 B 0.013072f
C474 VDD1.n46 B 0.012346f
C475 VDD1.n47 B 0.055304f
C476 VDD1.n48 B 0.053697f
C477 VDD1.t4 B 0.169032f
C478 VDD1.t8 B 0.169032f
C479 VDD1.n49 B 1.48163f
C480 VDD1.n50 B 0.464999f
C481 VDD1.n51 B 0.030899f
C482 VDD1.n52 B 0.022976f
C483 VDD1.n53 B 0.012346f
C484 VDD1.n54 B 0.029182f
C485 VDD1.n55 B 0.012709f
C486 VDD1.n56 B 0.022976f
C487 VDD1.n57 B 0.013072f
C488 VDD1.n58 B 0.029182f
C489 VDD1.n59 B 0.013072f
C490 VDD1.n60 B 0.022976f
C491 VDD1.n61 B 0.012346f
C492 VDD1.n62 B 0.029182f
C493 VDD1.n63 B 0.013072f
C494 VDD1.n64 B 0.88417f
C495 VDD1.n65 B 0.012346f
C496 VDD1.t6 B 0.048957f
C497 VDD1.n66 B 0.14193f
C498 VDD1.n67 B 0.020629f
C499 VDD1.n68 B 0.021886f
C500 VDD1.n69 B 0.029182f
C501 VDD1.n70 B 0.013072f
C502 VDD1.n71 B 0.012346f
C503 VDD1.n72 B 0.022976f
C504 VDD1.n73 B 0.022976f
C505 VDD1.n74 B 0.012346f
C506 VDD1.n75 B 0.013072f
C507 VDD1.n76 B 0.029182f
C508 VDD1.n77 B 0.029182f
C509 VDD1.n78 B 0.013072f
C510 VDD1.n79 B 0.012346f
C511 VDD1.n80 B 0.022976f
C512 VDD1.n81 B 0.022976f
C513 VDD1.n82 B 0.012346f
C514 VDD1.n83 B 0.012346f
C515 VDD1.n84 B 0.013072f
C516 VDD1.n85 B 0.029182f
C517 VDD1.n86 B 0.029182f
C518 VDD1.n87 B 0.029182f
C519 VDD1.n88 B 0.012709f
C520 VDD1.n89 B 0.012346f
C521 VDD1.n90 B 0.022976f
C522 VDD1.n91 B 0.022976f
C523 VDD1.n92 B 0.012346f
C524 VDD1.n93 B 0.013072f
C525 VDD1.n94 B 0.029182f
C526 VDD1.n95 B 0.060706f
C527 VDD1.n96 B 0.013072f
C528 VDD1.n97 B 0.012346f
C529 VDD1.n98 B 0.055304f
C530 VDD1.n99 B 0.053697f
C531 VDD1.t3 B 0.169032f
C532 VDD1.t0 B 0.169032f
C533 VDD1.n100 B 1.48162f
C534 VDD1.n101 B 0.4584f
C535 VDD1.t7 B 0.169032f
C536 VDD1.t2 B 0.169032f
C537 VDD1.n102 B 1.48732f
C538 VDD1.n103 B 1.97139f
C539 VDD1.t5 B 0.169032f
C540 VDD1.t9 B 0.169032f
C541 VDD1.n104 B 1.48162f
C542 VDD1.n105 B 2.22543f
C543 VP.n0 B 0.033443f
C544 VP.t2 B 1.09372f
C545 VP.n1 B 0.05605f
C546 VP.n2 B 0.033443f
C547 VP.t9 B 1.09372f
C548 VP.n3 B 0.440442f
C549 VP.n4 B 0.033443f
C550 VP.t1 B 1.09372f
C551 VP.n5 B 0.408885f
C552 VP.n6 B 0.033443f
C553 VP.t6 B 1.09372f
C554 VP.n7 B 0.470427f
C555 VP.n8 B 0.033443f
C556 VP.t3 B 1.09372f
C557 VP.n9 B 0.05605f
C558 VP.n10 B 0.033443f
C559 VP.t8 B 1.09372f
C560 VP.n11 B 0.440442f
C561 VP.n12 B 0.033443f
C562 VP.t0 B 1.09372f
C563 VP.n13 B 0.455969f
C564 VP.t5 B 1.16921f
C565 VP.n14 B 0.486764f
C566 VP.n15 B 0.1766f
C567 VP.n16 B 0.039558f
C568 VP.n17 B 0.042767f
C569 VP.n18 B 0.054882f
C570 VP.n19 B 0.033443f
C571 VP.n20 B 0.033443f
C572 VP.n21 B 0.033443f
C573 VP.n22 B 0.054882f
C574 VP.n23 B 0.042767f
C575 VP.t4 B 1.09372f
C576 VP.n24 B 0.408885f
C577 VP.n25 B 0.039558f
C578 VP.n26 B 0.033443f
C579 VP.n27 B 0.033443f
C580 VP.n28 B 0.033443f
C581 VP.n29 B 0.028359f
C582 VP.n30 B 0.052797f
C583 VP.n31 B 0.470427f
C584 VP.n32 B 1.49052f
C585 VP.n33 B 1.51789f
C586 VP.n34 B 0.033443f
C587 VP.n35 B 0.052797f
C588 VP.n36 B 0.028359f
C589 VP.n37 B 0.05605f
C590 VP.n38 B 0.033443f
C591 VP.n39 B 0.033443f
C592 VP.n40 B 0.039558f
C593 VP.n41 B 0.042767f
C594 VP.n42 B 0.054882f
C595 VP.n43 B 0.033443f
C596 VP.n44 B 0.033443f
C597 VP.n45 B 0.033443f
C598 VP.n46 B 0.054882f
C599 VP.n47 B 0.042767f
C600 VP.t7 B 1.09372f
C601 VP.n48 B 0.408885f
C602 VP.n49 B 0.039558f
C603 VP.n50 B 0.033443f
C604 VP.n51 B 0.033443f
C605 VP.n52 B 0.033443f
C606 VP.n53 B 0.028359f
C607 VP.n54 B 0.052797f
C608 VP.n55 B 0.470427f
C609 VP.n56 B 0.030398f
.ends

