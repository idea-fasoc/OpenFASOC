* NGSPICE file created from diff_pair_sample_0612.ext - technology: sky130A

.subckt diff_pair_sample_0612 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=4.641 ps=24.58 w=11.9 l=0.96
X1 VDD1.t1 VP.t0 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=4.641 ps=24.58 w=11.9 l=0.96
X2 B.t15 B.t13 B.t14 B.t10 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=0 ps=0 w=11.9 l=0.96
X3 B.t12 B.t9 B.t11 B.t10 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=0 ps=0 w=11.9 l=0.96
X4 B.t8 B.t6 B.t7 B.t3 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=0 ps=0 w=11.9 l=0.96
X5 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=0 ps=0 w=11.9 l=0.96
X6 VDD2.t0 VN.t1 VTAIL.t2 B.t1 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=4.641 ps=24.58 w=11.9 l=0.96
X7 VDD1.t0 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=4.641 pd=24.58 as=4.641 ps=24.58 w=11.9 l=0.96
R0 VN VN.t0 542.088
R1 VN VN.t1 501.514
R2 VTAIL.n262 VTAIL.n261 289.615
R3 VTAIL.n64 VTAIL.n63 289.615
R4 VTAIL.n196 VTAIL.n195 289.615
R5 VTAIL.n130 VTAIL.n129 289.615
R6 VTAIL.n221 VTAIL.n220 185
R7 VTAIL.n223 VTAIL.n222 185
R8 VTAIL.n216 VTAIL.n215 185
R9 VTAIL.n229 VTAIL.n228 185
R10 VTAIL.n231 VTAIL.n230 185
R11 VTAIL.n212 VTAIL.n211 185
R12 VTAIL.n237 VTAIL.n236 185
R13 VTAIL.n239 VTAIL.n238 185
R14 VTAIL.n208 VTAIL.n207 185
R15 VTAIL.n245 VTAIL.n244 185
R16 VTAIL.n247 VTAIL.n246 185
R17 VTAIL.n204 VTAIL.n203 185
R18 VTAIL.n253 VTAIL.n252 185
R19 VTAIL.n255 VTAIL.n254 185
R20 VTAIL.n200 VTAIL.n199 185
R21 VTAIL.n261 VTAIL.n260 185
R22 VTAIL.n23 VTAIL.n22 185
R23 VTAIL.n25 VTAIL.n24 185
R24 VTAIL.n18 VTAIL.n17 185
R25 VTAIL.n31 VTAIL.n30 185
R26 VTAIL.n33 VTAIL.n32 185
R27 VTAIL.n14 VTAIL.n13 185
R28 VTAIL.n39 VTAIL.n38 185
R29 VTAIL.n41 VTAIL.n40 185
R30 VTAIL.n10 VTAIL.n9 185
R31 VTAIL.n47 VTAIL.n46 185
R32 VTAIL.n49 VTAIL.n48 185
R33 VTAIL.n6 VTAIL.n5 185
R34 VTAIL.n55 VTAIL.n54 185
R35 VTAIL.n57 VTAIL.n56 185
R36 VTAIL.n2 VTAIL.n1 185
R37 VTAIL.n63 VTAIL.n62 185
R38 VTAIL.n195 VTAIL.n194 185
R39 VTAIL.n134 VTAIL.n133 185
R40 VTAIL.n189 VTAIL.n188 185
R41 VTAIL.n187 VTAIL.n186 185
R42 VTAIL.n138 VTAIL.n137 185
R43 VTAIL.n181 VTAIL.n180 185
R44 VTAIL.n179 VTAIL.n178 185
R45 VTAIL.n142 VTAIL.n141 185
R46 VTAIL.n173 VTAIL.n172 185
R47 VTAIL.n171 VTAIL.n170 185
R48 VTAIL.n146 VTAIL.n145 185
R49 VTAIL.n165 VTAIL.n164 185
R50 VTAIL.n163 VTAIL.n162 185
R51 VTAIL.n150 VTAIL.n149 185
R52 VTAIL.n157 VTAIL.n156 185
R53 VTAIL.n155 VTAIL.n154 185
R54 VTAIL.n129 VTAIL.n128 185
R55 VTAIL.n68 VTAIL.n67 185
R56 VTAIL.n123 VTAIL.n122 185
R57 VTAIL.n121 VTAIL.n120 185
R58 VTAIL.n72 VTAIL.n71 185
R59 VTAIL.n115 VTAIL.n114 185
R60 VTAIL.n113 VTAIL.n112 185
R61 VTAIL.n76 VTAIL.n75 185
R62 VTAIL.n107 VTAIL.n106 185
R63 VTAIL.n105 VTAIL.n104 185
R64 VTAIL.n80 VTAIL.n79 185
R65 VTAIL.n99 VTAIL.n98 185
R66 VTAIL.n97 VTAIL.n96 185
R67 VTAIL.n84 VTAIL.n83 185
R68 VTAIL.n91 VTAIL.n90 185
R69 VTAIL.n89 VTAIL.n88 185
R70 VTAIL.n87 VTAIL.t3 147.659
R71 VTAIL.n219 VTAIL.t2 147.659
R72 VTAIL.n21 VTAIL.t0 147.659
R73 VTAIL.n153 VTAIL.t1 147.659
R74 VTAIL.n222 VTAIL.n221 104.615
R75 VTAIL.n222 VTAIL.n215 104.615
R76 VTAIL.n229 VTAIL.n215 104.615
R77 VTAIL.n230 VTAIL.n229 104.615
R78 VTAIL.n230 VTAIL.n211 104.615
R79 VTAIL.n237 VTAIL.n211 104.615
R80 VTAIL.n238 VTAIL.n237 104.615
R81 VTAIL.n238 VTAIL.n207 104.615
R82 VTAIL.n245 VTAIL.n207 104.615
R83 VTAIL.n246 VTAIL.n245 104.615
R84 VTAIL.n246 VTAIL.n203 104.615
R85 VTAIL.n253 VTAIL.n203 104.615
R86 VTAIL.n254 VTAIL.n253 104.615
R87 VTAIL.n254 VTAIL.n199 104.615
R88 VTAIL.n261 VTAIL.n199 104.615
R89 VTAIL.n24 VTAIL.n23 104.615
R90 VTAIL.n24 VTAIL.n17 104.615
R91 VTAIL.n31 VTAIL.n17 104.615
R92 VTAIL.n32 VTAIL.n31 104.615
R93 VTAIL.n32 VTAIL.n13 104.615
R94 VTAIL.n39 VTAIL.n13 104.615
R95 VTAIL.n40 VTAIL.n39 104.615
R96 VTAIL.n40 VTAIL.n9 104.615
R97 VTAIL.n47 VTAIL.n9 104.615
R98 VTAIL.n48 VTAIL.n47 104.615
R99 VTAIL.n48 VTAIL.n5 104.615
R100 VTAIL.n55 VTAIL.n5 104.615
R101 VTAIL.n56 VTAIL.n55 104.615
R102 VTAIL.n56 VTAIL.n1 104.615
R103 VTAIL.n63 VTAIL.n1 104.615
R104 VTAIL.n195 VTAIL.n133 104.615
R105 VTAIL.n188 VTAIL.n133 104.615
R106 VTAIL.n188 VTAIL.n187 104.615
R107 VTAIL.n187 VTAIL.n137 104.615
R108 VTAIL.n180 VTAIL.n137 104.615
R109 VTAIL.n180 VTAIL.n179 104.615
R110 VTAIL.n179 VTAIL.n141 104.615
R111 VTAIL.n172 VTAIL.n141 104.615
R112 VTAIL.n172 VTAIL.n171 104.615
R113 VTAIL.n171 VTAIL.n145 104.615
R114 VTAIL.n164 VTAIL.n145 104.615
R115 VTAIL.n164 VTAIL.n163 104.615
R116 VTAIL.n163 VTAIL.n149 104.615
R117 VTAIL.n156 VTAIL.n149 104.615
R118 VTAIL.n156 VTAIL.n155 104.615
R119 VTAIL.n129 VTAIL.n67 104.615
R120 VTAIL.n122 VTAIL.n67 104.615
R121 VTAIL.n122 VTAIL.n121 104.615
R122 VTAIL.n121 VTAIL.n71 104.615
R123 VTAIL.n114 VTAIL.n71 104.615
R124 VTAIL.n114 VTAIL.n113 104.615
R125 VTAIL.n113 VTAIL.n75 104.615
R126 VTAIL.n106 VTAIL.n75 104.615
R127 VTAIL.n106 VTAIL.n105 104.615
R128 VTAIL.n105 VTAIL.n79 104.615
R129 VTAIL.n98 VTAIL.n79 104.615
R130 VTAIL.n98 VTAIL.n97 104.615
R131 VTAIL.n97 VTAIL.n83 104.615
R132 VTAIL.n90 VTAIL.n83 104.615
R133 VTAIL.n90 VTAIL.n89 104.615
R134 VTAIL.n221 VTAIL.t2 52.3082
R135 VTAIL.n23 VTAIL.t0 52.3082
R136 VTAIL.n155 VTAIL.t1 52.3082
R137 VTAIL.n89 VTAIL.t3 52.3082
R138 VTAIL.n263 VTAIL.n262 33.7369
R139 VTAIL.n65 VTAIL.n64 33.7369
R140 VTAIL.n197 VTAIL.n196 33.7369
R141 VTAIL.n131 VTAIL.n130 33.7369
R142 VTAIL.n131 VTAIL.n65 24.8669
R143 VTAIL.n263 VTAIL.n197 23.7548
R144 VTAIL.n220 VTAIL.n219 15.6677
R145 VTAIL.n22 VTAIL.n21 15.6677
R146 VTAIL.n154 VTAIL.n153 15.6677
R147 VTAIL.n88 VTAIL.n87 15.6677
R148 VTAIL.n223 VTAIL.n218 12.8005
R149 VTAIL.n25 VTAIL.n20 12.8005
R150 VTAIL.n157 VTAIL.n152 12.8005
R151 VTAIL.n91 VTAIL.n86 12.8005
R152 VTAIL.n224 VTAIL.n216 12.0247
R153 VTAIL.n260 VTAIL.n198 12.0247
R154 VTAIL.n26 VTAIL.n18 12.0247
R155 VTAIL.n62 VTAIL.n0 12.0247
R156 VTAIL.n194 VTAIL.n132 12.0247
R157 VTAIL.n158 VTAIL.n150 12.0247
R158 VTAIL.n128 VTAIL.n66 12.0247
R159 VTAIL.n92 VTAIL.n84 12.0247
R160 VTAIL.n228 VTAIL.n227 11.249
R161 VTAIL.n259 VTAIL.n200 11.249
R162 VTAIL.n30 VTAIL.n29 11.249
R163 VTAIL.n61 VTAIL.n2 11.249
R164 VTAIL.n193 VTAIL.n134 11.249
R165 VTAIL.n162 VTAIL.n161 11.249
R166 VTAIL.n127 VTAIL.n68 11.249
R167 VTAIL.n96 VTAIL.n95 11.249
R168 VTAIL.n231 VTAIL.n214 10.4732
R169 VTAIL.n256 VTAIL.n255 10.4732
R170 VTAIL.n33 VTAIL.n16 10.4732
R171 VTAIL.n58 VTAIL.n57 10.4732
R172 VTAIL.n190 VTAIL.n189 10.4732
R173 VTAIL.n165 VTAIL.n148 10.4732
R174 VTAIL.n124 VTAIL.n123 10.4732
R175 VTAIL.n99 VTAIL.n82 10.4732
R176 VTAIL.n232 VTAIL.n212 9.69747
R177 VTAIL.n252 VTAIL.n202 9.69747
R178 VTAIL.n34 VTAIL.n14 9.69747
R179 VTAIL.n54 VTAIL.n4 9.69747
R180 VTAIL.n186 VTAIL.n136 9.69747
R181 VTAIL.n166 VTAIL.n146 9.69747
R182 VTAIL.n120 VTAIL.n70 9.69747
R183 VTAIL.n100 VTAIL.n80 9.69747
R184 VTAIL.n258 VTAIL.n198 9.45567
R185 VTAIL.n60 VTAIL.n0 9.45567
R186 VTAIL.n192 VTAIL.n132 9.45567
R187 VTAIL.n126 VTAIL.n66 9.45567
R188 VTAIL.n243 VTAIL.n242 9.3005
R189 VTAIL.n206 VTAIL.n205 9.3005
R190 VTAIL.n249 VTAIL.n248 9.3005
R191 VTAIL.n251 VTAIL.n250 9.3005
R192 VTAIL.n202 VTAIL.n201 9.3005
R193 VTAIL.n257 VTAIL.n256 9.3005
R194 VTAIL.n259 VTAIL.n258 9.3005
R195 VTAIL.n210 VTAIL.n209 9.3005
R196 VTAIL.n235 VTAIL.n234 9.3005
R197 VTAIL.n233 VTAIL.n232 9.3005
R198 VTAIL.n214 VTAIL.n213 9.3005
R199 VTAIL.n227 VTAIL.n226 9.3005
R200 VTAIL.n225 VTAIL.n224 9.3005
R201 VTAIL.n218 VTAIL.n217 9.3005
R202 VTAIL.n241 VTAIL.n240 9.3005
R203 VTAIL.n45 VTAIL.n44 9.3005
R204 VTAIL.n8 VTAIL.n7 9.3005
R205 VTAIL.n51 VTAIL.n50 9.3005
R206 VTAIL.n53 VTAIL.n52 9.3005
R207 VTAIL.n4 VTAIL.n3 9.3005
R208 VTAIL.n59 VTAIL.n58 9.3005
R209 VTAIL.n61 VTAIL.n60 9.3005
R210 VTAIL.n12 VTAIL.n11 9.3005
R211 VTAIL.n37 VTAIL.n36 9.3005
R212 VTAIL.n35 VTAIL.n34 9.3005
R213 VTAIL.n16 VTAIL.n15 9.3005
R214 VTAIL.n29 VTAIL.n28 9.3005
R215 VTAIL.n27 VTAIL.n26 9.3005
R216 VTAIL.n20 VTAIL.n19 9.3005
R217 VTAIL.n43 VTAIL.n42 9.3005
R218 VTAIL.n193 VTAIL.n192 9.3005
R219 VTAIL.n191 VTAIL.n190 9.3005
R220 VTAIL.n136 VTAIL.n135 9.3005
R221 VTAIL.n185 VTAIL.n184 9.3005
R222 VTAIL.n183 VTAIL.n182 9.3005
R223 VTAIL.n140 VTAIL.n139 9.3005
R224 VTAIL.n177 VTAIL.n176 9.3005
R225 VTAIL.n175 VTAIL.n174 9.3005
R226 VTAIL.n144 VTAIL.n143 9.3005
R227 VTAIL.n169 VTAIL.n168 9.3005
R228 VTAIL.n167 VTAIL.n166 9.3005
R229 VTAIL.n148 VTAIL.n147 9.3005
R230 VTAIL.n161 VTAIL.n160 9.3005
R231 VTAIL.n159 VTAIL.n158 9.3005
R232 VTAIL.n152 VTAIL.n151 9.3005
R233 VTAIL.n74 VTAIL.n73 9.3005
R234 VTAIL.n117 VTAIL.n116 9.3005
R235 VTAIL.n119 VTAIL.n118 9.3005
R236 VTAIL.n70 VTAIL.n69 9.3005
R237 VTAIL.n125 VTAIL.n124 9.3005
R238 VTAIL.n127 VTAIL.n126 9.3005
R239 VTAIL.n111 VTAIL.n110 9.3005
R240 VTAIL.n109 VTAIL.n108 9.3005
R241 VTAIL.n78 VTAIL.n77 9.3005
R242 VTAIL.n103 VTAIL.n102 9.3005
R243 VTAIL.n101 VTAIL.n100 9.3005
R244 VTAIL.n82 VTAIL.n81 9.3005
R245 VTAIL.n95 VTAIL.n94 9.3005
R246 VTAIL.n93 VTAIL.n92 9.3005
R247 VTAIL.n86 VTAIL.n85 9.3005
R248 VTAIL.n236 VTAIL.n235 8.92171
R249 VTAIL.n251 VTAIL.n204 8.92171
R250 VTAIL.n38 VTAIL.n37 8.92171
R251 VTAIL.n53 VTAIL.n6 8.92171
R252 VTAIL.n185 VTAIL.n138 8.92171
R253 VTAIL.n170 VTAIL.n169 8.92171
R254 VTAIL.n119 VTAIL.n72 8.92171
R255 VTAIL.n104 VTAIL.n103 8.92171
R256 VTAIL.n239 VTAIL.n210 8.14595
R257 VTAIL.n248 VTAIL.n247 8.14595
R258 VTAIL.n41 VTAIL.n12 8.14595
R259 VTAIL.n50 VTAIL.n49 8.14595
R260 VTAIL.n182 VTAIL.n181 8.14595
R261 VTAIL.n173 VTAIL.n144 8.14595
R262 VTAIL.n116 VTAIL.n115 8.14595
R263 VTAIL.n107 VTAIL.n78 8.14595
R264 VTAIL.n240 VTAIL.n208 7.3702
R265 VTAIL.n244 VTAIL.n206 7.3702
R266 VTAIL.n42 VTAIL.n10 7.3702
R267 VTAIL.n46 VTAIL.n8 7.3702
R268 VTAIL.n178 VTAIL.n140 7.3702
R269 VTAIL.n174 VTAIL.n142 7.3702
R270 VTAIL.n112 VTAIL.n74 7.3702
R271 VTAIL.n108 VTAIL.n76 7.3702
R272 VTAIL.n243 VTAIL.n208 6.59444
R273 VTAIL.n244 VTAIL.n243 6.59444
R274 VTAIL.n45 VTAIL.n10 6.59444
R275 VTAIL.n46 VTAIL.n45 6.59444
R276 VTAIL.n178 VTAIL.n177 6.59444
R277 VTAIL.n177 VTAIL.n142 6.59444
R278 VTAIL.n112 VTAIL.n111 6.59444
R279 VTAIL.n111 VTAIL.n76 6.59444
R280 VTAIL.n240 VTAIL.n239 5.81868
R281 VTAIL.n247 VTAIL.n206 5.81868
R282 VTAIL.n42 VTAIL.n41 5.81868
R283 VTAIL.n49 VTAIL.n8 5.81868
R284 VTAIL.n181 VTAIL.n140 5.81868
R285 VTAIL.n174 VTAIL.n173 5.81868
R286 VTAIL.n115 VTAIL.n74 5.81868
R287 VTAIL.n108 VTAIL.n107 5.81868
R288 VTAIL.n236 VTAIL.n210 5.04292
R289 VTAIL.n248 VTAIL.n204 5.04292
R290 VTAIL.n38 VTAIL.n12 5.04292
R291 VTAIL.n50 VTAIL.n6 5.04292
R292 VTAIL.n182 VTAIL.n138 5.04292
R293 VTAIL.n170 VTAIL.n144 5.04292
R294 VTAIL.n116 VTAIL.n72 5.04292
R295 VTAIL.n104 VTAIL.n78 5.04292
R296 VTAIL.n87 VTAIL.n85 4.38563
R297 VTAIL.n219 VTAIL.n217 4.38563
R298 VTAIL.n21 VTAIL.n19 4.38563
R299 VTAIL.n153 VTAIL.n151 4.38563
R300 VTAIL.n235 VTAIL.n212 4.26717
R301 VTAIL.n252 VTAIL.n251 4.26717
R302 VTAIL.n37 VTAIL.n14 4.26717
R303 VTAIL.n54 VTAIL.n53 4.26717
R304 VTAIL.n186 VTAIL.n185 4.26717
R305 VTAIL.n169 VTAIL.n146 4.26717
R306 VTAIL.n120 VTAIL.n119 4.26717
R307 VTAIL.n103 VTAIL.n80 4.26717
R308 VTAIL.n232 VTAIL.n231 3.49141
R309 VTAIL.n255 VTAIL.n202 3.49141
R310 VTAIL.n34 VTAIL.n33 3.49141
R311 VTAIL.n57 VTAIL.n4 3.49141
R312 VTAIL.n189 VTAIL.n136 3.49141
R313 VTAIL.n166 VTAIL.n165 3.49141
R314 VTAIL.n123 VTAIL.n70 3.49141
R315 VTAIL.n100 VTAIL.n99 3.49141
R316 VTAIL.n228 VTAIL.n214 2.71565
R317 VTAIL.n256 VTAIL.n200 2.71565
R318 VTAIL.n30 VTAIL.n16 2.71565
R319 VTAIL.n58 VTAIL.n2 2.71565
R320 VTAIL.n190 VTAIL.n134 2.71565
R321 VTAIL.n162 VTAIL.n148 2.71565
R322 VTAIL.n124 VTAIL.n68 2.71565
R323 VTAIL.n96 VTAIL.n82 2.71565
R324 VTAIL.n227 VTAIL.n216 1.93989
R325 VTAIL.n260 VTAIL.n259 1.93989
R326 VTAIL.n29 VTAIL.n18 1.93989
R327 VTAIL.n62 VTAIL.n61 1.93989
R328 VTAIL.n194 VTAIL.n193 1.93989
R329 VTAIL.n161 VTAIL.n150 1.93989
R330 VTAIL.n128 VTAIL.n127 1.93989
R331 VTAIL.n95 VTAIL.n84 1.93989
R332 VTAIL.n224 VTAIL.n223 1.16414
R333 VTAIL.n262 VTAIL.n198 1.16414
R334 VTAIL.n26 VTAIL.n25 1.16414
R335 VTAIL.n64 VTAIL.n0 1.16414
R336 VTAIL.n196 VTAIL.n132 1.16414
R337 VTAIL.n158 VTAIL.n157 1.16414
R338 VTAIL.n130 VTAIL.n66 1.16414
R339 VTAIL.n92 VTAIL.n91 1.16414
R340 VTAIL.n197 VTAIL.n131 1.02636
R341 VTAIL VTAIL.n65 0.806535
R342 VTAIL.n220 VTAIL.n218 0.388379
R343 VTAIL.n22 VTAIL.n20 0.388379
R344 VTAIL.n154 VTAIL.n152 0.388379
R345 VTAIL.n88 VTAIL.n86 0.388379
R346 VTAIL VTAIL.n263 0.220328
R347 VTAIL.n225 VTAIL.n217 0.155672
R348 VTAIL.n226 VTAIL.n225 0.155672
R349 VTAIL.n226 VTAIL.n213 0.155672
R350 VTAIL.n233 VTAIL.n213 0.155672
R351 VTAIL.n234 VTAIL.n233 0.155672
R352 VTAIL.n234 VTAIL.n209 0.155672
R353 VTAIL.n241 VTAIL.n209 0.155672
R354 VTAIL.n242 VTAIL.n241 0.155672
R355 VTAIL.n242 VTAIL.n205 0.155672
R356 VTAIL.n249 VTAIL.n205 0.155672
R357 VTAIL.n250 VTAIL.n249 0.155672
R358 VTAIL.n250 VTAIL.n201 0.155672
R359 VTAIL.n257 VTAIL.n201 0.155672
R360 VTAIL.n258 VTAIL.n257 0.155672
R361 VTAIL.n27 VTAIL.n19 0.155672
R362 VTAIL.n28 VTAIL.n27 0.155672
R363 VTAIL.n28 VTAIL.n15 0.155672
R364 VTAIL.n35 VTAIL.n15 0.155672
R365 VTAIL.n36 VTAIL.n35 0.155672
R366 VTAIL.n36 VTAIL.n11 0.155672
R367 VTAIL.n43 VTAIL.n11 0.155672
R368 VTAIL.n44 VTAIL.n43 0.155672
R369 VTAIL.n44 VTAIL.n7 0.155672
R370 VTAIL.n51 VTAIL.n7 0.155672
R371 VTAIL.n52 VTAIL.n51 0.155672
R372 VTAIL.n52 VTAIL.n3 0.155672
R373 VTAIL.n59 VTAIL.n3 0.155672
R374 VTAIL.n60 VTAIL.n59 0.155672
R375 VTAIL.n192 VTAIL.n191 0.155672
R376 VTAIL.n191 VTAIL.n135 0.155672
R377 VTAIL.n184 VTAIL.n135 0.155672
R378 VTAIL.n184 VTAIL.n183 0.155672
R379 VTAIL.n183 VTAIL.n139 0.155672
R380 VTAIL.n176 VTAIL.n139 0.155672
R381 VTAIL.n176 VTAIL.n175 0.155672
R382 VTAIL.n175 VTAIL.n143 0.155672
R383 VTAIL.n168 VTAIL.n143 0.155672
R384 VTAIL.n168 VTAIL.n167 0.155672
R385 VTAIL.n167 VTAIL.n147 0.155672
R386 VTAIL.n160 VTAIL.n147 0.155672
R387 VTAIL.n160 VTAIL.n159 0.155672
R388 VTAIL.n159 VTAIL.n151 0.155672
R389 VTAIL.n126 VTAIL.n125 0.155672
R390 VTAIL.n125 VTAIL.n69 0.155672
R391 VTAIL.n118 VTAIL.n69 0.155672
R392 VTAIL.n118 VTAIL.n117 0.155672
R393 VTAIL.n117 VTAIL.n73 0.155672
R394 VTAIL.n110 VTAIL.n73 0.155672
R395 VTAIL.n110 VTAIL.n109 0.155672
R396 VTAIL.n109 VTAIL.n77 0.155672
R397 VTAIL.n102 VTAIL.n77 0.155672
R398 VTAIL.n102 VTAIL.n101 0.155672
R399 VTAIL.n101 VTAIL.n81 0.155672
R400 VTAIL.n94 VTAIL.n81 0.155672
R401 VTAIL.n94 VTAIL.n93 0.155672
R402 VTAIL.n93 VTAIL.n85 0.155672
R403 VDD2.n129 VDD2.n128 289.615
R404 VDD2.n64 VDD2.n63 289.615
R405 VDD2.n128 VDD2.n127 185
R406 VDD2.n67 VDD2.n66 185
R407 VDD2.n122 VDD2.n121 185
R408 VDD2.n120 VDD2.n119 185
R409 VDD2.n71 VDD2.n70 185
R410 VDD2.n114 VDD2.n113 185
R411 VDD2.n112 VDD2.n111 185
R412 VDD2.n75 VDD2.n74 185
R413 VDD2.n106 VDD2.n105 185
R414 VDD2.n104 VDD2.n103 185
R415 VDD2.n79 VDD2.n78 185
R416 VDD2.n98 VDD2.n97 185
R417 VDD2.n96 VDD2.n95 185
R418 VDD2.n83 VDD2.n82 185
R419 VDD2.n90 VDD2.n89 185
R420 VDD2.n88 VDD2.n87 185
R421 VDD2.n23 VDD2.n22 185
R422 VDD2.n25 VDD2.n24 185
R423 VDD2.n18 VDD2.n17 185
R424 VDD2.n31 VDD2.n30 185
R425 VDD2.n33 VDD2.n32 185
R426 VDD2.n14 VDD2.n13 185
R427 VDD2.n39 VDD2.n38 185
R428 VDD2.n41 VDD2.n40 185
R429 VDD2.n10 VDD2.n9 185
R430 VDD2.n47 VDD2.n46 185
R431 VDD2.n49 VDD2.n48 185
R432 VDD2.n6 VDD2.n5 185
R433 VDD2.n55 VDD2.n54 185
R434 VDD2.n57 VDD2.n56 185
R435 VDD2.n2 VDD2.n1 185
R436 VDD2.n63 VDD2.n62 185
R437 VDD2.n86 VDD2.t1 147.659
R438 VDD2.n21 VDD2.t0 147.659
R439 VDD2.n128 VDD2.n66 104.615
R440 VDD2.n121 VDD2.n66 104.615
R441 VDD2.n121 VDD2.n120 104.615
R442 VDD2.n120 VDD2.n70 104.615
R443 VDD2.n113 VDD2.n70 104.615
R444 VDD2.n113 VDD2.n112 104.615
R445 VDD2.n112 VDD2.n74 104.615
R446 VDD2.n105 VDD2.n74 104.615
R447 VDD2.n105 VDD2.n104 104.615
R448 VDD2.n104 VDD2.n78 104.615
R449 VDD2.n97 VDD2.n78 104.615
R450 VDD2.n97 VDD2.n96 104.615
R451 VDD2.n96 VDD2.n82 104.615
R452 VDD2.n89 VDD2.n82 104.615
R453 VDD2.n89 VDD2.n88 104.615
R454 VDD2.n24 VDD2.n23 104.615
R455 VDD2.n24 VDD2.n17 104.615
R456 VDD2.n31 VDD2.n17 104.615
R457 VDD2.n32 VDD2.n31 104.615
R458 VDD2.n32 VDD2.n13 104.615
R459 VDD2.n39 VDD2.n13 104.615
R460 VDD2.n40 VDD2.n39 104.615
R461 VDD2.n40 VDD2.n9 104.615
R462 VDD2.n47 VDD2.n9 104.615
R463 VDD2.n48 VDD2.n47 104.615
R464 VDD2.n48 VDD2.n5 104.615
R465 VDD2.n55 VDD2.n5 104.615
R466 VDD2.n56 VDD2.n55 104.615
R467 VDD2.n56 VDD2.n1 104.615
R468 VDD2.n63 VDD2.n1 104.615
R469 VDD2.n130 VDD2.n64 86.5751
R470 VDD2.n88 VDD2.t1 52.3082
R471 VDD2.n23 VDD2.t0 52.3082
R472 VDD2.n130 VDD2.n129 50.4157
R473 VDD2.n87 VDD2.n86 15.6677
R474 VDD2.n22 VDD2.n21 15.6677
R475 VDD2.n90 VDD2.n85 12.8005
R476 VDD2.n25 VDD2.n20 12.8005
R477 VDD2.n127 VDD2.n65 12.0247
R478 VDD2.n91 VDD2.n83 12.0247
R479 VDD2.n26 VDD2.n18 12.0247
R480 VDD2.n62 VDD2.n0 12.0247
R481 VDD2.n126 VDD2.n67 11.249
R482 VDD2.n95 VDD2.n94 11.249
R483 VDD2.n30 VDD2.n29 11.249
R484 VDD2.n61 VDD2.n2 11.249
R485 VDD2.n123 VDD2.n122 10.4732
R486 VDD2.n98 VDD2.n81 10.4732
R487 VDD2.n33 VDD2.n16 10.4732
R488 VDD2.n58 VDD2.n57 10.4732
R489 VDD2.n119 VDD2.n69 9.69747
R490 VDD2.n99 VDD2.n79 9.69747
R491 VDD2.n34 VDD2.n14 9.69747
R492 VDD2.n54 VDD2.n4 9.69747
R493 VDD2.n125 VDD2.n65 9.45567
R494 VDD2.n60 VDD2.n0 9.45567
R495 VDD2.n126 VDD2.n125 9.3005
R496 VDD2.n124 VDD2.n123 9.3005
R497 VDD2.n69 VDD2.n68 9.3005
R498 VDD2.n118 VDD2.n117 9.3005
R499 VDD2.n116 VDD2.n115 9.3005
R500 VDD2.n73 VDD2.n72 9.3005
R501 VDD2.n110 VDD2.n109 9.3005
R502 VDD2.n108 VDD2.n107 9.3005
R503 VDD2.n77 VDD2.n76 9.3005
R504 VDD2.n102 VDD2.n101 9.3005
R505 VDD2.n100 VDD2.n99 9.3005
R506 VDD2.n81 VDD2.n80 9.3005
R507 VDD2.n94 VDD2.n93 9.3005
R508 VDD2.n92 VDD2.n91 9.3005
R509 VDD2.n85 VDD2.n84 9.3005
R510 VDD2.n45 VDD2.n44 9.3005
R511 VDD2.n8 VDD2.n7 9.3005
R512 VDD2.n51 VDD2.n50 9.3005
R513 VDD2.n53 VDD2.n52 9.3005
R514 VDD2.n4 VDD2.n3 9.3005
R515 VDD2.n59 VDD2.n58 9.3005
R516 VDD2.n61 VDD2.n60 9.3005
R517 VDD2.n12 VDD2.n11 9.3005
R518 VDD2.n37 VDD2.n36 9.3005
R519 VDD2.n35 VDD2.n34 9.3005
R520 VDD2.n16 VDD2.n15 9.3005
R521 VDD2.n29 VDD2.n28 9.3005
R522 VDD2.n27 VDD2.n26 9.3005
R523 VDD2.n20 VDD2.n19 9.3005
R524 VDD2.n43 VDD2.n42 9.3005
R525 VDD2.n118 VDD2.n71 8.92171
R526 VDD2.n103 VDD2.n102 8.92171
R527 VDD2.n38 VDD2.n37 8.92171
R528 VDD2.n53 VDD2.n6 8.92171
R529 VDD2.n115 VDD2.n114 8.14595
R530 VDD2.n106 VDD2.n77 8.14595
R531 VDD2.n41 VDD2.n12 8.14595
R532 VDD2.n50 VDD2.n49 8.14595
R533 VDD2.n111 VDD2.n73 7.3702
R534 VDD2.n107 VDD2.n75 7.3702
R535 VDD2.n42 VDD2.n10 7.3702
R536 VDD2.n46 VDD2.n8 7.3702
R537 VDD2.n111 VDD2.n110 6.59444
R538 VDD2.n110 VDD2.n75 6.59444
R539 VDD2.n45 VDD2.n10 6.59444
R540 VDD2.n46 VDD2.n45 6.59444
R541 VDD2.n114 VDD2.n73 5.81868
R542 VDD2.n107 VDD2.n106 5.81868
R543 VDD2.n42 VDD2.n41 5.81868
R544 VDD2.n49 VDD2.n8 5.81868
R545 VDD2.n115 VDD2.n71 5.04292
R546 VDD2.n103 VDD2.n77 5.04292
R547 VDD2.n38 VDD2.n12 5.04292
R548 VDD2.n50 VDD2.n6 5.04292
R549 VDD2.n86 VDD2.n84 4.38563
R550 VDD2.n21 VDD2.n19 4.38563
R551 VDD2.n119 VDD2.n118 4.26717
R552 VDD2.n102 VDD2.n79 4.26717
R553 VDD2.n37 VDD2.n14 4.26717
R554 VDD2.n54 VDD2.n53 4.26717
R555 VDD2.n122 VDD2.n69 3.49141
R556 VDD2.n99 VDD2.n98 3.49141
R557 VDD2.n34 VDD2.n33 3.49141
R558 VDD2.n57 VDD2.n4 3.49141
R559 VDD2.n123 VDD2.n67 2.71565
R560 VDD2.n95 VDD2.n81 2.71565
R561 VDD2.n30 VDD2.n16 2.71565
R562 VDD2.n58 VDD2.n2 2.71565
R563 VDD2.n127 VDD2.n126 1.93989
R564 VDD2.n94 VDD2.n83 1.93989
R565 VDD2.n29 VDD2.n18 1.93989
R566 VDD2.n62 VDD2.n61 1.93989
R567 VDD2.n129 VDD2.n65 1.16414
R568 VDD2.n91 VDD2.n90 1.16414
R569 VDD2.n26 VDD2.n25 1.16414
R570 VDD2.n64 VDD2.n0 1.16414
R571 VDD2.n87 VDD2.n85 0.388379
R572 VDD2.n22 VDD2.n20 0.388379
R573 VDD2 VDD2.n130 0.336707
R574 VDD2.n125 VDD2.n124 0.155672
R575 VDD2.n124 VDD2.n68 0.155672
R576 VDD2.n117 VDD2.n68 0.155672
R577 VDD2.n117 VDD2.n116 0.155672
R578 VDD2.n116 VDD2.n72 0.155672
R579 VDD2.n109 VDD2.n72 0.155672
R580 VDD2.n109 VDD2.n108 0.155672
R581 VDD2.n108 VDD2.n76 0.155672
R582 VDD2.n101 VDD2.n76 0.155672
R583 VDD2.n101 VDD2.n100 0.155672
R584 VDD2.n100 VDD2.n80 0.155672
R585 VDD2.n93 VDD2.n80 0.155672
R586 VDD2.n93 VDD2.n92 0.155672
R587 VDD2.n92 VDD2.n84 0.155672
R588 VDD2.n27 VDD2.n19 0.155672
R589 VDD2.n28 VDD2.n27 0.155672
R590 VDD2.n28 VDD2.n15 0.155672
R591 VDD2.n35 VDD2.n15 0.155672
R592 VDD2.n36 VDD2.n35 0.155672
R593 VDD2.n36 VDD2.n11 0.155672
R594 VDD2.n43 VDD2.n11 0.155672
R595 VDD2.n44 VDD2.n43 0.155672
R596 VDD2.n44 VDD2.n7 0.155672
R597 VDD2.n51 VDD2.n7 0.155672
R598 VDD2.n52 VDD2.n51 0.155672
R599 VDD2.n52 VDD2.n3 0.155672
R600 VDD2.n59 VDD2.n3 0.155672
R601 VDD2.n60 VDD2.n59 0.155672
R602 B.n590 B.n589 585
R603 B.n261 B.n77 585
R604 B.n260 B.n259 585
R605 B.n258 B.n257 585
R606 B.n256 B.n255 585
R607 B.n254 B.n253 585
R608 B.n252 B.n251 585
R609 B.n250 B.n249 585
R610 B.n248 B.n247 585
R611 B.n246 B.n245 585
R612 B.n244 B.n243 585
R613 B.n242 B.n241 585
R614 B.n240 B.n239 585
R615 B.n238 B.n237 585
R616 B.n236 B.n235 585
R617 B.n234 B.n233 585
R618 B.n232 B.n231 585
R619 B.n230 B.n229 585
R620 B.n228 B.n227 585
R621 B.n226 B.n225 585
R622 B.n224 B.n223 585
R623 B.n222 B.n221 585
R624 B.n220 B.n219 585
R625 B.n218 B.n217 585
R626 B.n216 B.n215 585
R627 B.n214 B.n213 585
R628 B.n212 B.n211 585
R629 B.n210 B.n209 585
R630 B.n208 B.n207 585
R631 B.n206 B.n205 585
R632 B.n204 B.n203 585
R633 B.n202 B.n201 585
R634 B.n200 B.n199 585
R635 B.n198 B.n197 585
R636 B.n196 B.n195 585
R637 B.n194 B.n193 585
R638 B.n192 B.n191 585
R639 B.n190 B.n189 585
R640 B.n188 B.n187 585
R641 B.n186 B.n185 585
R642 B.n184 B.n183 585
R643 B.n181 B.n180 585
R644 B.n179 B.n178 585
R645 B.n177 B.n176 585
R646 B.n175 B.n174 585
R647 B.n173 B.n172 585
R648 B.n171 B.n170 585
R649 B.n169 B.n168 585
R650 B.n167 B.n166 585
R651 B.n165 B.n164 585
R652 B.n163 B.n162 585
R653 B.n160 B.n159 585
R654 B.n158 B.n157 585
R655 B.n156 B.n155 585
R656 B.n154 B.n153 585
R657 B.n152 B.n151 585
R658 B.n150 B.n149 585
R659 B.n148 B.n147 585
R660 B.n146 B.n145 585
R661 B.n144 B.n143 585
R662 B.n142 B.n141 585
R663 B.n140 B.n139 585
R664 B.n138 B.n137 585
R665 B.n136 B.n135 585
R666 B.n134 B.n133 585
R667 B.n132 B.n131 585
R668 B.n130 B.n129 585
R669 B.n128 B.n127 585
R670 B.n126 B.n125 585
R671 B.n124 B.n123 585
R672 B.n122 B.n121 585
R673 B.n120 B.n119 585
R674 B.n118 B.n117 585
R675 B.n116 B.n115 585
R676 B.n114 B.n113 585
R677 B.n112 B.n111 585
R678 B.n110 B.n109 585
R679 B.n108 B.n107 585
R680 B.n106 B.n105 585
R681 B.n104 B.n103 585
R682 B.n102 B.n101 585
R683 B.n100 B.n99 585
R684 B.n98 B.n97 585
R685 B.n96 B.n95 585
R686 B.n94 B.n93 585
R687 B.n92 B.n91 585
R688 B.n90 B.n89 585
R689 B.n88 B.n87 585
R690 B.n86 B.n85 585
R691 B.n84 B.n83 585
R692 B.n32 B.n31 585
R693 B.n595 B.n594 585
R694 B.n588 B.n78 585
R695 B.n78 B.n29 585
R696 B.n587 B.n28 585
R697 B.n599 B.n28 585
R698 B.n586 B.n27 585
R699 B.n600 B.n27 585
R700 B.n585 B.n26 585
R701 B.n601 B.n26 585
R702 B.n584 B.n583 585
R703 B.n583 B.n22 585
R704 B.n582 B.n21 585
R705 B.t10 B.n21 585
R706 B.n581 B.n20 585
R707 B.n607 B.n20 585
R708 B.n580 B.n19 585
R709 B.n608 B.n19 585
R710 B.n579 B.n578 585
R711 B.n578 B.n15 585
R712 B.n577 B.n14 585
R713 B.n614 B.n14 585
R714 B.n576 B.n13 585
R715 B.n615 B.n13 585
R716 B.n575 B.n12 585
R717 B.n616 B.n12 585
R718 B.n574 B.n573 585
R719 B.n573 B.t1 585
R720 B.n572 B.n571 585
R721 B.n572 B.n8 585
R722 B.n570 B.n7 585
R723 B.n623 B.n7 585
R724 B.n569 B.n6 585
R725 B.n624 B.n6 585
R726 B.n568 B.n5 585
R727 B.n625 B.n5 585
R728 B.n567 B.n566 585
R729 B.n566 B.n4 585
R730 B.n565 B.n262 585
R731 B.n565 B.n564 585
R732 B.n555 B.n263 585
R733 B.t0 B.n263 585
R734 B.n557 B.n556 585
R735 B.n558 B.n557 585
R736 B.n554 B.n268 585
R737 B.n268 B.n267 585
R738 B.n553 B.n552 585
R739 B.n552 B.n551 585
R740 B.n270 B.n269 585
R741 B.n271 B.n270 585
R742 B.n544 B.n543 585
R743 B.n545 B.n544 585
R744 B.n542 B.n276 585
R745 B.n276 B.n275 585
R746 B.n541 B.n540 585
R747 B.n540 B.t3 585
R748 B.n278 B.n277 585
R749 B.n279 B.n278 585
R750 B.n533 B.n532 585
R751 B.n534 B.n533 585
R752 B.n531 B.n284 585
R753 B.n284 B.n283 585
R754 B.n530 B.n529 585
R755 B.n529 B.n528 585
R756 B.n286 B.n285 585
R757 B.n287 B.n286 585
R758 B.n524 B.n523 585
R759 B.n290 B.n289 585
R760 B.n520 B.n519 585
R761 B.n521 B.n520 585
R762 B.n518 B.n336 585
R763 B.n517 B.n516 585
R764 B.n515 B.n514 585
R765 B.n513 B.n512 585
R766 B.n511 B.n510 585
R767 B.n509 B.n508 585
R768 B.n507 B.n506 585
R769 B.n505 B.n504 585
R770 B.n503 B.n502 585
R771 B.n501 B.n500 585
R772 B.n499 B.n498 585
R773 B.n497 B.n496 585
R774 B.n495 B.n494 585
R775 B.n493 B.n492 585
R776 B.n491 B.n490 585
R777 B.n489 B.n488 585
R778 B.n487 B.n486 585
R779 B.n485 B.n484 585
R780 B.n483 B.n482 585
R781 B.n481 B.n480 585
R782 B.n479 B.n478 585
R783 B.n477 B.n476 585
R784 B.n475 B.n474 585
R785 B.n473 B.n472 585
R786 B.n471 B.n470 585
R787 B.n469 B.n468 585
R788 B.n467 B.n466 585
R789 B.n465 B.n464 585
R790 B.n463 B.n462 585
R791 B.n461 B.n460 585
R792 B.n459 B.n458 585
R793 B.n457 B.n456 585
R794 B.n455 B.n454 585
R795 B.n453 B.n452 585
R796 B.n451 B.n450 585
R797 B.n449 B.n448 585
R798 B.n447 B.n446 585
R799 B.n445 B.n444 585
R800 B.n443 B.n442 585
R801 B.n441 B.n440 585
R802 B.n439 B.n438 585
R803 B.n437 B.n436 585
R804 B.n435 B.n434 585
R805 B.n433 B.n432 585
R806 B.n431 B.n430 585
R807 B.n429 B.n428 585
R808 B.n427 B.n426 585
R809 B.n425 B.n424 585
R810 B.n423 B.n422 585
R811 B.n421 B.n420 585
R812 B.n419 B.n418 585
R813 B.n417 B.n416 585
R814 B.n415 B.n414 585
R815 B.n413 B.n412 585
R816 B.n411 B.n410 585
R817 B.n409 B.n408 585
R818 B.n407 B.n406 585
R819 B.n405 B.n404 585
R820 B.n403 B.n402 585
R821 B.n401 B.n400 585
R822 B.n399 B.n398 585
R823 B.n397 B.n396 585
R824 B.n395 B.n394 585
R825 B.n393 B.n392 585
R826 B.n391 B.n390 585
R827 B.n389 B.n388 585
R828 B.n387 B.n386 585
R829 B.n385 B.n384 585
R830 B.n383 B.n382 585
R831 B.n381 B.n380 585
R832 B.n379 B.n378 585
R833 B.n377 B.n376 585
R834 B.n375 B.n374 585
R835 B.n373 B.n372 585
R836 B.n371 B.n370 585
R837 B.n369 B.n368 585
R838 B.n367 B.n366 585
R839 B.n365 B.n364 585
R840 B.n363 B.n362 585
R841 B.n361 B.n360 585
R842 B.n359 B.n358 585
R843 B.n357 B.n356 585
R844 B.n355 B.n354 585
R845 B.n353 B.n352 585
R846 B.n351 B.n350 585
R847 B.n349 B.n348 585
R848 B.n347 B.n346 585
R849 B.n345 B.n344 585
R850 B.n343 B.n335 585
R851 B.n521 B.n335 585
R852 B.n525 B.n288 585
R853 B.n288 B.n287 585
R854 B.n527 B.n526 585
R855 B.n528 B.n527 585
R856 B.n282 B.n281 585
R857 B.n283 B.n282 585
R858 B.n536 B.n535 585
R859 B.n535 B.n534 585
R860 B.n537 B.n280 585
R861 B.n280 B.n279 585
R862 B.n539 B.n538 585
R863 B.t3 B.n539 585
R864 B.n274 B.n273 585
R865 B.n275 B.n274 585
R866 B.n547 B.n546 585
R867 B.n546 B.n545 585
R868 B.n548 B.n272 585
R869 B.n272 B.n271 585
R870 B.n550 B.n549 585
R871 B.n551 B.n550 585
R872 B.n266 B.n265 585
R873 B.n267 B.n266 585
R874 B.n560 B.n559 585
R875 B.n559 B.n558 585
R876 B.n561 B.n264 585
R877 B.n264 B.t0 585
R878 B.n563 B.n562 585
R879 B.n564 B.n563 585
R880 B.n3 B.n0 585
R881 B.n4 B.n3 585
R882 B.n622 B.n1 585
R883 B.n623 B.n622 585
R884 B.n621 B.n620 585
R885 B.n621 B.n8 585
R886 B.n619 B.n9 585
R887 B.t1 B.n9 585
R888 B.n618 B.n617 585
R889 B.n617 B.n616 585
R890 B.n11 B.n10 585
R891 B.n615 B.n11 585
R892 B.n613 B.n612 585
R893 B.n614 B.n613 585
R894 B.n611 B.n16 585
R895 B.n16 B.n15 585
R896 B.n610 B.n609 585
R897 B.n609 B.n608 585
R898 B.n18 B.n17 585
R899 B.n607 B.n18 585
R900 B.n606 B.n605 585
R901 B.t10 B.n606 585
R902 B.n604 B.n23 585
R903 B.n23 B.n22 585
R904 B.n603 B.n602 585
R905 B.n602 B.n601 585
R906 B.n25 B.n24 585
R907 B.n600 B.n25 585
R908 B.n598 B.n597 585
R909 B.n599 B.n598 585
R910 B.n596 B.n30 585
R911 B.n30 B.n29 585
R912 B.n626 B.n625 585
R913 B.n624 B.n2 585
R914 B.n594 B.n30 559.769
R915 B.n590 B.n78 559.769
R916 B.n335 B.n286 559.769
R917 B.n523 B.n288 559.769
R918 B.n81 B.t13 501.385
R919 B.n79 B.t9 501.385
R920 B.n340 B.t2 501.385
R921 B.n337 B.t6 501.385
R922 B.n79 B.t11 305.087
R923 B.n340 B.t5 305.087
R924 B.n81 B.t14 305.087
R925 B.n337 B.t8 305.087
R926 B.n80 B.t12 280.068
R927 B.n341 B.t4 280.068
R928 B.n82 B.t15 280.068
R929 B.n338 B.t7 280.068
R930 B.n592 B.n591 256.663
R931 B.n592 B.n76 256.663
R932 B.n592 B.n75 256.663
R933 B.n592 B.n74 256.663
R934 B.n592 B.n73 256.663
R935 B.n592 B.n72 256.663
R936 B.n592 B.n71 256.663
R937 B.n592 B.n70 256.663
R938 B.n592 B.n69 256.663
R939 B.n592 B.n68 256.663
R940 B.n592 B.n67 256.663
R941 B.n592 B.n66 256.663
R942 B.n592 B.n65 256.663
R943 B.n592 B.n64 256.663
R944 B.n592 B.n63 256.663
R945 B.n592 B.n62 256.663
R946 B.n592 B.n61 256.663
R947 B.n592 B.n60 256.663
R948 B.n592 B.n59 256.663
R949 B.n592 B.n58 256.663
R950 B.n592 B.n57 256.663
R951 B.n592 B.n56 256.663
R952 B.n592 B.n55 256.663
R953 B.n592 B.n54 256.663
R954 B.n592 B.n53 256.663
R955 B.n592 B.n52 256.663
R956 B.n592 B.n51 256.663
R957 B.n592 B.n50 256.663
R958 B.n592 B.n49 256.663
R959 B.n592 B.n48 256.663
R960 B.n592 B.n47 256.663
R961 B.n592 B.n46 256.663
R962 B.n592 B.n45 256.663
R963 B.n592 B.n44 256.663
R964 B.n592 B.n43 256.663
R965 B.n592 B.n42 256.663
R966 B.n592 B.n41 256.663
R967 B.n592 B.n40 256.663
R968 B.n592 B.n39 256.663
R969 B.n592 B.n38 256.663
R970 B.n592 B.n37 256.663
R971 B.n592 B.n36 256.663
R972 B.n592 B.n35 256.663
R973 B.n592 B.n34 256.663
R974 B.n592 B.n33 256.663
R975 B.n593 B.n592 256.663
R976 B.n522 B.n521 256.663
R977 B.n521 B.n291 256.663
R978 B.n521 B.n292 256.663
R979 B.n521 B.n293 256.663
R980 B.n521 B.n294 256.663
R981 B.n521 B.n295 256.663
R982 B.n521 B.n296 256.663
R983 B.n521 B.n297 256.663
R984 B.n521 B.n298 256.663
R985 B.n521 B.n299 256.663
R986 B.n521 B.n300 256.663
R987 B.n521 B.n301 256.663
R988 B.n521 B.n302 256.663
R989 B.n521 B.n303 256.663
R990 B.n521 B.n304 256.663
R991 B.n521 B.n305 256.663
R992 B.n521 B.n306 256.663
R993 B.n521 B.n307 256.663
R994 B.n521 B.n308 256.663
R995 B.n521 B.n309 256.663
R996 B.n521 B.n310 256.663
R997 B.n521 B.n311 256.663
R998 B.n521 B.n312 256.663
R999 B.n521 B.n313 256.663
R1000 B.n521 B.n314 256.663
R1001 B.n521 B.n315 256.663
R1002 B.n521 B.n316 256.663
R1003 B.n521 B.n317 256.663
R1004 B.n521 B.n318 256.663
R1005 B.n521 B.n319 256.663
R1006 B.n521 B.n320 256.663
R1007 B.n521 B.n321 256.663
R1008 B.n521 B.n322 256.663
R1009 B.n521 B.n323 256.663
R1010 B.n521 B.n324 256.663
R1011 B.n521 B.n325 256.663
R1012 B.n521 B.n326 256.663
R1013 B.n521 B.n327 256.663
R1014 B.n521 B.n328 256.663
R1015 B.n521 B.n329 256.663
R1016 B.n521 B.n330 256.663
R1017 B.n521 B.n331 256.663
R1018 B.n521 B.n332 256.663
R1019 B.n521 B.n333 256.663
R1020 B.n521 B.n334 256.663
R1021 B.n628 B.n627 256.663
R1022 B.n83 B.n32 163.367
R1023 B.n87 B.n86 163.367
R1024 B.n91 B.n90 163.367
R1025 B.n95 B.n94 163.367
R1026 B.n99 B.n98 163.367
R1027 B.n103 B.n102 163.367
R1028 B.n107 B.n106 163.367
R1029 B.n111 B.n110 163.367
R1030 B.n115 B.n114 163.367
R1031 B.n119 B.n118 163.367
R1032 B.n123 B.n122 163.367
R1033 B.n127 B.n126 163.367
R1034 B.n131 B.n130 163.367
R1035 B.n135 B.n134 163.367
R1036 B.n139 B.n138 163.367
R1037 B.n143 B.n142 163.367
R1038 B.n147 B.n146 163.367
R1039 B.n151 B.n150 163.367
R1040 B.n155 B.n154 163.367
R1041 B.n159 B.n158 163.367
R1042 B.n164 B.n163 163.367
R1043 B.n168 B.n167 163.367
R1044 B.n172 B.n171 163.367
R1045 B.n176 B.n175 163.367
R1046 B.n180 B.n179 163.367
R1047 B.n185 B.n184 163.367
R1048 B.n189 B.n188 163.367
R1049 B.n193 B.n192 163.367
R1050 B.n197 B.n196 163.367
R1051 B.n201 B.n200 163.367
R1052 B.n205 B.n204 163.367
R1053 B.n209 B.n208 163.367
R1054 B.n213 B.n212 163.367
R1055 B.n217 B.n216 163.367
R1056 B.n221 B.n220 163.367
R1057 B.n225 B.n224 163.367
R1058 B.n229 B.n228 163.367
R1059 B.n233 B.n232 163.367
R1060 B.n237 B.n236 163.367
R1061 B.n241 B.n240 163.367
R1062 B.n245 B.n244 163.367
R1063 B.n249 B.n248 163.367
R1064 B.n253 B.n252 163.367
R1065 B.n257 B.n256 163.367
R1066 B.n259 B.n77 163.367
R1067 B.n529 B.n286 163.367
R1068 B.n529 B.n284 163.367
R1069 B.n533 B.n284 163.367
R1070 B.n533 B.n278 163.367
R1071 B.n540 B.n278 163.367
R1072 B.n540 B.n276 163.367
R1073 B.n544 B.n276 163.367
R1074 B.n544 B.n270 163.367
R1075 B.n552 B.n270 163.367
R1076 B.n552 B.n268 163.367
R1077 B.n557 B.n268 163.367
R1078 B.n557 B.n263 163.367
R1079 B.n565 B.n263 163.367
R1080 B.n566 B.n565 163.367
R1081 B.n566 B.n5 163.367
R1082 B.n6 B.n5 163.367
R1083 B.n7 B.n6 163.367
R1084 B.n572 B.n7 163.367
R1085 B.n573 B.n572 163.367
R1086 B.n573 B.n12 163.367
R1087 B.n13 B.n12 163.367
R1088 B.n14 B.n13 163.367
R1089 B.n578 B.n14 163.367
R1090 B.n578 B.n19 163.367
R1091 B.n20 B.n19 163.367
R1092 B.n21 B.n20 163.367
R1093 B.n583 B.n21 163.367
R1094 B.n583 B.n26 163.367
R1095 B.n27 B.n26 163.367
R1096 B.n28 B.n27 163.367
R1097 B.n78 B.n28 163.367
R1098 B.n520 B.n290 163.367
R1099 B.n520 B.n336 163.367
R1100 B.n516 B.n515 163.367
R1101 B.n512 B.n511 163.367
R1102 B.n508 B.n507 163.367
R1103 B.n504 B.n503 163.367
R1104 B.n500 B.n499 163.367
R1105 B.n496 B.n495 163.367
R1106 B.n492 B.n491 163.367
R1107 B.n488 B.n487 163.367
R1108 B.n484 B.n483 163.367
R1109 B.n480 B.n479 163.367
R1110 B.n476 B.n475 163.367
R1111 B.n472 B.n471 163.367
R1112 B.n468 B.n467 163.367
R1113 B.n464 B.n463 163.367
R1114 B.n460 B.n459 163.367
R1115 B.n456 B.n455 163.367
R1116 B.n452 B.n451 163.367
R1117 B.n448 B.n447 163.367
R1118 B.n444 B.n443 163.367
R1119 B.n440 B.n439 163.367
R1120 B.n436 B.n435 163.367
R1121 B.n432 B.n431 163.367
R1122 B.n428 B.n427 163.367
R1123 B.n424 B.n423 163.367
R1124 B.n420 B.n419 163.367
R1125 B.n416 B.n415 163.367
R1126 B.n412 B.n411 163.367
R1127 B.n408 B.n407 163.367
R1128 B.n404 B.n403 163.367
R1129 B.n400 B.n399 163.367
R1130 B.n396 B.n395 163.367
R1131 B.n392 B.n391 163.367
R1132 B.n388 B.n387 163.367
R1133 B.n384 B.n383 163.367
R1134 B.n380 B.n379 163.367
R1135 B.n376 B.n375 163.367
R1136 B.n372 B.n371 163.367
R1137 B.n368 B.n367 163.367
R1138 B.n364 B.n363 163.367
R1139 B.n360 B.n359 163.367
R1140 B.n356 B.n355 163.367
R1141 B.n352 B.n351 163.367
R1142 B.n348 B.n347 163.367
R1143 B.n344 B.n335 163.367
R1144 B.n527 B.n288 163.367
R1145 B.n527 B.n282 163.367
R1146 B.n535 B.n282 163.367
R1147 B.n535 B.n280 163.367
R1148 B.n539 B.n280 163.367
R1149 B.n539 B.n274 163.367
R1150 B.n546 B.n274 163.367
R1151 B.n546 B.n272 163.367
R1152 B.n550 B.n272 163.367
R1153 B.n550 B.n266 163.367
R1154 B.n559 B.n266 163.367
R1155 B.n559 B.n264 163.367
R1156 B.n563 B.n264 163.367
R1157 B.n563 B.n3 163.367
R1158 B.n626 B.n3 163.367
R1159 B.n622 B.n2 163.367
R1160 B.n622 B.n621 163.367
R1161 B.n621 B.n9 163.367
R1162 B.n617 B.n9 163.367
R1163 B.n617 B.n11 163.367
R1164 B.n613 B.n11 163.367
R1165 B.n613 B.n16 163.367
R1166 B.n609 B.n16 163.367
R1167 B.n609 B.n18 163.367
R1168 B.n606 B.n18 163.367
R1169 B.n606 B.n23 163.367
R1170 B.n602 B.n23 163.367
R1171 B.n602 B.n25 163.367
R1172 B.n598 B.n25 163.367
R1173 B.n598 B.n30 163.367
R1174 B.n521 B.n287 87.6423
R1175 B.n592 B.n29 87.6423
R1176 B.n594 B.n593 71.676
R1177 B.n83 B.n33 71.676
R1178 B.n87 B.n34 71.676
R1179 B.n91 B.n35 71.676
R1180 B.n95 B.n36 71.676
R1181 B.n99 B.n37 71.676
R1182 B.n103 B.n38 71.676
R1183 B.n107 B.n39 71.676
R1184 B.n111 B.n40 71.676
R1185 B.n115 B.n41 71.676
R1186 B.n119 B.n42 71.676
R1187 B.n123 B.n43 71.676
R1188 B.n127 B.n44 71.676
R1189 B.n131 B.n45 71.676
R1190 B.n135 B.n46 71.676
R1191 B.n139 B.n47 71.676
R1192 B.n143 B.n48 71.676
R1193 B.n147 B.n49 71.676
R1194 B.n151 B.n50 71.676
R1195 B.n155 B.n51 71.676
R1196 B.n159 B.n52 71.676
R1197 B.n164 B.n53 71.676
R1198 B.n168 B.n54 71.676
R1199 B.n172 B.n55 71.676
R1200 B.n176 B.n56 71.676
R1201 B.n180 B.n57 71.676
R1202 B.n185 B.n58 71.676
R1203 B.n189 B.n59 71.676
R1204 B.n193 B.n60 71.676
R1205 B.n197 B.n61 71.676
R1206 B.n201 B.n62 71.676
R1207 B.n205 B.n63 71.676
R1208 B.n209 B.n64 71.676
R1209 B.n213 B.n65 71.676
R1210 B.n217 B.n66 71.676
R1211 B.n221 B.n67 71.676
R1212 B.n225 B.n68 71.676
R1213 B.n229 B.n69 71.676
R1214 B.n233 B.n70 71.676
R1215 B.n237 B.n71 71.676
R1216 B.n241 B.n72 71.676
R1217 B.n245 B.n73 71.676
R1218 B.n249 B.n74 71.676
R1219 B.n253 B.n75 71.676
R1220 B.n257 B.n76 71.676
R1221 B.n591 B.n77 71.676
R1222 B.n591 B.n590 71.676
R1223 B.n259 B.n76 71.676
R1224 B.n256 B.n75 71.676
R1225 B.n252 B.n74 71.676
R1226 B.n248 B.n73 71.676
R1227 B.n244 B.n72 71.676
R1228 B.n240 B.n71 71.676
R1229 B.n236 B.n70 71.676
R1230 B.n232 B.n69 71.676
R1231 B.n228 B.n68 71.676
R1232 B.n224 B.n67 71.676
R1233 B.n220 B.n66 71.676
R1234 B.n216 B.n65 71.676
R1235 B.n212 B.n64 71.676
R1236 B.n208 B.n63 71.676
R1237 B.n204 B.n62 71.676
R1238 B.n200 B.n61 71.676
R1239 B.n196 B.n60 71.676
R1240 B.n192 B.n59 71.676
R1241 B.n188 B.n58 71.676
R1242 B.n184 B.n57 71.676
R1243 B.n179 B.n56 71.676
R1244 B.n175 B.n55 71.676
R1245 B.n171 B.n54 71.676
R1246 B.n167 B.n53 71.676
R1247 B.n163 B.n52 71.676
R1248 B.n158 B.n51 71.676
R1249 B.n154 B.n50 71.676
R1250 B.n150 B.n49 71.676
R1251 B.n146 B.n48 71.676
R1252 B.n142 B.n47 71.676
R1253 B.n138 B.n46 71.676
R1254 B.n134 B.n45 71.676
R1255 B.n130 B.n44 71.676
R1256 B.n126 B.n43 71.676
R1257 B.n122 B.n42 71.676
R1258 B.n118 B.n41 71.676
R1259 B.n114 B.n40 71.676
R1260 B.n110 B.n39 71.676
R1261 B.n106 B.n38 71.676
R1262 B.n102 B.n37 71.676
R1263 B.n98 B.n36 71.676
R1264 B.n94 B.n35 71.676
R1265 B.n90 B.n34 71.676
R1266 B.n86 B.n33 71.676
R1267 B.n593 B.n32 71.676
R1268 B.n523 B.n522 71.676
R1269 B.n336 B.n291 71.676
R1270 B.n515 B.n292 71.676
R1271 B.n511 B.n293 71.676
R1272 B.n507 B.n294 71.676
R1273 B.n503 B.n295 71.676
R1274 B.n499 B.n296 71.676
R1275 B.n495 B.n297 71.676
R1276 B.n491 B.n298 71.676
R1277 B.n487 B.n299 71.676
R1278 B.n483 B.n300 71.676
R1279 B.n479 B.n301 71.676
R1280 B.n475 B.n302 71.676
R1281 B.n471 B.n303 71.676
R1282 B.n467 B.n304 71.676
R1283 B.n463 B.n305 71.676
R1284 B.n459 B.n306 71.676
R1285 B.n455 B.n307 71.676
R1286 B.n451 B.n308 71.676
R1287 B.n447 B.n309 71.676
R1288 B.n443 B.n310 71.676
R1289 B.n439 B.n311 71.676
R1290 B.n435 B.n312 71.676
R1291 B.n431 B.n313 71.676
R1292 B.n427 B.n314 71.676
R1293 B.n423 B.n315 71.676
R1294 B.n419 B.n316 71.676
R1295 B.n415 B.n317 71.676
R1296 B.n411 B.n318 71.676
R1297 B.n407 B.n319 71.676
R1298 B.n403 B.n320 71.676
R1299 B.n399 B.n321 71.676
R1300 B.n395 B.n322 71.676
R1301 B.n391 B.n323 71.676
R1302 B.n387 B.n324 71.676
R1303 B.n383 B.n325 71.676
R1304 B.n379 B.n326 71.676
R1305 B.n375 B.n327 71.676
R1306 B.n371 B.n328 71.676
R1307 B.n367 B.n329 71.676
R1308 B.n363 B.n330 71.676
R1309 B.n359 B.n331 71.676
R1310 B.n355 B.n332 71.676
R1311 B.n351 B.n333 71.676
R1312 B.n347 B.n334 71.676
R1313 B.n522 B.n290 71.676
R1314 B.n516 B.n291 71.676
R1315 B.n512 B.n292 71.676
R1316 B.n508 B.n293 71.676
R1317 B.n504 B.n294 71.676
R1318 B.n500 B.n295 71.676
R1319 B.n496 B.n296 71.676
R1320 B.n492 B.n297 71.676
R1321 B.n488 B.n298 71.676
R1322 B.n484 B.n299 71.676
R1323 B.n480 B.n300 71.676
R1324 B.n476 B.n301 71.676
R1325 B.n472 B.n302 71.676
R1326 B.n468 B.n303 71.676
R1327 B.n464 B.n304 71.676
R1328 B.n460 B.n305 71.676
R1329 B.n456 B.n306 71.676
R1330 B.n452 B.n307 71.676
R1331 B.n448 B.n308 71.676
R1332 B.n444 B.n309 71.676
R1333 B.n440 B.n310 71.676
R1334 B.n436 B.n311 71.676
R1335 B.n432 B.n312 71.676
R1336 B.n428 B.n313 71.676
R1337 B.n424 B.n314 71.676
R1338 B.n420 B.n315 71.676
R1339 B.n416 B.n316 71.676
R1340 B.n412 B.n317 71.676
R1341 B.n408 B.n318 71.676
R1342 B.n404 B.n319 71.676
R1343 B.n400 B.n320 71.676
R1344 B.n396 B.n321 71.676
R1345 B.n392 B.n322 71.676
R1346 B.n388 B.n323 71.676
R1347 B.n384 B.n324 71.676
R1348 B.n380 B.n325 71.676
R1349 B.n376 B.n326 71.676
R1350 B.n372 B.n327 71.676
R1351 B.n368 B.n328 71.676
R1352 B.n364 B.n329 71.676
R1353 B.n360 B.n330 71.676
R1354 B.n356 B.n331 71.676
R1355 B.n352 B.n332 71.676
R1356 B.n348 B.n333 71.676
R1357 B.n344 B.n334 71.676
R1358 B.n627 B.n626 71.676
R1359 B.n627 B.n2 71.676
R1360 B.n161 B.n82 59.5399
R1361 B.n182 B.n80 59.5399
R1362 B.n342 B.n341 59.5399
R1363 B.n339 B.n338 59.5399
R1364 B.n528 B.n287 43.5015
R1365 B.n528 B.n283 43.5015
R1366 B.n534 B.n283 43.5015
R1367 B.n534 B.n279 43.5015
R1368 B.t3 B.n279 43.5015
R1369 B.t3 B.n275 43.5015
R1370 B.n545 B.n275 43.5015
R1371 B.n545 B.n271 43.5015
R1372 B.n551 B.n271 43.5015
R1373 B.n551 B.n267 43.5015
R1374 B.n558 B.n267 43.5015
R1375 B.n558 B.t0 43.5015
R1376 B.n564 B.t0 43.5015
R1377 B.n564 B.n4 43.5015
R1378 B.n625 B.n4 43.5015
R1379 B.n625 B.n624 43.5015
R1380 B.n624 B.n623 43.5015
R1381 B.n623 B.n8 43.5015
R1382 B.t1 B.n8 43.5015
R1383 B.n616 B.t1 43.5015
R1384 B.n616 B.n615 43.5015
R1385 B.n615 B.n614 43.5015
R1386 B.n614 B.n15 43.5015
R1387 B.n608 B.n15 43.5015
R1388 B.n608 B.n607 43.5015
R1389 B.n607 B.t10 43.5015
R1390 B.t10 B.n22 43.5015
R1391 B.n601 B.n22 43.5015
R1392 B.n601 B.n600 43.5015
R1393 B.n600 B.n599 43.5015
R1394 B.n599 B.n29 43.5015
R1395 B.n525 B.n524 36.3712
R1396 B.n343 B.n285 36.3712
R1397 B.n589 B.n588 36.3712
R1398 B.n596 B.n595 36.3712
R1399 B.n82 B.n81 25.0187
R1400 B.n80 B.n79 25.0187
R1401 B.n341 B.n340 25.0187
R1402 B.n338 B.n337 25.0187
R1403 B B.n628 18.0485
R1404 B.n526 B.n525 10.6151
R1405 B.n526 B.n281 10.6151
R1406 B.n536 B.n281 10.6151
R1407 B.n537 B.n536 10.6151
R1408 B.n538 B.n537 10.6151
R1409 B.n538 B.n273 10.6151
R1410 B.n547 B.n273 10.6151
R1411 B.n548 B.n547 10.6151
R1412 B.n549 B.n548 10.6151
R1413 B.n549 B.n265 10.6151
R1414 B.n560 B.n265 10.6151
R1415 B.n561 B.n560 10.6151
R1416 B.n562 B.n561 10.6151
R1417 B.n562 B.n0 10.6151
R1418 B.n524 B.n289 10.6151
R1419 B.n519 B.n289 10.6151
R1420 B.n519 B.n518 10.6151
R1421 B.n518 B.n517 10.6151
R1422 B.n517 B.n514 10.6151
R1423 B.n514 B.n513 10.6151
R1424 B.n513 B.n510 10.6151
R1425 B.n510 B.n509 10.6151
R1426 B.n509 B.n506 10.6151
R1427 B.n506 B.n505 10.6151
R1428 B.n505 B.n502 10.6151
R1429 B.n502 B.n501 10.6151
R1430 B.n501 B.n498 10.6151
R1431 B.n498 B.n497 10.6151
R1432 B.n497 B.n494 10.6151
R1433 B.n494 B.n493 10.6151
R1434 B.n493 B.n490 10.6151
R1435 B.n490 B.n489 10.6151
R1436 B.n489 B.n486 10.6151
R1437 B.n486 B.n485 10.6151
R1438 B.n485 B.n482 10.6151
R1439 B.n482 B.n481 10.6151
R1440 B.n481 B.n478 10.6151
R1441 B.n478 B.n477 10.6151
R1442 B.n477 B.n474 10.6151
R1443 B.n474 B.n473 10.6151
R1444 B.n473 B.n470 10.6151
R1445 B.n470 B.n469 10.6151
R1446 B.n469 B.n466 10.6151
R1447 B.n466 B.n465 10.6151
R1448 B.n465 B.n462 10.6151
R1449 B.n462 B.n461 10.6151
R1450 B.n461 B.n458 10.6151
R1451 B.n458 B.n457 10.6151
R1452 B.n457 B.n454 10.6151
R1453 B.n454 B.n453 10.6151
R1454 B.n453 B.n450 10.6151
R1455 B.n450 B.n449 10.6151
R1456 B.n449 B.n446 10.6151
R1457 B.n446 B.n445 10.6151
R1458 B.n442 B.n441 10.6151
R1459 B.n441 B.n438 10.6151
R1460 B.n438 B.n437 10.6151
R1461 B.n437 B.n434 10.6151
R1462 B.n434 B.n433 10.6151
R1463 B.n433 B.n430 10.6151
R1464 B.n430 B.n429 10.6151
R1465 B.n429 B.n426 10.6151
R1466 B.n426 B.n425 10.6151
R1467 B.n422 B.n421 10.6151
R1468 B.n421 B.n418 10.6151
R1469 B.n418 B.n417 10.6151
R1470 B.n417 B.n414 10.6151
R1471 B.n414 B.n413 10.6151
R1472 B.n413 B.n410 10.6151
R1473 B.n410 B.n409 10.6151
R1474 B.n409 B.n406 10.6151
R1475 B.n406 B.n405 10.6151
R1476 B.n405 B.n402 10.6151
R1477 B.n402 B.n401 10.6151
R1478 B.n401 B.n398 10.6151
R1479 B.n398 B.n397 10.6151
R1480 B.n397 B.n394 10.6151
R1481 B.n394 B.n393 10.6151
R1482 B.n393 B.n390 10.6151
R1483 B.n390 B.n389 10.6151
R1484 B.n389 B.n386 10.6151
R1485 B.n386 B.n385 10.6151
R1486 B.n385 B.n382 10.6151
R1487 B.n382 B.n381 10.6151
R1488 B.n381 B.n378 10.6151
R1489 B.n378 B.n377 10.6151
R1490 B.n377 B.n374 10.6151
R1491 B.n374 B.n373 10.6151
R1492 B.n373 B.n370 10.6151
R1493 B.n370 B.n369 10.6151
R1494 B.n369 B.n366 10.6151
R1495 B.n366 B.n365 10.6151
R1496 B.n365 B.n362 10.6151
R1497 B.n362 B.n361 10.6151
R1498 B.n361 B.n358 10.6151
R1499 B.n358 B.n357 10.6151
R1500 B.n357 B.n354 10.6151
R1501 B.n354 B.n353 10.6151
R1502 B.n353 B.n350 10.6151
R1503 B.n350 B.n349 10.6151
R1504 B.n349 B.n346 10.6151
R1505 B.n346 B.n345 10.6151
R1506 B.n345 B.n343 10.6151
R1507 B.n530 B.n285 10.6151
R1508 B.n531 B.n530 10.6151
R1509 B.n532 B.n531 10.6151
R1510 B.n532 B.n277 10.6151
R1511 B.n541 B.n277 10.6151
R1512 B.n542 B.n541 10.6151
R1513 B.n543 B.n542 10.6151
R1514 B.n543 B.n269 10.6151
R1515 B.n553 B.n269 10.6151
R1516 B.n554 B.n553 10.6151
R1517 B.n556 B.n554 10.6151
R1518 B.n556 B.n555 10.6151
R1519 B.n555 B.n262 10.6151
R1520 B.n567 B.n262 10.6151
R1521 B.n568 B.n567 10.6151
R1522 B.n569 B.n568 10.6151
R1523 B.n570 B.n569 10.6151
R1524 B.n571 B.n570 10.6151
R1525 B.n574 B.n571 10.6151
R1526 B.n575 B.n574 10.6151
R1527 B.n576 B.n575 10.6151
R1528 B.n577 B.n576 10.6151
R1529 B.n579 B.n577 10.6151
R1530 B.n580 B.n579 10.6151
R1531 B.n581 B.n580 10.6151
R1532 B.n582 B.n581 10.6151
R1533 B.n584 B.n582 10.6151
R1534 B.n585 B.n584 10.6151
R1535 B.n586 B.n585 10.6151
R1536 B.n587 B.n586 10.6151
R1537 B.n588 B.n587 10.6151
R1538 B.n620 B.n1 10.6151
R1539 B.n620 B.n619 10.6151
R1540 B.n619 B.n618 10.6151
R1541 B.n618 B.n10 10.6151
R1542 B.n612 B.n10 10.6151
R1543 B.n612 B.n611 10.6151
R1544 B.n611 B.n610 10.6151
R1545 B.n610 B.n17 10.6151
R1546 B.n605 B.n17 10.6151
R1547 B.n605 B.n604 10.6151
R1548 B.n604 B.n603 10.6151
R1549 B.n603 B.n24 10.6151
R1550 B.n597 B.n24 10.6151
R1551 B.n597 B.n596 10.6151
R1552 B.n595 B.n31 10.6151
R1553 B.n84 B.n31 10.6151
R1554 B.n85 B.n84 10.6151
R1555 B.n88 B.n85 10.6151
R1556 B.n89 B.n88 10.6151
R1557 B.n92 B.n89 10.6151
R1558 B.n93 B.n92 10.6151
R1559 B.n96 B.n93 10.6151
R1560 B.n97 B.n96 10.6151
R1561 B.n100 B.n97 10.6151
R1562 B.n101 B.n100 10.6151
R1563 B.n104 B.n101 10.6151
R1564 B.n105 B.n104 10.6151
R1565 B.n108 B.n105 10.6151
R1566 B.n109 B.n108 10.6151
R1567 B.n112 B.n109 10.6151
R1568 B.n113 B.n112 10.6151
R1569 B.n116 B.n113 10.6151
R1570 B.n117 B.n116 10.6151
R1571 B.n120 B.n117 10.6151
R1572 B.n121 B.n120 10.6151
R1573 B.n124 B.n121 10.6151
R1574 B.n125 B.n124 10.6151
R1575 B.n128 B.n125 10.6151
R1576 B.n129 B.n128 10.6151
R1577 B.n132 B.n129 10.6151
R1578 B.n133 B.n132 10.6151
R1579 B.n136 B.n133 10.6151
R1580 B.n137 B.n136 10.6151
R1581 B.n140 B.n137 10.6151
R1582 B.n141 B.n140 10.6151
R1583 B.n144 B.n141 10.6151
R1584 B.n145 B.n144 10.6151
R1585 B.n148 B.n145 10.6151
R1586 B.n149 B.n148 10.6151
R1587 B.n152 B.n149 10.6151
R1588 B.n153 B.n152 10.6151
R1589 B.n156 B.n153 10.6151
R1590 B.n157 B.n156 10.6151
R1591 B.n160 B.n157 10.6151
R1592 B.n165 B.n162 10.6151
R1593 B.n166 B.n165 10.6151
R1594 B.n169 B.n166 10.6151
R1595 B.n170 B.n169 10.6151
R1596 B.n173 B.n170 10.6151
R1597 B.n174 B.n173 10.6151
R1598 B.n177 B.n174 10.6151
R1599 B.n178 B.n177 10.6151
R1600 B.n181 B.n178 10.6151
R1601 B.n186 B.n183 10.6151
R1602 B.n187 B.n186 10.6151
R1603 B.n190 B.n187 10.6151
R1604 B.n191 B.n190 10.6151
R1605 B.n194 B.n191 10.6151
R1606 B.n195 B.n194 10.6151
R1607 B.n198 B.n195 10.6151
R1608 B.n199 B.n198 10.6151
R1609 B.n202 B.n199 10.6151
R1610 B.n203 B.n202 10.6151
R1611 B.n206 B.n203 10.6151
R1612 B.n207 B.n206 10.6151
R1613 B.n210 B.n207 10.6151
R1614 B.n211 B.n210 10.6151
R1615 B.n214 B.n211 10.6151
R1616 B.n215 B.n214 10.6151
R1617 B.n218 B.n215 10.6151
R1618 B.n219 B.n218 10.6151
R1619 B.n222 B.n219 10.6151
R1620 B.n223 B.n222 10.6151
R1621 B.n226 B.n223 10.6151
R1622 B.n227 B.n226 10.6151
R1623 B.n230 B.n227 10.6151
R1624 B.n231 B.n230 10.6151
R1625 B.n234 B.n231 10.6151
R1626 B.n235 B.n234 10.6151
R1627 B.n238 B.n235 10.6151
R1628 B.n239 B.n238 10.6151
R1629 B.n242 B.n239 10.6151
R1630 B.n243 B.n242 10.6151
R1631 B.n246 B.n243 10.6151
R1632 B.n247 B.n246 10.6151
R1633 B.n250 B.n247 10.6151
R1634 B.n251 B.n250 10.6151
R1635 B.n254 B.n251 10.6151
R1636 B.n255 B.n254 10.6151
R1637 B.n258 B.n255 10.6151
R1638 B.n260 B.n258 10.6151
R1639 B.n261 B.n260 10.6151
R1640 B.n589 B.n261 10.6151
R1641 B.n445 B.n339 8.74196
R1642 B.n422 B.n342 8.74196
R1643 B.n161 B.n160 8.74196
R1644 B.n183 B.n182 8.74196
R1645 B.n628 B.n0 8.11757
R1646 B.n628 B.n1 8.11757
R1647 B.n442 B.n339 1.87367
R1648 B.n425 B.n342 1.87367
R1649 B.n162 B.n161 1.87367
R1650 B.n182 B.n181 1.87367
R1651 VP.n0 VP.t1 541.708
R1652 VP.n0 VP.t0 501.462
R1653 VP VP.n0 0.0516364
R1654 VDD1.n64 VDD1.n63 289.615
R1655 VDD1.n129 VDD1.n128 289.615
R1656 VDD1.n63 VDD1.n62 185
R1657 VDD1.n2 VDD1.n1 185
R1658 VDD1.n57 VDD1.n56 185
R1659 VDD1.n55 VDD1.n54 185
R1660 VDD1.n6 VDD1.n5 185
R1661 VDD1.n49 VDD1.n48 185
R1662 VDD1.n47 VDD1.n46 185
R1663 VDD1.n10 VDD1.n9 185
R1664 VDD1.n41 VDD1.n40 185
R1665 VDD1.n39 VDD1.n38 185
R1666 VDD1.n14 VDD1.n13 185
R1667 VDD1.n33 VDD1.n32 185
R1668 VDD1.n31 VDD1.n30 185
R1669 VDD1.n18 VDD1.n17 185
R1670 VDD1.n25 VDD1.n24 185
R1671 VDD1.n23 VDD1.n22 185
R1672 VDD1.n88 VDD1.n87 185
R1673 VDD1.n90 VDD1.n89 185
R1674 VDD1.n83 VDD1.n82 185
R1675 VDD1.n96 VDD1.n95 185
R1676 VDD1.n98 VDD1.n97 185
R1677 VDD1.n79 VDD1.n78 185
R1678 VDD1.n104 VDD1.n103 185
R1679 VDD1.n106 VDD1.n105 185
R1680 VDD1.n75 VDD1.n74 185
R1681 VDD1.n112 VDD1.n111 185
R1682 VDD1.n114 VDD1.n113 185
R1683 VDD1.n71 VDD1.n70 185
R1684 VDD1.n120 VDD1.n119 185
R1685 VDD1.n122 VDD1.n121 185
R1686 VDD1.n67 VDD1.n66 185
R1687 VDD1.n128 VDD1.n127 185
R1688 VDD1.n21 VDD1.t0 147.659
R1689 VDD1.n86 VDD1.t1 147.659
R1690 VDD1.n63 VDD1.n1 104.615
R1691 VDD1.n56 VDD1.n1 104.615
R1692 VDD1.n56 VDD1.n55 104.615
R1693 VDD1.n55 VDD1.n5 104.615
R1694 VDD1.n48 VDD1.n5 104.615
R1695 VDD1.n48 VDD1.n47 104.615
R1696 VDD1.n47 VDD1.n9 104.615
R1697 VDD1.n40 VDD1.n9 104.615
R1698 VDD1.n40 VDD1.n39 104.615
R1699 VDD1.n39 VDD1.n13 104.615
R1700 VDD1.n32 VDD1.n13 104.615
R1701 VDD1.n32 VDD1.n31 104.615
R1702 VDD1.n31 VDD1.n17 104.615
R1703 VDD1.n24 VDD1.n17 104.615
R1704 VDD1.n24 VDD1.n23 104.615
R1705 VDD1.n89 VDD1.n88 104.615
R1706 VDD1.n89 VDD1.n82 104.615
R1707 VDD1.n96 VDD1.n82 104.615
R1708 VDD1.n97 VDD1.n96 104.615
R1709 VDD1.n97 VDD1.n78 104.615
R1710 VDD1.n104 VDD1.n78 104.615
R1711 VDD1.n105 VDD1.n104 104.615
R1712 VDD1.n105 VDD1.n74 104.615
R1713 VDD1.n112 VDD1.n74 104.615
R1714 VDD1.n113 VDD1.n112 104.615
R1715 VDD1.n113 VDD1.n70 104.615
R1716 VDD1.n120 VDD1.n70 104.615
R1717 VDD1.n121 VDD1.n120 104.615
R1718 VDD1.n121 VDD1.n66 104.615
R1719 VDD1.n128 VDD1.n66 104.615
R1720 VDD1 VDD1.n129 87.3779
R1721 VDD1.n23 VDD1.t0 52.3082
R1722 VDD1.n88 VDD1.t1 52.3082
R1723 VDD1 VDD1.n64 50.7519
R1724 VDD1.n22 VDD1.n21 15.6677
R1725 VDD1.n87 VDD1.n86 15.6677
R1726 VDD1.n25 VDD1.n20 12.8005
R1727 VDD1.n90 VDD1.n85 12.8005
R1728 VDD1.n62 VDD1.n0 12.0247
R1729 VDD1.n26 VDD1.n18 12.0247
R1730 VDD1.n91 VDD1.n83 12.0247
R1731 VDD1.n127 VDD1.n65 12.0247
R1732 VDD1.n61 VDD1.n2 11.249
R1733 VDD1.n30 VDD1.n29 11.249
R1734 VDD1.n95 VDD1.n94 11.249
R1735 VDD1.n126 VDD1.n67 11.249
R1736 VDD1.n58 VDD1.n57 10.4732
R1737 VDD1.n33 VDD1.n16 10.4732
R1738 VDD1.n98 VDD1.n81 10.4732
R1739 VDD1.n123 VDD1.n122 10.4732
R1740 VDD1.n54 VDD1.n4 9.69747
R1741 VDD1.n34 VDD1.n14 9.69747
R1742 VDD1.n99 VDD1.n79 9.69747
R1743 VDD1.n119 VDD1.n69 9.69747
R1744 VDD1.n60 VDD1.n0 9.45567
R1745 VDD1.n125 VDD1.n65 9.45567
R1746 VDD1.n61 VDD1.n60 9.3005
R1747 VDD1.n59 VDD1.n58 9.3005
R1748 VDD1.n4 VDD1.n3 9.3005
R1749 VDD1.n53 VDD1.n52 9.3005
R1750 VDD1.n51 VDD1.n50 9.3005
R1751 VDD1.n8 VDD1.n7 9.3005
R1752 VDD1.n45 VDD1.n44 9.3005
R1753 VDD1.n43 VDD1.n42 9.3005
R1754 VDD1.n12 VDD1.n11 9.3005
R1755 VDD1.n37 VDD1.n36 9.3005
R1756 VDD1.n35 VDD1.n34 9.3005
R1757 VDD1.n16 VDD1.n15 9.3005
R1758 VDD1.n29 VDD1.n28 9.3005
R1759 VDD1.n27 VDD1.n26 9.3005
R1760 VDD1.n20 VDD1.n19 9.3005
R1761 VDD1.n110 VDD1.n109 9.3005
R1762 VDD1.n73 VDD1.n72 9.3005
R1763 VDD1.n116 VDD1.n115 9.3005
R1764 VDD1.n118 VDD1.n117 9.3005
R1765 VDD1.n69 VDD1.n68 9.3005
R1766 VDD1.n124 VDD1.n123 9.3005
R1767 VDD1.n126 VDD1.n125 9.3005
R1768 VDD1.n77 VDD1.n76 9.3005
R1769 VDD1.n102 VDD1.n101 9.3005
R1770 VDD1.n100 VDD1.n99 9.3005
R1771 VDD1.n81 VDD1.n80 9.3005
R1772 VDD1.n94 VDD1.n93 9.3005
R1773 VDD1.n92 VDD1.n91 9.3005
R1774 VDD1.n85 VDD1.n84 9.3005
R1775 VDD1.n108 VDD1.n107 9.3005
R1776 VDD1.n53 VDD1.n6 8.92171
R1777 VDD1.n38 VDD1.n37 8.92171
R1778 VDD1.n103 VDD1.n102 8.92171
R1779 VDD1.n118 VDD1.n71 8.92171
R1780 VDD1.n50 VDD1.n49 8.14595
R1781 VDD1.n41 VDD1.n12 8.14595
R1782 VDD1.n106 VDD1.n77 8.14595
R1783 VDD1.n115 VDD1.n114 8.14595
R1784 VDD1.n46 VDD1.n8 7.3702
R1785 VDD1.n42 VDD1.n10 7.3702
R1786 VDD1.n107 VDD1.n75 7.3702
R1787 VDD1.n111 VDD1.n73 7.3702
R1788 VDD1.n46 VDD1.n45 6.59444
R1789 VDD1.n45 VDD1.n10 6.59444
R1790 VDD1.n110 VDD1.n75 6.59444
R1791 VDD1.n111 VDD1.n110 6.59444
R1792 VDD1.n49 VDD1.n8 5.81868
R1793 VDD1.n42 VDD1.n41 5.81868
R1794 VDD1.n107 VDD1.n106 5.81868
R1795 VDD1.n114 VDD1.n73 5.81868
R1796 VDD1.n50 VDD1.n6 5.04292
R1797 VDD1.n38 VDD1.n12 5.04292
R1798 VDD1.n103 VDD1.n77 5.04292
R1799 VDD1.n115 VDD1.n71 5.04292
R1800 VDD1.n21 VDD1.n19 4.38563
R1801 VDD1.n86 VDD1.n84 4.38563
R1802 VDD1.n54 VDD1.n53 4.26717
R1803 VDD1.n37 VDD1.n14 4.26717
R1804 VDD1.n102 VDD1.n79 4.26717
R1805 VDD1.n119 VDD1.n118 4.26717
R1806 VDD1.n57 VDD1.n4 3.49141
R1807 VDD1.n34 VDD1.n33 3.49141
R1808 VDD1.n99 VDD1.n98 3.49141
R1809 VDD1.n122 VDD1.n69 3.49141
R1810 VDD1.n58 VDD1.n2 2.71565
R1811 VDD1.n30 VDD1.n16 2.71565
R1812 VDD1.n95 VDD1.n81 2.71565
R1813 VDD1.n123 VDD1.n67 2.71565
R1814 VDD1.n62 VDD1.n61 1.93989
R1815 VDD1.n29 VDD1.n18 1.93989
R1816 VDD1.n94 VDD1.n83 1.93989
R1817 VDD1.n127 VDD1.n126 1.93989
R1818 VDD1.n64 VDD1.n0 1.16414
R1819 VDD1.n26 VDD1.n25 1.16414
R1820 VDD1.n91 VDD1.n90 1.16414
R1821 VDD1.n129 VDD1.n65 1.16414
R1822 VDD1.n22 VDD1.n20 0.388379
R1823 VDD1.n87 VDD1.n85 0.388379
R1824 VDD1.n60 VDD1.n59 0.155672
R1825 VDD1.n59 VDD1.n3 0.155672
R1826 VDD1.n52 VDD1.n3 0.155672
R1827 VDD1.n52 VDD1.n51 0.155672
R1828 VDD1.n51 VDD1.n7 0.155672
R1829 VDD1.n44 VDD1.n7 0.155672
R1830 VDD1.n44 VDD1.n43 0.155672
R1831 VDD1.n43 VDD1.n11 0.155672
R1832 VDD1.n36 VDD1.n11 0.155672
R1833 VDD1.n36 VDD1.n35 0.155672
R1834 VDD1.n35 VDD1.n15 0.155672
R1835 VDD1.n28 VDD1.n15 0.155672
R1836 VDD1.n28 VDD1.n27 0.155672
R1837 VDD1.n27 VDD1.n19 0.155672
R1838 VDD1.n92 VDD1.n84 0.155672
R1839 VDD1.n93 VDD1.n92 0.155672
R1840 VDD1.n93 VDD1.n80 0.155672
R1841 VDD1.n100 VDD1.n80 0.155672
R1842 VDD1.n101 VDD1.n100 0.155672
R1843 VDD1.n101 VDD1.n76 0.155672
R1844 VDD1.n108 VDD1.n76 0.155672
R1845 VDD1.n109 VDD1.n108 0.155672
R1846 VDD1.n109 VDD1.n72 0.155672
R1847 VDD1.n116 VDD1.n72 0.155672
R1848 VDD1.n117 VDD1.n116 0.155672
R1849 VDD1.n117 VDD1.n68 0.155672
R1850 VDD1.n124 VDD1.n68 0.155672
R1851 VDD1.n125 VDD1.n124 0.155672
C0 VDD2 VP 0.265459f
C1 VDD1 VN 0.148374f
C2 VDD2 VN 2.19138f
C3 VDD1 VTAIL 5.30205f
C4 VDD2 VTAIL 5.33861f
C5 VDD2 VDD1 0.487959f
C6 VN VP 4.66286f
C7 VTAIL VP 1.7424f
C8 VTAIL VN 1.72787f
C9 VDD1 VP 2.30455f
C10 VDD2 B 3.832699f
C11 VDD1 B 6.26253f
C12 VTAIL B 6.462572f
C13 VN B 8.19454f
C14 VP B 4.333629f
C15 VDD1.n0 B 0.011532f
C16 VDD1.n1 B 0.026043f
C17 VDD1.n2 B 0.011667f
C18 VDD1.n3 B 0.020505f
C19 VDD1.n4 B 0.011018f
C20 VDD1.n5 B 0.026043f
C21 VDD1.n6 B 0.011667f
C22 VDD1.n7 B 0.020505f
C23 VDD1.n8 B 0.011018f
C24 VDD1.n9 B 0.026043f
C25 VDD1.n10 B 0.011667f
C26 VDD1.n11 B 0.020505f
C27 VDD1.n12 B 0.011018f
C28 VDD1.n13 B 0.026043f
C29 VDD1.n14 B 0.011667f
C30 VDD1.n15 B 0.020505f
C31 VDD1.n16 B 0.011018f
C32 VDD1.n17 B 0.026043f
C33 VDD1.n18 B 0.011667f
C34 VDD1.n19 B 1.04275f
C35 VDD1.n20 B 0.011018f
C36 VDD1.t0 B 0.042724f
C37 VDD1.n21 B 0.117799f
C38 VDD1.n22 B 0.015385f
C39 VDD1.n23 B 0.019532f
C40 VDD1.n24 B 0.026043f
C41 VDD1.n25 B 0.011667f
C42 VDD1.n26 B 0.011018f
C43 VDD1.n27 B 0.020505f
C44 VDD1.n28 B 0.020505f
C45 VDD1.n29 B 0.011018f
C46 VDD1.n30 B 0.011667f
C47 VDD1.n31 B 0.026043f
C48 VDD1.n32 B 0.026043f
C49 VDD1.n33 B 0.011667f
C50 VDD1.n34 B 0.011018f
C51 VDD1.n35 B 0.020505f
C52 VDD1.n36 B 0.020505f
C53 VDD1.n37 B 0.011018f
C54 VDD1.n38 B 0.011667f
C55 VDD1.n39 B 0.026043f
C56 VDD1.n40 B 0.026043f
C57 VDD1.n41 B 0.011667f
C58 VDD1.n42 B 0.011018f
C59 VDD1.n43 B 0.020505f
C60 VDD1.n44 B 0.020505f
C61 VDD1.n45 B 0.011018f
C62 VDD1.n46 B 0.011667f
C63 VDD1.n47 B 0.026043f
C64 VDD1.n48 B 0.026043f
C65 VDD1.n49 B 0.011667f
C66 VDD1.n50 B 0.011018f
C67 VDD1.n51 B 0.020505f
C68 VDD1.n52 B 0.020505f
C69 VDD1.n53 B 0.011018f
C70 VDD1.n54 B 0.011667f
C71 VDD1.n55 B 0.026043f
C72 VDD1.n56 B 0.026043f
C73 VDD1.n57 B 0.011667f
C74 VDD1.n58 B 0.011018f
C75 VDD1.n59 B 0.020505f
C76 VDD1.n60 B 0.051317f
C77 VDD1.n61 B 0.011018f
C78 VDD1.n62 B 0.011667f
C79 VDD1.n63 B 0.050997f
C80 VDD1.n64 B 0.057205f
C81 VDD1.n65 B 0.011532f
C82 VDD1.n66 B 0.026043f
C83 VDD1.n67 B 0.011667f
C84 VDD1.n68 B 0.020505f
C85 VDD1.n69 B 0.011018f
C86 VDD1.n70 B 0.026043f
C87 VDD1.n71 B 0.011667f
C88 VDD1.n72 B 0.020505f
C89 VDD1.n73 B 0.011018f
C90 VDD1.n74 B 0.026043f
C91 VDD1.n75 B 0.011667f
C92 VDD1.n76 B 0.020505f
C93 VDD1.n77 B 0.011018f
C94 VDD1.n78 B 0.026043f
C95 VDD1.n79 B 0.011667f
C96 VDD1.n80 B 0.020505f
C97 VDD1.n81 B 0.011018f
C98 VDD1.n82 B 0.026043f
C99 VDD1.n83 B 0.011667f
C100 VDD1.n84 B 1.04275f
C101 VDD1.n85 B 0.011018f
C102 VDD1.t1 B 0.042724f
C103 VDD1.n86 B 0.117799f
C104 VDD1.n87 B 0.015385f
C105 VDD1.n88 B 0.019532f
C106 VDD1.n89 B 0.026043f
C107 VDD1.n90 B 0.011667f
C108 VDD1.n91 B 0.011018f
C109 VDD1.n92 B 0.020505f
C110 VDD1.n93 B 0.020505f
C111 VDD1.n94 B 0.011018f
C112 VDD1.n95 B 0.011667f
C113 VDD1.n96 B 0.026043f
C114 VDD1.n97 B 0.026043f
C115 VDD1.n98 B 0.011667f
C116 VDD1.n99 B 0.011018f
C117 VDD1.n100 B 0.020505f
C118 VDD1.n101 B 0.020505f
C119 VDD1.n102 B 0.011018f
C120 VDD1.n103 B 0.011667f
C121 VDD1.n104 B 0.026043f
C122 VDD1.n105 B 0.026043f
C123 VDD1.n106 B 0.011667f
C124 VDD1.n107 B 0.011018f
C125 VDD1.n108 B 0.020505f
C126 VDD1.n109 B 0.020505f
C127 VDD1.n110 B 0.011018f
C128 VDD1.n111 B 0.011667f
C129 VDD1.n112 B 0.026043f
C130 VDD1.n113 B 0.026043f
C131 VDD1.n114 B 0.011667f
C132 VDD1.n115 B 0.011018f
C133 VDD1.n116 B 0.020505f
C134 VDD1.n117 B 0.020505f
C135 VDD1.n118 B 0.011018f
C136 VDD1.n119 B 0.011667f
C137 VDD1.n120 B 0.026043f
C138 VDD1.n121 B 0.026043f
C139 VDD1.n122 B 0.011667f
C140 VDD1.n123 B 0.011018f
C141 VDD1.n124 B 0.020505f
C142 VDD1.n125 B 0.051317f
C143 VDD1.n126 B 0.011018f
C144 VDD1.n127 B 0.011667f
C145 VDD1.n128 B 0.050997f
C146 VDD1.n129 B 0.546165f
C147 VP.t1 B 1.66602f
C148 VP.t0 B 1.52032f
C149 VP.n0 B 3.79259f
C150 VDD2.n0 B 0.011495f
C151 VDD2.n1 B 0.025959f
C152 VDD2.n2 B 0.011629f
C153 VDD2.n3 B 0.020439f
C154 VDD2.n4 B 0.010983f
C155 VDD2.n5 B 0.025959f
C156 VDD2.n6 B 0.011629f
C157 VDD2.n7 B 0.020439f
C158 VDD2.n8 B 0.010983f
C159 VDD2.n9 B 0.025959f
C160 VDD2.n10 B 0.011629f
C161 VDD2.n11 B 0.020439f
C162 VDD2.n12 B 0.010983f
C163 VDD2.n13 B 0.025959f
C164 VDD2.n14 B 0.011629f
C165 VDD2.n15 B 0.020439f
C166 VDD2.n16 B 0.010983f
C167 VDD2.n17 B 0.025959f
C168 VDD2.n18 B 0.011629f
C169 VDD2.n19 B 1.03938f
C170 VDD2.n20 B 0.010983f
C171 VDD2.t0 B 0.042586f
C172 VDD2.n21 B 0.117419f
C173 VDD2.n22 B 0.015335f
C174 VDD2.n23 B 0.019469f
C175 VDD2.n24 B 0.025959f
C176 VDD2.n25 B 0.011629f
C177 VDD2.n26 B 0.010983f
C178 VDD2.n27 B 0.020439f
C179 VDD2.n28 B 0.020439f
C180 VDD2.n29 B 0.010983f
C181 VDD2.n30 B 0.011629f
C182 VDD2.n31 B 0.025959f
C183 VDD2.n32 B 0.025959f
C184 VDD2.n33 B 0.011629f
C185 VDD2.n34 B 0.010983f
C186 VDD2.n35 B 0.020439f
C187 VDD2.n36 B 0.020439f
C188 VDD2.n37 B 0.010983f
C189 VDD2.n38 B 0.011629f
C190 VDD2.n39 B 0.025959f
C191 VDD2.n40 B 0.025959f
C192 VDD2.n41 B 0.011629f
C193 VDD2.n42 B 0.010983f
C194 VDD2.n43 B 0.020439f
C195 VDD2.n44 B 0.020439f
C196 VDD2.n45 B 0.010983f
C197 VDD2.n46 B 0.011629f
C198 VDD2.n47 B 0.025959f
C199 VDD2.n48 B 0.025959f
C200 VDD2.n49 B 0.011629f
C201 VDD2.n50 B 0.010983f
C202 VDD2.n51 B 0.020439f
C203 VDD2.n52 B 0.020439f
C204 VDD2.n53 B 0.010983f
C205 VDD2.n54 B 0.011629f
C206 VDD2.n55 B 0.025959f
C207 VDD2.n56 B 0.025959f
C208 VDD2.n57 B 0.011629f
C209 VDD2.n58 B 0.010983f
C210 VDD2.n59 B 0.020439f
C211 VDD2.n60 B 0.051152f
C212 VDD2.n61 B 0.010983f
C213 VDD2.n62 B 0.011629f
C214 VDD2.n63 B 0.050833f
C215 VDD2.n64 B 0.515964f
C216 VDD2.n65 B 0.011495f
C217 VDD2.n66 B 0.025959f
C218 VDD2.n67 B 0.011629f
C219 VDD2.n68 B 0.020439f
C220 VDD2.n69 B 0.010983f
C221 VDD2.n70 B 0.025959f
C222 VDD2.n71 B 0.011629f
C223 VDD2.n72 B 0.020439f
C224 VDD2.n73 B 0.010983f
C225 VDD2.n74 B 0.025959f
C226 VDD2.n75 B 0.011629f
C227 VDD2.n76 B 0.020439f
C228 VDD2.n77 B 0.010983f
C229 VDD2.n78 B 0.025959f
C230 VDD2.n79 B 0.011629f
C231 VDD2.n80 B 0.020439f
C232 VDD2.n81 B 0.010983f
C233 VDD2.n82 B 0.025959f
C234 VDD2.n83 B 0.011629f
C235 VDD2.n84 B 1.03938f
C236 VDD2.n85 B 0.010983f
C237 VDD2.t1 B 0.042586f
C238 VDD2.n86 B 0.117419f
C239 VDD2.n87 B 0.015335f
C240 VDD2.n88 B 0.019469f
C241 VDD2.n89 B 0.025959f
C242 VDD2.n90 B 0.011629f
C243 VDD2.n91 B 0.010983f
C244 VDD2.n92 B 0.020439f
C245 VDD2.n93 B 0.020439f
C246 VDD2.n94 B 0.010983f
C247 VDD2.n95 B 0.011629f
C248 VDD2.n96 B 0.025959f
C249 VDD2.n97 B 0.025959f
C250 VDD2.n98 B 0.011629f
C251 VDD2.n99 B 0.010983f
C252 VDD2.n100 B 0.020439f
C253 VDD2.n101 B 0.020439f
C254 VDD2.n102 B 0.010983f
C255 VDD2.n103 B 0.011629f
C256 VDD2.n104 B 0.025959f
C257 VDD2.n105 B 0.025959f
C258 VDD2.n106 B 0.011629f
C259 VDD2.n107 B 0.010983f
C260 VDD2.n108 B 0.020439f
C261 VDD2.n109 B 0.020439f
C262 VDD2.n110 B 0.010983f
C263 VDD2.n111 B 0.011629f
C264 VDD2.n112 B 0.025959f
C265 VDD2.n113 B 0.025959f
C266 VDD2.n114 B 0.011629f
C267 VDD2.n115 B 0.010983f
C268 VDD2.n116 B 0.020439f
C269 VDD2.n117 B 0.020439f
C270 VDD2.n118 B 0.010983f
C271 VDD2.n119 B 0.011629f
C272 VDD2.n120 B 0.025959f
C273 VDD2.n121 B 0.025959f
C274 VDD2.n122 B 0.011629f
C275 VDD2.n123 B 0.010983f
C276 VDD2.n124 B 0.020439f
C277 VDD2.n125 B 0.051152f
C278 VDD2.n126 B 0.010983f
C279 VDD2.n127 B 0.011629f
C280 VDD2.n128 B 0.050833f
C281 VDD2.n129 B 0.056604f
C282 VDD2.n130 B 2.23615f
C283 VTAIL.n0 B 0.008681f
C284 VTAIL.n1 B 0.019605f
C285 VTAIL.n2 B 0.008782f
C286 VTAIL.n3 B 0.015435f
C287 VTAIL.n4 B 0.008294f
C288 VTAIL.n5 B 0.019605f
C289 VTAIL.n6 B 0.008782f
C290 VTAIL.n7 B 0.015435f
C291 VTAIL.n8 B 0.008294f
C292 VTAIL.n9 B 0.019605f
C293 VTAIL.n10 B 0.008782f
C294 VTAIL.n11 B 0.015435f
C295 VTAIL.n12 B 0.008294f
C296 VTAIL.n13 B 0.019605f
C297 VTAIL.n14 B 0.008782f
C298 VTAIL.n15 B 0.015435f
C299 VTAIL.n16 B 0.008294f
C300 VTAIL.n17 B 0.019605f
C301 VTAIL.n18 B 0.008782f
C302 VTAIL.n19 B 0.784943f
C303 VTAIL.n20 B 0.008294f
C304 VTAIL.t0 B 0.032161f
C305 VTAIL.n21 B 0.088675f
C306 VTAIL.n22 B 0.011581f
C307 VTAIL.n23 B 0.014703f
C308 VTAIL.n24 B 0.019605f
C309 VTAIL.n25 B 0.008782f
C310 VTAIL.n26 B 0.008294f
C311 VTAIL.n27 B 0.015435f
C312 VTAIL.n28 B 0.015435f
C313 VTAIL.n29 B 0.008294f
C314 VTAIL.n30 B 0.008782f
C315 VTAIL.n31 B 0.019605f
C316 VTAIL.n32 B 0.019605f
C317 VTAIL.n33 B 0.008782f
C318 VTAIL.n34 B 0.008294f
C319 VTAIL.n35 B 0.015435f
C320 VTAIL.n36 B 0.015435f
C321 VTAIL.n37 B 0.008294f
C322 VTAIL.n38 B 0.008782f
C323 VTAIL.n39 B 0.019605f
C324 VTAIL.n40 B 0.019605f
C325 VTAIL.n41 B 0.008782f
C326 VTAIL.n42 B 0.008294f
C327 VTAIL.n43 B 0.015435f
C328 VTAIL.n44 B 0.015435f
C329 VTAIL.n45 B 0.008294f
C330 VTAIL.n46 B 0.008782f
C331 VTAIL.n47 B 0.019605f
C332 VTAIL.n48 B 0.019605f
C333 VTAIL.n49 B 0.008782f
C334 VTAIL.n50 B 0.008294f
C335 VTAIL.n51 B 0.015435f
C336 VTAIL.n52 B 0.015435f
C337 VTAIL.n53 B 0.008294f
C338 VTAIL.n54 B 0.008782f
C339 VTAIL.n55 B 0.019605f
C340 VTAIL.n56 B 0.019605f
C341 VTAIL.n57 B 0.008782f
C342 VTAIL.n58 B 0.008294f
C343 VTAIL.n59 B 0.015435f
C344 VTAIL.n60 B 0.03863f
C345 VTAIL.n61 B 0.008294f
C346 VTAIL.n62 B 0.008782f
C347 VTAIL.n63 B 0.038389f
C348 VTAIL.n64 B 0.032103f
C349 VTAIL.n65 B 0.88559f
C350 VTAIL.n66 B 0.008681f
C351 VTAIL.n67 B 0.019605f
C352 VTAIL.n68 B 0.008782f
C353 VTAIL.n69 B 0.015435f
C354 VTAIL.n70 B 0.008294f
C355 VTAIL.n71 B 0.019605f
C356 VTAIL.n72 B 0.008782f
C357 VTAIL.n73 B 0.015435f
C358 VTAIL.n74 B 0.008294f
C359 VTAIL.n75 B 0.019605f
C360 VTAIL.n76 B 0.008782f
C361 VTAIL.n77 B 0.015435f
C362 VTAIL.n78 B 0.008294f
C363 VTAIL.n79 B 0.019605f
C364 VTAIL.n80 B 0.008782f
C365 VTAIL.n81 B 0.015435f
C366 VTAIL.n82 B 0.008294f
C367 VTAIL.n83 B 0.019605f
C368 VTAIL.n84 B 0.008782f
C369 VTAIL.n85 B 0.784943f
C370 VTAIL.n86 B 0.008294f
C371 VTAIL.t3 B 0.032161f
C372 VTAIL.n87 B 0.088675f
C373 VTAIL.n88 B 0.011581f
C374 VTAIL.n89 B 0.014703f
C375 VTAIL.n90 B 0.019605f
C376 VTAIL.n91 B 0.008782f
C377 VTAIL.n92 B 0.008294f
C378 VTAIL.n93 B 0.015435f
C379 VTAIL.n94 B 0.015435f
C380 VTAIL.n95 B 0.008294f
C381 VTAIL.n96 B 0.008782f
C382 VTAIL.n97 B 0.019605f
C383 VTAIL.n98 B 0.019605f
C384 VTAIL.n99 B 0.008782f
C385 VTAIL.n100 B 0.008294f
C386 VTAIL.n101 B 0.015435f
C387 VTAIL.n102 B 0.015435f
C388 VTAIL.n103 B 0.008294f
C389 VTAIL.n104 B 0.008782f
C390 VTAIL.n105 B 0.019605f
C391 VTAIL.n106 B 0.019605f
C392 VTAIL.n107 B 0.008782f
C393 VTAIL.n108 B 0.008294f
C394 VTAIL.n109 B 0.015435f
C395 VTAIL.n110 B 0.015435f
C396 VTAIL.n111 B 0.008294f
C397 VTAIL.n112 B 0.008782f
C398 VTAIL.n113 B 0.019605f
C399 VTAIL.n114 B 0.019605f
C400 VTAIL.n115 B 0.008782f
C401 VTAIL.n116 B 0.008294f
C402 VTAIL.n117 B 0.015435f
C403 VTAIL.n118 B 0.015435f
C404 VTAIL.n119 B 0.008294f
C405 VTAIL.n120 B 0.008782f
C406 VTAIL.n121 B 0.019605f
C407 VTAIL.n122 B 0.019605f
C408 VTAIL.n123 B 0.008782f
C409 VTAIL.n124 B 0.008294f
C410 VTAIL.n125 B 0.015435f
C411 VTAIL.n126 B 0.03863f
C412 VTAIL.n127 B 0.008294f
C413 VTAIL.n128 B 0.008782f
C414 VTAIL.n129 B 0.038389f
C415 VTAIL.n130 B 0.032103f
C416 VTAIL.n131 B 0.896523f
C417 VTAIL.n132 B 0.008681f
C418 VTAIL.n133 B 0.019605f
C419 VTAIL.n134 B 0.008782f
C420 VTAIL.n135 B 0.015435f
C421 VTAIL.n136 B 0.008294f
C422 VTAIL.n137 B 0.019605f
C423 VTAIL.n138 B 0.008782f
C424 VTAIL.n139 B 0.015435f
C425 VTAIL.n140 B 0.008294f
C426 VTAIL.n141 B 0.019605f
C427 VTAIL.n142 B 0.008782f
C428 VTAIL.n143 B 0.015435f
C429 VTAIL.n144 B 0.008294f
C430 VTAIL.n145 B 0.019605f
C431 VTAIL.n146 B 0.008782f
C432 VTAIL.n147 B 0.015435f
C433 VTAIL.n148 B 0.008294f
C434 VTAIL.n149 B 0.019605f
C435 VTAIL.n150 B 0.008782f
C436 VTAIL.n151 B 0.784943f
C437 VTAIL.n152 B 0.008294f
C438 VTAIL.t1 B 0.032161f
C439 VTAIL.n153 B 0.088675f
C440 VTAIL.n154 B 0.011581f
C441 VTAIL.n155 B 0.014703f
C442 VTAIL.n156 B 0.019605f
C443 VTAIL.n157 B 0.008782f
C444 VTAIL.n158 B 0.008294f
C445 VTAIL.n159 B 0.015435f
C446 VTAIL.n160 B 0.015435f
C447 VTAIL.n161 B 0.008294f
C448 VTAIL.n162 B 0.008782f
C449 VTAIL.n163 B 0.019605f
C450 VTAIL.n164 B 0.019605f
C451 VTAIL.n165 B 0.008782f
C452 VTAIL.n166 B 0.008294f
C453 VTAIL.n167 B 0.015435f
C454 VTAIL.n168 B 0.015435f
C455 VTAIL.n169 B 0.008294f
C456 VTAIL.n170 B 0.008782f
C457 VTAIL.n171 B 0.019605f
C458 VTAIL.n172 B 0.019605f
C459 VTAIL.n173 B 0.008782f
C460 VTAIL.n174 B 0.008294f
C461 VTAIL.n175 B 0.015435f
C462 VTAIL.n176 B 0.015435f
C463 VTAIL.n177 B 0.008294f
C464 VTAIL.n178 B 0.008782f
C465 VTAIL.n179 B 0.019605f
C466 VTAIL.n180 B 0.019605f
C467 VTAIL.n181 B 0.008782f
C468 VTAIL.n182 B 0.008294f
C469 VTAIL.n183 B 0.015435f
C470 VTAIL.n184 B 0.015435f
C471 VTAIL.n185 B 0.008294f
C472 VTAIL.n186 B 0.008782f
C473 VTAIL.n187 B 0.019605f
C474 VTAIL.n188 B 0.019605f
C475 VTAIL.n189 B 0.008782f
C476 VTAIL.n190 B 0.008294f
C477 VTAIL.n191 B 0.015435f
C478 VTAIL.n192 B 0.03863f
C479 VTAIL.n193 B 0.008294f
C480 VTAIL.n194 B 0.008782f
C481 VTAIL.n195 B 0.038389f
C482 VTAIL.n196 B 0.032103f
C483 VTAIL.n197 B 0.841214f
C484 VTAIL.n198 B 0.008681f
C485 VTAIL.n199 B 0.019605f
C486 VTAIL.n200 B 0.008782f
C487 VTAIL.n201 B 0.015435f
C488 VTAIL.n202 B 0.008294f
C489 VTAIL.n203 B 0.019605f
C490 VTAIL.n204 B 0.008782f
C491 VTAIL.n205 B 0.015435f
C492 VTAIL.n206 B 0.008294f
C493 VTAIL.n207 B 0.019605f
C494 VTAIL.n208 B 0.008782f
C495 VTAIL.n209 B 0.015435f
C496 VTAIL.n210 B 0.008294f
C497 VTAIL.n211 B 0.019605f
C498 VTAIL.n212 B 0.008782f
C499 VTAIL.n213 B 0.015435f
C500 VTAIL.n214 B 0.008294f
C501 VTAIL.n215 B 0.019605f
C502 VTAIL.n216 B 0.008782f
C503 VTAIL.n217 B 0.784943f
C504 VTAIL.n218 B 0.008294f
C505 VTAIL.t2 B 0.032161f
C506 VTAIL.n219 B 0.088675f
C507 VTAIL.n220 B 0.011581f
C508 VTAIL.n221 B 0.014703f
C509 VTAIL.n222 B 0.019605f
C510 VTAIL.n223 B 0.008782f
C511 VTAIL.n224 B 0.008294f
C512 VTAIL.n225 B 0.015435f
C513 VTAIL.n226 B 0.015435f
C514 VTAIL.n227 B 0.008294f
C515 VTAIL.n228 B 0.008782f
C516 VTAIL.n229 B 0.019605f
C517 VTAIL.n230 B 0.019605f
C518 VTAIL.n231 B 0.008782f
C519 VTAIL.n232 B 0.008294f
C520 VTAIL.n233 B 0.015435f
C521 VTAIL.n234 B 0.015435f
C522 VTAIL.n235 B 0.008294f
C523 VTAIL.n236 B 0.008782f
C524 VTAIL.n237 B 0.019605f
C525 VTAIL.n238 B 0.019605f
C526 VTAIL.n239 B 0.008782f
C527 VTAIL.n240 B 0.008294f
C528 VTAIL.n241 B 0.015435f
C529 VTAIL.n242 B 0.015435f
C530 VTAIL.n243 B 0.008294f
C531 VTAIL.n244 B 0.008782f
C532 VTAIL.n245 B 0.019605f
C533 VTAIL.n246 B 0.019605f
C534 VTAIL.n247 B 0.008782f
C535 VTAIL.n248 B 0.008294f
C536 VTAIL.n249 B 0.015435f
C537 VTAIL.n250 B 0.015435f
C538 VTAIL.n251 B 0.008294f
C539 VTAIL.n252 B 0.008782f
C540 VTAIL.n253 B 0.019605f
C541 VTAIL.n254 B 0.019605f
C542 VTAIL.n255 B 0.008782f
C543 VTAIL.n256 B 0.008294f
C544 VTAIL.n257 B 0.015435f
C545 VTAIL.n258 B 0.03863f
C546 VTAIL.n259 B 0.008294f
C547 VTAIL.n260 B 0.008782f
C548 VTAIL.n261 B 0.038389f
C549 VTAIL.n262 B 0.032103f
C550 VTAIL.n263 B 0.801125f
C551 VN.t1 B 1.48628f
C552 VN.t0 B 1.63191f
.ends

