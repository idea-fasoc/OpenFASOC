* NGSPICE file created from diff_pair_sample_1722.ext - technology: sky130A

.subckt diff_pair_sample_1722 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t7 VP.t0 VDD1.t1 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=1.76
X1 B.t11 B.t9 B.t10 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=1.76
X2 VDD1.t3 VP.t1 VTAIL.t6 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=1.76
X3 VTAIL.t1 VN.t0 VDD2.t3 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=1.76
X4 VDD2.t2 VN.t1 VTAIL.t2 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=1.76
X5 B.t8 B.t6 B.t7 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=1.76
X6 VTAIL.t3 VN.t2 VDD2.t1 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=1.76
X7 VTAIL.t5 VP.t2 VDD1.t2 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0.82335 ps=5.32 w=4.99 l=1.76
X8 VDD2.t0 VN.t3 VTAIL.t0 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=1.76
X9 VDD1.t0 VP.t3 VTAIL.t4 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=0.82335 pd=5.32 as=1.9461 ps=10.76 w=4.99 l=1.76
X10 B.t5 B.t3 B.t4 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=1.76
X11 B.t2 B.t0 B.t1 w_n2224_n1966# sky130_fd_pr__pfet_01v8 ad=1.9461 pd=10.76 as=0 ps=0 w=4.99 l=1.76
R0 VP.n5 VP.n4 183.565
R1 VP.n14 VP.n13 183.565
R2 VP.n12 VP.n0 161.3
R3 VP.n11 VP.n10 161.3
R4 VP.n9 VP.n1 161.3
R5 VP.n8 VP.n7 161.3
R6 VP.n6 VP.n2 161.3
R7 VP.n3 VP.t2 104.276
R8 VP.n3 VP.t3 103.85
R9 VP.n5 VP.t0 68.3295
R10 VP.n13 VP.t1 68.3295
R11 VP.n4 VP.n3 47.7203
R12 VP.n7 VP.n1 40.4934
R13 VP.n11 VP.n1 40.4934
R14 VP.n7 VP.n6 24.4675
R15 VP.n12 VP.n11 24.4675
R16 VP.n6 VP.n5 2.20253
R17 VP.n13 VP.n12 2.20253
R18 VP.n4 VP.n2 0.189894
R19 VP.n8 VP.n2 0.189894
R20 VP.n9 VP.n8 0.189894
R21 VP.n10 VP.n9 0.189894
R22 VP.n10 VP.n0 0.189894
R23 VP.n14 VP.n0 0.189894
R24 VP VP.n14 0.0516364
R25 VDD1 VDD1.n1 135.744
R26 VDD1 VDD1.n0 101.856
R27 VDD1.n0 VDD1.t2 6.51453
R28 VDD1.n0 VDD1.t0 6.51453
R29 VDD1.n1 VDD1.t1 6.51453
R30 VDD1.n1 VDD1.t3 6.51453
R31 VTAIL.n5 VTAIL.t5 91.6335
R32 VTAIL.n4 VTAIL.t2 91.6335
R33 VTAIL.n3 VTAIL.t1 91.6335
R34 VTAIL.n7 VTAIL.t0 91.6334
R35 VTAIL.n0 VTAIL.t3 91.6334
R36 VTAIL.n1 VTAIL.t6 91.6334
R37 VTAIL.n2 VTAIL.t7 91.6334
R38 VTAIL.n6 VTAIL.t4 91.6334
R39 VTAIL.n7 VTAIL.n6 18.4703
R40 VTAIL.n3 VTAIL.n2 18.4703
R41 VTAIL.n4 VTAIL.n3 1.80222
R42 VTAIL.n6 VTAIL.n5 1.80222
R43 VTAIL.n2 VTAIL.n1 1.80222
R44 VTAIL VTAIL.n0 0.959552
R45 VTAIL VTAIL.n7 0.843172
R46 VTAIL.n5 VTAIL.n4 0.470328
R47 VTAIL.n1 VTAIL.n0 0.470328
R48 B.n232 B.n73 585
R49 B.n231 B.n230 585
R50 B.n229 B.n74 585
R51 B.n228 B.n227 585
R52 B.n226 B.n75 585
R53 B.n225 B.n224 585
R54 B.n223 B.n76 585
R55 B.n222 B.n221 585
R56 B.n220 B.n77 585
R57 B.n219 B.n218 585
R58 B.n217 B.n78 585
R59 B.n216 B.n215 585
R60 B.n214 B.n79 585
R61 B.n213 B.n212 585
R62 B.n211 B.n80 585
R63 B.n210 B.n209 585
R64 B.n208 B.n81 585
R65 B.n207 B.n206 585
R66 B.n205 B.n82 585
R67 B.n204 B.n203 585
R68 B.n202 B.n83 585
R69 B.n201 B.n200 585
R70 B.n196 B.n84 585
R71 B.n195 B.n194 585
R72 B.n193 B.n85 585
R73 B.n192 B.n191 585
R74 B.n190 B.n86 585
R75 B.n189 B.n188 585
R76 B.n187 B.n87 585
R77 B.n186 B.n185 585
R78 B.n184 B.n88 585
R79 B.n182 B.n181 585
R80 B.n180 B.n91 585
R81 B.n179 B.n178 585
R82 B.n177 B.n92 585
R83 B.n176 B.n175 585
R84 B.n174 B.n93 585
R85 B.n173 B.n172 585
R86 B.n171 B.n94 585
R87 B.n170 B.n169 585
R88 B.n168 B.n95 585
R89 B.n167 B.n166 585
R90 B.n165 B.n96 585
R91 B.n164 B.n163 585
R92 B.n162 B.n97 585
R93 B.n161 B.n160 585
R94 B.n159 B.n98 585
R95 B.n158 B.n157 585
R96 B.n156 B.n99 585
R97 B.n155 B.n154 585
R98 B.n153 B.n100 585
R99 B.n152 B.n151 585
R100 B.n234 B.n233 585
R101 B.n235 B.n72 585
R102 B.n237 B.n236 585
R103 B.n238 B.n71 585
R104 B.n240 B.n239 585
R105 B.n241 B.n70 585
R106 B.n243 B.n242 585
R107 B.n244 B.n69 585
R108 B.n246 B.n245 585
R109 B.n247 B.n68 585
R110 B.n249 B.n248 585
R111 B.n250 B.n67 585
R112 B.n252 B.n251 585
R113 B.n253 B.n66 585
R114 B.n255 B.n254 585
R115 B.n256 B.n65 585
R116 B.n258 B.n257 585
R117 B.n259 B.n64 585
R118 B.n261 B.n260 585
R119 B.n262 B.n63 585
R120 B.n264 B.n263 585
R121 B.n265 B.n62 585
R122 B.n267 B.n266 585
R123 B.n268 B.n61 585
R124 B.n270 B.n269 585
R125 B.n271 B.n60 585
R126 B.n273 B.n272 585
R127 B.n274 B.n59 585
R128 B.n276 B.n275 585
R129 B.n277 B.n58 585
R130 B.n279 B.n278 585
R131 B.n280 B.n57 585
R132 B.n282 B.n281 585
R133 B.n283 B.n56 585
R134 B.n285 B.n284 585
R135 B.n286 B.n55 585
R136 B.n288 B.n287 585
R137 B.n289 B.n54 585
R138 B.n291 B.n290 585
R139 B.n292 B.n53 585
R140 B.n294 B.n293 585
R141 B.n295 B.n52 585
R142 B.n297 B.n296 585
R143 B.n298 B.n51 585
R144 B.n300 B.n299 585
R145 B.n301 B.n50 585
R146 B.n303 B.n302 585
R147 B.n304 B.n49 585
R148 B.n306 B.n305 585
R149 B.n307 B.n48 585
R150 B.n309 B.n308 585
R151 B.n310 B.n47 585
R152 B.n312 B.n311 585
R153 B.n313 B.n46 585
R154 B.n392 B.n15 585
R155 B.n391 B.n390 585
R156 B.n389 B.n16 585
R157 B.n388 B.n387 585
R158 B.n386 B.n17 585
R159 B.n385 B.n384 585
R160 B.n383 B.n18 585
R161 B.n382 B.n381 585
R162 B.n380 B.n19 585
R163 B.n379 B.n378 585
R164 B.n377 B.n20 585
R165 B.n376 B.n375 585
R166 B.n374 B.n21 585
R167 B.n373 B.n372 585
R168 B.n371 B.n22 585
R169 B.n370 B.n369 585
R170 B.n368 B.n23 585
R171 B.n367 B.n366 585
R172 B.n365 B.n24 585
R173 B.n364 B.n363 585
R174 B.n362 B.n25 585
R175 B.n360 B.n359 585
R176 B.n358 B.n28 585
R177 B.n357 B.n356 585
R178 B.n355 B.n29 585
R179 B.n354 B.n353 585
R180 B.n352 B.n30 585
R181 B.n351 B.n350 585
R182 B.n349 B.n31 585
R183 B.n348 B.n347 585
R184 B.n346 B.n32 585
R185 B.n345 B.n344 585
R186 B.n343 B.n33 585
R187 B.n342 B.n341 585
R188 B.n340 B.n37 585
R189 B.n339 B.n338 585
R190 B.n337 B.n38 585
R191 B.n336 B.n335 585
R192 B.n334 B.n39 585
R193 B.n333 B.n332 585
R194 B.n331 B.n40 585
R195 B.n330 B.n329 585
R196 B.n328 B.n41 585
R197 B.n327 B.n326 585
R198 B.n325 B.n42 585
R199 B.n324 B.n323 585
R200 B.n322 B.n43 585
R201 B.n321 B.n320 585
R202 B.n319 B.n44 585
R203 B.n318 B.n317 585
R204 B.n316 B.n45 585
R205 B.n315 B.n314 585
R206 B.n394 B.n393 585
R207 B.n395 B.n14 585
R208 B.n397 B.n396 585
R209 B.n398 B.n13 585
R210 B.n400 B.n399 585
R211 B.n401 B.n12 585
R212 B.n403 B.n402 585
R213 B.n404 B.n11 585
R214 B.n406 B.n405 585
R215 B.n407 B.n10 585
R216 B.n409 B.n408 585
R217 B.n410 B.n9 585
R218 B.n412 B.n411 585
R219 B.n413 B.n8 585
R220 B.n415 B.n414 585
R221 B.n416 B.n7 585
R222 B.n418 B.n417 585
R223 B.n419 B.n6 585
R224 B.n421 B.n420 585
R225 B.n422 B.n5 585
R226 B.n424 B.n423 585
R227 B.n425 B.n4 585
R228 B.n427 B.n426 585
R229 B.n428 B.n3 585
R230 B.n430 B.n429 585
R231 B.n431 B.n0 585
R232 B.n2 B.n1 585
R233 B.n114 B.n113 585
R234 B.n116 B.n115 585
R235 B.n117 B.n112 585
R236 B.n119 B.n118 585
R237 B.n120 B.n111 585
R238 B.n122 B.n121 585
R239 B.n123 B.n110 585
R240 B.n125 B.n124 585
R241 B.n126 B.n109 585
R242 B.n128 B.n127 585
R243 B.n129 B.n108 585
R244 B.n131 B.n130 585
R245 B.n132 B.n107 585
R246 B.n134 B.n133 585
R247 B.n135 B.n106 585
R248 B.n137 B.n136 585
R249 B.n138 B.n105 585
R250 B.n140 B.n139 585
R251 B.n141 B.n104 585
R252 B.n143 B.n142 585
R253 B.n144 B.n103 585
R254 B.n146 B.n145 585
R255 B.n147 B.n102 585
R256 B.n149 B.n148 585
R257 B.n150 B.n101 585
R258 B.n151 B.n150 473.281
R259 B.n233 B.n232 473.281
R260 B.n315 B.n46 473.281
R261 B.n394 B.n15 473.281
R262 B.n89 B.t9 274.622
R263 B.n197 B.t6 274.622
R264 B.n34 B.t3 274.622
R265 B.n26 B.t0 274.622
R266 B.n433 B.n432 256.663
R267 B.n432 B.n431 235.042
R268 B.n432 B.n2 235.042
R269 B.n151 B.n100 163.367
R270 B.n155 B.n100 163.367
R271 B.n156 B.n155 163.367
R272 B.n157 B.n156 163.367
R273 B.n157 B.n98 163.367
R274 B.n161 B.n98 163.367
R275 B.n162 B.n161 163.367
R276 B.n163 B.n162 163.367
R277 B.n163 B.n96 163.367
R278 B.n167 B.n96 163.367
R279 B.n168 B.n167 163.367
R280 B.n169 B.n168 163.367
R281 B.n169 B.n94 163.367
R282 B.n173 B.n94 163.367
R283 B.n174 B.n173 163.367
R284 B.n175 B.n174 163.367
R285 B.n175 B.n92 163.367
R286 B.n179 B.n92 163.367
R287 B.n180 B.n179 163.367
R288 B.n181 B.n180 163.367
R289 B.n181 B.n88 163.367
R290 B.n186 B.n88 163.367
R291 B.n187 B.n186 163.367
R292 B.n188 B.n187 163.367
R293 B.n188 B.n86 163.367
R294 B.n192 B.n86 163.367
R295 B.n193 B.n192 163.367
R296 B.n194 B.n193 163.367
R297 B.n194 B.n84 163.367
R298 B.n201 B.n84 163.367
R299 B.n202 B.n201 163.367
R300 B.n203 B.n202 163.367
R301 B.n203 B.n82 163.367
R302 B.n207 B.n82 163.367
R303 B.n208 B.n207 163.367
R304 B.n209 B.n208 163.367
R305 B.n209 B.n80 163.367
R306 B.n213 B.n80 163.367
R307 B.n214 B.n213 163.367
R308 B.n215 B.n214 163.367
R309 B.n215 B.n78 163.367
R310 B.n219 B.n78 163.367
R311 B.n220 B.n219 163.367
R312 B.n221 B.n220 163.367
R313 B.n221 B.n76 163.367
R314 B.n225 B.n76 163.367
R315 B.n226 B.n225 163.367
R316 B.n227 B.n226 163.367
R317 B.n227 B.n74 163.367
R318 B.n231 B.n74 163.367
R319 B.n232 B.n231 163.367
R320 B.n311 B.n46 163.367
R321 B.n311 B.n310 163.367
R322 B.n310 B.n309 163.367
R323 B.n309 B.n48 163.367
R324 B.n305 B.n48 163.367
R325 B.n305 B.n304 163.367
R326 B.n304 B.n303 163.367
R327 B.n303 B.n50 163.367
R328 B.n299 B.n50 163.367
R329 B.n299 B.n298 163.367
R330 B.n298 B.n297 163.367
R331 B.n297 B.n52 163.367
R332 B.n293 B.n52 163.367
R333 B.n293 B.n292 163.367
R334 B.n292 B.n291 163.367
R335 B.n291 B.n54 163.367
R336 B.n287 B.n54 163.367
R337 B.n287 B.n286 163.367
R338 B.n286 B.n285 163.367
R339 B.n285 B.n56 163.367
R340 B.n281 B.n56 163.367
R341 B.n281 B.n280 163.367
R342 B.n280 B.n279 163.367
R343 B.n279 B.n58 163.367
R344 B.n275 B.n58 163.367
R345 B.n275 B.n274 163.367
R346 B.n274 B.n273 163.367
R347 B.n273 B.n60 163.367
R348 B.n269 B.n60 163.367
R349 B.n269 B.n268 163.367
R350 B.n268 B.n267 163.367
R351 B.n267 B.n62 163.367
R352 B.n263 B.n62 163.367
R353 B.n263 B.n262 163.367
R354 B.n262 B.n261 163.367
R355 B.n261 B.n64 163.367
R356 B.n257 B.n64 163.367
R357 B.n257 B.n256 163.367
R358 B.n256 B.n255 163.367
R359 B.n255 B.n66 163.367
R360 B.n251 B.n66 163.367
R361 B.n251 B.n250 163.367
R362 B.n250 B.n249 163.367
R363 B.n249 B.n68 163.367
R364 B.n245 B.n68 163.367
R365 B.n245 B.n244 163.367
R366 B.n244 B.n243 163.367
R367 B.n243 B.n70 163.367
R368 B.n239 B.n70 163.367
R369 B.n239 B.n238 163.367
R370 B.n238 B.n237 163.367
R371 B.n237 B.n72 163.367
R372 B.n233 B.n72 163.367
R373 B.n390 B.n15 163.367
R374 B.n390 B.n389 163.367
R375 B.n389 B.n388 163.367
R376 B.n388 B.n17 163.367
R377 B.n384 B.n17 163.367
R378 B.n384 B.n383 163.367
R379 B.n383 B.n382 163.367
R380 B.n382 B.n19 163.367
R381 B.n378 B.n19 163.367
R382 B.n378 B.n377 163.367
R383 B.n377 B.n376 163.367
R384 B.n376 B.n21 163.367
R385 B.n372 B.n21 163.367
R386 B.n372 B.n371 163.367
R387 B.n371 B.n370 163.367
R388 B.n370 B.n23 163.367
R389 B.n366 B.n23 163.367
R390 B.n366 B.n365 163.367
R391 B.n365 B.n364 163.367
R392 B.n364 B.n25 163.367
R393 B.n359 B.n25 163.367
R394 B.n359 B.n358 163.367
R395 B.n358 B.n357 163.367
R396 B.n357 B.n29 163.367
R397 B.n353 B.n29 163.367
R398 B.n353 B.n352 163.367
R399 B.n352 B.n351 163.367
R400 B.n351 B.n31 163.367
R401 B.n347 B.n31 163.367
R402 B.n347 B.n346 163.367
R403 B.n346 B.n345 163.367
R404 B.n345 B.n33 163.367
R405 B.n341 B.n33 163.367
R406 B.n341 B.n340 163.367
R407 B.n340 B.n339 163.367
R408 B.n339 B.n38 163.367
R409 B.n335 B.n38 163.367
R410 B.n335 B.n334 163.367
R411 B.n334 B.n333 163.367
R412 B.n333 B.n40 163.367
R413 B.n329 B.n40 163.367
R414 B.n329 B.n328 163.367
R415 B.n328 B.n327 163.367
R416 B.n327 B.n42 163.367
R417 B.n323 B.n42 163.367
R418 B.n323 B.n322 163.367
R419 B.n322 B.n321 163.367
R420 B.n321 B.n44 163.367
R421 B.n317 B.n44 163.367
R422 B.n317 B.n316 163.367
R423 B.n316 B.n315 163.367
R424 B.n395 B.n394 163.367
R425 B.n396 B.n395 163.367
R426 B.n396 B.n13 163.367
R427 B.n400 B.n13 163.367
R428 B.n401 B.n400 163.367
R429 B.n402 B.n401 163.367
R430 B.n402 B.n11 163.367
R431 B.n406 B.n11 163.367
R432 B.n407 B.n406 163.367
R433 B.n408 B.n407 163.367
R434 B.n408 B.n9 163.367
R435 B.n412 B.n9 163.367
R436 B.n413 B.n412 163.367
R437 B.n414 B.n413 163.367
R438 B.n414 B.n7 163.367
R439 B.n418 B.n7 163.367
R440 B.n419 B.n418 163.367
R441 B.n420 B.n419 163.367
R442 B.n420 B.n5 163.367
R443 B.n424 B.n5 163.367
R444 B.n425 B.n424 163.367
R445 B.n426 B.n425 163.367
R446 B.n426 B.n3 163.367
R447 B.n430 B.n3 163.367
R448 B.n431 B.n430 163.367
R449 B.n114 B.n2 163.367
R450 B.n115 B.n114 163.367
R451 B.n115 B.n112 163.367
R452 B.n119 B.n112 163.367
R453 B.n120 B.n119 163.367
R454 B.n121 B.n120 163.367
R455 B.n121 B.n110 163.367
R456 B.n125 B.n110 163.367
R457 B.n126 B.n125 163.367
R458 B.n127 B.n126 163.367
R459 B.n127 B.n108 163.367
R460 B.n131 B.n108 163.367
R461 B.n132 B.n131 163.367
R462 B.n133 B.n132 163.367
R463 B.n133 B.n106 163.367
R464 B.n137 B.n106 163.367
R465 B.n138 B.n137 163.367
R466 B.n139 B.n138 163.367
R467 B.n139 B.n104 163.367
R468 B.n143 B.n104 163.367
R469 B.n144 B.n143 163.367
R470 B.n145 B.n144 163.367
R471 B.n145 B.n102 163.367
R472 B.n149 B.n102 163.367
R473 B.n150 B.n149 163.367
R474 B.n197 B.t7 159.526
R475 B.n34 B.t5 159.526
R476 B.n89 B.t10 159.522
R477 B.n26 B.t2 159.522
R478 B.n198 B.t8 118.993
R479 B.n35 B.t4 118.993
R480 B.n90 B.t11 118.989
R481 B.n27 B.t1 118.989
R482 B.n183 B.n90 59.5399
R483 B.n199 B.n198 59.5399
R484 B.n36 B.n35 59.5399
R485 B.n361 B.n27 59.5399
R486 B.n90 B.n89 40.5338
R487 B.n198 B.n197 40.5338
R488 B.n35 B.n34 40.5338
R489 B.n27 B.n26 40.5338
R490 B.n234 B.n73 30.7517
R491 B.n393 B.n392 30.7517
R492 B.n314 B.n313 30.7517
R493 B.n152 B.n101 30.7517
R494 B B.n433 18.0485
R495 B.n393 B.n14 10.6151
R496 B.n397 B.n14 10.6151
R497 B.n398 B.n397 10.6151
R498 B.n399 B.n398 10.6151
R499 B.n399 B.n12 10.6151
R500 B.n403 B.n12 10.6151
R501 B.n404 B.n403 10.6151
R502 B.n405 B.n404 10.6151
R503 B.n405 B.n10 10.6151
R504 B.n409 B.n10 10.6151
R505 B.n410 B.n409 10.6151
R506 B.n411 B.n410 10.6151
R507 B.n411 B.n8 10.6151
R508 B.n415 B.n8 10.6151
R509 B.n416 B.n415 10.6151
R510 B.n417 B.n416 10.6151
R511 B.n417 B.n6 10.6151
R512 B.n421 B.n6 10.6151
R513 B.n422 B.n421 10.6151
R514 B.n423 B.n422 10.6151
R515 B.n423 B.n4 10.6151
R516 B.n427 B.n4 10.6151
R517 B.n428 B.n427 10.6151
R518 B.n429 B.n428 10.6151
R519 B.n429 B.n0 10.6151
R520 B.n392 B.n391 10.6151
R521 B.n391 B.n16 10.6151
R522 B.n387 B.n16 10.6151
R523 B.n387 B.n386 10.6151
R524 B.n386 B.n385 10.6151
R525 B.n385 B.n18 10.6151
R526 B.n381 B.n18 10.6151
R527 B.n381 B.n380 10.6151
R528 B.n380 B.n379 10.6151
R529 B.n379 B.n20 10.6151
R530 B.n375 B.n20 10.6151
R531 B.n375 B.n374 10.6151
R532 B.n374 B.n373 10.6151
R533 B.n373 B.n22 10.6151
R534 B.n369 B.n22 10.6151
R535 B.n369 B.n368 10.6151
R536 B.n368 B.n367 10.6151
R537 B.n367 B.n24 10.6151
R538 B.n363 B.n24 10.6151
R539 B.n363 B.n362 10.6151
R540 B.n360 B.n28 10.6151
R541 B.n356 B.n28 10.6151
R542 B.n356 B.n355 10.6151
R543 B.n355 B.n354 10.6151
R544 B.n354 B.n30 10.6151
R545 B.n350 B.n30 10.6151
R546 B.n350 B.n349 10.6151
R547 B.n349 B.n348 10.6151
R548 B.n348 B.n32 10.6151
R549 B.n344 B.n343 10.6151
R550 B.n343 B.n342 10.6151
R551 B.n342 B.n37 10.6151
R552 B.n338 B.n37 10.6151
R553 B.n338 B.n337 10.6151
R554 B.n337 B.n336 10.6151
R555 B.n336 B.n39 10.6151
R556 B.n332 B.n39 10.6151
R557 B.n332 B.n331 10.6151
R558 B.n331 B.n330 10.6151
R559 B.n330 B.n41 10.6151
R560 B.n326 B.n41 10.6151
R561 B.n326 B.n325 10.6151
R562 B.n325 B.n324 10.6151
R563 B.n324 B.n43 10.6151
R564 B.n320 B.n43 10.6151
R565 B.n320 B.n319 10.6151
R566 B.n319 B.n318 10.6151
R567 B.n318 B.n45 10.6151
R568 B.n314 B.n45 10.6151
R569 B.n313 B.n312 10.6151
R570 B.n312 B.n47 10.6151
R571 B.n308 B.n47 10.6151
R572 B.n308 B.n307 10.6151
R573 B.n307 B.n306 10.6151
R574 B.n306 B.n49 10.6151
R575 B.n302 B.n49 10.6151
R576 B.n302 B.n301 10.6151
R577 B.n301 B.n300 10.6151
R578 B.n300 B.n51 10.6151
R579 B.n296 B.n51 10.6151
R580 B.n296 B.n295 10.6151
R581 B.n295 B.n294 10.6151
R582 B.n294 B.n53 10.6151
R583 B.n290 B.n53 10.6151
R584 B.n290 B.n289 10.6151
R585 B.n289 B.n288 10.6151
R586 B.n288 B.n55 10.6151
R587 B.n284 B.n55 10.6151
R588 B.n284 B.n283 10.6151
R589 B.n283 B.n282 10.6151
R590 B.n282 B.n57 10.6151
R591 B.n278 B.n57 10.6151
R592 B.n278 B.n277 10.6151
R593 B.n277 B.n276 10.6151
R594 B.n276 B.n59 10.6151
R595 B.n272 B.n59 10.6151
R596 B.n272 B.n271 10.6151
R597 B.n271 B.n270 10.6151
R598 B.n270 B.n61 10.6151
R599 B.n266 B.n61 10.6151
R600 B.n266 B.n265 10.6151
R601 B.n265 B.n264 10.6151
R602 B.n264 B.n63 10.6151
R603 B.n260 B.n63 10.6151
R604 B.n260 B.n259 10.6151
R605 B.n259 B.n258 10.6151
R606 B.n258 B.n65 10.6151
R607 B.n254 B.n65 10.6151
R608 B.n254 B.n253 10.6151
R609 B.n253 B.n252 10.6151
R610 B.n252 B.n67 10.6151
R611 B.n248 B.n67 10.6151
R612 B.n248 B.n247 10.6151
R613 B.n247 B.n246 10.6151
R614 B.n246 B.n69 10.6151
R615 B.n242 B.n69 10.6151
R616 B.n242 B.n241 10.6151
R617 B.n241 B.n240 10.6151
R618 B.n240 B.n71 10.6151
R619 B.n236 B.n71 10.6151
R620 B.n236 B.n235 10.6151
R621 B.n235 B.n234 10.6151
R622 B.n113 B.n1 10.6151
R623 B.n116 B.n113 10.6151
R624 B.n117 B.n116 10.6151
R625 B.n118 B.n117 10.6151
R626 B.n118 B.n111 10.6151
R627 B.n122 B.n111 10.6151
R628 B.n123 B.n122 10.6151
R629 B.n124 B.n123 10.6151
R630 B.n124 B.n109 10.6151
R631 B.n128 B.n109 10.6151
R632 B.n129 B.n128 10.6151
R633 B.n130 B.n129 10.6151
R634 B.n130 B.n107 10.6151
R635 B.n134 B.n107 10.6151
R636 B.n135 B.n134 10.6151
R637 B.n136 B.n135 10.6151
R638 B.n136 B.n105 10.6151
R639 B.n140 B.n105 10.6151
R640 B.n141 B.n140 10.6151
R641 B.n142 B.n141 10.6151
R642 B.n142 B.n103 10.6151
R643 B.n146 B.n103 10.6151
R644 B.n147 B.n146 10.6151
R645 B.n148 B.n147 10.6151
R646 B.n148 B.n101 10.6151
R647 B.n153 B.n152 10.6151
R648 B.n154 B.n153 10.6151
R649 B.n154 B.n99 10.6151
R650 B.n158 B.n99 10.6151
R651 B.n159 B.n158 10.6151
R652 B.n160 B.n159 10.6151
R653 B.n160 B.n97 10.6151
R654 B.n164 B.n97 10.6151
R655 B.n165 B.n164 10.6151
R656 B.n166 B.n165 10.6151
R657 B.n166 B.n95 10.6151
R658 B.n170 B.n95 10.6151
R659 B.n171 B.n170 10.6151
R660 B.n172 B.n171 10.6151
R661 B.n172 B.n93 10.6151
R662 B.n176 B.n93 10.6151
R663 B.n177 B.n176 10.6151
R664 B.n178 B.n177 10.6151
R665 B.n178 B.n91 10.6151
R666 B.n182 B.n91 10.6151
R667 B.n185 B.n184 10.6151
R668 B.n185 B.n87 10.6151
R669 B.n189 B.n87 10.6151
R670 B.n190 B.n189 10.6151
R671 B.n191 B.n190 10.6151
R672 B.n191 B.n85 10.6151
R673 B.n195 B.n85 10.6151
R674 B.n196 B.n195 10.6151
R675 B.n200 B.n196 10.6151
R676 B.n204 B.n83 10.6151
R677 B.n205 B.n204 10.6151
R678 B.n206 B.n205 10.6151
R679 B.n206 B.n81 10.6151
R680 B.n210 B.n81 10.6151
R681 B.n211 B.n210 10.6151
R682 B.n212 B.n211 10.6151
R683 B.n212 B.n79 10.6151
R684 B.n216 B.n79 10.6151
R685 B.n217 B.n216 10.6151
R686 B.n218 B.n217 10.6151
R687 B.n218 B.n77 10.6151
R688 B.n222 B.n77 10.6151
R689 B.n223 B.n222 10.6151
R690 B.n224 B.n223 10.6151
R691 B.n224 B.n75 10.6151
R692 B.n228 B.n75 10.6151
R693 B.n229 B.n228 10.6151
R694 B.n230 B.n229 10.6151
R695 B.n230 B.n73 10.6151
R696 B.n362 B.n361 9.36635
R697 B.n344 B.n36 9.36635
R698 B.n183 B.n182 9.36635
R699 B.n199 B.n83 9.36635
R700 B.n433 B.n0 8.11757
R701 B.n433 B.n1 8.11757
R702 B.n361 B.n360 1.24928
R703 B.n36 B.n32 1.24928
R704 B.n184 B.n183 1.24928
R705 B.n200 B.n199 1.24928
R706 VN.n0 VN.t2 104.276
R707 VN.n1 VN.t1 104.276
R708 VN.n0 VN.t3 103.85
R709 VN.n1 VN.t0 103.85
R710 VN VN.n1 48.1009
R711 VN VN.n0 9.41534
R712 VDD2.n2 VDD2.n0 135.22
R713 VDD2.n2 VDD2.n1 101.799
R714 VDD2.n1 VDD2.t3 6.51453
R715 VDD2.n1 VDD2.t2 6.51453
R716 VDD2.n0 VDD2.t1 6.51453
R717 VDD2.n0 VDD2.t0 6.51453
R718 VDD2 VDD2.n2 0.0586897
C0 VN VDD1 0.148062f
C1 VP VTAIL 2.19018f
C2 VP B 1.3397f
C3 VN VTAIL 2.17607f
C4 VN B 0.872755f
C5 VTAIL VDD1 3.46411f
C6 B VDD1 0.925396f
C7 B VTAIL 2.34651f
C8 w_n2224_n1966# VDD2 1.13387f
C9 w_n2224_n1966# VP 3.76698f
C10 w_n2224_n1966# VN 3.48329f
C11 w_n2224_n1966# VDD1 1.09682f
C12 w_n2224_n1966# VTAIL 2.33632f
C13 w_n2224_n1966# B 6.25377f
C14 VP VDD2 0.344767f
C15 VN VDD2 2.00256f
C16 VDD2 VDD1 0.821847f
C17 VN VP 4.28831f
C18 VDD2 VTAIL 3.51269f
C19 VDD2 B 0.963887f
C20 VP VDD1 2.1946f
C21 VDD2 VSUBS 0.639987f
C22 VDD1 VSUBS 4.315526f
C23 VTAIL VSUBS 0.585678f
C24 VN VSUBS 4.930009f
C25 VP VSUBS 1.451366f
C26 B VSUBS 2.814513f
C27 w_n2224_n1966# VSUBS 54.7905f
C28 VDD2.t1 VSUBS 0.107201f
C29 VDD2.t0 VSUBS 0.107201f
C30 VDD2.n0 VSUBS 1.01216f
C31 VDD2.t3 VSUBS 0.107201f
C32 VDD2.t2 VSUBS 0.107201f
C33 VDD2.n1 VSUBS 0.673902f
C34 VDD2.n2 VSUBS 3.22146f
C35 VN.t2 VSUBS 1.40473f
C36 VN.t3 VSUBS 1.40185f
C37 VN.n0 VSUBS 1.01532f
C38 VN.t1 VSUBS 1.40473f
C39 VN.t0 VSUBS 1.40185f
C40 VN.n1 VSUBS 2.74818f
C41 B.n0 VSUBS 0.008007f
C42 B.n1 VSUBS 0.008007f
C43 B.n2 VSUBS 0.011842f
C44 B.n3 VSUBS 0.009074f
C45 B.n4 VSUBS 0.009074f
C46 B.n5 VSUBS 0.009074f
C47 B.n6 VSUBS 0.009074f
C48 B.n7 VSUBS 0.009074f
C49 B.n8 VSUBS 0.009074f
C50 B.n9 VSUBS 0.009074f
C51 B.n10 VSUBS 0.009074f
C52 B.n11 VSUBS 0.009074f
C53 B.n12 VSUBS 0.009074f
C54 B.n13 VSUBS 0.009074f
C55 B.n14 VSUBS 0.009074f
C56 B.n15 VSUBS 0.021209f
C57 B.n16 VSUBS 0.009074f
C58 B.n17 VSUBS 0.009074f
C59 B.n18 VSUBS 0.009074f
C60 B.n19 VSUBS 0.009074f
C61 B.n20 VSUBS 0.009074f
C62 B.n21 VSUBS 0.009074f
C63 B.n22 VSUBS 0.009074f
C64 B.n23 VSUBS 0.009074f
C65 B.n24 VSUBS 0.009074f
C66 B.n25 VSUBS 0.009074f
C67 B.t1 VSUBS 0.180427f
C68 B.t2 VSUBS 0.199125f
C69 B.t0 VSUBS 0.532568f
C70 B.n26 VSUBS 0.123551f
C71 B.n27 VSUBS 0.086529f
C72 B.n28 VSUBS 0.009074f
C73 B.n29 VSUBS 0.009074f
C74 B.n30 VSUBS 0.009074f
C75 B.n31 VSUBS 0.009074f
C76 B.n32 VSUBS 0.005071f
C77 B.n33 VSUBS 0.009074f
C78 B.t4 VSUBS 0.180427f
C79 B.t5 VSUBS 0.199124f
C80 B.t3 VSUBS 0.532568f
C81 B.n34 VSUBS 0.123551f
C82 B.n35 VSUBS 0.086529f
C83 B.n36 VSUBS 0.021024f
C84 B.n37 VSUBS 0.009074f
C85 B.n38 VSUBS 0.009074f
C86 B.n39 VSUBS 0.009074f
C87 B.n40 VSUBS 0.009074f
C88 B.n41 VSUBS 0.009074f
C89 B.n42 VSUBS 0.009074f
C90 B.n43 VSUBS 0.009074f
C91 B.n44 VSUBS 0.009074f
C92 B.n45 VSUBS 0.009074f
C93 B.n46 VSUBS 0.019626f
C94 B.n47 VSUBS 0.009074f
C95 B.n48 VSUBS 0.009074f
C96 B.n49 VSUBS 0.009074f
C97 B.n50 VSUBS 0.009074f
C98 B.n51 VSUBS 0.009074f
C99 B.n52 VSUBS 0.009074f
C100 B.n53 VSUBS 0.009074f
C101 B.n54 VSUBS 0.009074f
C102 B.n55 VSUBS 0.009074f
C103 B.n56 VSUBS 0.009074f
C104 B.n57 VSUBS 0.009074f
C105 B.n58 VSUBS 0.009074f
C106 B.n59 VSUBS 0.009074f
C107 B.n60 VSUBS 0.009074f
C108 B.n61 VSUBS 0.009074f
C109 B.n62 VSUBS 0.009074f
C110 B.n63 VSUBS 0.009074f
C111 B.n64 VSUBS 0.009074f
C112 B.n65 VSUBS 0.009074f
C113 B.n66 VSUBS 0.009074f
C114 B.n67 VSUBS 0.009074f
C115 B.n68 VSUBS 0.009074f
C116 B.n69 VSUBS 0.009074f
C117 B.n70 VSUBS 0.009074f
C118 B.n71 VSUBS 0.009074f
C119 B.n72 VSUBS 0.009074f
C120 B.n73 VSUBS 0.02007f
C121 B.n74 VSUBS 0.009074f
C122 B.n75 VSUBS 0.009074f
C123 B.n76 VSUBS 0.009074f
C124 B.n77 VSUBS 0.009074f
C125 B.n78 VSUBS 0.009074f
C126 B.n79 VSUBS 0.009074f
C127 B.n80 VSUBS 0.009074f
C128 B.n81 VSUBS 0.009074f
C129 B.n82 VSUBS 0.009074f
C130 B.n83 VSUBS 0.00854f
C131 B.n84 VSUBS 0.009074f
C132 B.n85 VSUBS 0.009074f
C133 B.n86 VSUBS 0.009074f
C134 B.n87 VSUBS 0.009074f
C135 B.n88 VSUBS 0.009074f
C136 B.t11 VSUBS 0.180427f
C137 B.t10 VSUBS 0.199125f
C138 B.t9 VSUBS 0.532568f
C139 B.n89 VSUBS 0.123551f
C140 B.n90 VSUBS 0.086529f
C141 B.n91 VSUBS 0.009074f
C142 B.n92 VSUBS 0.009074f
C143 B.n93 VSUBS 0.009074f
C144 B.n94 VSUBS 0.009074f
C145 B.n95 VSUBS 0.009074f
C146 B.n96 VSUBS 0.009074f
C147 B.n97 VSUBS 0.009074f
C148 B.n98 VSUBS 0.009074f
C149 B.n99 VSUBS 0.009074f
C150 B.n100 VSUBS 0.009074f
C151 B.n101 VSUBS 0.019626f
C152 B.n102 VSUBS 0.009074f
C153 B.n103 VSUBS 0.009074f
C154 B.n104 VSUBS 0.009074f
C155 B.n105 VSUBS 0.009074f
C156 B.n106 VSUBS 0.009074f
C157 B.n107 VSUBS 0.009074f
C158 B.n108 VSUBS 0.009074f
C159 B.n109 VSUBS 0.009074f
C160 B.n110 VSUBS 0.009074f
C161 B.n111 VSUBS 0.009074f
C162 B.n112 VSUBS 0.009074f
C163 B.n113 VSUBS 0.009074f
C164 B.n114 VSUBS 0.009074f
C165 B.n115 VSUBS 0.009074f
C166 B.n116 VSUBS 0.009074f
C167 B.n117 VSUBS 0.009074f
C168 B.n118 VSUBS 0.009074f
C169 B.n119 VSUBS 0.009074f
C170 B.n120 VSUBS 0.009074f
C171 B.n121 VSUBS 0.009074f
C172 B.n122 VSUBS 0.009074f
C173 B.n123 VSUBS 0.009074f
C174 B.n124 VSUBS 0.009074f
C175 B.n125 VSUBS 0.009074f
C176 B.n126 VSUBS 0.009074f
C177 B.n127 VSUBS 0.009074f
C178 B.n128 VSUBS 0.009074f
C179 B.n129 VSUBS 0.009074f
C180 B.n130 VSUBS 0.009074f
C181 B.n131 VSUBS 0.009074f
C182 B.n132 VSUBS 0.009074f
C183 B.n133 VSUBS 0.009074f
C184 B.n134 VSUBS 0.009074f
C185 B.n135 VSUBS 0.009074f
C186 B.n136 VSUBS 0.009074f
C187 B.n137 VSUBS 0.009074f
C188 B.n138 VSUBS 0.009074f
C189 B.n139 VSUBS 0.009074f
C190 B.n140 VSUBS 0.009074f
C191 B.n141 VSUBS 0.009074f
C192 B.n142 VSUBS 0.009074f
C193 B.n143 VSUBS 0.009074f
C194 B.n144 VSUBS 0.009074f
C195 B.n145 VSUBS 0.009074f
C196 B.n146 VSUBS 0.009074f
C197 B.n147 VSUBS 0.009074f
C198 B.n148 VSUBS 0.009074f
C199 B.n149 VSUBS 0.009074f
C200 B.n150 VSUBS 0.019626f
C201 B.n151 VSUBS 0.021209f
C202 B.n152 VSUBS 0.021209f
C203 B.n153 VSUBS 0.009074f
C204 B.n154 VSUBS 0.009074f
C205 B.n155 VSUBS 0.009074f
C206 B.n156 VSUBS 0.009074f
C207 B.n157 VSUBS 0.009074f
C208 B.n158 VSUBS 0.009074f
C209 B.n159 VSUBS 0.009074f
C210 B.n160 VSUBS 0.009074f
C211 B.n161 VSUBS 0.009074f
C212 B.n162 VSUBS 0.009074f
C213 B.n163 VSUBS 0.009074f
C214 B.n164 VSUBS 0.009074f
C215 B.n165 VSUBS 0.009074f
C216 B.n166 VSUBS 0.009074f
C217 B.n167 VSUBS 0.009074f
C218 B.n168 VSUBS 0.009074f
C219 B.n169 VSUBS 0.009074f
C220 B.n170 VSUBS 0.009074f
C221 B.n171 VSUBS 0.009074f
C222 B.n172 VSUBS 0.009074f
C223 B.n173 VSUBS 0.009074f
C224 B.n174 VSUBS 0.009074f
C225 B.n175 VSUBS 0.009074f
C226 B.n176 VSUBS 0.009074f
C227 B.n177 VSUBS 0.009074f
C228 B.n178 VSUBS 0.009074f
C229 B.n179 VSUBS 0.009074f
C230 B.n180 VSUBS 0.009074f
C231 B.n181 VSUBS 0.009074f
C232 B.n182 VSUBS 0.00854f
C233 B.n183 VSUBS 0.021024f
C234 B.n184 VSUBS 0.005071f
C235 B.n185 VSUBS 0.009074f
C236 B.n186 VSUBS 0.009074f
C237 B.n187 VSUBS 0.009074f
C238 B.n188 VSUBS 0.009074f
C239 B.n189 VSUBS 0.009074f
C240 B.n190 VSUBS 0.009074f
C241 B.n191 VSUBS 0.009074f
C242 B.n192 VSUBS 0.009074f
C243 B.n193 VSUBS 0.009074f
C244 B.n194 VSUBS 0.009074f
C245 B.n195 VSUBS 0.009074f
C246 B.n196 VSUBS 0.009074f
C247 B.t8 VSUBS 0.180427f
C248 B.t7 VSUBS 0.199124f
C249 B.t6 VSUBS 0.532568f
C250 B.n197 VSUBS 0.123551f
C251 B.n198 VSUBS 0.086529f
C252 B.n199 VSUBS 0.021024f
C253 B.n200 VSUBS 0.005071f
C254 B.n201 VSUBS 0.009074f
C255 B.n202 VSUBS 0.009074f
C256 B.n203 VSUBS 0.009074f
C257 B.n204 VSUBS 0.009074f
C258 B.n205 VSUBS 0.009074f
C259 B.n206 VSUBS 0.009074f
C260 B.n207 VSUBS 0.009074f
C261 B.n208 VSUBS 0.009074f
C262 B.n209 VSUBS 0.009074f
C263 B.n210 VSUBS 0.009074f
C264 B.n211 VSUBS 0.009074f
C265 B.n212 VSUBS 0.009074f
C266 B.n213 VSUBS 0.009074f
C267 B.n214 VSUBS 0.009074f
C268 B.n215 VSUBS 0.009074f
C269 B.n216 VSUBS 0.009074f
C270 B.n217 VSUBS 0.009074f
C271 B.n218 VSUBS 0.009074f
C272 B.n219 VSUBS 0.009074f
C273 B.n220 VSUBS 0.009074f
C274 B.n221 VSUBS 0.009074f
C275 B.n222 VSUBS 0.009074f
C276 B.n223 VSUBS 0.009074f
C277 B.n224 VSUBS 0.009074f
C278 B.n225 VSUBS 0.009074f
C279 B.n226 VSUBS 0.009074f
C280 B.n227 VSUBS 0.009074f
C281 B.n228 VSUBS 0.009074f
C282 B.n229 VSUBS 0.009074f
C283 B.n230 VSUBS 0.009074f
C284 B.n231 VSUBS 0.009074f
C285 B.n232 VSUBS 0.021209f
C286 B.n233 VSUBS 0.019626f
C287 B.n234 VSUBS 0.020764f
C288 B.n235 VSUBS 0.009074f
C289 B.n236 VSUBS 0.009074f
C290 B.n237 VSUBS 0.009074f
C291 B.n238 VSUBS 0.009074f
C292 B.n239 VSUBS 0.009074f
C293 B.n240 VSUBS 0.009074f
C294 B.n241 VSUBS 0.009074f
C295 B.n242 VSUBS 0.009074f
C296 B.n243 VSUBS 0.009074f
C297 B.n244 VSUBS 0.009074f
C298 B.n245 VSUBS 0.009074f
C299 B.n246 VSUBS 0.009074f
C300 B.n247 VSUBS 0.009074f
C301 B.n248 VSUBS 0.009074f
C302 B.n249 VSUBS 0.009074f
C303 B.n250 VSUBS 0.009074f
C304 B.n251 VSUBS 0.009074f
C305 B.n252 VSUBS 0.009074f
C306 B.n253 VSUBS 0.009074f
C307 B.n254 VSUBS 0.009074f
C308 B.n255 VSUBS 0.009074f
C309 B.n256 VSUBS 0.009074f
C310 B.n257 VSUBS 0.009074f
C311 B.n258 VSUBS 0.009074f
C312 B.n259 VSUBS 0.009074f
C313 B.n260 VSUBS 0.009074f
C314 B.n261 VSUBS 0.009074f
C315 B.n262 VSUBS 0.009074f
C316 B.n263 VSUBS 0.009074f
C317 B.n264 VSUBS 0.009074f
C318 B.n265 VSUBS 0.009074f
C319 B.n266 VSUBS 0.009074f
C320 B.n267 VSUBS 0.009074f
C321 B.n268 VSUBS 0.009074f
C322 B.n269 VSUBS 0.009074f
C323 B.n270 VSUBS 0.009074f
C324 B.n271 VSUBS 0.009074f
C325 B.n272 VSUBS 0.009074f
C326 B.n273 VSUBS 0.009074f
C327 B.n274 VSUBS 0.009074f
C328 B.n275 VSUBS 0.009074f
C329 B.n276 VSUBS 0.009074f
C330 B.n277 VSUBS 0.009074f
C331 B.n278 VSUBS 0.009074f
C332 B.n279 VSUBS 0.009074f
C333 B.n280 VSUBS 0.009074f
C334 B.n281 VSUBS 0.009074f
C335 B.n282 VSUBS 0.009074f
C336 B.n283 VSUBS 0.009074f
C337 B.n284 VSUBS 0.009074f
C338 B.n285 VSUBS 0.009074f
C339 B.n286 VSUBS 0.009074f
C340 B.n287 VSUBS 0.009074f
C341 B.n288 VSUBS 0.009074f
C342 B.n289 VSUBS 0.009074f
C343 B.n290 VSUBS 0.009074f
C344 B.n291 VSUBS 0.009074f
C345 B.n292 VSUBS 0.009074f
C346 B.n293 VSUBS 0.009074f
C347 B.n294 VSUBS 0.009074f
C348 B.n295 VSUBS 0.009074f
C349 B.n296 VSUBS 0.009074f
C350 B.n297 VSUBS 0.009074f
C351 B.n298 VSUBS 0.009074f
C352 B.n299 VSUBS 0.009074f
C353 B.n300 VSUBS 0.009074f
C354 B.n301 VSUBS 0.009074f
C355 B.n302 VSUBS 0.009074f
C356 B.n303 VSUBS 0.009074f
C357 B.n304 VSUBS 0.009074f
C358 B.n305 VSUBS 0.009074f
C359 B.n306 VSUBS 0.009074f
C360 B.n307 VSUBS 0.009074f
C361 B.n308 VSUBS 0.009074f
C362 B.n309 VSUBS 0.009074f
C363 B.n310 VSUBS 0.009074f
C364 B.n311 VSUBS 0.009074f
C365 B.n312 VSUBS 0.009074f
C366 B.n313 VSUBS 0.019626f
C367 B.n314 VSUBS 0.021209f
C368 B.n315 VSUBS 0.021209f
C369 B.n316 VSUBS 0.009074f
C370 B.n317 VSUBS 0.009074f
C371 B.n318 VSUBS 0.009074f
C372 B.n319 VSUBS 0.009074f
C373 B.n320 VSUBS 0.009074f
C374 B.n321 VSUBS 0.009074f
C375 B.n322 VSUBS 0.009074f
C376 B.n323 VSUBS 0.009074f
C377 B.n324 VSUBS 0.009074f
C378 B.n325 VSUBS 0.009074f
C379 B.n326 VSUBS 0.009074f
C380 B.n327 VSUBS 0.009074f
C381 B.n328 VSUBS 0.009074f
C382 B.n329 VSUBS 0.009074f
C383 B.n330 VSUBS 0.009074f
C384 B.n331 VSUBS 0.009074f
C385 B.n332 VSUBS 0.009074f
C386 B.n333 VSUBS 0.009074f
C387 B.n334 VSUBS 0.009074f
C388 B.n335 VSUBS 0.009074f
C389 B.n336 VSUBS 0.009074f
C390 B.n337 VSUBS 0.009074f
C391 B.n338 VSUBS 0.009074f
C392 B.n339 VSUBS 0.009074f
C393 B.n340 VSUBS 0.009074f
C394 B.n341 VSUBS 0.009074f
C395 B.n342 VSUBS 0.009074f
C396 B.n343 VSUBS 0.009074f
C397 B.n344 VSUBS 0.00854f
C398 B.n345 VSUBS 0.009074f
C399 B.n346 VSUBS 0.009074f
C400 B.n347 VSUBS 0.009074f
C401 B.n348 VSUBS 0.009074f
C402 B.n349 VSUBS 0.009074f
C403 B.n350 VSUBS 0.009074f
C404 B.n351 VSUBS 0.009074f
C405 B.n352 VSUBS 0.009074f
C406 B.n353 VSUBS 0.009074f
C407 B.n354 VSUBS 0.009074f
C408 B.n355 VSUBS 0.009074f
C409 B.n356 VSUBS 0.009074f
C410 B.n357 VSUBS 0.009074f
C411 B.n358 VSUBS 0.009074f
C412 B.n359 VSUBS 0.009074f
C413 B.n360 VSUBS 0.005071f
C414 B.n361 VSUBS 0.021024f
C415 B.n362 VSUBS 0.00854f
C416 B.n363 VSUBS 0.009074f
C417 B.n364 VSUBS 0.009074f
C418 B.n365 VSUBS 0.009074f
C419 B.n366 VSUBS 0.009074f
C420 B.n367 VSUBS 0.009074f
C421 B.n368 VSUBS 0.009074f
C422 B.n369 VSUBS 0.009074f
C423 B.n370 VSUBS 0.009074f
C424 B.n371 VSUBS 0.009074f
C425 B.n372 VSUBS 0.009074f
C426 B.n373 VSUBS 0.009074f
C427 B.n374 VSUBS 0.009074f
C428 B.n375 VSUBS 0.009074f
C429 B.n376 VSUBS 0.009074f
C430 B.n377 VSUBS 0.009074f
C431 B.n378 VSUBS 0.009074f
C432 B.n379 VSUBS 0.009074f
C433 B.n380 VSUBS 0.009074f
C434 B.n381 VSUBS 0.009074f
C435 B.n382 VSUBS 0.009074f
C436 B.n383 VSUBS 0.009074f
C437 B.n384 VSUBS 0.009074f
C438 B.n385 VSUBS 0.009074f
C439 B.n386 VSUBS 0.009074f
C440 B.n387 VSUBS 0.009074f
C441 B.n388 VSUBS 0.009074f
C442 B.n389 VSUBS 0.009074f
C443 B.n390 VSUBS 0.009074f
C444 B.n391 VSUBS 0.009074f
C445 B.n392 VSUBS 0.021209f
C446 B.n393 VSUBS 0.019626f
C447 B.n394 VSUBS 0.019626f
C448 B.n395 VSUBS 0.009074f
C449 B.n396 VSUBS 0.009074f
C450 B.n397 VSUBS 0.009074f
C451 B.n398 VSUBS 0.009074f
C452 B.n399 VSUBS 0.009074f
C453 B.n400 VSUBS 0.009074f
C454 B.n401 VSUBS 0.009074f
C455 B.n402 VSUBS 0.009074f
C456 B.n403 VSUBS 0.009074f
C457 B.n404 VSUBS 0.009074f
C458 B.n405 VSUBS 0.009074f
C459 B.n406 VSUBS 0.009074f
C460 B.n407 VSUBS 0.009074f
C461 B.n408 VSUBS 0.009074f
C462 B.n409 VSUBS 0.009074f
C463 B.n410 VSUBS 0.009074f
C464 B.n411 VSUBS 0.009074f
C465 B.n412 VSUBS 0.009074f
C466 B.n413 VSUBS 0.009074f
C467 B.n414 VSUBS 0.009074f
C468 B.n415 VSUBS 0.009074f
C469 B.n416 VSUBS 0.009074f
C470 B.n417 VSUBS 0.009074f
C471 B.n418 VSUBS 0.009074f
C472 B.n419 VSUBS 0.009074f
C473 B.n420 VSUBS 0.009074f
C474 B.n421 VSUBS 0.009074f
C475 B.n422 VSUBS 0.009074f
C476 B.n423 VSUBS 0.009074f
C477 B.n424 VSUBS 0.009074f
C478 B.n425 VSUBS 0.009074f
C479 B.n426 VSUBS 0.009074f
C480 B.n427 VSUBS 0.009074f
C481 B.n428 VSUBS 0.009074f
C482 B.n429 VSUBS 0.009074f
C483 B.n430 VSUBS 0.009074f
C484 B.n431 VSUBS 0.011842f
C485 B.n432 VSUBS 0.012614f
C486 B.n433 VSUBS 0.025084f
C487 VTAIL.t3 VSUBS 0.841059f
C488 VTAIL.n0 VSUBS 0.647335f
C489 VTAIL.t6 VSUBS 0.841059f
C490 VTAIL.n1 VSUBS 0.722087f
C491 VTAIL.t7 VSUBS 0.841059f
C492 VTAIL.n2 VSUBS 1.5958f
C493 VTAIL.t1 VSUBS 0.841063f
C494 VTAIL.n3 VSUBS 1.59579f
C495 VTAIL.t2 VSUBS 0.841063f
C496 VTAIL.n4 VSUBS 0.722082f
C497 VTAIL.t5 VSUBS 0.841063f
C498 VTAIL.n5 VSUBS 0.722082f
C499 VTAIL.t4 VSUBS 0.841059f
C500 VTAIL.n6 VSUBS 1.5958f
C501 VTAIL.t0 VSUBS 0.841059f
C502 VTAIL.n7 VSUBS 1.51072f
C503 VDD1.t2 VSUBS 0.109107f
C504 VDD1.t0 VSUBS 0.109107f
C505 VDD1.n0 VSUBS 0.686228f
C506 VDD1.t1 VSUBS 0.109107f
C507 VDD1.t3 VSUBS 0.109107f
C508 VDD1.n1 VSUBS 1.04828f
C509 VP.n0 VSUBS 0.053028f
C510 VP.t1 VSUBS 1.21797f
C511 VP.n1 VSUBS 0.042868f
C512 VP.n2 VSUBS 0.053028f
C513 VP.t0 VSUBS 1.21797f
C514 VP.t2 VSUBS 1.47199f
C515 VP.t3 VSUBS 1.46897f
C516 VP.n3 VSUBS 2.84811f
C517 VP.n4 VSUBS 2.3736f
C518 VP.n5 VSUBS 0.596837f
C519 VP.n6 VSUBS 0.054427f
C520 VP.n7 VSUBS 0.105393f
C521 VP.n8 VSUBS 0.053028f
C522 VP.n9 VSUBS 0.053028f
C523 VP.n10 VSUBS 0.053028f
C524 VP.n11 VSUBS 0.105393f
C525 VP.n12 VSUBS 0.054427f
C526 VP.n13 VSUBS 0.596837f
C527 VP.n14 VSUBS 0.056692f
.ends

