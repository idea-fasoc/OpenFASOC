* NGSPICE file created from diff_pair_sample_0844.ext - technology: sky130A

.subckt diff_pair_sample_0844 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t8 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=2.95185 ps=18.22 w=17.89 l=3.78
X1 VTAIL.t1 VN.t0 VDD2.t5 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=2.95185 ps=18.22 w=17.89 l=3.78
X2 VTAIL.t10 VP.t1 VDD1.t4 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=2.95185 ps=18.22 w=17.89 l=3.78
X3 VDD1.t3 VP.t2 VTAIL.t11 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=2.95185 ps=18.22 w=17.89 l=3.78
X4 VDD2.t4 VN.t1 VTAIL.t5 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=6.9771 ps=36.56 w=17.89 l=3.78
X5 VDD2.t3 VN.t2 VTAIL.t4 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=2.95185 ps=18.22 w=17.89 l=3.78
X6 B.t11 B.t9 B.t10 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=0 ps=0 w=17.89 l=3.78
X7 B.t8 B.t6 B.t7 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=0 ps=0 w=17.89 l=3.78
X8 B.t5 B.t3 B.t4 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=0 ps=0 w=17.89 l=3.78
X9 VDD2.t2 VN.t3 VTAIL.t0 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=2.95185 ps=18.22 w=17.89 l=3.78
X10 VTAIL.t9 VP.t3 VDD1.t2 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=2.95185 ps=18.22 w=17.89 l=3.78
X11 VDD1.t1 VP.t4 VTAIL.t6 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=6.9771 ps=36.56 w=17.89 l=3.78
X12 VTAIL.t3 VN.t4 VDD2.t1 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=2.95185 ps=18.22 w=17.89 l=3.78
X13 B.t2 B.t0 B.t1 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=6.9771 pd=36.56 as=0 ps=0 w=17.89 l=3.78
X14 VDD2.t0 VN.t5 VTAIL.t2 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=6.9771 ps=36.56 w=17.89 l=3.78
X15 VDD1.t0 VP.t5 VTAIL.t7 w_n4258_n4546# sky130_fd_pr__pfet_01v8 ad=2.95185 pd=18.22 as=6.9771 ps=36.56 w=17.89 l=3.78
R0 VP.n16 VP.n13 161.3
R1 VP.n18 VP.n17 161.3
R2 VP.n19 VP.n12 161.3
R3 VP.n21 VP.n20 161.3
R4 VP.n22 VP.n11 161.3
R5 VP.n24 VP.n23 161.3
R6 VP.n25 VP.n10 161.3
R7 VP.n27 VP.n26 161.3
R8 VP.n56 VP.n55 161.3
R9 VP.n54 VP.n1 161.3
R10 VP.n53 VP.n52 161.3
R11 VP.n51 VP.n2 161.3
R12 VP.n50 VP.n49 161.3
R13 VP.n48 VP.n3 161.3
R14 VP.n47 VP.n46 161.3
R15 VP.n45 VP.n4 161.3
R16 VP.n44 VP.n43 161.3
R17 VP.n42 VP.n5 161.3
R18 VP.n41 VP.n40 161.3
R19 VP.n39 VP.n6 161.3
R20 VP.n38 VP.n37 161.3
R21 VP.n36 VP.n7 161.3
R22 VP.n35 VP.n34 161.3
R23 VP.n33 VP.n8 161.3
R24 VP.n32 VP.n31 161.3
R25 VP.n15 VP.t0 147.559
R26 VP.n43 VP.t1 114.061
R27 VP.n30 VP.t2 114.061
R28 VP.n0 VP.t5 114.061
R29 VP.n14 VP.t3 114.061
R30 VP.n9 VP.t4 114.061
R31 VP.n30 VP.n29 84.6847
R32 VP.n57 VP.n0 84.6847
R33 VP.n28 VP.n9 84.6847
R34 VP.n29 VP.n28 57.8516
R35 VP.n15 VP.n14 50.4867
R36 VP.n37 VP.n36 45.8354
R37 VP.n49 VP.n2 45.8354
R38 VP.n20 VP.n11 45.8354
R39 VP.n37 VP.n6 35.1514
R40 VP.n49 VP.n48 35.1514
R41 VP.n20 VP.n19 35.1514
R42 VP.n31 VP.n8 24.4675
R43 VP.n35 VP.n8 24.4675
R44 VP.n36 VP.n35 24.4675
R45 VP.n41 VP.n6 24.4675
R46 VP.n42 VP.n41 24.4675
R47 VP.n43 VP.n42 24.4675
R48 VP.n43 VP.n4 24.4675
R49 VP.n47 VP.n4 24.4675
R50 VP.n48 VP.n47 24.4675
R51 VP.n53 VP.n2 24.4675
R52 VP.n54 VP.n53 24.4675
R53 VP.n55 VP.n54 24.4675
R54 VP.n24 VP.n11 24.4675
R55 VP.n25 VP.n24 24.4675
R56 VP.n26 VP.n25 24.4675
R57 VP.n14 VP.n13 24.4675
R58 VP.n18 VP.n13 24.4675
R59 VP.n19 VP.n18 24.4675
R60 VP.n31 VP.n30 5.38324
R61 VP.n55 VP.n0 5.38324
R62 VP.n26 VP.n9 5.38324
R63 VP.n16 VP.n15 2.4101
R64 VP.n28 VP.n27 0.354971
R65 VP.n32 VP.n29 0.354971
R66 VP.n57 VP.n56 0.354971
R67 VP VP.n57 0.26696
R68 VP.n17 VP.n16 0.189894
R69 VP.n17 VP.n12 0.189894
R70 VP.n21 VP.n12 0.189894
R71 VP.n22 VP.n21 0.189894
R72 VP.n23 VP.n22 0.189894
R73 VP.n23 VP.n10 0.189894
R74 VP.n27 VP.n10 0.189894
R75 VP.n33 VP.n32 0.189894
R76 VP.n34 VP.n33 0.189894
R77 VP.n34 VP.n7 0.189894
R78 VP.n38 VP.n7 0.189894
R79 VP.n39 VP.n38 0.189894
R80 VP.n40 VP.n39 0.189894
R81 VP.n40 VP.n5 0.189894
R82 VP.n44 VP.n5 0.189894
R83 VP.n45 VP.n44 0.189894
R84 VP.n46 VP.n45 0.189894
R85 VP.n46 VP.n3 0.189894
R86 VP.n50 VP.n3 0.189894
R87 VP.n51 VP.n50 0.189894
R88 VP.n52 VP.n51 0.189894
R89 VP.n52 VP.n1 0.189894
R90 VP.n56 VP.n1 0.189894
R91 VTAIL.n7 VTAIL.t5 54.1828
R92 VTAIL.n11 VTAIL.t2 54.1825
R93 VTAIL.n2 VTAIL.t7 54.1825
R94 VTAIL.n10 VTAIL.t6 54.1825
R95 VTAIL.n9 VTAIL.n8 52.3658
R96 VTAIL.n6 VTAIL.n5 52.3658
R97 VTAIL.n1 VTAIL.n0 52.3656
R98 VTAIL.n4 VTAIL.n3 52.3656
R99 VTAIL.n6 VTAIL.n4 34.8755
R100 VTAIL.n11 VTAIL.n10 31.3324
R101 VTAIL.n7 VTAIL.n6 3.5436
R102 VTAIL.n10 VTAIL.n9 3.5436
R103 VTAIL.n4 VTAIL.n2 3.5436
R104 VTAIL VTAIL.n11 2.59964
R105 VTAIL.n9 VTAIL.n7 2.24188
R106 VTAIL.n2 VTAIL.n1 2.24188
R107 VTAIL.n0 VTAIL.t0 1.81744
R108 VTAIL.n0 VTAIL.t1 1.81744
R109 VTAIL.n3 VTAIL.t11 1.81744
R110 VTAIL.n3 VTAIL.t10 1.81744
R111 VTAIL.n8 VTAIL.t8 1.81744
R112 VTAIL.n8 VTAIL.t9 1.81744
R113 VTAIL.n5 VTAIL.t4 1.81744
R114 VTAIL.n5 VTAIL.t3 1.81744
R115 VTAIL VTAIL.n1 0.944465
R116 VDD1 VDD1.t5 73.5771
R117 VDD1.n1 VDD1.t3 73.4633
R118 VDD1.n1 VDD1.n0 69.8748
R119 VDD1.n3 VDD1.n2 69.0444
R120 VDD1.n3 VDD1.n1 53.0074
R121 VDD1.n2 VDD1.t2 1.81744
R122 VDD1.n2 VDD1.t1 1.81744
R123 VDD1.n0 VDD1.t4 1.81744
R124 VDD1.n0 VDD1.t0 1.81744
R125 VDD1 VDD1.n3 0.828086
R126 VN.n38 VN.n37 161.3
R127 VN.n36 VN.n21 161.3
R128 VN.n35 VN.n34 161.3
R129 VN.n33 VN.n22 161.3
R130 VN.n32 VN.n31 161.3
R131 VN.n30 VN.n23 161.3
R132 VN.n29 VN.n28 161.3
R133 VN.n27 VN.n24 161.3
R134 VN.n18 VN.n17 161.3
R135 VN.n16 VN.n1 161.3
R136 VN.n15 VN.n14 161.3
R137 VN.n13 VN.n2 161.3
R138 VN.n12 VN.n11 161.3
R139 VN.n10 VN.n3 161.3
R140 VN.n9 VN.n8 161.3
R141 VN.n7 VN.n4 161.3
R142 VN.n26 VN.t1 147.56
R143 VN.n6 VN.t3 147.56
R144 VN.n5 VN.t0 114.061
R145 VN.n0 VN.t5 114.061
R146 VN.n25 VN.t4 114.061
R147 VN.n20 VN.t2 114.061
R148 VN.n19 VN.n0 84.6847
R149 VN.n39 VN.n20 84.6847
R150 VN VN.n39 58.017
R151 VN.n26 VN.n25 50.4867
R152 VN.n6 VN.n5 50.4867
R153 VN.n11 VN.n2 45.8354
R154 VN.n31 VN.n22 45.8354
R155 VN.n11 VN.n10 35.1514
R156 VN.n31 VN.n30 35.1514
R157 VN.n5 VN.n4 24.4675
R158 VN.n9 VN.n4 24.4675
R159 VN.n10 VN.n9 24.4675
R160 VN.n15 VN.n2 24.4675
R161 VN.n16 VN.n15 24.4675
R162 VN.n17 VN.n16 24.4675
R163 VN.n30 VN.n29 24.4675
R164 VN.n29 VN.n24 24.4675
R165 VN.n25 VN.n24 24.4675
R166 VN.n37 VN.n36 24.4675
R167 VN.n36 VN.n35 24.4675
R168 VN.n35 VN.n22 24.4675
R169 VN.n17 VN.n0 5.38324
R170 VN.n37 VN.n20 5.38324
R171 VN.n27 VN.n26 2.41011
R172 VN.n7 VN.n6 2.41011
R173 VN.n39 VN.n38 0.354971
R174 VN.n19 VN.n18 0.354971
R175 VN VN.n19 0.26696
R176 VN.n38 VN.n21 0.189894
R177 VN.n34 VN.n21 0.189894
R178 VN.n34 VN.n33 0.189894
R179 VN.n33 VN.n32 0.189894
R180 VN.n32 VN.n23 0.189894
R181 VN.n28 VN.n23 0.189894
R182 VN.n28 VN.n27 0.189894
R183 VN.n8 VN.n7 0.189894
R184 VN.n8 VN.n3 0.189894
R185 VN.n12 VN.n3 0.189894
R186 VN.n13 VN.n12 0.189894
R187 VN.n14 VN.n13 0.189894
R188 VN.n14 VN.n1 0.189894
R189 VN.n18 VN.n1 0.189894
R190 VDD2.n1 VDD2.t2 73.4633
R191 VDD2.n2 VDD2.t3 70.8616
R192 VDD2.n1 VDD2.n0 69.8748
R193 VDD2 VDD2.n3 69.872
R194 VDD2.n2 VDD2.n1 50.6528
R195 VDD2 VDD2.n2 2.71602
R196 VDD2.n3 VDD2.t1 1.81744
R197 VDD2.n3 VDD2.t4 1.81744
R198 VDD2.n0 VDD2.t5 1.81744
R199 VDD2.n0 VDD2.t0 1.81744
R200 B.n524 B.n155 585
R201 B.n523 B.n522 585
R202 B.n521 B.n156 585
R203 B.n520 B.n519 585
R204 B.n518 B.n157 585
R205 B.n517 B.n516 585
R206 B.n515 B.n158 585
R207 B.n514 B.n513 585
R208 B.n512 B.n159 585
R209 B.n511 B.n510 585
R210 B.n509 B.n160 585
R211 B.n508 B.n507 585
R212 B.n506 B.n161 585
R213 B.n505 B.n504 585
R214 B.n503 B.n162 585
R215 B.n502 B.n501 585
R216 B.n500 B.n163 585
R217 B.n499 B.n498 585
R218 B.n497 B.n164 585
R219 B.n496 B.n495 585
R220 B.n494 B.n165 585
R221 B.n493 B.n492 585
R222 B.n491 B.n166 585
R223 B.n490 B.n489 585
R224 B.n488 B.n167 585
R225 B.n487 B.n486 585
R226 B.n485 B.n168 585
R227 B.n484 B.n483 585
R228 B.n482 B.n169 585
R229 B.n481 B.n480 585
R230 B.n479 B.n170 585
R231 B.n478 B.n477 585
R232 B.n476 B.n171 585
R233 B.n475 B.n474 585
R234 B.n473 B.n172 585
R235 B.n472 B.n471 585
R236 B.n470 B.n173 585
R237 B.n469 B.n468 585
R238 B.n467 B.n174 585
R239 B.n466 B.n465 585
R240 B.n464 B.n175 585
R241 B.n463 B.n462 585
R242 B.n461 B.n176 585
R243 B.n460 B.n459 585
R244 B.n458 B.n177 585
R245 B.n457 B.n456 585
R246 B.n455 B.n178 585
R247 B.n454 B.n453 585
R248 B.n452 B.n179 585
R249 B.n451 B.n450 585
R250 B.n449 B.n180 585
R251 B.n448 B.n447 585
R252 B.n446 B.n181 585
R253 B.n445 B.n444 585
R254 B.n443 B.n182 585
R255 B.n442 B.n441 585
R256 B.n440 B.n183 585
R257 B.n439 B.n438 585
R258 B.n437 B.n184 585
R259 B.n436 B.n435 585
R260 B.n431 B.n185 585
R261 B.n430 B.n429 585
R262 B.n428 B.n186 585
R263 B.n427 B.n426 585
R264 B.n425 B.n187 585
R265 B.n424 B.n423 585
R266 B.n422 B.n188 585
R267 B.n421 B.n420 585
R268 B.n418 B.n189 585
R269 B.n417 B.n416 585
R270 B.n415 B.n192 585
R271 B.n414 B.n413 585
R272 B.n412 B.n193 585
R273 B.n411 B.n410 585
R274 B.n409 B.n194 585
R275 B.n408 B.n407 585
R276 B.n406 B.n195 585
R277 B.n405 B.n404 585
R278 B.n403 B.n196 585
R279 B.n402 B.n401 585
R280 B.n400 B.n197 585
R281 B.n399 B.n398 585
R282 B.n397 B.n198 585
R283 B.n396 B.n395 585
R284 B.n394 B.n199 585
R285 B.n393 B.n392 585
R286 B.n391 B.n200 585
R287 B.n390 B.n389 585
R288 B.n388 B.n201 585
R289 B.n387 B.n386 585
R290 B.n385 B.n202 585
R291 B.n384 B.n383 585
R292 B.n382 B.n203 585
R293 B.n381 B.n380 585
R294 B.n379 B.n204 585
R295 B.n378 B.n377 585
R296 B.n376 B.n205 585
R297 B.n375 B.n374 585
R298 B.n373 B.n206 585
R299 B.n372 B.n371 585
R300 B.n370 B.n207 585
R301 B.n369 B.n368 585
R302 B.n367 B.n208 585
R303 B.n366 B.n365 585
R304 B.n364 B.n209 585
R305 B.n363 B.n362 585
R306 B.n361 B.n210 585
R307 B.n360 B.n359 585
R308 B.n358 B.n211 585
R309 B.n357 B.n356 585
R310 B.n355 B.n212 585
R311 B.n354 B.n353 585
R312 B.n352 B.n213 585
R313 B.n351 B.n350 585
R314 B.n349 B.n214 585
R315 B.n348 B.n347 585
R316 B.n346 B.n215 585
R317 B.n345 B.n344 585
R318 B.n343 B.n216 585
R319 B.n342 B.n341 585
R320 B.n340 B.n217 585
R321 B.n339 B.n338 585
R322 B.n337 B.n218 585
R323 B.n336 B.n335 585
R324 B.n334 B.n219 585
R325 B.n333 B.n332 585
R326 B.n331 B.n220 585
R327 B.n526 B.n525 585
R328 B.n527 B.n154 585
R329 B.n529 B.n528 585
R330 B.n530 B.n153 585
R331 B.n532 B.n531 585
R332 B.n533 B.n152 585
R333 B.n535 B.n534 585
R334 B.n536 B.n151 585
R335 B.n538 B.n537 585
R336 B.n539 B.n150 585
R337 B.n541 B.n540 585
R338 B.n542 B.n149 585
R339 B.n544 B.n543 585
R340 B.n545 B.n148 585
R341 B.n547 B.n546 585
R342 B.n548 B.n147 585
R343 B.n550 B.n549 585
R344 B.n551 B.n146 585
R345 B.n553 B.n552 585
R346 B.n554 B.n145 585
R347 B.n556 B.n555 585
R348 B.n557 B.n144 585
R349 B.n559 B.n558 585
R350 B.n560 B.n143 585
R351 B.n562 B.n561 585
R352 B.n563 B.n142 585
R353 B.n565 B.n564 585
R354 B.n566 B.n141 585
R355 B.n568 B.n567 585
R356 B.n569 B.n140 585
R357 B.n571 B.n570 585
R358 B.n572 B.n139 585
R359 B.n574 B.n573 585
R360 B.n575 B.n138 585
R361 B.n577 B.n576 585
R362 B.n578 B.n137 585
R363 B.n580 B.n579 585
R364 B.n581 B.n136 585
R365 B.n583 B.n582 585
R366 B.n584 B.n135 585
R367 B.n586 B.n585 585
R368 B.n587 B.n134 585
R369 B.n589 B.n588 585
R370 B.n590 B.n133 585
R371 B.n592 B.n591 585
R372 B.n593 B.n132 585
R373 B.n595 B.n594 585
R374 B.n596 B.n131 585
R375 B.n598 B.n597 585
R376 B.n599 B.n130 585
R377 B.n601 B.n600 585
R378 B.n602 B.n129 585
R379 B.n604 B.n603 585
R380 B.n605 B.n128 585
R381 B.n607 B.n606 585
R382 B.n608 B.n127 585
R383 B.n610 B.n609 585
R384 B.n611 B.n126 585
R385 B.n613 B.n612 585
R386 B.n614 B.n125 585
R387 B.n616 B.n615 585
R388 B.n617 B.n124 585
R389 B.n619 B.n618 585
R390 B.n620 B.n123 585
R391 B.n622 B.n621 585
R392 B.n623 B.n122 585
R393 B.n625 B.n624 585
R394 B.n626 B.n121 585
R395 B.n628 B.n627 585
R396 B.n629 B.n120 585
R397 B.n631 B.n630 585
R398 B.n632 B.n119 585
R399 B.n634 B.n633 585
R400 B.n635 B.n118 585
R401 B.n637 B.n636 585
R402 B.n638 B.n117 585
R403 B.n640 B.n639 585
R404 B.n641 B.n116 585
R405 B.n643 B.n642 585
R406 B.n644 B.n115 585
R407 B.n646 B.n645 585
R408 B.n647 B.n114 585
R409 B.n649 B.n648 585
R410 B.n650 B.n113 585
R411 B.n652 B.n651 585
R412 B.n653 B.n112 585
R413 B.n655 B.n654 585
R414 B.n656 B.n111 585
R415 B.n658 B.n657 585
R416 B.n659 B.n110 585
R417 B.n661 B.n660 585
R418 B.n662 B.n109 585
R419 B.n664 B.n663 585
R420 B.n665 B.n108 585
R421 B.n667 B.n666 585
R422 B.n668 B.n107 585
R423 B.n670 B.n669 585
R424 B.n671 B.n106 585
R425 B.n673 B.n672 585
R426 B.n674 B.n105 585
R427 B.n676 B.n675 585
R428 B.n677 B.n104 585
R429 B.n679 B.n678 585
R430 B.n680 B.n103 585
R431 B.n682 B.n681 585
R432 B.n683 B.n102 585
R433 B.n685 B.n684 585
R434 B.n686 B.n101 585
R435 B.n688 B.n687 585
R436 B.n689 B.n100 585
R437 B.n691 B.n690 585
R438 B.n692 B.n99 585
R439 B.n694 B.n693 585
R440 B.n695 B.n98 585
R441 B.n887 B.n30 585
R442 B.n886 B.n885 585
R443 B.n884 B.n31 585
R444 B.n883 B.n882 585
R445 B.n881 B.n32 585
R446 B.n880 B.n879 585
R447 B.n878 B.n33 585
R448 B.n877 B.n876 585
R449 B.n875 B.n34 585
R450 B.n874 B.n873 585
R451 B.n872 B.n35 585
R452 B.n871 B.n870 585
R453 B.n869 B.n36 585
R454 B.n868 B.n867 585
R455 B.n866 B.n37 585
R456 B.n865 B.n864 585
R457 B.n863 B.n38 585
R458 B.n862 B.n861 585
R459 B.n860 B.n39 585
R460 B.n859 B.n858 585
R461 B.n857 B.n40 585
R462 B.n856 B.n855 585
R463 B.n854 B.n41 585
R464 B.n853 B.n852 585
R465 B.n851 B.n42 585
R466 B.n850 B.n849 585
R467 B.n848 B.n43 585
R468 B.n847 B.n846 585
R469 B.n845 B.n44 585
R470 B.n844 B.n843 585
R471 B.n842 B.n45 585
R472 B.n841 B.n840 585
R473 B.n839 B.n46 585
R474 B.n838 B.n837 585
R475 B.n836 B.n47 585
R476 B.n835 B.n834 585
R477 B.n833 B.n48 585
R478 B.n832 B.n831 585
R479 B.n830 B.n49 585
R480 B.n829 B.n828 585
R481 B.n827 B.n50 585
R482 B.n826 B.n825 585
R483 B.n824 B.n51 585
R484 B.n823 B.n822 585
R485 B.n821 B.n52 585
R486 B.n820 B.n819 585
R487 B.n818 B.n53 585
R488 B.n817 B.n816 585
R489 B.n815 B.n54 585
R490 B.n814 B.n813 585
R491 B.n812 B.n55 585
R492 B.n811 B.n810 585
R493 B.n809 B.n56 585
R494 B.n808 B.n807 585
R495 B.n806 B.n57 585
R496 B.n805 B.n804 585
R497 B.n803 B.n58 585
R498 B.n802 B.n801 585
R499 B.n800 B.n59 585
R500 B.n798 B.n797 585
R501 B.n796 B.n62 585
R502 B.n795 B.n794 585
R503 B.n793 B.n63 585
R504 B.n792 B.n791 585
R505 B.n790 B.n64 585
R506 B.n789 B.n788 585
R507 B.n787 B.n65 585
R508 B.n786 B.n785 585
R509 B.n784 B.n783 585
R510 B.n782 B.n69 585
R511 B.n781 B.n780 585
R512 B.n779 B.n70 585
R513 B.n778 B.n777 585
R514 B.n776 B.n71 585
R515 B.n775 B.n774 585
R516 B.n773 B.n72 585
R517 B.n772 B.n771 585
R518 B.n770 B.n73 585
R519 B.n769 B.n768 585
R520 B.n767 B.n74 585
R521 B.n766 B.n765 585
R522 B.n764 B.n75 585
R523 B.n763 B.n762 585
R524 B.n761 B.n76 585
R525 B.n760 B.n759 585
R526 B.n758 B.n77 585
R527 B.n757 B.n756 585
R528 B.n755 B.n78 585
R529 B.n754 B.n753 585
R530 B.n752 B.n79 585
R531 B.n751 B.n750 585
R532 B.n749 B.n80 585
R533 B.n748 B.n747 585
R534 B.n746 B.n81 585
R535 B.n745 B.n744 585
R536 B.n743 B.n82 585
R537 B.n742 B.n741 585
R538 B.n740 B.n83 585
R539 B.n739 B.n738 585
R540 B.n737 B.n84 585
R541 B.n736 B.n735 585
R542 B.n734 B.n85 585
R543 B.n733 B.n732 585
R544 B.n731 B.n86 585
R545 B.n730 B.n729 585
R546 B.n728 B.n87 585
R547 B.n727 B.n726 585
R548 B.n725 B.n88 585
R549 B.n724 B.n723 585
R550 B.n722 B.n89 585
R551 B.n721 B.n720 585
R552 B.n719 B.n90 585
R553 B.n718 B.n717 585
R554 B.n716 B.n91 585
R555 B.n715 B.n714 585
R556 B.n713 B.n92 585
R557 B.n712 B.n711 585
R558 B.n710 B.n93 585
R559 B.n709 B.n708 585
R560 B.n707 B.n94 585
R561 B.n706 B.n705 585
R562 B.n704 B.n95 585
R563 B.n703 B.n702 585
R564 B.n701 B.n96 585
R565 B.n700 B.n699 585
R566 B.n698 B.n97 585
R567 B.n697 B.n696 585
R568 B.n889 B.n888 585
R569 B.n890 B.n29 585
R570 B.n892 B.n891 585
R571 B.n893 B.n28 585
R572 B.n895 B.n894 585
R573 B.n896 B.n27 585
R574 B.n898 B.n897 585
R575 B.n899 B.n26 585
R576 B.n901 B.n900 585
R577 B.n902 B.n25 585
R578 B.n904 B.n903 585
R579 B.n905 B.n24 585
R580 B.n907 B.n906 585
R581 B.n908 B.n23 585
R582 B.n910 B.n909 585
R583 B.n911 B.n22 585
R584 B.n913 B.n912 585
R585 B.n914 B.n21 585
R586 B.n916 B.n915 585
R587 B.n917 B.n20 585
R588 B.n919 B.n918 585
R589 B.n920 B.n19 585
R590 B.n922 B.n921 585
R591 B.n923 B.n18 585
R592 B.n925 B.n924 585
R593 B.n926 B.n17 585
R594 B.n928 B.n927 585
R595 B.n929 B.n16 585
R596 B.n931 B.n930 585
R597 B.n932 B.n15 585
R598 B.n934 B.n933 585
R599 B.n935 B.n14 585
R600 B.n937 B.n936 585
R601 B.n938 B.n13 585
R602 B.n940 B.n939 585
R603 B.n941 B.n12 585
R604 B.n943 B.n942 585
R605 B.n944 B.n11 585
R606 B.n946 B.n945 585
R607 B.n947 B.n10 585
R608 B.n949 B.n948 585
R609 B.n950 B.n9 585
R610 B.n952 B.n951 585
R611 B.n953 B.n8 585
R612 B.n955 B.n954 585
R613 B.n956 B.n7 585
R614 B.n958 B.n957 585
R615 B.n959 B.n6 585
R616 B.n961 B.n960 585
R617 B.n962 B.n5 585
R618 B.n964 B.n963 585
R619 B.n965 B.n4 585
R620 B.n967 B.n966 585
R621 B.n968 B.n3 585
R622 B.n970 B.n969 585
R623 B.n971 B.n0 585
R624 B.n2 B.n1 585
R625 B.n249 B.n248 585
R626 B.n250 B.n247 585
R627 B.n252 B.n251 585
R628 B.n253 B.n246 585
R629 B.n255 B.n254 585
R630 B.n256 B.n245 585
R631 B.n258 B.n257 585
R632 B.n259 B.n244 585
R633 B.n261 B.n260 585
R634 B.n262 B.n243 585
R635 B.n264 B.n263 585
R636 B.n265 B.n242 585
R637 B.n267 B.n266 585
R638 B.n268 B.n241 585
R639 B.n270 B.n269 585
R640 B.n271 B.n240 585
R641 B.n273 B.n272 585
R642 B.n274 B.n239 585
R643 B.n276 B.n275 585
R644 B.n277 B.n238 585
R645 B.n279 B.n278 585
R646 B.n280 B.n237 585
R647 B.n282 B.n281 585
R648 B.n283 B.n236 585
R649 B.n285 B.n284 585
R650 B.n286 B.n235 585
R651 B.n288 B.n287 585
R652 B.n289 B.n234 585
R653 B.n291 B.n290 585
R654 B.n292 B.n233 585
R655 B.n294 B.n293 585
R656 B.n295 B.n232 585
R657 B.n297 B.n296 585
R658 B.n298 B.n231 585
R659 B.n300 B.n299 585
R660 B.n301 B.n230 585
R661 B.n303 B.n302 585
R662 B.n304 B.n229 585
R663 B.n306 B.n305 585
R664 B.n307 B.n228 585
R665 B.n309 B.n308 585
R666 B.n310 B.n227 585
R667 B.n312 B.n311 585
R668 B.n313 B.n226 585
R669 B.n315 B.n314 585
R670 B.n316 B.n225 585
R671 B.n318 B.n317 585
R672 B.n319 B.n224 585
R673 B.n321 B.n320 585
R674 B.n322 B.n223 585
R675 B.n324 B.n323 585
R676 B.n325 B.n222 585
R677 B.n327 B.n326 585
R678 B.n328 B.n221 585
R679 B.n330 B.n329 585
R680 B.n331 B.n330 530.939
R681 B.n526 B.n155 530.939
R682 B.n696 B.n695 530.939
R683 B.n888 B.n887 530.939
R684 B.n190 B.t3 323.389
R685 B.n432 B.t0 323.389
R686 B.n66 B.t6 323.389
R687 B.n60 B.t9 323.389
R688 B.n973 B.n972 256.663
R689 B.n972 B.n971 235.042
R690 B.n972 B.n2 235.042
R691 B.n432 B.t1 189.996
R692 B.n66 B.t8 189.996
R693 B.n190 B.t4 189.974
R694 B.n60 B.t11 189.974
R695 B.n332 B.n331 163.367
R696 B.n332 B.n219 163.367
R697 B.n336 B.n219 163.367
R698 B.n337 B.n336 163.367
R699 B.n338 B.n337 163.367
R700 B.n338 B.n217 163.367
R701 B.n342 B.n217 163.367
R702 B.n343 B.n342 163.367
R703 B.n344 B.n343 163.367
R704 B.n344 B.n215 163.367
R705 B.n348 B.n215 163.367
R706 B.n349 B.n348 163.367
R707 B.n350 B.n349 163.367
R708 B.n350 B.n213 163.367
R709 B.n354 B.n213 163.367
R710 B.n355 B.n354 163.367
R711 B.n356 B.n355 163.367
R712 B.n356 B.n211 163.367
R713 B.n360 B.n211 163.367
R714 B.n361 B.n360 163.367
R715 B.n362 B.n361 163.367
R716 B.n362 B.n209 163.367
R717 B.n366 B.n209 163.367
R718 B.n367 B.n366 163.367
R719 B.n368 B.n367 163.367
R720 B.n368 B.n207 163.367
R721 B.n372 B.n207 163.367
R722 B.n373 B.n372 163.367
R723 B.n374 B.n373 163.367
R724 B.n374 B.n205 163.367
R725 B.n378 B.n205 163.367
R726 B.n379 B.n378 163.367
R727 B.n380 B.n379 163.367
R728 B.n380 B.n203 163.367
R729 B.n384 B.n203 163.367
R730 B.n385 B.n384 163.367
R731 B.n386 B.n385 163.367
R732 B.n386 B.n201 163.367
R733 B.n390 B.n201 163.367
R734 B.n391 B.n390 163.367
R735 B.n392 B.n391 163.367
R736 B.n392 B.n199 163.367
R737 B.n396 B.n199 163.367
R738 B.n397 B.n396 163.367
R739 B.n398 B.n397 163.367
R740 B.n398 B.n197 163.367
R741 B.n402 B.n197 163.367
R742 B.n403 B.n402 163.367
R743 B.n404 B.n403 163.367
R744 B.n404 B.n195 163.367
R745 B.n408 B.n195 163.367
R746 B.n409 B.n408 163.367
R747 B.n410 B.n409 163.367
R748 B.n410 B.n193 163.367
R749 B.n414 B.n193 163.367
R750 B.n415 B.n414 163.367
R751 B.n416 B.n415 163.367
R752 B.n416 B.n189 163.367
R753 B.n421 B.n189 163.367
R754 B.n422 B.n421 163.367
R755 B.n423 B.n422 163.367
R756 B.n423 B.n187 163.367
R757 B.n427 B.n187 163.367
R758 B.n428 B.n427 163.367
R759 B.n429 B.n428 163.367
R760 B.n429 B.n185 163.367
R761 B.n436 B.n185 163.367
R762 B.n437 B.n436 163.367
R763 B.n438 B.n437 163.367
R764 B.n438 B.n183 163.367
R765 B.n442 B.n183 163.367
R766 B.n443 B.n442 163.367
R767 B.n444 B.n443 163.367
R768 B.n444 B.n181 163.367
R769 B.n448 B.n181 163.367
R770 B.n449 B.n448 163.367
R771 B.n450 B.n449 163.367
R772 B.n450 B.n179 163.367
R773 B.n454 B.n179 163.367
R774 B.n455 B.n454 163.367
R775 B.n456 B.n455 163.367
R776 B.n456 B.n177 163.367
R777 B.n460 B.n177 163.367
R778 B.n461 B.n460 163.367
R779 B.n462 B.n461 163.367
R780 B.n462 B.n175 163.367
R781 B.n466 B.n175 163.367
R782 B.n467 B.n466 163.367
R783 B.n468 B.n467 163.367
R784 B.n468 B.n173 163.367
R785 B.n472 B.n173 163.367
R786 B.n473 B.n472 163.367
R787 B.n474 B.n473 163.367
R788 B.n474 B.n171 163.367
R789 B.n478 B.n171 163.367
R790 B.n479 B.n478 163.367
R791 B.n480 B.n479 163.367
R792 B.n480 B.n169 163.367
R793 B.n484 B.n169 163.367
R794 B.n485 B.n484 163.367
R795 B.n486 B.n485 163.367
R796 B.n486 B.n167 163.367
R797 B.n490 B.n167 163.367
R798 B.n491 B.n490 163.367
R799 B.n492 B.n491 163.367
R800 B.n492 B.n165 163.367
R801 B.n496 B.n165 163.367
R802 B.n497 B.n496 163.367
R803 B.n498 B.n497 163.367
R804 B.n498 B.n163 163.367
R805 B.n502 B.n163 163.367
R806 B.n503 B.n502 163.367
R807 B.n504 B.n503 163.367
R808 B.n504 B.n161 163.367
R809 B.n508 B.n161 163.367
R810 B.n509 B.n508 163.367
R811 B.n510 B.n509 163.367
R812 B.n510 B.n159 163.367
R813 B.n514 B.n159 163.367
R814 B.n515 B.n514 163.367
R815 B.n516 B.n515 163.367
R816 B.n516 B.n157 163.367
R817 B.n520 B.n157 163.367
R818 B.n521 B.n520 163.367
R819 B.n522 B.n521 163.367
R820 B.n522 B.n155 163.367
R821 B.n695 B.n694 163.367
R822 B.n694 B.n99 163.367
R823 B.n690 B.n99 163.367
R824 B.n690 B.n689 163.367
R825 B.n689 B.n688 163.367
R826 B.n688 B.n101 163.367
R827 B.n684 B.n101 163.367
R828 B.n684 B.n683 163.367
R829 B.n683 B.n682 163.367
R830 B.n682 B.n103 163.367
R831 B.n678 B.n103 163.367
R832 B.n678 B.n677 163.367
R833 B.n677 B.n676 163.367
R834 B.n676 B.n105 163.367
R835 B.n672 B.n105 163.367
R836 B.n672 B.n671 163.367
R837 B.n671 B.n670 163.367
R838 B.n670 B.n107 163.367
R839 B.n666 B.n107 163.367
R840 B.n666 B.n665 163.367
R841 B.n665 B.n664 163.367
R842 B.n664 B.n109 163.367
R843 B.n660 B.n109 163.367
R844 B.n660 B.n659 163.367
R845 B.n659 B.n658 163.367
R846 B.n658 B.n111 163.367
R847 B.n654 B.n111 163.367
R848 B.n654 B.n653 163.367
R849 B.n653 B.n652 163.367
R850 B.n652 B.n113 163.367
R851 B.n648 B.n113 163.367
R852 B.n648 B.n647 163.367
R853 B.n647 B.n646 163.367
R854 B.n646 B.n115 163.367
R855 B.n642 B.n115 163.367
R856 B.n642 B.n641 163.367
R857 B.n641 B.n640 163.367
R858 B.n640 B.n117 163.367
R859 B.n636 B.n117 163.367
R860 B.n636 B.n635 163.367
R861 B.n635 B.n634 163.367
R862 B.n634 B.n119 163.367
R863 B.n630 B.n119 163.367
R864 B.n630 B.n629 163.367
R865 B.n629 B.n628 163.367
R866 B.n628 B.n121 163.367
R867 B.n624 B.n121 163.367
R868 B.n624 B.n623 163.367
R869 B.n623 B.n622 163.367
R870 B.n622 B.n123 163.367
R871 B.n618 B.n123 163.367
R872 B.n618 B.n617 163.367
R873 B.n617 B.n616 163.367
R874 B.n616 B.n125 163.367
R875 B.n612 B.n125 163.367
R876 B.n612 B.n611 163.367
R877 B.n611 B.n610 163.367
R878 B.n610 B.n127 163.367
R879 B.n606 B.n127 163.367
R880 B.n606 B.n605 163.367
R881 B.n605 B.n604 163.367
R882 B.n604 B.n129 163.367
R883 B.n600 B.n129 163.367
R884 B.n600 B.n599 163.367
R885 B.n599 B.n598 163.367
R886 B.n598 B.n131 163.367
R887 B.n594 B.n131 163.367
R888 B.n594 B.n593 163.367
R889 B.n593 B.n592 163.367
R890 B.n592 B.n133 163.367
R891 B.n588 B.n133 163.367
R892 B.n588 B.n587 163.367
R893 B.n587 B.n586 163.367
R894 B.n586 B.n135 163.367
R895 B.n582 B.n135 163.367
R896 B.n582 B.n581 163.367
R897 B.n581 B.n580 163.367
R898 B.n580 B.n137 163.367
R899 B.n576 B.n137 163.367
R900 B.n576 B.n575 163.367
R901 B.n575 B.n574 163.367
R902 B.n574 B.n139 163.367
R903 B.n570 B.n139 163.367
R904 B.n570 B.n569 163.367
R905 B.n569 B.n568 163.367
R906 B.n568 B.n141 163.367
R907 B.n564 B.n141 163.367
R908 B.n564 B.n563 163.367
R909 B.n563 B.n562 163.367
R910 B.n562 B.n143 163.367
R911 B.n558 B.n143 163.367
R912 B.n558 B.n557 163.367
R913 B.n557 B.n556 163.367
R914 B.n556 B.n145 163.367
R915 B.n552 B.n145 163.367
R916 B.n552 B.n551 163.367
R917 B.n551 B.n550 163.367
R918 B.n550 B.n147 163.367
R919 B.n546 B.n147 163.367
R920 B.n546 B.n545 163.367
R921 B.n545 B.n544 163.367
R922 B.n544 B.n149 163.367
R923 B.n540 B.n149 163.367
R924 B.n540 B.n539 163.367
R925 B.n539 B.n538 163.367
R926 B.n538 B.n151 163.367
R927 B.n534 B.n151 163.367
R928 B.n534 B.n533 163.367
R929 B.n533 B.n532 163.367
R930 B.n532 B.n153 163.367
R931 B.n528 B.n153 163.367
R932 B.n528 B.n527 163.367
R933 B.n527 B.n526 163.367
R934 B.n887 B.n886 163.367
R935 B.n886 B.n31 163.367
R936 B.n882 B.n31 163.367
R937 B.n882 B.n881 163.367
R938 B.n881 B.n880 163.367
R939 B.n880 B.n33 163.367
R940 B.n876 B.n33 163.367
R941 B.n876 B.n875 163.367
R942 B.n875 B.n874 163.367
R943 B.n874 B.n35 163.367
R944 B.n870 B.n35 163.367
R945 B.n870 B.n869 163.367
R946 B.n869 B.n868 163.367
R947 B.n868 B.n37 163.367
R948 B.n864 B.n37 163.367
R949 B.n864 B.n863 163.367
R950 B.n863 B.n862 163.367
R951 B.n862 B.n39 163.367
R952 B.n858 B.n39 163.367
R953 B.n858 B.n857 163.367
R954 B.n857 B.n856 163.367
R955 B.n856 B.n41 163.367
R956 B.n852 B.n41 163.367
R957 B.n852 B.n851 163.367
R958 B.n851 B.n850 163.367
R959 B.n850 B.n43 163.367
R960 B.n846 B.n43 163.367
R961 B.n846 B.n845 163.367
R962 B.n845 B.n844 163.367
R963 B.n844 B.n45 163.367
R964 B.n840 B.n45 163.367
R965 B.n840 B.n839 163.367
R966 B.n839 B.n838 163.367
R967 B.n838 B.n47 163.367
R968 B.n834 B.n47 163.367
R969 B.n834 B.n833 163.367
R970 B.n833 B.n832 163.367
R971 B.n832 B.n49 163.367
R972 B.n828 B.n49 163.367
R973 B.n828 B.n827 163.367
R974 B.n827 B.n826 163.367
R975 B.n826 B.n51 163.367
R976 B.n822 B.n51 163.367
R977 B.n822 B.n821 163.367
R978 B.n821 B.n820 163.367
R979 B.n820 B.n53 163.367
R980 B.n816 B.n53 163.367
R981 B.n816 B.n815 163.367
R982 B.n815 B.n814 163.367
R983 B.n814 B.n55 163.367
R984 B.n810 B.n55 163.367
R985 B.n810 B.n809 163.367
R986 B.n809 B.n808 163.367
R987 B.n808 B.n57 163.367
R988 B.n804 B.n57 163.367
R989 B.n804 B.n803 163.367
R990 B.n803 B.n802 163.367
R991 B.n802 B.n59 163.367
R992 B.n797 B.n59 163.367
R993 B.n797 B.n796 163.367
R994 B.n796 B.n795 163.367
R995 B.n795 B.n63 163.367
R996 B.n791 B.n63 163.367
R997 B.n791 B.n790 163.367
R998 B.n790 B.n789 163.367
R999 B.n789 B.n65 163.367
R1000 B.n785 B.n65 163.367
R1001 B.n785 B.n784 163.367
R1002 B.n784 B.n69 163.367
R1003 B.n780 B.n69 163.367
R1004 B.n780 B.n779 163.367
R1005 B.n779 B.n778 163.367
R1006 B.n778 B.n71 163.367
R1007 B.n774 B.n71 163.367
R1008 B.n774 B.n773 163.367
R1009 B.n773 B.n772 163.367
R1010 B.n772 B.n73 163.367
R1011 B.n768 B.n73 163.367
R1012 B.n768 B.n767 163.367
R1013 B.n767 B.n766 163.367
R1014 B.n766 B.n75 163.367
R1015 B.n762 B.n75 163.367
R1016 B.n762 B.n761 163.367
R1017 B.n761 B.n760 163.367
R1018 B.n760 B.n77 163.367
R1019 B.n756 B.n77 163.367
R1020 B.n756 B.n755 163.367
R1021 B.n755 B.n754 163.367
R1022 B.n754 B.n79 163.367
R1023 B.n750 B.n79 163.367
R1024 B.n750 B.n749 163.367
R1025 B.n749 B.n748 163.367
R1026 B.n748 B.n81 163.367
R1027 B.n744 B.n81 163.367
R1028 B.n744 B.n743 163.367
R1029 B.n743 B.n742 163.367
R1030 B.n742 B.n83 163.367
R1031 B.n738 B.n83 163.367
R1032 B.n738 B.n737 163.367
R1033 B.n737 B.n736 163.367
R1034 B.n736 B.n85 163.367
R1035 B.n732 B.n85 163.367
R1036 B.n732 B.n731 163.367
R1037 B.n731 B.n730 163.367
R1038 B.n730 B.n87 163.367
R1039 B.n726 B.n87 163.367
R1040 B.n726 B.n725 163.367
R1041 B.n725 B.n724 163.367
R1042 B.n724 B.n89 163.367
R1043 B.n720 B.n89 163.367
R1044 B.n720 B.n719 163.367
R1045 B.n719 B.n718 163.367
R1046 B.n718 B.n91 163.367
R1047 B.n714 B.n91 163.367
R1048 B.n714 B.n713 163.367
R1049 B.n713 B.n712 163.367
R1050 B.n712 B.n93 163.367
R1051 B.n708 B.n93 163.367
R1052 B.n708 B.n707 163.367
R1053 B.n707 B.n706 163.367
R1054 B.n706 B.n95 163.367
R1055 B.n702 B.n95 163.367
R1056 B.n702 B.n701 163.367
R1057 B.n701 B.n700 163.367
R1058 B.n700 B.n97 163.367
R1059 B.n696 B.n97 163.367
R1060 B.n888 B.n29 163.367
R1061 B.n892 B.n29 163.367
R1062 B.n893 B.n892 163.367
R1063 B.n894 B.n893 163.367
R1064 B.n894 B.n27 163.367
R1065 B.n898 B.n27 163.367
R1066 B.n899 B.n898 163.367
R1067 B.n900 B.n899 163.367
R1068 B.n900 B.n25 163.367
R1069 B.n904 B.n25 163.367
R1070 B.n905 B.n904 163.367
R1071 B.n906 B.n905 163.367
R1072 B.n906 B.n23 163.367
R1073 B.n910 B.n23 163.367
R1074 B.n911 B.n910 163.367
R1075 B.n912 B.n911 163.367
R1076 B.n912 B.n21 163.367
R1077 B.n916 B.n21 163.367
R1078 B.n917 B.n916 163.367
R1079 B.n918 B.n917 163.367
R1080 B.n918 B.n19 163.367
R1081 B.n922 B.n19 163.367
R1082 B.n923 B.n922 163.367
R1083 B.n924 B.n923 163.367
R1084 B.n924 B.n17 163.367
R1085 B.n928 B.n17 163.367
R1086 B.n929 B.n928 163.367
R1087 B.n930 B.n929 163.367
R1088 B.n930 B.n15 163.367
R1089 B.n934 B.n15 163.367
R1090 B.n935 B.n934 163.367
R1091 B.n936 B.n935 163.367
R1092 B.n936 B.n13 163.367
R1093 B.n940 B.n13 163.367
R1094 B.n941 B.n940 163.367
R1095 B.n942 B.n941 163.367
R1096 B.n942 B.n11 163.367
R1097 B.n946 B.n11 163.367
R1098 B.n947 B.n946 163.367
R1099 B.n948 B.n947 163.367
R1100 B.n948 B.n9 163.367
R1101 B.n952 B.n9 163.367
R1102 B.n953 B.n952 163.367
R1103 B.n954 B.n953 163.367
R1104 B.n954 B.n7 163.367
R1105 B.n958 B.n7 163.367
R1106 B.n959 B.n958 163.367
R1107 B.n960 B.n959 163.367
R1108 B.n960 B.n5 163.367
R1109 B.n964 B.n5 163.367
R1110 B.n965 B.n964 163.367
R1111 B.n966 B.n965 163.367
R1112 B.n966 B.n3 163.367
R1113 B.n970 B.n3 163.367
R1114 B.n971 B.n970 163.367
R1115 B.n248 B.n2 163.367
R1116 B.n248 B.n247 163.367
R1117 B.n252 B.n247 163.367
R1118 B.n253 B.n252 163.367
R1119 B.n254 B.n253 163.367
R1120 B.n254 B.n245 163.367
R1121 B.n258 B.n245 163.367
R1122 B.n259 B.n258 163.367
R1123 B.n260 B.n259 163.367
R1124 B.n260 B.n243 163.367
R1125 B.n264 B.n243 163.367
R1126 B.n265 B.n264 163.367
R1127 B.n266 B.n265 163.367
R1128 B.n266 B.n241 163.367
R1129 B.n270 B.n241 163.367
R1130 B.n271 B.n270 163.367
R1131 B.n272 B.n271 163.367
R1132 B.n272 B.n239 163.367
R1133 B.n276 B.n239 163.367
R1134 B.n277 B.n276 163.367
R1135 B.n278 B.n277 163.367
R1136 B.n278 B.n237 163.367
R1137 B.n282 B.n237 163.367
R1138 B.n283 B.n282 163.367
R1139 B.n284 B.n283 163.367
R1140 B.n284 B.n235 163.367
R1141 B.n288 B.n235 163.367
R1142 B.n289 B.n288 163.367
R1143 B.n290 B.n289 163.367
R1144 B.n290 B.n233 163.367
R1145 B.n294 B.n233 163.367
R1146 B.n295 B.n294 163.367
R1147 B.n296 B.n295 163.367
R1148 B.n296 B.n231 163.367
R1149 B.n300 B.n231 163.367
R1150 B.n301 B.n300 163.367
R1151 B.n302 B.n301 163.367
R1152 B.n302 B.n229 163.367
R1153 B.n306 B.n229 163.367
R1154 B.n307 B.n306 163.367
R1155 B.n308 B.n307 163.367
R1156 B.n308 B.n227 163.367
R1157 B.n312 B.n227 163.367
R1158 B.n313 B.n312 163.367
R1159 B.n314 B.n313 163.367
R1160 B.n314 B.n225 163.367
R1161 B.n318 B.n225 163.367
R1162 B.n319 B.n318 163.367
R1163 B.n320 B.n319 163.367
R1164 B.n320 B.n223 163.367
R1165 B.n324 B.n223 163.367
R1166 B.n325 B.n324 163.367
R1167 B.n326 B.n325 163.367
R1168 B.n326 B.n221 163.367
R1169 B.n330 B.n221 163.367
R1170 B.n433 B.t2 110.287
R1171 B.n67 B.t7 110.287
R1172 B.n191 B.t5 110.264
R1173 B.n61 B.t10 110.264
R1174 B.n191 B.n190 79.7096
R1175 B.n433 B.n432 79.7096
R1176 B.n67 B.n66 79.7096
R1177 B.n61 B.n60 79.7096
R1178 B.n419 B.n191 59.5399
R1179 B.n434 B.n433 59.5399
R1180 B.n68 B.n67 59.5399
R1181 B.n799 B.n61 59.5399
R1182 B.n889 B.n30 34.4981
R1183 B.n697 B.n98 34.4981
R1184 B.n525 B.n524 34.4981
R1185 B.n329 B.n220 34.4981
R1186 B B.n973 18.0485
R1187 B.n890 B.n889 10.6151
R1188 B.n891 B.n890 10.6151
R1189 B.n891 B.n28 10.6151
R1190 B.n895 B.n28 10.6151
R1191 B.n896 B.n895 10.6151
R1192 B.n897 B.n896 10.6151
R1193 B.n897 B.n26 10.6151
R1194 B.n901 B.n26 10.6151
R1195 B.n902 B.n901 10.6151
R1196 B.n903 B.n902 10.6151
R1197 B.n903 B.n24 10.6151
R1198 B.n907 B.n24 10.6151
R1199 B.n908 B.n907 10.6151
R1200 B.n909 B.n908 10.6151
R1201 B.n909 B.n22 10.6151
R1202 B.n913 B.n22 10.6151
R1203 B.n914 B.n913 10.6151
R1204 B.n915 B.n914 10.6151
R1205 B.n915 B.n20 10.6151
R1206 B.n919 B.n20 10.6151
R1207 B.n920 B.n919 10.6151
R1208 B.n921 B.n920 10.6151
R1209 B.n921 B.n18 10.6151
R1210 B.n925 B.n18 10.6151
R1211 B.n926 B.n925 10.6151
R1212 B.n927 B.n926 10.6151
R1213 B.n927 B.n16 10.6151
R1214 B.n931 B.n16 10.6151
R1215 B.n932 B.n931 10.6151
R1216 B.n933 B.n932 10.6151
R1217 B.n933 B.n14 10.6151
R1218 B.n937 B.n14 10.6151
R1219 B.n938 B.n937 10.6151
R1220 B.n939 B.n938 10.6151
R1221 B.n939 B.n12 10.6151
R1222 B.n943 B.n12 10.6151
R1223 B.n944 B.n943 10.6151
R1224 B.n945 B.n944 10.6151
R1225 B.n945 B.n10 10.6151
R1226 B.n949 B.n10 10.6151
R1227 B.n950 B.n949 10.6151
R1228 B.n951 B.n950 10.6151
R1229 B.n951 B.n8 10.6151
R1230 B.n955 B.n8 10.6151
R1231 B.n956 B.n955 10.6151
R1232 B.n957 B.n956 10.6151
R1233 B.n957 B.n6 10.6151
R1234 B.n961 B.n6 10.6151
R1235 B.n962 B.n961 10.6151
R1236 B.n963 B.n962 10.6151
R1237 B.n963 B.n4 10.6151
R1238 B.n967 B.n4 10.6151
R1239 B.n968 B.n967 10.6151
R1240 B.n969 B.n968 10.6151
R1241 B.n969 B.n0 10.6151
R1242 B.n885 B.n30 10.6151
R1243 B.n885 B.n884 10.6151
R1244 B.n884 B.n883 10.6151
R1245 B.n883 B.n32 10.6151
R1246 B.n879 B.n32 10.6151
R1247 B.n879 B.n878 10.6151
R1248 B.n878 B.n877 10.6151
R1249 B.n877 B.n34 10.6151
R1250 B.n873 B.n34 10.6151
R1251 B.n873 B.n872 10.6151
R1252 B.n872 B.n871 10.6151
R1253 B.n871 B.n36 10.6151
R1254 B.n867 B.n36 10.6151
R1255 B.n867 B.n866 10.6151
R1256 B.n866 B.n865 10.6151
R1257 B.n865 B.n38 10.6151
R1258 B.n861 B.n38 10.6151
R1259 B.n861 B.n860 10.6151
R1260 B.n860 B.n859 10.6151
R1261 B.n859 B.n40 10.6151
R1262 B.n855 B.n40 10.6151
R1263 B.n855 B.n854 10.6151
R1264 B.n854 B.n853 10.6151
R1265 B.n853 B.n42 10.6151
R1266 B.n849 B.n42 10.6151
R1267 B.n849 B.n848 10.6151
R1268 B.n848 B.n847 10.6151
R1269 B.n847 B.n44 10.6151
R1270 B.n843 B.n44 10.6151
R1271 B.n843 B.n842 10.6151
R1272 B.n842 B.n841 10.6151
R1273 B.n841 B.n46 10.6151
R1274 B.n837 B.n46 10.6151
R1275 B.n837 B.n836 10.6151
R1276 B.n836 B.n835 10.6151
R1277 B.n835 B.n48 10.6151
R1278 B.n831 B.n48 10.6151
R1279 B.n831 B.n830 10.6151
R1280 B.n830 B.n829 10.6151
R1281 B.n829 B.n50 10.6151
R1282 B.n825 B.n50 10.6151
R1283 B.n825 B.n824 10.6151
R1284 B.n824 B.n823 10.6151
R1285 B.n823 B.n52 10.6151
R1286 B.n819 B.n52 10.6151
R1287 B.n819 B.n818 10.6151
R1288 B.n818 B.n817 10.6151
R1289 B.n817 B.n54 10.6151
R1290 B.n813 B.n54 10.6151
R1291 B.n813 B.n812 10.6151
R1292 B.n812 B.n811 10.6151
R1293 B.n811 B.n56 10.6151
R1294 B.n807 B.n56 10.6151
R1295 B.n807 B.n806 10.6151
R1296 B.n806 B.n805 10.6151
R1297 B.n805 B.n58 10.6151
R1298 B.n801 B.n58 10.6151
R1299 B.n801 B.n800 10.6151
R1300 B.n798 B.n62 10.6151
R1301 B.n794 B.n62 10.6151
R1302 B.n794 B.n793 10.6151
R1303 B.n793 B.n792 10.6151
R1304 B.n792 B.n64 10.6151
R1305 B.n788 B.n64 10.6151
R1306 B.n788 B.n787 10.6151
R1307 B.n787 B.n786 10.6151
R1308 B.n783 B.n782 10.6151
R1309 B.n782 B.n781 10.6151
R1310 B.n781 B.n70 10.6151
R1311 B.n777 B.n70 10.6151
R1312 B.n777 B.n776 10.6151
R1313 B.n776 B.n775 10.6151
R1314 B.n775 B.n72 10.6151
R1315 B.n771 B.n72 10.6151
R1316 B.n771 B.n770 10.6151
R1317 B.n770 B.n769 10.6151
R1318 B.n769 B.n74 10.6151
R1319 B.n765 B.n74 10.6151
R1320 B.n765 B.n764 10.6151
R1321 B.n764 B.n763 10.6151
R1322 B.n763 B.n76 10.6151
R1323 B.n759 B.n76 10.6151
R1324 B.n759 B.n758 10.6151
R1325 B.n758 B.n757 10.6151
R1326 B.n757 B.n78 10.6151
R1327 B.n753 B.n78 10.6151
R1328 B.n753 B.n752 10.6151
R1329 B.n752 B.n751 10.6151
R1330 B.n751 B.n80 10.6151
R1331 B.n747 B.n80 10.6151
R1332 B.n747 B.n746 10.6151
R1333 B.n746 B.n745 10.6151
R1334 B.n745 B.n82 10.6151
R1335 B.n741 B.n82 10.6151
R1336 B.n741 B.n740 10.6151
R1337 B.n740 B.n739 10.6151
R1338 B.n739 B.n84 10.6151
R1339 B.n735 B.n84 10.6151
R1340 B.n735 B.n734 10.6151
R1341 B.n734 B.n733 10.6151
R1342 B.n733 B.n86 10.6151
R1343 B.n729 B.n86 10.6151
R1344 B.n729 B.n728 10.6151
R1345 B.n728 B.n727 10.6151
R1346 B.n727 B.n88 10.6151
R1347 B.n723 B.n88 10.6151
R1348 B.n723 B.n722 10.6151
R1349 B.n722 B.n721 10.6151
R1350 B.n721 B.n90 10.6151
R1351 B.n717 B.n90 10.6151
R1352 B.n717 B.n716 10.6151
R1353 B.n716 B.n715 10.6151
R1354 B.n715 B.n92 10.6151
R1355 B.n711 B.n92 10.6151
R1356 B.n711 B.n710 10.6151
R1357 B.n710 B.n709 10.6151
R1358 B.n709 B.n94 10.6151
R1359 B.n705 B.n94 10.6151
R1360 B.n705 B.n704 10.6151
R1361 B.n704 B.n703 10.6151
R1362 B.n703 B.n96 10.6151
R1363 B.n699 B.n96 10.6151
R1364 B.n699 B.n698 10.6151
R1365 B.n698 B.n697 10.6151
R1366 B.n693 B.n98 10.6151
R1367 B.n693 B.n692 10.6151
R1368 B.n692 B.n691 10.6151
R1369 B.n691 B.n100 10.6151
R1370 B.n687 B.n100 10.6151
R1371 B.n687 B.n686 10.6151
R1372 B.n686 B.n685 10.6151
R1373 B.n685 B.n102 10.6151
R1374 B.n681 B.n102 10.6151
R1375 B.n681 B.n680 10.6151
R1376 B.n680 B.n679 10.6151
R1377 B.n679 B.n104 10.6151
R1378 B.n675 B.n104 10.6151
R1379 B.n675 B.n674 10.6151
R1380 B.n674 B.n673 10.6151
R1381 B.n673 B.n106 10.6151
R1382 B.n669 B.n106 10.6151
R1383 B.n669 B.n668 10.6151
R1384 B.n668 B.n667 10.6151
R1385 B.n667 B.n108 10.6151
R1386 B.n663 B.n108 10.6151
R1387 B.n663 B.n662 10.6151
R1388 B.n662 B.n661 10.6151
R1389 B.n661 B.n110 10.6151
R1390 B.n657 B.n110 10.6151
R1391 B.n657 B.n656 10.6151
R1392 B.n656 B.n655 10.6151
R1393 B.n655 B.n112 10.6151
R1394 B.n651 B.n112 10.6151
R1395 B.n651 B.n650 10.6151
R1396 B.n650 B.n649 10.6151
R1397 B.n649 B.n114 10.6151
R1398 B.n645 B.n114 10.6151
R1399 B.n645 B.n644 10.6151
R1400 B.n644 B.n643 10.6151
R1401 B.n643 B.n116 10.6151
R1402 B.n639 B.n116 10.6151
R1403 B.n639 B.n638 10.6151
R1404 B.n638 B.n637 10.6151
R1405 B.n637 B.n118 10.6151
R1406 B.n633 B.n118 10.6151
R1407 B.n633 B.n632 10.6151
R1408 B.n632 B.n631 10.6151
R1409 B.n631 B.n120 10.6151
R1410 B.n627 B.n120 10.6151
R1411 B.n627 B.n626 10.6151
R1412 B.n626 B.n625 10.6151
R1413 B.n625 B.n122 10.6151
R1414 B.n621 B.n122 10.6151
R1415 B.n621 B.n620 10.6151
R1416 B.n620 B.n619 10.6151
R1417 B.n619 B.n124 10.6151
R1418 B.n615 B.n124 10.6151
R1419 B.n615 B.n614 10.6151
R1420 B.n614 B.n613 10.6151
R1421 B.n613 B.n126 10.6151
R1422 B.n609 B.n126 10.6151
R1423 B.n609 B.n608 10.6151
R1424 B.n608 B.n607 10.6151
R1425 B.n607 B.n128 10.6151
R1426 B.n603 B.n128 10.6151
R1427 B.n603 B.n602 10.6151
R1428 B.n602 B.n601 10.6151
R1429 B.n601 B.n130 10.6151
R1430 B.n597 B.n130 10.6151
R1431 B.n597 B.n596 10.6151
R1432 B.n596 B.n595 10.6151
R1433 B.n595 B.n132 10.6151
R1434 B.n591 B.n132 10.6151
R1435 B.n591 B.n590 10.6151
R1436 B.n590 B.n589 10.6151
R1437 B.n589 B.n134 10.6151
R1438 B.n585 B.n134 10.6151
R1439 B.n585 B.n584 10.6151
R1440 B.n584 B.n583 10.6151
R1441 B.n583 B.n136 10.6151
R1442 B.n579 B.n136 10.6151
R1443 B.n579 B.n578 10.6151
R1444 B.n578 B.n577 10.6151
R1445 B.n577 B.n138 10.6151
R1446 B.n573 B.n138 10.6151
R1447 B.n573 B.n572 10.6151
R1448 B.n572 B.n571 10.6151
R1449 B.n571 B.n140 10.6151
R1450 B.n567 B.n140 10.6151
R1451 B.n567 B.n566 10.6151
R1452 B.n566 B.n565 10.6151
R1453 B.n565 B.n142 10.6151
R1454 B.n561 B.n142 10.6151
R1455 B.n561 B.n560 10.6151
R1456 B.n560 B.n559 10.6151
R1457 B.n559 B.n144 10.6151
R1458 B.n555 B.n144 10.6151
R1459 B.n555 B.n554 10.6151
R1460 B.n554 B.n553 10.6151
R1461 B.n553 B.n146 10.6151
R1462 B.n549 B.n146 10.6151
R1463 B.n549 B.n548 10.6151
R1464 B.n548 B.n547 10.6151
R1465 B.n547 B.n148 10.6151
R1466 B.n543 B.n148 10.6151
R1467 B.n543 B.n542 10.6151
R1468 B.n542 B.n541 10.6151
R1469 B.n541 B.n150 10.6151
R1470 B.n537 B.n150 10.6151
R1471 B.n537 B.n536 10.6151
R1472 B.n536 B.n535 10.6151
R1473 B.n535 B.n152 10.6151
R1474 B.n531 B.n152 10.6151
R1475 B.n531 B.n530 10.6151
R1476 B.n530 B.n529 10.6151
R1477 B.n529 B.n154 10.6151
R1478 B.n525 B.n154 10.6151
R1479 B.n249 B.n1 10.6151
R1480 B.n250 B.n249 10.6151
R1481 B.n251 B.n250 10.6151
R1482 B.n251 B.n246 10.6151
R1483 B.n255 B.n246 10.6151
R1484 B.n256 B.n255 10.6151
R1485 B.n257 B.n256 10.6151
R1486 B.n257 B.n244 10.6151
R1487 B.n261 B.n244 10.6151
R1488 B.n262 B.n261 10.6151
R1489 B.n263 B.n262 10.6151
R1490 B.n263 B.n242 10.6151
R1491 B.n267 B.n242 10.6151
R1492 B.n268 B.n267 10.6151
R1493 B.n269 B.n268 10.6151
R1494 B.n269 B.n240 10.6151
R1495 B.n273 B.n240 10.6151
R1496 B.n274 B.n273 10.6151
R1497 B.n275 B.n274 10.6151
R1498 B.n275 B.n238 10.6151
R1499 B.n279 B.n238 10.6151
R1500 B.n280 B.n279 10.6151
R1501 B.n281 B.n280 10.6151
R1502 B.n281 B.n236 10.6151
R1503 B.n285 B.n236 10.6151
R1504 B.n286 B.n285 10.6151
R1505 B.n287 B.n286 10.6151
R1506 B.n287 B.n234 10.6151
R1507 B.n291 B.n234 10.6151
R1508 B.n292 B.n291 10.6151
R1509 B.n293 B.n292 10.6151
R1510 B.n293 B.n232 10.6151
R1511 B.n297 B.n232 10.6151
R1512 B.n298 B.n297 10.6151
R1513 B.n299 B.n298 10.6151
R1514 B.n299 B.n230 10.6151
R1515 B.n303 B.n230 10.6151
R1516 B.n304 B.n303 10.6151
R1517 B.n305 B.n304 10.6151
R1518 B.n305 B.n228 10.6151
R1519 B.n309 B.n228 10.6151
R1520 B.n310 B.n309 10.6151
R1521 B.n311 B.n310 10.6151
R1522 B.n311 B.n226 10.6151
R1523 B.n315 B.n226 10.6151
R1524 B.n316 B.n315 10.6151
R1525 B.n317 B.n316 10.6151
R1526 B.n317 B.n224 10.6151
R1527 B.n321 B.n224 10.6151
R1528 B.n322 B.n321 10.6151
R1529 B.n323 B.n322 10.6151
R1530 B.n323 B.n222 10.6151
R1531 B.n327 B.n222 10.6151
R1532 B.n328 B.n327 10.6151
R1533 B.n329 B.n328 10.6151
R1534 B.n333 B.n220 10.6151
R1535 B.n334 B.n333 10.6151
R1536 B.n335 B.n334 10.6151
R1537 B.n335 B.n218 10.6151
R1538 B.n339 B.n218 10.6151
R1539 B.n340 B.n339 10.6151
R1540 B.n341 B.n340 10.6151
R1541 B.n341 B.n216 10.6151
R1542 B.n345 B.n216 10.6151
R1543 B.n346 B.n345 10.6151
R1544 B.n347 B.n346 10.6151
R1545 B.n347 B.n214 10.6151
R1546 B.n351 B.n214 10.6151
R1547 B.n352 B.n351 10.6151
R1548 B.n353 B.n352 10.6151
R1549 B.n353 B.n212 10.6151
R1550 B.n357 B.n212 10.6151
R1551 B.n358 B.n357 10.6151
R1552 B.n359 B.n358 10.6151
R1553 B.n359 B.n210 10.6151
R1554 B.n363 B.n210 10.6151
R1555 B.n364 B.n363 10.6151
R1556 B.n365 B.n364 10.6151
R1557 B.n365 B.n208 10.6151
R1558 B.n369 B.n208 10.6151
R1559 B.n370 B.n369 10.6151
R1560 B.n371 B.n370 10.6151
R1561 B.n371 B.n206 10.6151
R1562 B.n375 B.n206 10.6151
R1563 B.n376 B.n375 10.6151
R1564 B.n377 B.n376 10.6151
R1565 B.n377 B.n204 10.6151
R1566 B.n381 B.n204 10.6151
R1567 B.n382 B.n381 10.6151
R1568 B.n383 B.n382 10.6151
R1569 B.n383 B.n202 10.6151
R1570 B.n387 B.n202 10.6151
R1571 B.n388 B.n387 10.6151
R1572 B.n389 B.n388 10.6151
R1573 B.n389 B.n200 10.6151
R1574 B.n393 B.n200 10.6151
R1575 B.n394 B.n393 10.6151
R1576 B.n395 B.n394 10.6151
R1577 B.n395 B.n198 10.6151
R1578 B.n399 B.n198 10.6151
R1579 B.n400 B.n399 10.6151
R1580 B.n401 B.n400 10.6151
R1581 B.n401 B.n196 10.6151
R1582 B.n405 B.n196 10.6151
R1583 B.n406 B.n405 10.6151
R1584 B.n407 B.n406 10.6151
R1585 B.n407 B.n194 10.6151
R1586 B.n411 B.n194 10.6151
R1587 B.n412 B.n411 10.6151
R1588 B.n413 B.n412 10.6151
R1589 B.n413 B.n192 10.6151
R1590 B.n417 B.n192 10.6151
R1591 B.n418 B.n417 10.6151
R1592 B.n420 B.n188 10.6151
R1593 B.n424 B.n188 10.6151
R1594 B.n425 B.n424 10.6151
R1595 B.n426 B.n425 10.6151
R1596 B.n426 B.n186 10.6151
R1597 B.n430 B.n186 10.6151
R1598 B.n431 B.n430 10.6151
R1599 B.n435 B.n431 10.6151
R1600 B.n439 B.n184 10.6151
R1601 B.n440 B.n439 10.6151
R1602 B.n441 B.n440 10.6151
R1603 B.n441 B.n182 10.6151
R1604 B.n445 B.n182 10.6151
R1605 B.n446 B.n445 10.6151
R1606 B.n447 B.n446 10.6151
R1607 B.n447 B.n180 10.6151
R1608 B.n451 B.n180 10.6151
R1609 B.n452 B.n451 10.6151
R1610 B.n453 B.n452 10.6151
R1611 B.n453 B.n178 10.6151
R1612 B.n457 B.n178 10.6151
R1613 B.n458 B.n457 10.6151
R1614 B.n459 B.n458 10.6151
R1615 B.n459 B.n176 10.6151
R1616 B.n463 B.n176 10.6151
R1617 B.n464 B.n463 10.6151
R1618 B.n465 B.n464 10.6151
R1619 B.n465 B.n174 10.6151
R1620 B.n469 B.n174 10.6151
R1621 B.n470 B.n469 10.6151
R1622 B.n471 B.n470 10.6151
R1623 B.n471 B.n172 10.6151
R1624 B.n475 B.n172 10.6151
R1625 B.n476 B.n475 10.6151
R1626 B.n477 B.n476 10.6151
R1627 B.n477 B.n170 10.6151
R1628 B.n481 B.n170 10.6151
R1629 B.n482 B.n481 10.6151
R1630 B.n483 B.n482 10.6151
R1631 B.n483 B.n168 10.6151
R1632 B.n487 B.n168 10.6151
R1633 B.n488 B.n487 10.6151
R1634 B.n489 B.n488 10.6151
R1635 B.n489 B.n166 10.6151
R1636 B.n493 B.n166 10.6151
R1637 B.n494 B.n493 10.6151
R1638 B.n495 B.n494 10.6151
R1639 B.n495 B.n164 10.6151
R1640 B.n499 B.n164 10.6151
R1641 B.n500 B.n499 10.6151
R1642 B.n501 B.n500 10.6151
R1643 B.n501 B.n162 10.6151
R1644 B.n505 B.n162 10.6151
R1645 B.n506 B.n505 10.6151
R1646 B.n507 B.n506 10.6151
R1647 B.n507 B.n160 10.6151
R1648 B.n511 B.n160 10.6151
R1649 B.n512 B.n511 10.6151
R1650 B.n513 B.n512 10.6151
R1651 B.n513 B.n158 10.6151
R1652 B.n517 B.n158 10.6151
R1653 B.n518 B.n517 10.6151
R1654 B.n519 B.n518 10.6151
R1655 B.n519 B.n156 10.6151
R1656 B.n523 B.n156 10.6151
R1657 B.n524 B.n523 10.6151
R1658 B.n973 B.n0 8.11757
R1659 B.n973 B.n1 8.11757
R1660 B.n799 B.n798 6.5566
R1661 B.n786 B.n68 6.5566
R1662 B.n420 B.n419 6.5566
R1663 B.n435 B.n434 6.5566
R1664 B.n800 B.n799 4.05904
R1665 B.n783 B.n68 4.05904
R1666 B.n419 B.n418 4.05904
R1667 B.n434 B.n184 4.05904
C0 VP w_n4258_n4546# 9.015611f
C1 VN w_n4258_n4546# 8.461821f
C2 VP VTAIL 10.628901f
C3 VN VTAIL 10.6139f
C4 w_n4258_n4546# B 12.9572f
C5 VTAIL B 5.53599f
C6 VN VP 9.16381f
C7 VDD1 w_n4258_n4546# 2.97482f
C8 VDD1 VTAIL 10.0295f
C9 VP B 2.41591f
C10 VN B 1.48536f
C11 w_n4258_n4546# VDD2 3.09762f
C12 VDD1 VP 10.8557f
C13 VTAIL VDD2 10.0883f
C14 VDD1 VN 0.152248f
C15 VDD1 B 2.87513f
C16 VP VDD2 0.557953f
C17 VN VDD2 10.4531f
C18 VDD2 B 2.97752f
C19 VDD1 VDD2 1.86719f
C20 VTAIL w_n4258_n4546# 3.8658f
C21 VDD2 VSUBS 2.37364f
C22 VDD1 VSUBS 2.97046f
C23 VTAIL VSUBS 1.625984f
C24 VN VSUBS 7.20254f
C25 VP VSUBS 4.061625f
C26 B VSUBS 6.299672f
C27 w_n4258_n4546# VSUBS 0.236728p
C28 B.n0 VSUBS 0.006338f
C29 B.n1 VSUBS 0.006338f
C30 B.n2 VSUBS 0.009373f
C31 B.n3 VSUBS 0.007183f
C32 B.n4 VSUBS 0.007183f
C33 B.n5 VSUBS 0.007183f
C34 B.n6 VSUBS 0.007183f
C35 B.n7 VSUBS 0.007183f
C36 B.n8 VSUBS 0.007183f
C37 B.n9 VSUBS 0.007183f
C38 B.n10 VSUBS 0.007183f
C39 B.n11 VSUBS 0.007183f
C40 B.n12 VSUBS 0.007183f
C41 B.n13 VSUBS 0.007183f
C42 B.n14 VSUBS 0.007183f
C43 B.n15 VSUBS 0.007183f
C44 B.n16 VSUBS 0.007183f
C45 B.n17 VSUBS 0.007183f
C46 B.n18 VSUBS 0.007183f
C47 B.n19 VSUBS 0.007183f
C48 B.n20 VSUBS 0.007183f
C49 B.n21 VSUBS 0.007183f
C50 B.n22 VSUBS 0.007183f
C51 B.n23 VSUBS 0.007183f
C52 B.n24 VSUBS 0.007183f
C53 B.n25 VSUBS 0.007183f
C54 B.n26 VSUBS 0.007183f
C55 B.n27 VSUBS 0.007183f
C56 B.n28 VSUBS 0.007183f
C57 B.n29 VSUBS 0.007183f
C58 B.n30 VSUBS 0.017635f
C59 B.n31 VSUBS 0.007183f
C60 B.n32 VSUBS 0.007183f
C61 B.n33 VSUBS 0.007183f
C62 B.n34 VSUBS 0.007183f
C63 B.n35 VSUBS 0.007183f
C64 B.n36 VSUBS 0.007183f
C65 B.n37 VSUBS 0.007183f
C66 B.n38 VSUBS 0.007183f
C67 B.n39 VSUBS 0.007183f
C68 B.n40 VSUBS 0.007183f
C69 B.n41 VSUBS 0.007183f
C70 B.n42 VSUBS 0.007183f
C71 B.n43 VSUBS 0.007183f
C72 B.n44 VSUBS 0.007183f
C73 B.n45 VSUBS 0.007183f
C74 B.n46 VSUBS 0.007183f
C75 B.n47 VSUBS 0.007183f
C76 B.n48 VSUBS 0.007183f
C77 B.n49 VSUBS 0.007183f
C78 B.n50 VSUBS 0.007183f
C79 B.n51 VSUBS 0.007183f
C80 B.n52 VSUBS 0.007183f
C81 B.n53 VSUBS 0.007183f
C82 B.n54 VSUBS 0.007183f
C83 B.n55 VSUBS 0.007183f
C84 B.n56 VSUBS 0.007183f
C85 B.n57 VSUBS 0.007183f
C86 B.n58 VSUBS 0.007183f
C87 B.n59 VSUBS 0.007183f
C88 B.t10 VSUBS 0.619481f
C89 B.t11 VSUBS 0.648327f
C90 B.t9 VSUBS 3.16204f
C91 B.n60 VSUBS 0.402855f
C92 B.n61 VSUBS 0.078993f
C93 B.n62 VSUBS 0.007183f
C94 B.n63 VSUBS 0.007183f
C95 B.n64 VSUBS 0.007183f
C96 B.n65 VSUBS 0.007183f
C97 B.t7 VSUBS 0.619459f
C98 B.t8 VSUBS 0.64831f
C99 B.t6 VSUBS 3.16204f
C100 B.n66 VSUBS 0.402871f
C101 B.n67 VSUBS 0.079015f
C102 B.n68 VSUBS 0.016642f
C103 B.n69 VSUBS 0.007183f
C104 B.n70 VSUBS 0.007183f
C105 B.n71 VSUBS 0.007183f
C106 B.n72 VSUBS 0.007183f
C107 B.n73 VSUBS 0.007183f
C108 B.n74 VSUBS 0.007183f
C109 B.n75 VSUBS 0.007183f
C110 B.n76 VSUBS 0.007183f
C111 B.n77 VSUBS 0.007183f
C112 B.n78 VSUBS 0.007183f
C113 B.n79 VSUBS 0.007183f
C114 B.n80 VSUBS 0.007183f
C115 B.n81 VSUBS 0.007183f
C116 B.n82 VSUBS 0.007183f
C117 B.n83 VSUBS 0.007183f
C118 B.n84 VSUBS 0.007183f
C119 B.n85 VSUBS 0.007183f
C120 B.n86 VSUBS 0.007183f
C121 B.n87 VSUBS 0.007183f
C122 B.n88 VSUBS 0.007183f
C123 B.n89 VSUBS 0.007183f
C124 B.n90 VSUBS 0.007183f
C125 B.n91 VSUBS 0.007183f
C126 B.n92 VSUBS 0.007183f
C127 B.n93 VSUBS 0.007183f
C128 B.n94 VSUBS 0.007183f
C129 B.n95 VSUBS 0.007183f
C130 B.n96 VSUBS 0.007183f
C131 B.n97 VSUBS 0.007183f
C132 B.n98 VSUBS 0.017223f
C133 B.n99 VSUBS 0.007183f
C134 B.n100 VSUBS 0.007183f
C135 B.n101 VSUBS 0.007183f
C136 B.n102 VSUBS 0.007183f
C137 B.n103 VSUBS 0.007183f
C138 B.n104 VSUBS 0.007183f
C139 B.n105 VSUBS 0.007183f
C140 B.n106 VSUBS 0.007183f
C141 B.n107 VSUBS 0.007183f
C142 B.n108 VSUBS 0.007183f
C143 B.n109 VSUBS 0.007183f
C144 B.n110 VSUBS 0.007183f
C145 B.n111 VSUBS 0.007183f
C146 B.n112 VSUBS 0.007183f
C147 B.n113 VSUBS 0.007183f
C148 B.n114 VSUBS 0.007183f
C149 B.n115 VSUBS 0.007183f
C150 B.n116 VSUBS 0.007183f
C151 B.n117 VSUBS 0.007183f
C152 B.n118 VSUBS 0.007183f
C153 B.n119 VSUBS 0.007183f
C154 B.n120 VSUBS 0.007183f
C155 B.n121 VSUBS 0.007183f
C156 B.n122 VSUBS 0.007183f
C157 B.n123 VSUBS 0.007183f
C158 B.n124 VSUBS 0.007183f
C159 B.n125 VSUBS 0.007183f
C160 B.n126 VSUBS 0.007183f
C161 B.n127 VSUBS 0.007183f
C162 B.n128 VSUBS 0.007183f
C163 B.n129 VSUBS 0.007183f
C164 B.n130 VSUBS 0.007183f
C165 B.n131 VSUBS 0.007183f
C166 B.n132 VSUBS 0.007183f
C167 B.n133 VSUBS 0.007183f
C168 B.n134 VSUBS 0.007183f
C169 B.n135 VSUBS 0.007183f
C170 B.n136 VSUBS 0.007183f
C171 B.n137 VSUBS 0.007183f
C172 B.n138 VSUBS 0.007183f
C173 B.n139 VSUBS 0.007183f
C174 B.n140 VSUBS 0.007183f
C175 B.n141 VSUBS 0.007183f
C176 B.n142 VSUBS 0.007183f
C177 B.n143 VSUBS 0.007183f
C178 B.n144 VSUBS 0.007183f
C179 B.n145 VSUBS 0.007183f
C180 B.n146 VSUBS 0.007183f
C181 B.n147 VSUBS 0.007183f
C182 B.n148 VSUBS 0.007183f
C183 B.n149 VSUBS 0.007183f
C184 B.n150 VSUBS 0.007183f
C185 B.n151 VSUBS 0.007183f
C186 B.n152 VSUBS 0.007183f
C187 B.n153 VSUBS 0.007183f
C188 B.n154 VSUBS 0.007183f
C189 B.n155 VSUBS 0.017635f
C190 B.n156 VSUBS 0.007183f
C191 B.n157 VSUBS 0.007183f
C192 B.n158 VSUBS 0.007183f
C193 B.n159 VSUBS 0.007183f
C194 B.n160 VSUBS 0.007183f
C195 B.n161 VSUBS 0.007183f
C196 B.n162 VSUBS 0.007183f
C197 B.n163 VSUBS 0.007183f
C198 B.n164 VSUBS 0.007183f
C199 B.n165 VSUBS 0.007183f
C200 B.n166 VSUBS 0.007183f
C201 B.n167 VSUBS 0.007183f
C202 B.n168 VSUBS 0.007183f
C203 B.n169 VSUBS 0.007183f
C204 B.n170 VSUBS 0.007183f
C205 B.n171 VSUBS 0.007183f
C206 B.n172 VSUBS 0.007183f
C207 B.n173 VSUBS 0.007183f
C208 B.n174 VSUBS 0.007183f
C209 B.n175 VSUBS 0.007183f
C210 B.n176 VSUBS 0.007183f
C211 B.n177 VSUBS 0.007183f
C212 B.n178 VSUBS 0.007183f
C213 B.n179 VSUBS 0.007183f
C214 B.n180 VSUBS 0.007183f
C215 B.n181 VSUBS 0.007183f
C216 B.n182 VSUBS 0.007183f
C217 B.n183 VSUBS 0.007183f
C218 B.n184 VSUBS 0.004965f
C219 B.n185 VSUBS 0.007183f
C220 B.n186 VSUBS 0.007183f
C221 B.n187 VSUBS 0.007183f
C222 B.n188 VSUBS 0.007183f
C223 B.n189 VSUBS 0.007183f
C224 B.t5 VSUBS 0.619481f
C225 B.t4 VSUBS 0.648327f
C226 B.t3 VSUBS 3.16204f
C227 B.n190 VSUBS 0.402855f
C228 B.n191 VSUBS 0.078993f
C229 B.n192 VSUBS 0.007183f
C230 B.n193 VSUBS 0.007183f
C231 B.n194 VSUBS 0.007183f
C232 B.n195 VSUBS 0.007183f
C233 B.n196 VSUBS 0.007183f
C234 B.n197 VSUBS 0.007183f
C235 B.n198 VSUBS 0.007183f
C236 B.n199 VSUBS 0.007183f
C237 B.n200 VSUBS 0.007183f
C238 B.n201 VSUBS 0.007183f
C239 B.n202 VSUBS 0.007183f
C240 B.n203 VSUBS 0.007183f
C241 B.n204 VSUBS 0.007183f
C242 B.n205 VSUBS 0.007183f
C243 B.n206 VSUBS 0.007183f
C244 B.n207 VSUBS 0.007183f
C245 B.n208 VSUBS 0.007183f
C246 B.n209 VSUBS 0.007183f
C247 B.n210 VSUBS 0.007183f
C248 B.n211 VSUBS 0.007183f
C249 B.n212 VSUBS 0.007183f
C250 B.n213 VSUBS 0.007183f
C251 B.n214 VSUBS 0.007183f
C252 B.n215 VSUBS 0.007183f
C253 B.n216 VSUBS 0.007183f
C254 B.n217 VSUBS 0.007183f
C255 B.n218 VSUBS 0.007183f
C256 B.n219 VSUBS 0.007183f
C257 B.n220 VSUBS 0.017635f
C258 B.n221 VSUBS 0.007183f
C259 B.n222 VSUBS 0.007183f
C260 B.n223 VSUBS 0.007183f
C261 B.n224 VSUBS 0.007183f
C262 B.n225 VSUBS 0.007183f
C263 B.n226 VSUBS 0.007183f
C264 B.n227 VSUBS 0.007183f
C265 B.n228 VSUBS 0.007183f
C266 B.n229 VSUBS 0.007183f
C267 B.n230 VSUBS 0.007183f
C268 B.n231 VSUBS 0.007183f
C269 B.n232 VSUBS 0.007183f
C270 B.n233 VSUBS 0.007183f
C271 B.n234 VSUBS 0.007183f
C272 B.n235 VSUBS 0.007183f
C273 B.n236 VSUBS 0.007183f
C274 B.n237 VSUBS 0.007183f
C275 B.n238 VSUBS 0.007183f
C276 B.n239 VSUBS 0.007183f
C277 B.n240 VSUBS 0.007183f
C278 B.n241 VSUBS 0.007183f
C279 B.n242 VSUBS 0.007183f
C280 B.n243 VSUBS 0.007183f
C281 B.n244 VSUBS 0.007183f
C282 B.n245 VSUBS 0.007183f
C283 B.n246 VSUBS 0.007183f
C284 B.n247 VSUBS 0.007183f
C285 B.n248 VSUBS 0.007183f
C286 B.n249 VSUBS 0.007183f
C287 B.n250 VSUBS 0.007183f
C288 B.n251 VSUBS 0.007183f
C289 B.n252 VSUBS 0.007183f
C290 B.n253 VSUBS 0.007183f
C291 B.n254 VSUBS 0.007183f
C292 B.n255 VSUBS 0.007183f
C293 B.n256 VSUBS 0.007183f
C294 B.n257 VSUBS 0.007183f
C295 B.n258 VSUBS 0.007183f
C296 B.n259 VSUBS 0.007183f
C297 B.n260 VSUBS 0.007183f
C298 B.n261 VSUBS 0.007183f
C299 B.n262 VSUBS 0.007183f
C300 B.n263 VSUBS 0.007183f
C301 B.n264 VSUBS 0.007183f
C302 B.n265 VSUBS 0.007183f
C303 B.n266 VSUBS 0.007183f
C304 B.n267 VSUBS 0.007183f
C305 B.n268 VSUBS 0.007183f
C306 B.n269 VSUBS 0.007183f
C307 B.n270 VSUBS 0.007183f
C308 B.n271 VSUBS 0.007183f
C309 B.n272 VSUBS 0.007183f
C310 B.n273 VSUBS 0.007183f
C311 B.n274 VSUBS 0.007183f
C312 B.n275 VSUBS 0.007183f
C313 B.n276 VSUBS 0.007183f
C314 B.n277 VSUBS 0.007183f
C315 B.n278 VSUBS 0.007183f
C316 B.n279 VSUBS 0.007183f
C317 B.n280 VSUBS 0.007183f
C318 B.n281 VSUBS 0.007183f
C319 B.n282 VSUBS 0.007183f
C320 B.n283 VSUBS 0.007183f
C321 B.n284 VSUBS 0.007183f
C322 B.n285 VSUBS 0.007183f
C323 B.n286 VSUBS 0.007183f
C324 B.n287 VSUBS 0.007183f
C325 B.n288 VSUBS 0.007183f
C326 B.n289 VSUBS 0.007183f
C327 B.n290 VSUBS 0.007183f
C328 B.n291 VSUBS 0.007183f
C329 B.n292 VSUBS 0.007183f
C330 B.n293 VSUBS 0.007183f
C331 B.n294 VSUBS 0.007183f
C332 B.n295 VSUBS 0.007183f
C333 B.n296 VSUBS 0.007183f
C334 B.n297 VSUBS 0.007183f
C335 B.n298 VSUBS 0.007183f
C336 B.n299 VSUBS 0.007183f
C337 B.n300 VSUBS 0.007183f
C338 B.n301 VSUBS 0.007183f
C339 B.n302 VSUBS 0.007183f
C340 B.n303 VSUBS 0.007183f
C341 B.n304 VSUBS 0.007183f
C342 B.n305 VSUBS 0.007183f
C343 B.n306 VSUBS 0.007183f
C344 B.n307 VSUBS 0.007183f
C345 B.n308 VSUBS 0.007183f
C346 B.n309 VSUBS 0.007183f
C347 B.n310 VSUBS 0.007183f
C348 B.n311 VSUBS 0.007183f
C349 B.n312 VSUBS 0.007183f
C350 B.n313 VSUBS 0.007183f
C351 B.n314 VSUBS 0.007183f
C352 B.n315 VSUBS 0.007183f
C353 B.n316 VSUBS 0.007183f
C354 B.n317 VSUBS 0.007183f
C355 B.n318 VSUBS 0.007183f
C356 B.n319 VSUBS 0.007183f
C357 B.n320 VSUBS 0.007183f
C358 B.n321 VSUBS 0.007183f
C359 B.n322 VSUBS 0.007183f
C360 B.n323 VSUBS 0.007183f
C361 B.n324 VSUBS 0.007183f
C362 B.n325 VSUBS 0.007183f
C363 B.n326 VSUBS 0.007183f
C364 B.n327 VSUBS 0.007183f
C365 B.n328 VSUBS 0.007183f
C366 B.n329 VSUBS 0.017223f
C367 B.n330 VSUBS 0.017223f
C368 B.n331 VSUBS 0.017635f
C369 B.n332 VSUBS 0.007183f
C370 B.n333 VSUBS 0.007183f
C371 B.n334 VSUBS 0.007183f
C372 B.n335 VSUBS 0.007183f
C373 B.n336 VSUBS 0.007183f
C374 B.n337 VSUBS 0.007183f
C375 B.n338 VSUBS 0.007183f
C376 B.n339 VSUBS 0.007183f
C377 B.n340 VSUBS 0.007183f
C378 B.n341 VSUBS 0.007183f
C379 B.n342 VSUBS 0.007183f
C380 B.n343 VSUBS 0.007183f
C381 B.n344 VSUBS 0.007183f
C382 B.n345 VSUBS 0.007183f
C383 B.n346 VSUBS 0.007183f
C384 B.n347 VSUBS 0.007183f
C385 B.n348 VSUBS 0.007183f
C386 B.n349 VSUBS 0.007183f
C387 B.n350 VSUBS 0.007183f
C388 B.n351 VSUBS 0.007183f
C389 B.n352 VSUBS 0.007183f
C390 B.n353 VSUBS 0.007183f
C391 B.n354 VSUBS 0.007183f
C392 B.n355 VSUBS 0.007183f
C393 B.n356 VSUBS 0.007183f
C394 B.n357 VSUBS 0.007183f
C395 B.n358 VSUBS 0.007183f
C396 B.n359 VSUBS 0.007183f
C397 B.n360 VSUBS 0.007183f
C398 B.n361 VSUBS 0.007183f
C399 B.n362 VSUBS 0.007183f
C400 B.n363 VSUBS 0.007183f
C401 B.n364 VSUBS 0.007183f
C402 B.n365 VSUBS 0.007183f
C403 B.n366 VSUBS 0.007183f
C404 B.n367 VSUBS 0.007183f
C405 B.n368 VSUBS 0.007183f
C406 B.n369 VSUBS 0.007183f
C407 B.n370 VSUBS 0.007183f
C408 B.n371 VSUBS 0.007183f
C409 B.n372 VSUBS 0.007183f
C410 B.n373 VSUBS 0.007183f
C411 B.n374 VSUBS 0.007183f
C412 B.n375 VSUBS 0.007183f
C413 B.n376 VSUBS 0.007183f
C414 B.n377 VSUBS 0.007183f
C415 B.n378 VSUBS 0.007183f
C416 B.n379 VSUBS 0.007183f
C417 B.n380 VSUBS 0.007183f
C418 B.n381 VSUBS 0.007183f
C419 B.n382 VSUBS 0.007183f
C420 B.n383 VSUBS 0.007183f
C421 B.n384 VSUBS 0.007183f
C422 B.n385 VSUBS 0.007183f
C423 B.n386 VSUBS 0.007183f
C424 B.n387 VSUBS 0.007183f
C425 B.n388 VSUBS 0.007183f
C426 B.n389 VSUBS 0.007183f
C427 B.n390 VSUBS 0.007183f
C428 B.n391 VSUBS 0.007183f
C429 B.n392 VSUBS 0.007183f
C430 B.n393 VSUBS 0.007183f
C431 B.n394 VSUBS 0.007183f
C432 B.n395 VSUBS 0.007183f
C433 B.n396 VSUBS 0.007183f
C434 B.n397 VSUBS 0.007183f
C435 B.n398 VSUBS 0.007183f
C436 B.n399 VSUBS 0.007183f
C437 B.n400 VSUBS 0.007183f
C438 B.n401 VSUBS 0.007183f
C439 B.n402 VSUBS 0.007183f
C440 B.n403 VSUBS 0.007183f
C441 B.n404 VSUBS 0.007183f
C442 B.n405 VSUBS 0.007183f
C443 B.n406 VSUBS 0.007183f
C444 B.n407 VSUBS 0.007183f
C445 B.n408 VSUBS 0.007183f
C446 B.n409 VSUBS 0.007183f
C447 B.n410 VSUBS 0.007183f
C448 B.n411 VSUBS 0.007183f
C449 B.n412 VSUBS 0.007183f
C450 B.n413 VSUBS 0.007183f
C451 B.n414 VSUBS 0.007183f
C452 B.n415 VSUBS 0.007183f
C453 B.n416 VSUBS 0.007183f
C454 B.n417 VSUBS 0.007183f
C455 B.n418 VSUBS 0.004965f
C456 B.n419 VSUBS 0.016642f
C457 B.n420 VSUBS 0.00581f
C458 B.n421 VSUBS 0.007183f
C459 B.n422 VSUBS 0.007183f
C460 B.n423 VSUBS 0.007183f
C461 B.n424 VSUBS 0.007183f
C462 B.n425 VSUBS 0.007183f
C463 B.n426 VSUBS 0.007183f
C464 B.n427 VSUBS 0.007183f
C465 B.n428 VSUBS 0.007183f
C466 B.n429 VSUBS 0.007183f
C467 B.n430 VSUBS 0.007183f
C468 B.n431 VSUBS 0.007183f
C469 B.t2 VSUBS 0.619459f
C470 B.t1 VSUBS 0.64831f
C471 B.t0 VSUBS 3.16204f
C472 B.n432 VSUBS 0.402871f
C473 B.n433 VSUBS 0.079015f
C474 B.n434 VSUBS 0.016642f
C475 B.n435 VSUBS 0.00581f
C476 B.n436 VSUBS 0.007183f
C477 B.n437 VSUBS 0.007183f
C478 B.n438 VSUBS 0.007183f
C479 B.n439 VSUBS 0.007183f
C480 B.n440 VSUBS 0.007183f
C481 B.n441 VSUBS 0.007183f
C482 B.n442 VSUBS 0.007183f
C483 B.n443 VSUBS 0.007183f
C484 B.n444 VSUBS 0.007183f
C485 B.n445 VSUBS 0.007183f
C486 B.n446 VSUBS 0.007183f
C487 B.n447 VSUBS 0.007183f
C488 B.n448 VSUBS 0.007183f
C489 B.n449 VSUBS 0.007183f
C490 B.n450 VSUBS 0.007183f
C491 B.n451 VSUBS 0.007183f
C492 B.n452 VSUBS 0.007183f
C493 B.n453 VSUBS 0.007183f
C494 B.n454 VSUBS 0.007183f
C495 B.n455 VSUBS 0.007183f
C496 B.n456 VSUBS 0.007183f
C497 B.n457 VSUBS 0.007183f
C498 B.n458 VSUBS 0.007183f
C499 B.n459 VSUBS 0.007183f
C500 B.n460 VSUBS 0.007183f
C501 B.n461 VSUBS 0.007183f
C502 B.n462 VSUBS 0.007183f
C503 B.n463 VSUBS 0.007183f
C504 B.n464 VSUBS 0.007183f
C505 B.n465 VSUBS 0.007183f
C506 B.n466 VSUBS 0.007183f
C507 B.n467 VSUBS 0.007183f
C508 B.n468 VSUBS 0.007183f
C509 B.n469 VSUBS 0.007183f
C510 B.n470 VSUBS 0.007183f
C511 B.n471 VSUBS 0.007183f
C512 B.n472 VSUBS 0.007183f
C513 B.n473 VSUBS 0.007183f
C514 B.n474 VSUBS 0.007183f
C515 B.n475 VSUBS 0.007183f
C516 B.n476 VSUBS 0.007183f
C517 B.n477 VSUBS 0.007183f
C518 B.n478 VSUBS 0.007183f
C519 B.n479 VSUBS 0.007183f
C520 B.n480 VSUBS 0.007183f
C521 B.n481 VSUBS 0.007183f
C522 B.n482 VSUBS 0.007183f
C523 B.n483 VSUBS 0.007183f
C524 B.n484 VSUBS 0.007183f
C525 B.n485 VSUBS 0.007183f
C526 B.n486 VSUBS 0.007183f
C527 B.n487 VSUBS 0.007183f
C528 B.n488 VSUBS 0.007183f
C529 B.n489 VSUBS 0.007183f
C530 B.n490 VSUBS 0.007183f
C531 B.n491 VSUBS 0.007183f
C532 B.n492 VSUBS 0.007183f
C533 B.n493 VSUBS 0.007183f
C534 B.n494 VSUBS 0.007183f
C535 B.n495 VSUBS 0.007183f
C536 B.n496 VSUBS 0.007183f
C537 B.n497 VSUBS 0.007183f
C538 B.n498 VSUBS 0.007183f
C539 B.n499 VSUBS 0.007183f
C540 B.n500 VSUBS 0.007183f
C541 B.n501 VSUBS 0.007183f
C542 B.n502 VSUBS 0.007183f
C543 B.n503 VSUBS 0.007183f
C544 B.n504 VSUBS 0.007183f
C545 B.n505 VSUBS 0.007183f
C546 B.n506 VSUBS 0.007183f
C547 B.n507 VSUBS 0.007183f
C548 B.n508 VSUBS 0.007183f
C549 B.n509 VSUBS 0.007183f
C550 B.n510 VSUBS 0.007183f
C551 B.n511 VSUBS 0.007183f
C552 B.n512 VSUBS 0.007183f
C553 B.n513 VSUBS 0.007183f
C554 B.n514 VSUBS 0.007183f
C555 B.n515 VSUBS 0.007183f
C556 B.n516 VSUBS 0.007183f
C557 B.n517 VSUBS 0.007183f
C558 B.n518 VSUBS 0.007183f
C559 B.n519 VSUBS 0.007183f
C560 B.n520 VSUBS 0.007183f
C561 B.n521 VSUBS 0.007183f
C562 B.n522 VSUBS 0.007183f
C563 B.n523 VSUBS 0.007183f
C564 B.n524 VSUBS 0.016831f
C565 B.n525 VSUBS 0.018027f
C566 B.n526 VSUBS 0.017223f
C567 B.n527 VSUBS 0.007183f
C568 B.n528 VSUBS 0.007183f
C569 B.n529 VSUBS 0.007183f
C570 B.n530 VSUBS 0.007183f
C571 B.n531 VSUBS 0.007183f
C572 B.n532 VSUBS 0.007183f
C573 B.n533 VSUBS 0.007183f
C574 B.n534 VSUBS 0.007183f
C575 B.n535 VSUBS 0.007183f
C576 B.n536 VSUBS 0.007183f
C577 B.n537 VSUBS 0.007183f
C578 B.n538 VSUBS 0.007183f
C579 B.n539 VSUBS 0.007183f
C580 B.n540 VSUBS 0.007183f
C581 B.n541 VSUBS 0.007183f
C582 B.n542 VSUBS 0.007183f
C583 B.n543 VSUBS 0.007183f
C584 B.n544 VSUBS 0.007183f
C585 B.n545 VSUBS 0.007183f
C586 B.n546 VSUBS 0.007183f
C587 B.n547 VSUBS 0.007183f
C588 B.n548 VSUBS 0.007183f
C589 B.n549 VSUBS 0.007183f
C590 B.n550 VSUBS 0.007183f
C591 B.n551 VSUBS 0.007183f
C592 B.n552 VSUBS 0.007183f
C593 B.n553 VSUBS 0.007183f
C594 B.n554 VSUBS 0.007183f
C595 B.n555 VSUBS 0.007183f
C596 B.n556 VSUBS 0.007183f
C597 B.n557 VSUBS 0.007183f
C598 B.n558 VSUBS 0.007183f
C599 B.n559 VSUBS 0.007183f
C600 B.n560 VSUBS 0.007183f
C601 B.n561 VSUBS 0.007183f
C602 B.n562 VSUBS 0.007183f
C603 B.n563 VSUBS 0.007183f
C604 B.n564 VSUBS 0.007183f
C605 B.n565 VSUBS 0.007183f
C606 B.n566 VSUBS 0.007183f
C607 B.n567 VSUBS 0.007183f
C608 B.n568 VSUBS 0.007183f
C609 B.n569 VSUBS 0.007183f
C610 B.n570 VSUBS 0.007183f
C611 B.n571 VSUBS 0.007183f
C612 B.n572 VSUBS 0.007183f
C613 B.n573 VSUBS 0.007183f
C614 B.n574 VSUBS 0.007183f
C615 B.n575 VSUBS 0.007183f
C616 B.n576 VSUBS 0.007183f
C617 B.n577 VSUBS 0.007183f
C618 B.n578 VSUBS 0.007183f
C619 B.n579 VSUBS 0.007183f
C620 B.n580 VSUBS 0.007183f
C621 B.n581 VSUBS 0.007183f
C622 B.n582 VSUBS 0.007183f
C623 B.n583 VSUBS 0.007183f
C624 B.n584 VSUBS 0.007183f
C625 B.n585 VSUBS 0.007183f
C626 B.n586 VSUBS 0.007183f
C627 B.n587 VSUBS 0.007183f
C628 B.n588 VSUBS 0.007183f
C629 B.n589 VSUBS 0.007183f
C630 B.n590 VSUBS 0.007183f
C631 B.n591 VSUBS 0.007183f
C632 B.n592 VSUBS 0.007183f
C633 B.n593 VSUBS 0.007183f
C634 B.n594 VSUBS 0.007183f
C635 B.n595 VSUBS 0.007183f
C636 B.n596 VSUBS 0.007183f
C637 B.n597 VSUBS 0.007183f
C638 B.n598 VSUBS 0.007183f
C639 B.n599 VSUBS 0.007183f
C640 B.n600 VSUBS 0.007183f
C641 B.n601 VSUBS 0.007183f
C642 B.n602 VSUBS 0.007183f
C643 B.n603 VSUBS 0.007183f
C644 B.n604 VSUBS 0.007183f
C645 B.n605 VSUBS 0.007183f
C646 B.n606 VSUBS 0.007183f
C647 B.n607 VSUBS 0.007183f
C648 B.n608 VSUBS 0.007183f
C649 B.n609 VSUBS 0.007183f
C650 B.n610 VSUBS 0.007183f
C651 B.n611 VSUBS 0.007183f
C652 B.n612 VSUBS 0.007183f
C653 B.n613 VSUBS 0.007183f
C654 B.n614 VSUBS 0.007183f
C655 B.n615 VSUBS 0.007183f
C656 B.n616 VSUBS 0.007183f
C657 B.n617 VSUBS 0.007183f
C658 B.n618 VSUBS 0.007183f
C659 B.n619 VSUBS 0.007183f
C660 B.n620 VSUBS 0.007183f
C661 B.n621 VSUBS 0.007183f
C662 B.n622 VSUBS 0.007183f
C663 B.n623 VSUBS 0.007183f
C664 B.n624 VSUBS 0.007183f
C665 B.n625 VSUBS 0.007183f
C666 B.n626 VSUBS 0.007183f
C667 B.n627 VSUBS 0.007183f
C668 B.n628 VSUBS 0.007183f
C669 B.n629 VSUBS 0.007183f
C670 B.n630 VSUBS 0.007183f
C671 B.n631 VSUBS 0.007183f
C672 B.n632 VSUBS 0.007183f
C673 B.n633 VSUBS 0.007183f
C674 B.n634 VSUBS 0.007183f
C675 B.n635 VSUBS 0.007183f
C676 B.n636 VSUBS 0.007183f
C677 B.n637 VSUBS 0.007183f
C678 B.n638 VSUBS 0.007183f
C679 B.n639 VSUBS 0.007183f
C680 B.n640 VSUBS 0.007183f
C681 B.n641 VSUBS 0.007183f
C682 B.n642 VSUBS 0.007183f
C683 B.n643 VSUBS 0.007183f
C684 B.n644 VSUBS 0.007183f
C685 B.n645 VSUBS 0.007183f
C686 B.n646 VSUBS 0.007183f
C687 B.n647 VSUBS 0.007183f
C688 B.n648 VSUBS 0.007183f
C689 B.n649 VSUBS 0.007183f
C690 B.n650 VSUBS 0.007183f
C691 B.n651 VSUBS 0.007183f
C692 B.n652 VSUBS 0.007183f
C693 B.n653 VSUBS 0.007183f
C694 B.n654 VSUBS 0.007183f
C695 B.n655 VSUBS 0.007183f
C696 B.n656 VSUBS 0.007183f
C697 B.n657 VSUBS 0.007183f
C698 B.n658 VSUBS 0.007183f
C699 B.n659 VSUBS 0.007183f
C700 B.n660 VSUBS 0.007183f
C701 B.n661 VSUBS 0.007183f
C702 B.n662 VSUBS 0.007183f
C703 B.n663 VSUBS 0.007183f
C704 B.n664 VSUBS 0.007183f
C705 B.n665 VSUBS 0.007183f
C706 B.n666 VSUBS 0.007183f
C707 B.n667 VSUBS 0.007183f
C708 B.n668 VSUBS 0.007183f
C709 B.n669 VSUBS 0.007183f
C710 B.n670 VSUBS 0.007183f
C711 B.n671 VSUBS 0.007183f
C712 B.n672 VSUBS 0.007183f
C713 B.n673 VSUBS 0.007183f
C714 B.n674 VSUBS 0.007183f
C715 B.n675 VSUBS 0.007183f
C716 B.n676 VSUBS 0.007183f
C717 B.n677 VSUBS 0.007183f
C718 B.n678 VSUBS 0.007183f
C719 B.n679 VSUBS 0.007183f
C720 B.n680 VSUBS 0.007183f
C721 B.n681 VSUBS 0.007183f
C722 B.n682 VSUBS 0.007183f
C723 B.n683 VSUBS 0.007183f
C724 B.n684 VSUBS 0.007183f
C725 B.n685 VSUBS 0.007183f
C726 B.n686 VSUBS 0.007183f
C727 B.n687 VSUBS 0.007183f
C728 B.n688 VSUBS 0.007183f
C729 B.n689 VSUBS 0.007183f
C730 B.n690 VSUBS 0.007183f
C731 B.n691 VSUBS 0.007183f
C732 B.n692 VSUBS 0.007183f
C733 B.n693 VSUBS 0.007183f
C734 B.n694 VSUBS 0.007183f
C735 B.n695 VSUBS 0.017223f
C736 B.n696 VSUBS 0.017635f
C737 B.n697 VSUBS 0.017635f
C738 B.n698 VSUBS 0.007183f
C739 B.n699 VSUBS 0.007183f
C740 B.n700 VSUBS 0.007183f
C741 B.n701 VSUBS 0.007183f
C742 B.n702 VSUBS 0.007183f
C743 B.n703 VSUBS 0.007183f
C744 B.n704 VSUBS 0.007183f
C745 B.n705 VSUBS 0.007183f
C746 B.n706 VSUBS 0.007183f
C747 B.n707 VSUBS 0.007183f
C748 B.n708 VSUBS 0.007183f
C749 B.n709 VSUBS 0.007183f
C750 B.n710 VSUBS 0.007183f
C751 B.n711 VSUBS 0.007183f
C752 B.n712 VSUBS 0.007183f
C753 B.n713 VSUBS 0.007183f
C754 B.n714 VSUBS 0.007183f
C755 B.n715 VSUBS 0.007183f
C756 B.n716 VSUBS 0.007183f
C757 B.n717 VSUBS 0.007183f
C758 B.n718 VSUBS 0.007183f
C759 B.n719 VSUBS 0.007183f
C760 B.n720 VSUBS 0.007183f
C761 B.n721 VSUBS 0.007183f
C762 B.n722 VSUBS 0.007183f
C763 B.n723 VSUBS 0.007183f
C764 B.n724 VSUBS 0.007183f
C765 B.n725 VSUBS 0.007183f
C766 B.n726 VSUBS 0.007183f
C767 B.n727 VSUBS 0.007183f
C768 B.n728 VSUBS 0.007183f
C769 B.n729 VSUBS 0.007183f
C770 B.n730 VSUBS 0.007183f
C771 B.n731 VSUBS 0.007183f
C772 B.n732 VSUBS 0.007183f
C773 B.n733 VSUBS 0.007183f
C774 B.n734 VSUBS 0.007183f
C775 B.n735 VSUBS 0.007183f
C776 B.n736 VSUBS 0.007183f
C777 B.n737 VSUBS 0.007183f
C778 B.n738 VSUBS 0.007183f
C779 B.n739 VSUBS 0.007183f
C780 B.n740 VSUBS 0.007183f
C781 B.n741 VSUBS 0.007183f
C782 B.n742 VSUBS 0.007183f
C783 B.n743 VSUBS 0.007183f
C784 B.n744 VSUBS 0.007183f
C785 B.n745 VSUBS 0.007183f
C786 B.n746 VSUBS 0.007183f
C787 B.n747 VSUBS 0.007183f
C788 B.n748 VSUBS 0.007183f
C789 B.n749 VSUBS 0.007183f
C790 B.n750 VSUBS 0.007183f
C791 B.n751 VSUBS 0.007183f
C792 B.n752 VSUBS 0.007183f
C793 B.n753 VSUBS 0.007183f
C794 B.n754 VSUBS 0.007183f
C795 B.n755 VSUBS 0.007183f
C796 B.n756 VSUBS 0.007183f
C797 B.n757 VSUBS 0.007183f
C798 B.n758 VSUBS 0.007183f
C799 B.n759 VSUBS 0.007183f
C800 B.n760 VSUBS 0.007183f
C801 B.n761 VSUBS 0.007183f
C802 B.n762 VSUBS 0.007183f
C803 B.n763 VSUBS 0.007183f
C804 B.n764 VSUBS 0.007183f
C805 B.n765 VSUBS 0.007183f
C806 B.n766 VSUBS 0.007183f
C807 B.n767 VSUBS 0.007183f
C808 B.n768 VSUBS 0.007183f
C809 B.n769 VSUBS 0.007183f
C810 B.n770 VSUBS 0.007183f
C811 B.n771 VSUBS 0.007183f
C812 B.n772 VSUBS 0.007183f
C813 B.n773 VSUBS 0.007183f
C814 B.n774 VSUBS 0.007183f
C815 B.n775 VSUBS 0.007183f
C816 B.n776 VSUBS 0.007183f
C817 B.n777 VSUBS 0.007183f
C818 B.n778 VSUBS 0.007183f
C819 B.n779 VSUBS 0.007183f
C820 B.n780 VSUBS 0.007183f
C821 B.n781 VSUBS 0.007183f
C822 B.n782 VSUBS 0.007183f
C823 B.n783 VSUBS 0.004965f
C824 B.n784 VSUBS 0.007183f
C825 B.n785 VSUBS 0.007183f
C826 B.n786 VSUBS 0.00581f
C827 B.n787 VSUBS 0.007183f
C828 B.n788 VSUBS 0.007183f
C829 B.n789 VSUBS 0.007183f
C830 B.n790 VSUBS 0.007183f
C831 B.n791 VSUBS 0.007183f
C832 B.n792 VSUBS 0.007183f
C833 B.n793 VSUBS 0.007183f
C834 B.n794 VSUBS 0.007183f
C835 B.n795 VSUBS 0.007183f
C836 B.n796 VSUBS 0.007183f
C837 B.n797 VSUBS 0.007183f
C838 B.n798 VSUBS 0.00581f
C839 B.n799 VSUBS 0.016642f
C840 B.n800 VSUBS 0.004965f
C841 B.n801 VSUBS 0.007183f
C842 B.n802 VSUBS 0.007183f
C843 B.n803 VSUBS 0.007183f
C844 B.n804 VSUBS 0.007183f
C845 B.n805 VSUBS 0.007183f
C846 B.n806 VSUBS 0.007183f
C847 B.n807 VSUBS 0.007183f
C848 B.n808 VSUBS 0.007183f
C849 B.n809 VSUBS 0.007183f
C850 B.n810 VSUBS 0.007183f
C851 B.n811 VSUBS 0.007183f
C852 B.n812 VSUBS 0.007183f
C853 B.n813 VSUBS 0.007183f
C854 B.n814 VSUBS 0.007183f
C855 B.n815 VSUBS 0.007183f
C856 B.n816 VSUBS 0.007183f
C857 B.n817 VSUBS 0.007183f
C858 B.n818 VSUBS 0.007183f
C859 B.n819 VSUBS 0.007183f
C860 B.n820 VSUBS 0.007183f
C861 B.n821 VSUBS 0.007183f
C862 B.n822 VSUBS 0.007183f
C863 B.n823 VSUBS 0.007183f
C864 B.n824 VSUBS 0.007183f
C865 B.n825 VSUBS 0.007183f
C866 B.n826 VSUBS 0.007183f
C867 B.n827 VSUBS 0.007183f
C868 B.n828 VSUBS 0.007183f
C869 B.n829 VSUBS 0.007183f
C870 B.n830 VSUBS 0.007183f
C871 B.n831 VSUBS 0.007183f
C872 B.n832 VSUBS 0.007183f
C873 B.n833 VSUBS 0.007183f
C874 B.n834 VSUBS 0.007183f
C875 B.n835 VSUBS 0.007183f
C876 B.n836 VSUBS 0.007183f
C877 B.n837 VSUBS 0.007183f
C878 B.n838 VSUBS 0.007183f
C879 B.n839 VSUBS 0.007183f
C880 B.n840 VSUBS 0.007183f
C881 B.n841 VSUBS 0.007183f
C882 B.n842 VSUBS 0.007183f
C883 B.n843 VSUBS 0.007183f
C884 B.n844 VSUBS 0.007183f
C885 B.n845 VSUBS 0.007183f
C886 B.n846 VSUBS 0.007183f
C887 B.n847 VSUBS 0.007183f
C888 B.n848 VSUBS 0.007183f
C889 B.n849 VSUBS 0.007183f
C890 B.n850 VSUBS 0.007183f
C891 B.n851 VSUBS 0.007183f
C892 B.n852 VSUBS 0.007183f
C893 B.n853 VSUBS 0.007183f
C894 B.n854 VSUBS 0.007183f
C895 B.n855 VSUBS 0.007183f
C896 B.n856 VSUBS 0.007183f
C897 B.n857 VSUBS 0.007183f
C898 B.n858 VSUBS 0.007183f
C899 B.n859 VSUBS 0.007183f
C900 B.n860 VSUBS 0.007183f
C901 B.n861 VSUBS 0.007183f
C902 B.n862 VSUBS 0.007183f
C903 B.n863 VSUBS 0.007183f
C904 B.n864 VSUBS 0.007183f
C905 B.n865 VSUBS 0.007183f
C906 B.n866 VSUBS 0.007183f
C907 B.n867 VSUBS 0.007183f
C908 B.n868 VSUBS 0.007183f
C909 B.n869 VSUBS 0.007183f
C910 B.n870 VSUBS 0.007183f
C911 B.n871 VSUBS 0.007183f
C912 B.n872 VSUBS 0.007183f
C913 B.n873 VSUBS 0.007183f
C914 B.n874 VSUBS 0.007183f
C915 B.n875 VSUBS 0.007183f
C916 B.n876 VSUBS 0.007183f
C917 B.n877 VSUBS 0.007183f
C918 B.n878 VSUBS 0.007183f
C919 B.n879 VSUBS 0.007183f
C920 B.n880 VSUBS 0.007183f
C921 B.n881 VSUBS 0.007183f
C922 B.n882 VSUBS 0.007183f
C923 B.n883 VSUBS 0.007183f
C924 B.n884 VSUBS 0.007183f
C925 B.n885 VSUBS 0.007183f
C926 B.n886 VSUBS 0.007183f
C927 B.n887 VSUBS 0.017635f
C928 B.n888 VSUBS 0.017223f
C929 B.n889 VSUBS 0.017223f
C930 B.n890 VSUBS 0.007183f
C931 B.n891 VSUBS 0.007183f
C932 B.n892 VSUBS 0.007183f
C933 B.n893 VSUBS 0.007183f
C934 B.n894 VSUBS 0.007183f
C935 B.n895 VSUBS 0.007183f
C936 B.n896 VSUBS 0.007183f
C937 B.n897 VSUBS 0.007183f
C938 B.n898 VSUBS 0.007183f
C939 B.n899 VSUBS 0.007183f
C940 B.n900 VSUBS 0.007183f
C941 B.n901 VSUBS 0.007183f
C942 B.n902 VSUBS 0.007183f
C943 B.n903 VSUBS 0.007183f
C944 B.n904 VSUBS 0.007183f
C945 B.n905 VSUBS 0.007183f
C946 B.n906 VSUBS 0.007183f
C947 B.n907 VSUBS 0.007183f
C948 B.n908 VSUBS 0.007183f
C949 B.n909 VSUBS 0.007183f
C950 B.n910 VSUBS 0.007183f
C951 B.n911 VSUBS 0.007183f
C952 B.n912 VSUBS 0.007183f
C953 B.n913 VSUBS 0.007183f
C954 B.n914 VSUBS 0.007183f
C955 B.n915 VSUBS 0.007183f
C956 B.n916 VSUBS 0.007183f
C957 B.n917 VSUBS 0.007183f
C958 B.n918 VSUBS 0.007183f
C959 B.n919 VSUBS 0.007183f
C960 B.n920 VSUBS 0.007183f
C961 B.n921 VSUBS 0.007183f
C962 B.n922 VSUBS 0.007183f
C963 B.n923 VSUBS 0.007183f
C964 B.n924 VSUBS 0.007183f
C965 B.n925 VSUBS 0.007183f
C966 B.n926 VSUBS 0.007183f
C967 B.n927 VSUBS 0.007183f
C968 B.n928 VSUBS 0.007183f
C969 B.n929 VSUBS 0.007183f
C970 B.n930 VSUBS 0.007183f
C971 B.n931 VSUBS 0.007183f
C972 B.n932 VSUBS 0.007183f
C973 B.n933 VSUBS 0.007183f
C974 B.n934 VSUBS 0.007183f
C975 B.n935 VSUBS 0.007183f
C976 B.n936 VSUBS 0.007183f
C977 B.n937 VSUBS 0.007183f
C978 B.n938 VSUBS 0.007183f
C979 B.n939 VSUBS 0.007183f
C980 B.n940 VSUBS 0.007183f
C981 B.n941 VSUBS 0.007183f
C982 B.n942 VSUBS 0.007183f
C983 B.n943 VSUBS 0.007183f
C984 B.n944 VSUBS 0.007183f
C985 B.n945 VSUBS 0.007183f
C986 B.n946 VSUBS 0.007183f
C987 B.n947 VSUBS 0.007183f
C988 B.n948 VSUBS 0.007183f
C989 B.n949 VSUBS 0.007183f
C990 B.n950 VSUBS 0.007183f
C991 B.n951 VSUBS 0.007183f
C992 B.n952 VSUBS 0.007183f
C993 B.n953 VSUBS 0.007183f
C994 B.n954 VSUBS 0.007183f
C995 B.n955 VSUBS 0.007183f
C996 B.n956 VSUBS 0.007183f
C997 B.n957 VSUBS 0.007183f
C998 B.n958 VSUBS 0.007183f
C999 B.n959 VSUBS 0.007183f
C1000 B.n960 VSUBS 0.007183f
C1001 B.n961 VSUBS 0.007183f
C1002 B.n962 VSUBS 0.007183f
C1003 B.n963 VSUBS 0.007183f
C1004 B.n964 VSUBS 0.007183f
C1005 B.n965 VSUBS 0.007183f
C1006 B.n966 VSUBS 0.007183f
C1007 B.n967 VSUBS 0.007183f
C1008 B.n968 VSUBS 0.007183f
C1009 B.n969 VSUBS 0.007183f
C1010 B.n970 VSUBS 0.007183f
C1011 B.n971 VSUBS 0.009373f
C1012 B.n972 VSUBS 0.009985f
C1013 B.n973 VSUBS 0.019856f
C1014 VDD2.t2 VSUBS 4.21044f
C1015 VDD2.t5 VSUBS 0.387983f
C1016 VDD2.t0 VSUBS 0.387983f
C1017 VDD2.n0 VSUBS 3.232f
C1018 VDD2.n1 VSUBS 4.79774f
C1019 VDD2.t3 VSUBS 4.17921f
C1020 VDD2.n2 VSUBS 4.25623f
C1021 VDD2.t1 VSUBS 0.387983f
C1022 VDD2.t4 VSUBS 0.387983f
C1023 VDD2.n3 VSUBS 3.23195f
C1024 VN.t5 VSUBS 4.09836f
C1025 VN.n0 VSUBS 1.49762f
C1026 VN.n1 VSUBS 0.022036f
C1027 VN.n2 VSUBS 0.042204f
C1028 VN.n3 VSUBS 0.022036f
C1029 VN.n4 VSUBS 0.04107f
C1030 VN.t0 VSUBS 4.09836f
C1031 VN.n5 VSUBS 1.503f
C1032 VN.t3 VSUBS 4.45896f
C1033 VN.n6 VSUBS 1.42757f
C1034 VN.n7 VSUBS 0.281517f
C1035 VN.n8 VSUBS 0.022036f
C1036 VN.n9 VSUBS 0.04107f
C1037 VN.n10 VSUBS 0.044521f
C1038 VN.n11 VSUBS 0.018686f
C1039 VN.n12 VSUBS 0.022036f
C1040 VN.n13 VSUBS 0.022036f
C1041 VN.n14 VSUBS 0.022036f
C1042 VN.n15 VSUBS 0.04107f
C1043 VN.n16 VSUBS 0.04107f
C1044 VN.n17 VSUBS 0.025254f
C1045 VN.n18 VSUBS 0.035566f
C1046 VN.n19 VSUBS 0.065748f
C1047 VN.t2 VSUBS 4.09836f
C1048 VN.n20 VSUBS 1.49762f
C1049 VN.n21 VSUBS 0.022036f
C1050 VN.n22 VSUBS 0.042204f
C1051 VN.n23 VSUBS 0.022036f
C1052 VN.n24 VSUBS 0.04107f
C1053 VN.t1 VSUBS 4.45896f
C1054 VN.t4 VSUBS 4.09836f
C1055 VN.n25 VSUBS 1.503f
C1056 VN.n26 VSUBS 1.42757f
C1057 VN.n27 VSUBS 0.281517f
C1058 VN.n28 VSUBS 0.022036f
C1059 VN.n29 VSUBS 0.04107f
C1060 VN.n30 VSUBS 0.044521f
C1061 VN.n31 VSUBS 0.018686f
C1062 VN.n32 VSUBS 0.022036f
C1063 VN.n33 VSUBS 0.022036f
C1064 VN.n34 VSUBS 0.022036f
C1065 VN.n35 VSUBS 0.04107f
C1066 VN.n36 VSUBS 0.04107f
C1067 VN.n37 VSUBS 0.025254f
C1068 VN.n38 VSUBS 0.035566f
C1069 VN.n39 VSUBS 1.55815f
C1070 VDD1.t5 VSUBS 4.21191f
C1071 VDD1.t3 VSUBS 4.21023f
C1072 VDD1.t4 VSUBS 0.387963f
C1073 VDD1.t0 VSUBS 0.387963f
C1074 VDD1.n0 VSUBS 3.23184f
C1075 VDD1.n1 VSUBS 4.97365f
C1076 VDD1.t2 VSUBS 0.387963f
C1077 VDD1.t1 VSUBS 0.387963f
C1078 VDD1.n2 VSUBS 3.22067f
C1079 VDD1.n3 VSUBS 4.22783f
C1080 VTAIL.t0 VSUBS 0.399356f
C1081 VTAIL.t1 VSUBS 0.399356f
C1082 VTAIL.n0 VSUBS 3.1397f
C1083 VTAIL.n1 VSUBS 0.983661f
C1084 VTAIL.t7 VSUBS 4.10043f
C1085 VTAIL.n2 VSUBS 1.34866f
C1086 VTAIL.t11 VSUBS 0.399356f
C1087 VTAIL.t10 VSUBS 0.399356f
C1088 VTAIL.n3 VSUBS 3.1397f
C1089 VTAIL.n4 VSUBS 3.44875f
C1090 VTAIL.t4 VSUBS 0.399356f
C1091 VTAIL.t3 VSUBS 0.399356f
C1092 VTAIL.n5 VSUBS 3.1397f
C1093 VTAIL.n6 VSUBS 3.44875f
C1094 VTAIL.t5 VSUBS 4.10044f
C1095 VTAIL.n7 VSUBS 1.34865f
C1096 VTAIL.t8 VSUBS 0.399356f
C1097 VTAIL.t9 VSUBS 0.399356f
C1098 VTAIL.n8 VSUBS 3.1397f
C1099 VTAIL.n9 VSUBS 1.22024f
C1100 VTAIL.t6 VSUBS 4.10043f
C1101 VTAIL.n10 VSUBS 3.25467f
C1102 VTAIL.t2 VSUBS 4.10043f
C1103 VTAIL.n11 VSUBS 3.16874f
C1104 VP.t5 VSUBS 4.45048f
C1105 VP.n0 VSUBS 1.6263f
C1106 VP.n1 VSUBS 0.023929f
C1107 VP.n2 VSUBS 0.04583f
C1108 VP.n3 VSUBS 0.023929f
C1109 VP.n4 VSUBS 0.044598f
C1110 VP.n5 VSUBS 0.023929f
C1111 VP.t1 VSUBS 4.45048f
C1112 VP.n6 VSUBS 0.048346f
C1113 VP.n7 VSUBS 0.023929f
C1114 VP.n8 VSUBS 0.044598f
C1115 VP.t4 VSUBS 4.45048f
C1116 VP.n9 VSUBS 1.6263f
C1117 VP.n10 VSUBS 0.023929f
C1118 VP.n11 VSUBS 0.04583f
C1119 VP.n12 VSUBS 0.023929f
C1120 VP.n13 VSUBS 0.044598f
C1121 VP.t0 VSUBS 4.84206f
C1122 VP.t3 VSUBS 4.45048f
C1123 VP.n14 VSUBS 1.63214f
C1124 VP.n15 VSUBS 1.55023f
C1125 VP.n16 VSUBS 0.305705f
C1126 VP.n17 VSUBS 0.023929f
C1127 VP.n18 VSUBS 0.044598f
C1128 VP.n19 VSUBS 0.048346f
C1129 VP.n20 VSUBS 0.020292f
C1130 VP.n21 VSUBS 0.023929f
C1131 VP.n22 VSUBS 0.023929f
C1132 VP.n23 VSUBS 0.023929f
C1133 VP.n24 VSUBS 0.044598f
C1134 VP.n25 VSUBS 0.044598f
C1135 VP.n26 VSUBS 0.027424f
C1136 VP.n27 VSUBS 0.038622f
C1137 VP.n28 VSUBS 1.68269f
C1138 VP.n29 VSUBS 1.69756f
C1139 VP.t2 VSUBS 4.45048f
C1140 VP.n30 VSUBS 1.6263f
C1141 VP.n31 VSUBS 0.027424f
C1142 VP.n32 VSUBS 0.038622f
C1143 VP.n33 VSUBS 0.023929f
C1144 VP.n34 VSUBS 0.023929f
C1145 VP.n35 VSUBS 0.044598f
C1146 VP.n36 VSUBS 0.04583f
C1147 VP.n37 VSUBS 0.020292f
C1148 VP.n38 VSUBS 0.023929f
C1149 VP.n39 VSUBS 0.023929f
C1150 VP.n40 VSUBS 0.023929f
C1151 VP.n41 VSUBS 0.044598f
C1152 VP.n42 VSUBS 0.044598f
C1153 VP.n43 VSUBS 1.55626f
C1154 VP.n44 VSUBS 0.023929f
C1155 VP.n45 VSUBS 0.023929f
C1156 VP.n46 VSUBS 0.023929f
C1157 VP.n47 VSUBS 0.044598f
C1158 VP.n48 VSUBS 0.048346f
C1159 VP.n49 VSUBS 0.020292f
C1160 VP.n50 VSUBS 0.023929f
C1161 VP.n51 VSUBS 0.023929f
C1162 VP.n52 VSUBS 0.023929f
C1163 VP.n53 VSUBS 0.044598f
C1164 VP.n54 VSUBS 0.044598f
C1165 VP.n55 VSUBS 0.027424f
C1166 VP.n56 VSUBS 0.038622f
C1167 VP.n57 VSUBS 0.071397f
.ends

