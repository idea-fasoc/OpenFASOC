* NGSPICE file created from diff_pair_sample_0115.ext - technology: sky130A

.subckt diff_pair_sample_0115 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=0 ps=0 w=14.64 l=1.79
X1 VTAIL.t7 VP.t0 VDD1.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=2.4156 ps=14.97 w=14.64 l=1.79
X2 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=0 ps=0 w=14.64 l=1.79
X3 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=0 ps=0 w=14.64 l=1.79
X4 VDD1.t2 VP.t1 VTAIL.t6 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4156 pd=14.97 as=5.7096 ps=30.06 w=14.64 l=1.79
X5 VDD2.t3 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=2.4156 pd=14.97 as=5.7096 ps=30.06 w=14.64 l=1.79
X6 VTAIL.t2 VN.t1 VDD2.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=2.4156 ps=14.97 w=14.64 l=1.79
X7 VTAIL.t5 VP.t2 VDD1.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=2.4156 ps=14.97 w=14.64 l=1.79
X8 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=0 ps=0 w=14.64 l=1.79
X9 VTAIL.t1 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=5.7096 pd=30.06 as=2.4156 ps=14.97 w=14.64 l=1.79
X10 VDD1.t0 VP.t3 VTAIL.t4 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4156 pd=14.97 as=5.7096 ps=30.06 w=14.64 l=1.79
X11 VDD2.t0 VN.t3 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.4156 pd=14.97 as=5.7096 ps=30.06 w=14.64 l=1.79
R0 B.n766 B.n765 585
R1 B.n322 B.n106 585
R2 B.n321 B.n320 585
R3 B.n319 B.n318 585
R4 B.n317 B.n316 585
R5 B.n315 B.n314 585
R6 B.n313 B.n312 585
R7 B.n311 B.n310 585
R8 B.n309 B.n308 585
R9 B.n307 B.n306 585
R10 B.n305 B.n304 585
R11 B.n303 B.n302 585
R12 B.n301 B.n300 585
R13 B.n299 B.n298 585
R14 B.n297 B.n296 585
R15 B.n295 B.n294 585
R16 B.n293 B.n292 585
R17 B.n291 B.n290 585
R18 B.n289 B.n288 585
R19 B.n287 B.n286 585
R20 B.n285 B.n284 585
R21 B.n283 B.n282 585
R22 B.n281 B.n280 585
R23 B.n279 B.n278 585
R24 B.n277 B.n276 585
R25 B.n275 B.n274 585
R26 B.n273 B.n272 585
R27 B.n271 B.n270 585
R28 B.n269 B.n268 585
R29 B.n267 B.n266 585
R30 B.n265 B.n264 585
R31 B.n263 B.n262 585
R32 B.n261 B.n260 585
R33 B.n259 B.n258 585
R34 B.n257 B.n256 585
R35 B.n255 B.n254 585
R36 B.n253 B.n252 585
R37 B.n251 B.n250 585
R38 B.n249 B.n248 585
R39 B.n247 B.n246 585
R40 B.n245 B.n244 585
R41 B.n243 B.n242 585
R42 B.n241 B.n240 585
R43 B.n239 B.n238 585
R44 B.n237 B.n236 585
R45 B.n235 B.n234 585
R46 B.n233 B.n232 585
R47 B.n231 B.n230 585
R48 B.n229 B.n228 585
R49 B.n226 B.n225 585
R50 B.n224 B.n223 585
R51 B.n222 B.n221 585
R52 B.n220 B.n219 585
R53 B.n218 B.n217 585
R54 B.n216 B.n215 585
R55 B.n214 B.n213 585
R56 B.n212 B.n211 585
R57 B.n210 B.n209 585
R58 B.n208 B.n207 585
R59 B.n205 B.n204 585
R60 B.n203 B.n202 585
R61 B.n201 B.n200 585
R62 B.n199 B.n198 585
R63 B.n197 B.n196 585
R64 B.n195 B.n194 585
R65 B.n193 B.n192 585
R66 B.n191 B.n190 585
R67 B.n189 B.n188 585
R68 B.n187 B.n186 585
R69 B.n185 B.n184 585
R70 B.n183 B.n182 585
R71 B.n181 B.n180 585
R72 B.n179 B.n178 585
R73 B.n177 B.n176 585
R74 B.n175 B.n174 585
R75 B.n173 B.n172 585
R76 B.n171 B.n170 585
R77 B.n169 B.n168 585
R78 B.n167 B.n166 585
R79 B.n165 B.n164 585
R80 B.n163 B.n162 585
R81 B.n161 B.n160 585
R82 B.n159 B.n158 585
R83 B.n157 B.n156 585
R84 B.n155 B.n154 585
R85 B.n153 B.n152 585
R86 B.n151 B.n150 585
R87 B.n149 B.n148 585
R88 B.n147 B.n146 585
R89 B.n145 B.n144 585
R90 B.n143 B.n142 585
R91 B.n141 B.n140 585
R92 B.n139 B.n138 585
R93 B.n137 B.n136 585
R94 B.n135 B.n134 585
R95 B.n133 B.n132 585
R96 B.n131 B.n130 585
R97 B.n129 B.n128 585
R98 B.n127 B.n126 585
R99 B.n125 B.n124 585
R100 B.n123 B.n122 585
R101 B.n121 B.n120 585
R102 B.n119 B.n118 585
R103 B.n117 B.n116 585
R104 B.n115 B.n114 585
R105 B.n113 B.n112 585
R106 B.n53 B.n52 585
R107 B.n771 B.n770 585
R108 B.n764 B.n107 585
R109 B.n107 B.n50 585
R110 B.n763 B.n49 585
R111 B.n775 B.n49 585
R112 B.n762 B.n48 585
R113 B.n776 B.n48 585
R114 B.n761 B.n47 585
R115 B.n777 B.n47 585
R116 B.n760 B.n759 585
R117 B.n759 B.n43 585
R118 B.n758 B.n42 585
R119 B.n783 B.n42 585
R120 B.n757 B.n41 585
R121 B.n784 B.n41 585
R122 B.n756 B.n40 585
R123 B.n785 B.n40 585
R124 B.n755 B.n754 585
R125 B.n754 B.n36 585
R126 B.n753 B.n35 585
R127 B.n791 B.n35 585
R128 B.n752 B.n34 585
R129 B.n792 B.n34 585
R130 B.n751 B.n33 585
R131 B.n793 B.n33 585
R132 B.n750 B.n749 585
R133 B.n749 B.n29 585
R134 B.n748 B.n28 585
R135 B.n799 B.n28 585
R136 B.n747 B.n27 585
R137 B.n800 B.n27 585
R138 B.n746 B.n26 585
R139 B.n801 B.n26 585
R140 B.n745 B.n744 585
R141 B.n744 B.n25 585
R142 B.n743 B.n21 585
R143 B.n807 B.n21 585
R144 B.n742 B.n20 585
R145 B.n808 B.n20 585
R146 B.n741 B.n19 585
R147 B.n809 B.n19 585
R148 B.n740 B.n739 585
R149 B.n739 B.n15 585
R150 B.n738 B.n14 585
R151 B.n815 B.n14 585
R152 B.n737 B.n13 585
R153 B.n816 B.n13 585
R154 B.n736 B.n12 585
R155 B.n817 B.n12 585
R156 B.n735 B.n734 585
R157 B.n734 B.n8 585
R158 B.n733 B.n7 585
R159 B.n823 B.n7 585
R160 B.n732 B.n6 585
R161 B.n824 B.n6 585
R162 B.n731 B.n5 585
R163 B.n825 B.n5 585
R164 B.n730 B.n729 585
R165 B.n729 B.n4 585
R166 B.n728 B.n323 585
R167 B.n728 B.n727 585
R168 B.n718 B.n324 585
R169 B.n325 B.n324 585
R170 B.n720 B.n719 585
R171 B.n721 B.n720 585
R172 B.n717 B.n329 585
R173 B.n333 B.n329 585
R174 B.n716 B.n715 585
R175 B.n715 B.n714 585
R176 B.n331 B.n330 585
R177 B.n332 B.n331 585
R178 B.n707 B.n706 585
R179 B.n708 B.n707 585
R180 B.n705 B.n338 585
R181 B.n338 B.n337 585
R182 B.n704 B.n703 585
R183 B.n703 B.n702 585
R184 B.n340 B.n339 585
R185 B.n695 B.n340 585
R186 B.n694 B.n693 585
R187 B.n696 B.n694 585
R188 B.n692 B.n345 585
R189 B.n345 B.n344 585
R190 B.n691 B.n690 585
R191 B.n690 B.n689 585
R192 B.n347 B.n346 585
R193 B.n348 B.n347 585
R194 B.n682 B.n681 585
R195 B.n683 B.n682 585
R196 B.n680 B.n353 585
R197 B.n353 B.n352 585
R198 B.n679 B.n678 585
R199 B.n678 B.n677 585
R200 B.n355 B.n354 585
R201 B.n356 B.n355 585
R202 B.n670 B.n669 585
R203 B.n671 B.n670 585
R204 B.n668 B.n360 585
R205 B.n364 B.n360 585
R206 B.n667 B.n666 585
R207 B.n666 B.n665 585
R208 B.n362 B.n361 585
R209 B.n363 B.n362 585
R210 B.n658 B.n657 585
R211 B.n659 B.n658 585
R212 B.n656 B.n369 585
R213 B.n369 B.n368 585
R214 B.n655 B.n654 585
R215 B.n654 B.n653 585
R216 B.n371 B.n370 585
R217 B.n372 B.n371 585
R218 B.n649 B.n648 585
R219 B.n375 B.n374 585
R220 B.n645 B.n644 585
R221 B.n646 B.n645 585
R222 B.n643 B.n429 585
R223 B.n642 B.n641 585
R224 B.n640 B.n639 585
R225 B.n638 B.n637 585
R226 B.n636 B.n635 585
R227 B.n634 B.n633 585
R228 B.n632 B.n631 585
R229 B.n630 B.n629 585
R230 B.n628 B.n627 585
R231 B.n626 B.n625 585
R232 B.n624 B.n623 585
R233 B.n622 B.n621 585
R234 B.n620 B.n619 585
R235 B.n618 B.n617 585
R236 B.n616 B.n615 585
R237 B.n614 B.n613 585
R238 B.n612 B.n611 585
R239 B.n610 B.n609 585
R240 B.n608 B.n607 585
R241 B.n606 B.n605 585
R242 B.n604 B.n603 585
R243 B.n602 B.n601 585
R244 B.n600 B.n599 585
R245 B.n598 B.n597 585
R246 B.n596 B.n595 585
R247 B.n594 B.n593 585
R248 B.n592 B.n591 585
R249 B.n590 B.n589 585
R250 B.n588 B.n587 585
R251 B.n586 B.n585 585
R252 B.n584 B.n583 585
R253 B.n582 B.n581 585
R254 B.n580 B.n579 585
R255 B.n578 B.n577 585
R256 B.n576 B.n575 585
R257 B.n574 B.n573 585
R258 B.n572 B.n571 585
R259 B.n570 B.n569 585
R260 B.n568 B.n567 585
R261 B.n566 B.n565 585
R262 B.n564 B.n563 585
R263 B.n562 B.n561 585
R264 B.n560 B.n559 585
R265 B.n558 B.n557 585
R266 B.n556 B.n555 585
R267 B.n554 B.n553 585
R268 B.n552 B.n551 585
R269 B.n550 B.n549 585
R270 B.n548 B.n547 585
R271 B.n546 B.n545 585
R272 B.n544 B.n543 585
R273 B.n542 B.n541 585
R274 B.n540 B.n539 585
R275 B.n538 B.n537 585
R276 B.n536 B.n535 585
R277 B.n534 B.n533 585
R278 B.n532 B.n531 585
R279 B.n530 B.n529 585
R280 B.n528 B.n527 585
R281 B.n526 B.n525 585
R282 B.n524 B.n523 585
R283 B.n522 B.n521 585
R284 B.n520 B.n519 585
R285 B.n518 B.n517 585
R286 B.n516 B.n515 585
R287 B.n514 B.n513 585
R288 B.n512 B.n511 585
R289 B.n510 B.n509 585
R290 B.n508 B.n507 585
R291 B.n506 B.n505 585
R292 B.n504 B.n503 585
R293 B.n502 B.n501 585
R294 B.n500 B.n499 585
R295 B.n498 B.n497 585
R296 B.n496 B.n495 585
R297 B.n494 B.n493 585
R298 B.n492 B.n491 585
R299 B.n490 B.n489 585
R300 B.n488 B.n487 585
R301 B.n486 B.n485 585
R302 B.n484 B.n483 585
R303 B.n482 B.n481 585
R304 B.n480 B.n479 585
R305 B.n478 B.n477 585
R306 B.n476 B.n475 585
R307 B.n474 B.n473 585
R308 B.n472 B.n471 585
R309 B.n470 B.n469 585
R310 B.n468 B.n467 585
R311 B.n466 B.n465 585
R312 B.n464 B.n463 585
R313 B.n462 B.n461 585
R314 B.n460 B.n459 585
R315 B.n458 B.n457 585
R316 B.n456 B.n455 585
R317 B.n454 B.n453 585
R318 B.n452 B.n451 585
R319 B.n450 B.n449 585
R320 B.n448 B.n447 585
R321 B.n446 B.n445 585
R322 B.n444 B.n443 585
R323 B.n442 B.n441 585
R324 B.n440 B.n439 585
R325 B.n438 B.n437 585
R326 B.n436 B.n428 585
R327 B.n646 B.n428 585
R328 B.n650 B.n373 585
R329 B.n373 B.n372 585
R330 B.n652 B.n651 585
R331 B.n653 B.n652 585
R332 B.n367 B.n366 585
R333 B.n368 B.n367 585
R334 B.n661 B.n660 585
R335 B.n660 B.n659 585
R336 B.n662 B.n365 585
R337 B.n365 B.n363 585
R338 B.n664 B.n663 585
R339 B.n665 B.n664 585
R340 B.n359 B.n358 585
R341 B.n364 B.n359 585
R342 B.n673 B.n672 585
R343 B.n672 B.n671 585
R344 B.n674 B.n357 585
R345 B.n357 B.n356 585
R346 B.n676 B.n675 585
R347 B.n677 B.n676 585
R348 B.n351 B.n350 585
R349 B.n352 B.n351 585
R350 B.n685 B.n684 585
R351 B.n684 B.n683 585
R352 B.n686 B.n349 585
R353 B.n349 B.n348 585
R354 B.n688 B.n687 585
R355 B.n689 B.n688 585
R356 B.n343 B.n342 585
R357 B.n344 B.n343 585
R358 B.n698 B.n697 585
R359 B.n697 B.n696 585
R360 B.n699 B.n341 585
R361 B.n695 B.n341 585
R362 B.n701 B.n700 585
R363 B.n702 B.n701 585
R364 B.n336 B.n335 585
R365 B.n337 B.n336 585
R366 B.n710 B.n709 585
R367 B.n709 B.n708 585
R368 B.n711 B.n334 585
R369 B.n334 B.n332 585
R370 B.n713 B.n712 585
R371 B.n714 B.n713 585
R372 B.n328 B.n327 585
R373 B.n333 B.n328 585
R374 B.n723 B.n722 585
R375 B.n722 B.n721 585
R376 B.n724 B.n326 585
R377 B.n326 B.n325 585
R378 B.n726 B.n725 585
R379 B.n727 B.n726 585
R380 B.n2 B.n0 585
R381 B.n4 B.n2 585
R382 B.n3 B.n1 585
R383 B.n824 B.n3 585
R384 B.n822 B.n821 585
R385 B.n823 B.n822 585
R386 B.n820 B.n9 585
R387 B.n9 B.n8 585
R388 B.n819 B.n818 585
R389 B.n818 B.n817 585
R390 B.n11 B.n10 585
R391 B.n816 B.n11 585
R392 B.n814 B.n813 585
R393 B.n815 B.n814 585
R394 B.n812 B.n16 585
R395 B.n16 B.n15 585
R396 B.n811 B.n810 585
R397 B.n810 B.n809 585
R398 B.n18 B.n17 585
R399 B.n808 B.n18 585
R400 B.n806 B.n805 585
R401 B.n807 B.n806 585
R402 B.n804 B.n22 585
R403 B.n25 B.n22 585
R404 B.n803 B.n802 585
R405 B.n802 B.n801 585
R406 B.n24 B.n23 585
R407 B.n800 B.n24 585
R408 B.n798 B.n797 585
R409 B.n799 B.n798 585
R410 B.n796 B.n30 585
R411 B.n30 B.n29 585
R412 B.n795 B.n794 585
R413 B.n794 B.n793 585
R414 B.n32 B.n31 585
R415 B.n792 B.n32 585
R416 B.n790 B.n789 585
R417 B.n791 B.n790 585
R418 B.n788 B.n37 585
R419 B.n37 B.n36 585
R420 B.n787 B.n786 585
R421 B.n786 B.n785 585
R422 B.n39 B.n38 585
R423 B.n784 B.n39 585
R424 B.n782 B.n781 585
R425 B.n783 B.n782 585
R426 B.n780 B.n44 585
R427 B.n44 B.n43 585
R428 B.n779 B.n778 585
R429 B.n778 B.n777 585
R430 B.n46 B.n45 585
R431 B.n776 B.n46 585
R432 B.n774 B.n773 585
R433 B.n775 B.n774 585
R434 B.n772 B.n51 585
R435 B.n51 B.n50 585
R436 B.n827 B.n826 585
R437 B.n826 B.n825 585
R438 B.n648 B.n373 497.305
R439 B.n770 B.n51 497.305
R440 B.n428 B.n371 497.305
R441 B.n766 B.n107 497.305
R442 B.n433 B.t8 403.486
R443 B.n430 B.t12 403.486
R444 B.n110 B.t15 403.486
R445 B.n108 B.t4 403.486
R446 B.n433 B.t11 368.421
R447 B.n108 B.t6 368.421
R448 B.n430 B.t14 368.421
R449 B.n110 B.t16 368.421
R450 B.n434 B.t10 327.307
R451 B.n109 B.t7 327.307
R452 B.n431 B.t13 327.307
R453 B.n111 B.t17 327.307
R454 B.n768 B.n767 256.663
R455 B.n768 B.n105 256.663
R456 B.n768 B.n104 256.663
R457 B.n768 B.n103 256.663
R458 B.n768 B.n102 256.663
R459 B.n768 B.n101 256.663
R460 B.n768 B.n100 256.663
R461 B.n768 B.n99 256.663
R462 B.n768 B.n98 256.663
R463 B.n768 B.n97 256.663
R464 B.n768 B.n96 256.663
R465 B.n768 B.n95 256.663
R466 B.n768 B.n94 256.663
R467 B.n768 B.n93 256.663
R468 B.n768 B.n92 256.663
R469 B.n768 B.n91 256.663
R470 B.n768 B.n90 256.663
R471 B.n768 B.n89 256.663
R472 B.n768 B.n88 256.663
R473 B.n768 B.n87 256.663
R474 B.n768 B.n86 256.663
R475 B.n768 B.n85 256.663
R476 B.n768 B.n84 256.663
R477 B.n768 B.n83 256.663
R478 B.n768 B.n82 256.663
R479 B.n768 B.n81 256.663
R480 B.n768 B.n80 256.663
R481 B.n768 B.n79 256.663
R482 B.n768 B.n78 256.663
R483 B.n768 B.n77 256.663
R484 B.n768 B.n76 256.663
R485 B.n768 B.n75 256.663
R486 B.n768 B.n74 256.663
R487 B.n768 B.n73 256.663
R488 B.n768 B.n72 256.663
R489 B.n768 B.n71 256.663
R490 B.n768 B.n70 256.663
R491 B.n768 B.n69 256.663
R492 B.n768 B.n68 256.663
R493 B.n768 B.n67 256.663
R494 B.n768 B.n66 256.663
R495 B.n768 B.n65 256.663
R496 B.n768 B.n64 256.663
R497 B.n768 B.n63 256.663
R498 B.n768 B.n62 256.663
R499 B.n768 B.n61 256.663
R500 B.n768 B.n60 256.663
R501 B.n768 B.n59 256.663
R502 B.n768 B.n58 256.663
R503 B.n768 B.n57 256.663
R504 B.n768 B.n56 256.663
R505 B.n768 B.n55 256.663
R506 B.n768 B.n54 256.663
R507 B.n769 B.n768 256.663
R508 B.n647 B.n646 256.663
R509 B.n646 B.n376 256.663
R510 B.n646 B.n377 256.663
R511 B.n646 B.n378 256.663
R512 B.n646 B.n379 256.663
R513 B.n646 B.n380 256.663
R514 B.n646 B.n381 256.663
R515 B.n646 B.n382 256.663
R516 B.n646 B.n383 256.663
R517 B.n646 B.n384 256.663
R518 B.n646 B.n385 256.663
R519 B.n646 B.n386 256.663
R520 B.n646 B.n387 256.663
R521 B.n646 B.n388 256.663
R522 B.n646 B.n389 256.663
R523 B.n646 B.n390 256.663
R524 B.n646 B.n391 256.663
R525 B.n646 B.n392 256.663
R526 B.n646 B.n393 256.663
R527 B.n646 B.n394 256.663
R528 B.n646 B.n395 256.663
R529 B.n646 B.n396 256.663
R530 B.n646 B.n397 256.663
R531 B.n646 B.n398 256.663
R532 B.n646 B.n399 256.663
R533 B.n646 B.n400 256.663
R534 B.n646 B.n401 256.663
R535 B.n646 B.n402 256.663
R536 B.n646 B.n403 256.663
R537 B.n646 B.n404 256.663
R538 B.n646 B.n405 256.663
R539 B.n646 B.n406 256.663
R540 B.n646 B.n407 256.663
R541 B.n646 B.n408 256.663
R542 B.n646 B.n409 256.663
R543 B.n646 B.n410 256.663
R544 B.n646 B.n411 256.663
R545 B.n646 B.n412 256.663
R546 B.n646 B.n413 256.663
R547 B.n646 B.n414 256.663
R548 B.n646 B.n415 256.663
R549 B.n646 B.n416 256.663
R550 B.n646 B.n417 256.663
R551 B.n646 B.n418 256.663
R552 B.n646 B.n419 256.663
R553 B.n646 B.n420 256.663
R554 B.n646 B.n421 256.663
R555 B.n646 B.n422 256.663
R556 B.n646 B.n423 256.663
R557 B.n646 B.n424 256.663
R558 B.n646 B.n425 256.663
R559 B.n646 B.n426 256.663
R560 B.n646 B.n427 256.663
R561 B.n652 B.n373 163.367
R562 B.n652 B.n367 163.367
R563 B.n660 B.n367 163.367
R564 B.n660 B.n365 163.367
R565 B.n664 B.n365 163.367
R566 B.n664 B.n359 163.367
R567 B.n672 B.n359 163.367
R568 B.n672 B.n357 163.367
R569 B.n676 B.n357 163.367
R570 B.n676 B.n351 163.367
R571 B.n684 B.n351 163.367
R572 B.n684 B.n349 163.367
R573 B.n688 B.n349 163.367
R574 B.n688 B.n343 163.367
R575 B.n697 B.n343 163.367
R576 B.n697 B.n341 163.367
R577 B.n701 B.n341 163.367
R578 B.n701 B.n336 163.367
R579 B.n709 B.n336 163.367
R580 B.n709 B.n334 163.367
R581 B.n713 B.n334 163.367
R582 B.n713 B.n328 163.367
R583 B.n722 B.n328 163.367
R584 B.n722 B.n326 163.367
R585 B.n726 B.n326 163.367
R586 B.n726 B.n2 163.367
R587 B.n826 B.n2 163.367
R588 B.n826 B.n3 163.367
R589 B.n822 B.n3 163.367
R590 B.n822 B.n9 163.367
R591 B.n818 B.n9 163.367
R592 B.n818 B.n11 163.367
R593 B.n814 B.n11 163.367
R594 B.n814 B.n16 163.367
R595 B.n810 B.n16 163.367
R596 B.n810 B.n18 163.367
R597 B.n806 B.n18 163.367
R598 B.n806 B.n22 163.367
R599 B.n802 B.n22 163.367
R600 B.n802 B.n24 163.367
R601 B.n798 B.n24 163.367
R602 B.n798 B.n30 163.367
R603 B.n794 B.n30 163.367
R604 B.n794 B.n32 163.367
R605 B.n790 B.n32 163.367
R606 B.n790 B.n37 163.367
R607 B.n786 B.n37 163.367
R608 B.n786 B.n39 163.367
R609 B.n782 B.n39 163.367
R610 B.n782 B.n44 163.367
R611 B.n778 B.n44 163.367
R612 B.n778 B.n46 163.367
R613 B.n774 B.n46 163.367
R614 B.n774 B.n51 163.367
R615 B.n645 B.n375 163.367
R616 B.n645 B.n429 163.367
R617 B.n641 B.n640 163.367
R618 B.n637 B.n636 163.367
R619 B.n633 B.n632 163.367
R620 B.n629 B.n628 163.367
R621 B.n625 B.n624 163.367
R622 B.n621 B.n620 163.367
R623 B.n617 B.n616 163.367
R624 B.n613 B.n612 163.367
R625 B.n609 B.n608 163.367
R626 B.n605 B.n604 163.367
R627 B.n601 B.n600 163.367
R628 B.n597 B.n596 163.367
R629 B.n593 B.n592 163.367
R630 B.n589 B.n588 163.367
R631 B.n585 B.n584 163.367
R632 B.n581 B.n580 163.367
R633 B.n577 B.n576 163.367
R634 B.n573 B.n572 163.367
R635 B.n569 B.n568 163.367
R636 B.n565 B.n564 163.367
R637 B.n561 B.n560 163.367
R638 B.n557 B.n556 163.367
R639 B.n553 B.n552 163.367
R640 B.n549 B.n548 163.367
R641 B.n545 B.n544 163.367
R642 B.n541 B.n540 163.367
R643 B.n537 B.n536 163.367
R644 B.n533 B.n532 163.367
R645 B.n529 B.n528 163.367
R646 B.n525 B.n524 163.367
R647 B.n521 B.n520 163.367
R648 B.n517 B.n516 163.367
R649 B.n513 B.n512 163.367
R650 B.n509 B.n508 163.367
R651 B.n505 B.n504 163.367
R652 B.n501 B.n500 163.367
R653 B.n497 B.n496 163.367
R654 B.n493 B.n492 163.367
R655 B.n489 B.n488 163.367
R656 B.n485 B.n484 163.367
R657 B.n481 B.n480 163.367
R658 B.n477 B.n476 163.367
R659 B.n473 B.n472 163.367
R660 B.n469 B.n468 163.367
R661 B.n465 B.n464 163.367
R662 B.n461 B.n460 163.367
R663 B.n457 B.n456 163.367
R664 B.n453 B.n452 163.367
R665 B.n449 B.n448 163.367
R666 B.n445 B.n444 163.367
R667 B.n441 B.n440 163.367
R668 B.n437 B.n428 163.367
R669 B.n654 B.n371 163.367
R670 B.n654 B.n369 163.367
R671 B.n658 B.n369 163.367
R672 B.n658 B.n362 163.367
R673 B.n666 B.n362 163.367
R674 B.n666 B.n360 163.367
R675 B.n670 B.n360 163.367
R676 B.n670 B.n355 163.367
R677 B.n678 B.n355 163.367
R678 B.n678 B.n353 163.367
R679 B.n682 B.n353 163.367
R680 B.n682 B.n347 163.367
R681 B.n690 B.n347 163.367
R682 B.n690 B.n345 163.367
R683 B.n694 B.n345 163.367
R684 B.n694 B.n340 163.367
R685 B.n703 B.n340 163.367
R686 B.n703 B.n338 163.367
R687 B.n707 B.n338 163.367
R688 B.n707 B.n331 163.367
R689 B.n715 B.n331 163.367
R690 B.n715 B.n329 163.367
R691 B.n720 B.n329 163.367
R692 B.n720 B.n324 163.367
R693 B.n728 B.n324 163.367
R694 B.n729 B.n728 163.367
R695 B.n729 B.n5 163.367
R696 B.n6 B.n5 163.367
R697 B.n7 B.n6 163.367
R698 B.n734 B.n7 163.367
R699 B.n734 B.n12 163.367
R700 B.n13 B.n12 163.367
R701 B.n14 B.n13 163.367
R702 B.n739 B.n14 163.367
R703 B.n739 B.n19 163.367
R704 B.n20 B.n19 163.367
R705 B.n21 B.n20 163.367
R706 B.n744 B.n21 163.367
R707 B.n744 B.n26 163.367
R708 B.n27 B.n26 163.367
R709 B.n28 B.n27 163.367
R710 B.n749 B.n28 163.367
R711 B.n749 B.n33 163.367
R712 B.n34 B.n33 163.367
R713 B.n35 B.n34 163.367
R714 B.n754 B.n35 163.367
R715 B.n754 B.n40 163.367
R716 B.n41 B.n40 163.367
R717 B.n42 B.n41 163.367
R718 B.n759 B.n42 163.367
R719 B.n759 B.n47 163.367
R720 B.n48 B.n47 163.367
R721 B.n49 B.n48 163.367
R722 B.n107 B.n49 163.367
R723 B.n112 B.n53 163.367
R724 B.n116 B.n115 163.367
R725 B.n120 B.n119 163.367
R726 B.n124 B.n123 163.367
R727 B.n128 B.n127 163.367
R728 B.n132 B.n131 163.367
R729 B.n136 B.n135 163.367
R730 B.n140 B.n139 163.367
R731 B.n144 B.n143 163.367
R732 B.n148 B.n147 163.367
R733 B.n152 B.n151 163.367
R734 B.n156 B.n155 163.367
R735 B.n160 B.n159 163.367
R736 B.n164 B.n163 163.367
R737 B.n168 B.n167 163.367
R738 B.n172 B.n171 163.367
R739 B.n176 B.n175 163.367
R740 B.n180 B.n179 163.367
R741 B.n184 B.n183 163.367
R742 B.n188 B.n187 163.367
R743 B.n192 B.n191 163.367
R744 B.n196 B.n195 163.367
R745 B.n200 B.n199 163.367
R746 B.n204 B.n203 163.367
R747 B.n209 B.n208 163.367
R748 B.n213 B.n212 163.367
R749 B.n217 B.n216 163.367
R750 B.n221 B.n220 163.367
R751 B.n225 B.n224 163.367
R752 B.n230 B.n229 163.367
R753 B.n234 B.n233 163.367
R754 B.n238 B.n237 163.367
R755 B.n242 B.n241 163.367
R756 B.n246 B.n245 163.367
R757 B.n250 B.n249 163.367
R758 B.n254 B.n253 163.367
R759 B.n258 B.n257 163.367
R760 B.n262 B.n261 163.367
R761 B.n266 B.n265 163.367
R762 B.n270 B.n269 163.367
R763 B.n274 B.n273 163.367
R764 B.n278 B.n277 163.367
R765 B.n282 B.n281 163.367
R766 B.n286 B.n285 163.367
R767 B.n290 B.n289 163.367
R768 B.n294 B.n293 163.367
R769 B.n298 B.n297 163.367
R770 B.n302 B.n301 163.367
R771 B.n306 B.n305 163.367
R772 B.n310 B.n309 163.367
R773 B.n314 B.n313 163.367
R774 B.n318 B.n317 163.367
R775 B.n320 B.n106 163.367
R776 B.n648 B.n647 71.676
R777 B.n429 B.n376 71.676
R778 B.n640 B.n377 71.676
R779 B.n636 B.n378 71.676
R780 B.n632 B.n379 71.676
R781 B.n628 B.n380 71.676
R782 B.n624 B.n381 71.676
R783 B.n620 B.n382 71.676
R784 B.n616 B.n383 71.676
R785 B.n612 B.n384 71.676
R786 B.n608 B.n385 71.676
R787 B.n604 B.n386 71.676
R788 B.n600 B.n387 71.676
R789 B.n596 B.n388 71.676
R790 B.n592 B.n389 71.676
R791 B.n588 B.n390 71.676
R792 B.n584 B.n391 71.676
R793 B.n580 B.n392 71.676
R794 B.n576 B.n393 71.676
R795 B.n572 B.n394 71.676
R796 B.n568 B.n395 71.676
R797 B.n564 B.n396 71.676
R798 B.n560 B.n397 71.676
R799 B.n556 B.n398 71.676
R800 B.n552 B.n399 71.676
R801 B.n548 B.n400 71.676
R802 B.n544 B.n401 71.676
R803 B.n540 B.n402 71.676
R804 B.n536 B.n403 71.676
R805 B.n532 B.n404 71.676
R806 B.n528 B.n405 71.676
R807 B.n524 B.n406 71.676
R808 B.n520 B.n407 71.676
R809 B.n516 B.n408 71.676
R810 B.n512 B.n409 71.676
R811 B.n508 B.n410 71.676
R812 B.n504 B.n411 71.676
R813 B.n500 B.n412 71.676
R814 B.n496 B.n413 71.676
R815 B.n492 B.n414 71.676
R816 B.n488 B.n415 71.676
R817 B.n484 B.n416 71.676
R818 B.n480 B.n417 71.676
R819 B.n476 B.n418 71.676
R820 B.n472 B.n419 71.676
R821 B.n468 B.n420 71.676
R822 B.n464 B.n421 71.676
R823 B.n460 B.n422 71.676
R824 B.n456 B.n423 71.676
R825 B.n452 B.n424 71.676
R826 B.n448 B.n425 71.676
R827 B.n444 B.n426 71.676
R828 B.n440 B.n427 71.676
R829 B.n770 B.n769 71.676
R830 B.n112 B.n54 71.676
R831 B.n116 B.n55 71.676
R832 B.n120 B.n56 71.676
R833 B.n124 B.n57 71.676
R834 B.n128 B.n58 71.676
R835 B.n132 B.n59 71.676
R836 B.n136 B.n60 71.676
R837 B.n140 B.n61 71.676
R838 B.n144 B.n62 71.676
R839 B.n148 B.n63 71.676
R840 B.n152 B.n64 71.676
R841 B.n156 B.n65 71.676
R842 B.n160 B.n66 71.676
R843 B.n164 B.n67 71.676
R844 B.n168 B.n68 71.676
R845 B.n172 B.n69 71.676
R846 B.n176 B.n70 71.676
R847 B.n180 B.n71 71.676
R848 B.n184 B.n72 71.676
R849 B.n188 B.n73 71.676
R850 B.n192 B.n74 71.676
R851 B.n196 B.n75 71.676
R852 B.n200 B.n76 71.676
R853 B.n204 B.n77 71.676
R854 B.n209 B.n78 71.676
R855 B.n213 B.n79 71.676
R856 B.n217 B.n80 71.676
R857 B.n221 B.n81 71.676
R858 B.n225 B.n82 71.676
R859 B.n230 B.n83 71.676
R860 B.n234 B.n84 71.676
R861 B.n238 B.n85 71.676
R862 B.n242 B.n86 71.676
R863 B.n246 B.n87 71.676
R864 B.n250 B.n88 71.676
R865 B.n254 B.n89 71.676
R866 B.n258 B.n90 71.676
R867 B.n262 B.n91 71.676
R868 B.n266 B.n92 71.676
R869 B.n270 B.n93 71.676
R870 B.n274 B.n94 71.676
R871 B.n278 B.n95 71.676
R872 B.n282 B.n96 71.676
R873 B.n286 B.n97 71.676
R874 B.n290 B.n98 71.676
R875 B.n294 B.n99 71.676
R876 B.n298 B.n100 71.676
R877 B.n302 B.n101 71.676
R878 B.n306 B.n102 71.676
R879 B.n310 B.n103 71.676
R880 B.n314 B.n104 71.676
R881 B.n318 B.n105 71.676
R882 B.n767 B.n106 71.676
R883 B.n767 B.n766 71.676
R884 B.n320 B.n105 71.676
R885 B.n317 B.n104 71.676
R886 B.n313 B.n103 71.676
R887 B.n309 B.n102 71.676
R888 B.n305 B.n101 71.676
R889 B.n301 B.n100 71.676
R890 B.n297 B.n99 71.676
R891 B.n293 B.n98 71.676
R892 B.n289 B.n97 71.676
R893 B.n285 B.n96 71.676
R894 B.n281 B.n95 71.676
R895 B.n277 B.n94 71.676
R896 B.n273 B.n93 71.676
R897 B.n269 B.n92 71.676
R898 B.n265 B.n91 71.676
R899 B.n261 B.n90 71.676
R900 B.n257 B.n89 71.676
R901 B.n253 B.n88 71.676
R902 B.n249 B.n87 71.676
R903 B.n245 B.n86 71.676
R904 B.n241 B.n85 71.676
R905 B.n237 B.n84 71.676
R906 B.n233 B.n83 71.676
R907 B.n229 B.n82 71.676
R908 B.n224 B.n81 71.676
R909 B.n220 B.n80 71.676
R910 B.n216 B.n79 71.676
R911 B.n212 B.n78 71.676
R912 B.n208 B.n77 71.676
R913 B.n203 B.n76 71.676
R914 B.n199 B.n75 71.676
R915 B.n195 B.n74 71.676
R916 B.n191 B.n73 71.676
R917 B.n187 B.n72 71.676
R918 B.n183 B.n71 71.676
R919 B.n179 B.n70 71.676
R920 B.n175 B.n69 71.676
R921 B.n171 B.n68 71.676
R922 B.n167 B.n67 71.676
R923 B.n163 B.n66 71.676
R924 B.n159 B.n65 71.676
R925 B.n155 B.n64 71.676
R926 B.n151 B.n63 71.676
R927 B.n147 B.n62 71.676
R928 B.n143 B.n61 71.676
R929 B.n139 B.n60 71.676
R930 B.n135 B.n59 71.676
R931 B.n131 B.n58 71.676
R932 B.n127 B.n57 71.676
R933 B.n123 B.n56 71.676
R934 B.n119 B.n55 71.676
R935 B.n115 B.n54 71.676
R936 B.n769 B.n53 71.676
R937 B.n647 B.n375 71.676
R938 B.n641 B.n376 71.676
R939 B.n637 B.n377 71.676
R940 B.n633 B.n378 71.676
R941 B.n629 B.n379 71.676
R942 B.n625 B.n380 71.676
R943 B.n621 B.n381 71.676
R944 B.n617 B.n382 71.676
R945 B.n613 B.n383 71.676
R946 B.n609 B.n384 71.676
R947 B.n605 B.n385 71.676
R948 B.n601 B.n386 71.676
R949 B.n597 B.n387 71.676
R950 B.n593 B.n388 71.676
R951 B.n589 B.n389 71.676
R952 B.n585 B.n390 71.676
R953 B.n581 B.n391 71.676
R954 B.n577 B.n392 71.676
R955 B.n573 B.n393 71.676
R956 B.n569 B.n394 71.676
R957 B.n565 B.n395 71.676
R958 B.n561 B.n396 71.676
R959 B.n557 B.n397 71.676
R960 B.n553 B.n398 71.676
R961 B.n549 B.n399 71.676
R962 B.n545 B.n400 71.676
R963 B.n541 B.n401 71.676
R964 B.n537 B.n402 71.676
R965 B.n533 B.n403 71.676
R966 B.n529 B.n404 71.676
R967 B.n525 B.n405 71.676
R968 B.n521 B.n406 71.676
R969 B.n517 B.n407 71.676
R970 B.n513 B.n408 71.676
R971 B.n509 B.n409 71.676
R972 B.n505 B.n410 71.676
R973 B.n501 B.n411 71.676
R974 B.n497 B.n412 71.676
R975 B.n493 B.n413 71.676
R976 B.n489 B.n414 71.676
R977 B.n485 B.n415 71.676
R978 B.n481 B.n416 71.676
R979 B.n477 B.n417 71.676
R980 B.n473 B.n418 71.676
R981 B.n469 B.n419 71.676
R982 B.n465 B.n420 71.676
R983 B.n461 B.n421 71.676
R984 B.n457 B.n422 71.676
R985 B.n453 B.n423 71.676
R986 B.n449 B.n424 71.676
R987 B.n445 B.n425 71.676
R988 B.n441 B.n426 71.676
R989 B.n437 B.n427 71.676
R990 B.n646 B.n372 61.3111
R991 B.n768 B.n50 61.3111
R992 B.n435 B.n434 59.5399
R993 B.n432 B.n431 59.5399
R994 B.n206 B.n111 59.5399
R995 B.n227 B.n109 59.5399
R996 B.n434 B.n433 41.1157
R997 B.n431 B.n430 41.1157
R998 B.n111 B.n110 41.1157
R999 B.n109 B.n108 41.1157
R1000 B.n653 B.n372 37.5601
R1001 B.n653 B.n368 37.5601
R1002 B.n659 B.n368 37.5601
R1003 B.n659 B.n363 37.5601
R1004 B.n665 B.n363 37.5601
R1005 B.n665 B.n364 37.5601
R1006 B.n671 B.n356 37.5601
R1007 B.n677 B.n356 37.5601
R1008 B.n677 B.n352 37.5601
R1009 B.n683 B.n352 37.5601
R1010 B.n683 B.n348 37.5601
R1011 B.n689 B.n348 37.5601
R1012 B.n689 B.n344 37.5601
R1013 B.n696 B.n344 37.5601
R1014 B.n696 B.n695 37.5601
R1015 B.n702 B.n337 37.5601
R1016 B.n708 B.n337 37.5601
R1017 B.n708 B.n332 37.5601
R1018 B.n714 B.n332 37.5601
R1019 B.n714 B.n333 37.5601
R1020 B.n721 B.n325 37.5601
R1021 B.n727 B.n325 37.5601
R1022 B.n727 B.n4 37.5601
R1023 B.n825 B.n4 37.5601
R1024 B.n825 B.n824 37.5601
R1025 B.n824 B.n823 37.5601
R1026 B.n823 B.n8 37.5601
R1027 B.n817 B.n8 37.5601
R1028 B.n816 B.n815 37.5601
R1029 B.n815 B.n15 37.5601
R1030 B.n809 B.n15 37.5601
R1031 B.n809 B.n808 37.5601
R1032 B.n808 B.n807 37.5601
R1033 B.n801 B.n25 37.5601
R1034 B.n801 B.n800 37.5601
R1035 B.n800 B.n799 37.5601
R1036 B.n799 B.n29 37.5601
R1037 B.n793 B.n29 37.5601
R1038 B.n793 B.n792 37.5601
R1039 B.n792 B.n791 37.5601
R1040 B.n791 B.n36 37.5601
R1041 B.n785 B.n36 37.5601
R1042 B.n784 B.n783 37.5601
R1043 B.n783 B.n43 37.5601
R1044 B.n777 B.n43 37.5601
R1045 B.n777 B.n776 37.5601
R1046 B.n776 B.n775 37.5601
R1047 B.n775 B.n50 37.5601
R1048 B.n702 B.t3 35.9031
R1049 B.n807 B.t0 35.9031
R1050 B.n772 B.n771 32.3127
R1051 B.n765 B.n764 32.3127
R1052 B.n436 B.n370 32.3127
R1053 B.n650 B.n649 32.3127
R1054 B.n721 B.t1 27.0655
R1055 B.n817 B.t2 27.0655
R1056 B.n364 B.t9 22.6467
R1057 B.t5 B.n784 22.6467
R1058 B B.n827 18.0485
R1059 B.n671 B.t9 14.9139
R1060 B.n785 B.t5 14.9139
R1061 B.n771 B.n52 10.6151
R1062 B.n113 B.n52 10.6151
R1063 B.n114 B.n113 10.6151
R1064 B.n117 B.n114 10.6151
R1065 B.n118 B.n117 10.6151
R1066 B.n121 B.n118 10.6151
R1067 B.n122 B.n121 10.6151
R1068 B.n125 B.n122 10.6151
R1069 B.n126 B.n125 10.6151
R1070 B.n129 B.n126 10.6151
R1071 B.n130 B.n129 10.6151
R1072 B.n133 B.n130 10.6151
R1073 B.n134 B.n133 10.6151
R1074 B.n137 B.n134 10.6151
R1075 B.n138 B.n137 10.6151
R1076 B.n141 B.n138 10.6151
R1077 B.n142 B.n141 10.6151
R1078 B.n145 B.n142 10.6151
R1079 B.n146 B.n145 10.6151
R1080 B.n149 B.n146 10.6151
R1081 B.n150 B.n149 10.6151
R1082 B.n153 B.n150 10.6151
R1083 B.n154 B.n153 10.6151
R1084 B.n157 B.n154 10.6151
R1085 B.n158 B.n157 10.6151
R1086 B.n161 B.n158 10.6151
R1087 B.n162 B.n161 10.6151
R1088 B.n165 B.n162 10.6151
R1089 B.n166 B.n165 10.6151
R1090 B.n169 B.n166 10.6151
R1091 B.n170 B.n169 10.6151
R1092 B.n173 B.n170 10.6151
R1093 B.n174 B.n173 10.6151
R1094 B.n177 B.n174 10.6151
R1095 B.n178 B.n177 10.6151
R1096 B.n181 B.n178 10.6151
R1097 B.n182 B.n181 10.6151
R1098 B.n185 B.n182 10.6151
R1099 B.n186 B.n185 10.6151
R1100 B.n189 B.n186 10.6151
R1101 B.n190 B.n189 10.6151
R1102 B.n193 B.n190 10.6151
R1103 B.n194 B.n193 10.6151
R1104 B.n197 B.n194 10.6151
R1105 B.n198 B.n197 10.6151
R1106 B.n201 B.n198 10.6151
R1107 B.n202 B.n201 10.6151
R1108 B.n205 B.n202 10.6151
R1109 B.n210 B.n207 10.6151
R1110 B.n211 B.n210 10.6151
R1111 B.n214 B.n211 10.6151
R1112 B.n215 B.n214 10.6151
R1113 B.n218 B.n215 10.6151
R1114 B.n219 B.n218 10.6151
R1115 B.n222 B.n219 10.6151
R1116 B.n223 B.n222 10.6151
R1117 B.n226 B.n223 10.6151
R1118 B.n231 B.n228 10.6151
R1119 B.n232 B.n231 10.6151
R1120 B.n235 B.n232 10.6151
R1121 B.n236 B.n235 10.6151
R1122 B.n239 B.n236 10.6151
R1123 B.n240 B.n239 10.6151
R1124 B.n243 B.n240 10.6151
R1125 B.n244 B.n243 10.6151
R1126 B.n247 B.n244 10.6151
R1127 B.n248 B.n247 10.6151
R1128 B.n251 B.n248 10.6151
R1129 B.n252 B.n251 10.6151
R1130 B.n255 B.n252 10.6151
R1131 B.n256 B.n255 10.6151
R1132 B.n259 B.n256 10.6151
R1133 B.n260 B.n259 10.6151
R1134 B.n263 B.n260 10.6151
R1135 B.n264 B.n263 10.6151
R1136 B.n267 B.n264 10.6151
R1137 B.n268 B.n267 10.6151
R1138 B.n271 B.n268 10.6151
R1139 B.n272 B.n271 10.6151
R1140 B.n275 B.n272 10.6151
R1141 B.n276 B.n275 10.6151
R1142 B.n279 B.n276 10.6151
R1143 B.n280 B.n279 10.6151
R1144 B.n283 B.n280 10.6151
R1145 B.n284 B.n283 10.6151
R1146 B.n287 B.n284 10.6151
R1147 B.n288 B.n287 10.6151
R1148 B.n291 B.n288 10.6151
R1149 B.n292 B.n291 10.6151
R1150 B.n295 B.n292 10.6151
R1151 B.n296 B.n295 10.6151
R1152 B.n299 B.n296 10.6151
R1153 B.n300 B.n299 10.6151
R1154 B.n303 B.n300 10.6151
R1155 B.n304 B.n303 10.6151
R1156 B.n307 B.n304 10.6151
R1157 B.n308 B.n307 10.6151
R1158 B.n311 B.n308 10.6151
R1159 B.n312 B.n311 10.6151
R1160 B.n315 B.n312 10.6151
R1161 B.n316 B.n315 10.6151
R1162 B.n319 B.n316 10.6151
R1163 B.n321 B.n319 10.6151
R1164 B.n322 B.n321 10.6151
R1165 B.n765 B.n322 10.6151
R1166 B.n655 B.n370 10.6151
R1167 B.n656 B.n655 10.6151
R1168 B.n657 B.n656 10.6151
R1169 B.n657 B.n361 10.6151
R1170 B.n667 B.n361 10.6151
R1171 B.n668 B.n667 10.6151
R1172 B.n669 B.n668 10.6151
R1173 B.n669 B.n354 10.6151
R1174 B.n679 B.n354 10.6151
R1175 B.n680 B.n679 10.6151
R1176 B.n681 B.n680 10.6151
R1177 B.n681 B.n346 10.6151
R1178 B.n691 B.n346 10.6151
R1179 B.n692 B.n691 10.6151
R1180 B.n693 B.n692 10.6151
R1181 B.n693 B.n339 10.6151
R1182 B.n704 B.n339 10.6151
R1183 B.n705 B.n704 10.6151
R1184 B.n706 B.n705 10.6151
R1185 B.n706 B.n330 10.6151
R1186 B.n716 B.n330 10.6151
R1187 B.n717 B.n716 10.6151
R1188 B.n719 B.n717 10.6151
R1189 B.n719 B.n718 10.6151
R1190 B.n718 B.n323 10.6151
R1191 B.n730 B.n323 10.6151
R1192 B.n731 B.n730 10.6151
R1193 B.n732 B.n731 10.6151
R1194 B.n733 B.n732 10.6151
R1195 B.n735 B.n733 10.6151
R1196 B.n736 B.n735 10.6151
R1197 B.n737 B.n736 10.6151
R1198 B.n738 B.n737 10.6151
R1199 B.n740 B.n738 10.6151
R1200 B.n741 B.n740 10.6151
R1201 B.n742 B.n741 10.6151
R1202 B.n743 B.n742 10.6151
R1203 B.n745 B.n743 10.6151
R1204 B.n746 B.n745 10.6151
R1205 B.n747 B.n746 10.6151
R1206 B.n748 B.n747 10.6151
R1207 B.n750 B.n748 10.6151
R1208 B.n751 B.n750 10.6151
R1209 B.n752 B.n751 10.6151
R1210 B.n753 B.n752 10.6151
R1211 B.n755 B.n753 10.6151
R1212 B.n756 B.n755 10.6151
R1213 B.n757 B.n756 10.6151
R1214 B.n758 B.n757 10.6151
R1215 B.n760 B.n758 10.6151
R1216 B.n761 B.n760 10.6151
R1217 B.n762 B.n761 10.6151
R1218 B.n763 B.n762 10.6151
R1219 B.n764 B.n763 10.6151
R1220 B.n649 B.n374 10.6151
R1221 B.n644 B.n374 10.6151
R1222 B.n644 B.n643 10.6151
R1223 B.n643 B.n642 10.6151
R1224 B.n642 B.n639 10.6151
R1225 B.n639 B.n638 10.6151
R1226 B.n638 B.n635 10.6151
R1227 B.n635 B.n634 10.6151
R1228 B.n634 B.n631 10.6151
R1229 B.n631 B.n630 10.6151
R1230 B.n630 B.n627 10.6151
R1231 B.n627 B.n626 10.6151
R1232 B.n626 B.n623 10.6151
R1233 B.n623 B.n622 10.6151
R1234 B.n622 B.n619 10.6151
R1235 B.n619 B.n618 10.6151
R1236 B.n618 B.n615 10.6151
R1237 B.n615 B.n614 10.6151
R1238 B.n614 B.n611 10.6151
R1239 B.n611 B.n610 10.6151
R1240 B.n610 B.n607 10.6151
R1241 B.n607 B.n606 10.6151
R1242 B.n606 B.n603 10.6151
R1243 B.n603 B.n602 10.6151
R1244 B.n602 B.n599 10.6151
R1245 B.n599 B.n598 10.6151
R1246 B.n598 B.n595 10.6151
R1247 B.n595 B.n594 10.6151
R1248 B.n594 B.n591 10.6151
R1249 B.n591 B.n590 10.6151
R1250 B.n590 B.n587 10.6151
R1251 B.n587 B.n586 10.6151
R1252 B.n586 B.n583 10.6151
R1253 B.n583 B.n582 10.6151
R1254 B.n582 B.n579 10.6151
R1255 B.n579 B.n578 10.6151
R1256 B.n578 B.n575 10.6151
R1257 B.n575 B.n574 10.6151
R1258 B.n574 B.n571 10.6151
R1259 B.n571 B.n570 10.6151
R1260 B.n570 B.n567 10.6151
R1261 B.n567 B.n566 10.6151
R1262 B.n566 B.n563 10.6151
R1263 B.n563 B.n562 10.6151
R1264 B.n562 B.n559 10.6151
R1265 B.n559 B.n558 10.6151
R1266 B.n558 B.n555 10.6151
R1267 B.n555 B.n554 10.6151
R1268 B.n551 B.n550 10.6151
R1269 B.n550 B.n547 10.6151
R1270 B.n547 B.n546 10.6151
R1271 B.n546 B.n543 10.6151
R1272 B.n543 B.n542 10.6151
R1273 B.n542 B.n539 10.6151
R1274 B.n539 B.n538 10.6151
R1275 B.n538 B.n535 10.6151
R1276 B.n535 B.n534 10.6151
R1277 B.n531 B.n530 10.6151
R1278 B.n530 B.n527 10.6151
R1279 B.n527 B.n526 10.6151
R1280 B.n526 B.n523 10.6151
R1281 B.n523 B.n522 10.6151
R1282 B.n522 B.n519 10.6151
R1283 B.n519 B.n518 10.6151
R1284 B.n518 B.n515 10.6151
R1285 B.n515 B.n514 10.6151
R1286 B.n514 B.n511 10.6151
R1287 B.n511 B.n510 10.6151
R1288 B.n510 B.n507 10.6151
R1289 B.n507 B.n506 10.6151
R1290 B.n506 B.n503 10.6151
R1291 B.n503 B.n502 10.6151
R1292 B.n502 B.n499 10.6151
R1293 B.n499 B.n498 10.6151
R1294 B.n498 B.n495 10.6151
R1295 B.n495 B.n494 10.6151
R1296 B.n494 B.n491 10.6151
R1297 B.n491 B.n490 10.6151
R1298 B.n490 B.n487 10.6151
R1299 B.n487 B.n486 10.6151
R1300 B.n486 B.n483 10.6151
R1301 B.n483 B.n482 10.6151
R1302 B.n482 B.n479 10.6151
R1303 B.n479 B.n478 10.6151
R1304 B.n478 B.n475 10.6151
R1305 B.n475 B.n474 10.6151
R1306 B.n474 B.n471 10.6151
R1307 B.n471 B.n470 10.6151
R1308 B.n470 B.n467 10.6151
R1309 B.n467 B.n466 10.6151
R1310 B.n466 B.n463 10.6151
R1311 B.n463 B.n462 10.6151
R1312 B.n462 B.n459 10.6151
R1313 B.n459 B.n458 10.6151
R1314 B.n458 B.n455 10.6151
R1315 B.n455 B.n454 10.6151
R1316 B.n454 B.n451 10.6151
R1317 B.n451 B.n450 10.6151
R1318 B.n450 B.n447 10.6151
R1319 B.n447 B.n446 10.6151
R1320 B.n446 B.n443 10.6151
R1321 B.n443 B.n442 10.6151
R1322 B.n442 B.n439 10.6151
R1323 B.n439 B.n438 10.6151
R1324 B.n438 B.n436 10.6151
R1325 B.n651 B.n650 10.6151
R1326 B.n651 B.n366 10.6151
R1327 B.n661 B.n366 10.6151
R1328 B.n662 B.n661 10.6151
R1329 B.n663 B.n662 10.6151
R1330 B.n663 B.n358 10.6151
R1331 B.n673 B.n358 10.6151
R1332 B.n674 B.n673 10.6151
R1333 B.n675 B.n674 10.6151
R1334 B.n675 B.n350 10.6151
R1335 B.n685 B.n350 10.6151
R1336 B.n686 B.n685 10.6151
R1337 B.n687 B.n686 10.6151
R1338 B.n687 B.n342 10.6151
R1339 B.n698 B.n342 10.6151
R1340 B.n699 B.n698 10.6151
R1341 B.n700 B.n699 10.6151
R1342 B.n700 B.n335 10.6151
R1343 B.n710 B.n335 10.6151
R1344 B.n711 B.n710 10.6151
R1345 B.n712 B.n711 10.6151
R1346 B.n712 B.n327 10.6151
R1347 B.n723 B.n327 10.6151
R1348 B.n724 B.n723 10.6151
R1349 B.n725 B.n724 10.6151
R1350 B.n725 B.n0 10.6151
R1351 B.n821 B.n1 10.6151
R1352 B.n821 B.n820 10.6151
R1353 B.n820 B.n819 10.6151
R1354 B.n819 B.n10 10.6151
R1355 B.n813 B.n10 10.6151
R1356 B.n813 B.n812 10.6151
R1357 B.n812 B.n811 10.6151
R1358 B.n811 B.n17 10.6151
R1359 B.n805 B.n17 10.6151
R1360 B.n805 B.n804 10.6151
R1361 B.n804 B.n803 10.6151
R1362 B.n803 B.n23 10.6151
R1363 B.n797 B.n23 10.6151
R1364 B.n797 B.n796 10.6151
R1365 B.n796 B.n795 10.6151
R1366 B.n795 B.n31 10.6151
R1367 B.n789 B.n31 10.6151
R1368 B.n789 B.n788 10.6151
R1369 B.n788 B.n787 10.6151
R1370 B.n787 B.n38 10.6151
R1371 B.n781 B.n38 10.6151
R1372 B.n781 B.n780 10.6151
R1373 B.n780 B.n779 10.6151
R1374 B.n779 B.n45 10.6151
R1375 B.n773 B.n45 10.6151
R1376 B.n773 B.n772 10.6151
R1377 B.n333 B.t1 10.4951
R1378 B.t2 B.n816 10.4951
R1379 B.n206 B.n205 9.36635
R1380 B.n228 B.n227 9.36635
R1381 B.n554 B.n432 9.36635
R1382 B.n531 B.n435 9.36635
R1383 B.n827 B.n0 2.81026
R1384 B.n827 B.n1 2.81026
R1385 B.n695 B.t3 1.65754
R1386 B.n25 B.t0 1.65754
R1387 B.n207 B.n206 1.24928
R1388 B.n227 B.n226 1.24928
R1389 B.n551 B.n432 1.24928
R1390 B.n534 B.n435 1.24928
R1391 VP.n3 VP.t2 233.428
R1392 VP.n3 VP.t3 232.999
R1393 VP.n5 VP.t0 197.108
R1394 VP.n13 VP.t1 197.108
R1395 VP.n5 VP.n4 182.722
R1396 VP.n14 VP.n13 182.722
R1397 VP.n12 VP.n0 161.3
R1398 VP.n11 VP.n10 161.3
R1399 VP.n9 VP.n1 161.3
R1400 VP.n8 VP.n7 161.3
R1401 VP.n6 VP.n2 161.3
R1402 VP.n4 VP.n3 55.0913
R1403 VP.n7 VP.n1 40.4106
R1404 VP.n11 VP.n1 40.4106
R1405 VP.n7 VP.n6 24.3439
R1406 VP.n12 VP.n11 24.3439
R1407 VP.n6 VP.n5 2.92171
R1408 VP.n13 VP.n12 2.92171
R1409 VP.n4 VP.n2 0.189894
R1410 VP.n8 VP.n2 0.189894
R1411 VP.n9 VP.n8 0.189894
R1412 VP.n10 VP.n9 0.189894
R1413 VP.n10 VP.n0 0.189894
R1414 VP.n14 VP.n0 0.189894
R1415 VP VP.n14 0.0516364
R1416 VDD1 VDD1.n1 103.263
R1417 VDD1 VDD1.n0 60.9791
R1418 VDD1.n0 VDD1.t1 1.35296
R1419 VDD1.n0 VDD1.t0 1.35296
R1420 VDD1.n1 VDD1.t3 1.35296
R1421 VDD1.n1 VDD1.t2 1.35296
R1422 VTAIL.n650 VTAIL.n574 289.615
R1423 VTAIL.n76 VTAIL.n0 289.615
R1424 VTAIL.n158 VTAIL.n82 289.615
R1425 VTAIL.n240 VTAIL.n164 289.615
R1426 VTAIL.n568 VTAIL.n492 289.615
R1427 VTAIL.n486 VTAIL.n410 289.615
R1428 VTAIL.n404 VTAIL.n328 289.615
R1429 VTAIL.n322 VTAIL.n246 289.615
R1430 VTAIL.n601 VTAIL.n600 185
R1431 VTAIL.n598 VTAIL.n597 185
R1432 VTAIL.n607 VTAIL.n606 185
R1433 VTAIL.n609 VTAIL.n608 185
R1434 VTAIL.n594 VTAIL.n593 185
R1435 VTAIL.n615 VTAIL.n614 185
R1436 VTAIL.n617 VTAIL.n616 185
R1437 VTAIL.n590 VTAIL.n589 185
R1438 VTAIL.n623 VTAIL.n622 185
R1439 VTAIL.n625 VTAIL.n624 185
R1440 VTAIL.n586 VTAIL.n585 185
R1441 VTAIL.n631 VTAIL.n630 185
R1442 VTAIL.n633 VTAIL.n632 185
R1443 VTAIL.n582 VTAIL.n581 185
R1444 VTAIL.n639 VTAIL.n638 185
R1445 VTAIL.n642 VTAIL.n641 185
R1446 VTAIL.n640 VTAIL.n578 185
R1447 VTAIL.n647 VTAIL.n577 185
R1448 VTAIL.n649 VTAIL.n648 185
R1449 VTAIL.n651 VTAIL.n650 185
R1450 VTAIL.n27 VTAIL.n26 185
R1451 VTAIL.n24 VTAIL.n23 185
R1452 VTAIL.n33 VTAIL.n32 185
R1453 VTAIL.n35 VTAIL.n34 185
R1454 VTAIL.n20 VTAIL.n19 185
R1455 VTAIL.n41 VTAIL.n40 185
R1456 VTAIL.n43 VTAIL.n42 185
R1457 VTAIL.n16 VTAIL.n15 185
R1458 VTAIL.n49 VTAIL.n48 185
R1459 VTAIL.n51 VTAIL.n50 185
R1460 VTAIL.n12 VTAIL.n11 185
R1461 VTAIL.n57 VTAIL.n56 185
R1462 VTAIL.n59 VTAIL.n58 185
R1463 VTAIL.n8 VTAIL.n7 185
R1464 VTAIL.n65 VTAIL.n64 185
R1465 VTAIL.n68 VTAIL.n67 185
R1466 VTAIL.n66 VTAIL.n4 185
R1467 VTAIL.n73 VTAIL.n3 185
R1468 VTAIL.n75 VTAIL.n74 185
R1469 VTAIL.n77 VTAIL.n76 185
R1470 VTAIL.n109 VTAIL.n108 185
R1471 VTAIL.n106 VTAIL.n105 185
R1472 VTAIL.n115 VTAIL.n114 185
R1473 VTAIL.n117 VTAIL.n116 185
R1474 VTAIL.n102 VTAIL.n101 185
R1475 VTAIL.n123 VTAIL.n122 185
R1476 VTAIL.n125 VTAIL.n124 185
R1477 VTAIL.n98 VTAIL.n97 185
R1478 VTAIL.n131 VTAIL.n130 185
R1479 VTAIL.n133 VTAIL.n132 185
R1480 VTAIL.n94 VTAIL.n93 185
R1481 VTAIL.n139 VTAIL.n138 185
R1482 VTAIL.n141 VTAIL.n140 185
R1483 VTAIL.n90 VTAIL.n89 185
R1484 VTAIL.n147 VTAIL.n146 185
R1485 VTAIL.n150 VTAIL.n149 185
R1486 VTAIL.n148 VTAIL.n86 185
R1487 VTAIL.n155 VTAIL.n85 185
R1488 VTAIL.n157 VTAIL.n156 185
R1489 VTAIL.n159 VTAIL.n158 185
R1490 VTAIL.n191 VTAIL.n190 185
R1491 VTAIL.n188 VTAIL.n187 185
R1492 VTAIL.n197 VTAIL.n196 185
R1493 VTAIL.n199 VTAIL.n198 185
R1494 VTAIL.n184 VTAIL.n183 185
R1495 VTAIL.n205 VTAIL.n204 185
R1496 VTAIL.n207 VTAIL.n206 185
R1497 VTAIL.n180 VTAIL.n179 185
R1498 VTAIL.n213 VTAIL.n212 185
R1499 VTAIL.n215 VTAIL.n214 185
R1500 VTAIL.n176 VTAIL.n175 185
R1501 VTAIL.n221 VTAIL.n220 185
R1502 VTAIL.n223 VTAIL.n222 185
R1503 VTAIL.n172 VTAIL.n171 185
R1504 VTAIL.n229 VTAIL.n228 185
R1505 VTAIL.n232 VTAIL.n231 185
R1506 VTAIL.n230 VTAIL.n168 185
R1507 VTAIL.n237 VTAIL.n167 185
R1508 VTAIL.n239 VTAIL.n238 185
R1509 VTAIL.n241 VTAIL.n240 185
R1510 VTAIL.n569 VTAIL.n568 185
R1511 VTAIL.n567 VTAIL.n566 185
R1512 VTAIL.n565 VTAIL.n495 185
R1513 VTAIL.n499 VTAIL.n496 185
R1514 VTAIL.n560 VTAIL.n559 185
R1515 VTAIL.n558 VTAIL.n557 185
R1516 VTAIL.n501 VTAIL.n500 185
R1517 VTAIL.n552 VTAIL.n551 185
R1518 VTAIL.n550 VTAIL.n549 185
R1519 VTAIL.n505 VTAIL.n504 185
R1520 VTAIL.n544 VTAIL.n543 185
R1521 VTAIL.n542 VTAIL.n541 185
R1522 VTAIL.n509 VTAIL.n508 185
R1523 VTAIL.n536 VTAIL.n535 185
R1524 VTAIL.n534 VTAIL.n533 185
R1525 VTAIL.n513 VTAIL.n512 185
R1526 VTAIL.n528 VTAIL.n527 185
R1527 VTAIL.n526 VTAIL.n525 185
R1528 VTAIL.n517 VTAIL.n516 185
R1529 VTAIL.n520 VTAIL.n519 185
R1530 VTAIL.n487 VTAIL.n486 185
R1531 VTAIL.n485 VTAIL.n484 185
R1532 VTAIL.n483 VTAIL.n413 185
R1533 VTAIL.n417 VTAIL.n414 185
R1534 VTAIL.n478 VTAIL.n477 185
R1535 VTAIL.n476 VTAIL.n475 185
R1536 VTAIL.n419 VTAIL.n418 185
R1537 VTAIL.n470 VTAIL.n469 185
R1538 VTAIL.n468 VTAIL.n467 185
R1539 VTAIL.n423 VTAIL.n422 185
R1540 VTAIL.n462 VTAIL.n461 185
R1541 VTAIL.n460 VTAIL.n459 185
R1542 VTAIL.n427 VTAIL.n426 185
R1543 VTAIL.n454 VTAIL.n453 185
R1544 VTAIL.n452 VTAIL.n451 185
R1545 VTAIL.n431 VTAIL.n430 185
R1546 VTAIL.n446 VTAIL.n445 185
R1547 VTAIL.n444 VTAIL.n443 185
R1548 VTAIL.n435 VTAIL.n434 185
R1549 VTAIL.n438 VTAIL.n437 185
R1550 VTAIL.n405 VTAIL.n404 185
R1551 VTAIL.n403 VTAIL.n402 185
R1552 VTAIL.n401 VTAIL.n331 185
R1553 VTAIL.n335 VTAIL.n332 185
R1554 VTAIL.n396 VTAIL.n395 185
R1555 VTAIL.n394 VTAIL.n393 185
R1556 VTAIL.n337 VTAIL.n336 185
R1557 VTAIL.n388 VTAIL.n387 185
R1558 VTAIL.n386 VTAIL.n385 185
R1559 VTAIL.n341 VTAIL.n340 185
R1560 VTAIL.n380 VTAIL.n379 185
R1561 VTAIL.n378 VTAIL.n377 185
R1562 VTAIL.n345 VTAIL.n344 185
R1563 VTAIL.n372 VTAIL.n371 185
R1564 VTAIL.n370 VTAIL.n369 185
R1565 VTAIL.n349 VTAIL.n348 185
R1566 VTAIL.n364 VTAIL.n363 185
R1567 VTAIL.n362 VTAIL.n361 185
R1568 VTAIL.n353 VTAIL.n352 185
R1569 VTAIL.n356 VTAIL.n355 185
R1570 VTAIL.n323 VTAIL.n322 185
R1571 VTAIL.n321 VTAIL.n320 185
R1572 VTAIL.n319 VTAIL.n249 185
R1573 VTAIL.n253 VTAIL.n250 185
R1574 VTAIL.n314 VTAIL.n313 185
R1575 VTAIL.n312 VTAIL.n311 185
R1576 VTAIL.n255 VTAIL.n254 185
R1577 VTAIL.n306 VTAIL.n305 185
R1578 VTAIL.n304 VTAIL.n303 185
R1579 VTAIL.n259 VTAIL.n258 185
R1580 VTAIL.n298 VTAIL.n297 185
R1581 VTAIL.n296 VTAIL.n295 185
R1582 VTAIL.n263 VTAIL.n262 185
R1583 VTAIL.n290 VTAIL.n289 185
R1584 VTAIL.n288 VTAIL.n287 185
R1585 VTAIL.n267 VTAIL.n266 185
R1586 VTAIL.n282 VTAIL.n281 185
R1587 VTAIL.n280 VTAIL.n279 185
R1588 VTAIL.n271 VTAIL.n270 185
R1589 VTAIL.n274 VTAIL.n273 185
R1590 VTAIL.t4 VTAIL.n518 147.659
R1591 VTAIL.t5 VTAIL.n436 147.659
R1592 VTAIL.t3 VTAIL.n354 147.659
R1593 VTAIL.t2 VTAIL.n272 147.659
R1594 VTAIL.t0 VTAIL.n599 147.659
R1595 VTAIL.t1 VTAIL.n25 147.659
R1596 VTAIL.t6 VTAIL.n107 147.659
R1597 VTAIL.t7 VTAIL.n189 147.659
R1598 VTAIL.n600 VTAIL.n597 104.615
R1599 VTAIL.n607 VTAIL.n597 104.615
R1600 VTAIL.n608 VTAIL.n607 104.615
R1601 VTAIL.n608 VTAIL.n593 104.615
R1602 VTAIL.n615 VTAIL.n593 104.615
R1603 VTAIL.n616 VTAIL.n615 104.615
R1604 VTAIL.n616 VTAIL.n589 104.615
R1605 VTAIL.n623 VTAIL.n589 104.615
R1606 VTAIL.n624 VTAIL.n623 104.615
R1607 VTAIL.n624 VTAIL.n585 104.615
R1608 VTAIL.n631 VTAIL.n585 104.615
R1609 VTAIL.n632 VTAIL.n631 104.615
R1610 VTAIL.n632 VTAIL.n581 104.615
R1611 VTAIL.n639 VTAIL.n581 104.615
R1612 VTAIL.n641 VTAIL.n639 104.615
R1613 VTAIL.n641 VTAIL.n640 104.615
R1614 VTAIL.n640 VTAIL.n577 104.615
R1615 VTAIL.n649 VTAIL.n577 104.615
R1616 VTAIL.n650 VTAIL.n649 104.615
R1617 VTAIL.n26 VTAIL.n23 104.615
R1618 VTAIL.n33 VTAIL.n23 104.615
R1619 VTAIL.n34 VTAIL.n33 104.615
R1620 VTAIL.n34 VTAIL.n19 104.615
R1621 VTAIL.n41 VTAIL.n19 104.615
R1622 VTAIL.n42 VTAIL.n41 104.615
R1623 VTAIL.n42 VTAIL.n15 104.615
R1624 VTAIL.n49 VTAIL.n15 104.615
R1625 VTAIL.n50 VTAIL.n49 104.615
R1626 VTAIL.n50 VTAIL.n11 104.615
R1627 VTAIL.n57 VTAIL.n11 104.615
R1628 VTAIL.n58 VTAIL.n57 104.615
R1629 VTAIL.n58 VTAIL.n7 104.615
R1630 VTAIL.n65 VTAIL.n7 104.615
R1631 VTAIL.n67 VTAIL.n65 104.615
R1632 VTAIL.n67 VTAIL.n66 104.615
R1633 VTAIL.n66 VTAIL.n3 104.615
R1634 VTAIL.n75 VTAIL.n3 104.615
R1635 VTAIL.n76 VTAIL.n75 104.615
R1636 VTAIL.n108 VTAIL.n105 104.615
R1637 VTAIL.n115 VTAIL.n105 104.615
R1638 VTAIL.n116 VTAIL.n115 104.615
R1639 VTAIL.n116 VTAIL.n101 104.615
R1640 VTAIL.n123 VTAIL.n101 104.615
R1641 VTAIL.n124 VTAIL.n123 104.615
R1642 VTAIL.n124 VTAIL.n97 104.615
R1643 VTAIL.n131 VTAIL.n97 104.615
R1644 VTAIL.n132 VTAIL.n131 104.615
R1645 VTAIL.n132 VTAIL.n93 104.615
R1646 VTAIL.n139 VTAIL.n93 104.615
R1647 VTAIL.n140 VTAIL.n139 104.615
R1648 VTAIL.n140 VTAIL.n89 104.615
R1649 VTAIL.n147 VTAIL.n89 104.615
R1650 VTAIL.n149 VTAIL.n147 104.615
R1651 VTAIL.n149 VTAIL.n148 104.615
R1652 VTAIL.n148 VTAIL.n85 104.615
R1653 VTAIL.n157 VTAIL.n85 104.615
R1654 VTAIL.n158 VTAIL.n157 104.615
R1655 VTAIL.n190 VTAIL.n187 104.615
R1656 VTAIL.n197 VTAIL.n187 104.615
R1657 VTAIL.n198 VTAIL.n197 104.615
R1658 VTAIL.n198 VTAIL.n183 104.615
R1659 VTAIL.n205 VTAIL.n183 104.615
R1660 VTAIL.n206 VTAIL.n205 104.615
R1661 VTAIL.n206 VTAIL.n179 104.615
R1662 VTAIL.n213 VTAIL.n179 104.615
R1663 VTAIL.n214 VTAIL.n213 104.615
R1664 VTAIL.n214 VTAIL.n175 104.615
R1665 VTAIL.n221 VTAIL.n175 104.615
R1666 VTAIL.n222 VTAIL.n221 104.615
R1667 VTAIL.n222 VTAIL.n171 104.615
R1668 VTAIL.n229 VTAIL.n171 104.615
R1669 VTAIL.n231 VTAIL.n229 104.615
R1670 VTAIL.n231 VTAIL.n230 104.615
R1671 VTAIL.n230 VTAIL.n167 104.615
R1672 VTAIL.n239 VTAIL.n167 104.615
R1673 VTAIL.n240 VTAIL.n239 104.615
R1674 VTAIL.n568 VTAIL.n567 104.615
R1675 VTAIL.n567 VTAIL.n495 104.615
R1676 VTAIL.n499 VTAIL.n495 104.615
R1677 VTAIL.n559 VTAIL.n499 104.615
R1678 VTAIL.n559 VTAIL.n558 104.615
R1679 VTAIL.n558 VTAIL.n500 104.615
R1680 VTAIL.n551 VTAIL.n500 104.615
R1681 VTAIL.n551 VTAIL.n550 104.615
R1682 VTAIL.n550 VTAIL.n504 104.615
R1683 VTAIL.n543 VTAIL.n504 104.615
R1684 VTAIL.n543 VTAIL.n542 104.615
R1685 VTAIL.n542 VTAIL.n508 104.615
R1686 VTAIL.n535 VTAIL.n508 104.615
R1687 VTAIL.n535 VTAIL.n534 104.615
R1688 VTAIL.n534 VTAIL.n512 104.615
R1689 VTAIL.n527 VTAIL.n512 104.615
R1690 VTAIL.n527 VTAIL.n526 104.615
R1691 VTAIL.n526 VTAIL.n516 104.615
R1692 VTAIL.n519 VTAIL.n516 104.615
R1693 VTAIL.n486 VTAIL.n485 104.615
R1694 VTAIL.n485 VTAIL.n413 104.615
R1695 VTAIL.n417 VTAIL.n413 104.615
R1696 VTAIL.n477 VTAIL.n417 104.615
R1697 VTAIL.n477 VTAIL.n476 104.615
R1698 VTAIL.n476 VTAIL.n418 104.615
R1699 VTAIL.n469 VTAIL.n418 104.615
R1700 VTAIL.n469 VTAIL.n468 104.615
R1701 VTAIL.n468 VTAIL.n422 104.615
R1702 VTAIL.n461 VTAIL.n422 104.615
R1703 VTAIL.n461 VTAIL.n460 104.615
R1704 VTAIL.n460 VTAIL.n426 104.615
R1705 VTAIL.n453 VTAIL.n426 104.615
R1706 VTAIL.n453 VTAIL.n452 104.615
R1707 VTAIL.n452 VTAIL.n430 104.615
R1708 VTAIL.n445 VTAIL.n430 104.615
R1709 VTAIL.n445 VTAIL.n444 104.615
R1710 VTAIL.n444 VTAIL.n434 104.615
R1711 VTAIL.n437 VTAIL.n434 104.615
R1712 VTAIL.n404 VTAIL.n403 104.615
R1713 VTAIL.n403 VTAIL.n331 104.615
R1714 VTAIL.n335 VTAIL.n331 104.615
R1715 VTAIL.n395 VTAIL.n335 104.615
R1716 VTAIL.n395 VTAIL.n394 104.615
R1717 VTAIL.n394 VTAIL.n336 104.615
R1718 VTAIL.n387 VTAIL.n336 104.615
R1719 VTAIL.n387 VTAIL.n386 104.615
R1720 VTAIL.n386 VTAIL.n340 104.615
R1721 VTAIL.n379 VTAIL.n340 104.615
R1722 VTAIL.n379 VTAIL.n378 104.615
R1723 VTAIL.n378 VTAIL.n344 104.615
R1724 VTAIL.n371 VTAIL.n344 104.615
R1725 VTAIL.n371 VTAIL.n370 104.615
R1726 VTAIL.n370 VTAIL.n348 104.615
R1727 VTAIL.n363 VTAIL.n348 104.615
R1728 VTAIL.n363 VTAIL.n362 104.615
R1729 VTAIL.n362 VTAIL.n352 104.615
R1730 VTAIL.n355 VTAIL.n352 104.615
R1731 VTAIL.n322 VTAIL.n321 104.615
R1732 VTAIL.n321 VTAIL.n249 104.615
R1733 VTAIL.n253 VTAIL.n249 104.615
R1734 VTAIL.n313 VTAIL.n253 104.615
R1735 VTAIL.n313 VTAIL.n312 104.615
R1736 VTAIL.n312 VTAIL.n254 104.615
R1737 VTAIL.n305 VTAIL.n254 104.615
R1738 VTAIL.n305 VTAIL.n304 104.615
R1739 VTAIL.n304 VTAIL.n258 104.615
R1740 VTAIL.n297 VTAIL.n258 104.615
R1741 VTAIL.n297 VTAIL.n296 104.615
R1742 VTAIL.n296 VTAIL.n262 104.615
R1743 VTAIL.n289 VTAIL.n262 104.615
R1744 VTAIL.n289 VTAIL.n288 104.615
R1745 VTAIL.n288 VTAIL.n266 104.615
R1746 VTAIL.n281 VTAIL.n266 104.615
R1747 VTAIL.n281 VTAIL.n280 104.615
R1748 VTAIL.n280 VTAIL.n270 104.615
R1749 VTAIL.n273 VTAIL.n270 104.615
R1750 VTAIL.n600 VTAIL.t0 52.3082
R1751 VTAIL.n26 VTAIL.t1 52.3082
R1752 VTAIL.n108 VTAIL.t6 52.3082
R1753 VTAIL.n190 VTAIL.t7 52.3082
R1754 VTAIL.n519 VTAIL.t4 52.3082
R1755 VTAIL.n437 VTAIL.t5 52.3082
R1756 VTAIL.n355 VTAIL.t3 52.3082
R1757 VTAIL.n273 VTAIL.t2 52.3082
R1758 VTAIL.n655 VTAIL.n654 32.1853
R1759 VTAIL.n81 VTAIL.n80 32.1853
R1760 VTAIL.n163 VTAIL.n162 32.1853
R1761 VTAIL.n245 VTAIL.n244 32.1853
R1762 VTAIL.n573 VTAIL.n572 32.1853
R1763 VTAIL.n491 VTAIL.n490 32.1853
R1764 VTAIL.n409 VTAIL.n408 32.1853
R1765 VTAIL.n327 VTAIL.n326 32.1853
R1766 VTAIL.n655 VTAIL.n573 26.8152
R1767 VTAIL.n327 VTAIL.n245 26.8152
R1768 VTAIL.n601 VTAIL.n599 15.6677
R1769 VTAIL.n27 VTAIL.n25 15.6677
R1770 VTAIL.n109 VTAIL.n107 15.6677
R1771 VTAIL.n191 VTAIL.n189 15.6677
R1772 VTAIL.n520 VTAIL.n518 15.6677
R1773 VTAIL.n438 VTAIL.n436 15.6677
R1774 VTAIL.n356 VTAIL.n354 15.6677
R1775 VTAIL.n274 VTAIL.n272 15.6677
R1776 VTAIL.n648 VTAIL.n647 13.1884
R1777 VTAIL.n74 VTAIL.n73 13.1884
R1778 VTAIL.n156 VTAIL.n155 13.1884
R1779 VTAIL.n238 VTAIL.n237 13.1884
R1780 VTAIL.n566 VTAIL.n565 13.1884
R1781 VTAIL.n484 VTAIL.n483 13.1884
R1782 VTAIL.n402 VTAIL.n401 13.1884
R1783 VTAIL.n320 VTAIL.n319 13.1884
R1784 VTAIL.n602 VTAIL.n598 12.8005
R1785 VTAIL.n646 VTAIL.n578 12.8005
R1786 VTAIL.n651 VTAIL.n576 12.8005
R1787 VTAIL.n28 VTAIL.n24 12.8005
R1788 VTAIL.n72 VTAIL.n4 12.8005
R1789 VTAIL.n77 VTAIL.n2 12.8005
R1790 VTAIL.n110 VTAIL.n106 12.8005
R1791 VTAIL.n154 VTAIL.n86 12.8005
R1792 VTAIL.n159 VTAIL.n84 12.8005
R1793 VTAIL.n192 VTAIL.n188 12.8005
R1794 VTAIL.n236 VTAIL.n168 12.8005
R1795 VTAIL.n241 VTAIL.n166 12.8005
R1796 VTAIL.n569 VTAIL.n494 12.8005
R1797 VTAIL.n564 VTAIL.n496 12.8005
R1798 VTAIL.n521 VTAIL.n517 12.8005
R1799 VTAIL.n487 VTAIL.n412 12.8005
R1800 VTAIL.n482 VTAIL.n414 12.8005
R1801 VTAIL.n439 VTAIL.n435 12.8005
R1802 VTAIL.n405 VTAIL.n330 12.8005
R1803 VTAIL.n400 VTAIL.n332 12.8005
R1804 VTAIL.n357 VTAIL.n353 12.8005
R1805 VTAIL.n323 VTAIL.n248 12.8005
R1806 VTAIL.n318 VTAIL.n250 12.8005
R1807 VTAIL.n275 VTAIL.n271 12.8005
R1808 VTAIL.n606 VTAIL.n605 12.0247
R1809 VTAIL.n643 VTAIL.n642 12.0247
R1810 VTAIL.n652 VTAIL.n574 12.0247
R1811 VTAIL.n32 VTAIL.n31 12.0247
R1812 VTAIL.n69 VTAIL.n68 12.0247
R1813 VTAIL.n78 VTAIL.n0 12.0247
R1814 VTAIL.n114 VTAIL.n113 12.0247
R1815 VTAIL.n151 VTAIL.n150 12.0247
R1816 VTAIL.n160 VTAIL.n82 12.0247
R1817 VTAIL.n196 VTAIL.n195 12.0247
R1818 VTAIL.n233 VTAIL.n232 12.0247
R1819 VTAIL.n242 VTAIL.n164 12.0247
R1820 VTAIL.n570 VTAIL.n492 12.0247
R1821 VTAIL.n561 VTAIL.n560 12.0247
R1822 VTAIL.n525 VTAIL.n524 12.0247
R1823 VTAIL.n488 VTAIL.n410 12.0247
R1824 VTAIL.n479 VTAIL.n478 12.0247
R1825 VTAIL.n443 VTAIL.n442 12.0247
R1826 VTAIL.n406 VTAIL.n328 12.0247
R1827 VTAIL.n397 VTAIL.n396 12.0247
R1828 VTAIL.n361 VTAIL.n360 12.0247
R1829 VTAIL.n324 VTAIL.n246 12.0247
R1830 VTAIL.n315 VTAIL.n314 12.0247
R1831 VTAIL.n279 VTAIL.n278 12.0247
R1832 VTAIL.n609 VTAIL.n596 11.249
R1833 VTAIL.n638 VTAIL.n580 11.249
R1834 VTAIL.n35 VTAIL.n22 11.249
R1835 VTAIL.n64 VTAIL.n6 11.249
R1836 VTAIL.n117 VTAIL.n104 11.249
R1837 VTAIL.n146 VTAIL.n88 11.249
R1838 VTAIL.n199 VTAIL.n186 11.249
R1839 VTAIL.n228 VTAIL.n170 11.249
R1840 VTAIL.n557 VTAIL.n498 11.249
R1841 VTAIL.n528 VTAIL.n515 11.249
R1842 VTAIL.n475 VTAIL.n416 11.249
R1843 VTAIL.n446 VTAIL.n433 11.249
R1844 VTAIL.n393 VTAIL.n334 11.249
R1845 VTAIL.n364 VTAIL.n351 11.249
R1846 VTAIL.n311 VTAIL.n252 11.249
R1847 VTAIL.n282 VTAIL.n269 11.249
R1848 VTAIL.n610 VTAIL.n594 10.4732
R1849 VTAIL.n637 VTAIL.n582 10.4732
R1850 VTAIL.n36 VTAIL.n20 10.4732
R1851 VTAIL.n63 VTAIL.n8 10.4732
R1852 VTAIL.n118 VTAIL.n102 10.4732
R1853 VTAIL.n145 VTAIL.n90 10.4732
R1854 VTAIL.n200 VTAIL.n184 10.4732
R1855 VTAIL.n227 VTAIL.n172 10.4732
R1856 VTAIL.n556 VTAIL.n501 10.4732
R1857 VTAIL.n529 VTAIL.n513 10.4732
R1858 VTAIL.n474 VTAIL.n419 10.4732
R1859 VTAIL.n447 VTAIL.n431 10.4732
R1860 VTAIL.n392 VTAIL.n337 10.4732
R1861 VTAIL.n365 VTAIL.n349 10.4732
R1862 VTAIL.n310 VTAIL.n255 10.4732
R1863 VTAIL.n283 VTAIL.n267 10.4732
R1864 VTAIL.n614 VTAIL.n613 9.69747
R1865 VTAIL.n634 VTAIL.n633 9.69747
R1866 VTAIL.n40 VTAIL.n39 9.69747
R1867 VTAIL.n60 VTAIL.n59 9.69747
R1868 VTAIL.n122 VTAIL.n121 9.69747
R1869 VTAIL.n142 VTAIL.n141 9.69747
R1870 VTAIL.n204 VTAIL.n203 9.69747
R1871 VTAIL.n224 VTAIL.n223 9.69747
R1872 VTAIL.n553 VTAIL.n552 9.69747
R1873 VTAIL.n533 VTAIL.n532 9.69747
R1874 VTAIL.n471 VTAIL.n470 9.69747
R1875 VTAIL.n451 VTAIL.n450 9.69747
R1876 VTAIL.n389 VTAIL.n388 9.69747
R1877 VTAIL.n369 VTAIL.n368 9.69747
R1878 VTAIL.n307 VTAIL.n306 9.69747
R1879 VTAIL.n287 VTAIL.n286 9.69747
R1880 VTAIL.n654 VTAIL.n653 9.45567
R1881 VTAIL.n80 VTAIL.n79 9.45567
R1882 VTAIL.n162 VTAIL.n161 9.45567
R1883 VTAIL.n244 VTAIL.n243 9.45567
R1884 VTAIL.n572 VTAIL.n571 9.45567
R1885 VTAIL.n490 VTAIL.n489 9.45567
R1886 VTAIL.n408 VTAIL.n407 9.45567
R1887 VTAIL.n326 VTAIL.n325 9.45567
R1888 VTAIL.n653 VTAIL.n652 9.3005
R1889 VTAIL.n576 VTAIL.n575 9.3005
R1890 VTAIL.n621 VTAIL.n620 9.3005
R1891 VTAIL.n619 VTAIL.n618 9.3005
R1892 VTAIL.n592 VTAIL.n591 9.3005
R1893 VTAIL.n613 VTAIL.n612 9.3005
R1894 VTAIL.n611 VTAIL.n610 9.3005
R1895 VTAIL.n596 VTAIL.n595 9.3005
R1896 VTAIL.n605 VTAIL.n604 9.3005
R1897 VTAIL.n603 VTAIL.n602 9.3005
R1898 VTAIL.n588 VTAIL.n587 9.3005
R1899 VTAIL.n627 VTAIL.n626 9.3005
R1900 VTAIL.n629 VTAIL.n628 9.3005
R1901 VTAIL.n584 VTAIL.n583 9.3005
R1902 VTAIL.n635 VTAIL.n634 9.3005
R1903 VTAIL.n637 VTAIL.n636 9.3005
R1904 VTAIL.n580 VTAIL.n579 9.3005
R1905 VTAIL.n644 VTAIL.n643 9.3005
R1906 VTAIL.n646 VTAIL.n645 9.3005
R1907 VTAIL.n79 VTAIL.n78 9.3005
R1908 VTAIL.n2 VTAIL.n1 9.3005
R1909 VTAIL.n47 VTAIL.n46 9.3005
R1910 VTAIL.n45 VTAIL.n44 9.3005
R1911 VTAIL.n18 VTAIL.n17 9.3005
R1912 VTAIL.n39 VTAIL.n38 9.3005
R1913 VTAIL.n37 VTAIL.n36 9.3005
R1914 VTAIL.n22 VTAIL.n21 9.3005
R1915 VTAIL.n31 VTAIL.n30 9.3005
R1916 VTAIL.n29 VTAIL.n28 9.3005
R1917 VTAIL.n14 VTAIL.n13 9.3005
R1918 VTAIL.n53 VTAIL.n52 9.3005
R1919 VTAIL.n55 VTAIL.n54 9.3005
R1920 VTAIL.n10 VTAIL.n9 9.3005
R1921 VTAIL.n61 VTAIL.n60 9.3005
R1922 VTAIL.n63 VTAIL.n62 9.3005
R1923 VTAIL.n6 VTAIL.n5 9.3005
R1924 VTAIL.n70 VTAIL.n69 9.3005
R1925 VTAIL.n72 VTAIL.n71 9.3005
R1926 VTAIL.n161 VTAIL.n160 9.3005
R1927 VTAIL.n84 VTAIL.n83 9.3005
R1928 VTAIL.n129 VTAIL.n128 9.3005
R1929 VTAIL.n127 VTAIL.n126 9.3005
R1930 VTAIL.n100 VTAIL.n99 9.3005
R1931 VTAIL.n121 VTAIL.n120 9.3005
R1932 VTAIL.n119 VTAIL.n118 9.3005
R1933 VTAIL.n104 VTAIL.n103 9.3005
R1934 VTAIL.n113 VTAIL.n112 9.3005
R1935 VTAIL.n111 VTAIL.n110 9.3005
R1936 VTAIL.n96 VTAIL.n95 9.3005
R1937 VTAIL.n135 VTAIL.n134 9.3005
R1938 VTAIL.n137 VTAIL.n136 9.3005
R1939 VTAIL.n92 VTAIL.n91 9.3005
R1940 VTAIL.n143 VTAIL.n142 9.3005
R1941 VTAIL.n145 VTAIL.n144 9.3005
R1942 VTAIL.n88 VTAIL.n87 9.3005
R1943 VTAIL.n152 VTAIL.n151 9.3005
R1944 VTAIL.n154 VTAIL.n153 9.3005
R1945 VTAIL.n243 VTAIL.n242 9.3005
R1946 VTAIL.n166 VTAIL.n165 9.3005
R1947 VTAIL.n211 VTAIL.n210 9.3005
R1948 VTAIL.n209 VTAIL.n208 9.3005
R1949 VTAIL.n182 VTAIL.n181 9.3005
R1950 VTAIL.n203 VTAIL.n202 9.3005
R1951 VTAIL.n201 VTAIL.n200 9.3005
R1952 VTAIL.n186 VTAIL.n185 9.3005
R1953 VTAIL.n195 VTAIL.n194 9.3005
R1954 VTAIL.n193 VTAIL.n192 9.3005
R1955 VTAIL.n178 VTAIL.n177 9.3005
R1956 VTAIL.n217 VTAIL.n216 9.3005
R1957 VTAIL.n219 VTAIL.n218 9.3005
R1958 VTAIL.n174 VTAIL.n173 9.3005
R1959 VTAIL.n225 VTAIL.n224 9.3005
R1960 VTAIL.n227 VTAIL.n226 9.3005
R1961 VTAIL.n170 VTAIL.n169 9.3005
R1962 VTAIL.n234 VTAIL.n233 9.3005
R1963 VTAIL.n236 VTAIL.n235 9.3005
R1964 VTAIL.n546 VTAIL.n545 9.3005
R1965 VTAIL.n548 VTAIL.n547 9.3005
R1966 VTAIL.n503 VTAIL.n502 9.3005
R1967 VTAIL.n554 VTAIL.n553 9.3005
R1968 VTAIL.n556 VTAIL.n555 9.3005
R1969 VTAIL.n498 VTAIL.n497 9.3005
R1970 VTAIL.n562 VTAIL.n561 9.3005
R1971 VTAIL.n564 VTAIL.n563 9.3005
R1972 VTAIL.n571 VTAIL.n570 9.3005
R1973 VTAIL.n494 VTAIL.n493 9.3005
R1974 VTAIL.n507 VTAIL.n506 9.3005
R1975 VTAIL.n540 VTAIL.n539 9.3005
R1976 VTAIL.n538 VTAIL.n537 9.3005
R1977 VTAIL.n511 VTAIL.n510 9.3005
R1978 VTAIL.n532 VTAIL.n531 9.3005
R1979 VTAIL.n530 VTAIL.n529 9.3005
R1980 VTAIL.n515 VTAIL.n514 9.3005
R1981 VTAIL.n524 VTAIL.n523 9.3005
R1982 VTAIL.n522 VTAIL.n521 9.3005
R1983 VTAIL.n464 VTAIL.n463 9.3005
R1984 VTAIL.n466 VTAIL.n465 9.3005
R1985 VTAIL.n421 VTAIL.n420 9.3005
R1986 VTAIL.n472 VTAIL.n471 9.3005
R1987 VTAIL.n474 VTAIL.n473 9.3005
R1988 VTAIL.n416 VTAIL.n415 9.3005
R1989 VTAIL.n480 VTAIL.n479 9.3005
R1990 VTAIL.n482 VTAIL.n481 9.3005
R1991 VTAIL.n489 VTAIL.n488 9.3005
R1992 VTAIL.n412 VTAIL.n411 9.3005
R1993 VTAIL.n425 VTAIL.n424 9.3005
R1994 VTAIL.n458 VTAIL.n457 9.3005
R1995 VTAIL.n456 VTAIL.n455 9.3005
R1996 VTAIL.n429 VTAIL.n428 9.3005
R1997 VTAIL.n450 VTAIL.n449 9.3005
R1998 VTAIL.n448 VTAIL.n447 9.3005
R1999 VTAIL.n433 VTAIL.n432 9.3005
R2000 VTAIL.n442 VTAIL.n441 9.3005
R2001 VTAIL.n440 VTAIL.n439 9.3005
R2002 VTAIL.n382 VTAIL.n381 9.3005
R2003 VTAIL.n384 VTAIL.n383 9.3005
R2004 VTAIL.n339 VTAIL.n338 9.3005
R2005 VTAIL.n390 VTAIL.n389 9.3005
R2006 VTAIL.n392 VTAIL.n391 9.3005
R2007 VTAIL.n334 VTAIL.n333 9.3005
R2008 VTAIL.n398 VTAIL.n397 9.3005
R2009 VTAIL.n400 VTAIL.n399 9.3005
R2010 VTAIL.n407 VTAIL.n406 9.3005
R2011 VTAIL.n330 VTAIL.n329 9.3005
R2012 VTAIL.n343 VTAIL.n342 9.3005
R2013 VTAIL.n376 VTAIL.n375 9.3005
R2014 VTAIL.n374 VTAIL.n373 9.3005
R2015 VTAIL.n347 VTAIL.n346 9.3005
R2016 VTAIL.n368 VTAIL.n367 9.3005
R2017 VTAIL.n366 VTAIL.n365 9.3005
R2018 VTAIL.n351 VTAIL.n350 9.3005
R2019 VTAIL.n360 VTAIL.n359 9.3005
R2020 VTAIL.n358 VTAIL.n357 9.3005
R2021 VTAIL.n300 VTAIL.n299 9.3005
R2022 VTAIL.n302 VTAIL.n301 9.3005
R2023 VTAIL.n257 VTAIL.n256 9.3005
R2024 VTAIL.n308 VTAIL.n307 9.3005
R2025 VTAIL.n310 VTAIL.n309 9.3005
R2026 VTAIL.n252 VTAIL.n251 9.3005
R2027 VTAIL.n316 VTAIL.n315 9.3005
R2028 VTAIL.n318 VTAIL.n317 9.3005
R2029 VTAIL.n325 VTAIL.n324 9.3005
R2030 VTAIL.n248 VTAIL.n247 9.3005
R2031 VTAIL.n261 VTAIL.n260 9.3005
R2032 VTAIL.n294 VTAIL.n293 9.3005
R2033 VTAIL.n292 VTAIL.n291 9.3005
R2034 VTAIL.n265 VTAIL.n264 9.3005
R2035 VTAIL.n286 VTAIL.n285 9.3005
R2036 VTAIL.n284 VTAIL.n283 9.3005
R2037 VTAIL.n269 VTAIL.n268 9.3005
R2038 VTAIL.n278 VTAIL.n277 9.3005
R2039 VTAIL.n276 VTAIL.n275 9.3005
R2040 VTAIL.n617 VTAIL.n592 8.92171
R2041 VTAIL.n630 VTAIL.n584 8.92171
R2042 VTAIL.n43 VTAIL.n18 8.92171
R2043 VTAIL.n56 VTAIL.n10 8.92171
R2044 VTAIL.n125 VTAIL.n100 8.92171
R2045 VTAIL.n138 VTAIL.n92 8.92171
R2046 VTAIL.n207 VTAIL.n182 8.92171
R2047 VTAIL.n220 VTAIL.n174 8.92171
R2048 VTAIL.n549 VTAIL.n503 8.92171
R2049 VTAIL.n536 VTAIL.n511 8.92171
R2050 VTAIL.n467 VTAIL.n421 8.92171
R2051 VTAIL.n454 VTAIL.n429 8.92171
R2052 VTAIL.n385 VTAIL.n339 8.92171
R2053 VTAIL.n372 VTAIL.n347 8.92171
R2054 VTAIL.n303 VTAIL.n257 8.92171
R2055 VTAIL.n290 VTAIL.n265 8.92171
R2056 VTAIL.n618 VTAIL.n590 8.14595
R2057 VTAIL.n629 VTAIL.n586 8.14595
R2058 VTAIL.n44 VTAIL.n16 8.14595
R2059 VTAIL.n55 VTAIL.n12 8.14595
R2060 VTAIL.n126 VTAIL.n98 8.14595
R2061 VTAIL.n137 VTAIL.n94 8.14595
R2062 VTAIL.n208 VTAIL.n180 8.14595
R2063 VTAIL.n219 VTAIL.n176 8.14595
R2064 VTAIL.n548 VTAIL.n505 8.14595
R2065 VTAIL.n537 VTAIL.n509 8.14595
R2066 VTAIL.n466 VTAIL.n423 8.14595
R2067 VTAIL.n455 VTAIL.n427 8.14595
R2068 VTAIL.n384 VTAIL.n341 8.14595
R2069 VTAIL.n373 VTAIL.n345 8.14595
R2070 VTAIL.n302 VTAIL.n259 8.14595
R2071 VTAIL.n291 VTAIL.n263 8.14595
R2072 VTAIL.n622 VTAIL.n621 7.3702
R2073 VTAIL.n626 VTAIL.n625 7.3702
R2074 VTAIL.n48 VTAIL.n47 7.3702
R2075 VTAIL.n52 VTAIL.n51 7.3702
R2076 VTAIL.n130 VTAIL.n129 7.3702
R2077 VTAIL.n134 VTAIL.n133 7.3702
R2078 VTAIL.n212 VTAIL.n211 7.3702
R2079 VTAIL.n216 VTAIL.n215 7.3702
R2080 VTAIL.n545 VTAIL.n544 7.3702
R2081 VTAIL.n541 VTAIL.n540 7.3702
R2082 VTAIL.n463 VTAIL.n462 7.3702
R2083 VTAIL.n459 VTAIL.n458 7.3702
R2084 VTAIL.n381 VTAIL.n380 7.3702
R2085 VTAIL.n377 VTAIL.n376 7.3702
R2086 VTAIL.n299 VTAIL.n298 7.3702
R2087 VTAIL.n295 VTAIL.n294 7.3702
R2088 VTAIL.n622 VTAIL.n588 6.59444
R2089 VTAIL.n625 VTAIL.n588 6.59444
R2090 VTAIL.n48 VTAIL.n14 6.59444
R2091 VTAIL.n51 VTAIL.n14 6.59444
R2092 VTAIL.n130 VTAIL.n96 6.59444
R2093 VTAIL.n133 VTAIL.n96 6.59444
R2094 VTAIL.n212 VTAIL.n178 6.59444
R2095 VTAIL.n215 VTAIL.n178 6.59444
R2096 VTAIL.n544 VTAIL.n507 6.59444
R2097 VTAIL.n541 VTAIL.n507 6.59444
R2098 VTAIL.n462 VTAIL.n425 6.59444
R2099 VTAIL.n459 VTAIL.n425 6.59444
R2100 VTAIL.n380 VTAIL.n343 6.59444
R2101 VTAIL.n377 VTAIL.n343 6.59444
R2102 VTAIL.n298 VTAIL.n261 6.59444
R2103 VTAIL.n295 VTAIL.n261 6.59444
R2104 VTAIL.n621 VTAIL.n590 5.81868
R2105 VTAIL.n626 VTAIL.n586 5.81868
R2106 VTAIL.n47 VTAIL.n16 5.81868
R2107 VTAIL.n52 VTAIL.n12 5.81868
R2108 VTAIL.n129 VTAIL.n98 5.81868
R2109 VTAIL.n134 VTAIL.n94 5.81868
R2110 VTAIL.n211 VTAIL.n180 5.81868
R2111 VTAIL.n216 VTAIL.n176 5.81868
R2112 VTAIL.n545 VTAIL.n505 5.81868
R2113 VTAIL.n540 VTAIL.n509 5.81868
R2114 VTAIL.n463 VTAIL.n423 5.81868
R2115 VTAIL.n458 VTAIL.n427 5.81868
R2116 VTAIL.n381 VTAIL.n341 5.81868
R2117 VTAIL.n376 VTAIL.n345 5.81868
R2118 VTAIL.n299 VTAIL.n259 5.81868
R2119 VTAIL.n294 VTAIL.n263 5.81868
R2120 VTAIL.n618 VTAIL.n617 5.04292
R2121 VTAIL.n630 VTAIL.n629 5.04292
R2122 VTAIL.n44 VTAIL.n43 5.04292
R2123 VTAIL.n56 VTAIL.n55 5.04292
R2124 VTAIL.n126 VTAIL.n125 5.04292
R2125 VTAIL.n138 VTAIL.n137 5.04292
R2126 VTAIL.n208 VTAIL.n207 5.04292
R2127 VTAIL.n220 VTAIL.n219 5.04292
R2128 VTAIL.n549 VTAIL.n548 5.04292
R2129 VTAIL.n537 VTAIL.n536 5.04292
R2130 VTAIL.n467 VTAIL.n466 5.04292
R2131 VTAIL.n455 VTAIL.n454 5.04292
R2132 VTAIL.n385 VTAIL.n384 5.04292
R2133 VTAIL.n373 VTAIL.n372 5.04292
R2134 VTAIL.n303 VTAIL.n302 5.04292
R2135 VTAIL.n291 VTAIL.n290 5.04292
R2136 VTAIL.n522 VTAIL.n518 4.38563
R2137 VTAIL.n440 VTAIL.n436 4.38563
R2138 VTAIL.n358 VTAIL.n354 4.38563
R2139 VTAIL.n276 VTAIL.n272 4.38563
R2140 VTAIL.n603 VTAIL.n599 4.38563
R2141 VTAIL.n29 VTAIL.n25 4.38563
R2142 VTAIL.n111 VTAIL.n107 4.38563
R2143 VTAIL.n193 VTAIL.n189 4.38563
R2144 VTAIL.n614 VTAIL.n592 4.26717
R2145 VTAIL.n633 VTAIL.n584 4.26717
R2146 VTAIL.n40 VTAIL.n18 4.26717
R2147 VTAIL.n59 VTAIL.n10 4.26717
R2148 VTAIL.n122 VTAIL.n100 4.26717
R2149 VTAIL.n141 VTAIL.n92 4.26717
R2150 VTAIL.n204 VTAIL.n182 4.26717
R2151 VTAIL.n223 VTAIL.n174 4.26717
R2152 VTAIL.n552 VTAIL.n503 4.26717
R2153 VTAIL.n533 VTAIL.n511 4.26717
R2154 VTAIL.n470 VTAIL.n421 4.26717
R2155 VTAIL.n451 VTAIL.n429 4.26717
R2156 VTAIL.n388 VTAIL.n339 4.26717
R2157 VTAIL.n369 VTAIL.n347 4.26717
R2158 VTAIL.n306 VTAIL.n257 4.26717
R2159 VTAIL.n287 VTAIL.n265 4.26717
R2160 VTAIL.n613 VTAIL.n594 3.49141
R2161 VTAIL.n634 VTAIL.n582 3.49141
R2162 VTAIL.n39 VTAIL.n20 3.49141
R2163 VTAIL.n60 VTAIL.n8 3.49141
R2164 VTAIL.n121 VTAIL.n102 3.49141
R2165 VTAIL.n142 VTAIL.n90 3.49141
R2166 VTAIL.n203 VTAIL.n184 3.49141
R2167 VTAIL.n224 VTAIL.n172 3.49141
R2168 VTAIL.n553 VTAIL.n501 3.49141
R2169 VTAIL.n532 VTAIL.n513 3.49141
R2170 VTAIL.n471 VTAIL.n419 3.49141
R2171 VTAIL.n450 VTAIL.n431 3.49141
R2172 VTAIL.n389 VTAIL.n337 3.49141
R2173 VTAIL.n368 VTAIL.n349 3.49141
R2174 VTAIL.n307 VTAIL.n255 3.49141
R2175 VTAIL.n286 VTAIL.n267 3.49141
R2176 VTAIL.n610 VTAIL.n609 2.71565
R2177 VTAIL.n638 VTAIL.n637 2.71565
R2178 VTAIL.n36 VTAIL.n35 2.71565
R2179 VTAIL.n64 VTAIL.n63 2.71565
R2180 VTAIL.n118 VTAIL.n117 2.71565
R2181 VTAIL.n146 VTAIL.n145 2.71565
R2182 VTAIL.n200 VTAIL.n199 2.71565
R2183 VTAIL.n228 VTAIL.n227 2.71565
R2184 VTAIL.n557 VTAIL.n556 2.71565
R2185 VTAIL.n529 VTAIL.n528 2.71565
R2186 VTAIL.n475 VTAIL.n474 2.71565
R2187 VTAIL.n447 VTAIL.n446 2.71565
R2188 VTAIL.n393 VTAIL.n392 2.71565
R2189 VTAIL.n365 VTAIL.n364 2.71565
R2190 VTAIL.n311 VTAIL.n310 2.71565
R2191 VTAIL.n283 VTAIL.n282 2.71565
R2192 VTAIL.n606 VTAIL.n596 1.93989
R2193 VTAIL.n642 VTAIL.n580 1.93989
R2194 VTAIL.n654 VTAIL.n574 1.93989
R2195 VTAIL.n32 VTAIL.n22 1.93989
R2196 VTAIL.n68 VTAIL.n6 1.93989
R2197 VTAIL.n80 VTAIL.n0 1.93989
R2198 VTAIL.n114 VTAIL.n104 1.93989
R2199 VTAIL.n150 VTAIL.n88 1.93989
R2200 VTAIL.n162 VTAIL.n82 1.93989
R2201 VTAIL.n196 VTAIL.n186 1.93989
R2202 VTAIL.n232 VTAIL.n170 1.93989
R2203 VTAIL.n244 VTAIL.n164 1.93989
R2204 VTAIL.n572 VTAIL.n492 1.93989
R2205 VTAIL.n560 VTAIL.n498 1.93989
R2206 VTAIL.n525 VTAIL.n515 1.93989
R2207 VTAIL.n490 VTAIL.n410 1.93989
R2208 VTAIL.n478 VTAIL.n416 1.93989
R2209 VTAIL.n443 VTAIL.n433 1.93989
R2210 VTAIL.n408 VTAIL.n328 1.93989
R2211 VTAIL.n396 VTAIL.n334 1.93989
R2212 VTAIL.n361 VTAIL.n351 1.93989
R2213 VTAIL.n326 VTAIL.n246 1.93989
R2214 VTAIL.n314 VTAIL.n252 1.93989
R2215 VTAIL.n279 VTAIL.n269 1.93989
R2216 VTAIL.n409 VTAIL.n327 1.82809
R2217 VTAIL.n573 VTAIL.n491 1.82809
R2218 VTAIL.n245 VTAIL.n163 1.82809
R2219 VTAIL.n605 VTAIL.n598 1.16414
R2220 VTAIL.n643 VTAIL.n578 1.16414
R2221 VTAIL.n652 VTAIL.n651 1.16414
R2222 VTAIL.n31 VTAIL.n24 1.16414
R2223 VTAIL.n69 VTAIL.n4 1.16414
R2224 VTAIL.n78 VTAIL.n77 1.16414
R2225 VTAIL.n113 VTAIL.n106 1.16414
R2226 VTAIL.n151 VTAIL.n86 1.16414
R2227 VTAIL.n160 VTAIL.n159 1.16414
R2228 VTAIL.n195 VTAIL.n188 1.16414
R2229 VTAIL.n233 VTAIL.n168 1.16414
R2230 VTAIL.n242 VTAIL.n241 1.16414
R2231 VTAIL.n570 VTAIL.n569 1.16414
R2232 VTAIL.n561 VTAIL.n496 1.16414
R2233 VTAIL.n524 VTAIL.n517 1.16414
R2234 VTAIL.n488 VTAIL.n487 1.16414
R2235 VTAIL.n479 VTAIL.n414 1.16414
R2236 VTAIL.n442 VTAIL.n435 1.16414
R2237 VTAIL.n406 VTAIL.n405 1.16414
R2238 VTAIL.n397 VTAIL.n332 1.16414
R2239 VTAIL.n360 VTAIL.n353 1.16414
R2240 VTAIL.n324 VTAIL.n323 1.16414
R2241 VTAIL.n315 VTAIL.n250 1.16414
R2242 VTAIL.n278 VTAIL.n271 1.16414
R2243 VTAIL VTAIL.n81 0.972483
R2244 VTAIL VTAIL.n655 0.856103
R2245 VTAIL.n491 VTAIL.n409 0.470328
R2246 VTAIL.n163 VTAIL.n81 0.470328
R2247 VTAIL.n602 VTAIL.n601 0.388379
R2248 VTAIL.n647 VTAIL.n646 0.388379
R2249 VTAIL.n648 VTAIL.n576 0.388379
R2250 VTAIL.n28 VTAIL.n27 0.388379
R2251 VTAIL.n73 VTAIL.n72 0.388379
R2252 VTAIL.n74 VTAIL.n2 0.388379
R2253 VTAIL.n110 VTAIL.n109 0.388379
R2254 VTAIL.n155 VTAIL.n154 0.388379
R2255 VTAIL.n156 VTAIL.n84 0.388379
R2256 VTAIL.n192 VTAIL.n191 0.388379
R2257 VTAIL.n237 VTAIL.n236 0.388379
R2258 VTAIL.n238 VTAIL.n166 0.388379
R2259 VTAIL.n566 VTAIL.n494 0.388379
R2260 VTAIL.n565 VTAIL.n564 0.388379
R2261 VTAIL.n521 VTAIL.n520 0.388379
R2262 VTAIL.n484 VTAIL.n412 0.388379
R2263 VTAIL.n483 VTAIL.n482 0.388379
R2264 VTAIL.n439 VTAIL.n438 0.388379
R2265 VTAIL.n402 VTAIL.n330 0.388379
R2266 VTAIL.n401 VTAIL.n400 0.388379
R2267 VTAIL.n357 VTAIL.n356 0.388379
R2268 VTAIL.n320 VTAIL.n248 0.388379
R2269 VTAIL.n319 VTAIL.n318 0.388379
R2270 VTAIL.n275 VTAIL.n274 0.388379
R2271 VTAIL.n604 VTAIL.n603 0.155672
R2272 VTAIL.n604 VTAIL.n595 0.155672
R2273 VTAIL.n611 VTAIL.n595 0.155672
R2274 VTAIL.n612 VTAIL.n611 0.155672
R2275 VTAIL.n612 VTAIL.n591 0.155672
R2276 VTAIL.n619 VTAIL.n591 0.155672
R2277 VTAIL.n620 VTAIL.n619 0.155672
R2278 VTAIL.n620 VTAIL.n587 0.155672
R2279 VTAIL.n627 VTAIL.n587 0.155672
R2280 VTAIL.n628 VTAIL.n627 0.155672
R2281 VTAIL.n628 VTAIL.n583 0.155672
R2282 VTAIL.n635 VTAIL.n583 0.155672
R2283 VTAIL.n636 VTAIL.n635 0.155672
R2284 VTAIL.n636 VTAIL.n579 0.155672
R2285 VTAIL.n644 VTAIL.n579 0.155672
R2286 VTAIL.n645 VTAIL.n644 0.155672
R2287 VTAIL.n645 VTAIL.n575 0.155672
R2288 VTAIL.n653 VTAIL.n575 0.155672
R2289 VTAIL.n30 VTAIL.n29 0.155672
R2290 VTAIL.n30 VTAIL.n21 0.155672
R2291 VTAIL.n37 VTAIL.n21 0.155672
R2292 VTAIL.n38 VTAIL.n37 0.155672
R2293 VTAIL.n38 VTAIL.n17 0.155672
R2294 VTAIL.n45 VTAIL.n17 0.155672
R2295 VTAIL.n46 VTAIL.n45 0.155672
R2296 VTAIL.n46 VTAIL.n13 0.155672
R2297 VTAIL.n53 VTAIL.n13 0.155672
R2298 VTAIL.n54 VTAIL.n53 0.155672
R2299 VTAIL.n54 VTAIL.n9 0.155672
R2300 VTAIL.n61 VTAIL.n9 0.155672
R2301 VTAIL.n62 VTAIL.n61 0.155672
R2302 VTAIL.n62 VTAIL.n5 0.155672
R2303 VTAIL.n70 VTAIL.n5 0.155672
R2304 VTAIL.n71 VTAIL.n70 0.155672
R2305 VTAIL.n71 VTAIL.n1 0.155672
R2306 VTAIL.n79 VTAIL.n1 0.155672
R2307 VTAIL.n112 VTAIL.n111 0.155672
R2308 VTAIL.n112 VTAIL.n103 0.155672
R2309 VTAIL.n119 VTAIL.n103 0.155672
R2310 VTAIL.n120 VTAIL.n119 0.155672
R2311 VTAIL.n120 VTAIL.n99 0.155672
R2312 VTAIL.n127 VTAIL.n99 0.155672
R2313 VTAIL.n128 VTAIL.n127 0.155672
R2314 VTAIL.n128 VTAIL.n95 0.155672
R2315 VTAIL.n135 VTAIL.n95 0.155672
R2316 VTAIL.n136 VTAIL.n135 0.155672
R2317 VTAIL.n136 VTAIL.n91 0.155672
R2318 VTAIL.n143 VTAIL.n91 0.155672
R2319 VTAIL.n144 VTAIL.n143 0.155672
R2320 VTAIL.n144 VTAIL.n87 0.155672
R2321 VTAIL.n152 VTAIL.n87 0.155672
R2322 VTAIL.n153 VTAIL.n152 0.155672
R2323 VTAIL.n153 VTAIL.n83 0.155672
R2324 VTAIL.n161 VTAIL.n83 0.155672
R2325 VTAIL.n194 VTAIL.n193 0.155672
R2326 VTAIL.n194 VTAIL.n185 0.155672
R2327 VTAIL.n201 VTAIL.n185 0.155672
R2328 VTAIL.n202 VTAIL.n201 0.155672
R2329 VTAIL.n202 VTAIL.n181 0.155672
R2330 VTAIL.n209 VTAIL.n181 0.155672
R2331 VTAIL.n210 VTAIL.n209 0.155672
R2332 VTAIL.n210 VTAIL.n177 0.155672
R2333 VTAIL.n217 VTAIL.n177 0.155672
R2334 VTAIL.n218 VTAIL.n217 0.155672
R2335 VTAIL.n218 VTAIL.n173 0.155672
R2336 VTAIL.n225 VTAIL.n173 0.155672
R2337 VTAIL.n226 VTAIL.n225 0.155672
R2338 VTAIL.n226 VTAIL.n169 0.155672
R2339 VTAIL.n234 VTAIL.n169 0.155672
R2340 VTAIL.n235 VTAIL.n234 0.155672
R2341 VTAIL.n235 VTAIL.n165 0.155672
R2342 VTAIL.n243 VTAIL.n165 0.155672
R2343 VTAIL.n571 VTAIL.n493 0.155672
R2344 VTAIL.n563 VTAIL.n493 0.155672
R2345 VTAIL.n563 VTAIL.n562 0.155672
R2346 VTAIL.n562 VTAIL.n497 0.155672
R2347 VTAIL.n555 VTAIL.n497 0.155672
R2348 VTAIL.n555 VTAIL.n554 0.155672
R2349 VTAIL.n554 VTAIL.n502 0.155672
R2350 VTAIL.n547 VTAIL.n502 0.155672
R2351 VTAIL.n547 VTAIL.n546 0.155672
R2352 VTAIL.n546 VTAIL.n506 0.155672
R2353 VTAIL.n539 VTAIL.n506 0.155672
R2354 VTAIL.n539 VTAIL.n538 0.155672
R2355 VTAIL.n538 VTAIL.n510 0.155672
R2356 VTAIL.n531 VTAIL.n510 0.155672
R2357 VTAIL.n531 VTAIL.n530 0.155672
R2358 VTAIL.n530 VTAIL.n514 0.155672
R2359 VTAIL.n523 VTAIL.n514 0.155672
R2360 VTAIL.n523 VTAIL.n522 0.155672
R2361 VTAIL.n489 VTAIL.n411 0.155672
R2362 VTAIL.n481 VTAIL.n411 0.155672
R2363 VTAIL.n481 VTAIL.n480 0.155672
R2364 VTAIL.n480 VTAIL.n415 0.155672
R2365 VTAIL.n473 VTAIL.n415 0.155672
R2366 VTAIL.n473 VTAIL.n472 0.155672
R2367 VTAIL.n472 VTAIL.n420 0.155672
R2368 VTAIL.n465 VTAIL.n420 0.155672
R2369 VTAIL.n465 VTAIL.n464 0.155672
R2370 VTAIL.n464 VTAIL.n424 0.155672
R2371 VTAIL.n457 VTAIL.n424 0.155672
R2372 VTAIL.n457 VTAIL.n456 0.155672
R2373 VTAIL.n456 VTAIL.n428 0.155672
R2374 VTAIL.n449 VTAIL.n428 0.155672
R2375 VTAIL.n449 VTAIL.n448 0.155672
R2376 VTAIL.n448 VTAIL.n432 0.155672
R2377 VTAIL.n441 VTAIL.n432 0.155672
R2378 VTAIL.n441 VTAIL.n440 0.155672
R2379 VTAIL.n407 VTAIL.n329 0.155672
R2380 VTAIL.n399 VTAIL.n329 0.155672
R2381 VTAIL.n399 VTAIL.n398 0.155672
R2382 VTAIL.n398 VTAIL.n333 0.155672
R2383 VTAIL.n391 VTAIL.n333 0.155672
R2384 VTAIL.n391 VTAIL.n390 0.155672
R2385 VTAIL.n390 VTAIL.n338 0.155672
R2386 VTAIL.n383 VTAIL.n338 0.155672
R2387 VTAIL.n383 VTAIL.n382 0.155672
R2388 VTAIL.n382 VTAIL.n342 0.155672
R2389 VTAIL.n375 VTAIL.n342 0.155672
R2390 VTAIL.n375 VTAIL.n374 0.155672
R2391 VTAIL.n374 VTAIL.n346 0.155672
R2392 VTAIL.n367 VTAIL.n346 0.155672
R2393 VTAIL.n367 VTAIL.n366 0.155672
R2394 VTAIL.n366 VTAIL.n350 0.155672
R2395 VTAIL.n359 VTAIL.n350 0.155672
R2396 VTAIL.n359 VTAIL.n358 0.155672
R2397 VTAIL.n325 VTAIL.n247 0.155672
R2398 VTAIL.n317 VTAIL.n247 0.155672
R2399 VTAIL.n317 VTAIL.n316 0.155672
R2400 VTAIL.n316 VTAIL.n251 0.155672
R2401 VTAIL.n309 VTAIL.n251 0.155672
R2402 VTAIL.n309 VTAIL.n308 0.155672
R2403 VTAIL.n308 VTAIL.n256 0.155672
R2404 VTAIL.n301 VTAIL.n256 0.155672
R2405 VTAIL.n301 VTAIL.n300 0.155672
R2406 VTAIL.n300 VTAIL.n260 0.155672
R2407 VTAIL.n293 VTAIL.n260 0.155672
R2408 VTAIL.n293 VTAIL.n292 0.155672
R2409 VTAIL.n292 VTAIL.n264 0.155672
R2410 VTAIL.n285 VTAIL.n264 0.155672
R2411 VTAIL.n285 VTAIL.n284 0.155672
R2412 VTAIL.n284 VTAIL.n268 0.155672
R2413 VTAIL.n277 VTAIL.n268 0.155672
R2414 VTAIL.n277 VTAIL.n276 0.155672
R2415 VN.n0 VN.t2 233.428
R2416 VN.n1 VN.t0 233.428
R2417 VN.n0 VN.t3 232.999
R2418 VN.n1 VN.t1 232.999
R2419 VN VN.n1 55.472
R2420 VN VN.n0 9.36218
R2421 VDD2.n2 VDD2.n0 102.74
R2422 VDD2.n2 VDD2.n1 60.9209
R2423 VDD2.n1 VDD2.t2 1.35296
R2424 VDD2.n1 VDD2.t3 1.35296
R2425 VDD2.n0 VDD2.t1 1.35296
R2426 VDD2.n0 VDD2.t0 1.35296
R2427 VDD2 VDD2.n2 0.0586897
C0 VP VTAIL 4.99187f
C1 VTAIL VDD1 6.15155f
C2 VP VN 6.09936f
C3 VTAIL VDD2 6.20032f
C4 VN VDD1 0.147755f
C5 VN VDD2 5.29054f
C6 VP VDD1 5.4845f
C7 VP VDD2 0.342251f
C8 VN VTAIL 4.97777f
C9 VDD1 VDD2 0.8293f
C10 VDD2 B 3.51303f
C11 VDD1 B 7.67032f
C12 VTAIL B 11.144942f
C13 VN B 9.52396f
C14 VP B 7.380359f
C15 VDD2.t1 B 0.307998f
C16 VDD2.t0 B 0.307998f
C17 VDD2.n0 B 3.50542f
C18 VDD2.t2 B 0.307998f
C19 VDD2.t3 B 0.307998f
C20 VDD2.n1 B 2.78078f
C21 VDD2.n2 B 3.8193f
C22 VN.t2 B 2.40163f
C23 VN.t3 B 2.39987f
C24 VN.n0 B 1.66626f
C25 VN.t0 B 2.40163f
C26 VN.t1 B 2.39987f
C27 VN.n1 B 3.09601f
C28 VTAIL.n0 B 0.019817f
C29 VTAIL.n1 B 0.015596f
C30 VTAIL.n2 B 0.008381f
C31 VTAIL.n3 B 0.019809f
C32 VTAIL.n4 B 0.008874f
C33 VTAIL.n5 B 0.015596f
C34 VTAIL.n6 B 0.008381f
C35 VTAIL.n7 B 0.019809f
C36 VTAIL.n8 B 0.008874f
C37 VTAIL.n9 B 0.015596f
C38 VTAIL.n10 B 0.008381f
C39 VTAIL.n11 B 0.019809f
C40 VTAIL.n12 B 0.008874f
C41 VTAIL.n13 B 0.015596f
C42 VTAIL.n14 B 0.008381f
C43 VTAIL.n15 B 0.019809f
C44 VTAIL.n16 B 0.008874f
C45 VTAIL.n17 B 0.015596f
C46 VTAIL.n18 B 0.008381f
C47 VTAIL.n19 B 0.019809f
C48 VTAIL.n20 B 0.008874f
C49 VTAIL.n21 B 0.015596f
C50 VTAIL.n22 B 0.008381f
C51 VTAIL.n23 B 0.019809f
C52 VTAIL.n24 B 0.008874f
C53 VTAIL.n25 B 0.100313f
C54 VTAIL.t1 B 0.032643f
C55 VTAIL.n26 B 0.014856f
C56 VTAIL.n27 B 0.011702f
C57 VTAIL.n28 B 0.008381f
C58 VTAIL.n29 B 0.988967f
C59 VTAIL.n30 B 0.015596f
C60 VTAIL.n31 B 0.008381f
C61 VTAIL.n32 B 0.008874f
C62 VTAIL.n33 B 0.019809f
C63 VTAIL.n34 B 0.019809f
C64 VTAIL.n35 B 0.008874f
C65 VTAIL.n36 B 0.008381f
C66 VTAIL.n37 B 0.015596f
C67 VTAIL.n38 B 0.015596f
C68 VTAIL.n39 B 0.008381f
C69 VTAIL.n40 B 0.008874f
C70 VTAIL.n41 B 0.019809f
C71 VTAIL.n42 B 0.019809f
C72 VTAIL.n43 B 0.008874f
C73 VTAIL.n44 B 0.008381f
C74 VTAIL.n45 B 0.015596f
C75 VTAIL.n46 B 0.015596f
C76 VTAIL.n47 B 0.008381f
C77 VTAIL.n48 B 0.008874f
C78 VTAIL.n49 B 0.019809f
C79 VTAIL.n50 B 0.019809f
C80 VTAIL.n51 B 0.008874f
C81 VTAIL.n52 B 0.008381f
C82 VTAIL.n53 B 0.015596f
C83 VTAIL.n54 B 0.015596f
C84 VTAIL.n55 B 0.008381f
C85 VTAIL.n56 B 0.008874f
C86 VTAIL.n57 B 0.019809f
C87 VTAIL.n58 B 0.019809f
C88 VTAIL.n59 B 0.008874f
C89 VTAIL.n60 B 0.008381f
C90 VTAIL.n61 B 0.015596f
C91 VTAIL.n62 B 0.015596f
C92 VTAIL.n63 B 0.008381f
C93 VTAIL.n64 B 0.008874f
C94 VTAIL.n65 B 0.019809f
C95 VTAIL.n66 B 0.019809f
C96 VTAIL.n67 B 0.019809f
C97 VTAIL.n68 B 0.008874f
C98 VTAIL.n69 B 0.008381f
C99 VTAIL.n70 B 0.015596f
C100 VTAIL.n71 B 0.015596f
C101 VTAIL.n72 B 0.008381f
C102 VTAIL.n73 B 0.008627f
C103 VTAIL.n74 B 0.008627f
C104 VTAIL.n75 B 0.019809f
C105 VTAIL.n76 B 0.039161f
C106 VTAIL.n77 B 0.008874f
C107 VTAIL.n78 B 0.008381f
C108 VTAIL.n79 B 0.036049f
C109 VTAIL.n80 B 0.02153f
C110 VTAIL.n81 B 0.085777f
C111 VTAIL.n82 B 0.019817f
C112 VTAIL.n83 B 0.015596f
C113 VTAIL.n84 B 0.008381f
C114 VTAIL.n85 B 0.019809f
C115 VTAIL.n86 B 0.008874f
C116 VTAIL.n87 B 0.015596f
C117 VTAIL.n88 B 0.008381f
C118 VTAIL.n89 B 0.019809f
C119 VTAIL.n90 B 0.008874f
C120 VTAIL.n91 B 0.015596f
C121 VTAIL.n92 B 0.008381f
C122 VTAIL.n93 B 0.019809f
C123 VTAIL.n94 B 0.008874f
C124 VTAIL.n95 B 0.015596f
C125 VTAIL.n96 B 0.008381f
C126 VTAIL.n97 B 0.019809f
C127 VTAIL.n98 B 0.008874f
C128 VTAIL.n99 B 0.015596f
C129 VTAIL.n100 B 0.008381f
C130 VTAIL.n101 B 0.019809f
C131 VTAIL.n102 B 0.008874f
C132 VTAIL.n103 B 0.015596f
C133 VTAIL.n104 B 0.008381f
C134 VTAIL.n105 B 0.019809f
C135 VTAIL.n106 B 0.008874f
C136 VTAIL.n107 B 0.100313f
C137 VTAIL.t6 B 0.032643f
C138 VTAIL.n108 B 0.014856f
C139 VTAIL.n109 B 0.011702f
C140 VTAIL.n110 B 0.008381f
C141 VTAIL.n111 B 0.988967f
C142 VTAIL.n112 B 0.015596f
C143 VTAIL.n113 B 0.008381f
C144 VTAIL.n114 B 0.008874f
C145 VTAIL.n115 B 0.019809f
C146 VTAIL.n116 B 0.019809f
C147 VTAIL.n117 B 0.008874f
C148 VTAIL.n118 B 0.008381f
C149 VTAIL.n119 B 0.015596f
C150 VTAIL.n120 B 0.015596f
C151 VTAIL.n121 B 0.008381f
C152 VTAIL.n122 B 0.008874f
C153 VTAIL.n123 B 0.019809f
C154 VTAIL.n124 B 0.019809f
C155 VTAIL.n125 B 0.008874f
C156 VTAIL.n126 B 0.008381f
C157 VTAIL.n127 B 0.015596f
C158 VTAIL.n128 B 0.015596f
C159 VTAIL.n129 B 0.008381f
C160 VTAIL.n130 B 0.008874f
C161 VTAIL.n131 B 0.019809f
C162 VTAIL.n132 B 0.019809f
C163 VTAIL.n133 B 0.008874f
C164 VTAIL.n134 B 0.008381f
C165 VTAIL.n135 B 0.015596f
C166 VTAIL.n136 B 0.015596f
C167 VTAIL.n137 B 0.008381f
C168 VTAIL.n138 B 0.008874f
C169 VTAIL.n139 B 0.019809f
C170 VTAIL.n140 B 0.019809f
C171 VTAIL.n141 B 0.008874f
C172 VTAIL.n142 B 0.008381f
C173 VTAIL.n143 B 0.015596f
C174 VTAIL.n144 B 0.015596f
C175 VTAIL.n145 B 0.008381f
C176 VTAIL.n146 B 0.008874f
C177 VTAIL.n147 B 0.019809f
C178 VTAIL.n148 B 0.019809f
C179 VTAIL.n149 B 0.019809f
C180 VTAIL.n150 B 0.008874f
C181 VTAIL.n151 B 0.008381f
C182 VTAIL.n152 B 0.015596f
C183 VTAIL.n153 B 0.015596f
C184 VTAIL.n154 B 0.008381f
C185 VTAIL.n155 B 0.008627f
C186 VTAIL.n156 B 0.008627f
C187 VTAIL.n157 B 0.019809f
C188 VTAIL.n158 B 0.039161f
C189 VTAIL.n159 B 0.008874f
C190 VTAIL.n160 B 0.008381f
C191 VTAIL.n161 B 0.036049f
C192 VTAIL.n162 B 0.02153f
C193 VTAIL.n163 B 0.128774f
C194 VTAIL.n164 B 0.019817f
C195 VTAIL.n165 B 0.015596f
C196 VTAIL.n166 B 0.008381f
C197 VTAIL.n167 B 0.019809f
C198 VTAIL.n168 B 0.008874f
C199 VTAIL.n169 B 0.015596f
C200 VTAIL.n170 B 0.008381f
C201 VTAIL.n171 B 0.019809f
C202 VTAIL.n172 B 0.008874f
C203 VTAIL.n173 B 0.015596f
C204 VTAIL.n174 B 0.008381f
C205 VTAIL.n175 B 0.019809f
C206 VTAIL.n176 B 0.008874f
C207 VTAIL.n177 B 0.015596f
C208 VTAIL.n178 B 0.008381f
C209 VTAIL.n179 B 0.019809f
C210 VTAIL.n180 B 0.008874f
C211 VTAIL.n181 B 0.015596f
C212 VTAIL.n182 B 0.008381f
C213 VTAIL.n183 B 0.019809f
C214 VTAIL.n184 B 0.008874f
C215 VTAIL.n185 B 0.015596f
C216 VTAIL.n186 B 0.008381f
C217 VTAIL.n187 B 0.019809f
C218 VTAIL.n188 B 0.008874f
C219 VTAIL.n189 B 0.100313f
C220 VTAIL.t7 B 0.032643f
C221 VTAIL.n190 B 0.014856f
C222 VTAIL.n191 B 0.011702f
C223 VTAIL.n192 B 0.008381f
C224 VTAIL.n193 B 0.988967f
C225 VTAIL.n194 B 0.015596f
C226 VTAIL.n195 B 0.008381f
C227 VTAIL.n196 B 0.008874f
C228 VTAIL.n197 B 0.019809f
C229 VTAIL.n198 B 0.019809f
C230 VTAIL.n199 B 0.008874f
C231 VTAIL.n200 B 0.008381f
C232 VTAIL.n201 B 0.015596f
C233 VTAIL.n202 B 0.015596f
C234 VTAIL.n203 B 0.008381f
C235 VTAIL.n204 B 0.008874f
C236 VTAIL.n205 B 0.019809f
C237 VTAIL.n206 B 0.019809f
C238 VTAIL.n207 B 0.008874f
C239 VTAIL.n208 B 0.008381f
C240 VTAIL.n209 B 0.015596f
C241 VTAIL.n210 B 0.015596f
C242 VTAIL.n211 B 0.008381f
C243 VTAIL.n212 B 0.008874f
C244 VTAIL.n213 B 0.019809f
C245 VTAIL.n214 B 0.019809f
C246 VTAIL.n215 B 0.008874f
C247 VTAIL.n216 B 0.008381f
C248 VTAIL.n217 B 0.015596f
C249 VTAIL.n218 B 0.015596f
C250 VTAIL.n219 B 0.008381f
C251 VTAIL.n220 B 0.008874f
C252 VTAIL.n221 B 0.019809f
C253 VTAIL.n222 B 0.019809f
C254 VTAIL.n223 B 0.008874f
C255 VTAIL.n224 B 0.008381f
C256 VTAIL.n225 B 0.015596f
C257 VTAIL.n226 B 0.015596f
C258 VTAIL.n227 B 0.008381f
C259 VTAIL.n228 B 0.008874f
C260 VTAIL.n229 B 0.019809f
C261 VTAIL.n230 B 0.019809f
C262 VTAIL.n231 B 0.019809f
C263 VTAIL.n232 B 0.008874f
C264 VTAIL.n233 B 0.008381f
C265 VTAIL.n234 B 0.015596f
C266 VTAIL.n235 B 0.015596f
C267 VTAIL.n236 B 0.008381f
C268 VTAIL.n237 B 0.008627f
C269 VTAIL.n238 B 0.008627f
C270 VTAIL.n239 B 0.019809f
C271 VTAIL.n240 B 0.039161f
C272 VTAIL.n241 B 0.008874f
C273 VTAIL.n242 B 0.008381f
C274 VTAIL.n243 B 0.036049f
C275 VTAIL.n244 B 0.02153f
C276 VTAIL.n245 B 1.0431f
C277 VTAIL.n246 B 0.019817f
C278 VTAIL.n247 B 0.015596f
C279 VTAIL.n248 B 0.008381f
C280 VTAIL.n249 B 0.019809f
C281 VTAIL.n250 B 0.008874f
C282 VTAIL.n251 B 0.015596f
C283 VTAIL.n252 B 0.008381f
C284 VTAIL.n253 B 0.019809f
C285 VTAIL.n254 B 0.019809f
C286 VTAIL.n255 B 0.008874f
C287 VTAIL.n256 B 0.015596f
C288 VTAIL.n257 B 0.008381f
C289 VTAIL.n258 B 0.019809f
C290 VTAIL.n259 B 0.008874f
C291 VTAIL.n260 B 0.015596f
C292 VTAIL.n261 B 0.008381f
C293 VTAIL.n262 B 0.019809f
C294 VTAIL.n263 B 0.008874f
C295 VTAIL.n264 B 0.015596f
C296 VTAIL.n265 B 0.008381f
C297 VTAIL.n266 B 0.019809f
C298 VTAIL.n267 B 0.008874f
C299 VTAIL.n268 B 0.015596f
C300 VTAIL.n269 B 0.008381f
C301 VTAIL.n270 B 0.019809f
C302 VTAIL.n271 B 0.008874f
C303 VTAIL.n272 B 0.100313f
C304 VTAIL.t2 B 0.032643f
C305 VTAIL.n273 B 0.014856f
C306 VTAIL.n274 B 0.011702f
C307 VTAIL.n275 B 0.008381f
C308 VTAIL.n276 B 0.988967f
C309 VTAIL.n277 B 0.015596f
C310 VTAIL.n278 B 0.008381f
C311 VTAIL.n279 B 0.008874f
C312 VTAIL.n280 B 0.019809f
C313 VTAIL.n281 B 0.019809f
C314 VTAIL.n282 B 0.008874f
C315 VTAIL.n283 B 0.008381f
C316 VTAIL.n284 B 0.015596f
C317 VTAIL.n285 B 0.015596f
C318 VTAIL.n286 B 0.008381f
C319 VTAIL.n287 B 0.008874f
C320 VTAIL.n288 B 0.019809f
C321 VTAIL.n289 B 0.019809f
C322 VTAIL.n290 B 0.008874f
C323 VTAIL.n291 B 0.008381f
C324 VTAIL.n292 B 0.015596f
C325 VTAIL.n293 B 0.015596f
C326 VTAIL.n294 B 0.008381f
C327 VTAIL.n295 B 0.008874f
C328 VTAIL.n296 B 0.019809f
C329 VTAIL.n297 B 0.019809f
C330 VTAIL.n298 B 0.008874f
C331 VTAIL.n299 B 0.008381f
C332 VTAIL.n300 B 0.015596f
C333 VTAIL.n301 B 0.015596f
C334 VTAIL.n302 B 0.008381f
C335 VTAIL.n303 B 0.008874f
C336 VTAIL.n304 B 0.019809f
C337 VTAIL.n305 B 0.019809f
C338 VTAIL.n306 B 0.008874f
C339 VTAIL.n307 B 0.008381f
C340 VTAIL.n308 B 0.015596f
C341 VTAIL.n309 B 0.015596f
C342 VTAIL.n310 B 0.008381f
C343 VTAIL.n311 B 0.008874f
C344 VTAIL.n312 B 0.019809f
C345 VTAIL.n313 B 0.019809f
C346 VTAIL.n314 B 0.008874f
C347 VTAIL.n315 B 0.008381f
C348 VTAIL.n316 B 0.015596f
C349 VTAIL.n317 B 0.015596f
C350 VTAIL.n318 B 0.008381f
C351 VTAIL.n319 B 0.008627f
C352 VTAIL.n320 B 0.008627f
C353 VTAIL.n321 B 0.019809f
C354 VTAIL.n322 B 0.039161f
C355 VTAIL.n323 B 0.008874f
C356 VTAIL.n324 B 0.008381f
C357 VTAIL.n325 B 0.036049f
C358 VTAIL.n326 B 0.02153f
C359 VTAIL.n327 B 1.0431f
C360 VTAIL.n328 B 0.019817f
C361 VTAIL.n329 B 0.015596f
C362 VTAIL.n330 B 0.008381f
C363 VTAIL.n331 B 0.019809f
C364 VTAIL.n332 B 0.008874f
C365 VTAIL.n333 B 0.015596f
C366 VTAIL.n334 B 0.008381f
C367 VTAIL.n335 B 0.019809f
C368 VTAIL.n336 B 0.019809f
C369 VTAIL.n337 B 0.008874f
C370 VTAIL.n338 B 0.015596f
C371 VTAIL.n339 B 0.008381f
C372 VTAIL.n340 B 0.019809f
C373 VTAIL.n341 B 0.008874f
C374 VTAIL.n342 B 0.015596f
C375 VTAIL.n343 B 0.008381f
C376 VTAIL.n344 B 0.019809f
C377 VTAIL.n345 B 0.008874f
C378 VTAIL.n346 B 0.015596f
C379 VTAIL.n347 B 0.008381f
C380 VTAIL.n348 B 0.019809f
C381 VTAIL.n349 B 0.008874f
C382 VTAIL.n350 B 0.015596f
C383 VTAIL.n351 B 0.008381f
C384 VTAIL.n352 B 0.019809f
C385 VTAIL.n353 B 0.008874f
C386 VTAIL.n354 B 0.100313f
C387 VTAIL.t3 B 0.032643f
C388 VTAIL.n355 B 0.014856f
C389 VTAIL.n356 B 0.011702f
C390 VTAIL.n357 B 0.008381f
C391 VTAIL.n358 B 0.988967f
C392 VTAIL.n359 B 0.015596f
C393 VTAIL.n360 B 0.008381f
C394 VTAIL.n361 B 0.008874f
C395 VTAIL.n362 B 0.019809f
C396 VTAIL.n363 B 0.019809f
C397 VTAIL.n364 B 0.008874f
C398 VTAIL.n365 B 0.008381f
C399 VTAIL.n366 B 0.015596f
C400 VTAIL.n367 B 0.015596f
C401 VTAIL.n368 B 0.008381f
C402 VTAIL.n369 B 0.008874f
C403 VTAIL.n370 B 0.019809f
C404 VTAIL.n371 B 0.019809f
C405 VTAIL.n372 B 0.008874f
C406 VTAIL.n373 B 0.008381f
C407 VTAIL.n374 B 0.015596f
C408 VTAIL.n375 B 0.015596f
C409 VTAIL.n376 B 0.008381f
C410 VTAIL.n377 B 0.008874f
C411 VTAIL.n378 B 0.019809f
C412 VTAIL.n379 B 0.019809f
C413 VTAIL.n380 B 0.008874f
C414 VTAIL.n381 B 0.008381f
C415 VTAIL.n382 B 0.015596f
C416 VTAIL.n383 B 0.015596f
C417 VTAIL.n384 B 0.008381f
C418 VTAIL.n385 B 0.008874f
C419 VTAIL.n386 B 0.019809f
C420 VTAIL.n387 B 0.019809f
C421 VTAIL.n388 B 0.008874f
C422 VTAIL.n389 B 0.008381f
C423 VTAIL.n390 B 0.015596f
C424 VTAIL.n391 B 0.015596f
C425 VTAIL.n392 B 0.008381f
C426 VTAIL.n393 B 0.008874f
C427 VTAIL.n394 B 0.019809f
C428 VTAIL.n395 B 0.019809f
C429 VTAIL.n396 B 0.008874f
C430 VTAIL.n397 B 0.008381f
C431 VTAIL.n398 B 0.015596f
C432 VTAIL.n399 B 0.015596f
C433 VTAIL.n400 B 0.008381f
C434 VTAIL.n401 B 0.008627f
C435 VTAIL.n402 B 0.008627f
C436 VTAIL.n403 B 0.019809f
C437 VTAIL.n404 B 0.039161f
C438 VTAIL.n405 B 0.008874f
C439 VTAIL.n406 B 0.008381f
C440 VTAIL.n407 B 0.036049f
C441 VTAIL.n408 B 0.02153f
C442 VTAIL.n409 B 0.128774f
C443 VTAIL.n410 B 0.019817f
C444 VTAIL.n411 B 0.015596f
C445 VTAIL.n412 B 0.008381f
C446 VTAIL.n413 B 0.019809f
C447 VTAIL.n414 B 0.008874f
C448 VTAIL.n415 B 0.015596f
C449 VTAIL.n416 B 0.008381f
C450 VTAIL.n417 B 0.019809f
C451 VTAIL.n418 B 0.019809f
C452 VTAIL.n419 B 0.008874f
C453 VTAIL.n420 B 0.015596f
C454 VTAIL.n421 B 0.008381f
C455 VTAIL.n422 B 0.019809f
C456 VTAIL.n423 B 0.008874f
C457 VTAIL.n424 B 0.015596f
C458 VTAIL.n425 B 0.008381f
C459 VTAIL.n426 B 0.019809f
C460 VTAIL.n427 B 0.008874f
C461 VTAIL.n428 B 0.015596f
C462 VTAIL.n429 B 0.008381f
C463 VTAIL.n430 B 0.019809f
C464 VTAIL.n431 B 0.008874f
C465 VTAIL.n432 B 0.015596f
C466 VTAIL.n433 B 0.008381f
C467 VTAIL.n434 B 0.019809f
C468 VTAIL.n435 B 0.008874f
C469 VTAIL.n436 B 0.100313f
C470 VTAIL.t5 B 0.032643f
C471 VTAIL.n437 B 0.014856f
C472 VTAIL.n438 B 0.011702f
C473 VTAIL.n439 B 0.008381f
C474 VTAIL.n440 B 0.988967f
C475 VTAIL.n441 B 0.015596f
C476 VTAIL.n442 B 0.008381f
C477 VTAIL.n443 B 0.008874f
C478 VTAIL.n444 B 0.019809f
C479 VTAIL.n445 B 0.019809f
C480 VTAIL.n446 B 0.008874f
C481 VTAIL.n447 B 0.008381f
C482 VTAIL.n448 B 0.015596f
C483 VTAIL.n449 B 0.015596f
C484 VTAIL.n450 B 0.008381f
C485 VTAIL.n451 B 0.008874f
C486 VTAIL.n452 B 0.019809f
C487 VTAIL.n453 B 0.019809f
C488 VTAIL.n454 B 0.008874f
C489 VTAIL.n455 B 0.008381f
C490 VTAIL.n456 B 0.015596f
C491 VTAIL.n457 B 0.015596f
C492 VTAIL.n458 B 0.008381f
C493 VTAIL.n459 B 0.008874f
C494 VTAIL.n460 B 0.019809f
C495 VTAIL.n461 B 0.019809f
C496 VTAIL.n462 B 0.008874f
C497 VTAIL.n463 B 0.008381f
C498 VTAIL.n464 B 0.015596f
C499 VTAIL.n465 B 0.015596f
C500 VTAIL.n466 B 0.008381f
C501 VTAIL.n467 B 0.008874f
C502 VTAIL.n468 B 0.019809f
C503 VTAIL.n469 B 0.019809f
C504 VTAIL.n470 B 0.008874f
C505 VTAIL.n471 B 0.008381f
C506 VTAIL.n472 B 0.015596f
C507 VTAIL.n473 B 0.015596f
C508 VTAIL.n474 B 0.008381f
C509 VTAIL.n475 B 0.008874f
C510 VTAIL.n476 B 0.019809f
C511 VTAIL.n477 B 0.019809f
C512 VTAIL.n478 B 0.008874f
C513 VTAIL.n479 B 0.008381f
C514 VTAIL.n480 B 0.015596f
C515 VTAIL.n481 B 0.015596f
C516 VTAIL.n482 B 0.008381f
C517 VTAIL.n483 B 0.008627f
C518 VTAIL.n484 B 0.008627f
C519 VTAIL.n485 B 0.019809f
C520 VTAIL.n486 B 0.039161f
C521 VTAIL.n487 B 0.008874f
C522 VTAIL.n488 B 0.008381f
C523 VTAIL.n489 B 0.036049f
C524 VTAIL.n490 B 0.02153f
C525 VTAIL.n491 B 0.128774f
C526 VTAIL.n492 B 0.019817f
C527 VTAIL.n493 B 0.015596f
C528 VTAIL.n494 B 0.008381f
C529 VTAIL.n495 B 0.019809f
C530 VTAIL.n496 B 0.008874f
C531 VTAIL.n497 B 0.015596f
C532 VTAIL.n498 B 0.008381f
C533 VTAIL.n499 B 0.019809f
C534 VTAIL.n500 B 0.019809f
C535 VTAIL.n501 B 0.008874f
C536 VTAIL.n502 B 0.015596f
C537 VTAIL.n503 B 0.008381f
C538 VTAIL.n504 B 0.019809f
C539 VTAIL.n505 B 0.008874f
C540 VTAIL.n506 B 0.015596f
C541 VTAIL.n507 B 0.008381f
C542 VTAIL.n508 B 0.019809f
C543 VTAIL.n509 B 0.008874f
C544 VTAIL.n510 B 0.015596f
C545 VTAIL.n511 B 0.008381f
C546 VTAIL.n512 B 0.019809f
C547 VTAIL.n513 B 0.008874f
C548 VTAIL.n514 B 0.015596f
C549 VTAIL.n515 B 0.008381f
C550 VTAIL.n516 B 0.019809f
C551 VTAIL.n517 B 0.008874f
C552 VTAIL.n518 B 0.100313f
C553 VTAIL.t4 B 0.032643f
C554 VTAIL.n519 B 0.014856f
C555 VTAIL.n520 B 0.011702f
C556 VTAIL.n521 B 0.008381f
C557 VTAIL.n522 B 0.988967f
C558 VTAIL.n523 B 0.015596f
C559 VTAIL.n524 B 0.008381f
C560 VTAIL.n525 B 0.008874f
C561 VTAIL.n526 B 0.019809f
C562 VTAIL.n527 B 0.019809f
C563 VTAIL.n528 B 0.008874f
C564 VTAIL.n529 B 0.008381f
C565 VTAIL.n530 B 0.015596f
C566 VTAIL.n531 B 0.015596f
C567 VTAIL.n532 B 0.008381f
C568 VTAIL.n533 B 0.008874f
C569 VTAIL.n534 B 0.019809f
C570 VTAIL.n535 B 0.019809f
C571 VTAIL.n536 B 0.008874f
C572 VTAIL.n537 B 0.008381f
C573 VTAIL.n538 B 0.015596f
C574 VTAIL.n539 B 0.015596f
C575 VTAIL.n540 B 0.008381f
C576 VTAIL.n541 B 0.008874f
C577 VTAIL.n542 B 0.019809f
C578 VTAIL.n543 B 0.019809f
C579 VTAIL.n544 B 0.008874f
C580 VTAIL.n545 B 0.008381f
C581 VTAIL.n546 B 0.015596f
C582 VTAIL.n547 B 0.015596f
C583 VTAIL.n548 B 0.008381f
C584 VTAIL.n549 B 0.008874f
C585 VTAIL.n550 B 0.019809f
C586 VTAIL.n551 B 0.019809f
C587 VTAIL.n552 B 0.008874f
C588 VTAIL.n553 B 0.008381f
C589 VTAIL.n554 B 0.015596f
C590 VTAIL.n555 B 0.015596f
C591 VTAIL.n556 B 0.008381f
C592 VTAIL.n557 B 0.008874f
C593 VTAIL.n558 B 0.019809f
C594 VTAIL.n559 B 0.019809f
C595 VTAIL.n560 B 0.008874f
C596 VTAIL.n561 B 0.008381f
C597 VTAIL.n562 B 0.015596f
C598 VTAIL.n563 B 0.015596f
C599 VTAIL.n564 B 0.008381f
C600 VTAIL.n565 B 0.008627f
C601 VTAIL.n566 B 0.008627f
C602 VTAIL.n567 B 0.019809f
C603 VTAIL.n568 B 0.039161f
C604 VTAIL.n569 B 0.008874f
C605 VTAIL.n570 B 0.008381f
C606 VTAIL.n571 B 0.036049f
C607 VTAIL.n572 B 0.02153f
C608 VTAIL.n573 B 1.0431f
C609 VTAIL.n574 B 0.019817f
C610 VTAIL.n575 B 0.015596f
C611 VTAIL.n576 B 0.008381f
C612 VTAIL.n577 B 0.019809f
C613 VTAIL.n578 B 0.008874f
C614 VTAIL.n579 B 0.015596f
C615 VTAIL.n580 B 0.008381f
C616 VTAIL.n581 B 0.019809f
C617 VTAIL.n582 B 0.008874f
C618 VTAIL.n583 B 0.015596f
C619 VTAIL.n584 B 0.008381f
C620 VTAIL.n585 B 0.019809f
C621 VTAIL.n586 B 0.008874f
C622 VTAIL.n587 B 0.015596f
C623 VTAIL.n588 B 0.008381f
C624 VTAIL.n589 B 0.019809f
C625 VTAIL.n590 B 0.008874f
C626 VTAIL.n591 B 0.015596f
C627 VTAIL.n592 B 0.008381f
C628 VTAIL.n593 B 0.019809f
C629 VTAIL.n594 B 0.008874f
C630 VTAIL.n595 B 0.015596f
C631 VTAIL.n596 B 0.008381f
C632 VTAIL.n597 B 0.019809f
C633 VTAIL.n598 B 0.008874f
C634 VTAIL.n599 B 0.100313f
C635 VTAIL.t0 B 0.032643f
C636 VTAIL.n600 B 0.014856f
C637 VTAIL.n601 B 0.011702f
C638 VTAIL.n602 B 0.008381f
C639 VTAIL.n603 B 0.988967f
C640 VTAIL.n604 B 0.015596f
C641 VTAIL.n605 B 0.008381f
C642 VTAIL.n606 B 0.008874f
C643 VTAIL.n607 B 0.019809f
C644 VTAIL.n608 B 0.019809f
C645 VTAIL.n609 B 0.008874f
C646 VTAIL.n610 B 0.008381f
C647 VTAIL.n611 B 0.015596f
C648 VTAIL.n612 B 0.015596f
C649 VTAIL.n613 B 0.008381f
C650 VTAIL.n614 B 0.008874f
C651 VTAIL.n615 B 0.019809f
C652 VTAIL.n616 B 0.019809f
C653 VTAIL.n617 B 0.008874f
C654 VTAIL.n618 B 0.008381f
C655 VTAIL.n619 B 0.015596f
C656 VTAIL.n620 B 0.015596f
C657 VTAIL.n621 B 0.008381f
C658 VTAIL.n622 B 0.008874f
C659 VTAIL.n623 B 0.019809f
C660 VTAIL.n624 B 0.019809f
C661 VTAIL.n625 B 0.008874f
C662 VTAIL.n626 B 0.008381f
C663 VTAIL.n627 B 0.015596f
C664 VTAIL.n628 B 0.015596f
C665 VTAIL.n629 B 0.008381f
C666 VTAIL.n630 B 0.008874f
C667 VTAIL.n631 B 0.019809f
C668 VTAIL.n632 B 0.019809f
C669 VTAIL.n633 B 0.008874f
C670 VTAIL.n634 B 0.008381f
C671 VTAIL.n635 B 0.015596f
C672 VTAIL.n636 B 0.015596f
C673 VTAIL.n637 B 0.008381f
C674 VTAIL.n638 B 0.008874f
C675 VTAIL.n639 B 0.019809f
C676 VTAIL.n640 B 0.019809f
C677 VTAIL.n641 B 0.019809f
C678 VTAIL.n642 B 0.008874f
C679 VTAIL.n643 B 0.008381f
C680 VTAIL.n644 B 0.015596f
C681 VTAIL.n645 B 0.015596f
C682 VTAIL.n646 B 0.008381f
C683 VTAIL.n647 B 0.008627f
C684 VTAIL.n648 B 0.008627f
C685 VTAIL.n649 B 0.019809f
C686 VTAIL.n650 B 0.039161f
C687 VTAIL.n651 B 0.008874f
C688 VTAIL.n652 B 0.008381f
C689 VTAIL.n653 B 0.036049f
C690 VTAIL.n654 B 0.02153f
C691 VTAIL.n655 B 0.994252f
C692 VDD1.t1 B 0.310698f
C693 VDD1.t0 B 0.310698f
C694 VDD1.n0 B 2.80553f
C695 VDD1.t3 B 0.310698f
C696 VDD1.t2 B 0.310698f
C697 VDD1.n1 B 3.56352f
C698 VP.n0 B 0.031871f
C699 VP.t1 B 2.28734f
C700 VP.n1 B 0.025791f
C701 VP.n2 B 0.031871f
C702 VP.t0 B 2.28734f
C703 VP.t2 B 2.43748f
C704 VP.t3 B 2.43569f
C705 VP.n3 B 3.1229f
C706 VP.n4 B 1.83866f
C707 VP.n5 B 0.8806f
C708 VP.n6 B 0.03376f
C709 VP.n7 B 0.063682f
C710 VP.n8 B 0.031871f
C711 VP.n9 B 0.031871f
C712 VP.n10 B 0.031871f
C713 VP.n11 B 0.063682f
C714 VP.n12 B 0.03376f
C715 VP.n13 B 0.8806f
C716 VP.n14 B 0.034117f
.ends

