* NGSPICE file created from diff_pair_sample_1108.ext - technology: sky130A

.subckt diff_pair_sample_1108 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t1 VN.t0 VTAIL.t3 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=2.379 ps=12.98 w=6.1 l=2.97
X1 VDD2.t0 VN.t1 VTAIL.t2 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=2.379 ps=12.98 w=6.1 l=2.97
X2 VDD1.t1 VP.t0 VTAIL.t1 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=2.379 ps=12.98 w=6.1 l=2.97
X3 VDD1.t0 VP.t1 VTAIL.t0 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=2.379 ps=12.98 w=6.1 l=2.97
X4 B.t11 B.t9 B.t10 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=0 ps=0 w=6.1 l=2.97
X5 B.t8 B.t6 B.t7 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=0 ps=0 w=6.1 l=2.97
X6 B.t5 B.t3 B.t4 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=0 ps=0 w=6.1 l=2.97
X7 B.t2 B.t0 B.t1 w_n2290_n2188# sky130_fd_pr__pfet_01v8 ad=2.379 pd=12.98 as=0 ps=0 w=6.1 l=2.97
R0 VN VN.t1 131.806
R1 VN VN.t0 91.0679
R2 VTAIL.n122 VTAIL.n96 756.745
R3 VTAIL.n26 VTAIL.n0 756.745
R4 VTAIL.n90 VTAIL.n64 756.745
R5 VTAIL.n58 VTAIL.n32 756.745
R6 VTAIL.n107 VTAIL.n106 585
R7 VTAIL.n104 VTAIL.n103 585
R8 VTAIL.n113 VTAIL.n112 585
R9 VTAIL.n115 VTAIL.n114 585
R10 VTAIL.n100 VTAIL.n99 585
R11 VTAIL.n121 VTAIL.n120 585
R12 VTAIL.n123 VTAIL.n122 585
R13 VTAIL.n11 VTAIL.n10 585
R14 VTAIL.n8 VTAIL.n7 585
R15 VTAIL.n17 VTAIL.n16 585
R16 VTAIL.n19 VTAIL.n18 585
R17 VTAIL.n4 VTAIL.n3 585
R18 VTAIL.n25 VTAIL.n24 585
R19 VTAIL.n27 VTAIL.n26 585
R20 VTAIL.n91 VTAIL.n90 585
R21 VTAIL.n89 VTAIL.n88 585
R22 VTAIL.n68 VTAIL.n67 585
R23 VTAIL.n83 VTAIL.n82 585
R24 VTAIL.n81 VTAIL.n80 585
R25 VTAIL.n72 VTAIL.n71 585
R26 VTAIL.n75 VTAIL.n74 585
R27 VTAIL.n59 VTAIL.n58 585
R28 VTAIL.n57 VTAIL.n56 585
R29 VTAIL.n36 VTAIL.n35 585
R30 VTAIL.n51 VTAIL.n50 585
R31 VTAIL.n49 VTAIL.n48 585
R32 VTAIL.n40 VTAIL.n39 585
R33 VTAIL.n43 VTAIL.n42 585
R34 VTAIL.t3 VTAIL.n105 327.601
R35 VTAIL.t0 VTAIL.n9 327.601
R36 VTAIL.t1 VTAIL.n73 327.601
R37 VTAIL.t2 VTAIL.n41 327.601
R38 VTAIL.n106 VTAIL.n103 171.744
R39 VTAIL.n113 VTAIL.n103 171.744
R40 VTAIL.n114 VTAIL.n113 171.744
R41 VTAIL.n114 VTAIL.n99 171.744
R42 VTAIL.n121 VTAIL.n99 171.744
R43 VTAIL.n122 VTAIL.n121 171.744
R44 VTAIL.n10 VTAIL.n7 171.744
R45 VTAIL.n17 VTAIL.n7 171.744
R46 VTAIL.n18 VTAIL.n17 171.744
R47 VTAIL.n18 VTAIL.n3 171.744
R48 VTAIL.n25 VTAIL.n3 171.744
R49 VTAIL.n26 VTAIL.n25 171.744
R50 VTAIL.n90 VTAIL.n89 171.744
R51 VTAIL.n89 VTAIL.n67 171.744
R52 VTAIL.n82 VTAIL.n67 171.744
R53 VTAIL.n82 VTAIL.n81 171.744
R54 VTAIL.n81 VTAIL.n71 171.744
R55 VTAIL.n74 VTAIL.n71 171.744
R56 VTAIL.n58 VTAIL.n57 171.744
R57 VTAIL.n57 VTAIL.n35 171.744
R58 VTAIL.n50 VTAIL.n35 171.744
R59 VTAIL.n50 VTAIL.n49 171.744
R60 VTAIL.n49 VTAIL.n39 171.744
R61 VTAIL.n42 VTAIL.n39 171.744
R62 VTAIL.n106 VTAIL.t3 85.8723
R63 VTAIL.n10 VTAIL.t0 85.8723
R64 VTAIL.n74 VTAIL.t1 85.8723
R65 VTAIL.n42 VTAIL.t2 85.8723
R66 VTAIL.n127 VTAIL.n126 34.1247
R67 VTAIL.n31 VTAIL.n30 34.1247
R68 VTAIL.n95 VTAIL.n94 34.1247
R69 VTAIL.n63 VTAIL.n62 34.1247
R70 VTAIL.n63 VTAIL.n31 23.3152
R71 VTAIL.n127 VTAIL.n95 20.4703
R72 VTAIL.n107 VTAIL.n105 16.3865
R73 VTAIL.n11 VTAIL.n9 16.3865
R74 VTAIL.n75 VTAIL.n73 16.3865
R75 VTAIL.n43 VTAIL.n41 16.3865
R76 VTAIL.n108 VTAIL.n104 12.8005
R77 VTAIL.n12 VTAIL.n8 12.8005
R78 VTAIL.n76 VTAIL.n72 12.8005
R79 VTAIL.n44 VTAIL.n40 12.8005
R80 VTAIL.n112 VTAIL.n111 12.0247
R81 VTAIL.n16 VTAIL.n15 12.0247
R82 VTAIL.n80 VTAIL.n79 12.0247
R83 VTAIL.n48 VTAIL.n47 12.0247
R84 VTAIL.n115 VTAIL.n102 11.249
R85 VTAIL.n19 VTAIL.n6 11.249
R86 VTAIL.n83 VTAIL.n70 11.249
R87 VTAIL.n51 VTAIL.n38 11.249
R88 VTAIL.n116 VTAIL.n100 10.4732
R89 VTAIL.n20 VTAIL.n4 10.4732
R90 VTAIL.n84 VTAIL.n68 10.4732
R91 VTAIL.n52 VTAIL.n36 10.4732
R92 VTAIL.n120 VTAIL.n119 9.69747
R93 VTAIL.n24 VTAIL.n23 9.69747
R94 VTAIL.n88 VTAIL.n87 9.69747
R95 VTAIL.n56 VTAIL.n55 9.69747
R96 VTAIL.n126 VTAIL.n125 9.45567
R97 VTAIL.n30 VTAIL.n29 9.45567
R98 VTAIL.n94 VTAIL.n93 9.45567
R99 VTAIL.n62 VTAIL.n61 9.45567
R100 VTAIL.n125 VTAIL.n124 9.3005
R101 VTAIL.n98 VTAIL.n97 9.3005
R102 VTAIL.n119 VTAIL.n118 9.3005
R103 VTAIL.n117 VTAIL.n116 9.3005
R104 VTAIL.n102 VTAIL.n101 9.3005
R105 VTAIL.n111 VTAIL.n110 9.3005
R106 VTAIL.n109 VTAIL.n108 9.3005
R107 VTAIL.n29 VTAIL.n28 9.3005
R108 VTAIL.n2 VTAIL.n1 9.3005
R109 VTAIL.n23 VTAIL.n22 9.3005
R110 VTAIL.n21 VTAIL.n20 9.3005
R111 VTAIL.n6 VTAIL.n5 9.3005
R112 VTAIL.n15 VTAIL.n14 9.3005
R113 VTAIL.n13 VTAIL.n12 9.3005
R114 VTAIL.n93 VTAIL.n92 9.3005
R115 VTAIL.n66 VTAIL.n65 9.3005
R116 VTAIL.n87 VTAIL.n86 9.3005
R117 VTAIL.n85 VTAIL.n84 9.3005
R118 VTAIL.n70 VTAIL.n69 9.3005
R119 VTAIL.n79 VTAIL.n78 9.3005
R120 VTAIL.n77 VTAIL.n76 9.3005
R121 VTAIL.n61 VTAIL.n60 9.3005
R122 VTAIL.n34 VTAIL.n33 9.3005
R123 VTAIL.n55 VTAIL.n54 9.3005
R124 VTAIL.n53 VTAIL.n52 9.3005
R125 VTAIL.n38 VTAIL.n37 9.3005
R126 VTAIL.n47 VTAIL.n46 9.3005
R127 VTAIL.n45 VTAIL.n44 9.3005
R128 VTAIL.n123 VTAIL.n98 8.92171
R129 VTAIL.n27 VTAIL.n2 8.92171
R130 VTAIL.n91 VTAIL.n66 8.92171
R131 VTAIL.n59 VTAIL.n34 8.92171
R132 VTAIL.n124 VTAIL.n96 8.14595
R133 VTAIL.n28 VTAIL.n0 8.14595
R134 VTAIL.n92 VTAIL.n64 8.14595
R135 VTAIL.n60 VTAIL.n32 8.14595
R136 VTAIL.n126 VTAIL.n96 5.81868
R137 VTAIL.n30 VTAIL.n0 5.81868
R138 VTAIL.n94 VTAIL.n64 5.81868
R139 VTAIL.n62 VTAIL.n32 5.81868
R140 VTAIL.n124 VTAIL.n123 5.04292
R141 VTAIL.n28 VTAIL.n27 5.04292
R142 VTAIL.n92 VTAIL.n91 5.04292
R143 VTAIL.n60 VTAIL.n59 5.04292
R144 VTAIL.n120 VTAIL.n98 4.26717
R145 VTAIL.n24 VTAIL.n2 4.26717
R146 VTAIL.n88 VTAIL.n66 4.26717
R147 VTAIL.n56 VTAIL.n34 4.26717
R148 VTAIL.n77 VTAIL.n73 3.71286
R149 VTAIL.n45 VTAIL.n41 3.71286
R150 VTAIL.n109 VTAIL.n105 3.71286
R151 VTAIL.n13 VTAIL.n9 3.71286
R152 VTAIL.n119 VTAIL.n100 3.49141
R153 VTAIL.n23 VTAIL.n4 3.49141
R154 VTAIL.n87 VTAIL.n68 3.49141
R155 VTAIL.n55 VTAIL.n36 3.49141
R156 VTAIL.n116 VTAIL.n115 2.71565
R157 VTAIL.n20 VTAIL.n19 2.71565
R158 VTAIL.n84 VTAIL.n83 2.71565
R159 VTAIL.n52 VTAIL.n51 2.71565
R160 VTAIL.n112 VTAIL.n102 1.93989
R161 VTAIL.n16 VTAIL.n6 1.93989
R162 VTAIL.n80 VTAIL.n70 1.93989
R163 VTAIL.n48 VTAIL.n38 1.93989
R164 VTAIL.n95 VTAIL.n63 1.89274
R165 VTAIL VTAIL.n31 1.23972
R166 VTAIL.n111 VTAIL.n104 1.16414
R167 VTAIL.n15 VTAIL.n8 1.16414
R168 VTAIL.n79 VTAIL.n72 1.16414
R169 VTAIL.n47 VTAIL.n40 1.16414
R170 VTAIL VTAIL.n127 0.653517
R171 VTAIL.n108 VTAIL.n107 0.388379
R172 VTAIL.n12 VTAIL.n11 0.388379
R173 VTAIL.n76 VTAIL.n75 0.388379
R174 VTAIL.n44 VTAIL.n43 0.388379
R175 VTAIL.n110 VTAIL.n109 0.155672
R176 VTAIL.n110 VTAIL.n101 0.155672
R177 VTAIL.n117 VTAIL.n101 0.155672
R178 VTAIL.n118 VTAIL.n117 0.155672
R179 VTAIL.n118 VTAIL.n97 0.155672
R180 VTAIL.n125 VTAIL.n97 0.155672
R181 VTAIL.n14 VTAIL.n13 0.155672
R182 VTAIL.n14 VTAIL.n5 0.155672
R183 VTAIL.n21 VTAIL.n5 0.155672
R184 VTAIL.n22 VTAIL.n21 0.155672
R185 VTAIL.n22 VTAIL.n1 0.155672
R186 VTAIL.n29 VTAIL.n1 0.155672
R187 VTAIL.n93 VTAIL.n65 0.155672
R188 VTAIL.n86 VTAIL.n65 0.155672
R189 VTAIL.n86 VTAIL.n85 0.155672
R190 VTAIL.n85 VTAIL.n69 0.155672
R191 VTAIL.n78 VTAIL.n69 0.155672
R192 VTAIL.n78 VTAIL.n77 0.155672
R193 VTAIL.n61 VTAIL.n33 0.155672
R194 VTAIL.n54 VTAIL.n33 0.155672
R195 VTAIL.n54 VTAIL.n53 0.155672
R196 VTAIL.n53 VTAIL.n37 0.155672
R197 VTAIL.n46 VTAIL.n37 0.155672
R198 VTAIL.n46 VTAIL.n45 0.155672
R199 VDD2.n57 VDD2.n31 756.745
R200 VDD2.n26 VDD2.n0 756.745
R201 VDD2.n58 VDD2.n57 585
R202 VDD2.n56 VDD2.n55 585
R203 VDD2.n35 VDD2.n34 585
R204 VDD2.n50 VDD2.n49 585
R205 VDD2.n48 VDD2.n47 585
R206 VDD2.n39 VDD2.n38 585
R207 VDD2.n42 VDD2.n41 585
R208 VDD2.n11 VDD2.n10 585
R209 VDD2.n8 VDD2.n7 585
R210 VDD2.n17 VDD2.n16 585
R211 VDD2.n19 VDD2.n18 585
R212 VDD2.n4 VDD2.n3 585
R213 VDD2.n25 VDD2.n24 585
R214 VDD2.n27 VDD2.n26 585
R215 VDD2.t0 VDD2.n40 327.601
R216 VDD2.t1 VDD2.n9 327.601
R217 VDD2.n57 VDD2.n56 171.744
R218 VDD2.n56 VDD2.n34 171.744
R219 VDD2.n49 VDD2.n34 171.744
R220 VDD2.n49 VDD2.n48 171.744
R221 VDD2.n48 VDD2.n38 171.744
R222 VDD2.n41 VDD2.n38 171.744
R223 VDD2.n10 VDD2.n7 171.744
R224 VDD2.n17 VDD2.n7 171.744
R225 VDD2.n18 VDD2.n17 171.744
R226 VDD2.n18 VDD2.n3 171.744
R227 VDD2.n25 VDD2.n3 171.744
R228 VDD2.n26 VDD2.n25 171.744
R229 VDD2.n41 VDD2.t0 85.8723
R230 VDD2.n10 VDD2.t1 85.8723
R231 VDD2.n62 VDD2.n30 85.4113
R232 VDD2.n62 VDD2.n61 50.8035
R233 VDD2.n42 VDD2.n40 16.3865
R234 VDD2.n11 VDD2.n9 16.3865
R235 VDD2.n43 VDD2.n39 12.8005
R236 VDD2.n12 VDD2.n8 12.8005
R237 VDD2.n47 VDD2.n46 12.0247
R238 VDD2.n16 VDD2.n15 12.0247
R239 VDD2.n50 VDD2.n37 11.249
R240 VDD2.n19 VDD2.n6 11.249
R241 VDD2.n51 VDD2.n35 10.4732
R242 VDD2.n20 VDD2.n4 10.4732
R243 VDD2.n55 VDD2.n54 9.69747
R244 VDD2.n24 VDD2.n23 9.69747
R245 VDD2.n61 VDD2.n60 9.45567
R246 VDD2.n30 VDD2.n29 9.45567
R247 VDD2.n60 VDD2.n59 9.3005
R248 VDD2.n33 VDD2.n32 9.3005
R249 VDD2.n54 VDD2.n53 9.3005
R250 VDD2.n52 VDD2.n51 9.3005
R251 VDD2.n37 VDD2.n36 9.3005
R252 VDD2.n46 VDD2.n45 9.3005
R253 VDD2.n44 VDD2.n43 9.3005
R254 VDD2.n29 VDD2.n28 9.3005
R255 VDD2.n2 VDD2.n1 9.3005
R256 VDD2.n23 VDD2.n22 9.3005
R257 VDD2.n21 VDD2.n20 9.3005
R258 VDD2.n6 VDD2.n5 9.3005
R259 VDD2.n15 VDD2.n14 9.3005
R260 VDD2.n13 VDD2.n12 9.3005
R261 VDD2.n58 VDD2.n33 8.92171
R262 VDD2.n27 VDD2.n2 8.92171
R263 VDD2.n59 VDD2.n31 8.14595
R264 VDD2.n28 VDD2.n0 8.14595
R265 VDD2.n61 VDD2.n31 5.81868
R266 VDD2.n30 VDD2.n0 5.81868
R267 VDD2.n59 VDD2.n58 5.04292
R268 VDD2.n28 VDD2.n27 5.04292
R269 VDD2.n55 VDD2.n33 4.26717
R270 VDD2.n24 VDD2.n2 4.26717
R271 VDD2.n44 VDD2.n40 3.71286
R272 VDD2.n13 VDD2.n9 3.71286
R273 VDD2.n54 VDD2.n35 3.49141
R274 VDD2.n23 VDD2.n4 3.49141
R275 VDD2.n51 VDD2.n50 2.71565
R276 VDD2.n20 VDD2.n19 2.71565
R277 VDD2.n47 VDD2.n37 1.93989
R278 VDD2.n16 VDD2.n6 1.93989
R279 VDD2.n46 VDD2.n39 1.16414
R280 VDD2.n15 VDD2.n8 1.16414
R281 VDD2 VDD2.n62 0.769897
R282 VDD2.n43 VDD2.n42 0.388379
R283 VDD2.n12 VDD2.n11 0.388379
R284 VDD2.n60 VDD2.n32 0.155672
R285 VDD2.n53 VDD2.n32 0.155672
R286 VDD2.n53 VDD2.n52 0.155672
R287 VDD2.n52 VDD2.n36 0.155672
R288 VDD2.n45 VDD2.n36 0.155672
R289 VDD2.n45 VDD2.n44 0.155672
R290 VDD2.n14 VDD2.n13 0.155672
R291 VDD2.n14 VDD2.n5 0.155672
R292 VDD2.n21 VDD2.n5 0.155672
R293 VDD2.n22 VDD2.n21 0.155672
R294 VDD2.n22 VDD2.n1 0.155672
R295 VDD2.n29 VDD2.n1 0.155672
R296 VP.n0 VP.t0 131.804
R297 VP.n0 VP.t1 90.6366
R298 VP VP.n0 0.431812
R299 VDD1.n26 VDD1.n0 756.745
R300 VDD1.n57 VDD1.n31 756.745
R301 VDD1.n27 VDD1.n26 585
R302 VDD1.n25 VDD1.n24 585
R303 VDD1.n4 VDD1.n3 585
R304 VDD1.n19 VDD1.n18 585
R305 VDD1.n17 VDD1.n16 585
R306 VDD1.n8 VDD1.n7 585
R307 VDD1.n11 VDD1.n10 585
R308 VDD1.n42 VDD1.n41 585
R309 VDD1.n39 VDD1.n38 585
R310 VDD1.n48 VDD1.n47 585
R311 VDD1.n50 VDD1.n49 585
R312 VDD1.n35 VDD1.n34 585
R313 VDD1.n56 VDD1.n55 585
R314 VDD1.n58 VDD1.n57 585
R315 VDD1.t1 VDD1.n9 327.601
R316 VDD1.t0 VDD1.n40 327.601
R317 VDD1.n26 VDD1.n25 171.744
R318 VDD1.n25 VDD1.n3 171.744
R319 VDD1.n18 VDD1.n3 171.744
R320 VDD1.n18 VDD1.n17 171.744
R321 VDD1.n17 VDD1.n7 171.744
R322 VDD1.n10 VDD1.n7 171.744
R323 VDD1.n41 VDD1.n38 171.744
R324 VDD1.n48 VDD1.n38 171.744
R325 VDD1.n49 VDD1.n48 171.744
R326 VDD1.n49 VDD1.n34 171.744
R327 VDD1.n56 VDD1.n34 171.744
R328 VDD1.n57 VDD1.n56 171.744
R329 VDD1 VDD1.n61 86.6473
R330 VDD1.n10 VDD1.t1 85.8723
R331 VDD1.n41 VDD1.t0 85.8723
R332 VDD1 VDD1.n30 51.5729
R333 VDD1.n11 VDD1.n9 16.3865
R334 VDD1.n42 VDD1.n40 16.3865
R335 VDD1.n12 VDD1.n8 12.8005
R336 VDD1.n43 VDD1.n39 12.8005
R337 VDD1.n16 VDD1.n15 12.0247
R338 VDD1.n47 VDD1.n46 12.0247
R339 VDD1.n19 VDD1.n6 11.249
R340 VDD1.n50 VDD1.n37 11.249
R341 VDD1.n20 VDD1.n4 10.4732
R342 VDD1.n51 VDD1.n35 10.4732
R343 VDD1.n24 VDD1.n23 9.69747
R344 VDD1.n55 VDD1.n54 9.69747
R345 VDD1.n30 VDD1.n29 9.45567
R346 VDD1.n61 VDD1.n60 9.45567
R347 VDD1.n29 VDD1.n28 9.3005
R348 VDD1.n2 VDD1.n1 9.3005
R349 VDD1.n23 VDD1.n22 9.3005
R350 VDD1.n21 VDD1.n20 9.3005
R351 VDD1.n6 VDD1.n5 9.3005
R352 VDD1.n15 VDD1.n14 9.3005
R353 VDD1.n13 VDD1.n12 9.3005
R354 VDD1.n60 VDD1.n59 9.3005
R355 VDD1.n33 VDD1.n32 9.3005
R356 VDD1.n54 VDD1.n53 9.3005
R357 VDD1.n52 VDD1.n51 9.3005
R358 VDD1.n37 VDD1.n36 9.3005
R359 VDD1.n46 VDD1.n45 9.3005
R360 VDD1.n44 VDD1.n43 9.3005
R361 VDD1.n27 VDD1.n2 8.92171
R362 VDD1.n58 VDD1.n33 8.92171
R363 VDD1.n28 VDD1.n0 8.14595
R364 VDD1.n59 VDD1.n31 8.14595
R365 VDD1.n30 VDD1.n0 5.81868
R366 VDD1.n61 VDD1.n31 5.81868
R367 VDD1.n28 VDD1.n27 5.04292
R368 VDD1.n59 VDD1.n58 5.04292
R369 VDD1.n24 VDD1.n2 4.26717
R370 VDD1.n55 VDD1.n33 4.26717
R371 VDD1.n13 VDD1.n9 3.71286
R372 VDD1.n44 VDD1.n40 3.71286
R373 VDD1.n23 VDD1.n4 3.49141
R374 VDD1.n54 VDD1.n35 3.49141
R375 VDD1.n20 VDD1.n19 2.71565
R376 VDD1.n51 VDD1.n50 2.71565
R377 VDD1.n16 VDD1.n6 1.93989
R378 VDD1.n47 VDD1.n37 1.93989
R379 VDD1.n15 VDD1.n8 1.16414
R380 VDD1.n46 VDD1.n39 1.16414
R381 VDD1.n12 VDD1.n11 0.388379
R382 VDD1.n43 VDD1.n42 0.388379
R383 VDD1.n29 VDD1.n1 0.155672
R384 VDD1.n22 VDD1.n1 0.155672
R385 VDD1.n22 VDD1.n21 0.155672
R386 VDD1.n21 VDD1.n5 0.155672
R387 VDD1.n14 VDD1.n5 0.155672
R388 VDD1.n14 VDD1.n13 0.155672
R389 VDD1.n45 VDD1.n44 0.155672
R390 VDD1.n45 VDD1.n36 0.155672
R391 VDD1.n52 VDD1.n36 0.155672
R392 VDD1.n53 VDD1.n52 0.155672
R393 VDD1.n53 VDD1.n32 0.155672
R394 VDD1.n60 VDD1.n32 0.155672
R395 B.n251 B.n250 585
R396 B.n249 B.n78 585
R397 B.n248 B.n247 585
R398 B.n246 B.n79 585
R399 B.n245 B.n244 585
R400 B.n243 B.n80 585
R401 B.n242 B.n241 585
R402 B.n240 B.n81 585
R403 B.n239 B.n238 585
R404 B.n237 B.n82 585
R405 B.n236 B.n235 585
R406 B.n234 B.n83 585
R407 B.n233 B.n232 585
R408 B.n231 B.n84 585
R409 B.n230 B.n229 585
R410 B.n228 B.n85 585
R411 B.n227 B.n226 585
R412 B.n225 B.n86 585
R413 B.n224 B.n223 585
R414 B.n222 B.n87 585
R415 B.n221 B.n220 585
R416 B.n219 B.n88 585
R417 B.n218 B.n217 585
R418 B.n216 B.n89 585
R419 B.n215 B.n214 585
R420 B.n210 B.n90 585
R421 B.n209 B.n208 585
R422 B.n207 B.n91 585
R423 B.n206 B.n205 585
R424 B.n204 B.n92 585
R425 B.n203 B.n202 585
R426 B.n201 B.n93 585
R427 B.n200 B.n199 585
R428 B.n198 B.n94 585
R429 B.n196 B.n195 585
R430 B.n194 B.n97 585
R431 B.n193 B.n192 585
R432 B.n191 B.n98 585
R433 B.n190 B.n189 585
R434 B.n188 B.n99 585
R435 B.n187 B.n186 585
R436 B.n185 B.n100 585
R437 B.n184 B.n183 585
R438 B.n182 B.n101 585
R439 B.n181 B.n180 585
R440 B.n179 B.n102 585
R441 B.n178 B.n177 585
R442 B.n176 B.n103 585
R443 B.n175 B.n174 585
R444 B.n173 B.n104 585
R445 B.n172 B.n171 585
R446 B.n170 B.n105 585
R447 B.n169 B.n168 585
R448 B.n167 B.n106 585
R449 B.n166 B.n165 585
R450 B.n164 B.n107 585
R451 B.n163 B.n162 585
R452 B.n161 B.n108 585
R453 B.n252 B.n77 585
R454 B.n254 B.n253 585
R455 B.n255 B.n76 585
R456 B.n257 B.n256 585
R457 B.n258 B.n75 585
R458 B.n260 B.n259 585
R459 B.n261 B.n74 585
R460 B.n263 B.n262 585
R461 B.n264 B.n73 585
R462 B.n266 B.n265 585
R463 B.n267 B.n72 585
R464 B.n269 B.n268 585
R465 B.n270 B.n71 585
R466 B.n272 B.n271 585
R467 B.n273 B.n70 585
R468 B.n275 B.n274 585
R469 B.n276 B.n69 585
R470 B.n278 B.n277 585
R471 B.n279 B.n68 585
R472 B.n281 B.n280 585
R473 B.n282 B.n67 585
R474 B.n284 B.n283 585
R475 B.n285 B.n66 585
R476 B.n287 B.n286 585
R477 B.n288 B.n65 585
R478 B.n290 B.n289 585
R479 B.n291 B.n64 585
R480 B.n293 B.n292 585
R481 B.n294 B.n63 585
R482 B.n296 B.n295 585
R483 B.n297 B.n62 585
R484 B.n299 B.n298 585
R485 B.n300 B.n61 585
R486 B.n302 B.n301 585
R487 B.n303 B.n60 585
R488 B.n305 B.n304 585
R489 B.n306 B.n59 585
R490 B.n308 B.n307 585
R491 B.n309 B.n58 585
R492 B.n311 B.n310 585
R493 B.n312 B.n57 585
R494 B.n314 B.n313 585
R495 B.n315 B.n56 585
R496 B.n317 B.n316 585
R497 B.n318 B.n55 585
R498 B.n320 B.n319 585
R499 B.n321 B.n54 585
R500 B.n323 B.n322 585
R501 B.n324 B.n53 585
R502 B.n326 B.n325 585
R503 B.n327 B.n52 585
R504 B.n329 B.n328 585
R505 B.n330 B.n51 585
R506 B.n332 B.n331 585
R507 B.n333 B.n50 585
R508 B.n335 B.n334 585
R509 B.n423 B.n422 585
R510 B.n421 B.n16 585
R511 B.n420 B.n419 585
R512 B.n418 B.n17 585
R513 B.n417 B.n416 585
R514 B.n415 B.n18 585
R515 B.n414 B.n413 585
R516 B.n412 B.n19 585
R517 B.n411 B.n410 585
R518 B.n409 B.n20 585
R519 B.n408 B.n407 585
R520 B.n406 B.n21 585
R521 B.n405 B.n404 585
R522 B.n403 B.n22 585
R523 B.n402 B.n401 585
R524 B.n400 B.n23 585
R525 B.n399 B.n398 585
R526 B.n397 B.n24 585
R527 B.n396 B.n395 585
R528 B.n394 B.n25 585
R529 B.n393 B.n392 585
R530 B.n391 B.n26 585
R531 B.n390 B.n389 585
R532 B.n388 B.n27 585
R533 B.n386 B.n385 585
R534 B.n384 B.n30 585
R535 B.n383 B.n382 585
R536 B.n381 B.n31 585
R537 B.n380 B.n379 585
R538 B.n378 B.n32 585
R539 B.n377 B.n376 585
R540 B.n375 B.n33 585
R541 B.n374 B.n373 585
R542 B.n372 B.n34 585
R543 B.n371 B.n370 585
R544 B.n369 B.n35 585
R545 B.n368 B.n367 585
R546 B.n366 B.n39 585
R547 B.n365 B.n364 585
R548 B.n363 B.n40 585
R549 B.n362 B.n361 585
R550 B.n360 B.n41 585
R551 B.n359 B.n358 585
R552 B.n357 B.n42 585
R553 B.n356 B.n355 585
R554 B.n354 B.n43 585
R555 B.n353 B.n352 585
R556 B.n351 B.n44 585
R557 B.n350 B.n349 585
R558 B.n348 B.n45 585
R559 B.n347 B.n346 585
R560 B.n345 B.n46 585
R561 B.n344 B.n343 585
R562 B.n342 B.n47 585
R563 B.n341 B.n340 585
R564 B.n339 B.n48 585
R565 B.n338 B.n337 585
R566 B.n336 B.n49 585
R567 B.n424 B.n15 585
R568 B.n426 B.n425 585
R569 B.n427 B.n14 585
R570 B.n429 B.n428 585
R571 B.n430 B.n13 585
R572 B.n432 B.n431 585
R573 B.n433 B.n12 585
R574 B.n435 B.n434 585
R575 B.n436 B.n11 585
R576 B.n438 B.n437 585
R577 B.n439 B.n10 585
R578 B.n441 B.n440 585
R579 B.n442 B.n9 585
R580 B.n444 B.n443 585
R581 B.n445 B.n8 585
R582 B.n447 B.n446 585
R583 B.n448 B.n7 585
R584 B.n450 B.n449 585
R585 B.n451 B.n6 585
R586 B.n453 B.n452 585
R587 B.n454 B.n5 585
R588 B.n456 B.n455 585
R589 B.n457 B.n4 585
R590 B.n459 B.n458 585
R591 B.n460 B.n3 585
R592 B.n462 B.n461 585
R593 B.n463 B.n0 585
R594 B.n2 B.n1 585
R595 B.n122 B.n121 585
R596 B.n124 B.n123 585
R597 B.n125 B.n120 585
R598 B.n127 B.n126 585
R599 B.n128 B.n119 585
R600 B.n130 B.n129 585
R601 B.n131 B.n118 585
R602 B.n133 B.n132 585
R603 B.n134 B.n117 585
R604 B.n136 B.n135 585
R605 B.n137 B.n116 585
R606 B.n139 B.n138 585
R607 B.n140 B.n115 585
R608 B.n142 B.n141 585
R609 B.n143 B.n114 585
R610 B.n145 B.n144 585
R611 B.n146 B.n113 585
R612 B.n148 B.n147 585
R613 B.n149 B.n112 585
R614 B.n151 B.n150 585
R615 B.n152 B.n111 585
R616 B.n154 B.n153 585
R617 B.n155 B.n110 585
R618 B.n157 B.n156 585
R619 B.n158 B.n109 585
R620 B.n160 B.n159 585
R621 B.n159 B.n108 511.721
R622 B.n252 B.n251 511.721
R623 B.n336 B.n335 511.721
R624 B.n422 B.n15 511.721
R625 B.n211 B.t10 334.132
R626 B.n36 B.t8 334.132
R627 B.n95 B.t4 334.132
R628 B.n28 B.t2 334.132
R629 B.n212 B.t11 270.132
R630 B.n37 B.t7 270.132
R631 B.n96 B.t5 270.132
R632 B.n29 B.t1 270.132
R633 B.n95 B.t3 258.043
R634 B.n211 B.t9 258.043
R635 B.n36 B.t6 258.043
R636 B.n28 B.t0 258.043
R637 B.n465 B.n464 256.663
R638 B.n464 B.n463 235.042
R639 B.n464 B.n2 235.042
R640 B.n163 B.n108 163.367
R641 B.n164 B.n163 163.367
R642 B.n165 B.n164 163.367
R643 B.n165 B.n106 163.367
R644 B.n169 B.n106 163.367
R645 B.n170 B.n169 163.367
R646 B.n171 B.n170 163.367
R647 B.n171 B.n104 163.367
R648 B.n175 B.n104 163.367
R649 B.n176 B.n175 163.367
R650 B.n177 B.n176 163.367
R651 B.n177 B.n102 163.367
R652 B.n181 B.n102 163.367
R653 B.n182 B.n181 163.367
R654 B.n183 B.n182 163.367
R655 B.n183 B.n100 163.367
R656 B.n187 B.n100 163.367
R657 B.n188 B.n187 163.367
R658 B.n189 B.n188 163.367
R659 B.n189 B.n98 163.367
R660 B.n193 B.n98 163.367
R661 B.n194 B.n193 163.367
R662 B.n195 B.n194 163.367
R663 B.n195 B.n94 163.367
R664 B.n200 B.n94 163.367
R665 B.n201 B.n200 163.367
R666 B.n202 B.n201 163.367
R667 B.n202 B.n92 163.367
R668 B.n206 B.n92 163.367
R669 B.n207 B.n206 163.367
R670 B.n208 B.n207 163.367
R671 B.n208 B.n90 163.367
R672 B.n215 B.n90 163.367
R673 B.n216 B.n215 163.367
R674 B.n217 B.n216 163.367
R675 B.n217 B.n88 163.367
R676 B.n221 B.n88 163.367
R677 B.n222 B.n221 163.367
R678 B.n223 B.n222 163.367
R679 B.n223 B.n86 163.367
R680 B.n227 B.n86 163.367
R681 B.n228 B.n227 163.367
R682 B.n229 B.n228 163.367
R683 B.n229 B.n84 163.367
R684 B.n233 B.n84 163.367
R685 B.n234 B.n233 163.367
R686 B.n235 B.n234 163.367
R687 B.n235 B.n82 163.367
R688 B.n239 B.n82 163.367
R689 B.n240 B.n239 163.367
R690 B.n241 B.n240 163.367
R691 B.n241 B.n80 163.367
R692 B.n245 B.n80 163.367
R693 B.n246 B.n245 163.367
R694 B.n247 B.n246 163.367
R695 B.n247 B.n78 163.367
R696 B.n251 B.n78 163.367
R697 B.n335 B.n50 163.367
R698 B.n331 B.n50 163.367
R699 B.n331 B.n330 163.367
R700 B.n330 B.n329 163.367
R701 B.n329 B.n52 163.367
R702 B.n325 B.n52 163.367
R703 B.n325 B.n324 163.367
R704 B.n324 B.n323 163.367
R705 B.n323 B.n54 163.367
R706 B.n319 B.n54 163.367
R707 B.n319 B.n318 163.367
R708 B.n318 B.n317 163.367
R709 B.n317 B.n56 163.367
R710 B.n313 B.n56 163.367
R711 B.n313 B.n312 163.367
R712 B.n312 B.n311 163.367
R713 B.n311 B.n58 163.367
R714 B.n307 B.n58 163.367
R715 B.n307 B.n306 163.367
R716 B.n306 B.n305 163.367
R717 B.n305 B.n60 163.367
R718 B.n301 B.n60 163.367
R719 B.n301 B.n300 163.367
R720 B.n300 B.n299 163.367
R721 B.n299 B.n62 163.367
R722 B.n295 B.n62 163.367
R723 B.n295 B.n294 163.367
R724 B.n294 B.n293 163.367
R725 B.n293 B.n64 163.367
R726 B.n289 B.n64 163.367
R727 B.n289 B.n288 163.367
R728 B.n288 B.n287 163.367
R729 B.n287 B.n66 163.367
R730 B.n283 B.n66 163.367
R731 B.n283 B.n282 163.367
R732 B.n282 B.n281 163.367
R733 B.n281 B.n68 163.367
R734 B.n277 B.n68 163.367
R735 B.n277 B.n276 163.367
R736 B.n276 B.n275 163.367
R737 B.n275 B.n70 163.367
R738 B.n271 B.n70 163.367
R739 B.n271 B.n270 163.367
R740 B.n270 B.n269 163.367
R741 B.n269 B.n72 163.367
R742 B.n265 B.n72 163.367
R743 B.n265 B.n264 163.367
R744 B.n264 B.n263 163.367
R745 B.n263 B.n74 163.367
R746 B.n259 B.n74 163.367
R747 B.n259 B.n258 163.367
R748 B.n258 B.n257 163.367
R749 B.n257 B.n76 163.367
R750 B.n253 B.n76 163.367
R751 B.n253 B.n252 163.367
R752 B.n422 B.n421 163.367
R753 B.n421 B.n420 163.367
R754 B.n420 B.n17 163.367
R755 B.n416 B.n17 163.367
R756 B.n416 B.n415 163.367
R757 B.n415 B.n414 163.367
R758 B.n414 B.n19 163.367
R759 B.n410 B.n19 163.367
R760 B.n410 B.n409 163.367
R761 B.n409 B.n408 163.367
R762 B.n408 B.n21 163.367
R763 B.n404 B.n21 163.367
R764 B.n404 B.n403 163.367
R765 B.n403 B.n402 163.367
R766 B.n402 B.n23 163.367
R767 B.n398 B.n23 163.367
R768 B.n398 B.n397 163.367
R769 B.n397 B.n396 163.367
R770 B.n396 B.n25 163.367
R771 B.n392 B.n25 163.367
R772 B.n392 B.n391 163.367
R773 B.n391 B.n390 163.367
R774 B.n390 B.n27 163.367
R775 B.n385 B.n27 163.367
R776 B.n385 B.n384 163.367
R777 B.n384 B.n383 163.367
R778 B.n383 B.n31 163.367
R779 B.n379 B.n31 163.367
R780 B.n379 B.n378 163.367
R781 B.n378 B.n377 163.367
R782 B.n377 B.n33 163.367
R783 B.n373 B.n33 163.367
R784 B.n373 B.n372 163.367
R785 B.n372 B.n371 163.367
R786 B.n371 B.n35 163.367
R787 B.n367 B.n35 163.367
R788 B.n367 B.n366 163.367
R789 B.n366 B.n365 163.367
R790 B.n365 B.n40 163.367
R791 B.n361 B.n40 163.367
R792 B.n361 B.n360 163.367
R793 B.n360 B.n359 163.367
R794 B.n359 B.n42 163.367
R795 B.n355 B.n42 163.367
R796 B.n355 B.n354 163.367
R797 B.n354 B.n353 163.367
R798 B.n353 B.n44 163.367
R799 B.n349 B.n44 163.367
R800 B.n349 B.n348 163.367
R801 B.n348 B.n347 163.367
R802 B.n347 B.n46 163.367
R803 B.n343 B.n46 163.367
R804 B.n343 B.n342 163.367
R805 B.n342 B.n341 163.367
R806 B.n341 B.n48 163.367
R807 B.n337 B.n48 163.367
R808 B.n337 B.n336 163.367
R809 B.n426 B.n15 163.367
R810 B.n427 B.n426 163.367
R811 B.n428 B.n427 163.367
R812 B.n428 B.n13 163.367
R813 B.n432 B.n13 163.367
R814 B.n433 B.n432 163.367
R815 B.n434 B.n433 163.367
R816 B.n434 B.n11 163.367
R817 B.n438 B.n11 163.367
R818 B.n439 B.n438 163.367
R819 B.n440 B.n439 163.367
R820 B.n440 B.n9 163.367
R821 B.n444 B.n9 163.367
R822 B.n445 B.n444 163.367
R823 B.n446 B.n445 163.367
R824 B.n446 B.n7 163.367
R825 B.n450 B.n7 163.367
R826 B.n451 B.n450 163.367
R827 B.n452 B.n451 163.367
R828 B.n452 B.n5 163.367
R829 B.n456 B.n5 163.367
R830 B.n457 B.n456 163.367
R831 B.n458 B.n457 163.367
R832 B.n458 B.n3 163.367
R833 B.n462 B.n3 163.367
R834 B.n463 B.n462 163.367
R835 B.n122 B.n2 163.367
R836 B.n123 B.n122 163.367
R837 B.n123 B.n120 163.367
R838 B.n127 B.n120 163.367
R839 B.n128 B.n127 163.367
R840 B.n129 B.n128 163.367
R841 B.n129 B.n118 163.367
R842 B.n133 B.n118 163.367
R843 B.n134 B.n133 163.367
R844 B.n135 B.n134 163.367
R845 B.n135 B.n116 163.367
R846 B.n139 B.n116 163.367
R847 B.n140 B.n139 163.367
R848 B.n141 B.n140 163.367
R849 B.n141 B.n114 163.367
R850 B.n145 B.n114 163.367
R851 B.n146 B.n145 163.367
R852 B.n147 B.n146 163.367
R853 B.n147 B.n112 163.367
R854 B.n151 B.n112 163.367
R855 B.n152 B.n151 163.367
R856 B.n153 B.n152 163.367
R857 B.n153 B.n110 163.367
R858 B.n157 B.n110 163.367
R859 B.n158 B.n157 163.367
R860 B.n159 B.n158 163.367
R861 B.n96 B.n95 64.0005
R862 B.n212 B.n211 64.0005
R863 B.n37 B.n36 64.0005
R864 B.n29 B.n28 64.0005
R865 B.n197 B.n96 59.5399
R866 B.n213 B.n212 59.5399
R867 B.n38 B.n37 59.5399
R868 B.n387 B.n29 59.5399
R869 B.n424 B.n423 33.2493
R870 B.n334 B.n49 33.2493
R871 B.n250 B.n77 33.2493
R872 B.n161 B.n160 33.2493
R873 B B.n465 18.0485
R874 B.n425 B.n424 10.6151
R875 B.n425 B.n14 10.6151
R876 B.n429 B.n14 10.6151
R877 B.n430 B.n429 10.6151
R878 B.n431 B.n430 10.6151
R879 B.n431 B.n12 10.6151
R880 B.n435 B.n12 10.6151
R881 B.n436 B.n435 10.6151
R882 B.n437 B.n436 10.6151
R883 B.n437 B.n10 10.6151
R884 B.n441 B.n10 10.6151
R885 B.n442 B.n441 10.6151
R886 B.n443 B.n442 10.6151
R887 B.n443 B.n8 10.6151
R888 B.n447 B.n8 10.6151
R889 B.n448 B.n447 10.6151
R890 B.n449 B.n448 10.6151
R891 B.n449 B.n6 10.6151
R892 B.n453 B.n6 10.6151
R893 B.n454 B.n453 10.6151
R894 B.n455 B.n454 10.6151
R895 B.n455 B.n4 10.6151
R896 B.n459 B.n4 10.6151
R897 B.n460 B.n459 10.6151
R898 B.n461 B.n460 10.6151
R899 B.n461 B.n0 10.6151
R900 B.n423 B.n16 10.6151
R901 B.n419 B.n16 10.6151
R902 B.n419 B.n418 10.6151
R903 B.n418 B.n417 10.6151
R904 B.n417 B.n18 10.6151
R905 B.n413 B.n18 10.6151
R906 B.n413 B.n412 10.6151
R907 B.n412 B.n411 10.6151
R908 B.n411 B.n20 10.6151
R909 B.n407 B.n20 10.6151
R910 B.n407 B.n406 10.6151
R911 B.n406 B.n405 10.6151
R912 B.n405 B.n22 10.6151
R913 B.n401 B.n22 10.6151
R914 B.n401 B.n400 10.6151
R915 B.n400 B.n399 10.6151
R916 B.n399 B.n24 10.6151
R917 B.n395 B.n24 10.6151
R918 B.n395 B.n394 10.6151
R919 B.n394 B.n393 10.6151
R920 B.n393 B.n26 10.6151
R921 B.n389 B.n26 10.6151
R922 B.n389 B.n388 10.6151
R923 B.n386 B.n30 10.6151
R924 B.n382 B.n30 10.6151
R925 B.n382 B.n381 10.6151
R926 B.n381 B.n380 10.6151
R927 B.n380 B.n32 10.6151
R928 B.n376 B.n32 10.6151
R929 B.n376 B.n375 10.6151
R930 B.n375 B.n374 10.6151
R931 B.n374 B.n34 10.6151
R932 B.n370 B.n369 10.6151
R933 B.n369 B.n368 10.6151
R934 B.n368 B.n39 10.6151
R935 B.n364 B.n39 10.6151
R936 B.n364 B.n363 10.6151
R937 B.n363 B.n362 10.6151
R938 B.n362 B.n41 10.6151
R939 B.n358 B.n41 10.6151
R940 B.n358 B.n357 10.6151
R941 B.n357 B.n356 10.6151
R942 B.n356 B.n43 10.6151
R943 B.n352 B.n43 10.6151
R944 B.n352 B.n351 10.6151
R945 B.n351 B.n350 10.6151
R946 B.n350 B.n45 10.6151
R947 B.n346 B.n45 10.6151
R948 B.n346 B.n345 10.6151
R949 B.n345 B.n344 10.6151
R950 B.n344 B.n47 10.6151
R951 B.n340 B.n47 10.6151
R952 B.n340 B.n339 10.6151
R953 B.n339 B.n338 10.6151
R954 B.n338 B.n49 10.6151
R955 B.n334 B.n333 10.6151
R956 B.n333 B.n332 10.6151
R957 B.n332 B.n51 10.6151
R958 B.n328 B.n51 10.6151
R959 B.n328 B.n327 10.6151
R960 B.n327 B.n326 10.6151
R961 B.n326 B.n53 10.6151
R962 B.n322 B.n53 10.6151
R963 B.n322 B.n321 10.6151
R964 B.n321 B.n320 10.6151
R965 B.n320 B.n55 10.6151
R966 B.n316 B.n55 10.6151
R967 B.n316 B.n315 10.6151
R968 B.n315 B.n314 10.6151
R969 B.n314 B.n57 10.6151
R970 B.n310 B.n57 10.6151
R971 B.n310 B.n309 10.6151
R972 B.n309 B.n308 10.6151
R973 B.n308 B.n59 10.6151
R974 B.n304 B.n59 10.6151
R975 B.n304 B.n303 10.6151
R976 B.n303 B.n302 10.6151
R977 B.n302 B.n61 10.6151
R978 B.n298 B.n61 10.6151
R979 B.n298 B.n297 10.6151
R980 B.n297 B.n296 10.6151
R981 B.n296 B.n63 10.6151
R982 B.n292 B.n63 10.6151
R983 B.n292 B.n291 10.6151
R984 B.n291 B.n290 10.6151
R985 B.n290 B.n65 10.6151
R986 B.n286 B.n65 10.6151
R987 B.n286 B.n285 10.6151
R988 B.n285 B.n284 10.6151
R989 B.n284 B.n67 10.6151
R990 B.n280 B.n67 10.6151
R991 B.n280 B.n279 10.6151
R992 B.n279 B.n278 10.6151
R993 B.n278 B.n69 10.6151
R994 B.n274 B.n69 10.6151
R995 B.n274 B.n273 10.6151
R996 B.n273 B.n272 10.6151
R997 B.n272 B.n71 10.6151
R998 B.n268 B.n71 10.6151
R999 B.n268 B.n267 10.6151
R1000 B.n267 B.n266 10.6151
R1001 B.n266 B.n73 10.6151
R1002 B.n262 B.n73 10.6151
R1003 B.n262 B.n261 10.6151
R1004 B.n261 B.n260 10.6151
R1005 B.n260 B.n75 10.6151
R1006 B.n256 B.n75 10.6151
R1007 B.n256 B.n255 10.6151
R1008 B.n255 B.n254 10.6151
R1009 B.n254 B.n77 10.6151
R1010 B.n121 B.n1 10.6151
R1011 B.n124 B.n121 10.6151
R1012 B.n125 B.n124 10.6151
R1013 B.n126 B.n125 10.6151
R1014 B.n126 B.n119 10.6151
R1015 B.n130 B.n119 10.6151
R1016 B.n131 B.n130 10.6151
R1017 B.n132 B.n131 10.6151
R1018 B.n132 B.n117 10.6151
R1019 B.n136 B.n117 10.6151
R1020 B.n137 B.n136 10.6151
R1021 B.n138 B.n137 10.6151
R1022 B.n138 B.n115 10.6151
R1023 B.n142 B.n115 10.6151
R1024 B.n143 B.n142 10.6151
R1025 B.n144 B.n143 10.6151
R1026 B.n144 B.n113 10.6151
R1027 B.n148 B.n113 10.6151
R1028 B.n149 B.n148 10.6151
R1029 B.n150 B.n149 10.6151
R1030 B.n150 B.n111 10.6151
R1031 B.n154 B.n111 10.6151
R1032 B.n155 B.n154 10.6151
R1033 B.n156 B.n155 10.6151
R1034 B.n156 B.n109 10.6151
R1035 B.n160 B.n109 10.6151
R1036 B.n162 B.n161 10.6151
R1037 B.n162 B.n107 10.6151
R1038 B.n166 B.n107 10.6151
R1039 B.n167 B.n166 10.6151
R1040 B.n168 B.n167 10.6151
R1041 B.n168 B.n105 10.6151
R1042 B.n172 B.n105 10.6151
R1043 B.n173 B.n172 10.6151
R1044 B.n174 B.n173 10.6151
R1045 B.n174 B.n103 10.6151
R1046 B.n178 B.n103 10.6151
R1047 B.n179 B.n178 10.6151
R1048 B.n180 B.n179 10.6151
R1049 B.n180 B.n101 10.6151
R1050 B.n184 B.n101 10.6151
R1051 B.n185 B.n184 10.6151
R1052 B.n186 B.n185 10.6151
R1053 B.n186 B.n99 10.6151
R1054 B.n190 B.n99 10.6151
R1055 B.n191 B.n190 10.6151
R1056 B.n192 B.n191 10.6151
R1057 B.n192 B.n97 10.6151
R1058 B.n196 B.n97 10.6151
R1059 B.n199 B.n198 10.6151
R1060 B.n199 B.n93 10.6151
R1061 B.n203 B.n93 10.6151
R1062 B.n204 B.n203 10.6151
R1063 B.n205 B.n204 10.6151
R1064 B.n205 B.n91 10.6151
R1065 B.n209 B.n91 10.6151
R1066 B.n210 B.n209 10.6151
R1067 B.n214 B.n210 10.6151
R1068 B.n218 B.n89 10.6151
R1069 B.n219 B.n218 10.6151
R1070 B.n220 B.n219 10.6151
R1071 B.n220 B.n87 10.6151
R1072 B.n224 B.n87 10.6151
R1073 B.n225 B.n224 10.6151
R1074 B.n226 B.n225 10.6151
R1075 B.n226 B.n85 10.6151
R1076 B.n230 B.n85 10.6151
R1077 B.n231 B.n230 10.6151
R1078 B.n232 B.n231 10.6151
R1079 B.n232 B.n83 10.6151
R1080 B.n236 B.n83 10.6151
R1081 B.n237 B.n236 10.6151
R1082 B.n238 B.n237 10.6151
R1083 B.n238 B.n81 10.6151
R1084 B.n242 B.n81 10.6151
R1085 B.n243 B.n242 10.6151
R1086 B.n244 B.n243 10.6151
R1087 B.n244 B.n79 10.6151
R1088 B.n248 B.n79 10.6151
R1089 B.n249 B.n248 10.6151
R1090 B.n250 B.n249 10.6151
R1091 B.n388 B.n387 9.36635
R1092 B.n370 B.n38 9.36635
R1093 B.n197 B.n196 9.36635
R1094 B.n213 B.n89 9.36635
R1095 B.n465 B.n0 8.11757
R1096 B.n465 B.n1 8.11757
R1097 B.n387 B.n386 1.24928
R1098 B.n38 B.n34 1.24928
R1099 B.n198 B.n197 1.24928
R1100 B.n214 B.n213 1.24928
C0 w_n2290_n2188# VN 3.08378f
C1 VP VTAIL 1.63917f
C2 VP VDD1 1.76603f
C3 B VP 1.52472f
C4 w_n2290_n2188# VDD2 1.44555f
C5 VN VDD2 1.56758f
C6 w_n2290_n2188# VTAIL 1.93083f
C7 w_n2290_n2188# VDD1 1.41511f
C8 w_n2290_n2188# B 7.56528f
C9 VN VTAIL 1.62498f
C10 VDD1 VN 0.148626f
C11 B VN 1.04236f
C12 VDD2 VTAIL 3.65801f
C13 VDD1 VDD2 0.718877f
C14 B VDD2 1.31893f
C15 w_n2290_n2188# VP 3.37628f
C16 VDD1 VTAIL 3.60335f
C17 B VTAIL 2.43713f
C18 B VDD1 1.28556f
C19 VP VN 4.53242f
C20 VP VDD2 0.348513f
C21 VDD2 VSUBS 0.692872f
C22 VDD1 VSUBS 2.435767f
C23 VTAIL VSUBS 0.556264f
C24 VN VSUBS 5.49905f
C25 VP VSUBS 1.456554f
C26 B VSUBS 3.682775f
C27 w_n2290_n2188# VSUBS 62.517002f
C28 B.n0 VSUBS 0.006752f
C29 B.n1 VSUBS 0.006752f
C30 B.n2 VSUBS 0.009986f
C31 B.n3 VSUBS 0.007652f
C32 B.n4 VSUBS 0.007652f
C33 B.n5 VSUBS 0.007652f
C34 B.n6 VSUBS 0.007652f
C35 B.n7 VSUBS 0.007652f
C36 B.n8 VSUBS 0.007652f
C37 B.n9 VSUBS 0.007652f
C38 B.n10 VSUBS 0.007652f
C39 B.n11 VSUBS 0.007652f
C40 B.n12 VSUBS 0.007652f
C41 B.n13 VSUBS 0.007652f
C42 B.n14 VSUBS 0.007652f
C43 B.n15 VSUBS 0.017717f
C44 B.n16 VSUBS 0.007652f
C45 B.n17 VSUBS 0.007652f
C46 B.n18 VSUBS 0.007652f
C47 B.n19 VSUBS 0.007652f
C48 B.n20 VSUBS 0.007652f
C49 B.n21 VSUBS 0.007652f
C50 B.n22 VSUBS 0.007652f
C51 B.n23 VSUBS 0.007652f
C52 B.n24 VSUBS 0.007652f
C53 B.n25 VSUBS 0.007652f
C54 B.n26 VSUBS 0.007652f
C55 B.n27 VSUBS 0.007652f
C56 B.t1 VSUBS 0.099984f
C57 B.t2 VSUBS 0.131316f
C58 B.t0 VSUBS 0.941915f
C59 B.n28 VSUBS 0.22073f
C60 B.n29 VSUBS 0.174492f
C61 B.n30 VSUBS 0.007652f
C62 B.n31 VSUBS 0.007652f
C63 B.n32 VSUBS 0.007652f
C64 B.n33 VSUBS 0.007652f
C65 B.n34 VSUBS 0.004276f
C66 B.n35 VSUBS 0.007652f
C67 B.t7 VSUBS 0.099986f
C68 B.t8 VSUBS 0.131317f
C69 B.t6 VSUBS 0.941915f
C70 B.n36 VSUBS 0.220728f
C71 B.n37 VSUBS 0.17449f
C72 B.n38 VSUBS 0.01773f
C73 B.n39 VSUBS 0.007652f
C74 B.n40 VSUBS 0.007652f
C75 B.n41 VSUBS 0.007652f
C76 B.n42 VSUBS 0.007652f
C77 B.n43 VSUBS 0.007652f
C78 B.n44 VSUBS 0.007652f
C79 B.n45 VSUBS 0.007652f
C80 B.n46 VSUBS 0.007652f
C81 B.n47 VSUBS 0.007652f
C82 B.n48 VSUBS 0.007652f
C83 B.n49 VSUBS 0.018519f
C84 B.n50 VSUBS 0.007652f
C85 B.n51 VSUBS 0.007652f
C86 B.n52 VSUBS 0.007652f
C87 B.n53 VSUBS 0.007652f
C88 B.n54 VSUBS 0.007652f
C89 B.n55 VSUBS 0.007652f
C90 B.n56 VSUBS 0.007652f
C91 B.n57 VSUBS 0.007652f
C92 B.n58 VSUBS 0.007652f
C93 B.n59 VSUBS 0.007652f
C94 B.n60 VSUBS 0.007652f
C95 B.n61 VSUBS 0.007652f
C96 B.n62 VSUBS 0.007652f
C97 B.n63 VSUBS 0.007652f
C98 B.n64 VSUBS 0.007652f
C99 B.n65 VSUBS 0.007652f
C100 B.n66 VSUBS 0.007652f
C101 B.n67 VSUBS 0.007652f
C102 B.n68 VSUBS 0.007652f
C103 B.n69 VSUBS 0.007652f
C104 B.n70 VSUBS 0.007652f
C105 B.n71 VSUBS 0.007652f
C106 B.n72 VSUBS 0.007652f
C107 B.n73 VSUBS 0.007652f
C108 B.n74 VSUBS 0.007652f
C109 B.n75 VSUBS 0.007652f
C110 B.n76 VSUBS 0.007652f
C111 B.n77 VSUBS 0.018605f
C112 B.n78 VSUBS 0.007652f
C113 B.n79 VSUBS 0.007652f
C114 B.n80 VSUBS 0.007652f
C115 B.n81 VSUBS 0.007652f
C116 B.n82 VSUBS 0.007652f
C117 B.n83 VSUBS 0.007652f
C118 B.n84 VSUBS 0.007652f
C119 B.n85 VSUBS 0.007652f
C120 B.n86 VSUBS 0.007652f
C121 B.n87 VSUBS 0.007652f
C122 B.n88 VSUBS 0.007652f
C123 B.n89 VSUBS 0.007202f
C124 B.n90 VSUBS 0.007652f
C125 B.n91 VSUBS 0.007652f
C126 B.n92 VSUBS 0.007652f
C127 B.n93 VSUBS 0.007652f
C128 B.n94 VSUBS 0.007652f
C129 B.t5 VSUBS 0.099984f
C130 B.t4 VSUBS 0.131316f
C131 B.t3 VSUBS 0.941915f
C132 B.n95 VSUBS 0.22073f
C133 B.n96 VSUBS 0.174492f
C134 B.n97 VSUBS 0.007652f
C135 B.n98 VSUBS 0.007652f
C136 B.n99 VSUBS 0.007652f
C137 B.n100 VSUBS 0.007652f
C138 B.n101 VSUBS 0.007652f
C139 B.n102 VSUBS 0.007652f
C140 B.n103 VSUBS 0.007652f
C141 B.n104 VSUBS 0.007652f
C142 B.n105 VSUBS 0.007652f
C143 B.n106 VSUBS 0.007652f
C144 B.n107 VSUBS 0.007652f
C145 B.n108 VSUBS 0.018519f
C146 B.n109 VSUBS 0.007652f
C147 B.n110 VSUBS 0.007652f
C148 B.n111 VSUBS 0.007652f
C149 B.n112 VSUBS 0.007652f
C150 B.n113 VSUBS 0.007652f
C151 B.n114 VSUBS 0.007652f
C152 B.n115 VSUBS 0.007652f
C153 B.n116 VSUBS 0.007652f
C154 B.n117 VSUBS 0.007652f
C155 B.n118 VSUBS 0.007652f
C156 B.n119 VSUBS 0.007652f
C157 B.n120 VSUBS 0.007652f
C158 B.n121 VSUBS 0.007652f
C159 B.n122 VSUBS 0.007652f
C160 B.n123 VSUBS 0.007652f
C161 B.n124 VSUBS 0.007652f
C162 B.n125 VSUBS 0.007652f
C163 B.n126 VSUBS 0.007652f
C164 B.n127 VSUBS 0.007652f
C165 B.n128 VSUBS 0.007652f
C166 B.n129 VSUBS 0.007652f
C167 B.n130 VSUBS 0.007652f
C168 B.n131 VSUBS 0.007652f
C169 B.n132 VSUBS 0.007652f
C170 B.n133 VSUBS 0.007652f
C171 B.n134 VSUBS 0.007652f
C172 B.n135 VSUBS 0.007652f
C173 B.n136 VSUBS 0.007652f
C174 B.n137 VSUBS 0.007652f
C175 B.n138 VSUBS 0.007652f
C176 B.n139 VSUBS 0.007652f
C177 B.n140 VSUBS 0.007652f
C178 B.n141 VSUBS 0.007652f
C179 B.n142 VSUBS 0.007652f
C180 B.n143 VSUBS 0.007652f
C181 B.n144 VSUBS 0.007652f
C182 B.n145 VSUBS 0.007652f
C183 B.n146 VSUBS 0.007652f
C184 B.n147 VSUBS 0.007652f
C185 B.n148 VSUBS 0.007652f
C186 B.n149 VSUBS 0.007652f
C187 B.n150 VSUBS 0.007652f
C188 B.n151 VSUBS 0.007652f
C189 B.n152 VSUBS 0.007652f
C190 B.n153 VSUBS 0.007652f
C191 B.n154 VSUBS 0.007652f
C192 B.n155 VSUBS 0.007652f
C193 B.n156 VSUBS 0.007652f
C194 B.n157 VSUBS 0.007652f
C195 B.n158 VSUBS 0.007652f
C196 B.n159 VSUBS 0.017717f
C197 B.n160 VSUBS 0.017717f
C198 B.n161 VSUBS 0.018519f
C199 B.n162 VSUBS 0.007652f
C200 B.n163 VSUBS 0.007652f
C201 B.n164 VSUBS 0.007652f
C202 B.n165 VSUBS 0.007652f
C203 B.n166 VSUBS 0.007652f
C204 B.n167 VSUBS 0.007652f
C205 B.n168 VSUBS 0.007652f
C206 B.n169 VSUBS 0.007652f
C207 B.n170 VSUBS 0.007652f
C208 B.n171 VSUBS 0.007652f
C209 B.n172 VSUBS 0.007652f
C210 B.n173 VSUBS 0.007652f
C211 B.n174 VSUBS 0.007652f
C212 B.n175 VSUBS 0.007652f
C213 B.n176 VSUBS 0.007652f
C214 B.n177 VSUBS 0.007652f
C215 B.n178 VSUBS 0.007652f
C216 B.n179 VSUBS 0.007652f
C217 B.n180 VSUBS 0.007652f
C218 B.n181 VSUBS 0.007652f
C219 B.n182 VSUBS 0.007652f
C220 B.n183 VSUBS 0.007652f
C221 B.n184 VSUBS 0.007652f
C222 B.n185 VSUBS 0.007652f
C223 B.n186 VSUBS 0.007652f
C224 B.n187 VSUBS 0.007652f
C225 B.n188 VSUBS 0.007652f
C226 B.n189 VSUBS 0.007652f
C227 B.n190 VSUBS 0.007652f
C228 B.n191 VSUBS 0.007652f
C229 B.n192 VSUBS 0.007652f
C230 B.n193 VSUBS 0.007652f
C231 B.n194 VSUBS 0.007652f
C232 B.n195 VSUBS 0.007652f
C233 B.n196 VSUBS 0.007202f
C234 B.n197 VSUBS 0.01773f
C235 B.n198 VSUBS 0.004276f
C236 B.n199 VSUBS 0.007652f
C237 B.n200 VSUBS 0.007652f
C238 B.n201 VSUBS 0.007652f
C239 B.n202 VSUBS 0.007652f
C240 B.n203 VSUBS 0.007652f
C241 B.n204 VSUBS 0.007652f
C242 B.n205 VSUBS 0.007652f
C243 B.n206 VSUBS 0.007652f
C244 B.n207 VSUBS 0.007652f
C245 B.n208 VSUBS 0.007652f
C246 B.n209 VSUBS 0.007652f
C247 B.n210 VSUBS 0.007652f
C248 B.t11 VSUBS 0.099986f
C249 B.t10 VSUBS 0.131317f
C250 B.t9 VSUBS 0.941915f
C251 B.n211 VSUBS 0.220728f
C252 B.n212 VSUBS 0.17449f
C253 B.n213 VSUBS 0.01773f
C254 B.n214 VSUBS 0.004276f
C255 B.n215 VSUBS 0.007652f
C256 B.n216 VSUBS 0.007652f
C257 B.n217 VSUBS 0.007652f
C258 B.n218 VSUBS 0.007652f
C259 B.n219 VSUBS 0.007652f
C260 B.n220 VSUBS 0.007652f
C261 B.n221 VSUBS 0.007652f
C262 B.n222 VSUBS 0.007652f
C263 B.n223 VSUBS 0.007652f
C264 B.n224 VSUBS 0.007652f
C265 B.n225 VSUBS 0.007652f
C266 B.n226 VSUBS 0.007652f
C267 B.n227 VSUBS 0.007652f
C268 B.n228 VSUBS 0.007652f
C269 B.n229 VSUBS 0.007652f
C270 B.n230 VSUBS 0.007652f
C271 B.n231 VSUBS 0.007652f
C272 B.n232 VSUBS 0.007652f
C273 B.n233 VSUBS 0.007652f
C274 B.n234 VSUBS 0.007652f
C275 B.n235 VSUBS 0.007652f
C276 B.n236 VSUBS 0.007652f
C277 B.n237 VSUBS 0.007652f
C278 B.n238 VSUBS 0.007652f
C279 B.n239 VSUBS 0.007652f
C280 B.n240 VSUBS 0.007652f
C281 B.n241 VSUBS 0.007652f
C282 B.n242 VSUBS 0.007652f
C283 B.n243 VSUBS 0.007652f
C284 B.n244 VSUBS 0.007652f
C285 B.n245 VSUBS 0.007652f
C286 B.n246 VSUBS 0.007652f
C287 B.n247 VSUBS 0.007652f
C288 B.n248 VSUBS 0.007652f
C289 B.n249 VSUBS 0.007652f
C290 B.n250 VSUBS 0.017631f
C291 B.n251 VSUBS 0.018519f
C292 B.n252 VSUBS 0.017717f
C293 B.n253 VSUBS 0.007652f
C294 B.n254 VSUBS 0.007652f
C295 B.n255 VSUBS 0.007652f
C296 B.n256 VSUBS 0.007652f
C297 B.n257 VSUBS 0.007652f
C298 B.n258 VSUBS 0.007652f
C299 B.n259 VSUBS 0.007652f
C300 B.n260 VSUBS 0.007652f
C301 B.n261 VSUBS 0.007652f
C302 B.n262 VSUBS 0.007652f
C303 B.n263 VSUBS 0.007652f
C304 B.n264 VSUBS 0.007652f
C305 B.n265 VSUBS 0.007652f
C306 B.n266 VSUBS 0.007652f
C307 B.n267 VSUBS 0.007652f
C308 B.n268 VSUBS 0.007652f
C309 B.n269 VSUBS 0.007652f
C310 B.n270 VSUBS 0.007652f
C311 B.n271 VSUBS 0.007652f
C312 B.n272 VSUBS 0.007652f
C313 B.n273 VSUBS 0.007652f
C314 B.n274 VSUBS 0.007652f
C315 B.n275 VSUBS 0.007652f
C316 B.n276 VSUBS 0.007652f
C317 B.n277 VSUBS 0.007652f
C318 B.n278 VSUBS 0.007652f
C319 B.n279 VSUBS 0.007652f
C320 B.n280 VSUBS 0.007652f
C321 B.n281 VSUBS 0.007652f
C322 B.n282 VSUBS 0.007652f
C323 B.n283 VSUBS 0.007652f
C324 B.n284 VSUBS 0.007652f
C325 B.n285 VSUBS 0.007652f
C326 B.n286 VSUBS 0.007652f
C327 B.n287 VSUBS 0.007652f
C328 B.n288 VSUBS 0.007652f
C329 B.n289 VSUBS 0.007652f
C330 B.n290 VSUBS 0.007652f
C331 B.n291 VSUBS 0.007652f
C332 B.n292 VSUBS 0.007652f
C333 B.n293 VSUBS 0.007652f
C334 B.n294 VSUBS 0.007652f
C335 B.n295 VSUBS 0.007652f
C336 B.n296 VSUBS 0.007652f
C337 B.n297 VSUBS 0.007652f
C338 B.n298 VSUBS 0.007652f
C339 B.n299 VSUBS 0.007652f
C340 B.n300 VSUBS 0.007652f
C341 B.n301 VSUBS 0.007652f
C342 B.n302 VSUBS 0.007652f
C343 B.n303 VSUBS 0.007652f
C344 B.n304 VSUBS 0.007652f
C345 B.n305 VSUBS 0.007652f
C346 B.n306 VSUBS 0.007652f
C347 B.n307 VSUBS 0.007652f
C348 B.n308 VSUBS 0.007652f
C349 B.n309 VSUBS 0.007652f
C350 B.n310 VSUBS 0.007652f
C351 B.n311 VSUBS 0.007652f
C352 B.n312 VSUBS 0.007652f
C353 B.n313 VSUBS 0.007652f
C354 B.n314 VSUBS 0.007652f
C355 B.n315 VSUBS 0.007652f
C356 B.n316 VSUBS 0.007652f
C357 B.n317 VSUBS 0.007652f
C358 B.n318 VSUBS 0.007652f
C359 B.n319 VSUBS 0.007652f
C360 B.n320 VSUBS 0.007652f
C361 B.n321 VSUBS 0.007652f
C362 B.n322 VSUBS 0.007652f
C363 B.n323 VSUBS 0.007652f
C364 B.n324 VSUBS 0.007652f
C365 B.n325 VSUBS 0.007652f
C366 B.n326 VSUBS 0.007652f
C367 B.n327 VSUBS 0.007652f
C368 B.n328 VSUBS 0.007652f
C369 B.n329 VSUBS 0.007652f
C370 B.n330 VSUBS 0.007652f
C371 B.n331 VSUBS 0.007652f
C372 B.n332 VSUBS 0.007652f
C373 B.n333 VSUBS 0.007652f
C374 B.n334 VSUBS 0.017717f
C375 B.n335 VSUBS 0.017717f
C376 B.n336 VSUBS 0.018519f
C377 B.n337 VSUBS 0.007652f
C378 B.n338 VSUBS 0.007652f
C379 B.n339 VSUBS 0.007652f
C380 B.n340 VSUBS 0.007652f
C381 B.n341 VSUBS 0.007652f
C382 B.n342 VSUBS 0.007652f
C383 B.n343 VSUBS 0.007652f
C384 B.n344 VSUBS 0.007652f
C385 B.n345 VSUBS 0.007652f
C386 B.n346 VSUBS 0.007652f
C387 B.n347 VSUBS 0.007652f
C388 B.n348 VSUBS 0.007652f
C389 B.n349 VSUBS 0.007652f
C390 B.n350 VSUBS 0.007652f
C391 B.n351 VSUBS 0.007652f
C392 B.n352 VSUBS 0.007652f
C393 B.n353 VSUBS 0.007652f
C394 B.n354 VSUBS 0.007652f
C395 B.n355 VSUBS 0.007652f
C396 B.n356 VSUBS 0.007652f
C397 B.n357 VSUBS 0.007652f
C398 B.n358 VSUBS 0.007652f
C399 B.n359 VSUBS 0.007652f
C400 B.n360 VSUBS 0.007652f
C401 B.n361 VSUBS 0.007652f
C402 B.n362 VSUBS 0.007652f
C403 B.n363 VSUBS 0.007652f
C404 B.n364 VSUBS 0.007652f
C405 B.n365 VSUBS 0.007652f
C406 B.n366 VSUBS 0.007652f
C407 B.n367 VSUBS 0.007652f
C408 B.n368 VSUBS 0.007652f
C409 B.n369 VSUBS 0.007652f
C410 B.n370 VSUBS 0.007202f
C411 B.n371 VSUBS 0.007652f
C412 B.n372 VSUBS 0.007652f
C413 B.n373 VSUBS 0.007652f
C414 B.n374 VSUBS 0.007652f
C415 B.n375 VSUBS 0.007652f
C416 B.n376 VSUBS 0.007652f
C417 B.n377 VSUBS 0.007652f
C418 B.n378 VSUBS 0.007652f
C419 B.n379 VSUBS 0.007652f
C420 B.n380 VSUBS 0.007652f
C421 B.n381 VSUBS 0.007652f
C422 B.n382 VSUBS 0.007652f
C423 B.n383 VSUBS 0.007652f
C424 B.n384 VSUBS 0.007652f
C425 B.n385 VSUBS 0.007652f
C426 B.n386 VSUBS 0.004276f
C427 B.n387 VSUBS 0.01773f
C428 B.n388 VSUBS 0.007202f
C429 B.n389 VSUBS 0.007652f
C430 B.n390 VSUBS 0.007652f
C431 B.n391 VSUBS 0.007652f
C432 B.n392 VSUBS 0.007652f
C433 B.n393 VSUBS 0.007652f
C434 B.n394 VSUBS 0.007652f
C435 B.n395 VSUBS 0.007652f
C436 B.n396 VSUBS 0.007652f
C437 B.n397 VSUBS 0.007652f
C438 B.n398 VSUBS 0.007652f
C439 B.n399 VSUBS 0.007652f
C440 B.n400 VSUBS 0.007652f
C441 B.n401 VSUBS 0.007652f
C442 B.n402 VSUBS 0.007652f
C443 B.n403 VSUBS 0.007652f
C444 B.n404 VSUBS 0.007652f
C445 B.n405 VSUBS 0.007652f
C446 B.n406 VSUBS 0.007652f
C447 B.n407 VSUBS 0.007652f
C448 B.n408 VSUBS 0.007652f
C449 B.n409 VSUBS 0.007652f
C450 B.n410 VSUBS 0.007652f
C451 B.n411 VSUBS 0.007652f
C452 B.n412 VSUBS 0.007652f
C453 B.n413 VSUBS 0.007652f
C454 B.n414 VSUBS 0.007652f
C455 B.n415 VSUBS 0.007652f
C456 B.n416 VSUBS 0.007652f
C457 B.n417 VSUBS 0.007652f
C458 B.n418 VSUBS 0.007652f
C459 B.n419 VSUBS 0.007652f
C460 B.n420 VSUBS 0.007652f
C461 B.n421 VSUBS 0.007652f
C462 B.n422 VSUBS 0.018519f
C463 B.n423 VSUBS 0.018519f
C464 B.n424 VSUBS 0.017717f
C465 B.n425 VSUBS 0.007652f
C466 B.n426 VSUBS 0.007652f
C467 B.n427 VSUBS 0.007652f
C468 B.n428 VSUBS 0.007652f
C469 B.n429 VSUBS 0.007652f
C470 B.n430 VSUBS 0.007652f
C471 B.n431 VSUBS 0.007652f
C472 B.n432 VSUBS 0.007652f
C473 B.n433 VSUBS 0.007652f
C474 B.n434 VSUBS 0.007652f
C475 B.n435 VSUBS 0.007652f
C476 B.n436 VSUBS 0.007652f
C477 B.n437 VSUBS 0.007652f
C478 B.n438 VSUBS 0.007652f
C479 B.n439 VSUBS 0.007652f
C480 B.n440 VSUBS 0.007652f
C481 B.n441 VSUBS 0.007652f
C482 B.n442 VSUBS 0.007652f
C483 B.n443 VSUBS 0.007652f
C484 B.n444 VSUBS 0.007652f
C485 B.n445 VSUBS 0.007652f
C486 B.n446 VSUBS 0.007652f
C487 B.n447 VSUBS 0.007652f
C488 B.n448 VSUBS 0.007652f
C489 B.n449 VSUBS 0.007652f
C490 B.n450 VSUBS 0.007652f
C491 B.n451 VSUBS 0.007652f
C492 B.n452 VSUBS 0.007652f
C493 B.n453 VSUBS 0.007652f
C494 B.n454 VSUBS 0.007652f
C495 B.n455 VSUBS 0.007652f
C496 B.n456 VSUBS 0.007652f
C497 B.n457 VSUBS 0.007652f
C498 B.n458 VSUBS 0.007652f
C499 B.n459 VSUBS 0.007652f
C500 B.n460 VSUBS 0.007652f
C501 B.n461 VSUBS 0.007652f
C502 B.n462 VSUBS 0.007652f
C503 B.n463 VSUBS 0.009986f
C504 B.n464 VSUBS 0.010637f
C505 B.n465 VSUBS 0.021154f
C506 VDD1.n0 VSUBS 0.016293f
C507 VDD1.n1 VSUBS 0.01433f
C508 VDD1.n2 VSUBS 0.0077f
C509 VDD1.n3 VSUBS 0.018201f
C510 VDD1.n4 VSUBS 0.008153f
C511 VDD1.n5 VSUBS 0.01433f
C512 VDD1.n6 VSUBS 0.0077f
C513 VDD1.n7 VSUBS 0.018201f
C514 VDD1.n8 VSUBS 0.008153f
C515 VDD1.n9 VSUBS 0.063861f
C516 VDD1.t1 VSUBS 0.039136f
C517 VDD1.n10 VSUBS 0.013651f
C518 VDD1.n11 VSUBS 0.011572f
C519 VDD1.n12 VSUBS 0.0077f
C520 VDD1.n13 VSUBS 0.335077f
C521 VDD1.n14 VSUBS 0.01433f
C522 VDD1.n15 VSUBS 0.0077f
C523 VDD1.n16 VSUBS 0.008153f
C524 VDD1.n17 VSUBS 0.018201f
C525 VDD1.n18 VSUBS 0.018201f
C526 VDD1.n19 VSUBS 0.008153f
C527 VDD1.n20 VSUBS 0.0077f
C528 VDD1.n21 VSUBS 0.01433f
C529 VDD1.n22 VSUBS 0.01433f
C530 VDD1.n23 VSUBS 0.0077f
C531 VDD1.n24 VSUBS 0.008153f
C532 VDD1.n25 VSUBS 0.018201f
C533 VDD1.n26 VSUBS 0.045928f
C534 VDD1.n27 VSUBS 0.008153f
C535 VDD1.n28 VSUBS 0.0077f
C536 VDD1.n29 VSUBS 0.035081f
C537 VDD1.n30 VSUBS 0.034077f
C538 VDD1.n31 VSUBS 0.016293f
C539 VDD1.n32 VSUBS 0.01433f
C540 VDD1.n33 VSUBS 0.0077f
C541 VDD1.n34 VSUBS 0.018201f
C542 VDD1.n35 VSUBS 0.008153f
C543 VDD1.n36 VSUBS 0.01433f
C544 VDD1.n37 VSUBS 0.0077f
C545 VDD1.n38 VSUBS 0.018201f
C546 VDD1.n39 VSUBS 0.008153f
C547 VDD1.n40 VSUBS 0.063861f
C548 VDD1.t0 VSUBS 0.039136f
C549 VDD1.n41 VSUBS 0.013651f
C550 VDD1.n42 VSUBS 0.011572f
C551 VDD1.n43 VSUBS 0.0077f
C552 VDD1.n44 VSUBS 0.335077f
C553 VDD1.n45 VSUBS 0.01433f
C554 VDD1.n46 VSUBS 0.0077f
C555 VDD1.n47 VSUBS 0.008153f
C556 VDD1.n48 VSUBS 0.018201f
C557 VDD1.n49 VSUBS 0.018201f
C558 VDD1.n50 VSUBS 0.008153f
C559 VDD1.n51 VSUBS 0.0077f
C560 VDD1.n52 VSUBS 0.01433f
C561 VDD1.n53 VSUBS 0.01433f
C562 VDD1.n54 VSUBS 0.0077f
C563 VDD1.n55 VSUBS 0.008153f
C564 VDD1.n56 VSUBS 0.018201f
C565 VDD1.n57 VSUBS 0.045928f
C566 VDD1.n58 VSUBS 0.008153f
C567 VDD1.n59 VSUBS 0.0077f
C568 VDD1.n60 VSUBS 0.035081f
C569 VDD1.n61 VSUBS 0.342289f
C570 VP.t1 VSUBS 1.96953f
C571 VP.t0 VSUBS 2.5836f
C572 VP.n0 VSUBS 3.24924f
C573 VDD2.n0 VSUBS 0.016996f
C574 VDD2.n1 VSUBS 0.014948f
C575 VDD2.n2 VSUBS 0.008032f
C576 VDD2.n3 VSUBS 0.018986f
C577 VDD2.n4 VSUBS 0.008505f
C578 VDD2.n5 VSUBS 0.014948f
C579 VDD2.n6 VSUBS 0.008032f
C580 VDD2.n7 VSUBS 0.018986f
C581 VDD2.n8 VSUBS 0.008505f
C582 VDD2.n9 VSUBS 0.066614f
C583 VDD2.t1 VSUBS 0.040823f
C584 VDD2.n10 VSUBS 0.014239f
C585 VDD2.n11 VSUBS 0.012071f
C586 VDD2.n12 VSUBS 0.008032f
C587 VDD2.n13 VSUBS 0.349524f
C588 VDD2.n14 VSUBS 0.014948f
C589 VDD2.n15 VSUBS 0.008032f
C590 VDD2.n16 VSUBS 0.008505f
C591 VDD2.n17 VSUBS 0.018986f
C592 VDD2.n18 VSUBS 0.018986f
C593 VDD2.n19 VSUBS 0.008505f
C594 VDD2.n20 VSUBS 0.008032f
C595 VDD2.n21 VSUBS 0.014948f
C596 VDD2.n22 VSUBS 0.014948f
C597 VDD2.n23 VSUBS 0.008032f
C598 VDD2.n24 VSUBS 0.008505f
C599 VDD2.n25 VSUBS 0.018986f
C600 VDD2.n26 VSUBS 0.047908f
C601 VDD2.n27 VSUBS 0.008505f
C602 VDD2.n28 VSUBS 0.008032f
C603 VDD2.n29 VSUBS 0.036594f
C604 VDD2.n30 VSUBS 0.329729f
C605 VDD2.n31 VSUBS 0.016996f
C606 VDD2.n32 VSUBS 0.014948f
C607 VDD2.n33 VSUBS 0.008032f
C608 VDD2.n34 VSUBS 0.018986f
C609 VDD2.n35 VSUBS 0.008505f
C610 VDD2.n36 VSUBS 0.014948f
C611 VDD2.n37 VSUBS 0.008032f
C612 VDD2.n38 VSUBS 0.018986f
C613 VDD2.n39 VSUBS 0.008505f
C614 VDD2.n40 VSUBS 0.066614f
C615 VDD2.t0 VSUBS 0.040823f
C616 VDD2.n41 VSUBS 0.014239f
C617 VDD2.n42 VSUBS 0.012071f
C618 VDD2.n43 VSUBS 0.008032f
C619 VDD2.n44 VSUBS 0.349524f
C620 VDD2.n45 VSUBS 0.014948f
C621 VDD2.n46 VSUBS 0.008032f
C622 VDD2.n47 VSUBS 0.008505f
C623 VDD2.n48 VSUBS 0.018986f
C624 VDD2.n49 VSUBS 0.018986f
C625 VDD2.n50 VSUBS 0.008505f
C626 VDD2.n51 VSUBS 0.008032f
C627 VDD2.n52 VSUBS 0.014948f
C628 VDD2.n53 VSUBS 0.014948f
C629 VDD2.n54 VSUBS 0.008032f
C630 VDD2.n55 VSUBS 0.008505f
C631 VDD2.n56 VSUBS 0.018986f
C632 VDD2.n57 VSUBS 0.047908f
C633 VDD2.n58 VSUBS 0.008505f
C634 VDD2.n59 VSUBS 0.008032f
C635 VDD2.n60 VSUBS 0.036594f
C636 VDD2.n61 VSUBS 0.034546f
C637 VDD2.n62 VSUBS 1.50635f
C638 VTAIL.n0 VSUBS 0.024935f
C639 VTAIL.n1 VSUBS 0.021931f
C640 VTAIL.n2 VSUBS 0.011785f
C641 VTAIL.n3 VSUBS 0.027855f
C642 VTAIL.n4 VSUBS 0.012478f
C643 VTAIL.n5 VSUBS 0.021931f
C644 VTAIL.n6 VSUBS 0.011785f
C645 VTAIL.n7 VSUBS 0.027855f
C646 VTAIL.n8 VSUBS 0.012478f
C647 VTAIL.n9 VSUBS 0.097733f
C648 VTAIL.t0 VSUBS 0.059893f
C649 VTAIL.n10 VSUBS 0.020891f
C650 VTAIL.n11 VSUBS 0.017711f
C651 VTAIL.n12 VSUBS 0.011785f
C652 VTAIL.n13 VSUBS 0.512801f
C653 VTAIL.n14 VSUBS 0.021931f
C654 VTAIL.n15 VSUBS 0.011785f
C655 VTAIL.n16 VSUBS 0.012478f
C656 VTAIL.n17 VSUBS 0.027855f
C657 VTAIL.n18 VSUBS 0.027855f
C658 VTAIL.n19 VSUBS 0.012478f
C659 VTAIL.n20 VSUBS 0.011785f
C660 VTAIL.n21 VSUBS 0.021931f
C661 VTAIL.n22 VSUBS 0.021931f
C662 VTAIL.n23 VSUBS 0.011785f
C663 VTAIL.n24 VSUBS 0.012478f
C664 VTAIL.n25 VSUBS 0.027855f
C665 VTAIL.n26 VSUBS 0.070288f
C666 VTAIL.n27 VSUBS 0.012478f
C667 VTAIL.n28 VSUBS 0.011785f
C668 VTAIL.n29 VSUBS 0.053688f
C669 VTAIL.n30 VSUBS 0.035564f
C670 VTAIL.n31 VSUBS 1.17958f
C671 VTAIL.n32 VSUBS 0.024935f
C672 VTAIL.n33 VSUBS 0.021931f
C673 VTAIL.n34 VSUBS 0.011785f
C674 VTAIL.n35 VSUBS 0.027855f
C675 VTAIL.n36 VSUBS 0.012478f
C676 VTAIL.n37 VSUBS 0.021931f
C677 VTAIL.n38 VSUBS 0.011785f
C678 VTAIL.n39 VSUBS 0.027855f
C679 VTAIL.n40 VSUBS 0.012478f
C680 VTAIL.n41 VSUBS 0.097733f
C681 VTAIL.t2 VSUBS 0.059893f
C682 VTAIL.n42 VSUBS 0.020891f
C683 VTAIL.n43 VSUBS 0.017711f
C684 VTAIL.n44 VSUBS 0.011785f
C685 VTAIL.n45 VSUBS 0.512801f
C686 VTAIL.n46 VSUBS 0.021931f
C687 VTAIL.n47 VSUBS 0.011785f
C688 VTAIL.n48 VSUBS 0.012478f
C689 VTAIL.n49 VSUBS 0.027855f
C690 VTAIL.n50 VSUBS 0.027855f
C691 VTAIL.n51 VSUBS 0.012478f
C692 VTAIL.n52 VSUBS 0.011785f
C693 VTAIL.n53 VSUBS 0.021931f
C694 VTAIL.n54 VSUBS 0.021931f
C695 VTAIL.n55 VSUBS 0.011785f
C696 VTAIL.n56 VSUBS 0.012478f
C697 VTAIL.n57 VSUBS 0.027855f
C698 VTAIL.n58 VSUBS 0.070288f
C699 VTAIL.n59 VSUBS 0.012478f
C700 VTAIL.n60 VSUBS 0.011785f
C701 VTAIL.n61 VSUBS 0.053688f
C702 VTAIL.n62 VSUBS 0.035564f
C703 VTAIL.n63 VSUBS 1.22572f
C704 VTAIL.n64 VSUBS 0.024935f
C705 VTAIL.n65 VSUBS 0.021931f
C706 VTAIL.n66 VSUBS 0.011785f
C707 VTAIL.n67 VSUBS 0.027855f
C708 VTAIL.n68 VSUBS 0.012478f
C709 VTAIL.n69 VSUBS 0.021931f
C710 VTAIL.n70 VSUBS 0.011785f
C711 VTAIL.n71 VSUBS 0.027855f
C712 VTAIL.n72 VSUBS 0.012478f
C713 VTAIL.n73 VSUBS 0.097733f
C714 VTAIL.t1 VSUBS 0.059893f
C715 VTAIL.n74 VSUBS 0.020891f
C716 VTAIL.n75 VSUBS 0.017711f
C717 VTAIL.n76 VSUBS 0.011785f
C718 VTAIL.n77 VSUBS 0.512801f
C719 VTAIL.n78 VSUBS 0.021931f
C720 VTAIL.n79 VSUBS 0.011785f
C721 VTAIL.n80 VSUBS 0.012478f
C722 VTAIL.n81 VSUBS 0.027855f
C723 VTAIL.n82 VSUBS 0.027855f
C724 VTAIL.n83 VSUBS 0.012478f
C725 VTAIL.n84 VSUBS 0.011785f
C726 VTAIL.n85 VSUBS 0.021931f
C727 VTAIL.n86 VSUBS 0.021931f
C728 VTAIL.n87 VSUBS 0.011785f
C729 VTAIL.n88 VSUBS 0.012478f
C730 VTAIL.n89 VSUBS 0.027855f
C731 VTAIL.n90 VSUBS 0.070288f
C732 VTAIL.n91 VSUBS 0.012478f
C733 VTAIL.n92 VSUBS 0.011785f
C734 VTAIL.n93 VSUBS 0.053688f
C735 VTAIL.n94 VSUBS 0.035564f
C736 VTAIL.n95 VSUBS 1.02469f
C737 VTAIL.n96 VSUBS 0.024935f
C738 VTAIL.n97 VSUBS 0.021931f
C739 VTAIL.n98 VSUBS 0.011785f
C740 VTAIL.n99 VSUBS 0.027855f
C741 VTAIL.n100 VSUBS 0.012478f
C742 VTAIL.n101 VSUBS 0.021931f
C743 VTAIL.n102 VSUBS 0.011785f
C744 VTAIL.n103 VSUBS 0.027855f
C745 VTAIL.n104 VSUBS 0.012478f
C746 VTAIL.n105 VSUBS 0.097733f
C747 VTAIL.t3 VSUBS 0.059893f
C748 VTAIL.n106 VSUBS 0.020891f
C749 VTAIL.n107 VSUBS 0.017711f
C750 VTAIL.n108 VSUBS 0.011785f
C751 VTAIL.n109 VSUBS 0.512801f
C752 VTAIL.n110 VSUBS 0.021931f
C753 VTAIL.n111 VSUBS 0.011785f
C754 VTAIL.n112 VSUBS 0.012478f
C755 VTAIL.n113 VSUBS 0.027855f
C756 VTAIL.n114 VSUBS 0.027855f
C757 VTAIL.n115 VSUBS 0.012478f
C758 VTAIL.n116 VSUBS 0.011785f
C759 VTAIL.n117 VSUBS 0.021931f
C760 VTAIL.n118 VSUBS 0.021931f
C761 VTAIL.n119 VSUBS 0.011785f
C762 VTAIL.n120 VSUBS 0.012478f
C763 VTAIL.n121 VSUBS 0.027855f
C764 VTAIL.n122 VSUBS 0.070288f
C765 VTAIL.n123 VSUBS 0.012478f
C766 VTAIL.n124 VSUBS 0.011785f
C767 VTAIL.n125 VSUBS 0.053688f
C768 VTAIL.n126 VSUBS 0.035564f
C769 VTAIL.n127 VSUBS 0.937119f
C770 VN.t0 VSUBS 1.8865f
C771 VN.t1 VSUBS 2.4736f
.ends

