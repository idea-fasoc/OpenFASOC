* NGSPICE file created from diff_pair_sample_1042.ext - technology: sky130A

.subckt diff_pair_sample_1042 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t1 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=2.55585 pd=15.82 as=6.0411 ps=31.76 w=15.49 l=2.66
X1 VTAIL.t0 VN.t0 VDD2.t3 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=2.55585 ps=15.82 w=15.49 l=2.66
X2 B.t11 B.t9 B.t10 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=0 ps=0 w=15.49 l=2.66
X3 VTAIL.t5 VN.t1 VDD2.t2 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=2.55585 ps=15.82 w=15.49 l=2.66
X4 VTAIL.t3 VP.t1 VDD1.t2 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=2.55585 ps=15.82 w=15.49 l=2.66
X5 VDD2.t1 VN.t2 VTAIL.t7 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=2.55585 pd=15.82 as=6.0411 ps=31.76 w=15.49 l=2.66
X6 VDD2.t0 VN.t3 VTAIL.t6 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=2.55585 pd=15.82 as=6.0411 ps=31.76 w=15.49 l=2.66
X7 B.t8 B.t6 B.t7 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=0 ps=0 w=15.49 l=2.66
X8 B.t5 B.t3 B.t4 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=0 ps=0 w=15.49 l=2.66
X9 VDD1.t1 VP.t2 VTAIL.t2 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=2.55585 pd=15.82 as=6.0411 ps=31.76 w=15.49 l=2.66
X10 VTAIL.t4 VP.t3 VDD1.t0 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=2.55585 ps=15.82 w=15.49 l=2.66
X11 B.t2 B.t0 B.t1 w_n2764_n4066# sky130_fd_pr__pfet_01v8 ad=6.0411 pd=31.76 as=0 ps=0 w=15.49 l=2.66
R0 VP.n3 VP.t1 174.055
R1 VP.n3 VP.t0 173.195
R2 VP.n13 VP.n12 161.3
R3 VP.n11 VP.n1 161.3
R4 VP.n10 VP.n9 161.3
R5 VP.n8 VP.n2 161.3
R6 VP.n7 VP.n6 161.3
R7 VP.n5 VP.t3 140.343
R8 VP.n0 VP.t2 140.343
R9 VP.n5 VP.n4 65.8451
R10 VP.n14 VP.n0 65.8451
R11 VP.n4 VP.n3 52.8483
R12 VP.n10 VP.n2 40.4934
R13 VP.n11 VP.n10 40.4934
R14 VP.n6 VP.n2 24.4675
R15 VP.n12 VP.n11 24.4675
R16 VP.n6 VP.n5 24.2228
R17 VP.n12 VP.n0 24.2228
R18 VP.n7 VP.n4 0.354971
R19 VP.n14 VP.n13 0.354971
R20 VP VP.n14 0.26696
R21 VP.n8 VP.n7 0.189894
R22 VP.n9 VP.n8 0.189894
R23 VP.n9 VP.n1 0.189894
R24 VP.n13 VP.n1 0.189894
R25 VTAIL.n682 VTAIL.n602 756.745
R26 VTAIL.n80 VTAIL.n0 756.745
R27 VTAIL.n166 VTAIL.n86 756.745
R28 VTAIL.n252 VTAIL.n172 756.745
R29 VTAIL.n596 VTAIL.n516 756.745
R30 VTAIL.n510 VTAIL.n430 756.745
R31 VTAIL.n424 VTAIL.n344 756.745
R32 VTAIL.n338 VTAIL.n258 756.745
R33 VTAIL.n631 VTAIL.n630 585
R34 VTAIL.n633 VTAIL.n632 585
R35 VTAIL.n626 VTAIL.n625 585
R36 VTAIL.n639 VTAIL.n638 585
R37 VTAIL.n641 VTAIL.n640 585
R38 VTAIL.n622 VTAIL.n621 585
R39 VTAIL.n647 VTAIL.n646 585
R40 VTAIL.n649 VTAIL.n648 585
R41 VTAIL.n618 VTAIL.n617 585
R42 VTAIL.n655 VTAIL.n654 585
R43 VTAIL.n657 VTAIL.n656 585
R44 VTAIL.n614 VTAIL.n613 585
R45 VTAIL.n663 VTAIL.n662 585
R46 VTAIL.n665 VTAIL.n664 585
R47 VTAIL.n610 VTAIL.n609 585
R48 VTAIL.n672 VTAIL.n671 585
R49 VTAIL.n673 VTAIL.n608 585
R50 VTAIL.n675 VTAIL.n674 585
R51 VTAIL.n606 VTAIL.n605 585
R52 VTAIL.n681 VTAIL.n680 585
R53 VTAIL.n683 VTAIL.n682 585
R54 VTAIL.n29 VTAIL.n28 585
R55 VTAIL.n31 VTAIL.n30 585
R56 VTAIL.n24 VTAIL.n23 585
R57 VTAIL.n37 VTAIL.n36 585
R58 VTAIL.n39 VTAIL.n38 585
R59 VTAIL.n20 VTAIL.n19 585
R60 VTAIL.n45 VTAIL.n44 585
R61 VTAIL.n47 VTAIL.n46 585
R62 VTAIL.n16 VTAIL.n15 585
R63 VTAIL.n53 VTAIL.n52 585
R64 VTAIL.n55 VTAIL.n54 585
R65 VTAIL.n12 VTAIL.n11 585
R66 VTAIL.n61 VTAIL.n60 585
R67 VTAIL.n63 VTAIL.n62 585
R68 VTAIL.n8 VTAIL.n7 585
R69 VTAIL.n70 VTAIL.n69 585
R70 VTAIL.n71 VTAIL.n6 585
R71 VTAIL.n73 VTAIL.n72 585
R72 VTAIL.n4 VTAIL.n3 585
R73 VTAIL.n79 VTAIL.n78 585
R74 VTAIL.n81 VTAIL.n80 585
R75 VTAIL.n115 VTAIL.n114 585
R76 VTAIL.n117 VTAIL.n116 585
R77 VTAIL.n110 VTAIL.n109 585
R78 VTAIL.n123 VTAIL.n122 585
R79 VTAIL.n125 VTAIL.n124 585
R80 VTAIL.n106 VTAIL.n105 585
R81 VTAIL.n131 VTAIL.n130 585
R82 VTAIL.n133 VTAIL.n132 585
R83 VTAIL.n102 VTAIL.n101 585
R84 VTAIL.n139 VTAIL.n138 585
R85 VTAIL.n141 VTAIL.n140 585
R86 VTAIL.n98 VTAIL.n97 585
R87 VTAIL.n147 VTAIL.n146 585
R88 VTAIL.n149 VTAIL.n148 585
R89 VTAIL.n94 VTAIL.n93 585
R90 VTAIL.n156 VTAIL.n155 585
R91 VTAIL.n157 VTAIL.n92 585
R92 VTAIL.n159 VTAIL.n158 585
R93 VTAIL.n90 VTAIL.n89 585
R94 VTAIL.n165 VTAIL.n164 585
R95 VTAIL.n167 VTAIL.n166 585
R96 VTAIL.n201 VTAIL.n200 585
R97 VTAIL.n203 VTAIL.n202 585
R98 VTAIL.n196 VTAIL.n195 585
R99 VTAIL.n209 VTAIL.n208 585
R100 VTAIL.n211 VTAIL.n210 585
R101 VTAIL.n192 VTAIL.n191 585
R102 VTAIL.n217 VTAIL.n216 585
R103 VTAIL.n219 VTAIL.n218 585
R104 VTAIL.n188 VTAIL.n187 585
R105 VTAIL.n225 VTAIL.n224 585
R106 VTAIL.n227 VTAIL.n226 585
R107 VTAIL.n184 VTAIL.n183 585
R108 VTAIL.n233 VTAIL.n232 585
R109 VTAIL.n235 VTAIL.n234 585
R110 VTAIL.n180 VTAIL.n179 585
R111 VTAIL.n242 VTAIL.n241 585
R112 VTAIL.n243 VTAIL.n178 585
R113 VTAIL.n245 VTAIL.n244 585
R114 VTAIL.n176 VTAIL.n175 585
R115 VTAIL.n251 VTAIL.n250 585
R116 VTAIL.n253 VTAIL.n252 585
R117 VTAIL.n597 VTAIL.n596 585
R118 VTAIL.n595 VTAIL.n594 585
R119 VTAIL.n520 VTAIL.n519 585
R120 VTAIL.n524 VTAIL.n522 585
R121 VTAIL.n589 VTAIL.n588 585
R122 VTAIL.n587 VTAIL.n586 585
R123 VTAIL.n526 VTAIL.n525 585
R124 VTAIL.n581 VTAIL.n580 585
R125 VTAIL.n579 VTAIL.n578 585
R126 VTAIL.n530 VTAIL.n529 585
R127 VTAIL.n573 VTAIL.n572 585
R128 VTAIL.n571 VTAIL.n570 585
R129 VTAIL.n534 VTAIL.n533 585
R130 VTAIL.n565 VTAIL.n564 585
R131 VTAIL.n563 VTAIL.n562 585
R132 VTAIL.n538 VTAIL.n537 585
R133 VTAIL.n557 VTAIL.n556 585
R134 VTAIL.n555 VTAIL.n554 585
R135 VTAIL.n542 VTAIL.n541 585
R136 VTAIL.n549 VTAIL.n548 585
R137 VTAIL.n547 VTAIL.n546 585
R138 VTAIL.n511 VTAIL.n510 585
R139 VTAIL.n509 VTAIL.n508 585
R140 VTAIL.n434 VTAIL.n433 585
R141 VTAIL.n438 VTAIL.n436 585
R142 VTAIL.n503 VTAIL.n502 585
R143 VTAIL.n501 VTAIL.n500 585
R144 VTAIL.n440 VTAIL.n439 585
R145 VTAIL.n495 VTAIL.n494 585
R146 VTAIL.n493 VTAIL.n492 585
R147 VTAIL.n444 VTAIL.n443 585
R148 VTAIL.n487 VTAIL.n486 585
R149 VTAIL.n485 VTAIL.n484 585
R150 VTAIL.n448 VTAIL.n447 585
R151 VTAIL.n479 VTAIL.n478 585
R152 VTAIL.n477 VTAIL.n476 585
R153 VTAIL.n452 VTAIL.n451 585
R154 VTAIL.n471 VTAIL.n470 585
R155 VTAIL.n469 VTAIL.n468 585
R156 VTAIL.n456 VTAIL.n455 585
R157 VTAIL.n463 VTAIL.n462 585
R158 VTAIL.n461 VTAIL.n460 585
R159 VTAIL.n425 VTAIL.n424 585
R160 VTAIL.n423 VTAIL.n422 585
R161 VTAIL.n348 VTAIL.n347 585
R162 VTAIL.n352 VTAIL.n350 585
R163 VTAIL.n417 VTAIL.n416 585
R164 VTAIL.n415 VTAIL.n414 585
R165 VTAIL.n354 VTAIL.n353 585
R166 VTAIL.n409 VTAIL.n408 585
R167 VTAIL.n407 VTAIL.n406 585
R168 VTAIL.n358 VTAIL.n357 585
R169 VTAIL.n401 VTAIL.n400 585
R170 VTAIL.n399 VTAIL.n398 585
R171 VTAIL.n362 VTAIL.n361 585
R172 VTAIL.n393 VTAIL.n392 585
R173 VTAIL.n391 VTAIL.n390 585
R174 VTAIL.n366 VTAIL.n365 585
R175 VTAIL.n385 VTAIL.n384 585
R176 VTAIL.n383 VTAIL.n382 585
R177 VTAIL.n370 VTAIL.n369 585
R178 VTAIL.n377 VTAIL.n376 585
R179 VTAIL.n375 VTAIL.n374 585
R180 VTAIL.n339 VTAIL.n338 585
R181 VTAIL.n337 VTAIL.n336 585
R182 VTAIL.n262 VTAIL.n261 585
R183 VTAIL.n266 VTAIL.n264 585
R184 VTAIL.n331 VTAIL.n330 585
R185 VTAIL.n329 VTAIL.n328 585
R186 VTAIL.n268 VTAIL.n267 585
R187 VTAIL.n323 VTAIL.n322 585
R188 VTAIL.n321 VTAIL.n320 585
R189 VTAIL.n272 VTAIL.n271 585
R190 VTAIL.n315 VTAIL.n314 585
R191 VTAIL.n313 VTAIL.n312 585
R192 VTAIL.n276 VTAIL.n275 585
R193 VTAIL.n307 VTAIL.n306 585
R194 VTAIL.n305 VTAIL.n304 585
R195 VTAIL.n280 VTAIL.n279 585
R196 VTAIL.n299 VTAIL.n298 585
R197 VTAIL.n297 VTAIL.n296 585
R198 VTAIL.n284 VTAIL.n283 585
R199 VTAIL.n291 VTAIL.n290 585
R200 VTAIL.n289 VTAIL.n288 585
R201 VTAIL.n629 VTAIL.t6 327.466
R202 VTAIL.n27 VTAIL.t5 327.466
R203 VTAIL.n113 VTAIL.t2 327.466
R204 VTAIL.n199 VTAIL.t4 327.466
R205 VTAIL.n545 VTAIL.t1 327.466
R206 VTAIL.n459 VTAIL.t3 327.466
R207 VTAIL.n373 VTAIL.t7 327.466
R208 VTAIL.n287 VTAIL.t0 327.466
R209 VTAIL.n632 VTAIL.n631 171.744
R210 VTAIL.n632 VTAIL.n625 171.744
R211 VTAIL.n639 VTAIL.n625 171.744
R212 VTAIL.n640 VTAIL.n639 171.744
R213 VTAIL.n640 VTAIL.n621 171.744
R214 VTAIL.n647 VTAIL.n621 171.744
R215 VTAIL.n648 VTAIL.n647 171.744
R216 VTAIL.n648 VTAIL.n617 171.744
R217 VTAIL.n655 VTAIL.n617 171.744
R218 VTAIL.n656 VTAIL.n655 171.744
R219 VTAIL.n656 VTAIL.n613 171.744
R220 VTAIL.n663 VTAIL.n613 171.744
R221 VTAIL.n664 VTAIL.n663 171.744
R222 VTAIL.n664 VTAIL.n609 171.744
R223 VTAIL.n672 VTAIL.n609 171.744
R224 VTAIL.n673 VTAIL.n672 171.744
R225 VTAIL.n674 VTAIL.n673 171.744
R226 VTAIL.n674 VTAIL.n605 171.744
R227 VTAIL.n681 VTAIL.n605 171.744
R228 VTAIL.n682 VTAIL.n681 171.744
R229 VTAIL.n30 VTAIL.n29 171.744
R230 VTAIL.n30 VTAIL.n23 171.744
R231 VTAIL.n37 VTAIL.n23 171.744
R232 VTAIL.n38 VTAIL.n37 171.744
R233 VTAIL.n38 VTAIL.n19 171.744
R234 VTAIL.n45 VTAIL.n19 171.744
R235 VTAIL.n46 VTAIL.n45 171.744
R236 VTAIL.n46 VTAIL.n15 171.744
R237 VTAIL.n53 VTAIL.n15 171.744
R238 VTAIL.n54 VTAIL.n53 171.744
R239 VTAIL.n54 VTAIL.n11 171.744
R240 VTAIL.n61 VTAIL.n11 171.744
R241 VTAIL.n62 VTAIL.n61 171.744
R242 VTAIL.n62 VTAIL.n7 171.744
R243 VTAIL.n70 VTAIL.n7 171.744
R244 VTAIL.n71 VTAIL.n70 171.744
R245 VTAIL.n72 VTAIL.n71 171.744
R246 VTAIL.n72 VTAIL.n3 171.744
R247 VTAIL.n79 VTAIL.n3 171.744
R248 VTAIL.n80 VTAIL.n79 171.744
R249 VTAIL.n116 VTAIL.n115 171.744
R250 VTAIL.n116 VTAIL.n109 171.744
R251 VTAIL.n123 VTAIL.n109 171.744
R252 VTAIL.n124 VTAIL.n123 171.744
R253 VTAIL.n124 VTAIL.n105 171.744
R254 VTAIL.n131 VTAIL.n105 171.744
R255 VTAIL.n132 VTAIL.n131 171.744
R256 VTAIL.n132 VTAIL.n101 171.744
R257 VTAIL.n139 VTAIL.n101 171.744
R258 VTAIL.n140 VTAIL.n139 171.744
R259 VTAIL.n140 VTAIL.n97 171.744
R260 VTAIL.n147 VTAIL.n97 171.744
R261 VTAIL.n148 VTAIL.n147 171.744
R262 VTAIL.n148 VTAIL.n93 171.744
R263 VTAIL.n156 VTAIL.n93 171.744
R264 VTAIL.n157 VTAIL.n156 171.744
R265 VTAIL.n158 VTAIL.n157 171.744
R266 VTAIL.n158 VTAIL.n89 171.744
R267 VTAIL.n165 VTAIL.n89 171.744
R268 VTAIL.n166 VTAIL.n165 171.744
R269 VTAIL.n202 VTAIL.n201 171.744
R270 VTAIL.n202 VTAIL.n195 171.744
R271 VTAIL.n209 VTAIL.n195 171.744
R272 VTAIL.n210 VTAIL.n209 171.744
R273 VTAIL.n210 VTAIL.n191 171.744
R274 VTAIL.n217 VTAIL.n191 171.744
R275 VTAIL.n218 VTAIL.n217 171.744
R276 VTAIL.n218 VTAIL.n187 171.744
R277 VTAIL.n225 VTAIL.n187 171.744
R278 VTAIL.n226 VTAIL.n225 171.744
R279 VTAIL.n226 VTAIL.n183 171.744
R280 VTAIL.n233 VTAIL.n183 171.744
R281 VTAIL.n234 VTAIL.n233 171.744
R282 VTAIL.n234 VTAIL.n179 171.744
R283 VTAIL.n242 VTAIL.n179 171.744
R284 VTAIL.n243 VTAIL.n242 171.744
R285 VTAIL.n244 VTAIL.n243 171.744
R286 VTAIL.n244 VTAIL.n175 171.744
R287 VTAIL.n251 VTAIL.n175 171.744
R288 VTAIL.n252 VTAIL.n251 171.744
R289 VTAIL.n596 VTAIL.n595 171.744
R290 VTAIL.n595 VTAIL.n519 171.744
R291 VTAIL.n524 VTAIL.n519 171.744
R292 VTAIL.n588 VTAIL.n524 171.744
R293 VTAIL.n588 VTAIL.n587 171.744
R294 VTAIL.n587 VTAIL.n525 171.744
R295 VTAIL.n580 VTAIL.n525 171.744
R296 VTAIL.n580 VTAIL.n579 171.744
R297 VTAIL.n579 VTAIL.n529 171.744
R298 VTAIL.n572 VTAIL.n529 171.744
R299 VTAIL.n572 VTAIL.n571 171.744
R300 VTAIL.n571 VTAIL.n533 171.744
R301 VTAIL.n564 VTAIL.n533 171.744
R302 VTAIL.n564 VTAIL.n563 171.744
R303 VTAIL.n563 VTAIL.n537 171.744
R304 VTAIL.n556 VTAIL.n537 171.744
R305 VTAIL.n556 VTAIL.n555 171.744
R306 VTAIL.n555 VTAIL.n541 171.744
R307 VTAIL.n548 VTAIL.n541 171.744
R308 VTAIL.n548 VTAIL.n547 171.744
R309 VTAIL.n510 VTAIL.n509 171.744
R310 VTAIL.n509 VTAIL.n433 171.744
R311 VTAIL.n438 VTAIL.n433 171.744
R312 VTAIL.n502 VTAIL.n438 171.744
R313 VTAIL.n502 VTAIL.n501 171.744
R314 VTAIL.n501 VTAIL.n439 171.744
R315 VTAIL.n494 VTAIL.n439 171.744
R316 VTAIL.n494 VTAIL.n493 171.744
R317 VTAIL.n493 VTAIL.n443 171.744
R318 VTAIL.n486 VTAIL.n443 171.744
R319 VTAIL.n486 VTAIL.n485 171.744
R320 VTAIL.n485 VTAIL.n447 171.744
R321 VTAIL.n478 VTAIL.n447 171.744
R322 VTAIL.n478 VTAIL.n477 171.744
R323 VTAIL.n477 VTAIL.n451 171.744
R324 VTAIL.n470 VTAIL.n451 171.744
R325 VTAIL.n470 VTAIL.n469 171.744
R326 VTAIL.n469 VTAIL.n455 171.744
R327 VTAIL.n462 VTAIL.n455 171.744
R328 VTAIL.n462 VTAIL.n461 171.744
R329 VTAIL.n424 VTAIL.n423 171.744
R330 VTAIL.n423 VTAIL.n347 171.744
R331 VTAIL.n352 VTAIL.n347 171.744
R332 VTAIL.n416 VTAIL.n352 171.744
R333 VTAIL.n416 VTAIL.n415 171.744
R334 VTAIL.n415 VTAIL.n353 171.744
R335 VTAIL.n408 VTAIL.n353 171.744
R336 VTAIL.n408 VTAIL.n407 171.744
R337 VTAIL.n407 VTAIL.n357 171.744
R338 VTAIL.n400 VTAIL.n357 171.744
R339 VTAIL.n400 VTAIL.n399 171.744
R340 VTAIL.n399 VTAIL.n361 171.744
R341 VTAIL.n392 VTAIL.n361 171.744
R342 VTAIL.n392 VTAIL.n391 171.744
R343 VTAIL.n391 VTAIL.n365 171.744
R344 VTAIL.n384 VTAIL.n365 171.744
R345 VTAIL.n384 VTAIL.n383 171.744
R346 VTAIL.n383 VTAIL.n369 171.744
R347 VTAIL.n376 VTAIL.n369 171.744
R348 VTAIL.n376 VTAIL.n375 171.744
R349 VTAIL.n338 VTAIL.n337 171.744
R350 VTAIL.n337 VTAIL.n261 171.744
R351 VTAIL.n266 VTAIL.n261 171.744
R352 VTAIL.n330 VTAIL.n266 171.744
R353 VTAIL.n330 VTAIL.n329 171.744
R354 VTAIL.n329 VTAIL.n267 171.744
R355 VTAIL.n322 VTAIL.n267 171.744
R356 VTAIL.n322 VTAIL.n321 171.744
R357 VTAIL.n321 VTAIL.n271 171.744
R358 VTAIL.n314 VTAIL.n271 171.744
R359 VTAIL.n314 VTAIL.n313 171.744
R360 VTAIL.n313 VTAIL.n275 171.744
R361 VTAIL.n306 VTAIL.n275 171.744
R362 VTAIL.n306 VTAIL.n305 171.744
R363 VTAIL.n305 VTAIL.n279 171.744
R364 VTAIL.n298 VTAIL.n279 171.744
R365 VTAIL.n298 VTAIL.n297 171.744
R366 VTAIL.n297 VTAIL.n283 171.744
R367 VTAIL.n290 VTAIL.n283 171.744
R368 VTAIL.n290 VTAIL.n289 171.744
R369 VTAIL.n631 VTAIL.t6 85.8723
R370 VTAIL.n29 VTAIL.t5 85.8723
R371 VTAIL.n115 VTAIL.t2 85.8723
R372 VTAIL.n201 VTAIL.t4 85.8723
R373 VTAIL.n547 VTAIL.t1 85.8723
R374 VTAIL.n461 VTAIL.t3 85.8723
R375 VTAIL.n375 VTAIL.t7 85.8723
R376 VTAIL.n289 VTAIL.t0 85.8723
R377 VTAIL.n687 VTAIL.n686 34.7066
R378 VTAIL.n85 VTAIL.n84 34.7066
R379 VTAIL.n171 VTAIL.n170 34.7066
R380 VTAIL.n257 VTAIL.n256 34.7066
R381 VTAIL.n601 VTAIL.n600 34.7066
R382 VTAIL.n515 VTAIL.n514 34.7066
R383 VTAIL.n429 VTAIL.n428 34.7066
R384 VTAIL.n343 VTAIL.n342 34.7066
R385 VTAIL.n687 VTAIL.n601 28.2979
R386 VTAIL.n343 VTAIL.n257 28.2979
R387 VTAIL.n630 VTAIL.n629 16.3895
R388 VTAIL.n28 VTAIL.n27 16.3895
R389 VTAIL.n114 VTAIL.n113 16.3895
R390 VTAIL.n200 VTAIL.n199 16.3895
R391 VTAIL.n546 VTAIL.n545 16.3895
R392 VTAIL.n460 VTAIL.n459 16.3895
R393 VTAIL.n374 VTAIL.n373 16.3895
R394 VTAIL.n288 VTAIL.n287 16.3895
R395 VTAIL.n675 VTAIL.n606 13.1884
R396 VTAIL.n73 VTAIL.n4 13.1884
R397 VTAIL.n159 VTAIL.n90 13.1884
R398 VTAIL.n245 VTAIL.n176 13.1884
R399 VTAIL.n522 VTAIL.n520 13.1884
R400 VTAIL.n436 VTAIL.n434 13.1884
R401 VTAIL.n350 VTAIL.n348 13.1884
R402 VTAIL.n264 VTAIL.n262 13.1884
R403 VTAIL.n633 VTAIL.n628 12.8005
R404 VTAIL.n676 VTAIL.n608 12.8005
R405 VTAIL.n680 VTAIL.n679 12.8005
R406 VTAIL.n31 VTAIL.n26 12.8005
R407 VTAIL.n74 VTAIL.n6 12.8005
R408 VTAIL.n78 VTAIL.n77 12.8005
R409 VTAIL.n117 VTAIL.n112 12.8005
R410 VTAIL.n160 VTAIL.n92 12.8005
R411 VTAIL.n164 VTAIL.n163 12.8005
R412 VTAIL.n203 VTAIL.n198 12.8005
R413 VTAIL.n246 VTAIL.n178 12.8005
R414 VTAIL.n250 VTAIL.n249 12.8005
R415 VTAIL.n594 VTAIL.n593 12.8005
R416 VTAIL.n590 VTAIL.n589 12.8005
R417 VTAIL.n549 VTAIL.n544 12.8005
R418 VTAIL.n508 VTAIL.n507 12.8005
R419 VTAIL.n504 VTAIL.n503 12.8005
R420 VTAIL.n463 VTAIL.n458 12.8005
R421 VTAIL.n422 VTAIL.n421 12.8005
R422 VTAIL.n418 VTAIL.n417 12.8005
R423 VTAIL.n377 VTAIL.n372 12.8005
R424 VTAIL.n336 VTAIL.n335 12.8005
R425 VTAIL.n332 VTAIL.n331 12.8005
R426 VTAIL.n291 VTAIL.n286 12.8005
R427 VTAIL.n634 VTAIL.n626 12.0247
R428 VTAIL.n671 VTAIL.n670 12.0247
R429 VTAIL.n683 VTAIL.n604 12.0247
R430 VTAIL.n32 VTAIL.n24 12.0247
R431 VTAIL.n69 VTAIL.n68 12.0247
R432 VTAIL.n81 VTAIL.n2 12.0247
R433 VTAIL.n118 VTAIL.n110 12.0247
R434 VTAIL.n155 VTAIL.n154 12.0247
R435 VTAIL.n167 VTAIL.n88 12.0247
R436 VTAIL.n204 VTAIL.n196 12.0247
R437 VTAIL.n241 VTAIL.n240 12.0247
R438 VTAIL.n253 VTAIL.n174 12.0247
R439 VTAIL.n597 VTAIL.n518 12.0247
R440 VTAIL.n586 VTAIL.n523 12.0247
R441 VTAIL.n550 VTAIL.n542 12.0247
R442 VTAIL.n511 VTAIL.n432 12.0247
R443 VTAIL.n500 VTAIL.n437 12.0247
R444 VTAIL.n464 VTAIL.n456 12.0247
R445 VTAIL.n425 VTAIL.n346 12.0247
R446 VTAIL.n414 VTAIL.n351 12.0247
R447 VTAIL.n378 VTAIL.n370 12.0247
R448 VTAIL.n339 VTAIL.n260 12.0247
R449 VTAIL.n328 VTAIL.n265 12.0247
R450 VTAIL.n292 VTAIL.n284 12.0247
R451 VTAIL.n638 VTAIL.n637 11.249
R452 VTAIL.n669 VTAIL.n610 11.249
R453 VTAIL.n684 VTAIL.n602 11.249
R454 VTAIL.n36 VTAIL.n35 11.249
R455 VTAIL.n67 VTAIL.n8 11.249
R456 VTAIL.n82 VTAIL.n0 11.249
R457 VTAIL.n122 VTAIL.n121 11.249
R458 VTAIL.n153 VTAIL.n94 11.249
R459 VTAIL.n168 VTAIL.n86 11.249
R460 VTAIL.n208 VTAIL.n207 11.249
R461 VTAIL.n239 VTAIL.n180 11.249
R462 VTAIL.n254 VTAIL.n172 11.249
R463 VTAIL.n598 VTAIL.n516 11.249
R464 VTAIL.n585 VTAIL.n526 11.249
R465 VTAIL.n554 VTAIL.n553 11.249
R466 VTAIL.n512 VTAIL.n430 11.249
R467 VTAIL.n499 VTAIL.n440 11.249
R468 VTAIL.n468 VTAIL.n467 11.249
R469 VTAIL.n426 VTAIL.n344 11.249
R470 VTAIL.n413 VTAIL.n354 11.249
R471 VTAIL.n382 VTAIL.n381 11.249
R472 VTAIL.n340 VTAIL.n258 11.249
R473 VTAIL.n327 VTAIL.n268 11.249
R474 VTAIL.n296 VTAIL.n295 11.249
R475 VTAIL.n641 VTAIL.n624 10.4732
R476 VTAIL.n666 VTAIL.n665 10.4732
R477 VTAIL.n39 VTAIL.n22 10.4732
R478 VTAIL.n64 VTAIL.n63 10.4732
R479 VTAIL.n125 VTAIL.n108 10.4732
R480 VTAIL.n150 VTAIL.n149 10.4732
R481 VTAIL.n211 VTAIL.n194 10.4732
R482 VTAIL.n236 VTAIL.n235 10.4732
R483 VTAIL.n582 VTAIL.n581 10.4732
R484 VTAIL.n557 VTAIL.n540 10.4732
R485 VTAIL.n496 VTAIL.n495 10.4732
R486 VTAIL.n471 VTAIL.n454 10.4732
R487 VTAIL.n410 VTAIL.n409 10.4732
R488 VTAIL.n385 VTAIL.n368 10.4732
R489 VTAIL.n324 VTAIL.n323 10.4732
R490 VTAIL.n299 VTAIL.n282 10.4732
R491 VTAIL.n642 VTAIL.n622 9.69747
R492 VTAIL.n662 VTAIL.n612 9.69747
R493 VTAIL.n40 VTAIL.n20 9.69747
R494 VTAIL.n60 VTAIL.n10 9.69747
R495 VTAIL.n126 VTAIL.n106 9.69747
R496 VTAIL.n146 VTAIL.n96 9.69747
R497 VTAIL.n212 VTAIL.n192 9.69747
R498 VTAIL.n232 VTAIL.n182 9.69747
R499 VTAIL.n578 VTAIL.n528 9.69747
R500 VTAIL.n558 VTAIL.n538 9.69747
R501 VTAIL.n492 VTAIL.n442 9.69747
R502 VTAIL.n472 VTAIL.n452 9.69747
R503 VTAIL.n406 VTAIL.n356 9.69747
R504 VTAIL.n386 VTAIL.n366 9.69747
R505 VTAIL.n320 VTAIL.n270 9.69747
R506 VTAIL.n300 VTAIL.n280 9.69747
R507 VTAIL.n686 VTAIL.n685 9.45567
R508 VTAIL.n84 VTAIL.n83 9.45567
R509 VTAIL.n170 VTAIL.n169 9.45567
R510 VTAIL.n256 VTAIL.n255 9.45567
R511 VTAIL.n600 VTAIL.n599 9.45567
R512 VTAIL.n514 VTAIL.n513 9.45567
R513 VTAIL.n428 VTAIL.n427 9.45567
R514 VTAIL.n342 VTAIL.n341 9.45567
R515 VTAIL.n685 VTAIL.n684 9.3005
R516 VTAIL.n604 VTAIL.n603 9.3005
R517 VTAIL.n679 VTAIL.n678 9.3005
R518 VTAIL.n651 VTAIL.n650 9.3005
R519 VTAIL.n620 VTAIL.n619 9.3005
R520 VTAIL.n645 VTAIL.n644 9.3005
R521 VTAIL.n643 VTAIL.n642 9.3005
R522 VTAIL.n624 VTAIL.n623 9.3005
R523 VTAIL.n637 VTAIL.n636 9.3005
R524 VTAIL.n635 VTAIL.n634 9.3005
R525 VTAIL.n628 VTAIL.n627 9.3005
R526 VTAIL.n653 VTAIL.n652 9.3005
R527 VTAIL.n616 VTAIL.n615 9.3005
R528 VTAIL.n659 VTAIL.n658 9.3005
R529 VTAIL.n661 VTAIL.n660 9.3005
R530 VTAIL.n612 VTAIL.n611 9.3005
R531 VTAIL.n667 VTAIL.n666 9.3005
R532 VTAIL.n669 VTAIL.n668 9.3005
R533 VTAIL.n670 VTAIL.n607 9.3005
R534 VTAIL.n677 VTAIL.n676 9.3005
R535 VTAIL.n83 VTAIL.n82 9.3005
R536 VTAIL.n2 VTAIL.n1 9.3005
R537 VTAIL.n77 VTAIL.n76 9.3005
R538 VTAIL.n49 VTAIL.n48 9.3005
R539 VTAIL.n18 VTAIL.n17 9.3005
R540 VTAIL.n43 VTAIL.n42 9.3005
R541 VTAIL.n41 VTAIL.n40 9.3005
R542 VTAIL.n22 VTAIL.n21 9.3005
R543 VTAIL.n35 VTAIL.n34 9.3005
R544 VTAIL.n33 VTAIL.n32 9.3005
R545 VTAIL.n26 VTAIL.n25 9.3005
R546 VTAIL.n51 VTAIL.n50 9.3005
R547 VTAIL.n14 VTAIL.n13 9.3005
R548 VTAIL.n57 VTAIL.n56 9.3005
R549 VTAIL.n59 VTAIL.n58 9.3005
R550 VTAIL.n10 VTAIL.n9 9.3005
R551 VTAIL.n65 VTAIL.n64 9.3005
R552 VTAIL.n67 VTAIL.n66 9.3005
R553 VTAIL.n68 VTAIL.n5 9.3005
R554 VTAIL.n75 VTAIL.n74 9.3005
R555 VTAIL.n169 VTAIL.n168 9.3005
R556 VTAIL.n88 VTAIL.n87 9.3005
R557 VTAIL.n163 VTAIL.n162 9.3005
R558 VTAIL.n135 VTAIL.n134 9.3005
R559 VTAIL.n104 VTAIL.n103 9.3005
R560 VTAIL.n129 VTAIL.n128 9.3005
R561 VTAIL.n127 VTAIL.n126 9.3005
R562 VTAIL.n108 VTAIL.n107 9.3005
R563 VTAIL.n121 VTAIL.n120 9.3005
R564 VTAIL.n119 VTAIL.n118 9.3005
R565 VTAIL.n112 VTAIL.n111 9.3005
R566 VTAIL.n137 VTAIL.n136 9.3005
R567 VTAIL.n100 VTAIL.n99 9.3005
R568 VTAIL.n143 VTAIL.n142 9.3005
R569 VTAIL.n145 VTAIL.n144 9.3005
R570 VTAIL.n96 VTAIL.n95 9.3005
R571 VTAIL.n151 VTAIL.n150 9.3005
R572 VTAIL.n153 VTAIL.n152 9.3005
R573 VTAIL.n154 VTAIL.n91 9.3005
R574 VTAIL.n161 VTAIL.n160 9.3005
R575 VTAIL.n255 VTAIL.n254 9.3005
R576 VTAIL.n174 VTAIL.n173 9.3005
R577 VTAIL.n249 VTAIL.n248 9.3005
R578 VTAIL.n221 VTAIL.n220 9.3005
R579 VTAIL.n190 VTAIL.n189 9.3005
R580 VTAIL.n215 VTAIL.n214 9.3005
R581 VTAIL.n213 VTAIL.n212 9.3005
R582 VTAIL.n194 VTAIL.n193 9.3005
R583 VTAIL.n207 VTAIL.n206 9.3005
R584 VTAIL.n205 VTAIL.n204 9.3005
R585 VTAIL.n198 VTAIL.n197 9.3005
R586 VTAIL.n223 VTAIL.n222 9.3005
R587 VTAIL.n186 VTAIL.n185 9.3005
R588 VTAIL.n229 VTAIL.n228 9.3005
R589 VTAIL.n231 VTAIL.n230 9.3005
R590 VTAIL.n182 VTAIL.n181 9.3005
R591 VTAIL.n237 VTAIL.n236 9.3005
R592 VTAIL.n239 VTAIL.n238 9.3005
R593 VTAIL.n240 VTAIL.n177 9.3005
R594 VTAIL.n247 VTAIL.n246 9.3005
R595 VTAIL.n532 VTAIL.n531 9.3005
R596 VTAIL.n575 VTAIL.n574 9.3005
R597 VTAIL.n577 VTAIL.n576 9.3005
R598 VTAIL.n528 VTAIL.n527 9.3005
R599 VTAIL.n583 VTAIL.n582 9.3005
R600 VTAIL.n585 VTAIL.n584 9.3005
R601 VTAIL.n523 VTAIL.n521 9.3005
R602 VTAIL.n591 VTAIL.n590 9.3005
R603 VTAIL.n599 VTAIL.n598 9.3005
R604 VTAIL.n518 VTAIL.n517 9.3005
R605 VTAIL.n593 VTAIL.n592 9.3005
R606 VTAIL.n569 VTAIL.n568 9.3005
R607 VTAIL.n567 VTAIL.n566 9.3005
R608 VTAIL.n536 VTAIL.n535 9.3005
R609 VTAIL.n561 VTAIL.n560 9.3005
R610 VTAIL.n559 VTAIL.n558 9.3005
R611 VTAIL.n540 VTAIL.n539 9.3005
R612 VTAIL.n553 VTAIL.n552 9.3005
R613 VTAIL.n551 VTAIL.n550 9.3005
R614 VTAIL.n544 VTAIL.n543 9.3005
R615 VTAIL.n446 VTAIL.n445 9.3005
R616 VTAIL.n489 VTAIL.n488 9.3005
R617 VTAIL.n491 VTAIL.n490 9.3005
R618 VTAIL.n442 VTAIL.n441 9.3005
R619 VTAIL.n497 VTAIL.n496 9.3005
R620 VTAIL.n499 VTAIL.n498 9.3005
R621 VTAIL.n437 VTAIL.n435 9.3005
R622 VTAIL.n505 VTAIL.n504 9.3005
R623 VTAIL.n513 VTAIL.n512 9.3005
R624 VTAIL.n432 VTAIL.n431 9.3005
R625 VTAIL.n507 VTAIL.n506 9.3005
R626 VTAIL.n483 VTAIL.n482 9.3005
R627 VTAIL.n481 VTAIL.n480 9.3005
R628 VTAIL.n450 VTAIL.n449 9.3005
R629 VTAIL.n475 VTAIL.n474 9.3005
R630 VTAIL.n473 VTAIL.n472 9.3005
R631 VTAIL.n454 VTAIL.n453 9.3005
R632 VTAIL.n467 VTAIL.n466 9.3005
R633 VTAIL.n465 VTAIL.n464 9.3005
R634 VTAIL.n458 VTAIL.n457 9.3005
R635 VTAIL.n360 VTAIL.n359 9.3005
R636 VTAIL.n403 VTAIL.n402 9.3005
R637 VTAIL.n405 VTAIL.n404 9.3005
R638 VTAIL.n356 VTAIL.n355 9.3005
R639 VTAIL.n411 VTAIL.n410 9.3005
R640 VTAIL.n413 VTAIL.n412 9.3005
R641 VTAIL.n351 VTAIL.n349 9.3005
R642 VTAIL.n419 VTAIL.n418 9.3005
R643 VTAIL.n427 VTAIL.n426 9.3005
R644 VTAIL.n346 VTAIL.n345 9.3005
R645 VTAIL.n421 VTAIL.n420 9.3005
R646 VTAIL.n397 VTAIL.n396 9.3005
R647 VTAIL.n395 VTAIL.n394 9.3005
R648 VTAIL.n364 VTAIL.n363 9.3005
R649 VTAIL.n389 VTAIL.n388 9.3005
R650 VTAIL.n387 VTAIL.n386 9.3005
R651 VTAIL.n368 VTAIL.n367 9.3005
R652 VTAIL.n381 VTAIL.n380 9.3005
R653 VTAIL.n379 VTAIL.n378 9.3005
R654 VTAIL.n372 VTAIL.n371 9.3005
R655 VTAIL.n274 VTAIL.n273 9.3005
R656 VTAIL.n317 VTAIL.n316 9.3005
R657 VTAIL.n319 VTAIL.n318 9.3005
R658 VTAIL.n270 VTAIL.n269 9.3005
R659 VTAIL.n325 VTAIL.n324 9.3005
R660 VTAIL.n327 VTAIL.n326 9.3005
R661 VTAIL.n265 VTAIL.n263 9.3005
R662 VTAIL.n333 VTAIL.n332 9.3005
R663 VTAIL.n341 VTAIL.n340 9.3005
R664 VTAIL.n260 VTAIL.n259 9.3005
R665 VTAIL.n335 VTAIL.n334 9.3005
R666 VTAIL.n311 VTAIL.n310 9.3005
R667 VTAIL.n309 VTAIL.n308 9.3005
R668 VTAIL.n278 VTAIL.n277 9.3005
R669 VTAIL.n303 VTAIL.n302 9.3005
R670 VTAIL.n301 VTAIL.n300 9.3005
R671 VTAIL.n282 VTAIL.n281 9.3005
R672 VTAIL.n295 VTAIL.n294 9.3005
R673 VTAIL.n293 VTAIL.n292 9.3005
R674 VTAIL.n286 VTAIL.n285 9.3005
R675 VTAIL.n646 VTAIL.n645 8.92171
R676 VTAIL.n661 VTAIL.n614 8.92171
R677 VTAIL.n44 VTAIL.n43 8.92171
R678 VTAIL.n59 VTAIL.n12 8.92171
R679 VTAIL.n130 VTAIL.n129 8.92171
R680 VTAIL.n145 VTAIL.n98 8.92171
R681 VTAIL.n216 VTAIL.n215 8.92171
R682 VTAIL.n231 VTAIL.n184 8.92171
R683 VTAIL.n577 VTAIL.n530 8.92171
R684 VTAIL.n562 VTAIL.n561 8.92171
R685 VTAIL.n491 VTAIL.n444 8.92171
R686 VTAIL.n476 VTAIL.n475 8.92171
R687 VTAIL.n405 VTAIL.n358 8.92171
R688 VTAIL.n390 VTAIL.n389 8.92171
R689 VTAIL.n319 VTAIL.n272 8.92171
R690 VTAIL.n304 VTAIL.n303 8.92171
R691 VTAIL.n649 VTAIL.n620 8.14595
R692 VTAIL.n658 VTAIL.n657 8.14595
R693 VTAIL.n47 VTAIL.n18 8.14595
R694 VTAIL.n56 VTAIL.n55 8.14595
R695 VTAIL.n133 VTAIL.n104 8.14595
R696 VTAIL.n142 VTAIL.n141 8.14595
R697 VTAIL.n219 VTAIL.n190 8.14595
R698 VTAIL.n228 VTAIL.n227 8.14595
R699 VTAIL.n574 VTAIL.n573 8.14595
R700 VTAIL.n565 VTAIL.n536 8.14595
R701 VTAIL.n488 VTAIL.n487 8.14595
R702 VTAIL.n479 VTAIL.n450 8.14595
R703 VTAIL.n402 VTAIL.n401 8.14595
R704 VTAIL.n393 VTAIL.n364 8.14595
R705 VTAIL.n316 VTAIL.n315 8.14595
R706 VTAIL.n307 VTAIL.n278 8.14595
R707 VTAIL.n650 VTAIL.n618 7.3702
R708 VTAIL.n654 VTAIL.n616 7.3702
R709 VTAIL.n48 VTAIL.n16 7.3702
R710 VTAIL.n52 VTAIL.n14 7.3702
R711 VTAIL.n134 VTAIL.n102 7.3702
R712 VTAIL.n138 VTAIL.n100 7.3702
R713 VTAIL.n220 VTAIL.n188 7.3702
R714 VTAIL.n224 VTAIL.n186 7.3702
R715 VTAIL.n570 VTAIL.n532 7.3702
R716 VTAIL.n566 VTAIL.n534 7.3702
R717 VTAIL.n484 VTAIL.n446 7.3702
R718 VTAIL.n480 VTAIL.n448 7.3702
R719 VTAIL.n398 VTAIL.n360 7.3702
R720 VTAIL.n394 VTAIL.n362 7.3702
R721 VTAIL.n312 VTAIL.n274 7.3702
R722 VTAIL.n308 VTAIL.n276 7.3702
R723 VTAIL.n653 VTAIL.n618 6.59444
R724 VTAIL.n654 VTAIL.n653 6.59444
R725 VTAIL.n51 VTAIL.n16 6.59444
R726 VTAIL.n52 VTAIL.n51 6.59444
R727 VTAIL.n137 VTAIL.n102 6.59444
R728 VTAIL.n138 VTAIL.n137 6.59444
R729 VTAIL.n223 VTAIL.n188 6.59444
R730 VTAIL.n224 VTAIL.n223 6.59444
R731 VTAIL.n570 VTAIL.n569 6.59444
R732 VTAIL.n569 VTAIL.n534 6.59444
R733 VTAIL.n484 VTAIL.n483 6.59444
R734 VTAIL.n483 VTAIL.n448 6.59444
R735 VTAIL.n398 VTAIL.n397 6.59444
R736 VTAIL.n397 VTAIL.n362 6.59444
R737 VTAIL.n312 VTAIL.n311 6.59444
R738 VTAIL.n311 VTAIL.n276 6.59444
R739 VTAIL.n650 VTAIL.n649 5.81868
R740 VTAIL.n657 VTAIL.n616 5.81868
R741 VTAIL.n48 VTAIL.n47 5.81868
R742 VTAIL.n55 VTAIL.n14 5.81868
R743 VTAIL.n134 VTAIL.n133 5.81868
R744 VTAIL.n141 VTAIL.n100 5.81868
R745 VTAIL.n220 VTAIL.n219 5.81868
R746 VTAIL.n227 VTAIL.n186 5.81868
R747 VTAIL.n573 VTAIL.n532 5.81868
R748 VTAIL.n566 VTAIL.n565 5.81868
R749 VTAIL.n487 VTAIL.n446 5.81868
R750 VTAIL.n480 VTAIL.n479 5.81868
R751 VTAIL.n401 VTAIL.n360 5.81868
R752 VTAIL.n394 VTAIL.n393 5.81868
R753 VTAIL.n315 VTAIL.n274 5.81868
R754 VTAIL.n308 VTAIL.n307 5.81868
R755 VTAIL.n646 VTAIL.n620 5.04292
R756 VTAIL.n658 VTAIL.n614 5.04292
R757 VTAIL.n44 VTAIL.n18 5.04292
R758 VTAIL.n56 VTAIL.n12 5.04292
R759 VTAIL.n130 VTAIL.n104 5.04292
R760 VTAIL.n142 VTAIL.n98 5.04292
R761 VTAIL.n216 VTAIL.n190 5.04292
R762 VTAIL.n228 VTAIL.n184 5.04292
R763 VTAIL.n574 VTAIL.n530 5.04292
R764 VTAIL.n562 VTAIL.n536 5.04292
R765 VTAIL.n488 VTAIL.n444 5.04292
R766 VTAIL.n476 VTAIL.n450 5.04292
R767 VTAIL.n402 VTAIL.n358 5.04292
R768 VTAIL.n390 VTAIL.n364 5.04292
R769 VTAIL.n316 VTAIL.n272 5.04292
R770 VTAIL.n304 VTAIL.n278 5.04292
R771 VTAIL.n645 VTAIL.n622 4.26717
R772 VTAIL.n662 VTAIL.n661 4.26717
R773 VTAIL.n43 VTAIL.n20 4.26717
R774 VTAIL.n60 VTAIL.n59 4.26717
R775 VTAIL.n129 VTAIL.n106 4.26717
R776 VTAIL.n146 VTAIL.n145 4.26717
R777 VTAIL.n215 VTAIL.n192 4.26717
R778 VTAIL.n232 VTAIL.n231 4.26717
R779 VTAIL.n578 VTAIL.n577 4.26717
R780 VTAIL.n561 VTAIL.n538 4.26717
R781 VTAIL.n492 VTAIL.n491 4.26717
R782 VTAIL.n475 VTAIL.n452 4.26717
R783 VTAIL.n406 VTAIL.n405 4.26717
R784 VTAIL.n389 VTAIL.n366 4.26717
R785 VTAIL.n320 VTAIL.n319 4.26717
R786 VTAIL.n303 VTAIL.n280 4.26717
R787 VTAIL.n629 VTAIL.n627 3.70982
R788 VTAIL.n27 VTAIL.n25 3.70982
R789 VTAIL.n113 VTAIL.n111 3.70982
R790 VTAIL.n199 VTAIL.n197 3.70982
R791 VTAIL.n545 VTAIL.n543 3.70982
R792 VTAIL.n459 VTAIL.n457 3.70982
R793 VTAIL.n373 VTAIL.n371 3.70982
R794 VTAIL.n287 VTAIL.n285 3.70982
R795 VTAIL.n642 VTAIL.n641 3.49141
R796 VTAIL.n665 VTAIL.n612 3.49141
R797 VTAIL.n40 VTAIL.n39 3.49141
R798 VTAIL.n63 VTAIL.n10 3.49141
R799 VTAIL.n126 VTAIL.n125 3.49141
R800 VTAIL.n149 VTAIL.n96 3.49141
R801 VTAIL.n212 VTAIL.n211 3.49141
R802 VTAIL.n235 VTAIL.n182 3.49141
R803 VTAIL.n581 VTAIL.n528 3.49141
R804 VTAIL.n558 VTAIL.n557 3.49141
R805 VTAIL.n495 VTAIL.n442 3.49141
R806 VTAIL.n472 VTAIL.n471 3.49141
R807 VTAIL.n409 VTAIL.n356 3.49141
R808 VTAIL.n386 VTAIL.n385 3.49141
R809 VTAIL.n323 VTAIL.n270 3.49141
R810 VTAIL.n300 VTAIL.n299 3.49141
R811 VTAIL.n638 VTAIL.n624 2.71565
R812 VTAIL.n666 VTAIL.n610 2.71565
R813 VTAIL.n686 VTAIL.n602 2.71565
R814 VTAIL.n36 VTAIL.n22 2.71565
R815 VTAIL.n64 VTAIL.n8 2.71565
R816 VTAIL.n84 VTAIL.n0 2.71565
R817 VTAIL.n122 VTAIL.n108 2.71565
R818 VTAIL.n150 VTAIL.n94 2.71565
R819 VTAIL.n170 VTAIL.n86 2.71565
R820 VTAIL.n208 VTAIL.n194 2.71565
R821 VTAIL.n236 VTAIL.n180 2.71565
R822 VTAIL.n256 VTAIL.n172 2.71565
R823 VTAIL.n600 VTAIL.n516 2.71565
R824 VTAIL.n582 VTAIL.n526 2.71565
R825 VTAIL.n554 VTAIL.n540 2.71565
R826 VTAIL.n514 VTAIL.n430 2.71565
R827 VTAIL.n496 VTAIL.n440 2.71565
R828 VTAIL.n468 VTAIL.n454 2.71565
R829 VTAIL.n428 VTAIL.n344 2.71565
R830 VTAIL.n410 VTAIL.n354 2.71565
R831 VTAIL.n382 VTAIL.n368 2.71565
R832 VTAIL.n342 VTAIL.n258 2.71565
R833 VTAIL.n324 VTAIL.n268 2.71565
R834 VTAIL.n296 VTAIL.n282 2.71565
R835 VTAIL.n429 VTAIL.n343 2.57809
R836 VTAIL.n601 VTAIL.n515 2.57809
R837 VTAIL.n257 VTAIL.n171 2.57809
R838 VTAIL.n637 VTAIL.n626 1.93989
R839 VTAIL.n671 VTAIL.n669 1.93989
R840 VTAIL.n684 VTAIL.n683 1.93989
R841 VTAIL.n35 VTAIL.n24 1.93989
R842 VTAIL.n69 VTAIL.n67 1.93989
R843 VTAIL.n82 VTAIL.n81 1.93989
R844 VTAIL.n121 VTAIL.n110 1.93989
R845 VTAIL.n155 VTAIL.n153 1.93989
R846 VTAIL.n168 VTAIL.n167 1.93989
R847 VTAIL.n207 VTAIL.n196 1.93989
R848 VTAIL.n241 VTAIL.n239 1.93989
R849 VTAIL.n254 VTAIL.n253 1.93989
R850 VTAIL.n598 VTAIL.n597 1.93989
R851 VTAIL.n586 VTAIL.n585 1.93989
R852 VTAIL.n553 VTAIL.n542 1.93989
R853 VTAIL.n512 VTAIL.n511 1.93989
R854 VTAIL.n500 VTAIL.n499 1.93989
R855 VTAIL.n467 VTAIL.n456 1.93989
R856 VTAIL.n426 VTAIL.n425 1.93989
R857 VTAIL.n414 VTAIL.n413 1.93989
R858 VTAIL.n381 VTAIL.n370 1.93989
R859 VTAIL.n340 VTAIL.n339 1.93989
R860 VTAIL.n328 VTAIL.n327 1.93989
R861 VTAIL.n295 VTAIL.n284 1.93989
R862 VTAIL VTAIL.n85 1.34748
R863 VTAIL VTAIL.n687 1.2311
R864 VTAIL.n634 VTAIL.n633 1.16414
R865 VTAIL.n670 VTAIL.n608 1.16414
R866 VTAIL.n680 VTAIL.n604 1.16414
R867 VTAIL.n32 VTAIL.n31 1.16414
R868 VTAIL.n68 VTAIL.n6 1.16414
R869 VTAIL.n78 VTAIL.n2 1.16414
R870 VTAIL.n118 VTAIL.n117 1.16414
R871 VTAIL.n154 VTAIL.n92 1.16414
R872 VTAIL.n164 VTAIL.n88 1.16414
R873 VTAIL.n204 VTAIL.n203 1.16414
R874 VTAIL.n240 VTAIL.n178 1.16414
R875 VTAIL.n250 VTAIL.n174 1.16414
R876 VTAIL.n594 VTAIL.n518 1.16414
R877 VTAIL.n589 VTAIL.n523 1.16414
R878 VTAIL.n550 VTAIL.n549 1.16414
R879 VTAIL.n508 VTAIL.n432 1.16414
R880 VTAIL.n503 VTAIL.n437 1.16414
R881 VTAIL.n464 VTAIL.n463 1.16414
R882 VTAIL.n422 VTAIL.n346 1.16414
R883 VTAIL.n417 VTAIL.n351 1.16414
R884 VTAIL.n378 VTAIL.n377 1.16414
R885 VTAIL.n336 VTAIL.n260 1.16414
R886 VTAIL.n331 VTAIL.n265 1.16414
R887 VTAIL.n292 VTAIL.n291 1.16414
R888 VTAIL.n515 VTAIL.n429 0.470328
R889 VTAIL.n171 VTAIL.n85 0.470328
R890 VTAIL.n630 VTAIL.n628 0.388379
R891 VTAIL.n676 VTAIL.n675 0.388379
R892 VTAIL.n679 VTAIL.n606 0.388379
R893 VTAIL.n28 VTAIL.n26 0.388379
R894 VTAIL.n74 VTAIL.n73 0.388379
R895 VTAIL.n77 VTAIL.n4 0.388379
R896 VTAIL.n114 VTAIL.n112 0.388379
R897 VTAIL.n160 VTAIL.n159 0.388379
R898 VTAIL.n163 VTAIL.n90 0.388379
R899 VTAIL.n200 VTAIL.n198 0.388379
R900 VTAIL.n246 VTAIL.n245 0.388379
R901 VTAIL.n249 VTAIL.n176 0.388379
R902 VTAIL.n593 VTAIL.n520 0.388379
R903 VTAIL.n590 VTAIL.n522 0.388379
R904 VTAIL.n546 VTAIL.n544 0.388379
R905 VTAIL.n507 VTAIL.n434 0.388379
R906 VTAIL.n504 VTAIL.n436 0.388379
R907 VTAIL.n460 VTAIL.n458 0.388379
R908 VTAIL.n421 VTAIL.n348 0.388379
R909 VTAIL.n418 VTAIL.n350 0.388379
R910 VTAIL.n374 VTAIL.n372 0.388379
R911 VTAIL.n335 VTAIL.n262 0.388379
R912 VTAIL.n332 VTAIL.n264 0.388379
R913 VTAIL.n288 VTAIL.n286 0.388379
R914 VTAIL.n635 VTAIL.n627 0.155672
R915 VTAIL.n636 VTAIL.n635 0.155672
R916 VTAIL.n636 VTAIL.n623 0.155672
R917 VTAIL.n643 VTAIL.n623 0.155672
R918 VTAIL.n644 VTAIL.n643 0.155672
R919 VTAIL.n644 VTAIL.n619 0.155672
R920 VTAIL.n651 VTAIL.n619 0.155672
R921 VTAIL.n652 VTAIL.n651 0.155672
R922 VTAIL.n652 VTAIL.n615 0.155672
R923 VTAIL.n659 VTAIL.n615 0.155672
R924 VTAIL.n660 VTAIL.n659 0.155672
R925 VTAIL.n660 VTAIL.n611 0.155672
R926 VTAIL.n667 VTAIL.n611 0.155672
R927 VTAIL.n668 VTAIL.n667 0.155672
R928 VTAIL.n668 VTAIL.n607 0.155672
R929 VTAIL.n677 VTAIL.n607 0.155672
R930 VTAIL.n678 VTAIL.n677 0.155672
R931 VTAIL.n678 VTAIL.n603 0.155672
R932 VTAIL.n685 VTAIL.n603 0.155672
R933 VTAIL.n33 VTAIL.n25 0.155672
R934 VTAIL.n34 VTAIL.n33 0.155672
R935 VTAIL.n34 VTAIL.n21 0.155672
R936 VTAIL.n41 VTAIL.n21 0.155672
R937 VTAIL.n42 VTAIL.n41 0.155672
R938 VTAIL.n42 VTAIL.n17 0.155672
R939 VTAIL.n49 VTAIL.n17 0.155672
R940 VTAIL.n50 VTAIL.n49 0.155672
R941 VTAIL.n50 VTAIL.n13 0.155672
R942 VTAIL.n57 VTAIL.n13 0.155672
R943 VTAIL.n58 VTAIL.n57 0.155672
R944 VTAIL.n58 VTAIL.n9 0.155672
R945 VTAIL.n65 VTAIL.n9 0.155672
R946 VTAIL.n66 VTAIL.n65 0.155672
R947 VTAIL.n66 VTAIL.n5 0.155672
R948 VTAIL.n75 VTAIL.n5 0.155672
R949 VTAIL.n76 VTAIL.n75 0.155672
R950 VTAIL.n76 VTAIL.n1 0.155672
R951 VTAIL.n83 VTAIL.n1 0.155672
R952 VTAIL.n119 VTAIL.n111 0.155672
R953 VTAIL.n120 VTAIL.n119 0.155672
R954 VTAIL.n120 VTAIL.n107 0.155672
R955 VTAIL.n127 VTAIL.n107 0.155672
R956 VTAIL.n128 VTAIL.n127 0.155672
R957 VTAIL.n128 VTAIL.n103 0.155672
R958 VTAIL.n135 VTAIL.n103 0.155672
R959 VTAIL.n136 VTAIL.n135 0.155672
R960 VTAIL.n136 VTAIL.n99 0.155672
R961 VTAIL.n143 VTAIL.n99 0.155672
R962 VTAIL.n144 VTAIL.n143 0.155672
R963 VTAIL.n144 VTAIL.n95 0.155672
R964 VTAIL.n151 VTAIL.n95 0.155672
R965 VTAIL.n152 VTAIL.n151 0.155672
R966 VTAIL.n152 VTAIL.n91 0.155672
R967 VTAIL.n161 VTAIL.n91 0.155672
R968 VTAIL.n162 VTAIL.n161 0.155672
R969 VTAIL.n162 VTAIL.n87 0.155672
R970 VTAIL.n169 VTAIL.n87 0.155672
R971 VTAIL.n205 VTAIL.n197 0.155672
R972 VTAIL.n206 VTAIL.n205 0.155672
R973 VTAIL.n206 VTAIL.n193 0.155672
R974 VTAIL.n213 VTAIL.n193 0.155672
R975 VTAIL.n214 VTAIL.n213 0.155672
R976 VTAIL.n214 VTAIL.n189 0.155672
R977 VTAIL.n221 VTAIL.n189 0.155672
R978 VTAIL.n222 VTAIL.n221 0.155672
R979 VTAIL.n222 VTAIL.n185 0.155672
R980 VTAIL.n229 VTAIL.n185 0.155672
R981 VTAIL.n230 VTAIL.n229 0.155672
R982 VTAIL.n230 VTAIL.n181 0.155672
R983 VTAIL.n237 VTAIL.n181 0.155672
R984 VTAIL.n238 VTAIL.n237 0.155672
R985 VTAIL.n238 VTAIL.n177 0.155672
R986 VTAIL.n247 VTAIL.n177 0.155672
R987 VTAIL.n248 VTAIL.n247 0.155672
R988 VTAIL.n248 VTAIL.n173 0.155672
R989 VTAIL.n255 VTAIL.n173 0.155672
R990 VTAIL.n599 VTAIL.n517 0.155672
R991 VTAIL.n592 VTAIL.n517 0.155672
R992 VTAIL.n592 VTAIL.n591 0.155672
R993 VTAIL.n591 VTAIL.n521 0.155672
R994 VTAIL.n584 VTAIL.n521 0.155672
R995 VTAIL.n584 VTAIL.n583 0.155672
R996 VTAIL.n583 VTAIL.n527 0.155672
R997 VTAIL.n576 VTAIL.n527 0.155672
R998 VTAIL.n576 VTAIL.n575 0.155672
R999 VTAIL.n575 VTAIL.n531 0.155672
R1000 VTAIL.n568 VTAIL.n531 0.155672
R1001 VTAIL.n568 VTAIL.n567 0.155672
R1002 VTAIL.n567 VTAIL.n535 0.155672
R1003 VTAIL.n560 VTAIL.n535 0.155672
R1004 VTAIL.n560 VTAIL.n559 0.155672
R1005 VTAIL.n559 VTAIL.n539 0.155672
R1006 VTAIL.n552 VTAIL.n539 0.155672
R1007 VTAIL.n552 VTAIL.n551 0.155672
R1008 VTAIL.n551 VTAIL.n543 0.155672
R1009 VTAIL.n513 VTAIL.n431 0.155672
R1010 VTAIL.n506 VTAIL.n431 0.155672
R1011 VTAIL.n506 VTAIL.n505 0.155672
R1012 VTAIL.n505 VTAIL.n435 0.155672
R1013 VTAIL.n498 VTAIL.n435 0.155672
R1014 VTAIL.n498 VTAIL.n497 0.155672
R1015 VTAIL.n497 VTAIL.n441 0.155672
R1016 VTAIL.n490 VTAIL.n441 0.155672
R1017 VTAIL.n490 VTAIL.n489 0.155672
R1018 VTAIL.n489 VTAIL.n445 0.155672
R1019 VTAIL.n482 VTAIL.n445 0.155672
R1020 VTAIL.n482 VTAIL.n481 0.155672
R1021 VTAIL.n481 VTAIL.n449 0.155672
R1022 VTAIL.n474 VTAIL.n449 0.155672
R1023 VTAIL.n474 VTAIL.n473 0.155672
R1024 VTAIL.n473 VTAIL.n453 0.155672
R1025 VTAIL.n466 VTAIL.n453 0.155672
R1026 VTAIL.n466 VTAIL.n465 0.155672
R1027 VTAIL.n465 VTAIL.n457 0.155672
R1028 VTAIL.n427 VTAIL.n345 0.155672
R1029 VTAIL.n420 VTAIL.n345 0.155672
R1030 VTAIL.n420 VTAIL.n419 0.155672
R1031 VTAIL.n419 VTAIL.n349 0.155672
R1032 VTAIL.n412 VTAIL.n349 0.155672
R1033 VTAIL.n412 VTAIL.n411 0.155672
R1034 VTAIL.n411 VTAIL.n355 0.155672
R1035 VTAIL.n404 VTAIL.n355 0.155672
R1036 VTAIL.n404 VTAIL.n403 0.155672
R1037 VTAIL.n403 VTAIL.n359 0.155672
R1038 VTAIL.n396 VTAIL.n359 0.155672
R1039 VTAIL.n396 VTAIL.n395 0.155672
R1040 VTAIL.n395 VTAIL.n363 0.155672
R1041 VTAIL.n388 VTAIL.n363 0.155672
R1042 VTAIL.n388 VTAIL.n387 0.155672
R1043 VTAIL.n387 VTAIL.n367 0.155672
R1044 VTAIL.n380 VTAIL.n367 0.155672
R1045 VTAIL.n380 VTAIL.n379 0.155672
R1046 VTAIL.n379 VTAIL.n371 0.155672
R1047 VTAIL.n341 VTAIL.n259 0.155672
R1048 VTAIL.n334 VTAIL.n259 0.155672
R1049 VTAIL.n334 VTAIL.n333 0.155672
R1050 VTAIL.n333 VTAIL.n263 0.155672
R1051 VTAIL.n326 VTAIL.n263 0.155672
R1052 VTAIL.n326 VTAIL.n325 0.155672
R1053 VTAIL.n325 VTAIL.n269 0.155672
R1054 VTAIL.n318 VTAIL.n269 0.155672
R1055 VTAIL.n318 VTAIL.n317 0.155672
R1056 VTAIL.n317 VTAIL.n273 0.155672
R1057 VTAIL.n310 VTAIL.n273 0.155672
R1058 VTAIL.n310 VTAIL.n309 0.155672
R1059 VTAIL.n309 VTAIL.n277 0.155672
R1060 VTAIL.n302 VTAIL.n277 0.155672
R1061 VTAIL.n302 VTAIL.n301 0.155672
R1062 VTAIL.n301 VTAIL.n281 0.155672
R1063 VTAIL.n294 VTAIL.n281 0.155672
R1064 VTAIL.n294 VTAIL.n293 0.155672
R1065 VTAIL.n293 VTAIL.n285 0.155672
R1066 VDD1 VDD1.n1 118.105
R1067 VDD1 VDD1.n0 72.8374
R1068 VDD1.n0 VDD1.t2 2.09895
R1069 VDD1.n0 VDD1.t3 2.09895
R1070 VDD1.n1 VDD1.t0 2.09895
R1071 VDD1.n1 VDD1.t1 2.09895
R1072 VN.n1 VN.t2 174.056
R1073 VN.n0 VN.t1 174.056
R1074 VN.n0 VN.t3 173.195
R1075 VN.n1 VN.t0 173.195
R1076 VN VN.n1 53.0136
R1077 VN VN.n0 3.72197
R1078 VDD2.n2 VDD2.n0 117.581
R1079 VDD2.n2 VDD2.n1 72.7792
R1080 VDD2.n1 VDD2.t3 2.09895
R1081 VDD2.n1 VDD2.t1 2.09895
R1082 VDD2.n0 VDD2.t2 2.09895
R1083 VDD2.n0 VDD2.t0 2.09895
R1084 VDD2 VDD2.n2 0.0586897
R1085 B.n412 B.n411 585
R1086 B.n410 B.n115 585
R1087 B.n409 B.n408 585
R1088 B.n407 B.n116 585
R1089 B.n406 B.n405 585
R1090 B.n404 B.n117 585
R1091 B.n403 B.n402 585
R1092 B.n401 B.n118 585
R1093 B.n400 B.n399 585
R1094 B.n398 B.n119 585
R1095 B.n397 B.n396 585
R1096 B.n395 B.n120 585
R1097 B.n394 B.n393 585
R1098 B.n392 B.n121 585
R1099 B.n391 B.n390 585
R1100 B.n389 B.n122 585
R1101 B.n388 B.n387 585
R1102 B.n386 B.n123 585
R1103 B.n385 B.n384 585
R1104 B.n383 B.n124 585
R1105 B.n382 B.n381 585
R1106 B.n380 B.n125 585
R1107 B.n379 B.n378 585
R1108 B.n377 B.n126 585
R1109 B.n376 B.n375 585
R1110 B.n374 B.n127 585
R1111 B.n373 B.n372 585
R1112 B.n371 B.n128 585
R1113 B.n370 B.n369 585
R1114 B.n368 B.n129 585
R1115 B.n367 B.n366 585
R1116 B.n365 B.n130 585
R1117 B.n364 B.n363 585
R1118 B.n362 B.n131 585
R1119 B.n361 B.n360 585
R1120 B.n359 B.n132 585
R1121 B.n358 B.n357 585
R1122 B.n356 B.n133 585
R1123 B.n355 B.n354 585
R1124 B.n353 B.n134 585
R1125 B.n352 B.n351 585
R1126 B.n350 B.n135 585
R1127 B.n349 B.n348 585
R1128 B.n347 B.n136 585
R1129 B.n346 B.n345 585
R1130 B.n344 B.n137 585
R1131 B.n343 B.n342 585
R1132 B.n341 B.n138 585
R1133 B.n340 B.n339 585
R1134 B.n338 B.n139 585
R1135 B.n337 B.n336 585
R1136 B.n335 B.n140 585
R1137 B.n334 B.n333 585
R1138 B.n329 B.n141 585
R1139 B.n328 B.n327 585
R1140 B.n326 B.n142 585
R1141 B.n325 B.n324 585
R1142 B.n323 B.n143 585
R1143 B.n322 B.n321 585
R1144 B.n320 B.n144 585
R1145 B.n319 B.n318 585
R1146 B.n316 B.n145 585
R1147 B.n315 B.n314 585
R1148 B.n313 B.n148 585
R1149 B.n312 B.n311 585
R1150 B.n310 B.n149 585
R1151 B.n309 B.n308 585
R1152 B.n307 B.n150 585
R1153 B.n306 B.n305 585
R1154 B.n304 B.n151 585
R1155 B.n303 B.n302 585
R1156 B.n301 B.n152 585
R1157 B.n300 B.n299 585
R1158 B.n298 B.n153 585
R1159 B.n297 B.n296 585
R1160 B.n295 B.n154 585
R1161 B.n294 B.n293 585
R1162 B.n292 B.n155 585
R1163 B.n291 B.n290 585
R1164 B.n289 B.n156 585
R1165 B.n288 B.n287 585
R1166 B.n286 B.n157 585
R1167 B.n285 B.n284 585
R1168 B.n283 B.n158 585
R1169 B.n282 B.n281 585
R1170 B.n280 B.n159 585
R1171 B.n279 B.n278 585
R1172 B.n277 B.n160 585
R1173 B.n276 B.n275 585
R1174 B.n274 B.n161 585
R1175 B.n273 B.n272 585
R1176 B.n271 B.n162 585
R1177 B.n270 B.n269 585
R1178 B.n268 B.n163 585
R1179 B.n267 B.n266 585
R1180 B.n265 B.n164 585
R1181 B.n264 B.n263 585
R1182 B.n262 B.n165 585
R1183 B.n261 B.n260 585
R1184 B.n259 B.n166 585
R1185 B.n258 B.n257 585
R1186 B.n256 B.n167 585
R1187 B.n255 B.n254 585
R1188 B.n253 B.n168 585
R1189 B.n252 B.n251 585
R1190 B.n250 B.n169 585
R1191 B.n249 B.n248 585
R1192 B.n247 B.n170 585
R1193 B.n246 B.n245 585
R1194 B.n244 B.n171 585
R1195 B.n243 B.n242 585
R1196 B.n241 B.n172 585
R1197 B.n240 B.n239 585
R1198 B.n413 B.n114 585
R1199 B.n415 B.n414 585
R1200 B.n416 B.n113 585
R1201 B.n418 B.n417 585
R1202 B.n419 B.n112 585
R1203 B.n421 B.n420 585
R1204 B.n422 B.n111 585
R1205 B.n424 B.n423 585
R1206 B.n425 B.n110 585
R1207 B.n427 B.n426 585
R1208 B.n428 B.n109 585
R1209 B.n430 B.n429 585
R1210 B.n431 B.n108 585
R1211 B.n433 B.n432 585
R1212 B.n434 B.n107 585
R1213 B.n436 B.n435 585
R1214 B.n437 B.n106 585
R1215 B.n439 B.n438 585
R1216 B.n440 B.n105 585
R1217 B.n442 B.n441 585
R1218 B.n443 B.n104 585
R1219 B.n445 B.n444 585
R1220 B.n446 B.n103 585
R1221 B.n448 B.n447 585
R1222 B.n449 B.n102 585
R1223 B.n451 B.n450 585
R1224 B.n452 B.n101 585
R1225 B.n454 B.n453 585
R1226 B.n455 B.n100 585
R1227 B.n457 B.n456 585
R1228 B.n458 B.n99 585
R1229 B.n460 B.n459 585
R1230 B.n461 B.n98 585
R1231 B.n463 B.n462 585
R1232 B.n464 B.n97 585
R1233 B.n466 B.n465 585
R1234 B.n467 B.n96 585
R1235 B.n469 B.n468 585
R1236 B.n470 B.n95 585
R1237 B.n472 B.n471 585
R1238 B.n473 B.n94 585
R1239 B.n475 B.n474 585
R1240 B.n476 B.n93 585
R1241 B.n478 B.n477 585
R1242 B.n479 B.n92 585
R1243 B.n481 B.n480 585
R1244 B.n482 B.n91 585
R1245 B.n484 B.n483 585
R1246 B.n485 B.n90 585
R1247 B.n487 B.n486 585
R1248 B.n488 B.n89 585
R1249 B.n490 B.n489 585
R1250 B.n491 B.n88 585
R1251 B.n493 B.n492 585
R1252 B.n494 B.n87 585
R1253 B.n496 B.n495 585
R1254 B.n497 B.n86 585
R1255 B.n499 B.n498 585
R1256 B.n500 B.n85 585
R1257 B.n502 B.n501 585
R1258 B.n503 B.n84 585
R1259 B.n505 B.n504 585
R1260 B.n506 B.n83 585
R1261 B.n508 B.n507 585
R1262 B.n509 B.n82 585
R1263 B.n511 B.n510 585
R1264 B.n512 B.n81 585
R1265 B.n514 B.n513 585
R1266 B.n515 B.n80 585
R1267 B.n517 B.n516 585
R1268 B.n688 B.n19 585
R1269 B.n687 B.n686 585
R1270 B.n685 B.n20 585
R1271 B.n684 B.n683 585
R1272 B.n682 B.n21 585
R1273 B.n681 B.n680 585
R1274 B.n679 B.n22 585
R1275 B.n678 B.n677 585
R1276 B.n676 B.n23 585
R1277 B.n675 B.n674 585
R1278 B.n673 B.n24 585
R1279 B.n672 B.n671 585
R1280 B.n670 B.n25 585
R1281 B.n669 B.n668 585
R1282 B.n667 B.n26 585
R1283 B.n666 B.n665 585
R1284 B.n664 B.n27 585
R1285 B.n663 B.n662 585
R1286 B.n661 B.n28 585
R1287 B.n660 B.n659 585
R1288 B.n658 B.n29 585
R1289 B.n657 B.n656 585
R1290 B.n655 B.n30 585
R1291 B.n654 B.n653 585
R1292 B.n652 B.n31 585
R1293 B.n651 B.n650 585
R1294 B.n649 B.n32 585
R1295 B.n648 B.n647 585
R1296 B.n646 B.n33 585
R1297 B.n645 B.n644 585
R1298 B.n643 B.n34 585
R1299 B.n642 B.n641 585
R1300 B.n640 B.n35 585
R1301 B.n639 B.n638 585
R1302 B.n637 B.n36 585
R1303 B.n636 B.n635 585
R1304 B.n634 B.n37 585
R1305 B.n633 B.n632 585
R1306 B.n631 B.n38 585
R1307 B.n630 B.n629 585
R1308 B.n628 B.n39 585
R1309 B.n627 B.n626 585
R1310 B.n625 B.n40 585
R1311 B.n624 B.n623 585
R1312 B.n622 B.n41 585
R1313 B.n621 B.n620 585
R1314 B.n619 B.n42 585
R1315 B.n618 B.n617 585
R1316 B.n616 B.n43 585
R1317 B.n615 B.n614 585
R1318 B.n613 B.n44 585
R1319 B.n612 B.n611 585
R1320 B.n609 B.n45 585
R1321 B.n608 B.n607 585
R1322 B.n606 B.n48 585
R1323 B.n605 B.n604 585
R1324 B.n603 B.n49 585
R1325 B.n602 B.n601 585
R1326 B.n600 B.n50 585
R1327 B.n599 B.n598 585
R1328 B.n597 B.n51 585
R1329 B.n595 B.n594 585
R1330 B.n593 B.n54 585
R1331 B.n592 B.n591 585
R1332 B.n590 B.n55 585
R1333 B.n589 B.n588 585
R1334 B.n587 B.n56 585
R1335 B.n586 B.n585 585
R1336 B.n584 B.n57 585
R1337 B.n583 B.n582 585
R1338 B.n581 B.n58 585
R1339 B.n580 B.n579 585
R1340 B.n578 B.n59 585
R1341 B.n577 B.n576 585
R1342 B.n575 B.n60 585
R1343 B.n574 B.n573 585
R1344 B.n572 B.n61 585
R1345 B.n571 B.n570 585
R1346 B.n569 B.n62 585
R1347 B.n568 B.n567 585
R1348 B.n566 B.n63 585
R1349 B.n565 B.n564 585
R1350 B.n563 B.n64 585
R1351 B.n562 B.n561 585
R1352 B.n560 B.n65 585
R1353 B.n559 B.n558 585
R1354 B.n557 B.n66 585
R1355 B.n556 B.n555 585
R1356 B.n554 B.n67 585
R1357 B.n553 B.n552 585
R1358 B.n551 B.n68 585
R1359 B.n550 B.n549 585
R1360 B.n548 B.n69 585
R1361 B.n547 B.n546 585
R1362 B.n545 B.n70 585
R1363 B.n544 B.n543 585
R1364 B.n542 B.n71 585
R1365 B.n541 B.n540 585
R1366 B.n539 B.n72 585
R1367 B.n538 B.n537 585
R1368 B.n536 B.n73 585
R1369 B.n535 B.n534 585
R1370 B.n533 B.n74 585
R1371 B.n532 B.n531 585
R1372 B.n530 B.n75 585
R1373 B.n529 B.n528 585
R1374 B.n527 B.n76 585
R1375 B.n526 B.n525 585
R1376 B.n524 B.n77 585
R1377 B.n523 B.n522 585
R1378 B.n521 B.n78 585
R1379 B.n520 B.n519 585
R1380 B.n518 B.n79 585
R1381 B.n690 B.n689 585
R1382 B.n691 B.n18 585
R1383 B.n693 B.n692 585
R1384 B.n694 B.n17 585
R1385 B.n696 B.n695 585
R1386 B.n697 B.n16 585
R1387 B.n699 B.n698 585
R1388 B.n700 B.n15 585
R1389 B.n702 B.n701 585
R1390 B.n703 B.n14 585
R1391 B.n705 B.n704 585
R1392 B.n706 B.n13 585
R1393 B.n708 B.n707 585
R1394 B.n709 B.n12 585
R1395 B.n711 B.n710 585
R1396 B.n712 B.n11 585
R1397 B.n714 B.n713 585
R1398 B.n715 B.n10 585
R1399 B.n717 B.n716 585
R1400 B.n718 B.n9 585
R1401 B.n720 B.n719 585
R1402 B.n721 B.n8 585
R1403 B.n723 B.n722 585
R1404 B.n724 B.n7 585
R1405 B.n726 B.n725 585
R1406 B.n727 B.n6 585
R1407 B.n729 B.n728 585
R1408 B.n730 B.n5 585
R1409 B.n732 B.n731 585
R1410 B.n733 B.n4 585
R1411 B.n735 B.n734 585
R1412 B.n736 B.n3 585
R1413 B.n738 B.n737 585
R1414 B.n739 B.n0 585
R1415 B.n2 B.n1 585
R1416 B.n190 B.n189 585
R1417 B.n192 B.n191 585
R1418 B.n193 B.n188 585
R1419 B.n195 B.n194 585
R1420 B.n196 B.n187 585
R1421 B.n198 B.n197 585
R1422 B.n199 B.n186 585
R1423 B.n201 B.n200 585
R1424 B.n202 B.n185 585
R1425 B.n204 B.n203 585
R1426 B.n205 B.n184 585
R1427 B.n207 B.n206 585
R1428 B.n208 B.n183 585
R1429 B.n210 B.n209 585
R1430 B.n211 B.n182 585
R1431 B.n213 B.n212 585
R1432 B.n214 B.n181 585
R1433 B.n216 B.n215 585
R1434 B.n217 B.n180 585
R1435 B.n219 B.n218 585
R1436 B.n220 B.n179 585
R1437 B.n222 B.n221 585
R1438 B.n223 B.n178 585
R1439 B.n225 B.n224 585
R1440 B.n226 B.n177 585
R1441 B.n228 B.n227 585
R1442 B.n229 B.n176 585
R1443 B.n231 B.n230 585
R1444 B.n232 B.n175 585
R1445 B.n234 B.n233 585
R1446 B.n235 B.n174 585
R1447 B.n237 B.n236 585
R1448 B.n238 B.n173 585
R1449 B.n240 B.n173 526.135
R1450 B.n413 B.n412 526.135
R1451 B.n516 B.n79 526.135
R1452 B.n690 B.n19 526.135
R1453 B.n330 B.t7 496.502
R1454 B.n52 B.t2 496.502
R1455 B.n146 B.t10 496.502
R1456 B.n46 B.t5 496.502
R1457 B.n331 B.t8 438.514
R1458 B.n53 B.t1 438.514
R1459 B.n147 B.t11 438.514
R1460 B.n47 B.t4 438.514
R1461 B.n146 B.t9 348.478
R1462 B.n330 B.t6 348.478
R1463 B.n52 B.t0 348.478
R1464 B.n46 B.t3 348.478
R1465 B.n741 B.n740 256.663
R1466 B.n740 B.n739 235.042
R1467 B.n740 B.n2 235.042
R1468 B.n241 B.n240 163.367
R1469 B.n242 B.n241 163.367
R1470 B.n242 B.n171 163.367
R1471 B.n246 B.n171 163.367
R1472 B.n247 B.n246 163.367
R1473 B.n248 B.n247 163.367
R1474 B.n248 B.n169 163.367
R1475 B.n252 B.n169 163.367
R1476 B.n253 B.n252 163.367
R1477 B.n254 B.n253 163.367
R1478 B.n254 B.n167 163.367
R1479 B.n258 B.n167 163.367
R1480 B.n259 B.n258 163.367
R1481 B.n260 B.n259 163.367
R1482 B.n260 B.n165 163.367
R1483 B.n264 B.n165 163.367
R1484 B.n265 B.n264 163.367
R1485 B.n266 B.n265 163.367
R1486 B.n266 B.n163 163.367
R1487 B.n270 B.n163 163.367
R1488 B.n271 B.n270 163.367
R1489 B.n272 B.n271 163.367
R1490 B.n272 B.n161 163.367
R1491 B.n276 B.n161 163.367
R1492 B.n277 B.n276 163.367
R1493 B.n278 B.n277 163.367
R1494 B.n278 B.n159 163.367
R1495 B.n282 B.n159 163.367
R1496 B.n283 B.n282 163.367
R1497 B.n284 B.n283 163.367
R1498 B.n284 B.n157 163.367
R1499 B.n288 B.n157 163.367
R1500 B.n289 B.n288 163.367
R1501 B.n290 B.n289 163.367
R1502 B.n290 B.n155 163.367
R1503 B.n294 B.n155 163.367
R1504 B.n295 B.n294 163.367
R1505 B.n296 B.n295 163.367
R1506 B.n296 B.n153 163.367
R1507 B.n300 B.n153 163.367
R1508 B.n301 B.n300 163.367
R1509 B.n302 B.n301 163.367
R1510 B.n302 B.n151 163.367
R1511 B.n306 B.n151 163.367
R1512 B.n307 B.n306 163.367
R1513 B.n308 B.n307 163.367
R1514 B.n308 B.n149 163.367
R1515 B.n312 B.n149 163.367
R1516 B.n313 B.n312 163.367
R1517 B.n314 B.n313 163.367
R1518 B.n314 B.n145 163.367
R1519 B.n319 B.n145 163.367
R1520 B.n320 B.n319 163.367
R1521 B.n321 B.n320 163.367
R1522 B.n321 B.n143 163.367
R1523 B.n325 B.n143 163.367
R1524 B.n326 B.n325 163.367
R1525 B.n327 B.n326 163.367
R1526 B.n327 B.n141 163.367
R1527 B.n334 B.n141 163.367
R1528 B.n335 B.n334 163.367
R1529 B.n336 B.n335 163.367
R1530 B.n336 B.n139 163.367
R1531 B.n340 B.n139 163.367
R1532 B.n341 B.n340 163.367
R1533 B.n342 B.n341 163.367
R1534 B.n342 B.n137 163.367
R1535 B.n346 B.n137 163.367
R1536 B.n347 B.n346 163.367
R1537 B.n348 B.n347 163.367
R1538 B.n348 B.n135 163.367
R1539 B.n352 B.n135 163.367
R1540 B.n353 B.n352 163.367
R1541 B.n354 B.n353 163.367
R1542 B.n354 B.n133 163.367
R1543 B.n358 B.n133 163.367
R1544 B.n359 B.n358 163.367
R1545 B.n360 B.n359 163.367
R1546 B.n360 B.n131 163.367
R1547 B.n364 B.n131 163.367
R1548 B.n365 B.n364 163.367
R1549 B.n366 B.n365 163.367
R1550 B.n366 B.n129 163.367
R1551 B.n370 B.n129 163.367
R1552 B.n371 B.n370 163.367
R1553 B.n372 B.n371 163.367
R1554 B.n372 B.n127 163.367
R1555 B.n376 B.n127 163.367
R1556 B.n377 B.n376 163.367
R1557 B.n378 B.n377 163.367
R1558 B.n378 B.n125 163.367
R1559 B.n382 B.n125 163.367
R1560 B.n383 B.n382 163.367
R1561 B.n384 B.n383 163.367
R1562 B.n384 B.n123 163.367
R1563 B.n388 B.n123 163.367
R1564 B.n389 B.n388 163.367
R1565 B.n390 B.n389 163.367
R1566 B.n390 B.n121 163.367
R1567 B.n394 B.n121 163.367
R1568 B.n395 B.n394 163.367
R1569 B.n396 B.n395 163.367
R1570 B.n396 B.n119 163.367
R1571 B.n400 B.n119 163.367
R1572 B.n401 B.n400 163.367
R1573 B.n402 B.n401 163.367
R1574 B.n402 B.n117 163.367
R1575 B.n406 B.n117 163.367
R1576 B.n407 B.n406 163.367
R1577 B.n408 B.n407 163.367
R1578 B.n408 B.n115 163.367
R1579 B.n412 B.n115 163.367
R1580 B.n516 B.n515 163.367
R1581 B.n515 B.n514 163.367
R1582 B.n514 B.n81 163.367
R1583 B.n510 B.n81 163.367
R1584 B.n510 B.n509 163.367
R1585 B.n509 B.n508 163.367
R1586 B.n508 B.n83 163.367
R1587 B.n504 B.n83 163.367
R1588 B.n504 B.n503 163.367
R1589 B.n503 B.n502 163.367
R1590 B.n502 B.n85 163.367
R1591 B.n498 B.n85 163.367
R1592 B.n498 B.n497 163.367
R1593 B.n497 B.n496 163.367
R1594 B.n496 B.n87 163.367
R1595 B.n492 B.n87 163.367
R1596 B.n492 B.n491 163.367
R1597 B.n491 B.n490 163.367
R1598 B.n490 B.n89 163.367
R1599 B.n486 B.n89 163.367
R1600 B.n486 B.n485 163.367
R1601 B.n485 B.n484 163.367
R1602 B.n484 B.n91 163.367
R1603 B.n480 B.n91 163.367
R1604 B.n480 B.n479 163.367
R1605 B.n479 B.n478 163.367
R1606 B.n478 B.n93 163.367
R1607 B.n474 B.n93 163.367
R1608 B.n474 B.n473 163.367
R1609 B.n473 B.n472 163.367
R1610 B.n472 B.n95 163.367
R1611 B.n468 B.n95 163.367
R1612 B.n468 B.n467 163.367
R1613 B.n467 B.n466 163.367
R1614 B.n466 B.n97 163.367
R1615 B.n462 B.n97 163.367
R1616 B.n462 B.n461 163.367
R1617 B.n461 B.n460 163.367
R1618 B.n460 B.n99 163.367
R1619 B.n456 B.n99 163.367
R1620 B.n456 B.n455 163.367
R1621 B.n455 B.n454 163.367
R1622 B.n454 B.n101 163.367
R1623 B.n450 B.n101 163.367
R1624 B.n450 B.n449 163.367
R1625 B.n449 B.n448 163.367
R1626 B.n448 B.n103 163.367
R1627 B.n444 B.n103 163.367
R1628 B.n444 B.n443 163.367
R1629 B.n443 B.n442 163.367
R1630 B.n442 B.n105 163.367
R1631 B.n438 B.n105 163.367
R1632 B.n438 B.n437 163.367
R1633 B.n437 B.n436 163.367
R1634 B.n436 B.n107 163.367
R1635 B.n432 B.n107 163.367
R1636 B.n432 B.n431 163.367
R1637 B.n431 B.n430 163.367
R1638 B.n430 B.n109 163.367
R1639 B.n426 B.n109 163.367
R1640 B.n426 B.n425 163.367
R1641 B.n425 B.n424 163.367
R1642 B.n424 B.n111 163.367
R1643 B.n420 B.n111 163.367
R1644 B.n420 B.n419 163.367
R1645 B.n419 B.n418 163.367
R1646 B.n418 B.n113 163.367
R1647 B.n414 B.n113 163.367
R1648 B.n414 B.n413 163.367
R1649 B.n686 B.n19 163.367
R1650 B.n686 B.n685 163.367
R1651 B.n685 B.n684 163.367
R1652 B.n684 B.n21 163.367
R1653 B.n680 B.n21 163.367
R1654 B.n680 B.n679 163.367
R1655 B.n679 B.n678 163.367
R1656 B.n678 B.n23 163.367
R1657 B.n674 B.n23 163.367
R1658 B.n674 B.n673 163.367
R1659 B.n673 B.n672 163.367
R1660 B.n672 B.n25 163.367
R1661 B.n668 B.n25 163.367
R1662 B.n668 B.n667 163.367
R1663 B.n667 B.n666 163.367
R1664 B.n666 B.n27 163.367
R1665 B.n662 B.n27 163.367
R1666 B.n662 B.n661 163.367
R1667 B.n661 B.n660 163.367
R1668 B.n660 B.n29 163.367
R1669 B.n656 B.n29 163.367
R1670 B.n656 B.n655 163.367
R1671 B.n655 B.n654 163.367
R1672 B.n654 B.n31 163.367
R1673 B.n650 B.n31 163.367
R1674 B.n650 B.n649 163.367
R1675 B.n649 B.n648 163.367
R1676 B.n648 B.n33 163.367
R1677 B.n644 B.n33 163.367
R1678 B.n644 B.n643 163.367
R1679 B.n643 B.n642 163.367
R1680 B.n642 B.n35 163.367
R1681 B.n638 B.n35 163.367
R1682 B.n638 B.n637 163.367
R1683 B.n637 B.n636 163.367
R1684 B.n636 B.n37 163.367
R1685 B.n632 B.n37 163.367
R1686 B.n632 B.n631 163.367
R1687 B.n631 B.n630 163.367
R1688 B.n630 B.n39 163.367
R1689 B.n626 B.n39 163.367
R1690 B.n626 B.n625 163.367
R1691 B.n625 B.n624 163.367
R1692 B.n624 B.n41 163.367
R1693 B.n620 B.n41 163.367
R1694 B.n620 B.n619 163.367
R1695 B.n619 B.n618 163.367
R1696 B.n618 B.n43 163.367
R1697 B.n614 B.n43 163.367
R1698 B.n614 B.n613 163.367
R1699 B.n613 B.n612 163.367
R1700 B.n612 B.n45 163.367
R1701 B.n607 B.n45 163.367
R1702 B.n607 B.n606 163.367
R1703 B.n606 B.n605 163.367
R1704 B.n605 B.n49 163.367
R1705 B.n601 B.n49 163.367
R1706 B.n601 B.n600 163.367
R1707 B.n600 B.n599 163.367
R1708 B.n599 B.n51 163.367
R1709 B.n594 B.n51 163.367
R1710 B.n594 B.n593 163.367
R1711 B.n593 B.n592 163.367
R1712 B.n592 B.n55 163.367
R1713 B.n588 B.n55 163.367
R1714 B.n588 B.n587 163.367
R1715 B.n587 B.n586 163.367
R1716 B.n586 B.n57 163.367
R1717 B.n582 B.n57 163.367
R1718 B.n582 B.n581 163.367
R1719 B.n581 B.n580 163.367
R1720 B.n580 B.n59 163.367
R1721 B.n576 B.n59 163.367
R1722 B.n576 B.n575 163.367
R1723 B.n575 B.n574 163.367
R1724 B.n574 B.n61 163.367
R1725 B.n570 B.n61 163.367
R1726 B.n570 B.n569 163.367
R1727 B.n569 B.n568 163.367
R1728 B.n568 B.n63 163.367
R1729 B.n564 B.n63 163.367
R1730 B.n564 B.n563 163.367
R1731 B.n563 B.n562 163.367
R1732 B.n562 B.n65 163.367
R1733 B.n558 B.n65 163.367
R1734 B.n558 B.n557 163.367
R1735 B.n557 B.n556 163.367
R1736 B.n556 B.n67 163.367
R1737 B.n552 B.n67 163.367
R1738 B.n552 B.n551 163.367
R1739 B.n551 B.n550 163.367
R1740 B.n550 B.n69 163.367
R1741 B.n546 B.n69 163.367
R1742 B.n546 B.n545 163.367
R1743 B.n545 B.n544 163.367
R1744 B.n544 B.n71 163.367
R1745 B.n540 B.n71 163.367
R1746 B.n540 B.n539 163.367
R1747 B.n539 B.n538 163.367
R1748 B.n538 B.n73 163.367
R1749 B.n534 B.n73 163.367
R1750 B.n534 B.n533 163.367
R1751 B.n533 B.n532 163.367
R1752 B.n532 B.n75 163.367
R1753 B.n528 B.n75 163.367
R1754 B.n528 B.n527 163.367
R1755 B.n527 B.n526 163.367
R1756 B.n526 B.n77 163.367
R1757 B.n522 B.n77 163.367
R1758 B.n522 B.n521 163.367
R1759 B.n521 B.n520 163.367
R1760 B.n520 B.n79 163.367
R1761 B.n691 B.n690 163.367
R1762 B.n692 B.n691 163.367
R1763 B.n692 B.n17 163.367
R1764 B.n696 B.n17 163.367
R1765 B.n697 B.n696 163.367
R1766 B.n698 B.n697 163.367
R1767 B.n698 B.n15 163.367
R1768 B.n702 B.n15 163.367
R1769 B.n703 B.n702 163.367
R1770 B.n704 B.n703 163.367
R1771 B.n704 B.n13 163.367
R1772 B.n708 B.n13 163.367
R1773 B.n709 B.n708 163.367
R1774 B.n710 B.n709 163.367
R1775 B.n710 B.n11 163.367
R1776 B.n714 B.n11 163.367
R1777 B.n715 B.n714 163.367
R1778 B.n716 B.n715 163.367
R1779 B.n716 B.n9 163.367
R1780 B.n720 B.n9 163.367
R1781 B.n721 B.n720 163.367
R1782 B.n722 B.n721 163.367
R1783 B.n722 B.n7 163.367
R1784 B.n726 B.n7 163.367
R1785 B.n727 B.n726 163.367
R1786 B.n728 B.n727 163.367
R1787 B.n728 B.n5 163.367
R1788 B.n732 B.n5 163.367
R1789 B.n733 B.n732 163.367
R1790 B.n734 B.n733 163.367
R1791 B.n734 B.n3 163.367
R1792 B.n738 B.n3 163.367
R1793 B.n739 B.n738 163.367
R1794 B.n189 B.n2 163.367
R1795 B.n192 B.n189 163.367
R1796 B.n193 B.n192 163.367
R1797 B.n194 B.n193 163.367
R1798 B.n194 B.n187 163.367
R1799 B.n198 B.n187 163.367
R1800 B.n199 B.n198 163.367
R1801 B.n200 B.n199 163.367
R1802 B.n200 B.n185 163.367
R1803 B.n204 B.n185 163.367
R1804 B.n205 B.n204 163.367
R1805 B.n206 B.n205 163.367
R1806 B.n206 B.n183 163.367
R1807 B.n210 B.n183 163.367
R1808 B.n211 B.n210 163.367
R1809 B.n212 B.n211 163.367
R1810 B.n212 B.n181 163.367
R1811 B.n216 B.n181 163.367
R1812 B.n217 B.n216 163.367
R1813 B.n218 B.n217 163.367
R1814 B.n218 B.n179 163.367
R1815 B.n222 B.n179 163.367
R1816 B.n223 B.n222 163.367
R1817 B.n224 B.n223 163.367
R1818 B.n224 B.n177 163.367
R1819 B.n228 B.n177 163.367
R1820 B.n229 B.n228 163.367
R1821 B.n230 B.n229 163.367
R1822 B.n230 B.n175 163.367
R1823 B.n234 B.n175 163.367
R1824 B.n235 B.n234 163.367
R1825 B.n236 B.n235 163.367
R1826 B.n236 B.n173 163.367
R1827 B.n317 B.n147 59.5399
R1828 B.n332 B.n331 59.5399
R1829 B.n596 B.n53 59.5399
R1830 B.n610 B.n47 59.5399
R1831 B.n147 B.n146 57.9884
R1832 B.n331 B.n330 57.9884
R1833 B.n53 B.n52 57.9884
R1834 B.n47 B.n46 57.9884
R1835 B.n689 B.n688 34.1859
R1836 B.n518 B.n517 34.1859
R1837 B.n411 B.n114 34.1859
R1838 B.n239 B.n238 34.1859
R1839 B B.n741 18.0485
R1840 B.n689 B.n18 10.6151
R1841 B.n693 B.n18 10.6151
R1842 B.n694 B.n693 10.6151
R1843 B.n695 B.n694 10.6151
R1844 B.n695 B.n16 10.6151
R1845 B.n699 B.n16 10.6151
R1846 B.n700 B.n699 10.6151
R1847 B.n701 B.n700 10.6151
R1848 B.n701 B.n14 10.6151
R1849 B.n705 B.n14 10.6151
R1850 B.n706 B.n705 10.6151
R1851 B.n707 B.n706 10.6151
R1852 B.n707 B.n12 10.6151
R1853 B.n711 B.n12 10.6151
R1854 B.n712 B.n711 10.6151
R1855 B.n713 B.n712 10.6151
R1856 B.n713 B.n10 10.6151
R1857 B.n717 B.n10 10.6151
R1858 B.n718 B.n717 10.6151
R1859 B.n719 B.n718 10.6151
R1860 B.n719 B.n8 10.6151
R1861 B.n723 B.n8 10.6151
R1862 B.n724 B.n723 10.6151
R1863 B.n725 B.n724 10.6151
R1864 B.n725 B.n6 10.6151
R1865 B.n729 B.n6 10.6151
R1866 B.n730 B.n729 10.6151
R1867 B.n731 B.n730 10.6151
R1868 B.n731 B.n4 10.6151
R1869 B.n735 B.n4 10.6151
R1870 B.n736 B.n735 10.6151
R1871 B.n737 B.n736 10.6151
R1872 B.n737 B.n0 10.6151
R1873 B.n688 B.n687 10.6151
R1874 B.n687 B.n20 10.6151
R1875 B.n683 B.n20 10.6151
R1876 B.n683 B.n682 10.6151
R1877 B.n682 B.n681 10.6151
R1878 B.n681 B.n22 10.6151
R1879 B.n677 B.n22 10.6151
R1880 B.n677 B.n676 10.6151
R1881 B.n676 B.n675 10.6151
R1882 B.n675 B.n24 10.6151
R1883 B.n671 B.n24 10.6151
R1884 B.n671 B.n670 10.6151
R1885 B.n670 B.n669 10.6151
R1886 B.n669 B.n26 10.6151
R1887 B.n665 B.n26 10.6151
R1888 B.n665 B.n664 10.6151
R1889 B.n664 B.n663 10.6151
R1890 B.n663 B.n28 10.6151
R1891 B.n659 B.n28 10.6151
R1892 B.n659 B.n658 10.6151
R1893 B.n658 B.n657 10.6151
R1894 B.n657 B.n30 10.6151
R1895 B.n653 B.n30 10.6151
R1896 B.n653 B.n652 10.6151
R1897 B.n652 B.n651 10.6151
R1898 B.n651 B.n32 10.6151
R1899 B.n647 B.n32 10.6151
R1900 B.n647 B.n646 10.6151
R1901 B.n646 B.n645 10.6151
R1902 B.n645 B.n34 10.6151
R1903 B.n641 B.n34 10.6151
R1904 B.n641 B.n640 10.6151
R1905 B.n640 B.n639 10.6151
R1906 B.n639 B.n36 10.6151
R1907 B.n635 B.n36 10.6151
R1908 B.n635 B.n634 10.6151
R1909 B.n634 B.n633 10.6151
R1910 B.n633 B.n38 10.6151
R1911 B.n629 B.n38 10.6151
R1912 B.n629 B.n628 10.6151
R1913 B.n628 B.n627 10.6151
R1914 B.n627 B.n40 10.6151
R1915 B.n623 B.n40 10.6151
R1916 B.n623 B.n622 10.6151
R1917 B.n622 B.n621 10.6151
R1918 B.n621 B.n42 10.6151
R1919 B.n617 B.n42 10.6151
R1920 B.n617 B.n616 10.6151
R1921 B.n616 B.n615 10.6151
R1922 B.n615 B.n44 10.6151
R1923 B.n611 B.n44 10.6151
R1924 B.n609 B.n608 10.6151
R1925 B.n608 B.n48 10.6151
R1926 B.n604 B.n48 10.6151
R1927 B.n604 B.n603 10.6151
R1928 B.n603 B.n602 10.6151
R1929 B.n602 B.n50 10.6151
R1930 B.n598 B.n50 10.6151
R1931 B.n598 B.n597 10.6151
R1932 B.n595 B.n54 10.6151
R1933 B.n591 B.n54 10.6151
R1934 B.n591 B.n590 10.6151
R1935 B.n590 B.n589 10.6151
R1936 B.n589 B.n56 10.6151
R1937 B.n585 B.n56 10.6151
R1938 B.n585 B.n584 10.6151
R1939 B.n584 B.n583 10.6151
R1940 B.n583 B.n58 10.6151
R1941 B.n579 B.n58 10.6151
R1942 B.n579 B.n578 10.6151
R1943 B.n578 B.n577 10.6151
R1944 B.n577 B.n60 10.6151
R1945 B.n573 B.n60 10.6151
R1946 B.n573 B.n572 10.6151
R1947 B.n572 B.n571 10.6151
R1948 B.n571 B.n62 10.6151
R1949 B.n567 B.n62 10.6151
R1950 B.n567 B.n566 10.6151
R1951 B.n566 B.n565 10.6151
R1952 B.n565 B.n64 10.6151
R1953 B.n561 B.n64 10.6151
R1954 B.n561 B.n560 10.6151
R1955 B.n560 B.n559 10.6151
R1956 B.n559 B.n66 10.6151
R1957 B.n555 B.n66 10.6151
R1958 B.n555 B.n554 10.6151
R1959 B.n554 B.n553 10.6151
R1960 B.n553 B.n68 10.6151
R1961 B.n549 B.n68 10.6151
R1962 B.n549 B.n548 10.6151
R1963 B.n548 B.n547 10.6151
R1964 B.n547 B.n70 10.6151
R1965 B.n543 B.n70 10.6151
R1966 B.n543 B.n542 10.6151
R1967 B.n542 B.n541 10.6151
R1968 B.n541 B.n72 10.6151
R1969 B.n537 B.n72 10.6151
R1970 B.n537 B.n536 10.6151
R1971 B.n536 B.n535 10.6151
R1972 B.n535 B.n74 10.6151
R1973 B.n531 B.n74 10.6151
R1974 B.n531 B.n530 10.6151
R1975 B.n530 B.n529 10.6151
R1976 B.n529 B.n76 10.6151
R1977 B.n525 B.n76 10.6151
R1978 B.n525 B.n524 10.6151
R1979 B.n524 B.n523 10.6151
R1980 B.n523 B.n78 10.6151
R1981 B.n519 B.n78 10.6151
R1982 B.n519 B.n518 10.6151
R1983 B.n517 B.n80 10.6151
R1984 B.n513 B.n80 10.6151
R1985 B.n513 B.n512 10.6151
R1986 B.n512 B.n511 10.6151
R1987 B.n511 B.n82 10.6151
R1988 B.n507 B.n82 10.6151
R1989 B.n507 B.n506 10.6151
R1990 B.n506 B.n505 10.6151
R1991 B.n505 B.n84 10.6151
R1992 B.n501 B.n84 10.6151
R1993 B.n501 B.n500 10.6151
R1994 B.n500 B.n499 10.6151
R1995 B.n499 B.n86 10.6151
R1996 B.n495 B.n86 10.6151
R1997 B.n495 B.n494 10.6151
R1998 B.n494 B.n493 10.6151
R1999 B.n493 B.n88 10.6151
R2000 B.n489 B.n88 10.6151
R2001 B.n489 B.n488 10.6151
R2002 B.n488 B.n487 10.6151
R2003 B.n487 B.n90 10.6151
R2004 B.n483 B.n90 10.6151
R2005 B.n483 B.n482 10.6151
R2006 B.n482 B.n481 10.6151
R2007 B.n481 B.n92 10.6151
R2008 B.n477 B.n92 10.6151
R2009 B.n477 B.n476 10.6151
R2010 B.n476 B.n475 10.6151
R2011 B.n475 B.n94 10.6151
R2012 B.n471 B.n94 10.6151
R2013 B.n471 B.n470 10.6151
R2014 B.n470 B.n469 10.6151
R2015 B.n469 B.n96 10.6151
R2016 B.n465 B.n96 10.6151
R2017 B.n465 B.n464 10.6151
R2018 B.n464 B.n463 10.6151
R2019 B.n463 B.n98 10.6151
R2020 B.n459 B.n98 10.6151
R2021 B.n459 B.n458 10.6151
R2022 B.n458 B.n457 10.6151
R2023 B.n457 B.n100 10.6151
R2024 B.n453 B.n100 10.6151
R2025 B.n453 B.n452 10.6151
R2026 B.n452 B.n451 10.6151
R2027 B.n451 B.n102 10.6151
R2028 B.n447 B.n102 10.6151
R2029 B.n447 B.n446 10.6151
R2030 B.n446 B.n445 10.6151
R2031 B.n445 B.n104 10.6151
R2032 B.n441 B.n104 10.6151
R2033 B.n441 B.n440 10.6151
R2034 B.n440 B.n439 10.6151
R2035 B.n439 B.n106 10.6151
R2036 B.n435 B.n106 10.6151
R2037 B.n435 B.n434 10.6151
R2038 B.n434 B.n433 10.6151
R2039 B.n433 B.n108 10.6151
R2040 B.n429 B.n108 10.6151
R2041 B.n429 B.n428 10.6151
R2042 B.n428 B.n427 10.6151
R2043 B.n427 B.n110 10.6151
R2044 B.n423 B.n110 10.6151
R2045 B.n423 B.n422 10.6151
R2046 B.n422 B.n421 10.6151
R2047 B.n421 B.n112 10.6151
R2048 B.n417 B.n112 10.6151
R2049 B.n417 B.n416 10.6151
R2050 B.n416 B.n415 10.6151
R2051 B.n415 B.n114 10.6151
R2052 B.n190 B.n1 10.6151
R2053 B.n191 B.n190 10.6151
R2054 B.n191 B.n188 10.6151
R2055 B.n195 B.n188 10.6151
R2056 B.n196 B.n195 10.6151
R2057 B.n197 B.n196 10.6151
R2058 B.n197 B.n186 10.6151
R2059 B.n201 B.n186 10.6151
R2060 B.n202 B.n201 10.6151
R2061 B.n203 B.n202 10.6151
R2062 B.n203 B.n184 10.6151
R2063 B.n207 B.n184 10.6151
R2064 B.n208 B.n207 10.6151
R2065 B.n209 B.n208 10.6151
R2066 B.n209 B.n182 10.6151
R2067 B.n213 B.n182 10.6151
R2068 B.n214 B.n213 10.6151
R2069 B.n215 B.n214 10.6151
R2070 B.n215 B.n180 10.6151
R2071 B.n219 B.n180 10.6151
R2072 B.n220 B.n219 10.6151
R2073 B.n221 B.n220 10.6151
R2074 B.n221 B.n178 10.6151
R2075 B.n225 B.n178 10.6151
R2076 B.n226 B.n225 10.6151
R2077 B.n227 B.n226 10.6151
R2078 B.n227 B.n176 10.6151
R2079 B.n231 B.n176 10.6151
R2080 B.n232 B.n231 10.6151
R2081 B.n233 B.n232 10.6151
R2082 B.n233 B.n174 10.6151
R2083 B.n237 B.n174 10.6151
R2084 B.n238 B.n237 10.6151
R2085 B.n239 B.n172 10.6151
R2086 B.n243 B.n172 10.6151
R2087 B.n244 B.n243 10.6151
R2088 B.n245 B.n244 10.6151
R2089 B.n245 B.n170 10.6151
R2090 B.n249 B.n170 10.6151
R2091 B.n250 B.n249 10.6151
R2092 B.n251 B.n250 10.6151
R2093 B.n251 B.n168 10.6151
R2094 B.n255 B.n168 10.6151
R2095 B.n256 B.n255 10.6151
R2096 B.n257 B.n256 10.6151
R2097 B.n257 B.n166 10.6151
R2098 B.n261 B.n166 10.6151
R2099 B.n262 B.n261 10.6151
R2100 B.n263 B.n262 10.6151
R2101 B.n263 B.n164 10.6151
R2102 B.n267 B.n164 10.6151
R2103 B.n268 B.n267 10.6151
R2104 B.n269 B.n268 10.6151
R2105 B.n269 B.n162 10.6151
R2106 B.n273 B.n162 10.6151
R2107 B.n274 B.n273 10.6151
R2108 B.n275 B.n274 10.6151
R2109 B.n275 B.n160 10.6151
R2110 B.n279 B.n160 10.6151
R2111 B.n280 B.n279 10.6151
R2112 B.n281 B.n280 10.6151
R2113 B.n281 B.n158 10.6151
R2114 B.n285 B.n158 10.6151
R2115 B.n286 B.n285 10.6151
R2116 B.n287 B.n286 10.6151
R2117 B.n287 B.n156 10.6151
R2118 B.n291 B.n156 10.6151
R2119 B.n292 B.n291 10.6151
R2120 B.n293 B.n292 10.6151
R2121 B.n293 B.n154 10.6151
R2122 B.n297 B.n154 10.6151
R2123 B.n298 B.n297 10.6151
R2124 B.n299 B.n298 10.6151
R2125 B.n299 B.n152 10.6151
R2126 B.n303 B.n152 10.6151
R2127 B.n304 B.n303 10.6151
R2128 B.n305 B.n304 10.6151
R2129 B.n305 B.n150 10.6151
R2130 B.n309 B.n150 10.6151
R2131 B.n310 B.n309 10.6151
R2132 B.n311 B.n310 10.6151
R2133 B.n311 B.n148 10.6151
R2134 B.n315 B.n148 10.6151
R2135 B.n316 B.n315 10.6151
R2136 B.n318 B.n144 10.6151
R2137 B.n322 B.n144 10.6151
R2138 B.n323 B.n322 10.6151
R2139 B.n324 B.n323 10.6151
R2140 B.n324 B.n142 10.6151
R2141 B.n328 B.n142 10.6151
R2142 B.n329 B.n328 10.6151
R2143 B.n333 B.n329 10.6151
R2144 B.n337 B.n140 10.6151
R2145 B.n338 B.n337 10.6151
R2146 B.n339 B.n338 10.6151
R2147 B.n339 B.n138 10.6151
R2148 B.n343 B.n138 10.6151
R2149 B.n344 B.n343 10.6151
R2150 B.n345 B.n344 10.6151
R2151 B.n345 B.n136 10.6151
R2152 B.n349 B.n136 10.6151
R2153 B.n350 B.n349 10.6151
R2154 B.n351 B.n350 10.6151
R2155 B.n351 B.n134 10.6151
R2156 B.n355 B.n134 10.6151
R2157 B.n356 B.n355 10.6151
R2158 B.n357 B.n356 10.6151
R2159 B.n357 B.n132 10.6151
R2160 B.n361 B.n132 10.6151
R2161 B.n362 B.n361 10.6151
R2162 B.n363 B.n362 10.6151
R2163 B.n363 B.n130 10.6151
R2164 B.n367 B.n130 10.6151
R2165 B.n368 B.n367 10.6151
R2166 B.n369 B.n368 10.6151
R2167 B.n369 B.n128 10.6151
R2168 B.n373 B.n128 10.6151
R2169 B.n374 B.n373 10.6151
R2170 B.n375 B.n374 10.6151
R2171 B.n375 B.n126 10.6151
R2172 B.n379 B.n126 10.6151
R2173 B.n380 B.n379 10.6151
R2174 B.n381 B.n380 10.6151
R2175 B.n381 B.n124 10.6151
R2176 B.n385 B.n124 10.6151
R2177 B.n386 B.n385 10.6151
R2178 B.n387 B.n386 10.6151
R2179 B.n387 B.n122 10.6151
R2180 B.n391 B.n122 10.6151
R2181 B.n392 B.n391 10.6151
R2182 B.n393 B.n392 10.6151
R2183 B.n393 B.n120 10.6151
R2184 B.n397 B.n120 10.6151
R2185 B.n398 B.n397 10.6151
R2186 B.n399 B.n398 10.6151
R2187 B.n399 B.n118 10.6151
R2188 B.n403 B.n118 10.6151
R2189 B.n404 B.n403 10.6151
R2190 B.n405 B.n404 10.6151
R2191 B.n405 B.n116 10.6151
R2192 B.n409 B.n116 10.6151
R2193 B.n410 B.n409 10.6151
R2194 B.n411 B.n410 10.6151
R2195 B.n741 B.n0 8.11757
R2196 B.n741 B.n1 8.11757
R2197 B.n610 B.n609 6.5566
R2198 B.n597 B.n596 6.5566
R2199 B.n318 B.n317 6.5566
R2200 B.n333 B.n332 6.5566
R2201 B.n611 B.n610 4.05904
R2202 B.n596 B.n595 4.05904
R2203 B.n317 B.n316 4.05904
R2204 B.n332 B.n140 4.05904
C0 VP VDD1 6.31777f
C1 VN VDD2 6.06945f
C2 VTAIL VDD1 6.24021f
C3 w_n2764_n4066# VDD2 1.61336f
C4 B VDD1 1.3655f
C5 VP VDD2 0.397959f
C6 VTAIL VDD2 6.29481f
C7 w_n2764_n4066# VN 4.77133f
C8 B VDD2 1.41863f
C9 VP VN 6.88508f
C10 VDD1 VDD2 1.03371f
C11 VN VTAIL 5.82642f
C12 w_n2764_n4066# VP 5.12681f
C13 w_n2764_n4066# VTAIL 4.75914f
C14 B VN 1.16103f
C15 VN VDD1 0.14889f
C16 w_n2764_n4066# B 10.298599f
C17 VP VTAIL 5.84053f
C18 w_n2764_n4066# VDD1 1.55591f
C19 B VP 1.7512f
C20 B VTAIL 6.12289f
C21 VDD2 VSUBS 1.046949f
C22 VDD1 VSUBS 6.18916f
C23 VTAIL VSUBS 1.385032f
C24 VN VSUBS 5.60431f
C25 VP VSUBS 2.45782f
C26 B VSUBS 4.623542f
C27 w_n2764_n4066# VSUBS 0.137747p
C28 B.n0 VSUBS 0.0055f
C29 B.n1 VSUBS 0.0055f
C30 B.n2 VSUBS 0.008134f
C31 B.n3 VSUBS 0.006233f
C32 B.n4 VSUBS 0.006233f
C33 B.n5 VSUBS 0.006233f
C34 B.n6 VSUBS 0.006233f
C35 B.n7 VSUBS 0.006233f
C36 B.n8 VSUBS 0.006233f
C37 B.n9 VSUBS 0.006233f
C38 B.n10 VSUBS 0.006233f
C39 B.n11 VSUBS 0.006233f
C40 B.n12 VSUBS 0.006233f
C41 B.n13 VSUBS 0.006233f
C42 B.n14 VSUBS 0.006233f
C43 B.n15 VSUBS 0.006233f
C44 B.n16 VSUBS 0.006233f
C45 B.n17 VSUBS 0.006233f
C46 B.n18 VSUBS 0.006233f
C47 B.n19 VSUBS 0.015265f
C48 B.n20 VSUBS 0.006233f
C49 B.n21 VSUBS 0.006233f
C50 B.n22 VSUBS 0.006233f
C51 B.n23 VSUBS 0.006233f
C52 B.n24 VSUBS 0.006233f
C53 B.n25 VSUBS 0.006233f
C54 B.n26 VSUBS 0.006233f
C55 B.n27 VSUBS 0.006233f
C56 B.n28 VSUBS 0.006233f
C57 B.n29 VSUBS 0.006233f
C58 B.n30 VSUBS 0.006233f
C59 B.n31 VSUBS 0.006233f
C60 B.n32 VSUBS 0.006233f
C61 B.n33 VSUBS 0.006233f
C62 B.n34 VSUBS 0.006233f
C63 B.n35 VSUBS 0.006233f
C64 B.n36 VSUBS 0.006233f
C65 B.n37 VSUBS 0.006233f
C66 B.n38 VSUBS 0.006233f
C67 B.n39 VSUBS 0.006233f
C68 B.n40 VSUBS 0.006233f
C69 B.n41 VSUBS 0.006233f
C70 B.n42 VSUBS 0.006233f
C71 B.n43 VSUBS 0.006233f
C72 B.n44 VSUBS 0.006233f
C73 B.n45 VSUBS 0.006233f
C74 B.t4 VSUBS 0.259266f
C75 B.t5 VSUBS 0.289234f
C76 B.t3 VSUBS 1.64675f
C77 B.n46 VSUBS 0.449238f
C78 B.n47 VSUBS 0.265484f
C79 B.n48 VSUBS 0.006233f
C80 B.n49 VSUBS 0.006233f
C81 B.n50 VSUBS 0.006233f
C82 B.n51 VSUBS 0.006233f
C83 B.t1 VSUBS 0.259269f
C84 B.t2 VSUBS 0.289237f
C85 B.t0 VSUBS 1.64675f
C86 B.n52 VSUBS 0.449235f
C87 B.n53 VSUBS 0.265481f
C88 B.n54 VSUBS 0.006233f
C89 B.n55 VSUBS 0.006233f
C90 B.n56 VSUBS 0.006233f
C91 B.n57 VSUBS 0.006233f
C92 B.n58 VSUBS 0.006233f
C93 B.n59 VSUBS 0.006233f
C94 B.n60 VSUBS 0.006233f
C95 B.n61 VSUBS 0.006233f
C96 B.n62 VSUBS 0.006233f
C97 B.n63 VSUBS 0.006233f
C98 B.n64 VSUBS 0.006233f
C99 B.n65 VSUBS 0.006233f
C100 B.n66 VSUBS 0.006233f
C101 B.n67 VSUBS 0.006233f
C102 B.n68 VSUBS 0.006233f
C103 B.n69 VSUBS 0.006233f
C104 B.n70 VSUBS 0.006233f
C105 B.n71 VSUBS 0.006233f
C106 B.n72 VSUBS 0.006233f
C107 B.n73 VSUBS 0.006233f
C108 B.n74 VSUBS 0.006233f
C109 B.n75 VSUBS 0.006233f
C110 B.n76 VSUBS 0.006233f
C111 B.n77 VSUBS 0.006233f
C112 B.n78 VSUBS 0.006233f
C113 B.n79 VSUBS 0.015265f
C114 B.n80 VSUBS 0.006233f
C115 B.n81 VSUBS 0.006233f
C116 B.n82 VSUBS 0.006233f
C117 B.n83 VSUBS 0.006233f
C118 B.n84 VSUBS 0.006233f
C119 B.n85 VSUBS 0.006233f
C120 B.n86 VSUBS 0.006233f
C121 B.n87 VSUBS 0.006233f
C122 B.n88 VSUBS 0.006233f
C123 B.n89 VSUBS 0.006233f
C124 B.n90 VSUBS 0.006233f
C125 B.n91 VSUBS 0.006233f
C126 B.n92 VSUBS 0.006233f
C127 B.n93 VSUBS 0.006233f
C128 B.n94 VSUBS 0.006233f
C129 B.n95 VSUBS 0.006233f
C130 B.n96 VSUBS 0.006233f
C131 B.n97 VSUBS 0.006233f
C132 B.n98 VSUBS 0.006233f
C133 B.n99 VSUBS 0.006233f
C134 B.n100 VSUBS 0.006233f
C135 B.n101 VSUBS 0.006233f
C136 B.n102 VSUBS 0.006233f
C137 B.n103 VSUBS 0.006233f
C138 B.n104 VSUBS 0.006233f
C139 B.n105 VSUBS 0.006233f
C140 B.n106 VSUBS 0.006233f
C141 B.n107 VSUBS 0.006233f
C142 B.n108 VSUBS 0.006233f
C143 B.n109 VSUBS 0.006233f
C144 B.n110 VSUBS 0.006233f
C145 B.n111 VSUBS 0.006233f
C146 B.n112 VSUBS 0.006233f
C147 B.n113 VSUBS 0.006233f
C148 B.n114 VSUBS 0.015505f
C149 B.n115 VSUBS 0.006233f
C150 B.n116 VSUBS 0.006233f
C151 B.n117 VSUBS 0.006233f
C152 B.n118 VSUBS 0.006233f
C153 B.n119 VSUBS 0.006233f
C154 B.n120 VSUBS 0.006233f
C155 B.n121 VSUBS 0.006233f
C156 B.n122 VSUBS 0.006233f
C157 B.n123 VSUBS 0.006233f
C158 B.n124 VSUBS 0.006233f
C159 B.n125 VSUBS 0.006233f
C160 B.n126 VSUBS 0.006233f
C161 B.n127 VSUBS 0.006233f
C162 B.n128 VSUBS 0.006233f
C163 B.n129 VSUBS 0.006233f
C164 B.n130 VSUBS 0.006233f
C165 B.n131 VSUBS 0.006233f
C166 B.n132 VSUBS 0.006233f
C167 B.n133 VSUBS 0.006233f
C168 B.n134 VSUBS 0.006233f
C169 B.n135 VSUBS 0.006233f
C170 B.n136 VSUBS 0.006233f
C171 B.n137 VSUBS 0.006233f
C172 B.n138 VSUBS 0.006233f
C173 B.n139 VSUBS 0.006233f
C174 B.n140 VSUBS 0.004308f
C175 B.n141 VSUBS 0.006233f
C176 B.n142 VSUBS 0.006233f
C177 B.n143 VSUBS 0.006233f
C178 B.n144 VSUBS 0.006233f
C179 B.n145 VSUBS 0.006233f
C180 B.t11 VSUBS 0.259266f
C181 B.t10 VSUBS 0.289234f
C182 B.t9 VSUBS 1.64675f
C183 B.n146 VSUBS 0.449238f
C184 B.n147 VSUBS 0.265484f
C185 B.n148 VSUBS 0.006233f
C186 B.n149 VSUBS 0.006233f
C187 B.n150 VSUBS 0.006233f
C188 B.n151 VSUBS 0.006233f
C189 B.n152 VSUBS 0.006233f
C190 B.n153 VSUBS 0.006233f
C191 B.n154 VSUBS 0.006233f
C192 B.n155 VSUBS 0.006233f
C193 B.n156 VSUBS 0.006233f
C194 B.n157 VSUBS 0.006233f
C195 B.n158 VSUBS 0.006233f
C196 B.n159 VSUBS 0.006233f
C197 B.n160 VSUBS 0.006233f
C198 B.n161 VSUBS 0.006233f
C199 B.n162 VSUBS 0.006233f
C200 B.n163 VSUBS 0.006233f
C201 B.n164 VSUBS 0.006233f
C202 B.n165 VSUBS 0.006233f
C203 B.n166 VSUBS 0.006233f
C204 B.n167 VSUBS 0.006233f
C205 B.n168 VSUBS 0.006233f
C206 B.n169 VSUBS 0.006233f
C207 B.n170 VSUBS 0.006233f
C208 B.n171 VSUBS 0.006233f
C209 B.n172 VSUBS 0.006233f
C210 B.n173 VSUBS 0.014802f
C211 B.n174 VSUBS 0.006233f
C212 B.n175 VSUBS 0.006233f
C213 B.n176 VSUBS 0.006233f
C214 B.n177 VSUBS 0.006233f
C215 B.n178 VSUBS 0.006233f
C216 B.n179 VSUBS 0.006233f
C217 B.n180 VSUBS 0.006233f
C218 B.n181 VSUBS 0.006233f
C219 B.n182 VSUBS 0.006233f
C220 B.n183 VSUBS 0.006233f
C221 B.n184 VSUBS 0.006233f
C222 B.n185 VSUBS 0.006233f
C223 B.n186 VSUBS 0.006233f
C224 B.n187 VSUBS 0.006233f
C225 B.n188 VSUBS 0.006233f
C226 B.n189 VSUBS 0.006233f
C227 B.n190 VSUBS 0.006233f
C228 B.n191 VSUBS 0.006233f
C229 B.n192 VSUBS 0.006233f
C230 B.n193 VSUBS 0.006233f
C231 B.n194 VSUBS 0.006233f
C232 B.n195 VSUBS 0.006233f
C233 B.n196 VSUBS 0.006233f
C234 B.n197 VSUBS 0.006233f
C235 B.n198 VSUBS 0.006233f
C236 B.n199 VSUBS 0.006233f
C237 B.n200 VSUBS 0.006233f
C238 B.n201 VSUBS 0.006233f
C239 B.n202 VSUBS 0.006233f
C240 B.n203 VSUBS 0.006233f
C241 B.n204 VSUBS 0.006233f
C242 B.n205 VSUBS 0.006233f
C243 B.n206 VSUBS 0.006233f
C244 B.n207 VSUBS 0.006233f
C245 B.n208 VSUBS 0.006233f
C246 B.n209 VSUBS 0.006233f
C247 B.n210 VSUBS 0.006233f
C248 B.n211 VSUBS 0.006233f
C249 B.n212 VSUBS 0.006233f
C250 B.n213 VSUBS 0.006233f
C251 B.n214 VSUBS 0.006233f
C252 B.n215 VSUBS 0.006233f
C253 B.n216 VSUBS 0.006233f
C254 B.n217 VSUBS 0.006233f
C255 B.n218 VSUBS 0.006233f
C256 B.n219 VSUBS 0.006233f
C257 B.n220 VSUBS 0.006233f
C258 B.n221 VSUBS 0.006233f
C259 B.n222 VSUBS 0.006233f
C260 B.n223 VSUBS 0.006233f
C261 B.n224 VSUBS 0.006233f
C262 B.n225 VSUBS 0.006233f
C263 B.n226 VSUBS 0.006233f
C264 B.n227 VSUBS 0.006233f
C265 B.n228 VSUBS 0.006233f
C266 B.n229 VSUBS 0.006233f
C267 B.n230 VSUBS 0.006233f
C268 B.n231 VSUBS 0.006233f
C269 B.n232 VSUBS 0.006233f
C270 B.n233 VSUBS 0.006233f
C271 B.n234 VSUBS 0.006233f
C272 B.n235 VSUBS 0.006233f
C273 B.n236 VSUBS 0.006233f
C274 B.n237 VSUBS 0.006233f
C275 B.n238 VSUBS 0.014802f
C276 B.n239 VSUBS 0.015265f
C277 B.n240 VSUBS 0.015265f
C278 B.n241 VSUBS 0.006233f
C279 B.n242 VSUBS 0.006233f
C280 B.n243 VSUBS 0.006233f
C281 B.n244 VSUBS 0.006233f
C282 B.n245 VSUBS 0.006233f
C283 B.n246 VSUBS 0.006233f
C284 B.n247 VSUBS 0.006233f
C285 B.n248 VSUBS 0.006233f
C286 B.n249 VSUBS 0.006233f
C287 B.n250 VSUBS 0.006233f
C288 B.n251 VSUBS 0.006233f
C289 B.n252 VSUBS 0.006233f
C290 B.n253 VSUBS 0.006233f
C291 B.n254 VSUBS 0.006233f
C292 B.n255 VSUBS 0.006233f
C293 B.n256 VSUBS 0.006233f
C294 B.n257 VSUBS 0.006233f
C295 B.n258 VSUBS 0.006233f
C296 B.n259 VSUBS 0.006233f
C297 B.n260 VSUBS 0.006233f
C298 B.n261 VSUBS 0.006233f
C299 B.n262 VSUBS 0.006233f
C300 B.n263 VSUBS 0.006233f
C301 B.n264 VSUBS 0.006233f
C302 B.n265 VSUBS 0.006233f
C303 B.n266 VSUBS 0.006233f
C304 B.n267 VSUBS 0.006233f
C305 B.n268 VSUBS 0.006233f
C306 B.n269 VSUBS 0.006233f
C307 B.n270 VSUBS 0.006233f
C308 B.n271 VSUBS 0.006233f
C309 B.n272 VSUBS 0.006233f
C310 B.n273 VSUBS 0.006233f
C311 B.n274 VSUBS 0.006233f
C312 B.n275 VSUBS 0.006233f
C313 B.n276 VSUBS 0.006233f
C314 B.n277 VSUBS 0.006233f
C315 B.n278 VSUBS 0.006233f
C316 B.n279 VSUBS 0.006233f
C317 B.n280 VSUBS 0.006233f
C318 B.n281 VSUBS 0.006233f
C319 B.n282 VSUBS 0.006233f
C320 B.n283 VSUBS 0.006233f
C321 B.n284 VSUBS 0.006233f
C322 B.n285 VSUBS 0.006233f
C323 B.n286 VSUBS 0.006233f
C324 B.n287 VSUBS 0.006233f
C325 B.n288 VSUBS 0.006233f
C326 B.n289 VSUBS 0.006233f
C327 B.n290 VSUBS 0.006233f
C328 B.n291 VSUBS 0.006233f
C329 B.n292 VSUBS 0.006233f
C330 B.n293 VSUBS 0.006233f
C331 B.n294 VSUBS 0.006233f
C332 B.n295 VSUBS 0.006233f
C333 B.n296 VSUBS 0.006233f
C334 B.n297 VSUBS 0.006233f
C335 B.n298 VSUBS 0.006233f
C336 B.n299 VSUBS 0.006233f
C337 B.n300 VSUBS 0.006233f
C338 B.n301 VSUBS 0.006233f
C339 B.n302 VSUBS 0.006233f
C340 B.n303 VSUBS 0.006233f
C341 B.n304 VSUBS 0.006233f
C342 B.n305 VSUBS 0.006233f
C343 B.n306 VSUBS 0.006233f
C344 B.n307 VSUBS 0.006233f
C345 B.n308 VSUBS 0.006233f
C346 B.n309 VSUBS 0.006233f
C347 B.n310 VSUBS 0.006233f
C348 B.n311 VSUBS 0.006233f
C349 B.n312 VSUBS 0.006233f
C350 B.n313 VSUBS 0.006233f
C351 B.n314 VSUBS 0.006233f
C352 B.n315 VSUBS 0.006233f
C353 B.n316 VSUBS 0.004308f
C354 B.n317 VSUBS 0.014442f
C355 B.n318 VSUBS 0.005042f
C356 B.n319 VSUBS 0.006233f
C357 B.n320 VSUBS 0.006233f
C358 B.n321 VSUBS 0.006233f
C359 B.n322 VSUBS 0.006233f
C360 B.n323 VSUBS 0.006233f
C361 B.n324 VSUBS 0.006233f
C362 B.n325 VSUBS 0.006233f
C363 B.n326 VSUBS 0.006233f
C364 B.n327 VSUBS 0.006233f
C365 B.n328 VSUBS 0.006233f
C366 B.n329 VSUBS 0.006233f
C367 B.t8 VSUBS 0.259269f
C368 B.t7 VSUBS 0.289237f
C369 B.t6 VSUBS 1.64675f
C370 B.n330 VSUBS 0.449235f
C371 B.n331 VSUBS 0.265481f
C372 B.n332 VSUBS 0.014442f
C373 B.n333 VSUBS 0.005042f
C374 B.n334 VSUBS 0.006233f
C375 B.n335 VSUBS 0.006233f
C376 B.n336 VSUBS 0.006233f
C377 B.n337 VSUBS 0.006233f
C378 B.n338 VSUBS 0.006233f
C379 B.n339 VSUBS 0.006233f
C380 B.n340 VSUBS 0.006233f
C381 B.n341 VSUBS 0.006233f
C382 B.n342 VSUBS 0.006233f
C383 B.n343 VSUBS 0.006233f
C384 B.n344 VSUBS 0.006233f
C385 B.n345 VSUBS 0.006233f
C386 B.n346 VSUBS 0.006233f
C387 B.n347 VSUBS 0.006233f
C388 B.n348 VSUBS 0.006233f
C389 B.n349 VSUBS 0.006233f
C390 B.n350 VSUBS 0.006233f
C391 B.n351 VSUBS 0.006233f
C392 B.n352 VSUBS 0.006233f
C393 B.n353 VSUBS 0.006233f
C394 B.n354 VSUBS 0.006233f
C395 B.n355 VSUBS 0.006233f
C396 B.n356 VSUBS 0.006233f
C397 B.n357 VSUBS 0.006233f
C398 B.n358 VSUBS 0.006233f
C399 B.n359 VSUBS 0.006233f
C400 B.n360 VSUBS 0.006233f
C401 B.n361 VSUBS 0.006233f
C402 B.n362 VSUBS 0.006233f
C403 B.n363 VSUBS 0.006233f
C404 B.n364 VSUBS 0.006233f
C405 B.n365 VSUBS 0.006233f
C406 B.n366 VSUBS 0.006233f
C407 B.n367 VSUBS 0.006233f
C408 B.n368 VSUBS 0.006233f
C409 B.n369 VSUBS 0.006233f
C410 B.n370 VSUBS 0.006233f
C411 B.n371 VSUBS 0.006233f
C412 B.n372 VSUBS 0.006233f
C413 B.n373 VSUBS 0.006233f
C414 B.n374 VSUBS 0.006233f
C415 B.n375 VSUBS 0.006233f
C416 B.n376 VSUBS 0.006233f
C417 B.n377 VSUBS 0.006233f
C418 B.n378 VSUBS 0.006233f
C419 B.n379 VSUBS 0.006233f
C420 B.n380 VSUBS 0.006233f
C421 B.n381 VSUBS 0.006233f
C422 B.n382 VSUBS 0.006233f
C423 B.n383 VSUBS 0.006233f
C424 B.n384 VSUBS 0.006233f
C425 B.n385 VSUBS 0.006233f
C426 B.n386 VSUBS 0.006233f
C427 B.n387 VSUBS 0.006233f
C428 B.n388 VSUBS 0.006233f
C429 B.n389 VSUBS 0.006233f
C430 B.n390 VSUBS 0.006233f
C431 B.n391 VSUBS 0.006233f
C432 B.n392 VSUBS 0.006233f
C433 B.n393 VSUBS 0.006233f
C434 B.n394 VSUBS 0.006233f
C435 B.n395 VSUBS 0.006233f
C436 B.n396 VSUBS 0.006233f
C437 B.n397 VSUBS 0.006233f
C438 B.n398 VSUBS 0.006233f
C439 B.n399 VSUBS 0.006233f
C440 B.n400 VSUBS 0.006233f
C441 B.n401 VSUBS 0.006233f
C442 B.n402 VSUBS 0.006233f
C443 B.n403 VSUBS 0.006233f
C444 B.n404 VSUBS 0.006233f
C445 B.n405 VSUBS 0.006233f
C446 B.n406 VSUBS 0.006233f
C447 B.n407 VSUBS 0.006233f
C448 B.n408 VSUBS 0.006233f
C449 B.n409 VSUBS 0.006233f
C450 B.n410 VSUBS 0.006233f
C451 B.n411 VSUBS 0.014561f
C452 B.n412 VSUBS 0.015265f
C453 B.n413 VSUBS 0.014802f
C454 B.n414 VSUBS 0.006233f
C455 B.n415 VSUBS 0.006233f
C456 B.n416 VSUBS 0.006233f
C457 B.n417 VSUBS 0.006233f
C458 B.n418 VSUBS 0.006233f
C459 B.n419 VSUBS 0.006233f
C460 B.n420 VSUBS 0.006233f
C461 B.n421 VSUBS 0.006233f
C462 B.n422 VSUBS 0.006233f
C463 B.n423 VSUBS 0.006233f
C464 B.n424 VSUBS 0.006233f
C465 B.n425 VSUBS 0.006233f
C466 B.n426 VSUBS 0.006233f
C467 B.n427 VSUBS 0.006233f
C468 B.n428 VSUBS 0.006233f
C469 B.n429 VSUBS 0.006233f
C470 B.n430 VSUBS 0.006233f
C471 B.n431 VSUBS 0.006233f
C472 B.n432 VSUBS 0.006233f
C473 B.n433 VSUBS 0.006233f
C474 B.n434 VSUBS 0.006233f
C475 B.n435 VSUBS 0.006233f
C476 B.n436 VSUBS 0.006233f
C477 B.n437 VSUBS 0.006233f
C478 B.n438 VSUBS 0.006233f
C479 B.n439 VSUBS 0.006233f
C480 B.n440 VSUBS 0.006233f
C481 B.n441 VSUBS 0.006233f
C482 B.n442 VSUBS 0.006233f
C483 B.n443 VSUBS 0.006233f
C484 B.n444 VSUBS 0.006233f
C485 B.n445 VSUBS 0.006233f
C486 B.n446 VSUBS 0.006233f
C487 B.n447 VSUBS 0.006233f
C488 B.n448 VSUBS 0.006233f
C489 B.n449 VSUBS 0.006233f
C490 B.n450 VSUBS 0.006233f
C491 B.n451 VSUBS 0.006233f
C492 B.n452 VSUBS 0.006233f
C493 B.n453 VSUBS 0.006233f
C494 B.n454 VSUBS 0.006233f
C495 B.n455 VSUBS 0.006233f
C496 B.n456 VSUBS 0.006233f
C497 B.n457 VSUBS 0.006233f
C498 B.n458 VSUBS 0.006233f
C499 B.n459 VSUBS 0.006233f
C500 B.n460 VSUBS 0.006233f
C501 B.n461 VSUBS 0.006233f
C502 B.n462 VSUBS 0.006233f
C503 B.n463 VSUBS 0.006233f
C504 B.n464 VSUBS 0.006233f
C505 B.n465 VSUBS 0.006233f
C506 B.n466 VSUBS 0.006233f
C507 B.n467 VSUBS 0.006233f
C508 B.n468 VSUBS 0.006233f
C509 B.n469 VSUBS 0.006233f
C510 B.n470 VSUBS 0.006233f
C511 B.n471 VSUBS 0.006233f
C512 B.n472 VSUBS 0.006233f
C513 B.n473 VSUBS 0.006233f
C514 B.n474 VSUBS 0.006233f
C515 B.n475 VSUBS 0.006233f
C516 B.n476 VSUBS 0.006233f
C517 B.n477 VSUBS 0.006233f
C518 B.n478 VSUBS 0.006233f
C519 B.n479 VSUBS 0.006233f
C520 B.n480 VSUBS 0.006233f
C521 B.n481 VSUBS 0.006233f
C522 B.n482 VSUBS 0.006233f
C523 B.n483 VSUBS 0.006233f
C524 B.n484 VSUBS 0.006233f
C525 B.n485 VSUBS 0.006233f
C526 B.n486 VSUBS 0.006233f
C527 B.n487 VSUBS 0.006233f
C528 B.n488 VSUBS 0.006233f
C529 B.n489 VSUBS 0.006233f
C530 B.n490 VSUBS 0.006233f
C531 B.n491 VSUBS 0.006233f
C532 B.n492 VSUBS 0.006233f
C533 B.n493 VSUBS 0.006233f
C534 B.n494 VSUBS 0.006233f
C535 B.n495 VSUBS 0.006233f
C536 B.n496 VSUBS 0.006233f
C537 B.n497 VSUBS 0.006233f
C538 B.n498 VSUBS 0.006233f
C539 B.n499 VSUBS 0.006233f
C540 B.n500 VSUBS 0.006233f
C541 B.n501 VSUBS 0.006233f
C542 B.n502 VSUBS 0.006233f
C543 B.n503 VSUBS 0.006233f
C544 B.n504 VSUBS 0.006233f
C545 B.n505 VSUBS 0.006233f
C546 B.n506 VSUBS 0.006233f
C547 B.n507 VSUBS 0.006233f
C548 B.n508 VSUBS 0.006233f
C549 B.n509 VSUBS 0.006233f
C550 B.n510 VSUBS 0.006233f
C551 B.n511 VSUBS 0.006233f
C552 B.n512 VSUBS 0.006233f
C553 B.n513 VSUBS 0.006233f
C554 B.n514 VSUBS 0.006233f
C555 B.n515 VSUBS 0.006233f
C556 B.n516 VSUBS 0.014802f
C557 B.n517 VSUBS 0.014802f
C558 B.n518 VSUBS 0.015265f
C559 B.n519 VSUBS 0.006233f
C560 B.n520 VSUBS 0.006233f
C561 B.n521 VSUBS 0.006233f
C562 B.n522 VSUBS 0.006233f
C563 B.n523 VSUBS 0.006233f
C564 B.n524 VSUBS 0.006233f
C565 B.n525 VSUBS 0.006233f
C566 B.n526 VSUBS 0.006233f
C567 B.n527 VSUBS 0.006233f
C568 B.n528 VSUBS 0.006233f
C569 B.n529 VSUBS 0.006233f
C570 B.n530 VSUBS 0.006233f
C571 B.n531 VSUBS 0.006233f
C572 B.n532 VSUBS 0.006233f
C573 B.n533 VSUBS 0.006233f
C574 B.n534 VSUBS 0.006233f
C575 B.n535 VSUBS 0.006233f
C576 B.n536 VSUBS 0.006233f
C577 B.n537 VSUBS 0.006233f
C578 B.n538 VSUBS 0.006233f
C579 B.n539 VSUBS 0.006233f
C580 B.n540 VSUBS 0.006233f
C581 B.n541 VSUBS 0.006233f
C582 B.n542 VSUBS 0.006233f
C583 B.n543 VSUBS 0.006233f
C584 B.n544 VSUBS 0.006233f
C585 B.n545 VSUBS 0.006233f
C586 B.n546 VSUBS 0.006233f
C587 B.n547 VSUBS 0.006233f
C588 B.n548 VSUBS 0.006233f
C589 B.n549 VSUBS 0.006233f
C590 B.n550 VSUBS 0.006233f
C591 B.n551 VSUBS 0.006233f
C592 B.n552 VSUBS 0.006233f
C593 B.n553 VSUBS 0.006233f
C594 B.n554 VSUBS 0.006233f
C595 B.n555 VSUBS 0.006233f
C596 B.n556 VSUBS 0.006233f
C597 B.n557 VSUBS 0.006233f
C598 B.n558 VSUBS 0.006233f
C599 B.n559 VSUBS 0.006233f
C600 B.n560 VSUBS 0.006233f
C601 B.n561 VSUBS 0.006233f
C602 B.n562 VSUBS 0.006233f
C603 B.n563 VSUBS 0.006233f
C604 B.n564 VSUBS 0.006233f
C605 B.n565 VSUBS 0.006233f
C606 B.n566 VSUBS 0.006233f
C607 B.n567 VSUBS 0.006233f
C608 B.n568 VSUBS 0.006233f
C609 B.n569 VSUBS 0.006233f
C610 B.n570 VSUBS 0.006233f
C611 B.n571 VSUBS 0.006233f
C612 B.n572 VSUBS 0.006233f
C613 B.n573 VSUBS 0.006233f
C614 B.n574 VSUBS 0.006233f
C615 B.n575 VSUBS 0.006233f
C616 B.n576 VSUBS 0.006233f
C617 B.n577 VSUBS 0.006233f
C618 B.n578 VSUBS 0.006233f
C619 B.n579 VSUBS 0.006233f
C620 B.n580 VSUBS 0.006233f
C621 B.n581 VSUBS 0.006233f
C622 B.n582 VSUBS 0.006233f
C623 B.n583 VSUBS 0.006233f
C624 B.n584 VSUBS 0.006233f
C625 B.n585 VSUBS 0.006233f
C626 B.n586 VSUBS 0.006233f
C627 B.n587 VSUBS 0.006233f
C628 B.n588 VSUBS 0.006233f
C629 B.n589 VSUBS 0.006233f
C630 B.n590 VSUBS 0.006233f
C631 B.n591 VSUBS 0.006233f
C632 B.n592 VSUBS 0.006233f
C633 B.n593 VSUBS 0.006233f
C634 B.n594 VSUBS 0.006233f
C635 B.n595 VSUBS 0.004308f
C636 B.n596 VSUBS 0.014442f
C637 B.n597 VSUBS 0.005042f
C638 B.n598 VSUBS 0.006233f
C639 B.n599 VSUBS 0.006233f
C640 B.n600 VSUBS 0.006233f
C641 B.n601 VSUBS 0.006233f
C642 B.n602 VSUBS 0.006233f
C643 B.n603 VSUBS 0.006233f
C644 B.n604 VSUBS 0.006233f
C645 B.n605 VSUBS 0.006233f
C646 B.n606 VSUBS 0.006233f
C647 B.n607 VSUBS 0.006233f
C648 B.n608 VSUBS 0.006233f
C649 B.n609 VSUBS 0.005042f
C650 B.n610 VSUBS 0.014442f
C651 B.n611 VSUBS 0.004308f
C652 B.n612 VSUBS 0.006233f
C653 B.n613 VSUBS 0.006233f
C654 B.n614 VSUBS 0.006233f
C655 B.n615 VSUBS 0.006233f
C656 B.n616 VSUBS 0.006233f
C657 B.n617 VSUBS 0.006233f
C658 B.n618 VSUBS 0.006233f
C659 B.n619 VSUBS 0.006233f
C660 B.n620 VSUBS 0.006233f
C661 B.n621 VSUBS 0.006233f
C662 B.n622 VSUBS 0.006233f
C663 B.n623 VSUBS 0.006233f
C664 B.n624 VSUBS 0.006233f
C665 B.n625 VSUBS 0.006233f
C666 B.n626 VSUBS 0.006233f
C667 B.n627 VSUBS 0.006233f
C668 B.n628 VSUBS 0.006233f
C669 B.n629 VSUBS 0.006233f
C670 B.n630 VSUBS 0.006233f
C671 B.n631 VSUBS 0.006233f
C672 B.n632 VSUBS 0.006233f
C673 B.n633 VSUBS 0.006233f
C674 B.n634 VSUBS 0.006233f
C675 B.n635 VSUBS 0.006233f
C676 B.n636 VSUBS 0.006233f
C677 B.n637 VSUBS 0.006233f
C678 B.n638 VSUBS 0.006233f
C679 B.n639 VSUBS 0.006233f
C680 B.n640 VSUBS 0.006233f
C681 B.n641 VSUBS 0.006233f
C682 B.n642 VSUBS 0.006233f
C683 B.n643 VSUBS 0.006233f
C684 B.n644 VSUBS 0.006233f
C685 B.n645 VSUBS 0.006233f
C686 B.n646 VSUBS 0.006233f
C687 B.n647 VSUBS 0.006233f
C688 B.n648 VSUBS 0.006233f
C689 B.n649 VSUBS 0.006233f
C690 B.n650 VSUBS 0.006233f
C691 B.n651 VSUBS 0.006233f
C692 B.n652 VSUBS 0.006233f
C693 B.n653 VSUBS 0.006233f
C694 B.n654 VSUBS 0.006233f
C695 B.n655 VSUBS 0.006233f
C696 B.n656 VSUBS 0.006233f
C697 B.n657 VSUBS 0.006233f
C698 B.n658 VSUBS 0.006233f
C699 B.n659 VSUBS 0.006233f
C700 B.n660 VSUBS 0.006233f
C701 B.n661 VSUBS 0.006233f
C702 B.n662 VSUBS 0.006233f
C703 B.n663 VSUBS 0.006233f
C704 B.n664 VSUBS 0.006233f
C705 B.n665 VSUBS 0.006233f
C706 B.n666 VSUBS 0.006233f
C707 B.n667 VSUBS 0.006233f
C708 B.n668 VSUBS 0.006233f
C709 B.n669 VSUBS 0.006233f
C710 B.n670 VSUBS 0.006233f
C711 B.n671 VSUBS 0.006233f
C712 B.n672 VSUBS 0.006233f
C713 B.n673 VSUBS 0.006233f
C714 B.n674 VSUBS 0.006233f
C715 B.n675 VSUBS 0.006233f
C716 B.n676 VSUBS 0.006233f
C717 B.n677 VSUBS 0.006233f
C718 B.n678 VSUBS 0.006233f
C719 B.n679 VSUBS 0.006233f
C720 B.n680 VSUBS 0.006233f
C721 B.n681 VSUBS 0.006233f
C722 B.n682 VSUBS 0.006233f
C723 B.n683 VSUBS 0.006233f
C724 B.n684 VSUBS 0.006233f
C725 B.n685 VSUBS 0.006233f
C726 B.n686 VSUBS 0.006233f
C727 B.n687 VSUBS 0.006233f
C728 B.n688 VSUBS 0.015265f
C729 B.n689 VSUBS 0.014802f
C730 B.n690 VSUBS 0.014802f
C731 B.n691 VSUBS 0.006233f
C732 B.n692 VSUBS 0.006233f
C733 B.n693 VSUBS 0.006233f
C734 B.n694 VSUBS 0.006233f
C735 B.n695 VSUBS 0.006233f
C736 B.n696 VSUBS 0.006233f
C737 B.n697 VSUBS 0.006233f
C738 B.n698 VSUBS 0.006233f
C739 B.n699 VSUBS 0.006233f
C740 B.n700 VSUBS 0.006233f
C741 B.n701 VSUBS 0.006233f
C742 B.n702 VSUBS 0.006233f
C743 B.n703 VSUBS 0.006233f
C744 B.n704 VSUBS 0.006233f
C745 B.n705 VSUBS 0.006233f
C746 B.n706 VSUBS 0.006233f
C747 B.n707 VSUBS 0.006233f
C748 B.n708 VSUBS 0.006233f
C749 B.n709 VSUBS 0.006233f
C750 B.n710 VSUBS 0.006233f
C751 B.n711 VSUBS 0.006233f
C752 B.n712 VSUBS 0.006233f
C753 B.n713 VSUBS 0.006233f
C754 B.n714 VSUBS 0.006233f
C755 B.n715 VSUBS 0.006233f
C756 B.n716 VSUBS 0.006233f
C757 B.n717 VSUBS 0.006233f
C758 B.n718 VSUBS 0.006233f
C759 B.n719 VSUBS 0.006233f
C760 B.n720 VSUBS 0.006233f
C761 B.n721 VSUBS 0.006233f
C762 B.n722 VSUBS 0.006233f
C763 B.n723 VSUBS 0.006233f
C764 B.n724 VSUBS 0.006233f
C765 B.n725 VSUBS 0.006233f
C766 B.n726 VSUBS 0.006233f
C767 B.n727 VSUBS 0.006233f
C768 B.n728 VSUBS 0.006233f
C769 B.n729 VSUBS 0.006233f
C770 B.n730 VSUBS 0.006233f
C771 B.n731 VSUBS 0.006233f
C772 B.n732 VSUBS 0.006233f
C773 B.n733 VSUBS 0.006233f
C774 B.n734 VSUBS 0.006233f
C775 B.n735 VSUBS 0.006233f
C776 B.n736 VSUBS 0.006233f
C777 B.n737 VSUBS 0.006233f
C778 B.n738 VSUBS 0.006233f
C779 B.n739 VSUBS 0.008134f
C780 B.n740 VSUBS 0.008665f
C781 B.n741 VSUBS 0.017231f
C782 VDD2.t2 VSUBS 0.326955f
C783 VDD2.t0 VSUBS 0.326955f
C784 VDD2.n0 VSUBS 3.50848f
C785 VDD2.t3 VSUBS 0.326955f
C786 VDD2.t1 VSUBS 0.326955f
C787 VDD2.n1 VSUBS 2.67467f
C788 VDD2.n2 VSUBS 4.68144f
C789 VN.t3 VSUBS 3.70977f
C790 VN.t1 VSUBS 3.71663f
C791 VN.n0 VSUBS 2.40531f
C792 VN.t0 VSUBS 3.70977f
C793 VN.t2 VSUBS 3.71663f
C794 VN.n1 VSUBS 4.22509f
C795 VDD1.t2 VSUBS 0.32699f
C796 VDD1.t3 VSUBS 0.32699f
C797 VDD1.n0 VSUBS 2.67555f
C798 VDD1.t0 VSUBS 0.32699f
C799 VDD1.t1 VSUBS 0.32699f
C800 VDD1.n1 VSUBS 3.53512f
C801 VTAIL.n0 VSUBS 0.02458f
C802 VTAIL.n1 VSUBS 0.02272f
C803 VTAIL.n2 VSUBS 0.012209f
C804 VTAIL.n3 VSUBS 0.028857f
C805 VTAIL.n4 VSUBS 0.012568f
C806 VTAIL.n5 VSUBS 0.02272f
C807 VTAIL.n6 VSUBS 0.012927f
C808 VTAIL.n7 VSUBS 0.028857f
C809 VTAIL.n8 VSUBS 0.012927f
C810 VTAIL.n9 VSUBS 0.02272f
C811 VTAIL.n10 VSUBS 0.012209f
C812 VTAIL.n11 VSUBS 0.028857f
C813 VTAIL.n12 VSUBS 0.012927f
C814 VTAIL.n13 VSUBS 0.02272f
C815 VTAIL.n14 VSUBS 0.012209f
C816 VTAIL.n15 VSUBS 0.028857f
C817 VTAIL.n16 VSUBS 0.012927f
C818 VTAIL.n17 VSUBS 0.02272f
C819 VTAIL.n18 VSUBS 0.012209f
C820 VTAIL.n19 VSUBS 0.028857f
C821 VTAIL.n20 VSUBS 0.012927f
C822 VTAIL.n21 VSUBS 0.02272f
C823 VTAIL.n22 VSUBS 0.012209f
C824 VTAIL.n23 VSUBS 0.028857f
C825 VTAIL.n24 VSUBS 0.012927f
C826 VTAIL.n25 VSUBS 1.50126f
C827 VTAIL.n26 VSUBS 0.012209f
C828 VTAIL.t5 VSUBS 0.061805f
C829 VTAIL.n27 VSUBS 0.16344f
C830 VTAIL.n28 VSUBS 0.018358f
C831 VTAIL.n29 VSUBS 0.021643f
C832 VTAIL.n30 VSUBS 0.028857f
C833 VTAIL.n31 VSUBS 0.012927f
C834 VTAIL.n32 VSUBS 0.012209f
C835 VTAIL.n33 VSUBS 0.02272f
C836 VTAIL.n34 VSUBS 0.02272f
C837 VTAIL.n35 VSUBS 0.012209f
C838 VTAIL.n36 VSUBS 0.012927f
C839 VTAIL.n37 VSUBS 0.028857f
C840 VTAIL.n38 VSUBS 0.028857f
C841 VTAIL.n39 VSUBS 0.012927f
C842 VTAIL.n40 VSUBS 0.012209f
C843 VTAIL.n41 VSUBS 0.02272f
C844 VTAIL.n42 VSUBS 0.02272f
C845 VTAIL.n43 VSUBS 0.012209f
C846 VTAIL.n44 VSUBS 0.012927f
C847 VTAIL.n45 VSUBS 0.028857f
C848 VTAIL.n46 VSUBS 0.028857f
C849 VTAIL.n47 VSUBS 0.012927f
C850 VTAIL.n48 VSUBS 0.012209f
C851 VTAIL.n49 VSUBS 0.02272f
C852 VTAIL.n50 VSUBS 0.02272f
C853 VTAIL.n51 VSUBS 0.012209f
C854 VTAIL.n52 VSUBS 0.012927f
C855 VTAIL.n53 VSUBS 0.028857f
C856 VTAIL.n54 VSUBS 0.028857f
C857 VTAIL.n55 VSUBS 0.012927f
C858 VTAIL.n56 VSUBS 0.012209f
C859 VTAIL.n57 VSUBS 0.02272f
C860 VTAIL.n58 VSUBS 0.02272f
C861 VTAIL.n59 VSUBS 0.012209f
C862 VTAIL.n60 VSUBS 0.012927f
C863 VTAIL.n61 VSUBS 0.028857f
C864 VTAIL.n62 VSUBS 0.028857f
C865 VTAIL.n63 VSUBS 0.012927f
C866 VTAIL.n64 VSUBS 0.012209f
C867 VTAIL.n65 VSUBS 0.02272f
C868 VTAIL.n66 VSUBS 0.02272f
C869 VTAIL.n67 VSUBS 0.012209f
C870 VTAIL.n68 VSUBS 0.012209f
C871 VTAIL.n69 VSUBS 0.012927f
C872 VTAIL.n70 VSUBS 0.028857f
C873 VTAIL.n71 VSUBS 0.028857f
C874 VTAIL.n72 VSUBS 0.028857f
C875 VTAIL.n73 VSUBS 0.012568f
C876 VTAIL.n74 VSUBS 0.012209f
C877 VTAIL.n75 VSUBS 0.02272f
C878 VTAIL.n76 VSUBS 0.02272f
C879 VTAIL.n77 VSUBS 0.012209f
C880 VTAIL.n78 VSUBS 0.012927f
C881 VTAIL.n79 VSUBS 0.028857f
C882 VTAIL.n80 VSUBS 0.068552f
C883 VTAIL.n81 VSUBS 0.012927f
C884 VTAIL.n82 VSUBS 0.012209f
C885 VTAIL.n83 VSUBS 0.056551f
C886 VTAIL.n84 VSUBS 0.034536f
C887 VTAIL.n85 VSUBS 0.154692f
C888 VTAIL.n86 VSUBS 0.02458f
C889 VTAIL.n87 VSUBS 0.02272f
C890 VTAIL.n88 VSUBS 0.012209f
C891 VTAIL.n89 VSUBS 0.028857f
C892 VTAIL.n90 VSUBS 0.012568f
C893 VTAIL.n91 VSUBS 0.02272f
C894 VTAIL.n92 VSUBS 0.012927f
C895 VTAIL.n93 VSUBS 0.028857f
C896 VTAIL.n94 VSUBS 0.012927f
C897 VTAIL.n95 VSUBS 0.02272f
C898 VTAIL.n96 VSUBS 0.012209f
C899 VTAIL.n97 VSUBS 0.028857f
C900 VTAIL.n98 VSUBS 0.012927f
C901 VTAIL.n99 VSUBS 0.02272f
C902 VTAIL.n100 VSUBS 0.012209f
C903 VTAIL.n101 VSUBS 0.028857f
C904 VTAIL.n102 VSUBS 0.012927f
C905 VTAIL.n103 VSUBS 0.02272f
C906 VTAIL.n104 VSUBS 0.012209f
C907 VTAIL.n105 VSUBS 0.028857f
C908 VTAIL.n106 VSUBS 0.012927f
C909 VTAIL.n107 VSUBS 0.02272f
C910 VTAIL.n108 VSUBS 0.012209f
C911 VTAIL.n109 VSUBS 0.028857f
C912 VTAIL.n110 VSUBS 0.012927f
C913 VTAIL.n111 VSUBS 1.50126f
C914 VTAIL.n112 VSUBS 0.012209f
C915 VTAIL.t2 VSUBS 0.061805f
C916 VTAIL.n113 VSUBS 0.16344f
C917 VTAIL.n114 VSUBS 0.018358f
C918 VTAIL.n115 VSUBS 0.021643f
C919 VTAIL.n116 VSUBS 0.028857f
C920 VTAIL.n117 VSUBS 0.012927f
C921 VTAIL.n118 VSUBS 0.012209f
C922 VTAIL.n119 VSUBS 0.02272f
C923 VTAIL.n120 VSUBS 0.02272f
C924 VTAIL.n121 VSUBS 0.012209f
C925 VTAIL.n122 VSUBS 0.012927f
C926 VTAIL.n123 VSUBS 0.028857f
C927 VTAIL.n124 VSUBS 0.028857f
C928 VTAIL.n125 VSUBS 0.012927f
C929 VTAIL.n126 VSUBS 0.012209f
C930 VTAIL.n127 VSUBS 0.02272f
C931 VTAIL.n128 VSUBS 0.02272f
C932 VTAIL.n129 VSUBS 0.012209f
C933 VTAIL.n130 VSUBS 0.012927f
C934 VTAIL.n131 VSUBS 0.028857f
C935 VTAIL.n132 VSUBS 0.028857f
C936 VTAIL.n133 VSUBS 0.012927f
C937 VTAIL.n134 VSUBS 0.012209f
C938 VTAIL.n135 VSUBS 0.02272f
C939 VTAIL.n136 VSUBS 0.02272f
C940 VTAIL.n137 VSUBS 0.012209f
C941 VTAIL.n138 VSUBS 0.012927f
C942 VTAIL.n139 VSUBS 0.028857f
C943 VTAIL.n140 VSUBS 0.028857f
C944 VTAIL.n141 VSUBS 0.012927f
C945 VTAIL.n142 VSUBS 0.012209f
C946 VTAIL.n143 VSUBS 0.02272f
C947 VTAIL.n144 VSUBS 0.02272f
C948 VTAIL.n145 VSUBS 0.012209f
C949 VTAIL.n146 VSUBS 0.012927f
C950 VTAIL.n147 VSUBS 0.028857f
C951 VTAIL.n148 VSUBS 0.028857f
C952 VTAIL.n149 VSUBS 0.012927f
C953 VTAIL.n150 VSUBS 0.012209f
C954 VTAIL.n151 VSUBS 0.02272f
C955 VTAIL.n152 VSUBS 0.02272f
C956 VTAIL.n153 VSUBS 0.012209f
C957 VTAIL.n154 VSUBS 0.012209f
C958 VTAIL.n155 VSUBS 0.012927f
C959 VTAIL.n156 VSUBS 0.028857f
C960 VTAIL.n157 VSUBS 0.028857f
C961 VTAIL.n158 VSUBS 0.028857f
C962 VTAIL.n159 VSUBS 0.012568f
C963 VTAIL.n160 VSUBS 0.012209f
C964 VTAIL.n161 VSUBS 0.02272f
C965 VTAIL.n162 VSUBS 0.02272f
C966 VTAIL.n163 VSUBS 0.012209f
C967 VTAIL.n164 VSUBS 0.012927f
C968 VTAIL.n165 VSUBS 0.028857f
C969 VTAIL.n166 VSUBS 0.068552f
C970 VTAIL.n167 VSUBS 0.012927f
C971 VTAIL.n168 VSUBS 0.012209f
C972 VTAIL.n169 VSUBS 0.056551f
C973 VTAIL.n170 VSUBS 0.034536f
C974 VTAIL.n171 VSUBS 0.244783f
C975 VTAIL.n172 VSUBS 0.02458f
C976 VTAIL.n173 VSUBS 0.02272f
C977 VTAIL.n174 VSUBS 0.012209f
C978 VTAIL.n175 VSUBS 0.028857f
C979 VTAIL.n176 VSUBS 0.012568f
C980 VTAIL.n177 VSUBS 0.02272f
C981 VTAIL.n178 VSUBS 0.012927f
C982 VTAIL.n179 VSUBS 0.028857f
C983 VTAIL.n180 VSUBS 0.012927f
C984 VTAIL.n181 VSUBS 0.02272f
C985 VTAIL.n182 VSUBS 0.012209f
C986 VTAIL.n183 VSUBS 0.028857f
C987 VTAIL.n184 VSUBS 0.012927f
C988 VTAIL.n185 VSUBS 0.02272f
C989 VTAIL.n186 VSUBS 0.012209f
C990 VTAIL.n187 VSUBS 0.028857f
C991 VTAIL.n188 VSUBS 0.012927f
C992 VTAIL.n189 VSUBS 0.02272f
C993 VTAIL.n190 VSUBS 0.012209f
C994 VTAIL.n191 VSUBS 0.028857f
C995 VTAIL.n192 VSUBS 0.012927f
C996 VTAIL.n193 VSUBS 0.02272f
C997 VTAIL.n194 VSUBS 0.012209f
C998 VTAIL.n195 VSUBS 0.028857f
C999 VTAIL.n196 VSUBS 0.012927f
C1000 VTAIL.n197 VSUBS 1.50126f
C1001 VTAIL.n198 VSUBS 0.012209f
C1002 VTAIL.t4 VSUBS 0.061805f
C1003 VTAIL.n199 VSUBS 0.16344f
C1004 VTAIL.n200 VSUBS 0.018358f
C1005 VTAIL.n201 VSUBS 0.021643f
C1006 VTAIL.n202 VSUBS 0.028857f
C1007 VTAIL.n203 VSUBS 0.012927f
C1008 VTAIL.n204 VSUBS 0.012209f
C1009 VTAIL.n205 VSUBS 0.02272f
C1010 VTAIL.n206 VSUBS 0.02272f
C1011 VTAIL.n207 VSUBS 0.012209f
C1012 VTAIL.n208 VSUBS 0.012927f
C1013 VTAIL.n209 VSUBS 0.028857f
C1014 VTAIL.n210 VSUBS 0.028857f
C1015 VTAIL.n211 VSUBS 0.012927f
C1016 VTAIL.n212 VSUBS 0.012209f
C1017 VTAIL.n213 VSUBS 0.02272f
C1018 VTAIL.n214 VSUBS 0.02272f
C1019 VTAIL.n215 VSUBS 0.012209f
C1020 VTAIL.n216 VSUBS 0.012927f
C1021 VTAIL.n217 VSUBS 0.028857f
C1022 VTAIL.n218 VSUBS 0.028857f
C1023 VTAIL.n219 VSUBS 0.012927f
C1024 VTAIL.n220 VSUBS 0.012209f
C1025 VTAIL.n221 VSUBS 0.02272f
C1026 VTAIL.n222 VSUBS 0.02272f
C1027 VTAIL.n223 VSUBS 0.012209f
C1028 VTAIL.n224 VSUBS 0.012927f
C1029 VTAIL.n225 VSUBS 0.028857f
C1030 VTAIL.n226 VSUBS 0.028857f
C1031 VTAIL.n227 VSUBS 0.012927f
C1032 VTAIL.n228 VSUBS 0.012209f
C1033 VTAIL.n229 VSUBS 0.02272f
C1034 VTAIL.n230 VSUBS 0.02272f
C1035 VTAIL.n231 VSUBS 0.012209f
C1036 VTAIL.n232 VSUBS 0.012927f
C1037 VTAIL.n233 VSUBS 0.028857f
C1038 VTAIL.n234 VSUBS 0.028857f
C1039 VTAIL.n235 VSUBS 0.012927f
C1040 VTAIL.n236 VSUBS 0.012209f
C1041 VTAIL.n237 VSUBS 0.02272f
C1042 VTAIL.n238 VSUBS 0.02272f
C1043 VTAIL.n239 VSUBS 0.012209f
C1044 VTAIL.n240 VSUBS 0.012209f
C1045 VTAIL.n241 VSUBS 0.012927f
C1046 VTAIL.n242 VSUBS 0.028857f
C1047 VTAIL.n243 VSUBS 0.028857f
C1048 VTAIL.n244 VSUBS 0.028857f
C1049 VTAIL.n245 VSUBS 0.012568f
C1050 VTAIL.n246 VSUBS 0.012209f
C1051 VTAIL.n247 VSUBS 0.02272f
C1052 VTAIL.n248 VSUBS 0.02272f
C1053 VTAIL.n249 VSUBS 0.012209f
C1054 VTAIL.n250 VSUBS 0.012927f
C1055 VTAIL.n251 VSUBS 0.028857f
C1056 VTAIL.n252 VSUBS 0.068552f
C1057 VTAIL.n253 VSUBS 0.012927f
C1058 VTAIL.n254 VSUBS 0.012209f
C1059 VTAIL.n255 VSUBS 0.056551f
C1060 VTAIL.n256 VSUBS 0.034536f
C1061 VTAIL.n257 VSUBS 1.6853f
C1062 VTAIL.n258 VSUBS 0.02458f
C1063 VTAIL.n259 VSUBS 0.02272f
C1064 VTAIL.n260 VSUBS 0.012209f
C1065 VTAIL.n261 VSUBS 0.028857f
C1066 VTAIL.n262 VSUBS 0.012568f
C1067 VTAIL.n263 VSUBS 0.02272f
C1068 VTAIL.n264 VSUBS 0.012568f
C1069 VTAIL.n265 VSUBS 0.012209f
C1070 VTAIL.n266 VSUBS 0.028857f
C1071 VTAIL.n267 VSUBS 0.028857f
C1072 VTAIL.n268 VSUBS 0.012927f
C1073 VTAIL.n269 VSUBS 0.02272f
C1074 VTAIL.n270 VSUBS 0.012209f
C1075 VTAIL.n271 VSUBS 0.028857f
C1076 VTAIL.n272 VSUBS 0.012927f
C1077 VTAIL.n273 VSUBS 0.02272f
C1078 VTAIL.n274 VSUBS 0.012209f
C1079 VTAIL.n275 VSUBS 0.028857f
C1080 VTAIL.n276 VSUBS 0.012927f
C1081 VTAIL.n277 VSUBS 0.02272f
C1082 VTAIL.n278 VSUBS 0.012209f
C1083 VTAIL.n279 VSUBS 0.028857f
C1084 VTAIL.n280 VSUBS 0.012927f
C1085 VTAIL.n281 VSUBS 0.02272f
C1086 VTAIL.n282 VSUBS 0.012209f
C1087 VTAIL.n283 VSUBS 0.028857f
C1088 VTAIL.n284 VSUBS 0.012927f
C1089 VTAIL.n285 VSUBS 1.50126f
C1090 VTAIL.n286 VSUBS 0.012209f
C1091 VTAIL.t0 VSUBS 0.061805f
C1092 VTAIL.n287 VSUBS 0.16344f
C1093 VTAIL.n288 VSUBS 0.018358f
C1094 VTAIL.n289 VSUBS 0.021643f
C1095 VTAIL.n290 VSUBS 0.028857f
C1096 VTAIL.n291 VSUBS 0.012927f
C1097 VTAIL.n292 VSUBS 0.012209f
C1098 VTAIL.n293 VSUBS 0.02272f
C1099 VTAIL.n294 VSUBS 0.02272f
C1100 VTAIL.n295 VSUBS 0.012209f
C1101 VTAIL.n296 VSUBS 0.012927f
C1102 VTAIL.n297 VSUBS 0.028857f
C1103 VTAIL.n298 VSUBS 0.028857f
C1104 VTAIL.n299 VSUBS 0.012927f
C1105 VTAIL.n300 VSUBS 0.012209f
C1106 VTAIL.n301 VSUBS 0.02272f
C1107 VTAIL.n302 VSUBS 0.02272f
C1108 VTAIL.n303 VSUBS 0.012209f
C1109 VTAIL.n304 VSUBS 0.012927f
C1110 VTAIL.n305 VSUBS 0.028857f
C1111 VTAIL.n306 VSUBS 0.028857f
C1112 VTAIL.n307 VSUBS 0.012927f
C1113 VTAIL.n308 VSUBS 0.012209f
C1114 VTAIL.n309 VSUBS 0.02272f
C1115 VTAIL.n310 VSUBS 0.02272f
C1116 VTAIL.n311 VSUBS 0.012209f
C1117 VTAIL.n312 VSUBS 0.012927f
C1118 VTAIL.n313 VSUBS 0.028857f
C1119 VTAIL.n314 VSUBS 0.028857f
C1120 VTAIL.n315 VSUBS 0.012927f
C1121 VTAIL.n316 VSUBS 0.012209f
C1122 VTAIL.n317 VSUBS 0.02272f
C1123 VTAIL.n318 VSUBS 0.02272f
C1124 VTAIL.n319 VSUBS 0.012209f
C1125 VTAIL.n320 VSUBS 0.012927f
C1126 VTAIL.n321 VSUBS 0.028857f
C1127 VTAIL.n322 VSUBS 0.028857f
C1128 VTAIL.n323 VSUBS 0.012927f
C1129 VTAIL.n324 VSUBS 0.012209f
C1130 VTAIL.n325 VSUBS 0.02272f
C1131 VTAIL.n326 VSUBS 0.02272f
C1132 VTAIL.n327 VSUBS 0.012209f
C1133 VTAIL.n328 VSUBS 0.012927f
C1134 VTAIL.n329 VSUBS 0.028857f
C1135 VTAIL.n330 VSUBS 0.028857f
C1136 VTAIL.n331 VSUBS 0.012927f
C1137 VTAIL.n332 VSUBS 0.012209f
C1138 VTAIL.n333 VSUBS 0.02272f
C1139 VTAIL.n334 VSUBS 0.02272f
C1140 VTAIL.n335 VSUBS 0.012209f
C1141 VTAIL.n336 VSUBS 0.012927f
C1142 VTAIL.n337 VSUBS 0.028857f
C1143 VTAIL.n338 VSUBS 0.068552f
C1144 VTAIL.n339 VSUBS 0.012927f
C1145 VTAIL.n340 VSUBS 0.012209f
C1146 VTAIL.n341 VSUBS 0.056551f
C1147 VTAIL.n342 VSUBS 0.034536f
C1148 VTAIL.n343 VSUBS 1.6853f
C1149 VTAIL.n344 VSUBS 0.02458f
C1150 VTAIL.n345 VSUBS 0.02272f
C1151 VTAIL.n346 VSUBS 0.012209f
C1152 VTAIL.n347 VSUBS 0.028857f
C1153 VTAIL.n348 VSUBS 0.012568f
C1154 VTAIL.n349 VSUBS 0.02272f
C1155 VTAIL.n350 VSUBS 0.012568f
C1156 VTAIL.n351 VSUBS 0.012209f
C1157 VTAIL.n352 VSUBS 0.028857f
C1158 VTAIL.n353 VSUBS 0.028857f
C1159 VTAIL.n354 VSUBS 0.012927f
C1160 VTAIL.n355 VSUBS 0.02272f
C1161 VTAIL.n356 VSUBS 0.012209f
C1162 VTAIL.n357 VSUBS 0.028857f
C1163 VTAIL.n358 VSUBS 0.012927f
C1164 VTAIL.n359 VSUBS 0.02272f
C1165 VTAIL.n360 VSUBS 0.012209f
C1166 VTAIL.n361 VSUBS 0.028857f
C1167 VTAIL.n362 VSUBS 0.012927f
C1168 VTAIL.n363 VSUBS 0.02272f
C1169 VTAIL.n364 VSUBS 0.012209f
C1170 VTAIL.n365 VSUBS 0.028857f
C1171 VTAIL.n366 VSUBS 0.012927f
C1172 VTAIL.n367 VSUBS 0.02272f
C1173 VTAIL.n368 VSUBS 0.012209f
C1174 VTAIL.n369 VSUBS 0.028857f
C1175 VTAIL.n370 VSUBS 0.012927f
C1176 VTAIL.n371 VSUBS 1.50126f
C1177 VTAIL.n372 VSUBS 0.012209f
C1178 VTAIL.t7 VSUBS 0.061805f
C1179 VTAIL.n373 VSUBS 0.16344f
C1180 VTAIL.n374 VSUBS 0.018358f
C1181 VTAIL.n375 VSUBS 0.021643f
C1182 VTAIL.n376 VSUBS 0.028857f
C1183 VTAIL.n377 VSUBS 0.012927f
C1184 VTAIL.n378 VSUBS 0.012209f
C1185 VTAIL.n379 VSUBS 0.02272f
C1186 VTAIL.n380 VSUBS 0.02272f
C1187 VTAIL.n381 VSUBS 0.012209f
C1188 VTAIL.n382 VSUBS 0.012927f
C1189 VTAIL.n383 VSUBS 0.028857f
C1190 VTAIL.n384 VSUBS 0.028857f
C1191 VTAIL.n385 VSUBS 0.012927f
C1192 VTAIL.n386 VSUBS 0.012209f
C1193 VTAIL.n387 VSUBS 0.02272f
C1194 VTAIL.n388 VSUBS 0.02272f
C1195 VTAIL.n389 VSUBS 0.012209f
C1196 VTAIL.n390 VSUBS 0.012927f
C1197 VTAIL.n391 VSUBS 0.028857f
C1198 VTAIL.n392 VSUBS 0.028857f
C1199 VTAIL.n393 VSUBS 0.012927f
C1200 VTAIL.n394 VSUBS 0.012209f
C1201 VTAIL.n395 VSUBS 0.02272f
C1202 VTAIL.n396 VSUBS 0.02272f
C1203 VTAIL.n397 VSUBS 0.012209f
C1204 VTAIL.n398 VSUBS 0.012927f
C1205 VTAIL.n399 VSUBS 0.028857f
C1206 VTAIL.n400 VSUBS 0.028857f
C1207 VTAIL.n401 VSUBS 0.012927f
C1208 VTAIL.n402 VSUBS 0.012209f
C1209 VTAIL.n403 VSUBS 0.02272f
C1210 VTAIL.n404 VSUBS 0.02272f
C1211 VTAIL.n405 VSUBS 0.012209f
C1212 VTAIL.n406 VSUBS 0.012927f
C1213 VTAIL.n407 VSUBS 0.028857f
C1214 VTAIL.n408 VSUBS 0.028857f
C1215 VTAIL.n409 VSUBS 0.012927f
C1216 VTAIL.n410 VSUBS 0.012209f
C1217 VTAIL.n411 VSUBS 0.02272f
C1218 VTAIL.n412 VSUBS 0.02272f
C1219 VTAIL.n413 VSUBS 0.012209f
C1220 VTAIL.n414 VSUBS 0.012927f
C1221 VTAIL.n415 VSUBS 0.028857f
C1222 VTAIL.n416 VSUBS 0.028857f
C1223 VTAIL.n417 VSUBS 0.012927f
C1224 VTAIL.n418 VSUBS 0.012209f
C1225 VTAIL.n419 VSUBS 0.02272f
C1226 VTAIL.n420 VSUBS 0.02272f
C1227 VTAIL.n421 VSUBS 0.012209f
C1228 VTAIL.n422 VSUBS 0.012927f
C1229 VTAIL.n423 VSUBS 0.028857f
C1230 VTAIL.n424 VSUBS 0.068552f
C1231 VTAIL.n425 VSUBS 0.012927f
C1232 VTAIL.n426 VSUBS 0.012209f
C1233 VTAIL.n427 VSUBS 0.056551f
C1234 VTAIL.n428 VSUBS 0.034536f
C1235 VTAIL.n429 VSUBS 0.244783f
C1236 VTAIL.n430 VSUBS 0.02458f
C1237 VTAIL.n431 VSUBS 0.02272f
C1238 VTAIL.n432 VSUBS 0.012209f
C1239 VTAIL.n433 VSUBS 0.028857f
C1240 VTAIL.n434 VSUBS 0.012568f
C1241 VTAIL.n435 VSUBS 0.02272f
C1242 VTAIL.n436 VSUBS 0.012568f
C1243 VTAIL.n437 VSUBS 0.012209f
C1244 VTAIL.n438 VSUBS 0.028857f
C1245 VTAIL.n439 VSUBS 0.028857f
C1246 VTAIL.n440 VSUBS 0.012927f
C1247 VTAIL.n441 VSUBS 0.02272f
C1248 VTAIL.n442 VSUBS 0.012209f
C1249 VTAIL.n443 VSUBS 0.028857f
C1250 VTAIL.n444 VSUBS 0.012927f
C1251 VTAIL.n445 VSUBS 0.02272f
C1252 VTAIL.n446 VSUBS 0.012209f
C1253 VTAIL.n447 VSUBS 0.028857f
C1254 VTAIL.n448 VSUBS 0.012927f
C1255 VTAIL.n449 VSUBS 0.02272f
C1256 VTAIL.n450 VSUBS 0.012209f
C1257 VTAIL.n451 VSUBS 0.028857f
C1258 VTAIL.n452 VSUBS 0.012927f
C1259 VTAIL.n453 VSUBS 0.02272f
C1260 VTAIL.n454 VSUBS 0.012209f
C1261 VTAIL.n455 VSUBS 0.028857f
C1262 VTAIL.n456 VSUBS 0.012927f
C1263 VTAIL.n457 VSUBS 1.50126f
C1264 VTAIL.n458 VSUBS 0.012209f
C1265 VTAIL.t3 VSUBS 0.061805f
C1266 VTAIL.n459 VSUBS 0.16344f
C1267 VTAIL.n460 VSUBS 0.018358f
C1268 VTAIL.n461 VSUBS 0.021643f
C1269 VTAIL.n462 VSUBS 0.028857f
C1270 VTAIL.n463 VSUBS 0.012927f
C1271 VTAIL.n464 VSUBS 0.012209f
C1272 VTAIL.n465 VSUBS 0.02272f
C1273 VTAIL.n466 VSUBS 0.02272f
C1274 VTAIL.n467 VSUBS 0.012209f
C1275 VTAIL.n468 VSUBS 0.012927f
C1276 VTAIL.n469 VSUBS 0.028857f
C1277 VTAIL.n470 VSUBS 0.028857f
C1278 VTAIL.n471 VSUBS 0.012927f
C1279 VTAIL.n472 VSUBS 0.012209f
C1280 VTAIL.n473 VSUBS 0.02272f
C1281 VTAIL.n474 VSUBS 0.02272f
C1282 VTAIL.n475 VSUBS 0.012209f
C1283 VTAIL.n476 VSUBS 0.012927f
C1284 VTAIL.n477 VSUBS 0.028857f
C1285 VTAIL.n478 VSUBS 0.028857f
C1286 VTAIL.n479 VSUBS 0.012927f
C1287 VTAIL.n480 VSUBS 0.012209f
C1288 VTAIL.n481 VSUBS 0.02272f
C1289 VTAIL.n482 VSUBS 0.02272f
C1290 VTAIL.n483 VSUBS 0.012209f
C1291 VTAIL.n484 VSUBS 0.012927f
C1292 VTAIL.n485 VSUBS 0.028857f
C1293 VTAIL.n486 VSUBS 0.028857f
C1294 VTAIL.n487 VSUBS 0.012927f
C1295 VTAIL.n488 VSUBS 0.012209f
C1296 VTAIL.n489 VSUBS 0.02272f
C1297 VTAIL.n490 VSUBS 0.02272f
C1298 VTAIL.n491 VSUBS 0.012209f
C1299 VTAIL.n492 VSUBS 0.012927f
C1300 VTAIL.n493 VSUBS 0.028857f
C1301 VTAIL.n494 VSUBS 0.028857f
C1302 VTAIL.n495 VSUBS 0.012927f
C1303 VTAIL.n496 VSUBS 0.012209f
C1304 VTAIL.n497 VSUBS 0.02272f
C1305 VTAIL.n498 VSUBS 0.02272f
C1306 VTAIL.n499 VSUBS 0.012209f
C1307 VTAIL.n500 VSUBS 0.012927f
C1308 VTAIL.n501 VSUBS 0.028857f
C1309 VTAIL.n502 VSUBS 0.028857f
C1310 VTAIL.n503 VSUBS 0.012927f
C1311 VTAIL.n504 VSUBS 0.012209f
C1312 VTAIL.n505 VSUBS 0.02272f
C1313 VTAIL.n506 VSUBS 0.02272f
C1314 VTAIL.n507 VSUBS 0.012209f
C1315 VTAIL.n508 VSUBS 0.012927f
C1316 VTAIL.n509 VSUBS 0.028857f
C1317 VTAIL.n510 VSUBS 0.068552f
C1318 VTAIL.n511 VSUBS 0.012927f
C1319 VTAIL.n512 VSUBS 0.012209f
C1320 VTAIL.n513 VSUBS 0.056551f
C1321 VTAIL.n514 VSUBS 0.034536f
C1322 VTAIL.n515 VSUBS 0.244783f
C1323 VTAIL.n516 VSUBS 0.02458f
C1324 VTAIL.n517 VSUBS 0.02272f
C1325 VTAIL.n518 VSUBS 0.012209f
C1326 VTAIL.n519 VSUBS 0.028857f
C1327 VTAIL.n520 VSUBS 0.012568f
C1328 VTAIL.n521 VSUBS 0.02272f
C1329 VTAIL.n522 VSUBS 0.012568f
C1330 VTAIL.n523 VSUBS 0.012209f
C1331 VTAIL.n524 VSUBS 0.028857f
C1332 VTAIL.n525 VSUBS 0.028857f
C1333 VTAIL.n526 VSUBS 0.012927f
C1334 VTAIL.n527 VSUBS 0.02272f
C1335 VTAIL.n528 VSUBS 0.012209f
C1336 VTAIL.n529 VSUBS 0.028857f
C1337 VTAIL.n530 VSUBS 0.012927f
C1338 VTAIL.n531 VSUBS 0.02272f
C1339 VTAIL.n532 VSUBS 0.012209f
C1340 VTAIL.n533 VSUBS 0.028857f
C1341 VTAIL.n534 VSUBS 0.012927f
C1342 VTAIL.n535 VSUBS 0.02272f
C1343 VTAIL.n536 VSUBS 0.012209f
C1344 VTAIL.n537 VSUBS 0.028857f
C1345 VTAIL.n538 VSUBS 0.012927f
C1346 VTAIL.n539 VSUBS 0.02272f
C1347 VTAIL.n540 VSUBS 0.012209f
C1348 VTAIL.n541 VSUBS 0.028857f
C1349 VTAIL.n542 VSUBS 0.012927f
C1350 VTAIL.n543 VSUBS 1.50126f
C1351 VTAIL.n544 VSUBS 0.012209f
C1352 VTAIL.t1 VSUBS 0.061805f
C1353 VTAIL.n545 VSUBS 0.16344f
C1354 VTAIL.n546 VSUBS 0.018358f
C1355 VTAIL.n547 VSUBS 0.021643f
C1356 VTAIL.n548 VSUBS 0.028857f
C1357 VTAIL.n549 VSUBS 0.012927f
C1358 VTAIL.n550 VSUBS 0.012209f
C1359 VTAIL.n551 VSUBS 0.02272f
C1360 VTAIL.n552 VSUBS 0.02272f
C1361 VTAIL.n553 VSUBS 0.012209f
C1362 VTAIL.n554 VSUBS 0.012927f
C1363 VTAIL.n555 VSUBS 0.028857f
C1364 VTAIL.n556 VSUBS 0.028857f
C1365 VTAIL.n557 VSUBS 0.012927f
C1366 VTAIL.n558 VSUBS 0.012209f
C1367 VTAIL.n559 VSUBS 0.02272f
C1368 VTAIL.n560 VSUBS 0.02272f
C1369 VTAIL.n561 VSUBS 0.012209f
C1370 VTAIL.n562 VSUBS 0.012927f
C1371 VTAIL.n563 VSUBS 0.028857f
C1372 VTAIL.n564 VSUBS 0.028857f
C1373 VTAIL.n565 VSUBS 0.012927f
C1374 VTAIL.n566 VSUBS 0.012209f
C1375 VTAIL.n567 VSUBS 0.02272f
C1376 VTAIL.n568 VSUBS 0.02272f
C1377 VTAIL.n569 VSUBS 0.012209f
C1378 VTAIL.n570 VSUBS 0.012927f
C1379 VTAIL.n571 VSUBS 0.028857f
C1380 VTAIL.n572 VSUBS 0.028857f
C1381 VTAIL.n573 VSUBS 0.012927f
C1382 VTAIL.n574 VSUBS 0.012209f
C1383 VTAIL.n575 VSUBS 0.02272f
C1384 VTAIL.n576 VSUBS 0.02272f
C1385 VTAIL.n577 VSUBS 0.012209f
C1386 VTAIL.n578 VSUBS 0.012927f
C1387 VTAIL.n579 VSUBS 0.028857f
C1388 VTAIL.n580 VSUBS 0.028857f
C1389 VTAIL.n581 VSUBS 0.012927f
C1390 VTAIL.n582 VSUBS 0.012209f
C1391 VTAIL.n583 VSUBS 0.02272f
C1392 VTAIL.n584 VSUBS 0.02272f
C1393 VTAIL.n585 VSUBS 0.012209f
C1394 VTAIL.n586 VSUBS 0.012927f
C1395 VTAIL.n587 VSUBS 0.028857f
C1396 VTAIL.n588 VSUBS 0.028857f
C1397 VTAIL.n589 VSUBS 0.012927f
C1398 VTAIL.n590 VSUBS 0.012209f
C1399 VTAIL.n591 VSUBS 0.02272f
C1400 VTAIL.n592 VSUBS 0.02272f
C1401 VTAIL.n593 VSUBS 0.012209f
C1402 VTAIL.n594 VSUBS 0.012927f
C1403 VTAIL.n595 VSUBS 0.028857f
C1404 VTAIL.n596 VSUBS 0.068552f
C1405 VTAIL.n597 VSUBS 0.012927f
C1406 VTAIL.n598 VSUBS 0.012209f
C1407 VTAIL.n599 VSUBS 0.056551f
C1408 VTAIL.n600 VSUBS 0.034536f
C1409 VTAIL.n601 VSUBS 1.6853f
C1410 VTAIL.n602 VSUBS 0.02458f
C1411 VTAIL.n603 VSUBS 0.02272f
C1412 VTAIL.n604 VSUBS 0.012209f
C1413 VTAIL.n605 VSUBS 0.028857f
C1414 VTAIL.n606 VSUBS 0.012568f
C1415 VTAIL.n607 VSUBS 0.02272f
C1416 VTAIL.n608 VSUBS 0.012927f
C1417 VTAIL.n609 VSUBS 0.028857f
C1418 VTAIL.n610 VSUBS 0.012927f
C1419 VTAIL.n611 VSUBS 0.02272f
C1420 VTAIL.n612 VSUBS 0.012209f
C1421 VTAIL.n613 VSUBS 0.028857f
C1422 VTAIL.n614 VSUBS 0.012927f
C1423 VTAIL.n615 VSUBS 0.02272f
C1424 VTAIL.n616 VSUBS 0.012209f
C1425 VTAIL.n617 VSUBS 0.028857f
C1426 VTAIL.n618 VSUBS 0.012927f
C1427 VTAIL.n619 VSUBS 0.02272f
C1428 VTAIL.n620 VSUBS 0.012209f
C1429 VTAIL.n621 VSUBS 0.028857f
C1430 VTAIL.n622 VSUBS 0.012927f
C1431 VTAIL.n623 VSUBS 0.02272f
C1432 VTAIL.n624 VSUBS 0.012209f
C1433 VTAIL.n625 VSUBS 0.028857f
C1434 VTAIL.n626 VSUBS 0.012927f
C1435 VTAIL.n627 VSUBS 1.50126f
C1436 VTAIL.n628 VSUBS 0.012209f
C1437 VTAIL.t6 VSUBS 0.061805f
C1438 VTAIL.n629 VSUBS 0.16344f
C1439 VTAIL.n630 VSUBS 0.018358f
C1440 VTAIL.n631 VSUBS 0.021643f
C1441 VTAIL.n632 VSUBS 0.028857f
C1442 VTAIL.n633 VSUBS 0.012927f
C1443 VTAIL.n634 VSUBS 0.012209f
C1444 VTAIL.n635 VSUBS 0.02272f
C1445 VTAIL.n636 VSUBS 0.02272f
C1446 VTAIL.n637 VSUBS 0.012209f
C1447 VTAIL.n638 VSUBS 0.012927f
C1448 VTAIL.n639 VSUBS 0.028857f
C1449 VTAIL.n640 VSUBS 0.028857f
C1450 VTAIL.n641 VSUBS 0.012927f
C1451 VTAIL.n642 VSUBS 0.012209f
C1452 VTAIL.n643 VSUBS 0.02272f
C1453 VTAIL.n644 VSUBS 0.02272f
C1454 VTAIL.n645 VSUBS 0.012209f
C1455 VTAIL.n646 VSUBS 0.012927f
C1456 VTAIL.n647 VSUBS 0.028857f
C1457 VTAIL.n648 VSUBS 0.028857f
C1458 VTAIL.n649 VSUBS 0.012927f
C1459 VTAIL.n650 VSUBS 0.012209f
C1460 VTAIL.n651 VSUBS 0.02272f
C1461 VTAIL.n652 VSUBS 0.02272f
C1462 VTAIL.n653 VSUBS 0.012209f
C1463 VTAIL.n654 VSUBS 0.012927f
C1464 VTAIL.n655 VSUBS 0.028857f
C1465 VTAIL.n656 VSUBS 0.028857f
C1466 VTAIL.n657 VSUBS 0.012927f
C1467 VTAIL.n658 VSUBS 0.012209f
C1468 VTAIL.n659 VSUBS 0.02272f
C1469 VTAIL.n660 VSUBS 0.02272f
C1470 VTAIL.n661 VSUBS 0.012209f
C1471 VTAIL.n662 VSUBS 0.012927f
C1472 VTAIL.n663 VSUBS 0.028857f
C1473 VTAIL.n664 VSUBS 0.028857f
C1474 VTAIL.n665 VSUBS 0.012927f
C1475 VTAIL.n666 VSUBS 0.012209f
C1476 VTAIL.n667 VSUBS 0.02272f
C1477 VTAIL.n668 VSUBS 0.02272f
C1478 VTAIL.n669 VSUBS 0.012209f
C1479 VTAIL.n670 VSUBS 0.012209f
C1480 VTAIL.n671 VSUBS 0.012927f
C1481 VTAIL.n672 VSUBS 0.028857f
C1482 VTAIL.n673 VSUBS 0.028857f
C1483 VTAIL.n674 VSUBS 0.028857f
C1484 VTAIL.n675 VSUBS 0.012568f
C1485 VTAIL.n676 VSUBS 0.012209f
C1486 VTAIL.n677 VSUBS 0.02272f
C1487 VTAIL.n678 VSUBS 0.02272f
C1488 VTAIL.n679 VSUBS 0.012209f
C1489 VTAIL.n680 VSUBS 0.012927f
C1490 VTAIL.n681 VSUBS 0.028857f
C1491 VTAIL.n682 VSUBS 0.068552f
C1492 VTAIL.n683 VSUBS 0.012927f
C1493 VTAIL.n684 VSUBS 0.012209f
C1494 VTAIL.n685 VSUBS 0.056551f
C1495 VTAIL.n686 VSUBS 0.034536f
C1496 VTAIL.n687 VSUBS 1.58669f
C1497 VP.t2 VSUBS 3.52416f
C1498 VP.n0 VSUBS 1.34896f
C1499 VP.n1 VSUBS 0.031191f
C1500 VP.n2 VSUBS 0.061992f
C1501 VP.t1 VSUBS 3.80228f
C1502 VP.t0 VSUBS 3.79525f
C1503 VP.n3 VSUBS 4.31006f
C1504 VP.n4 VSUBS 1.87482f
C1505 VP.t3 VSUBS 3.52416f
C1506 VP.n5 VSUBS 1.34896f
C1507 VP.n6 VSUBS 0.057844f
C1508 VP.n7 VSUBS 0.050342f
C1509 VP.n8 VSUBS 0.031191f
C1510 VP.n9 VSUBS 0.031191f
C1511 VP.n10 VSUBS 0.025215f
C1512 VP.n11 VSUBS 0.061992f
C1513 VP.n12 VSUBS 0.057844f
C1514 VP.n13 VSUBS 0.050342f
C1515 VP.n14 VSUBS 0.055668f
.ends

