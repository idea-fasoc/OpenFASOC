* NGSPICE file created from diff_pair_sample_0152.ext - technology: sky130A

.subckt diff_pair_sample_0152 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=0 ps=0 w=13.22 l=1.42
X1 VDD2.t5 VN.t0 VTAIL.t10 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=5.1558 ps=27.22 w=13.22 l=1.42
X2 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=0 ps=0 w=13.22 l=1.42
X3 VTAIL.t6 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=2.1813 ps=13.55 w=13.22 l=1.42
X4 VTAIL.t11 VN.t2 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=2.1813 ps=13.55 w=13.22 l=1.42
X5 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=0 ps=0 w=13.22 l=1.42
X6 VDD1.t5 VP.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=5.1558 ps=27.22 w=13.22 l=1.42
X7 VDD2.t2 VN.t3 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=2.1813 ps=13.55 w=13.22 l=1.42
X8 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=0 ps=0 w=13.22 l=1.42
X9 VDD2.t1 VN.t4 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=5.1558 ps=27.22 w=13.22 l=1.42
X10 VDD1.t4 VP.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=5.1558 ps=27.22 w=13.22 l=1.42
X11 VTAIL.t5 VP.t2 VDD1.t3 B.t4 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=2.1813 ps=13.55 w=13.22 l=1.42
X12 VDD2.t0 VN.t5 VTAIL.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=2.1813 ps=13.55 w=13.22 l=1.42
X13 VDD1.t2 VP.t3 VTAIL.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=2.1813 ps=13.55 w=13.22 l=1.42
X14 VDD1.t1 VP.t4 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=5.1558 pd=27.22 as=2.1813 ps=13.55 w=13.22 l=1.42
X15 VTAIL.t4 VP.t5 VDD1.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=2.1813 pd=13.55 as=2.1813 ps=13.55 w=13.22 l=1.42
R0 B.n739 B.n738 585
R1 B.n305 B.n104 585
R2 B.n304 B.n303 585
R3 B.n302 B.n301 585
R4 B.n300 B.n299 585
R5 B.n298 B.n297 585
R6 B.n296 B.n295 585
R7 B.n294 B.n293 585
R8 B.n292 B.n291 585
R9 B.n290 B.n289 585
R10 B.n288 B.n287 585
R11 B.n286 B.n285 585
R12 B.n284 B.n283 585
R13 B.n282 B.n281 585
R14 B.n280 B.n279 585
R15 B.n278 B.n277 585
R16 B.n276 B.n275 585
R17 B.n274 B.n273 585
R18 B.n272 B.n271 585
R19 B.n270 B.n269 585
R20 B.n268 B.n267 585
R21 B.n266 B.n265 585
R22 B.n264 B.n263 585
R23 B.n262 B.n261 585
R24 B.n260 B.n259 585
R25 B.n258 B.n257 585
R26 B.n256 B.n255 585
R27 B.n254 B.n253 585
R28 B.n252 B.n251 585
R29 B.n250 B.n249 585
R30 B.n248 B.n247 585
R31 B.n246 B.n245 585
R32 B.n244 B.n243 585
R33 B.n242 B.n241 585
R34 B.n240 B.n239 585
R35 B.n238 B.n237 585
R36 B.n236 B.n235 585
R37 B.n234 B.n233 585
R38 B.n232 B.n231 585
R39 B.n230 B.n229 585
R40 B.n228 B.n227 585
R41 B.n226 B.n225 585
R42 B.n224 B.n223 585
R43 B.n222 B.n221 585
R44 B.n220 B.n219 585
R45 B.n217 B.n216 585
R46 B.n215 B.n214 585
R47 B.n213 B.n212 585
R48 B.n211 B.n210 585
R49 B.n209 B.n208 585
R50 B.n207 B.n206 585
R51 B.n205 B.n204 585
R52 B.n203 B.n202 585
R53 B.n201 B.n200 585
R54 B.n199 B.n198 585
R55 B.n196 B.n195 585
R56 B.n194 B.n193 585
R57 B.n192 B.n191 585
R58 B.n190 B.n189 585
R59 B.n188 B.n187 585
R60 B.n186 B.n185 585
R61 B.n184 B.n183 585
R62 B.n182 B.n181 585
R63 B.n180 B.n179 585
R64 B.n178 B.n177 585
R65 B.n176 B.n175 585
R66 B.n174 B.n173 585
R67 B.n172 B.n171 585
R68 B.n170 B.n169 585
R69 B.n168 B.n167 585
R70 B.n166 B.n165 585
R71 B.n164 B.n163 585
R72 B.n162 B.n161 585
R73 B.n160 B.n159 585
R74 B.n158 B.n157 585
R75 B.n156 B.n155 585
R76 B.n154 B.n153 585
R77 B.n152 B.n151 585
R78 B.n150 B.n149 585
R79 B.n148 B.n147 585
R80 B.n146 B.n145 585
R81 B.n144 B.n143 585
R82 B.n142 B.n141 585
R83 B.n140 B.n139 585
R84 B.n138 B.n137 585
R85 B.n136 B.n135 585
R86 B.n134 B.n133 585
R87 B.n132 B.n131 585
R88 B.n130 B.n129 585
R89 B.n128 B.n127 585
R90 B.n126 B.n125 585
R91 B.n124 B.n123 585
R92 B.n122 B.n121 585
R93 B.n120 B.n119 585
R94 B.n118 B.n117 585
R95 B.n116 B.n115 585
R96 B.n114 B.n113 585
R97 B.n112 B.n111 585
R98 B.n110 B.n109 585
R99 B.n53 B.n52 585
R100 B.n737 B.n54 585
R101 B.n742 B.n54 585
R102 B.n736 B.n735 585
R103 B.n735 B.n50 585
R104 B.n734 B.n49 585
R105 B.n748 B.n49 585
R106 B.n733 B.n48 585
R107 B.n749 B.n48 585
R108 B.n732 B.n47 585
R109 B.n750 B.n47 585
R110 B.n731 B.n730 585
R111 B.n730 B.n46 585
R112 B.n729 B.n42 585
R113 B.n756 B.n42 585
R114 B.n728 B.n41 585
R115 B.n757 B.n41 585
R116 B.n727 B.n40 585
R117 B.n758 B.n40 585
R118 B.n726 B.n725 585
R119 B.n725 B.n36 585
R120 B.n724 B.n35 585
R121 B.n764 B.n35 585
R122 B.n723 B.n34 585
R123 B.n765 B.n34 585
R124 B.n722 B.n33 585
R125 B.n766 B.n33 585
R126 B.n721 B.n720 585
R127 B.n720 B.n29 585
R128 B.n719 B.n28 585
R129 B.n772 B.n28 585
R130 B.n718 B.n27 585
R131 B.n773 B.n27 585
R132 B.n717 B.n26 585
R133 B.n774 B.n26 585
R134 B.n716 B.n715 585
R135 B.n715 B.n22 585
R136 B.n714 B.n21 585
R137 B.n780 B.n21 585
R138 B.n713 B.n20 585
R139 B.n781 B.n20 585
R140 B.n712 B.n19 585
R141 B.n782 B.n19 585
R142 B.n711 B.n710 585
R143 B.n710 B.n15 585
R144 B.n709 B.n14 585
R145 B.n788 B.n14 585
R146 B.n708 B.n13 585
R147 B.n789 B.n13 585
R148 B.n707 B.n12 585
R149 B.n790 B.n12 585
R150 B.n706 B.n705 585
R151 B.n705 B.n704 585
R152 B.n703 B.n702 585
R153 B.n703 B.n8 585
R154 B.n701 B.n7 585
R155 B.n797 B.n7 585
R156 B.n700 B.n6 585
R157 B.n798 B.n6 585
R158 B.n699 B.n5 585
R159 B.n799 B.n5 585
R160 B.n698 B.n697 585
R161 B.n697 B.n4 585
R162 B.n696 B.n306 585
R163 B.n696 B.n695 585
R164 B.n686 B.n307 585
R165 B.n308 B.n307 585
R166 B.n688 B.n687 585
R167 B.n689 B.n688 585
R168 B.n685 B.n313 585
R169 B.n313 B.n312 585
R170 B.n684 B.n683 585
R171 B.n683 B.n682 585
R172 B.n315 B.n314 585
R173 B.n316 B.n315 585
R174 B.n675 B.n674 585
R175 B.n676 B.n675 585
R176 B.n673 B.n320 585
R177 B.n324 B.n320 585
R178 B.n672 B.n671 585
R179 B.n671 B.n670 585
R180 B.n322 B.n321 585
R181 B.n323 B.n322 585
R182 B.n663 B.n662 585
R183 B.n664 B.n663 585
R184 B.n661 B.n329 585
R185 B.n329 B.n328 585
R186 B.n660 B.n659 585
R187 B.n659 B.n658 585
R188 B.n331 B.n330 585
R189 B.n332 B.n331 585
R190 B.n651 B.n650 585
R191 B.n652 B.n651 585
R192 B.n649 B.n337 585
R193 B.n337 B.n336 585
R194 B.n648 B.n647 585
R195 B.n647 B.n646 585
R196 B.n339 B.n338 585
R197 B.n340 B.n339 585
R198 B.n639 B.n638 585
R199 B.n640 B.n639 585
R200 B.n637 B.n345 585
R201 B.n345 B.n344 585
R202 B.n636 B.n635 585
R203 B.n635 B.n634 585
R204 B.n347 B.n346 585
R205 B.n627 B.n347 585
R206 B.n626 B.n625 585
R207 B.n628 B.n626 585
R208 B.n624 B.n352 585
R209 B.n352 B.n351 585
R210 B.n623 B.n622 585
R211 B.n622 B.n621 585
R212 B.n354 B.n353 585
R213 B.n355 B.n354 585
R214 B.n614 B.n613 585
R215 B.n615 B.n614 585
R216 B.n358 B.n357 585
R217 B.n417 B.n416 585
R218 B.n418 B.n414 585
R219 B.n414 B.n359 585
R220 B.n420 B.n419 585
R221 B.n422 B.n413 585
R222 B.n425 B.n424 585
R223 B.n426 B.n412 585
R224 B.n428 B.n427 585
R225 B.n430 B.n411 585
R226 B.n433 B.n432 585
R227 B.n434 B.n410 585
R228 B.n436 B.n435 585
R229 B.n438 B.n409 585
R230 B.n441 B.n440 585
R231 B.n442 B.n408 585
R232 B.n444 B.n443 585
R233 B.n446 B.n407 585
R234 B.n449 B.n448 585
R235 B.n450 B.n406 585
R236 B.n452 B.n451 585
R237 B.n454 B.n405 585
R238 B.n457 B.n456 585
R239 B.n458 B.n404 585
R240 B.n460 B.n459 585
R241 B.n462 B.n403 585
R242 B.n465 B.n464 585
R243 B.n466 B.n402 585
R244 B.n468 B.n467 585
R245 B.n470 B.n401 585
R246 B.n473 B.n472 585
R247 B.n474 B.n400 585
R248 B.n476 B.n475 585
R249 B.n478 B.n399 585
R250 B.n481 B.n480 585
R251 B.n482 B.n398 585
R252 B.n484 B.n483 585
R253 B.n486 B.n397 585
R254 B.n489 B.n488 585
R255 B.n490 B.n396 585
R256 B.n492 B.n491 585
R257 B.n494 B.n395 585
R258 B.n497 B.n496 585
R259 B.n498 B.n394 585
R260 B.n500 B.n499 585
R261 B.n502 B.n393 585
R262 B.n505 B.n504 585
R263 B.n506 B.n389 585
R264 B.n508 B.n507 585
R265 B.n510 B.n388 585
R266 B.n513 B.n512 585
R267 B.n514 B.n387 585
R268 B.n516 B.n515 585
R269 B.n518 B.n386 585
R270 B.n521 B.n520 585
R271 B.n522 B.n383 585
R272 B.n525 B.n524 585
R273 B.n527 B.n382 585
R274 B.n530 B.n529 585
R275 B.n531 B.n381 585
R276 B.n533 B.n532 585
R277 B.n535 B.n380 585
R278 B.n538 B.n537 585
R279 B.n539 B.n379 585
R280 B.n541 B.n540 585
R281 B.n543 B.n378 585
R282 B.n546 B.n545 585
R283 B.n547 B.n377 585
R284 B.n549 B.n548 585
R285 B.n551 B.n376 585
R286 B.n554 B.n553 585
R287 B.n555 B.n375 585
R288 B.n557 B.n556 585
R289 B.n559 B.n374 585
R290 B.n562 B.n561 585
R291 B.n563 B.n373 585
R292 B.n565 B.n564 585
R293 B.n567 B.n372 585
R294 B.n570 B.n569 585
R295 B.n571 B.n371 585
R296 B.n573 B.n572 585
R297 B.n575 B.n370 585
R298 B.n578 B.n577 585
R299 B.n579 B.n369 585
R300 B.n581 B.n580 585
R301 B.n583 B.n368 585
R302 B.n586 B.n585 585
R303 B.n587 B.n367 585
R304 B.n589 B.n588 585
R305 B.n591 B.n366 585
R306 B.n594 B.n593 585
R307 B.n595 B.n365 585
R308 B.n597 B.n596 585
R309 B.n599 B.n364 585
R310 B.n602 B.n601 585
R311 B.n603 B.n363 585
R312 B.n605 B.n604 585
R313 B.n607 B.n362 585
R314 B.n608 B.n361 585
R315 B.n611 B.n610 585
R316 B.n612 B.n360 585
R317 B.n360 B.n359 585
R318 B.n617 B.n616 585
R319 B.n616 B.n615 585
R320 B.n618 B.n356 585
R321 B.n356 B.n355 585
R322 B.n620 B.n619 585
R323 B.n621 B.n620 585
R324 B.n350 B.n349 585
R325 B.n351 B.n350 585
R326 B.n630 B.n629 585
R327 B.n629 B.n628 585
R328 B.n631 B.n348 585
R329 B.n627 B.n348 585
R330 B.n633 B.n632 585
R331 B.n634 B.n633 585
R332 B.n343 B.n342 585
R333 B.n344 B.n343 585
R334 B.n642 B.n641 585
R335 B.n641 B.n640 585
R336 B.n643 B.n341 585
R337 B.n341 B.n340 585
R338 B.n645 B.n644 585
R339 B.n646 B.n645 585
R340 B.n335 B.n334 585
R341 B.n336 B.n335 585
R342 B.n654 B.n653 585
R343 B.n653 B.n652 585
R344 B.n655 B.n333 585
R345 B.n333 B.n332 585
R346 B.n657 B.n656 585
R347 B.n658 B.n657 585
R348 B.n327 B.n326 585
R349 B.n328 B.n327 585
R350 B.n666 B.n665 585
R351 B.n665 B.n664 585
R352 B.n667 B.n325 585
R353 B.n325 B.n323 585
R354 B.n669 B.n668 585
R355 B.n670 B.n669 585
R356 B.n319 B.n318 585
R357 B.n324 B.n319 585
R358 B.n678 B.n677 585
R359 B.n677 B.n676 585
R360 B.n679 B.n317 585
R361 B.n317 B.n316 585
R362 B.n681 B.n680 585
R363 B.n682 B.n681 585
R364 B.n311 B.n310 585
R365 B.n312 B.n311 585
R366 B.n691 B.n690 585
R367 B.n690 B.n689 585
R368 B.n692 B.n309 585
R369 B.n309 B.n308 585
R370 B.n694 B.n693 585
R371 B.n695 B.n694 585
R372 B.n3 B.n0 585
R373 B.n4 B.n3 585
R374 B.n796 B.n1 585
R375 B.n797 B.n796 585
R376 B.n795 B.n794 585
R377 B.n795 B.n8 585
R378 B.n793 B.n9 585
R379 B.n704 B.n9 585
R380 B.n792 B.n791 585
R381 B.n791 B.n790 585
R382 B.n11 B.n10 585
R383 B.n789 B.n11 585
R384 B.n787 B.n786 585
R385 B.n788 B.n787 585
R386 B.n785 B.n16 585
R387 B.n16 B.n15 585
R388 B.n784 B.n783 585
R389 B.n783 B.n782 585
R390 B.n18 B.n17 585
R391 B.n781 B.n18 585
R392 B.n779 B.n778 585
R393 B.n780 B.n779 585
R394 B.n777 B.n23 585
R395 B.n23 B.n22 585
R396 B.n776 B.n775 585
R397 B.n775 B.n774 585
R398 B.n25 B.n24 585
R399 B.n773 B.n25 585
R400 B.n771 B.n770 585
R401 B.n772 B.n771 585
R402 B.n769 B.n30 585
R403 B.n30 B.n29 585
R404 B.n768 B.n767 585
R405 B.n767 B.n766 585
R406 B.n32 B.n31 585
R407 B.n765 B.n32 585
R408 B.n763 B.n762 585
R409 B.n764 B.n763 585
R410 B.n761 B.n37 585
R411 B.n37 B.n36 585
R412 B.n760 B.n759 585
R413 B.n759 B.n758 585
R414 B.n39 B.n38 585
R415 B.n757 B.n39 585
R416 B.n755 B.n754 585
R417 B.n756 B.n755 585
R418 B.n753 B.n43 585
R419 B.n46 B.n43 585
R420 B.n752 B.n751 585
R421 B.n751 B.n750 585
R422 B.n45 B.n44 585
R423 B.n749 B.n45 585
R424 B.n747 B.n746 585
R425 B.n748 B.n747 585
R426 B.n745 B.n51 585
R427 B.n51 B.n50 585
R428 B.n744 B.n743 585
R429 B.n743 B.n742 585
R430 B.n800 B.n799 585
R431 B.n798 B.n2 585
R432 B.n743 B.n53 530.939
R433 B.n739 B.n54 530.939
R434 B.n614 B.n360 530.939
R435 B.n616 B.n358 530.939
R436 B.n107 B.t17 429.497
R437 B.n105 B.t6 429.497
R438 B.n384 B.t10 429.497
R439 B.n390 B.t14 429.497
R440 B.n741 B.n740 256.663
R441 B.n741 B.n103 256.663
R442 B.n741 B.n102 256.663
R443 B.n741 B.n101 256.663
R444 B.n741 B.n100 256.663
R445 B.n741 B.n99 256.663
R446 B.n741 B.n98 256.663
R447 B.n741 B.n97 256.663
R448 B.n741 B.n96 256.663
R449 B.n741 B.n95 256.663
R450 B.n741 B.n94 256.663
R451 B.n741 B.n93 256.663
R452 B.n741 B.n92 256.663
R453 B.n741 B.n91 256.663
R454 B.n741 B.n90 256.663
R455 B.n741 B.n89 256.663
R456 B.n741 B.n88 256.663
R457 B.n741 B.n87 256.663
R458 B.n741 B.n86 256.663
R459 B.n741 B.n85 256.663
R460 B.n741 B.n84 256.663
R461 B.n741 B.n83 256.663
R462 B.n741 B.n82 256.663
R463 B.n741 B.n81 256.663
R464 B.n741 B.n80 256.663
R465 B.n741 B.n79 256.663
R466 B.n741 B.n78 256.663
R467 B.n741 B.n77 256.663
R468 B.n741 B.n76 256.663
R469 B.n741 B.n75 256.663
R470 B.n741 B.n74 256.663
R471 B.n741 B.n73 256.663
R472 B.n741 B.n72 256.663
R473 B.n741 B.n71 256.663
R474 B.n741 B.n70 256.663
R475 B.n741 B.n69 256.663
R476 B.n741 B.n68 256.663
R477 B.n741 B.n67 256.663
R478 B.n741 B.n66 256.663
R479 B.n741 B.n65 256.663
R480 B.n741 B.n64 256.663
R481 B.n741 B.n63 256.663
R482 B.n741 B.n62 256.663
R483 B.n741 B.n61 256.663
R484 B.n741 B.n60 256.663
R485 B.n741 B.n59 256.663
R486 B.n741 B.n58 256.663
R487 B.n741 B.n57 256.663
R488 B.n741 B.n56 256.663
R489 B.n741 B.n55 256.663
R490 B.n415 B.n359 256.663
R491 B.n421 B.n359 256.663
R492 B.n423 B.n359 256.663
R493 B.n429 B.n359 256.663
R494 B.n431 B.n359 256.663
R495 B.n437 B.n359 256.663
R496 B.n439 B.n359 256.663
R497 B.n445 B.n359 256.663
R498 B.n447 B.n359 256.663
R499 B.n453 B.n359 256.663
R500 B.n455 B.n359 256.663
R501 B.n461 B.n359 256.663
R502 B.n463 B.n359 256.663
R503 B.n469 B.n359 256.663
R504 B.n471 B.n359 256.663
R505 B.n477 B.n359 256.663
R506 B.n479 B.n359 256.663
R507 B.n485 B.n359 256.663
R508 B.n487 B.n359 256.663
R509 B.n493 B.n359 256.663
R510 B.n495 B.n359 256.663
R511 B.n501 B.n359 256.663
R512 B.n503 B.n359 256.663
R513 B.n509 B.n359 256.663
R514 B.n511 B.n359 256.663
R515 B.n517 B.n359 256.663
R516 B.n519 B.n359 256.663
R517 B.n526 B.n359 256.663
R518 B.n528 B.n359 256.663
R519 B.n534 B.n359 256.663
R520 B.n536 B.n359 256.663
R521 B.n542 B.n359 256.663
R522 B.n544 B.n359 256.663
R523 B.n550 B.n359 256.663
R524 B.n552 B.n359 256.663
R525 B.n558 B.n359 256.663
R526 B.n560 B.n359 256.663
R527 B.n566 B.n359 256.663
R528 B.n568 B.n359 256.663
R529 B.n574 B.n359 256.663
R530 B.n576 B.n359 256.663
R531 B.n582 B.n359 256.663
R532 B.n584 B.n359 256.663
R533 B.n590 B.n359 256.663
R534 B.n592 B.n359 256.663
R535 B.n598 B.n359 256.663
R536 B.n600 B.n359 256.663
R537 B.n606 B.n359 256.663
R538 B.n609 B.n359 256.663
R539 B.n802 B.n801 256.663
R540 B.n111 B.n110 163.367
R541 B.n115 B.n114 163.367
R542 B.n119 B.n118 163.367
R543 B.n123 B.n122 163.367
R544 B.n127 B.n126 163.367
R545 B.n131 B.n130 163.367
R546 B.n135 B.n134 163.367
R547 B.n139 B.n138 163.367
R548 B.n143 B.n142 163.367
R549 B.n147 B.n146 163.367
R550 B.n151 B.n150 163.367
R551 B.n155 B.n154 163.367
R552 B.n159 B.n158 163.367
R553 B.n163 B.n162 163.367
R554 B.n167 B.n166 163.367
R555 B.n171 B.n170 163.367
R556 B.n175 B.n174 163.367
R557 B.n179 B.n178 163.367
R558 B.n183 B.n182 163.367
R559 B.n187 B.n186 163.367
R560 B.n191 B.n190 163.367
R561 B.n195 B.n194 163.367
R562 B.n200 B.n199 163.367
R563 B.n204 B.n203 163.367
R564 B.n208 B.n207 163.367
R565 B.n212 B.n211 163.367
R566 B.n216 B.n215 163.367
R567 B.n221 B.n220 163.367
R568 B.n225 B.n224 163.367
R569 B.n229 B.n228 163.367
R570 B.n233 B.n232 163.367
R571 B.n237 B.n236 163.367
R572 B.n241 B.n240 163.367
R573 B.n245 B.n244 163.367
R574 B.n249 B.n248 163.367
R575 B.n253 B.n252 163.367
R576 B.n257 B.n256 163.367
R577 B.n261 B.n260 163.367
R578 B.n265 B.n264 163.367
R579 B.n269 B.n268 163.367
R580 B.n273 B.n272 163.367
R581 B.n277 B.n276 163.367
R582 B.n281 B.n280 163.367
R583 B.n285 B.n284 163.367
R584 B.n289 B.n288 163.367
R585 B.n293 B.n292 163.367
R586 B.n297 B.n296 163.367
R587 B.n301 B.n300 163.367
R588 B.n303 B.n104 163.367
R589 B.n614 B.n354 163.367
R590 B.n622 B.n354 163.367
R591 B.n622 B.n352 163.367
R592 B.n626 B.n352 163.367
R593 B.n626 B.n347 163.367
R594 B.n635 B.n347 163.367
R595 B.n635 B.n345 163.367
R596 B.n639 B.n345 163.367
R597 B.n639 B.n339 163.367
R598 B.n647 B.n339 163.367
R599 B.n647 B.n337 163.367
R600 B.n651 B.n337 163.367
R601 B.n651 B.n331 163.367
R602 B.n659 B.n331 163.367
R603 B.n659 B.n329 163.367
R604 B.n663 B.n329 163.367
R605 B.n663 B.n322 163.367
R606 B.n671 B.n322 163.367
R607 B.n671 B.n320 163.367
R608 B.n675 B.n320 163.367
R609 B.n675 B.n315 163.367
R610 B.n683 B.n315 163.367
R611 B.n683 B.n313 163.367
R612 B.n688 B.n313 163.367
R613 B.n688 B.n307 163.367
R614 B.n696 B.n307 163.367
R615 B.n697 B.n696 163.367
R616 B.n697 B.n5 163.367
R617 B.n6 B.n5 163.367
R618 B.n7 B.n6 163.367
R619 B.n703 B.n7 163.367
R620 B.n705 B.n703 163.367
R621 B.n705 B.n12 163.367
R622 B.n13 B.n12 163.367
R623 B.n14 B.n13 163.367
R624 B.n710 B.n14 163.367
R625 B.n710 B.n19 163.367
R626 B.n20 B.n19 163.367
R627 B.n21 B.n20 163.367
R628 B.n715 B.n21 163.367
R629 B.n715 B.n26 163.367
R630 B.n27 B.n26 163.367
R631 B.n28 B.n27 163.367
R632 B.n720 B.n28 163.367
R633 B.n720 B.n33 163.367
R634 B.n34 B.n33 163.367
R635 B.n35 B.n34 163.367
R636 B.n725 B.n35 163.367
R637 B.n725 B.n40 163.367
R638 B.n41 B.n40 163.367
R639 B.n42 B.n41 163.367
R640 B.n730 B.n42 163.367
R641 B.n730 B.n47 163.367
R642 B.n48 B.n47 163.367
R643 B.n49 B.n48 163.367
R644 B.n735 B.n49 163.367
R645 B.n735 B.n54 163.367
R646 B.n416 B.n414 163.367
R647 B.n420 B.n414 163.367
R648 B.n424 B.n422 163.367
R649 B.n428 B.n412 163.367
R650 B.n432 B.n430 163.367
R651 B.n436 B.n410 163.367
R652 B.n440 B.n438 163.367
R653 B.n444 B.n408 163.367
R654 B.n448 B.n446 163.367
R655 B.n452 B.n406 163.367
R656 B.n456 B.n454 163.367
R657 B.n460 B.n404 163.367
R658 B.n464 B.n462 163.367
R659 B.n468 B.n402 163.367
R660 B.n472 B.n470 163.367
R661 B.n476 B.n400 163.367
R662 B.n480 B.n478 163.367
R663 B.n484 B.n398 163.367
R664 B.n488 B.n486 163.367
R665 B.n492 B.n396 163.367
R666 B.n496 B.n494 163.367
R667 B.n500 B.n394 163.367
R668 B.n504 B.n502 163.367
R669 B.n508 B.n389 163.367
R670 B.n512 B.n510 163.367
R671 B.n516 B.n387 163.367
R672 B.n520 B.n518 163.367
R673 B.n525 B.n383 163.367
R674 B.n529 B.n527 163.367
R675 B.n533 B.n381 163.367
R676 B.n537 B.n535 163.367
R677 B.n541 B.n379 163.367
R678 B.n545 B.n543 163.367
R679 B.n549 B.n377 163.367
R680 B.n553 B.n551 163.367
R681 B.n557 B.n375 163.367
R682 B.n561 B.n559 163.367
R683 B.n565 B.n373 163.367
R684 B.n569 B.n567 163.367
R685 B.n573 B.n371 163.367
R686 B.n577 B.n575 163.367
R687 B.n581 B.n369 163.367
R688 B.n585 B.n583 163.367
R689 B.n589 B.n367 163.367
R690 B.n593 B.n591 163.367
R691 B.n597 B.n365 163.367
R692 B.n601 B.n599 163.367
R693 B.n605 B.n363 163.367
R694 B.n608 B.n607 163.367
R695 B.n610 B.n360 163.367
R696 B.n616 B.n356 163.367
R697 B.n620 B.n356 163.367
R698 B.n620 B.n350 163.367
R699 B.n629 B.n350 163.367
R700 B.n629 B.n348 163.367
R701 B.n633 B.n348 163.367
R702 B.n633 B.n343 163.367
R703 B.n641 B.n343 163.367
R704 B.n641 B.n341 163.367
R705 B.n645 B.n341 163.367
R706 B.n645 B.n335 163.367
R707 B.n653 B.n335 163.367
R708 B.n653 B.n333 163.367
R709 B.n657 B.n333 163.367
R710 B.n657 B.n327 163.367
R711 B.n665 B.n327 163.367
R712 B.n665 B.n325 163.367
R713 B.n669 B.n325 163.367
R714 B.n669 B.n319 163.367
R715 B.n677 B.n319 163.367
R716 B.n677 B.n317 163.367
R717 B.n681 B.n317 163.367
R718 B.n681 B.n311 163.367
R719 B.n690 B.n311 163.367
R720 B.n690 B.n309 163.367
R721 B.n694 B.n309 163.367
R722 B.n694 B.n3 163.367
R723 B.n800 B.n3 163.367
R724 B.n796 B.n2 163.367
R725 B.n796 B.n795 163.367
R726 B.n795 B.n9 163.367
R727 B.n791 B.n9 163.367
R728 B.n791 B.n11 163.367
R729 B.n787 B.n11 163.367
R730 B.n787 B.n16 163.367
R731 B.n783 B.n16 163.367
R732 B.n783 B.n18 163.367
R733 B.n779 B.n18 163.367
R734 B.n779 B.n23 163.367
R735 B.n775 B.n23 163.367
R736 B.n775 B.n25 163.367
R737 B.n771 B.n25 163.367
R738 B.n771 B.n30 163.367
R739 B.n767 B.n30 163.367
R740 B.n767 B.n32 163.367
R741 B.n763 B.n32 163.367
R742 B.n763 B.n37 163.367
R743 B.n759 B.n37 163.367
R744 B.n759 B.n39 163.367
R745 B.n755 B.n39 163.367
R746 B.n755 B.n43 163.367
R747 B.n751 B.n43 163.367
R748 B.n751 B.n45 163.367
R749 B.n747 B.n45 163.367
R750 B.n747 B.n51 163.367
R751 B.n743 B.n51 163.367
R752 B.n105 B.t8 107.397
R753 B.n384 B.t13 107.397
R754 B.n107 B.t18 107.379
R755 B.n390 B.t16 107.379
R756 B.n615 B.n359 81.482
R757 B.n742 B.n741 81.482
R758 B.n106 B.t9 73.4573
R759 B.n385 B.t12 73.4573
R760 B.n108 B.t19 73.4406
R761 B.n391 B.t15 73.4406
R762 B.n55 B.n53 71.676
R763 B.n111 B.n56 71.676
R764 B.n115 B.n57 71.676
R765 B.n119 B.n58 71.676
R766 B.n123 B.n59 71.676
R767 B.n127 B.n60 71.676
R768 B.n131 B.n61 71.676
R769 B.n135 B.n62 71.676
R770 B.n139 B.n63 71.676
R771 B.n143 B.n64 71.676
R772 B.n147 B.n65 71.676
R773 B.n151 B.n66 71.676
R774 B.n155 B.n67 71.676
R775 B.n159 B.n68 71.676
R776 B.n163 B.n69 71.676
R777 B.n167 B.n70 71.676
R778 B.n171 B.n71 71.676
R779 B.n175 B.n72 71.676
R780 B.n179 B.n73 71.676
R781 B.n183 B.n74 71.676
R782 B.n187 B.n75 71.676
R783 B.n191 B.n76 71.676
R784 B.n195 B.n77 71.676
R785 B.n200 B.n78 71.676
R786 B.n204 B.n79 71.676
R787 B.n208 B.n80 71.676
R788 B.n212 B.n81 71.676
R789 B.n216 B.n82 71.676
R790 B.n221 B.n83 71.676
R791 B.n225 B.n84 71.676
R792 B.n229 B.n85 71.676
R793 B.n233 B.n86 71.676
R794 B.n237 B.n87 71.676
R795 B.n241 B.n88 71.676
R796 B.n245 B.n89 71.676
R797 B.n249 B.n90 71.676
R798 B.n253 B.n91 71.676
R799 B.n257 B.n92 71.676
R800 B.n261 B.n93 71.676
R801 B.n265 B.n94 71.676
R802 B.n269 B.n95 71.676
R803 B.n273 B.n96 71.676
R804 B.n277 B.n97 71.676
R805 B.n281 B.n98 71.676
R806 B.n285 B.n99 71.676
R807 B.n289 B.n100 71.676
R808 B.n293 B.n101 71.676
R809 B.n297 B.n102 71.676
R810 B.n301 B.n103 71.676
R811 B.n740 B.n104 71.676
R812 B.n740 B.n739 71.676
R813 B.n303 B.n103 71.676
R814 B.n300 B.n102 71.676
R815 B.n296 B.n101 71.676
R816 B.n292 B.n100 71.676
R817 B.n288 B.n99 71.676
R818 B.n284 B.n98 71.676
R819 B.n280 B.n97 71.676
R820 B.n276 B.n96 71.676
R821 B.n272 B.n95 71.676
R822 B.n268 B.n94 71.676
R823 B.n264 B.n93 71.676
R824 B.n260 B.n92 71.676
R825 B.n256 B.n91 71.676
R826 B.n252 B.n90 71.676
R827 B.n248 B.n89 71.676
R828 B.n244 B.n88 71.676
R829 B.n240 B.n87 71.676
R830 B.n236 B.n86 71.676
R831 B.n232 B.n85 71.676
R832 B.n228 B.n84 71.676
R833 B.n224 B.n83 71.676
R834 B.n220 B.n82 71.676
R835 B.n215 B.n81 71.676
R836 B.n211 B.n80 71.676
R837 B.n207 B.n79 71.676
R838 B.n203 B.n78 71.676
R839 B.n199 B.n77 71.676
R840 B.n194 B.n76 71.676
R841 B.n190 B.n75 71.676
R842 B.n186 B.n74 71.676
R843 B.n182 B.n73 71.676
R844 B.n178 B.n72 71.676
R845 B.n174 B.n71 71.676
R846 B.n170 B.n70 71.676
R847 B.n166 B.n69 71.676
R848 B.n162 B.n68 71.676
R849 B.n158 B.n67 71.676
R850 B.n154 B.n66 71.676
R851 B.n150 B.n65 71.676
R852 B.n146 B.n64 71.676
R853 B.n142 B.n63 71.676
R854 B.n138 B.n62 71.676
R855 B.n134 B.n61 71.676
R856 B.n130 B.n60 71.676
R857 B.n126 B.n59 71.676
R858 B.n122 B.n58 71.676
R859 B.n118 B.n57 71.676
R860 B.n114 B.n56 71.676
R861 B.n110 B.n55 71.676
R862 B.n415 B.n358 71.676
R863 B.n421 B.n420 71.676
R864 B.n424 B.n423 71.676
R865 B.n429 B.n428 71.676
R866 B.n432 B.n431 71.676
R867 B.n437 B.n436 71.676
R868 B.n440 B.n439 71.676
R869 B.n445 B.n444 71.676
R870 B.n448 B.n447 71.676
R871 B.n453 B.n452 71.676
R872 B.n456 B.n455 71.676
R873 B.n461 B.n460 71.676
R874 B.n464 B.n463 71.676
R875 B.n469 B.n468 71.676
R876 B.n472 B.n471 71.676
R877 B.n477 B.n476 71.676
R878 B.n480 B.n479 71.676
R879 B.n485 B.n484 71.676
R880 B.n488 B.n487 71.676
R881 B.n493 B.n492 71.676
R882 B.n496 B.n495 71.676
R883 B.n501 B.n500 71.676
R884 B.n504 B.n503 71.676
R885 B.n509 B.n508 71.676
R886 B.n512 B.n511 71.676
R887 B.n517 B.n516 71.676
R888 B.n520 B.n519 71.676
R889 B.n526 B.n525 71.676
R890 B.n529 B.n528 71.676
R891 B.n534 B.n533 71.676
R892 B.n537 B.n536 71.676
R893 B.n542 B.n541 71.676
R894 B.n545 B.n544 71.676
R895 B.n550 B.n549 71.676
R896 B.n553 B.n552 71.676
R897 B.n558 B.n557 71.676
R898 B.n561 B.n560 71.676
R899 B.n566 B.n565 71.676
R900 B.n569 B.n568 71.676
R901 B.n574 B.n573 71.676
R902 B.n577 B.n576 71.676
R903 B.n582 B.n581 71.676
R904 B.n585 B.n584 71.676
R905 B.n590 B.n589 71.676
R906 B.n593 B.n592 71.676
R907 B.n598 B.n597 71.676
R908 B.n601 B.n600 71.676
R909 B.n606 B.n605 71.676
R910 B.n609 B.n608 71.676
R911 B.n416 B.n415 71.676
R912 B.n422 B.n421 71.676
R913 B.n423 B.n412 71.676
R914 B.n430 B.n429 71.676
R915 B.n431 B.n410 71.676
R916 B.n438 B.n437 71.676
R917 B.n439 B.n408 71.676
R918 B.n446 B.n445 71.676
R919 B.n447 B.n406 71.676
R920 B.n454 B.n453 71.676
R921 B.n455 B.n404 71.676
R922 B.n462 B.n461 71.676
R923 B.n463 B.n402 71.676
R924 B.n470 B.n469 71.676
R925 B.n471 B.n400 71.676
R926 B.n478 B.n477 71.676
R927 B.n479 B.n398 71.676
R928 B.n486 B.n485 71.676
R929 B.n487 B.n396 71.676
R930 B.n494 B.n493 71.676
R931 B.n495 B.n394 71.676
R932 B.n502 B.n501 71.676
R933 B.n503 B.n389 71.676
R934 B.n510 B.n509 71.676
R935 B.n511 B.n387 71.676
R936 B.n518 B.n517 71.676
R937 B.n519 B.n383 71.676
R938 B.n527 B.n526 71.676
R939 B.n528 B.n381 71.676
R940 B.n535 B.n534 71.676
R941 B.n536 B.n379 71.676
R942 B.n543 B.n542 71.676
R943 B.n544 B.n377 71.676
R944 B.n551 B.n550 71.676
R945 B.n552 B.n375 71.676
R946 B.n559 B.n558 71.676
R947 B.n560 B.n373 71.676
R948 B.n567 B.n566 71.676
R949 B.n568 B.n371 71.676
R950 B.n575 B.n574 71.676
R951 B.n576 B.n369 71.676
R952 B.n583 B.n582 71.676
R953 B.n584 B.n367 71.676
R954 B.n591 B.n590 71.676
R955 B.n592 B.n365 71.676
R956 B.n599 B.n598 71.676
R957 B.n600 B.n363 71.676
R958 B.n607 B.n606 71.676
R959 B.n610 B.n609 71.676
R960 B.n801 B.n800 71.676
R961 B.n801 B.n2 71.676
R962 B.n197 B.n108 59.5399
R963 B.n218 B.n106 59.5399
R964 B.n523 B.n385 59.5399
R965 B.n392 B.n391 59.5399
R966 B.n615 B.n355 40.4439
R967 B.n621 B.n355 40.4439
R968 B.n621 B.n351 40.4439
R969 B.n628 B.n351 40.4439
R970 B.n628 B.n627 40.4439
R971 B.n634 B.n344 40.4439
R972 B.n640 B.n344 40.4439
R973 B.n640 B.n340 40.4439
R974 B.n646 B.n340 40.4439
R975 B.n646 B.n336 40.4439
R976 B.n652 B.n336 40.4439
R977 B.n652 B.n332 40.4439
R978 B.n658 B.n332 40.4439
R979 B.n664 B.n328 40.4439
R980 B.n664 B.n323 40.4439
R981 B.n670 B.n323 40.4439
R982 B.n670 B.n324 40.4439
R983 B.n676 B.n316 40.4439
R984 B.n682 B.n316 40.4439
R985 B.n682 B.n312 40.4439
R986 B.n689 B.n312 40.4439
R987 B.n695 B.n308 40.4439
R988 B.n695 B.n4 40.4439
R989 B.n799 B.n4 40.4439
R990 B.n799 B.n798 40.4439
R991 B.n798 B.n797 40.4439
R992 B.n797 B.n8 40.4439
R993 B.n704 B.n8 40.4439
R994 B.n790 B.n789 40.4439
R995 B.n789 B.n788 40.4439
R996 B.n788 B.n15 40.4439
R997 B.n782 B.n15 40.4439
R998 B.n781 B.n780 40.4439
R999 B.n780 B.n22 40.4439
R1000 B.n774 B.n22 40.4439
R1001 B.n774 B.n773 40.4439
R1002 B.n772 B.n29 40.4439
R1003 B.n766 B.n29 40.4439
R1004 B.n766 B.n765 40.4439
R1005 B.n765 B.n764 40.4439
R1006 B.n764 B.n36 40.4439
R1007 B.n758 B.n36 40.4439
R1008 B.n758 B.n757 40.4439
R1009 B.n757 B.n756 40.4439
R1010 B.n750 B.n46 40.4439
R1011 B.n750 B.n749 40.4439
R1012 B.n749 B.n748 40.4439
R1013 B.n748 B.n50 40.4439
R1014 B.n742 B.n50 40.4439
R1015 B.t0 B.n328 39.2544
R1016 B.n773 B.t1 39.2544
R1017 B.n617 B.n357 34.4981
R1018 B.n613 B.n612 34.4981
R1019 B.n738 B.n737 34.4981
R1020 B.n744 B.n52 34.4981
R1021 B.n108 B.n107 33.9399
R1022 B.n106 B.n105 33.9399
R1023 B.n385 B.n384 33.9399
R1024 B.n391 B.n390 33.9399
R1025 B.n676 B.t3 33.3068
R1026 B.n782 B.t4 33.3068
R1027 B.n627 B.t11 27.3592
R1028 B.t2 B.n308 27.3592
R1029 B.n704 B.t5 27.3592
R1030 B.n46 B.t7 27.3592
R1031 B B.n802 18.0485
R1032 B.n634 B.t11 13.0851
R1033 B.n689 B.t2 13.0851
R1034 B.n790 B.t5 13.0851
R1035 B.n756 B.t7 13.0851
R1036 B.n618 B.n617 10.6151
R1037 B.n619 B.n618 10.6151
R1038 B.n619 B.n349 10.6151
R1039 B.n630 B.n349 10.6151
R1040 B.n631 B.n630 10.6151
R1041 B.n632 B.n631 10.6151
R1042 B.n632 B.n342 10.6151
R1043 B.n642 B.n342 10.6151
R1044 B.n643 B.n642 10.6151
R1045 B.n644 B.n643 10.6151
R1046 B.n644 B.n334 10.6151
R1047 B.n654 B.n334 10.6151
R1048 B.n655 B.n654 10.6151
R1049 B.n656 B.n655 10.6151
R1050 B.n656 B.n326 10.6151
R1051 B.n666 B.n326 10.6151
R1052 B.n667 B.n666 10.6151
R1053 B.n668 B.n667 10.6151
R1054 B.n668 B.n318 10.6151
R1055 B.n678 B.n318 10.6151
R1056 B.n679 B.n678 10.6151
R1057 B.n680 B.n679 10.6151
R1058 B.n680 B.n310 10.6151
R1059 B.n691 B.n310 10.6151
R1060 B.n692 B.n691 10.6151
R1061 B.n693 B.n692 10.6151
R1062 B.n693 B.n0 10.6151
R1063 B.n417 B.n357 10.6151
R1064 B.n418 B.n417 10.6151
R1065 B.n419 B.n418 10.6151
R1066 B.n419 B.n413 10.6151
R1067 B.n425 B.n413 10.6151
R1068 B.n426 B.n425 10.6151
R1069 B.n427 B.n426 10.6151
R1070 B.n427 B.n411 10.6151
R1071 B.n433 B.n411 10.6151
R1072 B.n434 B.n433 10.6151
R1073 B.n435 B.n434 10.6151
R1074 B.n435 B.n409 10.6151
R1075 B.n441 B.n409 10.6151
R1076 B.n442 B.n441 10.6151
R1077 B.n443 B.n442 10.6151
R1078 B.n443 B.n407 10.6151
R1079 B.n449 B.n407 10.6151
R1080 B.n450 B.n449 10.6151
R1081 B.n451 B.n450 10.6151
R1082 B.n451 B.n405 10.6151
R1083 B.n457 B.n405 10.6151
R1084 B.n458 B.n457 10.6151
R1085 B.n459 B.n458 10.6151
R1086 B.n459 B.n403 10.6151
R1087 B.n465 B.n403 10.6151
R1088 B.n466 B.n465 10.6151
R1089 B.n467 B.n466 10.6151
R1090 B.n467 B.n401 10.6151
R1091 B.n473 B.n401 10.6151
R1092 B.n474 B.n473 10.6151
R1093 B.n475 B.n474 10.6151
R1094 B.n475 B.n399 10.6151
R1095 B.n481 B.n399 10.6151
R1096 B.n482 B.n481 10.6151
R1097 B.n483 B.n482 10.6151
R1098 B.n483 B.n397 10.6151
R1099 B.n489 B.n397 10.6151
R1100 B.n490 B.n489 10.6151
R1101 B.n491 B.n490 10.6151
R1102 B.n491 B.n395 10.6151
R1103 B.n497 B.n395 10.6151
R1104 B.n498 B.n497 10.6151
R1105 B.n499 B.n498 10.6151
R1106 B.n499 B.n393 10.6151
R1107 B.n506 B.n505 10.6151
R1108 B.n507 B.n506 10.6151
R1109 B.n507 B.n388 10.6151
R1110 B.n513 B.n388 10.6151
R1111 B.n514 B.n513 10.6151
R1112 B.n515 B.n514 10.6151
R1113 B.n515 B.n386 10.6151
R1114 B.n521 B.n386 10.6151
R1115 B.n522 B.n521 10.6151
R1116 B.n524 B.n382 10.6151
R1117 B.n530 B.n382 10.6151
R1118 B.n531 B.n530 10.6151
R1119 B.n532 B.n531 10.6151
R1120 B.n532 B.n380 10.6151
R1121 B.n538 B.n380 10.6151
R1122 B.n539 B.n538 10.6151
R1123 B.n540 B.n539 10.6151
R1124 B.n540 B.n378 10.6151
R1125 B.n546 B.n378 10.6151
R1126 B.n547 B.n546 10.6151
R1127 B.n548 B.n547 10.6151
R1128 B.n548 B.n376 10.6151
R1129 B.n554 B.n376 10.6151
R1130 B.n555 B.n554 10.6151
R1131 B.n556 B.n555 10.6151
R1132 B.n556 B.n374 10.6151
R1133 B.n562 B.n374 10.6151
R1134 B.n563 B.n562 10.6151
R1135 B.n564 B.n563 10.6151
R1136 B.n564 B.n372 10.6151
R1137 B.n570 B.n372 10.6151
R1138 B.n571 B.n570 10.6151
R1139 B.n572 B.n571 10.6151
R1140 B.n572 B.n370 10.6151
R1141 B.n578 B.n370 10.6151
R1142 B.n579 B.n578 10.6151
R1143 B.n580 B.n579 10.6151
R1144 B.n580 B.n368 10.6151
R1145 B.n586 B.n368 10.6151
R1146 B.n587 B.n586 10.6151
R1147 B.n588 B.n587 10.6151
R1148 B.n588 B.n366 10.6151
R1149 B.n594 B.n366 10.6151
R1150 B.n595 B.n594 10.6151
R1151 B.n596 B.n595 10.6151
R1152 B.n596 B.n364 10.6151
R1153 B.n602 B.n364 10.6151
R1154 B.n603 B.n602 10.6151
R1155 B.n604 B.n603 10.6151
R1156 B.n604 B.n362 10.6151
R1157 B.n362 B.n361 10.6151
R1158 B.n611 B.n361 10.6151
R1159 B.n612 B.n611 10.6151
R1160 B.n613 B.n353 10.6151
R1161 B.n623 B.n353 10.6151
R1162 B.n624 B.n623 10.6151
R1163 B.n625 B.n624 10.6151
R1164 B.n625 B.n346 10.6151
R1165 B.n636 B.n346 10.6151
R1166 B.n637 B.n636 10.6151
R1167 B.n638 B.n637 10.6151
R1168 B.n638 B.n338 10.6151
R1169 B.n648 B.n338 10.6151
R1170 B.n649 B.n648 10.6151
R1171 B.n650 B.n649 10.6151
R1172 B.n650 B.n330 10.6151
R1173 B.n660 B.n330 10.6151
R1174 B.n661 B.n660 10.6151
R1175 B.n662 B.n661 10.6151
R1176 B.n662 B.n321 10.6151
R1177 B.n672 B.n321 10.6151
R1178 B.n673 B.n672 10.6151
R1179 B.n674 B.n673 10.6151
R1180 B.n674 B.n314 10.6151
R1181 B.n684 B.n314 10.6151
R1182 B.n685 B.n684 10.6151
R1183 B.n687 B.n685 10.6151
R1184 B.n687 B.n686 10.6151
R1185 B.n686 B.n306 10.6151
R1186 B.n698 B.n306 10.6151
R1187 B.n699 B.n698 10.6151
R1188 B.n700 B.n699 10.6151
R1189 B.n701 B.n700 10.6151
R1190 B.n702 B.n701 10.6151
R1191 B.n706 B.n702 10.6151
R1192 B.n707 B.n706 10.6151
R1193 B.n708 B.n707 10.6151
R1194 B.n709 B.n708 10.6151
R1195 B.n711 B.n709 10.6151
R1196 B.n712 B.n711 10.6151
R1197 B.n713 B.n712 10.6151
R1198 B.n714 B.n713 10.6151
R1199 B.n716 B.n714 10.6151
R1200 B.n717 B.n716 10.6151
R1201 B.n718 B.n717 10.6151
R1202 B.n719 B.n718 10.6151
R1203 B.n721 B.n719 10.6151
R1204 B.n722 B.n721 10.6151
R1205 B.n723 B.n722 10.6151
R1206 B.n724 B.n723 10.6151
R1207 B.n726 B.n724 10.6151
R1208 B.n727 B.n726 10.6151
R1209 B.n728 B.n727 10.6151
R1210 B.n729 B.n728 10.6151
R1211 B.n731 B.n729 10.6151
R1212 B.n732 B.n731 10.6151
R1213 B.n733 B.n732 10.6151
R1214 B.n734 B.n733 10.6151
R1215 B.n736 B.n734 10.6151
R1216 B.n737 B.n736 10.6151
R1217 B.n794 B.n1 10.6151
R1218 B.n794 B.n793 10.6151
R1219 B.n793 B.n792 10.6151
R1220 B.n792 B.n10 10.6151
R1221 B.n786 B.n10 10.6151
R1222 B.n786 B.n785 10.6151
R1223 B.n785 B.n784 10.6151
R1224 B.n784 B.n17 10.6151
R1225 B.n778 B.n17 10.6151
R1226 B.n778 B.n777 10.6151
R1227 B.n777 B.n776 10.6151
R1228 B.n776 B.n24 10.6151
R1229 B.n770 B.n24 10.6151
R1230 B.n770 B.n769 10.6151
R1231 B.n769 B.n768 10.6151
R1232 B.n768 B.n31 10.6151
R1233 B.n762 B.n31 10.6151
R1234 B.n762 B.n761 10.6151
R1235 B.n761 B.n760 10.6151
R1236 B.n760 B.n38 10.6151
R1237 B.n754 B.n38 10.6151
R1238 B.n754 B.n753 10.6151
R1239 B.n753 B.n752 10.6151
R1240 B.n752 B.n44 10.6151
R1241 B.n746 B.n44 10.6151
R1242 B.n746 B.n745 10.6151
R1243 B.n745 B.n744 10.6151
R1244 B.n109 B.n52 10.6151
R1245 B.n112 B.n109 10.6151
R1246 B.n113 B.n112 10.6151
R1247 B.n116 B.n113 10.6151
R1248 B.n117 B.n116 10.6151
R1249 B.n120 B.n117 10.6151
R1250 B.n121 B.n120 10.6151
R1251 B.n124 B.n121 10.6151
R1252 B.n125 B.n124 10.6151
R1253 B.n128 B.n125 10.6151
R1254 B.n129 B.n128 10.6151
R1255 B.n132 B.n129 10.6151
R1256 B.n133 B.n132 10.6151
R1257 B.n136 B.n133 10.6151
R1258 B.n137 B.n136 10.6151
R1259 B.n140 B.n137 10.6151
R1260 B.n141 B.n140 10.6151
R1261 B.n144 B.n141 10.6151
R1262 B.n145 B.n144 10.6151
R1263 B.n148 B.n145 10.6151
R1264 B.n149 B.n148 10.6151
R1265 B.n152 B.n149 10.6151
R1266 B.n153 B.n152 10.6151
R1267 B.n156 B.n153 10.6151
R1268 B.n157 B.n156 10.6151
R1269 B.n160 B.n157 10.6151
R1270 B.n161 B.n160 10.6151
R1271 B.n164 B.n161 10.6151
R1272 B.n165 B.n164 10.6151
R1273 B.n168 B.n165 10.6151
R1274 B.n169 B.n168 10.6151
R1275 B.n172 B.n169 10.6151
R1276 B.n173 B.n172 10.6151
R1277 B.n176 B.n173 10.6151
R1278 B.n177 B.n176 10.6151
R1279 B.n180 B.n177 10.6151
R1280 B.n181 B.n180 10.6151
R1281 B.n184 B.n181 10.6151
R1282 B.n185 B.n184 10.6151
R1283 B.n188 B.n185 10.6151
R1284 B.n189 B.n188 10.6151
R1285 B.n192 B.n189 10.6151
R1286 B.n193 B.n192 10.6151
R1287 B.n196 B.n193 10.6151
R1288 B.n201 B.n198 10.6151
R1289 B.n202 B.n201 10.6151
R1290 B.n205 B.n202 10.6151
R1291 B.n206 B.n205 10.6151
R1292 B.n209 B.n206 10.6151
R1293 B.n210 B.n209 10.6151
R1294 B.n213 B.n210 10.6151
R1295 B.n214 B.n213 10.6151
R1296 B.n217 B.n214 10.6151
R1297 B.n222 B.n219 10.6151
R1298 B.n223 B.n222 10.6151
R1299 B.n226 B.n223 10.6151
R1300 B.n227 B.n226 10.6151
R1301 B.n230 B.n227 10.6151
R1302 B.n231 B.n230 10.6151
R1303 B.n234 B.n231 10.6151
R1304 B.n235 B.n234 10.6151
R1305 B.n238 B.n235 10.6151
R1306 B.n239 B.n238 10.6151
R1307 B.n242 B.n239 10.6151
R1308 B.n243 B.n242 10.6151
R1309 B.n246 B.n243 10.6151
R1310 B.n247 B.n246 10.6151
R1311 B.n250 B.n247 10.6151
R1312 B.n251 B.n250 10.6151
R1313 B.n254 B.n251 10.6151
R1314 B.n255 B.n254 10.6151
R1315 B.n258 B.n255 10.6151
R1316 B.n259 B.n258 10.6151
R1317 B.n262 B.n259 10.6151
R1318 B.n263 B.n262 10.6151
R1319 B.n266 B.n263 10.6151
R1320 B.n267 B.n266 10.6151
R1321 B.n270 B.n267 10.6151
R1322 B.n271 B.n270 10.6151
R1323 B.n274 B.n271 10.6151
R1324 B.n275 B.n274 10.6151
R1325 B.n278 B.n275 10.6151
R1326 B.n279 B.n278 10.6151
R1327 B.n282 B.n279 10.6151
R1328 B.n283 B.n282 10.6151
R1329 B.n286 B.n283 10.6151
R1330 B.n287 B.n286 10.6151
R1331 B.n290 B.n287 10.6151
R1332 B.n291 B.n290 10.6151
R1333 B.n294 B.n291 10.6151
R1334 B.n295 B.n294 10.6151
R1335 B.n298 B.n295 10.6151
R1336 B.n299 B.n298 10.6151
R1337 B.n302 B.n299 10.6151
R1338 B.n304 B.n302 10.6151
R1339 B.n305 B.n304 10.6151
R1340 B.n738 B.n305 10.6151
R1341 B.n393 B.n392 9.36635
R1342 B.n524 B.n523 9.36635
R1343 B.n197 B.n196 9.36635
R1344 B.n219 B.n218 9.36635
R1345 B.n802 B.n0 8.11757
R1346 B.n802 B.n1 8.11757
R1347 B.n324 B.t3 7.13756
R1348 B.t4 B.n781 7.13756
R1349 B.n505 B.n392 1.24928
R1350 B.n523 B.n522 1.24928
R1351 B.n198 B.n197 1.24928
R1352 B.n218 B.n217 1.24928
R1353 B.n658 B.t0 1.19001
R1354 B.t1 B.n772 1.19001
R1355 VN.n3 VN.t5 259.7
R1356 VN.n13 VN.t4 259.7
R1357 VN.n2 VN.t1 224.369
R1358 VN.n8 VN.t0 224.369
R1359 VN.n12 VN.t2 224.369
R1360 VN.n18 VN.t3 224.369
R1361 VN.n9 VN.n8 173.472
R1362 VN.n19 VN.n18 173.472
R1363 VN.n17 VN.n10 161.3
R1364 VN.n16 VN.n15 161.3
R1365 VN.n14 VN.n11 161.3
R1366 VN.n7 VN.n0 161.3
R1367 VN.n6 VN.n5 161.3
R1368 VN.n4 VN.n1 161.3
R1369 VN.n6 VN.n1 52.5823
R1370 VN.n16 VN.n11 52.5823
R1371 VN VN.n19 45.2941
R1372 VN.n3 VN.n2 41.7378
R1373 VN.n13 VN.n12 41.7378
R1374 VN.n7 VN.n6 28.2389
R1375 VN.n17 VN.n16 28.2389
R1376 VN.n2 VN.n1 24.3439
R1377 VN.n12 VN.n11 24.3439
R1378 VN.n14 VN.n13 17.5582
R1379 VN.n4 VN.n3 17.5582
R1380 VN.n8 VN.n7 12.1722
R1381 VN.n18 VN.n17 12.1722
R1382 VN.n19 VN.n10 0.189894
R1383 VN.n15 VN.n10 0.189894
R1384 VN.n15 VN.n14 0.189894
R1385 VN.n5 VN.n4 0.189894
R1386 VN.n5 VN.n0 0.189894
R1387 VN.n9 VN.n0 0.189894
R1388 VN VN.n9 0.0516364
R1389 VTAIL.n7 VTAIL.t8 46.8321
R1390 VTAIL.n11 VTAIL.t10 46.8319
R1391 VTAIL.n2 VTAIL.t2 46.8319
R1392 VTAIL.n10 VTAIL.t1 46.8319
R1393 VTAIL.n9 VTAIL.n8 45.3344
R1394 VTAIL.n6 VTAIL.n5 45.3344
R1395 VTAIL.n1 VTAIL.n0 45.3343
R1396 VTAIL.n4 VTAIL.n3 45.3343
R1397 VTAIL.n6 VTAIL.n4 26.7807
R1398 VTAIL.n11 VTAIL.n10 25.2721
R1399 VTAIL.n7 VTAIL.n6 1.50912
R1400 VTAIL.n10 VTAIL.n9 1.50912
R1401 VTAIL.n4 VTAIL.n2 1.50912
R1402 VTAIL.n0 VTAIL.t9 1.49823
R1403 VTAIL.n0 VTAIL.t6 1.49823
R1404 VTAIL.n3 VTAIL.t0 1.49823
R1405 VTAIL.n3 VTAIL.t4 1.49823
R1406 VTAIL.n8 VTAIL.t3 1.49823
R1407 VTAIL.n8 VTAIL.t5 1.49823
R1408 VTAIL.n5 VTAIL.t7 1.49823
R1409 VTAIL.n5 VTAIL.t11 1.49823
R1410 VTAIL.n9 VTAIL.n7 1.22464
R1411 VTAIL.n2 VTAIL.n1 1.22464
R1412 VTAIL VTAIL.n11 1.07378
R1413 VTAIL VTAIL.n1 0.435845
R1414 VDD2.n1 VDD2.t0 64.5868
R1415 VDD2.n2 VDD2.t2 63.5109
R1416 VDD2.n1 VDD2.n0 62.3349
R1417 VDD2 VDD2.n3 62.332
R1418 VDD2.n2 VDD2.n1 40.0149
R1419 VDD2.n3 VDD2.t3 1.49823
R1420 VDD2.n3 VDD2.t1 1.49823
R1421 VDD2.n0 VDD2.t4 1.49823
R1422 VDD2.n0 VDD2.t5 1.49823
R1423 VDD2 VDD2.n2 1.19016
R1424 VP.n7 VP.t3 259.7
R1425 VP.n20 VP.t5 224.369
R1426 VP.n14 VP.t4 224.369
R1427 VP.n26 VP.t0 224.369
R1428 VP.n6 VP.t2 224.369
R1429 VP.n12 VP.t1 224.369
R1430 VP.n15 VP.n14 173.472
R1431 VP.n27 VP.n26 173.472
R1432 VP.n13 VP.n12 173.472
R1433 VP.n8 VP.n5 161.3
R1434 VP.n10 VP.n9 161.3
R1435 VP.n11 VP.n4 161.3
R1436 VP.n25 VP.n0 161.3
R1437 VP.n24 VP.n23 161.3
R1438 VP.n22 VP.n1 161.3
R1439 VP.n21 VP.n20 161.3
R1440 VP.n19 VP.n2 161.3
R1441 VP.n18 VP.n17 161.3
R1442 VP.n16 VP.n3 161.3
R1443 VP.n19 VP.n18 52.5823
R1444 VP.n24 VP.n1 52.5823
R1445 VP.n10 VP.n5 52.5823
R1446 VP.n15 VP.n13 44.9134
R1447 VP.n7 VP.n6 41.7378
R1448 VP.n18 VP.n3 28.2389
R1449 VP.n25 VP.n24 28.2389
R1450 VP.n11 VP.n10 28.2389
R1451 VP.n20 VP.n19 24.3439
R1452 VP.n20 VP.n1 24.3439
R1453 VP.n6 VP.n5 24.3439
R1454 VP.n8 VP.n7 17.5582
R1455 VP.n14 VP.n3 12.1722
R1456 VP.n26 VP.n25 12.1722
R1457 VP.n12 VP.n11 12.1722
R1458 VP.n9 VP.n8 0.189894
R1459 VP.n9 VP.n4 0.189894
R1460 VP.n13 VP.n4 0.189894
R1461 VP.n16 VP.n15 0.189894
R1462 VP.n17 VP.n16 0.189894
R1463 VP.n17 VP.n2 0.189894
R1464 VP.n21 VP.n2 0.189894
R1465 VP.n22 VP.n21 0.189894
R1466 VP.n23 VP.n22 0.189894
R1467 VP.n23 VP.n0 0.189894
R1468 VP.n27 VP.n0 0.189894
R1469 VP VP.n27 0.0516364
R1470 VDD1 VDD1.t2 64.7006
R1471 VDD1.n1 VDD1.t1 64.5868
R1472 VDD1.n1 VDD1.n0 62.3349
R1473 VDD1.n3 VDD1.n2 62.013
R1474 VDD1.n3 VDD1.n1 41.3522
R1475 VDD1.n2 VDD1.t3 1.49823
R1476 VDD1.n2 VDD1.t4 1.49823
R1477 VDD1.n0 VDD1.t0 1.49823
R1478 VDD1.n0 VDD1.t5 1.49823
R1479 VDD1 VDD1.n3 0.319466
C0 VDD2 VTAIL 8.68705f
C1 VTAIL VP 6.18038f
C2 VDD2 VP 0.358214f
C3 VN VTAIL 6.16592f
C4 VDD1 VTAIL 8.64645f
C5 VDD2 VDD1 0.97716f
C6 VN VDD2 6.328681f
C7 VN VP 6.00907f
C8 VDD1 VP 6.53404f
C9 VN VDD1 0.148779f
C10 VDD2 B 5.27185f
C11 VDD1 B 5.536317f
C12 VTAIL B 7.443413f
C13 VN B 9.683001f
C14 VP B 8.016622f
C15 VDD1.t2 B 2.60807f
C16 VDD1.t1 B 2.60737f
C17 VDD1.t0 B 0.227517f
C18 VDD1.t5 B 0.227517f
C19 VDD1.n0 B 2.04049f
C20 VDD1.n1 B 2.23997f
C21 VDD1.t3 B 0.227517f
C22 VDD1.t4 B 0.227517f
C23 VDD1.n2 B 2.03883f
C24 VDD1.n3 B 2.22437f
C25 VP.n0 B 0.03364f
C26 VP.t0 B 1.72512f
C27 VP.n1 B 0.060337f
C28 VP.n2 B 0.03364f
C29 VP.t5 B 1.72512f
C30 VP.n3 B 0.051059f
C31 VP.n4 B 0.03364f
C32 VP.t1 B 1.72512f
C33 VP.n5 B 0.060337f
C34 VP.t3 B 1.82686f
C35 VP.t2 B 1.72512f
C36 VP.n6 B 0.698421f
C37 VP.n7 B 0.691978f
C38 VP.n8 B 0.212047f
C39 VP.n9 B 0.03364f
C40 VP.n10 B 0.034702f
C41 VP.n11 B 0.051059f
C42 VP.n12 B 0.68945f
C43 VP.n13 B 1.55419f
C44 VP.t4 B 1.72512f
C45 VP.n14 B 0.68945f
C46 VP.n15 B 1.58104f
C47 VP.n16 B 0.03364f
C48 VP.n17 B 0.03364f
C49 VP.n18 B 0.034702f
C50 VP.n19 B 0.060337f
C51 VP.n20 B 0.652926f
C52 VP.n21 B 0.03364f
C53 VP.n22 B 0.03364f
C54 VP.n23 B 0.03364f
C55 VP.n24 B 0.034702f
C56 VP.n25 B 0.051059f
C57 VP.n26 B 0.68945f
C58 VP.n27 B 0.031233f
C59 VDD2.t0 B 2.60398f
C60 VDD2.t4 B 0.227221f
C61 VDD2.t5 B 0.227221f
C62 VDD2.n0 B 2.03783f
C63 VDD2.n1 B 2.15448f
C64 VDD2.t2 B 2.5986f
C65 VDD2.n2 B 2.23626f
C66 VDD2.t3 B 0.227221f
C67 VDD2.t1 B 0.227221f
C68 VDD2.n3 B 2.0378f
C69 VTAIL.t9 B 0.241023f
C70 VTAIL.t6 B 0.241023f
C71 VTAIL.n0 B 2.09077f
C72 VTAIL.n1 B 0.353321f
C73 VTAIL.t2 B 2.66792f
C74 VTAIL.n2 B 0.513297f
C75 VTAIL.t0 B 0.241023f
C76 VTAIL.t4 B 0.241023f
C77 VTAIL.n3 B 2.09077f
C78 VTAIL.n4 B 1.72704f
C79 VTAIL.t7 B 0.241023f
C80 VTAIL.t11 B 0.241023f
C81 VTAIL.n5 B 2.09077f
C82 VTAIL.n6 B 1.72705f
C83 VTAIL.t8 B 2.66793f
C84 VTAIL.n7 B 0.513291f
C85 VTAIL.t3 B 0.241023f
C86 VTAIL.t5 B 0.241023f
C87 VTAIL.n8 B 2.09077f
C88 VTAIL.n9 B 0.433111f
C89 VTAIL.t1 B 2.66792f
C90 VTAIL.n10 B 1.69508f
C91 VTAIL.t10 B 2.66792f
C92 VTAIL.n11 B 1.66271f
C93 VN.n0 B 0.033196f
C94 VN.t0 B 1.70237f
C95 VN.n1 B 0.059541f
C96 VN.t5 B 1.80277f
C97 VN.t1 B 1.70237f
C98 VN.n2 B 0.689208f
C99 VN.n3 B 0.68285f
C100 VN.n4 B 0.20925f
C101 VN.n5 B 0.033196f
C102 VN.n6 B 0.034244f
C103 VN.n7 B 0.050386f
C104 VN.n8 B 0.680356f
C105 VN.n9 B 0.030821f
C106 VN.n10 B 0.033196f
C107 VN.t3 B 1.70237f
C108 VN.n11 B 0.059541f
C109 VN.t4 B 1.80277f
C110 VN.t2 B 1.70237f
C111 VN.n12 B 0.689208f
C112 VN.n13 B 0.68285f
C113 VN.n14 B 0.20925f
C114 VN.n15 B 0.033196f
C115 VN.n16 B 0.034244f
C116 VN.n17 B 0.050386f
C117 VN.n18 B 0.680356f
C118 VN.n19 B 1.5554f
.ends

