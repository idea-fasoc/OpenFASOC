* NGSPICE file created from tg_sample_0001.ext - technology: sky130A

.subckt tg_sample_0001 VIN VGN VGP VSS VCC VOUT
X0 VCC.t7 VCC.t4 VCC.t6 VCC.t5 sky130_fd_pr__pfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X1 VSS.t7 VSS.t4 VSS.t6 VSS.t5 sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
X2 VCC.t3 VCC.t0 VCC.t2 VCC.t1 sky130_fd_pr__pfet_01v8 ad=0.95 pd=4.95 as=0 ps=0 w=2 l=0.15
X3 VOUT.t1 VGN.t0 VIN.t1 VSS.t8 sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0.475 ps=2.95 w=1 l=0.15
X4 VOUT.t0 VGP.t0 VIN.t0 VCC.t8 sky130_fd_pr__pfet_01v8 ad=0.95 pd=4.95 as=0.95 ps=4.95 w=2 l=0.15
X5 VSS.t3 VSS.t0 VSS.t2 VSS.t1 sky130_fd_pr__nfet_01v8 ad=0.475 pd=2.95 as=0 ps=0 w=1 l=0.15
R0 VCC.n98 VCC.t0 577.768
R1 VCC.n42 VCC.t4 577.768
R2 VCC.n128 VCC.n9 362.928
R3 VCC.n126 VCC.n13 362.928
R4 VCC.n65 VCC.n32 362.928
R5 VCC.n62 VCC.n30 362.928
R6 VCC.n98 VCC.t2 223.349
R7 VCC.n42 VCC.t7 223.349
R8 VCC.n99 VCC.t3 210.743
R9 VCC.n43 VCC.t6 210.743
R10 VCC.n126 VCC.n125 185
R11 VCC.n127 VCC.n126 185
R12 VCC.n14 VCC.n12 185
R13 VCC.n12 VCC.n10 185
R14 VCC.n91 VCC.n90 185
R15 VCC.n90 VCC.n89 185
R16 VCC.n17 VCC.n16 185
R17 VCC.n88 VCC.n17 185
R18 VCC.n86 VCC.n85 185
R19 VCC.n87 VCC.n86 185
R20 VCC.n19 VCC.n18 185
R21 VCC.n24 VCC.n18 185
R22 VCC.n81 VCC.n80 185
R23 VCC.n80 VCC.n79 185
R24 VCC.n22 VCC.n21 185
R25 VCC.n23 VCC.n22 185
R26 VCC.n70 VCC.n69 185
R27 VCC.n71 VCC.n70 185
R28 VCC.n33 VCC.n32 185
R29 VCC.n32 VCC.n31 185
R30 VCC.n30 VCC.n29 185
R31 VCC.n31 VCC.n30 185
R32 VCC.n73 VCC.n72 185
R33 VCC.n72 VCC.n71 185
R34 VCC.n27 VCC.n25 185
R35 VCC.n25 VCC.n23 185
R36 VCC.n78 VCC.n77 185
R37 VCC.n79 VCC.n78 185
R38 VCC.n26 VCC.n2 185
R39 VCC.n26 VCC.n24 185
R40 VCC.n135 VCC.n3 185
R41 VCC.n87 VCC.n3 185
R42 VCC.n134 VCC.n4 185
R43 VCC.n88 VCC.n4 185
R44 VCC.n133 VCC.n5 185
R45 VCC.n89 VCC.n5 185
R46 VCC.n8 VCC.n6 185
R47 VCC.n10 VCC.n8 185
R48 VCC.n129 VCC.n128 185
R49 VCC.n128 VCC.n127 185
R50 VCC.n123 VCC.n13 185
R51 VCC.n122 VCC.n121 185
R52 VCC.n119 VCC.n94 185
R53 VCC.n117 VCC.n116 185
R54 VCC.n115 VCC.n95 185
R55 VCC.n114 VCC.n113 185
R56 VCC.n111 VCC.n96 185
R57 VCC.n109 VCC.n108 185
R58 VCC.n107 VCC.n97 185
R59 VCC.n106 VCC.n105 185
R60 VCC.n103 VCC.n102 185
R61 VCC.n9 VCC.n7 185
R62 VCC.n62 VCC.n61 185
R63 VCC.n60 VCC.n41 185
R64 VCC.n58 VCC.n40 185
R65 VCC.n64 VCC.n40 185
R66 VCC.n57 VCC.n56 185
R67 VCC.n55 VCC.n54 185
R68 VCC.n53 VCC.n52 185
R69 VCC.n51 VCC.n50 185
R70 VCC.n49 VCC.n48 185
R71 VCC.n47 VCC.n46 185
R72 VCC.n45 VCC.n44 185
R73 VCC.n35 VCC.n34 185
R74 VCC.n66 VCC.n65 185
R75 VCC.n65 VCC.n64 185
R76 VCC.n70 VCC.n32 146.341
R77 VCC.n70 VCC.n22 146.341
R78 VCC.n80 VCC.n22 146.341
R79 VCC.n80 VCC.n18 146.341
R80 VCC.n86 VCC.n18 146.341
R81 VCC.n86 VCC.n17 146.341
R82 VCC.n90 VCC.n17 146.341
R83 VCC.n90 VCC.n12 146.341
R84 VCC.n126 VCC.n12 146.341
R85 VCC.n72 VCC.n30 146.341
R86 VCC.n72 VCC.n25 146.341
R87 VCC.n78 VCC.n25 146.341
R88 VCC.n78 VCC.n26 146.341
R89 VCC.n26 VCC.n3 146.341
R90 VCC.n4 VCC.n3 146.341
R91 VCC.n5 VCC.n4 146.341
R92 VCC.n8 VCC.n5 146.341
R93 VCC.n128 VCC.n8 146.341
R94 VCC.n64 VCC.n31 120.499
R95 VCC.n127 VCC.n11 120.499
R96 VCC.n105 VCC.n103 99.5127
R97 VCC.n109 VCC.n97 99.5127
R98 VCC.n113 VCC.n111 99.5127
R99 VCC.n117 VCC.n95 99.5127
R100 VCC.n121 VCC.n119 99.5127
R101 VCC.n41 VCC.n40 99.5127
R102 VCC.n56 VCC.n40 99.5127
R103 VCC.n54 VCC.n53 99.5127
R104 VCC.n50 VCC.n49 99.5127
R105 VCC.n46 VCC.n45 99.5127
R106 VCC.n65 VCC.n35 99.5127
R107 VCC.n71 VCC.n31 77.7419
R108 VCC.n79 VCC.n23 77.7419
R109 VCC.n79 VCC.n24 77.7419
R110 VCC.n88 VCC.n87 77.7419
R111 VCC.n89 VCC.n88 77.7419
R112 VCC.n127 VCC.n10 77.7419
R113 VCC.t5 VCC.n23 76.1871
R114 VCC.n89 VCC.t1 76.1871
R115 VCC.n120 VCC.n11 72.8958
R116 VCC.n118 VCC.n11 72.8958
R117 VCC.n112 VCC.n11 72.8958
R118 VCC.n110 VCC.n11 72.8958
R119 VCC.n104 VCC.n11 72.8958
R120 VCC.n101 VCC.n11 72.8958
R121 VCC.n64 VCC.n63 72.8958
R122 VCC.n64 VCC.n36 72.8958
R123 VCC.n64 VCC.n37 72.8958
R124 VCC.n64 VCC.n38 72.8958
R125 VCC.n64 VCC.n39 72.8958
R126 VCC.n103 VCC.n101 39.2114
R127 VCC.n104 VCC.n97 39.2114
R128 VCC.n111 VCC.n110 39.2114
R129 VCC.n112 VCC.n95 39.2114
R130 VCC.n119 VCC.n118 39.2114
R131 VCC.n120 VCC.n13 39.2114
R132 VCC.n63 VCC.n62 39.2114
R133 VCC.n56 VCC.n36 39.2114
R134 VCC.n53 VCC.n37 39.2114
R135 VCC.n49 VCC.n38 39.2114
R136 VCC.n45 VCC.n39 39.2114
R137 VCC.n121 VCC.n120 39.2114
R138 VCC.n118 VCC.n117 39.2114
R139 VCC.n113 VCC.n112 39.2114
R140 VCC.n110 VCC.n109 39.2114
R141 VCC.n105 VCC.n104 39.2114
R142 VCC.n101 VCC.n9 39.2114
R143 VCC.n63 VCC.n41 39.2114
R144 VCC.n54 VCC.n36 39.2114
R145 VCC.n50 VCC.n37 39.2114
R146 VCC.n46 VCC.n38 39.2114
R147 VCC.n39 VCC.n35 39.2114
R148 VCC.n24 VCC.t8 38.8712
R149 VCC.n87 VCC.t8 38.8712
R150 VCC.n130 VCC.n7 30.4539
R151 VCC.n124 VCC.n123 30.4539
R152 VCC.n61 VCC.n28 30.4539
R153 VCC.n67 VCC.n66 30.4539
R154 VCC.n100 VCC.n99 29.2853
R155 VCC.n59 VCC.n43 29.2853
R156 VCC.n69 VCC.n33 19.3944
R157 VCC.n69 VCC.n21 19.3944
R158 VCC.n81 VCC.n21 19.3944
R159 VCC.n81 VCC.n19 19.3944
R160 VCC.n85 VCC.n19 19.3944
R161 VCC.n85 VCC.n16 19.3944
R162 VCC.n91 VCC.n16 19.3944
R163 VCC.n91 VCC.n14 19.3944
R164 VCC.n125 VCC.n14 19.3944
R165 VCC.n73 VCC.n29 19.3944
R166 VCC.n73 VCC.n27 19.3944
R167 VCC.n77 VCC.n27 19.3944
R168 VCC.n77 VCC.n2 19.3944
R169 VCC.n135 VCC.n2 19.3944
R170 VCC.n135 VCC.n134 19.3944
R171 VCC.n134 VCC.n133 19.3944
R172 VCC.n133 VCC.n6 19.3944
R173 VCC.n129 VCC.n6 19.3944
R174 VCC.n99 VCC.n98 12.6066
R175 VCC.n43 VCC.n42 12.6066
R176 VCC.n102 VCC.n7 10.6151
R177 VCC.n107 VCC.n106 10.6151
R178 VCC.n108 VCC.n107 10.6151
R179 VCC.n108 VCC.n96 10.6151
R180 VCC.n114 VCC.n96 10.6151
R181 VCC.n115 VCC.n114 10.6151
R182 VCC.n116 VCC.n115 10.6151
R183 VCC.n116 VCC.n94 10.6151
R184 VCC.n122 VCC.n94 10.6151
R185 VCC.n123 VCC.n122 10.6151
R186 VCC.n61 VCC.n60 10.6151
R187 VCC.n58 VCC.n57 10.6151
R188 VCC.n57 VCC.n55 10.6151
R189 VCC.n55 VCC.n52 10.6151
R190 VCC.n52 VCC.n51 10.6151
R191 VCC.n51 VCC.n48 10.6151
R192 VCC.n48 VCC.n47 10.6151
R193 VCC.n47 VCC.n44 10.6151
R194 VCC.n44 VCC.n34 10.6151
R195 VCC.n66 VCC.n34 10.6151
R196 VCC.n134 VCC.n0 9.3005
R197 VCC.n133 VCC.n132 9.3005
R198 VCC.n131 VCC.n6 9.3005
R199 VCC.n130 VCC.n129 9.3005
R200 VCC.n69 VCC.n68 9.3005
R201 VCC.n21 VCC.n20 9.3005
R202 VCC.n82 VCC.n81 9.3005
R203 VCC.n83 VCC.n19 9.3005
R204 VCC.n85 VCC.n84 9.3005
R205 VCC.n16 VCC.n15 9.3005
R206 VCC.n92 VCC.n91 9.3005
R207 VCC.n93 VCC.n14 9.3005
R208 VCC.n125 VCC.n124 9.3005
R209 VCC.n67 VCC.n33 9.3005
R210 VCC.n29 VCC.n28 9.3005
R211 VCC.n74 VCC.n73 9.3005
R212 VCC.n75 VCC.n27 9.3005
R213 VCC.n77 VCC.n76 9.3005
R214 VCC.n2 VCC.n1 9.3005
R215 VCC VCC.n135 9.3005
R216 VCC.n102 VCC.n100 5.77611
R217 VCC.n60 VCC.n59 5.77611
R218 VCC.n106 VCC.n100 4.83952
R219 VCC.n59 VCC.n58 4.83952
R220 VCC.n71 VCC.t5 1.55533
R221 VCC.t1 VCC.n10 1.55533
R222 VCC VCC.n0 0.152939
R223 VCC.n132 VCC.n0 0.152939
R224 VCC.n132 VCC.n131 0.152939
R225 VCC.n131 VCC.n130 0.152939
R226 VCC.n68 VCC.n67 0.152939
R227 VCC.n68 VCC.n20 0.152939
R228 VCC.n82 VCC.n20 0.152939
R229 VCC.n83 VCC.n82 0.152939
R230 VCC.n84 VCC.n83 0.152939
R231 VCC.n84 VCC.n15 0.152939
R232 VCC.n92 VCC.n15 0.152939
R233 VCC.n93 VCC.n92 0.152939
R234 VCC.n124 VCC.n93 0.152939
R235 VCC.n74 VCC.n28 0.152939
R236 VCC.n75 VCC.n74 0.152939
R237 VCC.n76 VCC.n75 0.152939
R238 VCC.n76 VCC.n1 0.152939
R239 VCC VCC.n1 0.1255
R240 VSS.n56 VSS.n29 712.345
R241 VSS.n117 VSS.n11 712.345
R242 VSS.n58 VSS.n30 643.855
R243 VSS.n37 VSS.n28 643.855
R244 VSS.n116 VSS.n13 643.855
R245 VSS.n118 VSS.n9 643.855
R246 VSS.n31 VSS.n30 585
R247 VSS.n30 VSS.n29 585
R248 VSS.n63 VSS.n62 585
R249 VSS.n64 VSS.n63 585
R250 VSS.n22 VSS.n21 585
R251 VSS.n23 VSS.n22 585
R252 VSS.n76 VSS.n75 585
R253 VSS.n75 VSS.n74 585
R254 VSS.n19 VSS.n18 585
R255 VSS.n73 VSS.n18 585
R256 VSS.n81 VSS.n80 585
R257 VSS.n82 VSS.n81 585
R258 VSS.n17 VSS.n16 585
R259 VSS.n83 VSS.n17 585
R260 VSS.n86 VSS.n85 585
R261 VSS.n85 VSS.n84 585
R262 VSS.n14 VSS.n12 585
R263 VSS.n12 VSS.n10 585
R264 VSS.n116 VSS.n115 585
R265 VSS.n117 VSS.n116 585
R266 VSS.n119 VSS.n118 585
R267 VSS.n118 VSS.n117 585
R268 VSS.n8 VSS.n6 585
R269 VSS.n10 VSS.n8 585
R270 VSS.n123 VSS.n5 585
R271 VSS.n84 VSS.n5 585
R272 VSS.n124 VSS.n4 585
R273 VSS.n83 VSS.n4 585
R274 VSS.n125 VSS.n3 585
R275 VSS.n82 VSS.n3 585
R276 VSS.n72 VSS.n2 585
R277 VSS.n73 VSS.n72 585
R278 VSS.n71 VSS.n70 585
R279 VSS.n74 VSS.n71 585
R280 VSS.n25 VSS.n24 585
R281 VSS.n24 VSS.n23 585
R282 VSS.n66 VSS.n65 585
R283 VSS.n65 VSS.n64 585
R284 VSS.n28 VSS.n27 585
R285 VSS.n29 VSS.n28 585
R286 VSS.n9 VSS.n7 585
R287 VSS.n99 VSS.n95 585
R288 VSS.n101 VSS.n100 585
R289 VSS.n103 VSS.n92 585
R290 VSS.n105 VSS.n104 585
R291 VSS.n106 VSS.n91 585
R292 VSS.n108 VSS.n107 585
R293 VSS.n110 VSS.n89 585
R294 VSS.n112 VSS.n111 585
R295 VSS.n113 VSS.n13 585
R296 VSS.n59 VSS.n58 585
R297 VSS.n33 VSS.n32 585
R298 VSS.n55 VSS.n54 585
R299 VSS.n56 VSS.n55 585
R300 VSS.n53 VSS.n38 585
R301 VSS.n52 VSS.n51 585
R302 VSS.n50 VSS.n49 585
R303 VSS.n48 VSS.n47 585
R304 VSS.n46 VSS.n45 585
R305 VSS.n44 VSS.n43 585
R306 VSS.n42 VSS.n37 585
R307 VSS.n56 VSS.n37 585
R308 VSS.n96 VSS.t4 417.101
R309 VSS.n39 VSS.t0 417.101
R310 VSS.n64 VSS.n29 393.56
R311 VSS.n74 VSS.n23 393.56
R312 VSS.n74 VSS.n73 393.56
R313 VSS.n83 VSS.n82 393.56
R314 VSS.n84 VSS.n83 393.56
R315 VSS.n117 VSS.n10 393.56
R316 VSS.t1 VSS.n23 385.69
R317 VSS.n84 VSS.t5 385.69
R318 VSS.n96 VSS.t6 256.697
R319 VSS.n39 VSS.t3 256.697
R320 VSS.n94 VSS.n11 256.663
R321 VSS.n102 VSS.n11 256.663
R322 VSS.n93 VSS.n11 256.663
R323 VSS.n109 VSS.n11 256.663
R324 VSS.n90 VSS.n11 256.663
R325 VSS.n57 VSS.n56 256.663
R326 VSS.n56 VSS.n34 256.663
R327 VSS.n56 VSS.n35 256.663
R328 VSS.n56 VSS.n36 256.663
R329 VSS.n97 VSS.t7 244.091
R330 VSS.n40 VSS.t2 244.091
R331 VSS.n63 VSS.n30 240.244
R332 VSS.n63 VSS.n22 240.244
R333 VSS.n75 VSS.n22 240.244
R334 VSS.n75 VSS.n18 240.244
R335 VSS.n81 VSS.n18 240.244
R336 VSS.n81 VSS.n17 240.244
R337 VSS.n85 VSS.n17 240.244
R338 VSS.n85 VSS.n12 240.244
R339 VSS.n116 VSS.n12 240.244
R340 VSS.n65 VSS.n28 240.244
R341 VSS.n65 VSS.n24 240.244
R342 VSS.n71 VSS.n24 240.244
R343 VSS.n72 VSS.n71 240.244
R344 VSS.n72 VSS.n3 240.244
R345 VSS.n4 VSS.n3 240.244
R346 VSS.n5 VSS.n4 240.244
R347 VSS.n8 VSS.n5 240.244
R348 VSS.n118 VSS.n8 240.244
R349 VSS.n73 VSS.t8 196.78
R350 VSS.n82 VSS.t8 196.78
R351 VSS.n55 VSS.n33 163.367
R352 VSS.n55 VSS.n38 163.367
R353 VSS.n51 VSS.n50 163.367
R354 VSS.n47 VSS.n46 163.367
R355 VSS.n43 VSS.n37 163.367
R356 VSS.n111 VSS.n110 163.367
R357 VSS.n108 VSS.n91 163.367
R358 VSS.n104 VSS.n103 163.367
R359 VSS.n101 VSS.n95 163.367
R360 VSS.n58 VSS.n57 71.676
R361 VSS.n38 VSS.n34 71.676
R362 VSS.n50 VSS.n35 71.676
R363 VSS.n46 VSS.n36 71.676
R364 VSS.n111 VSS.n90 71.676
R365 VSS.n109 VSS.n108 71.676
R366 VSS.n104 VSS.n93 71.676
R367 VSS.n102 VSS.n101 71.676
R368 VSS.n94 VSS.n9 71.676
R369 VSS.n95 VSS.n94 71.676
R370 VSS.n103 VSS.n102 71.676
R371 VSS.n93 VSS.n91 71.676
R372 VSS.n110 VSS.n109 71.676
R373 VSS.n90 VSS.n13 71.676
R374 VSS.n57 VSS.n33 71.676
R375 VSS.n51 VSS.n34 71.676
R376 VSS.n47 VSS.n35 71.676
R377 VSS.n43 VSS.n36 71.676
R378 VSS.n98 VSS.n97 34.3278
R379 VSS.n41 VSS.n40 34.3278
R380 VSS.n114 VSS.n113 29.5569
R381 VSS.n120 VSS.n7 29.5569
R382 VSS.n60 VSS.n59 29.5569
R383 VSS.n42 VSS.n26 29.5569
R384 VSS.n62 VSS.n31 19.3944
R385 VSS.n62 VSS.n21 19.3944
R386 VSS.n76 VSS.n21 19.3944
R387 VSS.n76 VSS.n19 19.3944
R388 VSS.n80 VSS.n19 19.3944
R389 VSS.n80 VSS.n16 19.3944
R390 VSS.n86 VSS.n16 19.3944
R391 VSS.n86 VSS.n14 19.3944
R392 VSS.n115 VSS.n14 19.3944
R393 VSS.n66 VSS.n27 19.3944
R394 VSS.n66 VSS.n25 19.3944
R395 VSS.n70 VSS.n25 19.3944
R396 VSS.n70 VSS.n2 19.3944
R397 VSS.n125 VSS.n2 19.3944
R398 VSS.n125 VSS.n124 19.3944
R399 VSS.n124 VSS.n123 19.3944
R400 VSS.n123 VSS.n6 19.3944
R401 VSS.n119 VSS.n6 19.3944
R402 VSS.n97 VSS.n96 12.6066
R403 VSS.n40 VSS.n39 12.6066
R404 VSS.n113 VSS.n112 10.6151
R405 VSS.n112 VSS.n89 10.6151
R406 VSS.n107 VSS.n89 10.6151
R407 VSS.n107 VSS.n106 10.6151
R408 VSS.n106 VSS.n105 10.6151
R409 VSS.n105 VSS.n92 10.6151
R410 VSS.n100 VSS.n99 10.6151
R411 VSS.n99 VSS.n7 10.6151
R412 VSS.n59 VSS.n32 10.6151
R413 VSS.n54 VSS.n32 10.6151
R414 VSS.n54 VSS.n53 10.6151
R415 VSS.n53 VSS.n52 10.6151
R416 VSS.n52 VSS.n49 10.6151
R417 VSS.n49 VSS.n48 10.6151
R418 VSS.n45 VSS.n44 10.6151
R419 VSS.n44 VSS.n42 10.6151
R420 VSS.n98 VSS.n92 10.459
R421 VSS.n48 VSS.n41 10.459
R422 VSS.n124 VSS.n0 9.3005
R423 VSS.n123 VSS.n122 9.3005
R424 VSS.n121 VSS.n6 9.3005
R425 VSS.n120 VSS.n119 9.3005
R426 VSS.n60 VSS.n31 9.3005
R427 VSS.n62 VSS.n61 9.3005
R428 VSS.n21 VSS.n20 9.3005
R429 VSS.n77 VSS.n76 9.3005
R430 VSS.n78 VSS.n19 9.3005
R431 VSS.n80 VSS.n79 9.3005
R432 VSS.n16 VSS.n15 9.3005
R433 VSS.n87 VSS.n86 9.3005
R434 VSS.n88 VSS.n14 9.3005
R435 VSS.n115 VSS.n114 9.3005
R436 VSS.n67 VSS.n66 9.3005
R437 VSS.n68 VSS.n25 9.3005
R438 VSS.n70 VSS.n69 9.3005
R439 VSS.n2 VSS.n1 9.3005
R440 VSS.n27 VSS.n26 9.3005
R441 VSS VSS.n125 9.3005
R442 VSS.n64 VSS.t1 7.8717
R443 VSS.t5 VSS.n10 7.8717
R444 VSS.n100 VSS.n98 0.156598
R445 VSS.n45 VSS.n41 0.156598
R446 VSS VSS.n0 0.152939
R447 VSS.n122 VSS.n0 0.152939
R448 VSS.n122 VSS.n121 0.152939
R449 VSS.n121 VSS.n120 0.152939
R450 VSS.n61 VSS.n60 0.152939
R451 VSS.n61 VSS.n20 0.152939
R452 VSS.n77 VSS.n20 0.152939
R453 VSS.n78 VSS.n77 0.152939
R454 VSS.n79 VSS.n78 0.152939
R455 VSS.n79 VSS.n15 0.152939
R456 VSS.n87 VSS.n15 0.152939
R457 VSS.n88 VSS.n87 0.152939
R458 VSS.n114 VSS.n88 0.152939
R459 VSS.n67 VSS.n26 0.152939
R460 VSS.n68 VSS.n67 0.152939
R461 VSS.n69 VSS.n68 0.152939
R462 VSS.n69 VSS.n1 0.152939
R463 VSS VSS.n1 0.1255
R464 VGN VGN.t0 554.946
R465 VIN VIN.t1 253.738
R466 VIN VIN.t0 220.423
R467 VOUT VOUT.t1 281.171
R468 VOUT VOUT.t0 225.857
R469 VGP VGP.t0 715.611
C0 VIN VOUT 0.900701f
C1 VGN VGP 6e-19
C2 VGN VCC 9.03e-19
C3 VOUT VGP 0.039324f
C4 VOUT VCC 0.590075f
C5 VIN VGP 0.045268f
C6 VIN VCC 0.482153f
C7 VGN VOUT 0.025611f
C8 VGN VIN 0.033741f
C9 VCC VGP 0.300445f
C10 VGN VSS 0.32606f
C11 VOUT VSS 0.67486f
C12 VIN VSS 0.63023f
C13 VGP VSS 0.035537f
C14 VCC VSS 6.31784f
.ends

