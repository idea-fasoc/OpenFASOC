* NGSPICE file created from diff_pair_sample_0602.ext - technology: sky130A

.subckt diff_pair_sample_0602 VTAIL VN VP B VDD2 VDD1
X0 B.t17 B.t15 B.t16 B.t12 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=0 ps=0 w=18.99 l=3.36
X1 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=0 ps=0 w=18.99 l=3.36
X2 VTAIL.t7 VN.t0 VDD2.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=3.13335 ps=19.32 w=18.99 l=3.36
X3 B.t10 B.t8 B.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=0 ps=0 w=18.99 l=3.36
X4 VTAIL.t1 VP.t0 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=3.13335 ps=19.32 w=18.99 l=3.36
X5 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=0 ps=0 w=18.99 l=3.36
X6 VDD2.t0 VN.t1 VTAIL.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=3.13335 pd=19.32 as=7.4061 ps=38.76 w=18.99 l=3.36
X7 VDD2.t3 VN.t2 VTAIL.t5 B.t0 sky130_fd_pr__nfet_01v8 ad=3.13335 pd=19.32 as=7.4061 ps=38.76 w=18.99 l=3.36
X8 VTAIL.t4 VN.t3 VDD2.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=3.13335 ps=19.32 w=18.99 l=3.36
X9 VDD1.t2 VP.t1 VTAIL.t2 B.t3 sky130_fd_pr__nfet_01v8 ad=3.13335 pd=19.32 as=7.4061 ps=38.76 w=18.99 l=3.36
X10 VTAIL.t0 VP.t2 VDD1.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=7.4061 pd=38.76 as=3.13335 ps=19.32 w=18.99 l=3.36
X11 VDD1.t0 VP.t3 VTAIL.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=3.13335 pd=19.32 as=7.4061 ps=38.76 w=18.99 l=3.36
R0 B.n1005 B.n1004 585
R1 B.n412 B.n143 585
R2 B.n411 B.n410 585
R3 B.n409 B.n408 585
R4 B.n407 B.n406 585
R5 B.n405 B.n404 585
R6 B.n403 B.n402 585
R7 B.n401 B.n400 585
R8 B.n399 B.n398 585
R9 B.n397 B.n396 585
R10 B.n395 B.n394 585
R11 B.n393 B.n392 585
R12 B.n391 B.n390 585
R13 B.n389 B.n388 585
R14 B.n387 B.n386 585
R15 B.n385 B.n384 585
R16 B.n383 B.n382 585
R17 B.n381 B.n380 585
R18 B.n379 B.n378 585
R19 B.n377 B.n376 585
R20 B.n375 B.n374 585
R21 B.n373 B.n372 585
R22 B.n371 B.n370 585
R23 B.n369 B.n368 585
R24 B.n367 B.n366 585
R25 B.n365 B.n364 585
R26 B.n363 B.n362 585
R27 B.n361 B.n360 585
R28 B.n359 B.n358 585
R29 B.n357 B.n356 585
R30 B.n355 B.n354 585
R31 B.n353 B.n352 585
R32 B.n351 B.n350 585
R33 B.n349 B.n348 585
R34 B.n347 B.n346 585
R35 B.n345 B.n344 585
R36 B.n343 B.n342 585
R37 B.n341 B.n340 585
R38 B.n339 B.n338 585
R39 B.n337 B.n336 585
R40 B.n335 B.n334 585
R41 B.n333 B.n332 585
R42 B.n331 B.n330 585
R43 B.n329 B.n328 585
R44 B.n327 B.n326 585
R45 B.n325 B.n324 585
R46 B.n323 B.n322 585
R47 B.n321 B.n320 585
R48 B.n319 B.n318 585
R49 B.n317 B.n316 585
R50 B.n315 B.n314 585
R51 B.n313 B.n312 585
R52 B.n311 B.n310 585
R53 B.n309 B.n308 585
R54 B.n307 B.n306 585
R55 B.n305 B.n304 585
R56 B.n303 B.n302 585
R57 B.n301 B.n300 585
R58 B.n299 B.n298 585
R59 B.n297 B.n296 585
R60 B.n295 B.n294 585
R61 B.n293 B.n292 585
R62 B.n291 B.n290 585
R63 B.n289 B.n288 585
R64 B.n287 B.n286 585
R65 B.n285 B.n284 585
R66 B.n283 B.n282 585
R67 B.n281 B.n280 585
R68 B.n279 B.n278 585
R69 B.n277 B.n276 585
R70 B.n275 B.n274 585
R71 B.n273 B.n272 585
R72 B.n271 B.n270 585
R73 B.n269 B.n268 585
R74 B.n267 B.n266 585
R75 B.n265 B.n264 585
R76 B.n263 B.n262 585
R77 B.n261 B.n260 585
R78 B.n259 B.n258 585
R79 B.n257 B.n256 585
R80 B.n255 B.n254 585
R81 B.n253 B.n252 585
R82 B.n251 B.n250 585
R83 B.n249 B.n248 585
R84 B.n247 B.n246 585
R85 B.n245 B.n244 585
R86 B.n243 B.n242 585
R87 B.n241 B.n240 585
R88 B.n239 B.n238 585
R89 B.n237 B.n236 585
R90 B.n235 B.n234 585
R91 B.n233 B.n232 585
R92 B.n231 B.n230 585
R93 B.n229 B.n228 585
R94 B.n227 B.n226 585
R95 B.n225 B.n224 585
R96 B.n223 B.n222 585
R97 B.n221 B.n220 585
R98 B.n219 B.n218 585
R99 B.n217 B.n216 585
R100 B.n215 B.n214 585
R101 B.n213 B.n212 585
R102 B.n211 B.n210 585
R103 B.n209 B.n208 585
R104 B.n207 B.n206 585
R105 B.n205 B.n204 585
R106 B.n203 B.n202 585
R107 B.n201 B.n200 585
R108 B.n199 B.n198 585
R109 B.n197 B.n196 585
R110 B.n195 B.n194 585
R111 B.n193 B.n192 585
R112 B.n191 B.n190 585
R113 B.n189 B.n188 585
R114 B.n187 B.n186 585
R115 B.n185 B.n184 585
R116 B.n183 B.n182 585
R117 B.n181 B.n180 585
R118 B.n179 B.n178 585
R119 B.n177 B.n176 585
R120 B.n175 B.n174 585
R121 B.n173 B.n172 585
R122 B.n171 B.n170 585
R123 B.n169 B.n168 585
R124 B.n167 B.n166 585
R125 B.n165 B.n164 585
R126 B.n163 B.n162 585
R127 B.n161 B.n160 585
R128 B.n159 B.n158 585
R129 B.n157 B.n156 585
R130 B.n155 B.n154 585
R131 B.n153 B.n152 585
R132 B.n151 B.n150 585
R133 B.n75 B.n74 585
R134 B.n1003 B.n76 585
R135 B.n1008 B.n76 585
R136 B.n1002 B.n1001 585
R137 B.n1001 B.n72 585
R138 B.n1000 B.n71 585
R139 B.n1014 B.n71 585
R140 B.n999 B.n70 585
R141 B.n1015 B.n70 585
R142 B.n998 B.n69 585
R143 B.n1016 B.n69 585
R144 B.n997 B.n996 585
R145 B.n996 B.n65 585
R146 B.n995 B.n64 585
R147 B.n1022 B.n64 585
R148 B.n994 B.n63 585
R149 B.n1023 B.n63 585
R150 B.n993 B.n62 585
R151 B.n1024 B.n62 585
R152 B.n992 B.n991 585
R153 B.n991 B.n58 585
R154 B.n990 B.n57 585
R155 B.n1030 B.n57 585
R156 B.n989 B.n56 585
R157 B.n1031 B.n56 585
R158 B.n988 B.n55 585
R159 B.n1032 B.n55 585
R160 B.n987 B.n986 585
R161 B.n986 B.n51 585
R162 B.n985 B.n50 585
R163 B.n1038 B.n50 585
R164 B.n984 B.n49 585
R165 B.n1039 B.n49 585
R166 B.n983 B.n48 585
R167 B.n1040 B.n48 585
R168 B.n982 B.n981 585
R169 B.n981 B.n44 585
R170 B.n980 B.n43 585
R171 B.n1046 B.n43 585
R172 B.n979 B.n42 585
R173 B.n1047 B.n42 585
R174 B.n978 B.n41 585
R175 B.n1048 B.n41 585
R176 B.n977 B.n976 585
R177 B.n976 B.n37 585
R178 B.n975 B.n36 585
R179 B.n1054 B.n36 585
R180 B.n974 B.n35 585
R181 B.n1055 B.n35 585
R182 B.n973 B.n34 585
R183 B.n1056 B.n34 585
R184 B.n972 B.n971 585
R185 B.n971 B.n30 585
R186 B.n970 B.n29 585
R187 B.n1062 B.n29 585
R188 B.n969 B.n28 585
R189 B.n1063 B.n28 585
R190 B.n968 B.n27 585
R191 B.n1064 B.n27 585
R192 B.n967 B.n966 585
R193 B.n966 B.n23 585
R194 B.n965 B.n22 585
R195 B.n1070 B.n22 585
R196 B.n964 B.n21 585
R197 B.n1071 B.n21 585
R198 B.n963 B.n20 585
R199 B.n1072 B.n20 585
R200 B.n962 B.n961 585
R201 B.n961 B.n19 585
R202 B.n960 B.n15 585
R203 B.n1078 B.n15 585
R204 B.n959 B.n14 585
R205 B.n1079 B.n14 585
R206 B.n958 B.n13 585
R207 B.n1080 B.n13 585
R208 B.n957 B.n956 585
R209 B.n956 B.n12 585
R210 B.n955 B.n954 585
R211 B.n955 B.n8 585
R212 B.n953 B.n7 585
R213 B.n1087 B.n7 585
R214 B.n952 B.n6 585
R215 B.n1088 B.n6 585
R216 B.n951 B.n5 585
R217 B.n1089 B.n5 585
R218 B.n950 B.n949 585
R219 B.n949 B.n4 585
R220 B.n948 B.n413 585
R221 B.n948 B.n947 585
R222 B.n938 B.n414 585
R223 B.n415 B.n414 585
R224 B.n940 B.n939 585
R225 B.n941 B.n940 585
R226 B.n937 B.n420 585
R227 B.n420 B.n419 585
R228 B.n936 B.n935 585
R229 B.n935 B.n934 585
R230 B.n422 B.n421 585
R231 B.n927 B.n422 585
R232 B.n926 B.n925 585
R233 B.n928 B.n926 585
R234 B.n924 B.n427 585
R235 B.n427 B.n426 585
R236 B.n923 B.n922 585
R237 B.n922 B.n921 585
R238 B.n429 B.n428 585
R239 B.n430 B.n429 585
R240 B.n914 B.n913 585
R241 B.n915 B.n914 585
R242 B.n912 B.n435 585
R243 B.n435 B.n434 585
R244 B.n911 B.n910 585
R245 B.n910 B.n909 585
R246 B.n437 B.n436 585
R247 B.n438 B.n437 585
R248 B.n902 B.n901 585
R249 B.n903 B.n902 585
R250 B.n900 B.n443 585
R251 B.n443 B.n442 585
R252 B.n899 B.n898 585
R253 B.n898 B.n897 585
R254 B.n445 B.n444 585
R255 B.n446 B.n445 585
R256 B.n890 B.n889 585
R257 B.n891 B.n890 585
R258 B.n888 B.n451 585
R259 B.n451 B.n450 585
R260 B.n887 B.n886 585
R261 B.n886 B.n885 585
R262 B.n453 B.n452 585
R263 B.n454 B.n453 585
R264 B.n878 B.n877 585
R265 B.n879 B.n878 585
R266 B.n876 B.n459 585
R267 B.n459 B.n458 585
R268 B.n875 B.n874 585
R269 B.n874 B.n873 585
R270 B.n461 B.n460 585
R271 B.n462 B.n461 585
R272 B.n866 B.n865 585
R273 B.n867 B.n866 585
R274 B.n864 B.n467 585
R275 B.n467 B.n466 585
R276 B.n863 B.n862 585
R277 B.n862 B.n861 585
R278 B.n469 B.n468 585
R279 B.n470 B.n469 585
R280 B.n854 B.n853 585
R281 B.n855 B.n854 585
R282 B.n852 B.n475 585
R283 B.n475 B.n474 585
R284 B.n851 B.n850 585
R285 B.n850 B.n849 585
R286 B.n477 B.n476 585
R287 B.n478 B.n477 585
R288 B.n842 B.n841 585
R289 B.n843 B.n842 585
R290 B.n840 B.n483 585
R291 B.n483 B.n482 585
R292 B.n839 B.n838 585
R293 B.n838 B.n837 585
R294 B.n485 B.n484 585
R295 B.n486 B.n485 585
R296 B.n830 B.n829 585
R297 B.n831 B.n830 585
R298 B.n489 B.n488 585
R299 B.n562 B.n560 585
R300 B.n563 B.n559 585
R301 B.n563 B.n490 585
R302 B.n566 B.n565 585
R303 B.n567 B.n558 585
R304 B.n569 B.n568 585
R305 B.n571 B.n557 585
R306 B.n574 B.n573 585
R307 B.n575 B.n556 585
R308 B.n577 B.n576 585
R309 B.n579 B.n555 585
R310 B.n582 B.n581 585
R311 B.n583 B.n554 585
R312 B.n585 B.n584 585
R313 B.n587 B.n553 585
R314 B.n590 B.n589 585
R315 B.n591 B.n552 585
R316 B.n593 B.n592 585
R317 B.n595 B.n551 585
R318 B.n598 B.n597 585
R319 B.n599 B.n550 585
R320 B.n601 B.n600 585
R321 B.n603 B.n549 585
R322 B.n606 B.n605 585
R323 B.n607 B.n548 585
R324 B.n609 B.n608 585
R325 B.n611 B.n547 585
R326 B.n614 B.n613 585
R327 B.n615 B.n546 585
R328 B.n617 B.n616 585
R329 B.n619 B.n545 585
R330 B.n622 B.n621 585
R331 B.n623 B.n544 585
R332 B.n625 B.n624 585
R333 B.n627 B.n543 585
R334 B.n630 B.n629 585
R335 B.n631 B.n542 585
R336 B.n633 B.n632 585
R337 B.n635 B.n541 585
R338 B.n638 B.n637 585
R339 B.n639 B.n540 585
R340 B.n641 B.n640 585
R341 B.n643 B.n539 585
R342 B.n646 B.n645 585
R343 B.n647 B.n538 585
R344 B.n649 B.n648 585
R345 B.n651 B.n537 585
R346 B.n654 B.n653 585
R347 B.n655 B.n536 585
R348 B.n657 B.n656 585
R349 B.n659 B.n535 585
R350 B.n662 B.n661 585
R351 B.n663 B.n534 585
R352 B.n665 B.n664 585
R353 B.n667 B.n533 585
R354 B.n670 B.n669 585
R355 B.n671 B.n532 585
R356 B.n673 B.n672 585
R357 B.n675 B.n531 585
R358 B.n678 B.n677 585
R359 B.n679 B.n530 585
R360 B.n684 B.n683 585
R361 B.n686 B.n529 585
R362 B.n689 B.n688 585
R363 B.n690 B.n528 585
R364 B.n692 B.n691 585
R365 B.n694 B.n527 585
R366 B.n697 B.n696 585
R367 B.n698 B.n526 585
R368 B.n700 B.n699 585
R369 B.n702 B.n525 585
R370 B.n705 B.n704 585
R371 B.n707 B.n522 585
R372 B.n709 B.n708 585
R373 B.n711 B.n521 585
R374 B.n714 B.n713 585
R375 B.n715 B.n520 585
R376 B.n717 B.n716 585
R377 B.n719 B.n519 585
R378 B.n722 B.n721 585
R379 B.n723 B.n518 585
R380 B.n725 B.n724 585
R381 B.n727 B.n517 585
R382 B.n730 B.n729 585
R383 B.n731 B.n516 585
R384 B.n733 B.n732 585
R385 B.n735 B.n515 585
R386 B.n738 B.n737 585
R387 B.n739 B.n514 585
R388 B.n741 B.n740 585
R389 B.n743 B.n513 585
R390 B.n746 B.n745 585
R391 B.n747 B.n512 585
R392 B.n749 B.n748 585
R393 B.n751 B.n511 585
R394 B.n754 B.n753 585
R395 B.n755 B.n510 585
R396 B.n757 B.n756 585
R397 B.n759 B.n509 585
R398 B.n762 B.n761 585
R399 B.n763 B.n508 585
R400 B.n765 B.n764 585
R401 B.n767 B.n507 585
R402 B.n770 B.n769 585
R403 B.n771 B.n506 585
R404 B.n773 B.n772 585
R405 B.n775 B.n505 585
R406 B.n778 B.n777 585
R407 B.n779 B.n504 585
R408 B.n781 B.n780 585
R409 B.n783 B.n503 585
R410 B.n786 B.n785 585
R411 B.n787 B.n502 585
R412 B.n789 B.n788 585
R413 B.n791 B.n501 585
R414 B.n794 B.n793 585
R415 B.n795 B.n500 585
R416 B.n797 B.n796 585
R417 B.n799 B.n499 585
R418 B.n802 B.n801 585
R419 B.n803 B.n498 585
R420 B.n805 B.n804 585
R421 B.n807 B.n497 585
R422 B.n810 B.n809 585
R423 B.n811 B.n496 585
R424 B.n813 B.n812 585
R425 B.n815 B.n495 585
R426 B.n818 B.n817 585
R427 B.n819 B.n494 585
R428 B.n821 B.n820 585
R429 B.n823 B.n493 585
R430 B.n824 B.n492 585
R431 B.n827 B.n826 585
R432 B.n828 B.n491 585
R433 B.n491 B.n490 585
R434 B.n833 B.n832 585
R435 B.n832 B.n831 585
R436 B.n834 B.n487 585
R437 B.n487 B.n486 585
R438 B.n836 B.n835 585
R439 B.n837 B.n836 585
R440 B.n481 B.n480 585
R441 B.n482 B.n481 585
R442 B.n845 B.n844 585
R443 B.n844 B.n843 585
R444 B.n846 B.n479 585
R445 B.n479 B.n478 585
R446 B.n848 B.n847 585
R447 B.n849 B.n848 585
R448 B.n473 B.n472 585
R449 B.n474 B.n473 585
R450 B.n857 B.n856 585
R451 B.n856 B.n855 585
R452 B.n858 B.n471 585
R453 B.n471 B.n470 585
R454 B.n860 B.n859 585
R455 B.n861 B.n860 585
R456 B.n465 B.n464 585
R457 B.n466 B.n465 585
R458 B.n869 B.n868 585
R459 B.n868 B.n867 585
R460 B.n870 B.n463 585
R461 B.n463 B.n462 585
R462 B.n872 B.n871 585
R463 B.n873 B.n872 585
R464 B.n457 B.n456 585
R465 B.n458 B.n457 585
R466 B.n881 B.n880 585
R467 B.n880 B.n879 585
R468 B.n882 B.n455 585
R469 B.n455 B.n454 585
R470 B.n884 B.n883 585
R471 B.n885 B.n884 585
R472 B.n449 B.n448 585
R473 B.n450 B.n449 585
R474 B.n893 B.n892 585
R475 B.n892 B.n891 585
R476 B.n894 B.n447 585
R477 B.n447 B.n446 585
R478 B.n896 B.n895 585
R479 B.n897 B.n896 585
R480 B.n441 B.n440 585
R481 B.n442 B.n441 585
R482 B.n905 B.n904 585
R483 B.n904 B.n903 585
R484 B.n906 B.n439 585
R485 B.n439 B.n438 585
R486 B.n908 B.n907 585
R487 B.n909 B.n908 585
R488 B.n433 B.n432 585
R489 B.n434 B.n433 585
R490 B.n917 B.n916 585
R491 B.n916 B.n915 585
R492 B.n918 B.n431 585
R493 B.n431 B.n430 585
R494 B.n920 B.n919 585
R495 B.n921 B.n920 585
R496 B.n425 B.n424 585
R497 B.n426 B.n425 585
R498 B.n930 B.n929 585
R499 B.n929 B.n928 585
R500 B.n931 B.n423 585
R501 B.n927 B.n423 585
R502 B.n933 B.n932 585
R503 B.n934 B.n933 585
R504 B.n418 B.n417 585
R505 B.n419 B.n418 585
R506 B.n943 B.n942 585
R507 B.n942 B.n941 585
R508 B.n944 B.n416 585
R509 B.n416 B.n415 585
R510 B.n946 B.n945 585
R511 B.n947 B.n946 585
R512 B.n3 B.n0 585
R513 B.n4 B.n3 585
R514 B.n1086 B.n1 585
R515 B.n1087 B.n1086 585
R516 B.n1085 B.n1084 585
R517 B.n1085 B.n8 585
R518 B.n1083 B.n9 585
R519 B.n12 B.n9 585
R520 B.n1082 B.n1081 585
R521 B.n1081 B.n1080 585
R522 B.n11 B.n10 585
R523 B.n1079 B.n11 585
R524 B.n1077 B.n1076 585
R525 B.n1078 B.n1077 585
R526 B.n1075 B.n16 585
R527 B.n19 B.n16 585
R528 B.n1074 B.n1073 585
R529 B.n1073 B.n1072 585
R530 B.n18 B.n17 585
R531 B.n1071 B.n18 585
R532 B.n1069 B.n1068 585
R533 B.n1070 B.n1069 585
R534 B.n1067 B.n24 585
R535 B.n24 B.n23 585
R536 B.n1066 B.n1065 585
R537 B.n1065 B.n1064 585
R538 B.n26 B.n25 585
R539 B.n1063 B.n26 585
R540 B.n1061 B.n1060 585
R541 B.n1062 B.n1061 585
R542 B.n1059 B.n31 585
R543 B.n31 B.n30 585
R544 B.n1058 B.n1057 585
R545 B.n1057 B.n1056 585
R546 B.n33 B.n32 585
R547 B.n1055 B.n33 585
R548 B.n1053 B.n1052 585
R549 B.n1054 B.n1053 585
R550 B.n1051 B.n38 585
R551 B.n38 B.n37 585
R552 B.n1050 B.n1049 585
R553 B.n1049 B.n1048 585
R554 B.n40 B.n39 585
R555 B.n1047 B.n40 585
R556 B.n1045 B.n1044 585
R557 B.n1046 B.n1045 585
R558 B.n1043 B.n45 585
R559 B.n45 B.n44 585
R560 B.n1042 B.n1041 585
R561 B.n1041 B.n1040 585
R562 B.n47 B.n46 585
R563 B.n1039 B.n47 585
R564 B.n1037 B.n1036 585
R565 B.n1038 B.n1037 585
R566 B.n1035 B.n52 585
R567 B.n52 B.n51 585
R568 B.n1034 B.n1033 585
R569 B.n1033 B.n1032 585
R570 B.n54 B.n53 585
R571 B.n1031 B.n54 585
R572 B.n1029 B.n1028 585
R573 B.n1030 B.n1029 585
R574 B.n1027 B.n59 585
R575 B.n59 B.n58 585
R576 B.n1026 B.n1025 585
R577 B.n1025 B.n1024 585
R578 B.n61 B.n60 585
R579 B.n1023 B.n61 585
R580 B.n1021 B.n1020 585
R581 B.n1022 B.n1021 585
R582 B.n1019 B.n66 585
R583 B.n66 B.n65 585
R584 B.n1018 B.n1017 585
R585 B.n1017 B.n1016 585
R586 B.n68 B.n67 585
R587 B.n1015 B.n68 585
R588 B.n1013 B.n1012 585
R589 B.n1014 B.n1013 585
R590 B.n1011 B.n73 585
R591 B.n73 B.n72 585
R592 B.n1010 B.n1009 585
R593 B.n1009 B.n1008 585
R594 B.n1090 B.n1089 585
R595 B.n1088 B.n2 585
R596 B.n1009 B.n75 521.33
R597 B.n1005 B.n76 521.33
R598 B.n830 B.n491 521.33
R599 B.n832 B.n489 521.33
R600 B.n147 B.t16 474.38
R601 B.n144 B.t13 474.38
R602 B.n523 B.t10 474.38
R603 B.n680 B.t7 474.38
R604 B.n145 B.t14 402.817
R605 B.n524 B.t9 402.817
R606 B.n148 B.t17 402.817
R607 B.n681 B.t6 402.817
R608 B.n147 B.t15 345.171
R609 B.n144 B.t11 345.171
R610 B.n523 B.t8 345.171
R611 B.n680 B.t4 345.171
R612 B.n1007 B.n1006 256.663
R613 B.n1007 B.n142 256.663
R614 B.n1007 B.n141 256.663
R615 B.n1007 B.n140 256.663
R616 B.n1007 B.n139 256.663
R617 B.n1007 B.n138 256.663
R618 B.n1007 B.n137 256.663
R619 B.n1007 B.n136 256.663
R620 B.n1007 B.n135 256.663
R621 B.n1007 B.n134 256.663
R622 B.n1007 B.n133 256.663
R623 B.n1007 B.n132 256.663
R624 B.n1007 B.n131 256.663
R625 B.n1007 B.n130 256.663
R626 B.n1007 B.n129 256.663
R627 B.n1007 B.n128 256.663
R628 B.n1007 B.n127 256.663
R629 B.n1007 B.n126 256.663
R630 B.n1007 B.n125 256.663
R631 B.n1007 B.n124 256.663
R632 B.n1007 B.n123 256.663
R633 B.n1007 B.n122 256.663
R634 B.n1007 B.n121 256.663
R635 B.n1007 B.n120 256.663
R636 B.n1007 B.n119 256.663
R637 B.n1007 B.n118 256.663
R638 B.n1007 B.n117 256.663
R639 B.n1007 B.n116 256.663
R640 B.n1007 B.n115 256.663
R641 B.n1007 B.n114 256.663
R642 B.n1007 B.n113 256.663
R643 B.n1007 B.n112 256.663
R644 B.n1007 B.n111 256.663
R645 B.n1007 B.n110 256.663
R646 B.n1007 B.n109 256.663
R647 B.n1007 B.n108 256.663
R648 B.n1007 B.n107 256.663
R649 B.n1007 B.n106 256.663
R650 B.n1007 B.n105 256.663
R651 B.n1007 B.n104 256.663
R652 B.n1007 B.n103 256.663
R653 B.n1007 B.n102 256.663
R654 B.n1007 B.n101 256.663
R655 B.n1007 B.n100 256.663
R656 B.n1007 B.n99 256.663
R657 B.n1007 B.n98 256.663
R658 B.n1007 B.n97 256.663
R659 B.n1007 B.n96 256.663
R660 B.n1007 B.n95 256.663
R661 B.n1007 B.n94 256.663
R662 B.n1007 B.n93 256.663
R663 B.n1007 B.n92 256.663
R664 B.n1007 B.n91 256.663
R665 B.n1007 B.n90 256.663
R666 B.n1007 B.n89 256.663
R667 B.n1007 B.n88 256.663
R668 B.n1007 B.n87 256.663
R669 B.n1007 B.n86 256.663
R670 B.n1007 B.n85 256.663
R671 B.n1007 B.n84 256.663
R672 B.n1007 B.n83 256.663
R673 B.n1007 B.n82 256.663
R674 B.n1007 B.n81 256.663
R675 B.n1007 B.n80 256.663
R676 B.n1007 B.n79 256.663
R677 B.n1007 B.n78 256.663
R678 B.n1007 B.n77 256.663
R679 B.n561 B.n490 256.663
R680 B.n564 B.n490 256.663
R681 B.n570 B.n490 256.663
R682 B.n572 B.n490 256.663
R683 B.n578 B.n490 256.663
R684 B.n580 B.n490 256.663
R685 B.n586 B.n490 256.663
R686 B.n588 B.n490 256.663
R687 B.n594 B.n490 256.663
R688 B.n596 B.n490 256.663
R689 B.n602 B.n490 256.663
R690 B.n604 B.n490 256.663
R691 B.n610 B.n490 256.663
R692 B.n612 B.n490 256.663
R693 B.n618 B.n490 256.663
R694 B.n620 B.n490 256.663
R695 B.n626 B.n490 256.663
R696 B.n628 B.n490 256.663
R697 B.n634 B.n490 256.663
R698 B.n636 B.n490 256.663
R699 B.n642 B.n490 256.663
R700 B.n644 B.n490 256.663
R701 B.n650 B.n490 256.663
R702 B.n652 B.n490 256.663
R703 B.n658 B.n490 256.663
R704 B.n660 B.n490 256.663
R705 B.n666 B.n490 256.663
R706 B.n668 B.n490 256.663
R707 B.n674 B.n490 256.663
R708 B.n676 B.n490 256.663
R709 B.n685 B.n490 256.663
R710 B.n687 B.n490 256.663
R711 B.n693 B.n490 256.663
R712 B.n695 B.n490 256.663
R713 B.n701 B.n490 256.663
R714 B.n703 B.n490 256.663
R715 B.n710 B.n490 256.663
R716 B.n712 B.n490 256.663
R717 B.n718 B.n490 256.663
R718 B.n720 B.n490 256.663
R719 B.n726 B.n490 256.663
R720 B.n728 B.n490 256.663
R721 B.n734 B.n490 256.663
R722 B.n736 B.n490 256.663
R723 B.n742 B.n490 256.663
R724 B.n744 B.n490 256.663
R725 B.n750 B.n490 256.663
R726 B.n752 B.n490 256.663
R727 B.n758 B.n490 256.663
R728 B.n760 B.n490 256.663
R729 B.n766 B.n490 256.663
R730 B.n768 B.n490 256.663
R731 B.n774 B.n490 256.663
R732 B.n776 B.n490 256.663
R733 B.n782 B.n490 256.663
R734 B.n784 B.n490 256.663
R735 B.n790 B.n490 256.663
R736 B.n792 B.n490 256.663
R737 B.n798 B.n490 256.663
R738 B.n800 B.n490 256.663
R739 B.n806 B.n490 256.663
R740 B.n808 B.n490 256.663
R741 B.n814 B.n490 256.663
R742 B.n816 B.n490 256.663
R743 B.n822 B.n490 256.663
R744 B.n825 B.n490 256.663
R745 B.n1092 B.n1091 256.663
R746 B.n152 B.n151 163.367
R747 B.n156 B.n155 163.367
R748 B.n160 B.n159 163.367
R749 B.n164 B.n163 163.367
R750 B.n168 B.n167 163.367
R751 B.n172 B.n171 163.367
R752 B.n176 B.n175 163.367
R753 B.n180 B.n179 163.367
R754 B.n184 B.n183 163.367
R755 B.n188 B.n187 163.367
R756 B.n192 B.n191 163.367
R757 B.n196 B.n195 163.367
R758 B.n200 B.n199 163.367
R759 B.n204 B.n203 163.367
R760 B.n208 B.n207 163.367
R761 B.n212 B.n211 163.367
R762 B.n216 B.n215 163.367
R763 B.n220 B.n219 163.367
R764 B.n224 B.n223 163.367
R765 B.n228 B.n227 163.367
R766 B.n232 B.n231 163.367
R767 B.n236 B.n235 163.367
R768 B.n240 B.n239 163.367
R769 B.n244 B.n243 163.367
R770 B.n248 B.n247 163.367
R771 B.n252 B.n251 163.367
R772 B.n256 B.n255 163.367
R773 B.n260 B.n259 163.367
R774 B.n264 B.n263 163.367
R775 B.n268 B.n267 163.367
R776 B.n272 B.n271 163.367
R777 B.n276 B.n275 163.367
R778 B.n280 B.n279 163.367
R779 B.n284 B.n283 163.367
R780 B.n288 B.n287 163.367
R781 B.n292 B.n291 163.367
R782 B.n296 B.n295 163.367
R783 B.n300 B.n299 163.367
R784 B.n304 B.n303 163.367
R785 B.n308 B.n307 163.367
R786 B.n312 B.n311 163.367
R787 B.n316 B.n315 163.367
R788 B.n320 B.n319 163.367
R789 B.n324 B.n323 163.367
R790 B.n328 B.n327 163.367
R791 B.n332 B.n331 163.367
R792 B.n336 B.n335 163.367
R793 B.n340 B.n339 163.367
R794 B.n344 B.n343 163.367
R795 B.n348 B.n347 163.367
R796 B.n352 B.n351 163.367
R797 B.n356 B.n355 163.367
R798 B.n360 B.n359 163.367
R799 B.n364 B.n363 163.367
R800 B.n368 B.n367 163.367
R801 B.n372 B.n371 163.367
R802 B.n376 B.n375 163.367
R803 B.n380 B.n379 163.367
R804 B.n384 B.n383 163.367
R805 B.n388 B.n387 163.367
R806 B.n392 B.n391 163.367
R807 B.n396 B.n395 163.367
R808 B.n400 B.n399 163.367
R809 B.n404 B.n403 163.367
R810 B.n408 B.n407 163.367
R811 B.n410 B.n143 163.367
R812 B.n830 B.n485 163.367
R813 B.n838 B.n485 163.367
R814 B.n838 B.n483 163.367
R815 B.n842 B.n483 163.367
R816 B.n842 B.n477 163.367
R817 B.n850 B.n477 163.367
R818 B.n850 B.n475 163.367
R819 B.n854 B.n475 163.367
R820 B.n854 B.n469 163.367
R821 B.n862 B.n469 163.367
R822 B.n862 B.n467 163.367
R823 B.n866 B.n467 163.367
R824 B.n866 B.n461 163.367
R825 B.n874 B.n461 163.367
R826 B.n874 B.n459 163.367
R827 B.n878 B.n459 163.367
R828 B.n878 B.n453 163.367
R829 B.n886 B.n453 163.367
R830 B.n886 B.n451 163.367
R831 B.n890 B.n451 163.367
R832 B.n890 B.n445 163.367
R833 B.n898 B.n445 163.367
R834 B.n898 B.n443 163.367
R835 B.n902 B.n443 163.367
R836 B.n902 B.n437 163.367
R837 B.n910 B.n437 163.367
R838 B.n910 B.n435 163.367
R839 B.n914 B.n435 163.367
R840 B.n914 B.n429 163.367
R841 B.n922 B.n429 163.367
R842 B.n922 B.n427 163.367
R843 B.n926 B.n427 163.367
R844 B.n926 B.n422 163.367
R845 B.n935 B.n422 163.367
R846 B.n935 B.n420 163.367
R847 B.n940 B.n420 163.367
R848 B.n940 B.n414 163.367
R849 B.n948 B.n414 163.367
R850 B.n949 B.n948 163.367
R851 B.n949 B.n5 163.367
R852 B.n6 B.n5 163.367
R853 B.n7 B.n6 163.367
R854 B.n955 B.n7 163.367
R855 B.n956 B.n955 163.367
R856 B.n956 B.n13 163.367
R857 B.n14 B.n13 163.367
R858 B.n15 B.n14 163.367
R859 B.n961 B.n15 163.367
R860 B.n961 B.n20 163.367
R861 B.n21 B.n20 163.367
R862 B.n22 B.n21 163.367
R863 B.n966 B.n22 163.367
R864 B.n966 B.n27 163.367
R865 B.n28 B.n27 163.367
R866 B.n29 B.n28 163.367
R867 B.n971 B.n29 163.367
R868 B.n971 B.n34 163.367
R869 B.n35 B.n34 163.367
R870 B.n36 B.n35 163.367
R871 B.n976 B.n36 163.367
R872 B.n976 B.n41 163.367
R873 B.n42 B.n41 163.367
R874 B.n43 B.n42 163.367
R875 B.n981 B.n43 163.367
R876 B.n981 B.n48 163.367
R877 B.n49 B.n48 163.367
R878 B.n50 B.n49 163.367
R879 B.n986 B.n50 163.367
R880 B.n986 B.n55 163.367
R881 B.n56 B.n55 163.367
R882 B.n57 B.n56 163.367
R883 B.n991 B.n57 163.367
R884 B.n991 B.n62 163.367
R885 B.n63 B.n62 163.367
R886 B.n64 B.n63 163.367
R887 B.n996 B.n64 163.367
R888 B.n996 B.n69 163.367
R889 B.n70 B.n69 163.367
R890 B.n71 B.n70 163.367
R891 B.n1001 B.n71 163.367
R892 B.n1001 B.n76 163.367
R893 B.n563 B.n562 163.367
R894 B.n565 B.n563 163.367
R895 B.n569 B.n558 163.367
R896 B.n573 B.n571 163.367
R897 B.n577 B.n556 163.367
R898 B.n581 B.n579 163.367
R899 B.n585 B.n554 163.367
R900 B.n589 B.n587 163.367
R901 B.n593 B.n552 163.367
R902 B.n597 B.n595 163.367
R903 B.n601 B.n550 163.367
R904 B.n605 B.n603 163.367
R905 B.n609 B.n548 163.367
R906 B.n613 B.n611 163.367
R907 B.n617 B.n546 163.367
R908 B.n621 B.n619 163.367
R909 B.n625 B.n544 163.367
R910 B.n629 B.n627 163.367
R911 B.n633 B.n542 163.367
R912 B.n637 B.n635 163.367
R913 B.n641 B.n540 163.367
R914 B.n645 B.n643 163.367
R915 B.n649 B.n538 163.367
R916 B.n653 B.n651 163.367
R917 B.n657 B.n536 163.367
R918 B.n661 B.n659 163.367
R919 B.n665 B.n534 163.367
R920 B.n669 B.n667 163.367
R921 B.n673 B.n532 163.367
R922 B.n677 B.n675 163.367
R923 B.n684 B.n530 163.367
R924 B.n688 B.n686 163.367
R925 B.n692 B.n528 163.367
R926 B.n696 B.n694 163.367
R927 B.n700 B.n526 163.367
R928 B.n704 B.n702 163.367
R929 B.n709 B.n522 163.367
R930 B.n713 B.n711 163.367
R931 B.n717 B.n520 163.367
R932 B.n721 B.n719 163.367
R933 B.n725 B.n518 163.367
R934 B.n729 B.n727 163.367
R935 B.n733 B.n516 163.367
R936 B.n737 B.n735 163.367
R937 B.n741 B.n514 163.367
R938 B.n745 B.n743 163.367
R939 B.n749 B.n512 163.367
R940 B.n753 B.n751 163.367
R941 B.n757 B.n510 163.367
R942 B.n761 B.n759 163.367
R943 B.n765 B.n508 163.367
R944 B.n769 B.n767 163.367
R945 B.n773 B.n506 163.367
R946 B.n777 B.n775 163.367
R947 B.n781 B.n504 163.367
R948 B.n785 B.n783 163.367
R949 B.n789 B.n502 163.367
R950 B.n793 B.n791 163.367
R951 B.n797 B.n500 163.367
R952 B.n801 B.n799 163.367
R953 B.n805 B.n498 163.367
R954 B.n809 B.n807 163.367
R955 B.n813 B.n496 163.367
R956 B.n817 B.n815 163.367
R957 B.n821 B.n494 163.367
R958 B.n824 B.n823 163.367
R959 B.n826 B.n491 163.367
R960 B.n832 B.n487 163.367
R961 B.n836 B.n487 163.367
R962 B.n836 B.n481 163.367
R963 B.n844 B.n481 163.367
R964 B.n844 B.n479 163.367
R965 B.n848 B.n479 163.367
R966 B.n848 B.n473 163.367
R967 B.n856 B.n473 163.367
R968 B.n856 B.n471 163.367
R969 B.n860 B.n471 163.367
R970 B.n860 B.n465 163.367
R971 B.n868 B.n465 163.367
R972 B.n868 B.n463 163.367
R973 B.n872 B.n463 163.367
R974 B.n872 B.n457 163.367
R975 B.n880 B.n457 163.367
R976 B.n880 B.n455 163.367
R977 B.n884 B.n455 163.367
R978 B.n884 B.n449 163.367
R979 B.n892 B.n449 163.367
R980 B.n892 B.n447 163.367
R981 B.n896 B.n447 163.367
R982 B.n896 B.n441 163.367
R983 B.n904 B.n441 163.367
R984 B.n904 B.n439 163.367
R985 B.n908 B.n439 163.367
R986 B.n908 B.n433 163.367
R987 B.n916 B.n433 163.367
R988 B.n916 B.n431 163.367
R989 B.n920 B.n431 163.367
R990 B.n920 B.n425 163.367
R991 B.n929 B.n425 163.367
R992 B.n929 B.n423 163.367
R993 B.n933 B.n423 163.367
R994 B.n933 B.n418 163.367
R995 B.n942 B.n418 163.367
R996 B.n942 B.n416 163.367
R997 B.n946 B.n416 163.367
R998 B.n946 B.n3 163.367
R999 B.n1090 B.n3 163.367
R1000 B.n1086 B.n2 163.367
R1001 B.n1086 B.n1085 163.367
R1002 B.n1085 B.n9 163.367
R1003 B.n1081 B.n9 163.367
R1004 B.n1081 B.n11 163.367
R1005 B.n1077 B.n11 163.367
R1006 B.n1077 B.n16 163.367
R1007 B.n1073 B.n16 163.367
R1008 B.n1073 B.n18 163.367
R1009 B.n1069 B.n18 163.367
R1010 B.n1069 B.n24 163.367
R1011 B.n1065 B.n24 163.367
R1012 B.n1065 B.n26 163.367
R1013 B.n1061 B.n26 163.367
R1014 B.n1061 B.n31 163.367
R1015 B.n1057 B.n31 163.367
R1016 B.n1057 B.n33 163.367
R1017 B.n1053 B.n33 163.367
R1018 B.n1053 B.n38 163.367
R1019 B.n1049 B.n38 163.367
R1020 B.n1049 B.n40 163.367
R1021 B.n1045 B.n40 163.367
R1022 B.n1045 B.n45 163.367
R1023 B.n1041 B.n45 163.367
R1024 B.n1041 B.n47 163.367
R1025 B.n1037 B.n47 163.367
R1026 B.n1037 B.n52 163.367
R1027 B.n1033 B.n52 163.367
R1028 B.n1033 B.n54 163.367
R1029 B.n1029 B.n54 163.367
R1030 B.n1029 B.n59 163.367
R1031 B.n1025 B.n59 163.367
R1032 B.n1025 B.n61 163.367
R1033 B.n1021 B.n61 163.367
R1034 B.n1021 B.n66 163.367
R1035 B.n1017 B.n66 163.367
R1036 B.n1017 B.n68 163.367
R1037 B.n1013 B.n68 163.367
R1038 B.n1013 B.n73 163.367
R1039 B.n1009 B.n73 163.367
R1040 B.n77 B.n75 71.676
R1041 B.n152 B.n78 71.676
R1042 B.n156 B.n79 71.676
R1043 B.n160 B.n80 71.676
R1044 B.n164 B.n81 71.676
R1045 B.n168 B.n82 71.676
R1046 B.n172 B.n83 71.676
R1047 B.n176 B.n84 71.676
R1048 B.n180 B.n85 71.676
R1049 B.n184 B.n86 71.676
R1050 B.n188 B.n87 71.676
R1051 B.n192 B.n88 71.676
R1052 B.n196 B.n89 71.676
R1053 B.n200 B.n90 71.676
R1054 B.n204 B.n91 71.676
R1055 B.n208 B.n92 71.676
R1056 B.n212 B.n93 71.676
R1057 B.n216 B.n94 71.676
R1058 B.n220 B.n95 71.676
R1059 B.n224 B.n96 71.676
R1060 B.n228 B.n97 71.676
R1061 B.n232 B.n98 71.676
R1062 B.n236 B.n99 71.676
R1063 B.n240 B.n100 71.676
R1064 B.n244 B.n101 71.676
R1065 B.n248 B.n102 71.676
R1066 B.n252 B.n103 71.676
R1067 B.n256 B.n104 71.676
R1068 B.n260 B.n105 71.676
R1069 B.n264 B.n106 71.676
R1070 B.n268 B.n107 71.676
R1071 B.n272 B.n108 71.676
R1072 B.n276 B.n109 71.676
R1073 B.n280 B.n110 71.676
R1074 B.n284 B.n111 71.676
R1075 B.n288 B.n112 71.676
R1076 B.n292 B.n113 71.676
R1077 B.n296 B.n114 71.676
R1078 B.n300 B.n115 71.676
R1079 B.n304 B.n116 71.676
R1080 B.n308 B.n117 71.676
R1081 B.n312 B.n118 71.676
R1082 B.n316 B.n119 71.676
R1083 B.n320 B.n120 71.676
R1084 B.n324 B.n121 71.676
R1085 B.n328 B.n122 71.676
R1086 B.n332 B.n123 71.676
R1087 B.n336 B.n124 71.676
R1088 B.n340 B.n125 71.676
R1089 B.n344 B.n126 71.676
R1090 B.n348 B.n127 71.676
R1091 B.n352 B.n128 71.676
R1092 B.n356 B.n129 71.676
R1093 B.n360 B.n130 71.676
R1094 B.n364 B.n131 71.676
R1095 B.n368 B.n132 71.676
R1096 B.n372 B.n133 71.676
R1097 B.n376 B.n134 71.676
R1098 B.n380 B.n135 71.676
R1099 B.n384 B.n136 71.676
R1100 B.n388 B.n137 71.676
R1101 B.n392 B.n138 71.676
R1102 B.n396 B.n139 71.676
R1103 B.n400 B.n140 71.676
R1104 B.n404 B.n141 71.676
R1105 B.n408 B.n142 71.676
R1106 B.n1006 B.n143 71.676
R1107 B.n1006 B.n1005 71.676
R1108 B.n410 B.n142 71.676
R1109 B.n407 B.n141 71.676
R1110 B.n403 B.n140 71.676
R1111 B.n399 B.n139 71.676
R1112 B.n395 B.n138 71.676
R1113 B.n391 B.n137 71.676
R1114 B.n387 B.n136 71.676
R1115 B.n383 B.n135 71.676
R1116 B.n379 B.n134 71.676
R1117 B.n375 B.n133 71.676
R1118 B.n371 B.n132 71.676
R1119 B.n367 B.n131 71.676
R1120 B.n363 B.n130 71.676
R1121 B.n359 B.n129 71.676
R1122 B.n355 B.n128 71.676
R1123 B.n351 B.n127 71.676
R1124 B.n347 B.n126 71.676
R1125 B.n343 B.n125 71.676
R1126 B.n339 B.n124 71.676
R1127 B.n335 B.n123 71.676
R1128 B.n331 B.n122 71.676
R1129 B.n327 B.n121 71.676
R1130 B.n323 B.n120 71.676
R1131 B.n319 B.n119 71.676
R1132 B.n315 B.n118 71.676
R1133 B.n311 B.n117 71.676
R1134 B.n307 B.n116 71.676
R1135 B.n303 B.n115 71.676
R1136 B.n299 B.n114 71.676
R1137 B.n295 B.n113 71.676
R1138 B.n291 B.n112 71.676
R1139 B.n287 B.n111 71.676
R1140 B.n283 B.n110 71.676
R1141 B.n279 B.n109 71.676
R1142 B.n275 B.n108 71.676
R1143 B.n271 B.n107 71.676
R1144 B.n267 B.n106 71.676
R1145 B.n263 B.n105 71.676
R1146 B.n259 B.n104 71.676
R1147 B.n255 B.n103 71.676
R1148 B.n251 B.n102 71.676
R1149 B.n247 B.n101 71.676
R1150 B.n243 B.n100 71.676
R1151 B.n239 B.n99 71.676
R1152 B.n235 B.n98 71.676
R1153 B.n231 B.n97 71.676
R1154 B.n227 B.n96 71.676
R1155 B.n223 B.n95 71.676
R1156 B.n219 B.n94 71.676
R1157 B.n215 B.n93 71.676
R1158 B.n211 B.n92 71.676
R1159 B.n207 B.n91 71.676
R1160 B.n203 B.n90 71.676
R1161 B.n199 B.n89 71.676
R1162 B.n195 B.n88 71.676
R1163 B.n191 B.n87 71.676
R1164 B.n187 B.n86 71.676
R1165 B.n183 B.n85 71.676
R1166 B.n179 B.n84 71.676
R1167 B.n175 B.n83 71.676
R1168 B.n171 B.n82 71.676
R1169 B.n167 B.n81 71.676
R1170 B.n163 B.n80 71.676
R1171 B.n159 B.n79 71.676
R1172 B.n155 B.n78 71.676
R1173 B.n151 B.n77 71.676
R1174 B.n561 B.n489 71.676
R1175 B.n565 B.n564 71.676
R1176 B.n570 B.n569 71.676
R1177 B.n573 B.n572 71.676
R1178 B.n578 B.n577 71.676
R1179 B.n581 B.n580 71.676
R1180 B.n586 B.n585 71.676
R1181 B.n589 B.n588 71.676
R1182 B.n594 B.n593 71.676
R1183 B.n597 B.n596 71.676
R1184 B.n602 B.n601 71.676
R1185 B.n605 B.n604 71.676
R1186 B.n610 B.n609 71.676
R1187 B.n613 B.n612 71.676
R1188 B.n618 B.n617 71.676
R1189 B.n621 B.n620 71.676
R1190 B.n626 B.n625 71.676
R1191 B.n629 B.n628 71.676
R1192 B.n634 B.n633 71.676
R1193 B.n637 B.n636 71.676
R1194 B.n642 B.n641 71.676
R1195 B.n645 B.n644 71.676
R1196 B.n650 B.n649 71.676
R1197 B.n653 B.n652 71.676
R1198 B.n658 B.n657 71.676
R1199 B.n661 B.n660 71.676
R1200 B.n666 B.n665 71.676
R1201 B.n669 B.n668 71.676
R1202 B.n674 B.n673 71.676
R1203 B.n677 B.n676 71.676
R1204 B.n685 B.n684 71.676
R1205 B.n688 B.n687 71.676
R1206 B.n693 B.n692 71.676
R1207 B.n696 B.n695 71.676
R1208 B.n701 B.n700 71.676
R1209 B.n704 B.n703 71.676
R1210 B.n710 B.n709 71.676
R1211 B.n713 B.n712 71.676
R1212 B.n718 B.n717 71.676
R1213 B.n721 B.n720 71.676
R1214 B.n726 B.n725 71.676
R1215 B.n729 B.n728 71.676
R1216 B.n734 B.n733 71.676
R1217 B.n737 B.n736 71.676
R1218 B.n742 B.n741 71.676
R1219 B.n745 B.n744 71.676
R1220 B.n750 B.n749 71.676
R1221 B.n753 B.n752 71.676
R1222 B.n758 B.n757 71.676
R1223 B.n761 B.n760 71.676
R1224 B.n766 B.n765 71.676
R1225 B.n769 B.n768 71.676
R1226 B.n774 B.n773 71.676
R1227 B.n777 B.n776 71.676
R1228 B.n782 B.n781 71.676
R1229 B.n785 B.n784 71.676
R1230 B.n790 B.n789 71.676
R1231 B.n793 B.n792 71.676
R1232 B.n798 B.n797 71.676
R1233 B.n801 B.n800 71.676
R1234 B.n806 B.n805 71.676
R1235 B.n809 B.n808 71.676
R1236 B.n814 B.n813 71.676
R1237 B.n817 B.n816 71.676
R1238 B.n822 B.n821 71.676
R1239 B.n825 B.n824 71.676
R1240 B.n562 B.n561 71.676
R1241 B.n564 B.n558 71.676
R1242 B.n571 B.n570 71.676
R1243 B.n572 B.n556 71.676
R1244 B.n579 B.n578 71.676
R1245 B.n580 B.n554 71.676
R1246 B.n587 B.n586 71.676
R1247 B.n588 B.n552 71.676
R1248 B.n595 B.n594 71.676
R1249 B.n596 B.n550 71.676
R1250 B.n603 B.n602 71.676
R1251 B.n604 B.n548 71.676
R1252 B.n611 B.n610 71.676
R1253 B.n612 B.n546 71.676
R1254 B.n619 B.n618 71.676
R1255 B.n620 B.n544 71.676
R1256 B.n627 B.n626 71.676
R1257 B.n628 B.n542 71.676
R1258 B.n635 B.n634 71.676
R1259 B.n636 B.n540 71.676
R1260 B.n643 B.n642 71.676
R1261 B.n644 B.n538 71.676
R1262 B.n651 B.n650 71.676
R1263 B.n652 B.n536 71.676
R1264 B.n659 B.n658 71.676
R1265 B.n660 B.n534 71.676
R1266 B.n667 B.n666 71.676
R1267 B.n668 B.n532 71.676
R1268 B.n675 B.n674 71.676
R1269 B.n676 B.n530 71.676
R1270 B.n686 B.n685 71.676
R1271 B.n687 B.n528 71.676
R1272 B.n694 B.n693 71.676
R1273 B.n695 B.n526 71.676
R1274 B.n702 B.n701 71.676
R1275 B.n703 B.n522 71.676
R1276 B.n711 B.n710 71.676
R1277 B.n712 B.n520 71.676
R1278 B.n719 B.n718 71.676
R1279 B.n720 B.n518 71.676
R1280 B.n727 B.n726 71.676
R1281 B.n728 B.n516 71.676
R1282 B.n735 B.n734 71.676
R1283 B.n736 B.n514 71.676
R1284 B.n743 B.n742 71.676
R1285 B.n744 B.n512 71.676
R1286 B.n751 B.n750 71.676
R1287 B.n752 B.n510 71.676
R1288 B.n759 B.n758 71.676
R1289 B.n760 B.n508 71.676
R1290 B.n767 B.n766 71.676
R1291 B.n768 B.n506 71.676
R1292 B.n775 B.n774 71.676
R1293 B.n776 B.n504 71.676
R1294 B.n783 B.n782 71.676
R1295 B.n784 B.n502 71.676
R1296 B.n791 B.n790 71.676
R1297 B.n792 B.n500 71.676
R1298 B.n799 B.n798 71.676
R1299 B.n800 B.n498 71.676
R1300 B.n807 B.n806 71.676
R1301 B.n808 B.n496 71.676
R1302 B.n815 B.n814 71.676
R1303 B.n816 B.n494 71.676
R1304 B.n823 B.n822 71.676
R1305 B.n826 B.n825 71.676
R1306 B.n1091 B.n1090 71.676
R1307 B.n1091 B.n2 71.676
R1308 B.n148 B.n147 71.5641
R1309 B.n145 B.n144 71.5641
R1310 B.n524 B.n523 71.5641
R1311 B.n681 B.n680 71.5641
R1312 B.n831 B.n490 61.1998
R1313 B.n1008 B.n1007 61.1998
R1314 B.n149 B.n148 59.5399
R1315 B.n146 B.n145 59.5399
R1316 B.n706 B.n524 59.5399
R1317 B.n682 B.n681 59.5399
R1318 B.n833 B.n488 33.8737
R1319 B.n829 B.n828 33.8737
R1320 B.n1004 B.n1003 33.8737
R1321 B.n1010 B.n74 33.8737
R1322 B.n831 B.n486 30.8268
R1323 B.n837 B.n486 30.8268
R1324 B.n837 B.n482 30.8268
R1325 B.n843 B.n482 30.8268
R1326 B.n843 B.n478 30.8268
R1327 B.n849 B.n478 30.8268
R1328 B.n849 B.n474 30.8268
R1329 B.n855 B.n474 30.8268
R1330 B.n861 B.n470 30.8268
R1331 B.n861 B.n466 30.8268
R1332 B.n867 B.n466 30.8268
R1333 B.n867 B.n462 30.8268
R1334 B.n873 B.n462 30.8268
R1335 B.n873 B.n458 30.8268
R1336 B.n879 B.n458 30.8268
R1337 B.n879 B.n454 30.8268
R1338 B.n885 B.n454 30.8268
R1339 B.n885 B.n450 30.8268
R1340 B.n891 B.n450 30.8268
R1341 B.n891 B.n446 30.8268
R1342 B.n897 B.n446 30.8268
R1343 B.n903 B.n442 30.8268
R1344 B.n903 B.n438 30.8268
R1345 B.n909 B.n438 30.8268
R1346 B.n909 B.n434 30.8268
R1347 B.n915 B.n434 30.8268
R1348 B.n915 B.n430 30.8268
R1349 B.n921 B.n430 30.8268
R1350 B.n921 B.n426 30.8268
R1351 B.n928 B.n426 30.8268
R1352 B.n928 B.n927 30.8268
R1353 B.n934 B.n419 30.8268
R1354 B.n941 B.n419 30.8268
R1355 B.n941 B.n415 30.8268
R1356 B.n947 B.n415 30.8268
R1357 B.n947 B.n4 30.8268
R1358 B.n1089 B.n4 30.8268
R1359 B.n1089 B.n1088 30.8268
R1360 B.n1088 B.n1087 30.8268
R1361 B.n1087 B.n8 30.8268
R1362 B.n12 B.n8 30.8268
R1363 B.n1080 B.n12 30.8268
R1364 B.n1080 B.n1079 30.8268
R1365 B.n1079 B.n1078 30.8268
R1366 B.n1072 B.n19 30.8268
R1367 B.n1072 B.n1071 30.8268
R1368 B.n1071 B.n1070 30.8268
R1369 B.n1070 B.n23 30.8268
R1370 B.n1064 B.n23 30.8268
R1371 B.n1064 B.n1063 30.8268
R1372 B.n1063 B.n1062 30.8268
R1373 B.n1062 B.n30 30.8268
R1374 B.n1056 B.n30 30.8268
R1375 B.n1056 B.n1055 30.8268
R1376 B.n1054 B.n37 30.8268
R1377 B.n1048 B.n37 30.8268
R1378 B.n1048 B.n1047 30.8268
R1379 B.n1047 B.n1046 30.8268
R1380 B.n1046 B.n44 30.8268
R1381 B.n1040 B.n44 30.8268
R1382 B.n1040 B.n1039 30.8268
R1383 B.n1039 B.n1038 30.8268
R1384 B.n1038 B.n51 30.8268
R1385 B.n1032 B.n51 30.8268
R1386 B.n1032 B.n1031 30.8268
R1387 B.n1031 B.n1030 30.8268
R1388 B.n1030 B.n58 30.8268
R1389 B.n1024 B.n1023 30.8268
R1390 B.n1023 B.n1022 30.8268
R1391 B.n1022 B.n65 30.8268
R1392 B.n1016 B.n65 30.8268
R1393 B.n1016 B.n1015 30.8268
R1394 B.n1015 B.n1014 30.8268
R1395 B.n1014 B.n72 30.8268
R1396 B.n1008 B.n72 30.8268
R1397 B.n897 B.t1 19.0403
R1398 B.t0 B.n1054 19.0403
R1399 B B.n1092 18.0485
R1400 B.n855 B.t5 17.227
R1401 B.n1024 B.t12 17.227
R1402 B.n934 B.t3 16.3203
R1403 B.n1078 B.t2 16.3203
R1404 B.n927 B.t3 14.507
R1405 B.n19 B.t2 14.507
R1406 B.t5 B.n470 13.6003
R1407 B.t12 B.n58 13.6003
R1408 B.t1 B.n442 11.787
R1409 B.n1055 B.t0 11.787
R1410 B.n834 B.n833 10.6151
R1411 B.n835 B.n834 10.6151
R1412 B.n835 B.n480 10.6151
R1413 B.n845 B.n480 10.6151
R1414 B.n846 B.n845 10.6151
R1415 B.n847 B.n846 10.6151
R1416 B.n847 B.n472 10.6151
R1417 B.n857 B.n472 10.6151
R1418 B.n858 B.n857 10.6151
R1419 B.n859 B.n858 10.6151
R1420 B.n859 B.n464 10.6151
R1421 B.n869 B.n464 10.6151
R1422 B.n870 B.n869 10.6151
R1423 B.n871 B.n870 10.6151
R1424 B.n871 B.n456 10.6151
R1425 B.n881 B.n456 10.6151
R1426 B.n882 B.n881 10.6151
R1427 B.n883 B.n882 10.6151
R1428 B.n883 B.n448 10.6151
R1429 B.n893 B.n448 10.6151
R1430 B.n894 B.n893 10.6151
R1431 B.n895 B.n894 10.6151
R1432 B.n895 B.n440 10.6151
R1433 B.n905 B.n440 10.6151
R1434 B.n906 B.n905 10.6151
R1435 B.n907 B.n906 10.6151
R1436 B.n907 B.n432 10.6151
R1437 B.n917 B.n432 10.6151
R1438 B.n918 B.n917 10.6151
R1439 B.n919 B.n918 10.6151
R1440 B.n919 B.n424 10.6151
R1441 B.n930 B.n424 10.6151
R1442 B.n931 B.n930 10.6151
R1443 B.n932 B.n931 10.6151
R1444 B.n932 B.n417 10.6151
R1445 B.n943 B.n417 10.6151
R1446 B.n944 B.n943 10.6151
R1447 B.n945 B.n944 10.6151
R1448 B.n945 B.n0 10.6151
R1449 B.n560 B.n488 10.6151
R1450 B.n560 B.n559 10.6151
R1451 B.n566 B.n559 10.6151
R1452 B.n567 B.n566 10.6151
R1453 B.n568 B.n567 10.6151
R1454 B.n568 B.n557 10.6151
R1455 B.n574 B.n557 10.6151
R1456 B.n575 B.n574 10.6151
R1457 B.n576 B.n575 10.6151
R1458 B.n576 B.n555 10.6151
R1459 B.n582 B.n555 10.6151
R1460 B.n583 B.n582 10.6151
R1461 B.n584 B.n583 10.6151
R1462 B.n584 B.n553 10.6151
R1463 B.n590 B.n553 10.6151
R1464 B.n591 B.n590 10.6151
R1465 B.n592 B.n591 10.6151
R1466 B.n592 B.n551 10.6151
R1467 B.n598 B.n551 10.6151
R1468 B.n599 B.n598 10.6151
R1469 B.n600 B.n599 10.6151
R1470 B.n600 B.n549 10.6151
R1471 B.n606 B.n549 10.6151
R1472 B.n607 B.n606 10.6151
R1473 B.n608 B.n607 10.6151
R1474 B.n608 B.n547 10.6151
R1475 B.n614 B.n547 10.6151
R1476 B.n615 B.n614 10.6151
R1477 B.n616 B.n615 10.6151
R1478 B.n616 B.n545 10.6151
R1479 B.n622 B.n545 10.6151
R1480 B.n623 B.n622 10.6151
R1481 B.n624 B.n623 10.6151
R1482 B.n624 B.n543 10.6151
R1483 B.n630 B.n543 10.6151
R1484 B.n631 B.n630 10.6151
R1485 B.n632 B.n631 10.6151
R1486 B.n632 B.n541 10.6151
R1487 B.n638 B.n541 10.6151
R1488 B.n639 B.n638 10.6151
R1489 B.n640 B.n639 10.6151
R1490 B.n640 B.n539 10.6151
R1491 B.n646 B.n539 10.6151
R1492 B.n647 B.n646 10.6151
R1493 B.n648 B.n647 10.6151
R1494 B.n648 B.n537 10.6151
R1495 B.n654 B.n537 10.6151
R1496 B.n655 B.n654 10.6151
R1497 B.n656 B.n655 10.6151
R1498 B.n656 B.n535 10.6151
R1499 B.n662 B.n535 10.6151
R1500 B.n663 B.n662 10.6151
R1501 B.n664 B.n663 10.6151
R1502 B.n664 B.n533 10.6151
R1503 B.n670 B.n533 10.6151
R1504 B.n671 B.n670 10.6151
R1505 B.n672 B.n671 10.6151
R1506 B.n672 B.n531 10.6151
R1507 B.n678 B.n531 10.6151
R1508 B.n679 B.n678 10.6151
R1509 B.n683 B.n679 10.6151
R1510 B.n689 B.n529 10.6151
R1511 B.n690 B.n689 10.6151
R1512 B.n691 B.n690 10.6151
R1513 B.n691 B.n527 10.6151
R1514 B.n697 B.n527 10.6151
R1515 B.n698 B.n697 10.6151
R1516 B.n699 B.n698 10.6151
R1517 B.n699 B.n525 10.6151
R1518 B.n705 B.n525 10.6151
R1519 B.n708 B.n707 10.6151
R1520 B.n708 B.n521 10.6151
R1521 B.n714 B.n521 10.6151
R1522 B.n715 B.n714 10.6151
R1523 B.n716 B.n715 10.6151
R1524 B.n716 B.n519 10.6151
R1525 B.n722 B.n519 10.6151
R1526 B.n723 B.n722 10.6151
R1527 B.n724 B.n723 10.6151
R1528 B.n724 B.n517 10.6151
R1529 B.n730 B.n517 10.6151
R1530 B.n731 B.n730 10.6151
R1531 B.n732 B.n731 10.6151
R1532 B.n732 B.n515 10.6151
R1533 B.n738 B.n515 10.6151
R1534 B.n739 B.n738 10.6151
R1535 B.n740 B.n739 10.6151
R1536 B.n740 B.n513 10.6151
R1537 B.n746 B.n513 10.6151
R1538 B.n747 B.n746 10.6151
R1539 B.n748 B.n747 10.6151
R1540 B.n748 B.n511 10.6151
R1541 B.n754 B.n511 10.6151
R1542 B.n755 B.n754 10.6151
R1543 B.n756 B.n755 10.6151
R1544 B.n756 B.n509 10.6151
R1545 B.n762 B.n509 10.6151
R1546 B.n763 B.n762 10.6151
R1547 B.n764 B.n763 10.6151
R1548 B.n764 B.n507 10.6151
R1549 B.n770 B.n507 10.6151
R1550 B.n771 B.n770 10.6151
R1551 B.n772 B.n771 10.6151
R1552 B.n772 B.n505 10.6151
R1553 B.n778 B.n505 10.6151
R1554 B.n779 B.n778 10.6151
R1555 B.n780 B.n779 10.6151
R1556 B.n780 B.n503 10.6151
R1557 B.n786 B.n503 10.6151
R1558 B.n787 B.n786 10.6151
R1559 B.n788 B.n787 10.6151
R1560 B.n788 B.n501 10.6151
R1561 B.n794 B.n501 10.6151
R1562 B.n795 B.n794 10.6151
R1563 B.n796 B.n795 10.6151
R1564 B.n796 B.n499 10.6151
R1565 B.n802 B.n499 10.6151
R1566 B.n803 B.n802 10.6151
R1567 B.n804 B.n803 10.6151
R1568 B.n804 B.n497 10.6151
R1569 B.n810 B.n497 10.6151
R1570 B.n811 B.n810 10.6151
R1571 B.n812 B.n811 10.6151
R1572 B.n812 B.n495 10.6151
R1573 B.n818 B.n495 10.6151
R1574 B.n819 B.n818 10.6151
R1575 B.n820 B.n819 10.6151
R1576 B.n820 B.n493 10.6151
R1577 B.n493 B.n492 10.6151
R1578 B.n827 B.n492 10.6151
R1579 B.n828 B.n827 10.6151
R1580 B.n829 B.n484 10.6151
R1581 B.n839 B.n484 10.6151
R1582 B.n840 B.n839 10.6151
R1583 B.n841 B.n840 10.6151
R1584 B.n841 B.n476 10.6151
R1585 B.n851 B.n476 10.6151
R1586 B.n852 B.n851 10.6151
R1587 B.n853 B.n852 10.6151
R1588 B.n853 B.n468 10.6151
R1589 B.n863 B.n468 10.6151
R1590 B.n864 B.n863 10.6151
R1591 B.n865 B.n864 10.6151
R1592 B.n865 B.n460 10.6151
R1593 B.n875 B.n460 10.6151
R1594 B.n876 B.n875 10.6151
R1595 B.n877 B.n876 10.6151
R1596 B.n877 B.n452 10.6151
R1597 B.n887 B.n452 10.6151
R1598 B.n888 B.n887 10.6151
R1599 B.n889 B.n888 10.6151
R1600 B.n889 B.n444 10.6151
R1601 B.n899 B.n444 10.6151
R1602 B.n900 B.n899 10.6151
R1603 B.n901 B.n900 10.6151
R1604 B.n901 B.n436 10.6151
R1605 B.n911 B.n436 10.6151
R1606 B.n912 B.n911 10.6151
R1607 B.n913 B.n912 10.6151
R1608 B.n913 B.n428 10.6151
R1609 B.n923 B.n428 10.6151
R1610 B.n924 B.n923 10.6151
R1611 B.n925 B.n924 10.6151
R1612 B.n925 B.n421 10.6151
R1613 B.n936 B.n421 10.6151
R1614 B.n937 B.n936 10.6151
R1615 B.n939 B.n937 10.6151
R1616 B.n939 B.n938 10.6151
R1617 B.n938 B.n413 10.6151
R1618 B.n950 B.n413 10.6151
R1619 B.n951 B.n950 10.6151
R1620 B.n952 B.n951 10.6151
R1621 B.n953 B.n952 10.6151
R1622 B.n954 B.n953 10.6151
R1623 B.n957 B.n954 10.6151
R1624 B.n958 B.n957 10.6151
R1625 B.n959 B.n958 10.6151
R1626 B.n960 B.n959 10.6151
R1627 B.n962 B.n960 10.6151
R1628 B.n963 B.n962 10.6151
R1629 B.n964 B.n963 10.6151
R1630 B.n965 B.n964 10.6151
R1631 B.n967 B.n965 10.6151
R1632 B.n968 B.n967 10.6151
R1633 B.n969 B.n968 10.6151
R1634 B.n970 B.n969 10.6151
R1635 B.n972 B.n970 10.6151
R1636 B.n973 B.n972 10.6151
R1637 B.n974 B.n973 10.6151
R1638 B.n975 B.n974 10.6151
R1639 B.n977 B.n975 10.6151
R1640 B.n978 B.n977 10.6151
R1641 B.n979 B.n978 10.6151
R1642 B.n980 B.n979 10.6151
R1643 B.n982 B.n980 10.6151
R1644 B.n983 B.n982 10.6151
R1645 B.n984 B.n983 10.6151
R1646 B.n985 B.n984 10.6151
R1647 B.n987 B.n985 10.6151
R1648 B.n988 B.n987 10.6151
R1649 B.n989 B.n988 10.6151
R1650 B.n990 B.n989 10.6151
R1651 B.n992 B.n990 10.6151
R1652 B.n993 B.n992 10.6151
R1653 B.n994 B.n993 10.6151
R1654 B.n995 B.n994 10.6151
R1655 B.n997 B.n995 10.6151
R1656 B.n998 B.n997 10.6151
R1657 B.n999 B.n998 10.6151
R1658 B.n1000 B.n999 10.6151
R1659 B.n1002 B.n1000 10.6151
R1660 B.n1003 B.n1002 10.6151
R1661 B.n1084 B.n1 10.6151
R1662 B.n1084 B.n1083 10.6151
R1663 B.n1083 B.n1082 10.6151
R1664 B.n1082 B.n10 10.6151
R1665 B.n1076 B.n10 10.6151
R1666 B.n1076 B.n1075 10.6151
R1667 B.n1075 B.n1074 10.6151
R1668 B.n1074 B.n17 10.6151
R1669 B.n1068 B.n17 10.6151
R1670 B.n1068 B.n1067 10.6151
R1671 B.n1067 B.n1066 10.6151
R1672 B.n1066 B.n25 10.6151
R1673 B.n1060 B.n25 10.6151
R1674 B.n1060 B.n1059 10.6151
R1675 B.n1059 B.n1058 10.6151
R1676 B.n1058 B.n32 10.6151
R1677 B.n1052 B.n32 10.6151
R1678 B.n1052 B.n1051 10.6151
R1679 B.n1051 B.n1050 10.6151
R1680 B.n1050 B.n39 10.6151
R1681 B.n1044 B.n39 10.6151
R1682 B.n1044 B.n1043 10.6151
R1683 B.n1043 B.n1042 10.6151
R1684 B.n1042 B.n46 10.6151
R1685 B.n1036 B.n46 10.6151
R1686 B.n1036 B.n1035 10.6151
R1687 B.n1035 B.n1034 10.6151
R1688 B.n1034 B.n53 10.6151
R1689 B.n1028 B.n53 10.6151
R1690 B.n1028 B.n1027 10.6151
R1691 B.n1027 B.n1026 10.6151
R1692 B.n1026 B.n60 10.6151
R1693 B.n1020 B.n60 10.6151
R1694 B.n1020 B.n1019 10.6151
R1695 B.n1019 B.n1018 10.6151
R1696 B.n1018 B.n67 10.6151
R1697 B.n1012 B.n67 10.6151
R1698 B.n1012 B.n1011 10.6151
R1699 B.n1011 B.n1010 10.6151
R1700 B.n150 B.n74 10.6151
R1701 B.n153 B.n150 10.6151
R1702 B.n154 B.n153 10.6151
R1703 B.n157 B.n154 10.6151
R1704 B.n158 B.n157 10.6151
R1705 B.n161 B.n158 10.6151
R1706 B.n162 B.n161 10.6151
R1707 B.n165 B.n162 10.6151
R1708 B.n166 B.n165 10.6151
R1709 B.n169 B.n166 10.6151
R1710 B.n170 B.n169 10.6151
R1711 B.n173 B.n170 10.6151
R1712 B.n174 B.n173 10.6151
R1713 B.n177 B.n174 10.6151
R1714 B.n178 B.n177 10.6151
R1715 B.n181 B.n178 10.6151
R1716 B.n182 B.n181 10.6151
R1717 B.n185 B.n182 10.6151
R1718 B.n186 B.n185 10.6151
R1719 B.n189 B.n186 10.6151
R1720 B.n190 B.n189 10.6151
R1721 B.n193 B.n190 10.6151
R1722 B.n194 B.n193 10.6151
R1723 B.n197 B.n194 10.6151
R1724 B.n198 B.n197 10.6151
R1725 B.n201 B.n198 10.6151
R1726 B.n202 B.n201 10.6151
R1727 B.n205 B.n202 10.6151
R1728 B.n206 B.n205 10.6151
R1729 B.n209 B.n206 10.6151
R1730 B.n210 B.n209 10.6151
R1731 B.n213 B.n210 10.6151
R1732 B.n214 B.n213 10.6151
R1733 B.n217 B.n214 10.6151
R1734 B.n218 B.n217 10.6151
R1735 B.n221 B.n218 10.6151
R1736 B.n222 B.n221 10.6151
R1737 B.n225 B.n222 10.6151
R1738 B.n226 B.n225 10.6151
R1739 B.n229 B.n226 10.6151
R1740 B.n230 B.n229 10.6151
R1741 B.n233 B.n230 10.6151
R1742 B.n234 B.n233 10.6151
R1743 B.n237 B.n234 10.6151
R1744 B.n238 B.n237 10.6151
R1745 B.n241 B.n238 10.6151
R1746 B.n242 B.n241 10.6151
R1747 B.n245 B.n242 10.6151
R1748 B.n246 B.n245 10.6151
R1749 B.n249 B.n246 10.6151
R1750 B.n250 B.n249 10.6151
R1751 B.n253 B.n250 10.6151
R1752 B.n254 B.n253 10.6151
R1753 B.n257 B.n254 10.6151
R1754 B.n258 B.n257 10.6151
R1755 B.n261 B.n258 10.6151
R1756 B.n262 B.n261 10.6151
R1757 B.n265 B.n262 10.6151
R1758 B.n266 B.n265 10.6151
R1759 B.n269 B.n266 10.6151
R1760 B.n270 B.n269 10.6151
R1761 B.n274 B.n273 10.6151
R1762 B.n277 B.n274 10.6151
R1763 B.n278 B.n277 10.6151
R1764 B.n281 B.n278 10.6151
R1765 B.n282 B.n281 10.6151
R1766 B.n285 B.n282 10.6151
R1767 B.n286 B.n285 10.6151
R1768 B.n289 B.n286 10.6151
R1769 B.n290 B.n289 10.6151
R1770 B.n294 B.n293 10.6151
R1771 B.n297 B.n294 10.6151
R1772 B.n298 B.n297 10.6151
R1773 B.n301 B.n298 10.6151
R1774 B.n302 B.n301 10.6151
R1775 B.n305 B.n302 10.6151
R1776 B.n306 B.n305 10.6151
R1777 B.n309 B.n306 10.6151
R1778 B.n310 B.n309 10.6151
R1779 B.n313 B.n310 10.6151
R1780 B.n314 B.n313 10.6151
R1781 B.n317 B.n314 10.6151
R1782 B.n318 B.n317 10.6151
R1783 B.n321 B.n318 10.6151
R1784 B.n322 B.n321 10.6151
R1785 B.n325 B.n322 10.6151
R1786 B.n326 B.n325 10.6151
R1787 B.n329 B.n326 10.6151
R1788 B.n330 B.n329 10.6151
R1789 B.n333 B.n330 10.6151
R1790 B.n334 B.n333 10.6151
R1791 B.n337 B.n334 10.6151
R1792 B.n338 B.n337 10.6151
R1793 B.n341 B.n338 10.6151
R1794 B.n342 B.n341 10.6151
R1795 B.n345 B.n342 10.6151
R1796 B.n346 B.n345 10.6151
R1797 B.n349 B.n346 10.6151
R1798 B.n350 B.n349 10.6151
R1799 B.n353 B.n350 10.6151
R1800 B.n354 B.n353 10.6151
R1801 B.n357 B.n354 10.6151
R1802 B.n358 B.n357 10.6151
R1803 B.n361 B.n358 10.6151
R1804 B.n362 B.n361 10.6151
R1805 B.n365 B.n362 10.6151
R1806 B.n366 B.n365 10.6151
R1807 B.n369 B.n366 10.6151
R1808 B.n370 B.n369 10.6151
R1809 B.n373 B.n370 10.6151
R1810 B.n374 B.n373 10.6151
R1811 B.n377 B.n374 10.6151
R1812 B.n378 B.n377 10.6151
R1813 B.n381 B.n378 10.6151
R1814 B.n382 B.n381 10.6151
R1815 B.n385 B.n382 10.6151
R1816 B.n386 B.n385 10.6151
R1817 B.n389 B.n386 10.6151
R1818 B.n390 B.n389 10.6151
R1819 B.n393 B.n390 10.6151
R1820 B.n394 B.n393 10.6151
R1821 B.n397 B.n394 10.6151
R1822 B.n398 B.n397 10.6151
R1823 B.n401 B.n398 10.6151
R1824 B.n402 B.n401 10.6151
R1825 B.n405 B.n402 10.6151
R1826 B.n406 B.n405 10.6151
R1827 B.n409 B.n406 10.6151
R1828 B.n411 B.n409 10.6151
R1829 B.n412 B.n411 10.6151
R1830 B.n1004 B.n412 10.6151
R1831 B.n683 B.n682 9.36635
R1832 B.n707 B.n706 9.36635
R1833 B.n270 B.n149 9.36635
R1834 B.n293 B.n146 9.36635
R1835 B.n1092 B.n0 8.11757
R1836 B.n1092 B.n1 8.11757
R1837 B.n682 B.n529 1.24928
R1838 B.n706 B.n705 1.24928
R1839 B.n273 B.n149 1.24928
R1840 B.n290 B.n146 1.24928
R1841 VN.n1 VN.t1 171.273
R1842 VN.n0 VN.t3 171.273
R1843 VN.n0 VN.t2 170.139
R1844 VN.n1 VN.t0 170.139
R1845 VN VN.n1 56.6228
R1846 VN VN.n0 2.40691
R1847 VDD2.n2 VDD2.n0 110.832
R1848 VDD2.n2 VDD2.n1 61.2036
R1849 VDD2.n1 VDD2.t1 1.04315
R1850 VDD2.n1 VDD2.t0 1.04315
R1851 VDD2.n0 VDD2.t2 1.04315
R1852 VDD2.n0 VDD2.t3 1.04315
R1853 VDD2 VDD2.n2 0.0586897
R1854 VTAIL.n842 VTAIL.n742 289.615
R1855 VTAIL.n100 VTAIL.n0 289.615
R1856 VTAIL.n206 VTAIL.n106 289.615
R1857 VTAIL.n312 VTAIL.n212 289.615
R1858 VTAIL.n736 VTAIL.n636 289.615
R1859 VTAIL.n630 VTAIL.n530 289.615
R1860 VTAIL.n524 VTAIL.n424 289.615
R1861 VTAIL.n418 VTAIL.n318 289.615
R1862 VTAIL.n777 VTAIL.n776 185
R1863 VTAIL.n774 VTAIL.n773 185
R1864 VTAIL.n783 VTAIL.n782 185
R1865 VTAIL.n785 VTAIL.n784 185
R1866 VTAIL.n770 VTAIL.n769 185
R1867 VTAIL.n791 VTAIL.n790 185
R1868 VTAIL.n793 VTAIL.n792 185
R1869 VTAIL.n766 VTAIL.n765 185
R1870 VTAIL.n799 VTAIL.n798 185
R1871 VTAIL.n801 VTAIL.n800 185
R1872 VTAIL.n762 VTAIL.n761 185
R1873 VTAIL.n807 VTAIL.n806 185
R1874 VTAIL.n809 VTAIL.n808 185
R1875 VTAIL.n758 VTAIL.n757 185
R1876 VTAIL.n815 VTAIL.n814 185
R1877 VTAIL.n818 VTAIL.n817 185
R1878 VTAIL.n816 VTAIL.n754 185
R1879 VTAIL.n823 VTAIL.n753 185
R1880 VTAIL.n825 VTAIL.n824 185
R1881 VTAIL.n827 VTAIL.n826 185
R1882 VTAIL.n750 VTAIL.n749 185
R1883 VTAIL.n833 VTAIL.n832 185
R1884 VTAIL.n835 VTAIL.n834 185
R1885 VTAIL.n746 VTAIL.n745 185
R1886 VTAIL.n841 VTAIL.n840 185
R1887 VTAIL.n843 VTAIL.n842 185
R1888 VTAIL.n35 VTAIL.n34 185
R1889 VTAIL.n32 VTAIL.n31 185
R1890 VTAIL.n41 VTAIL.n40 185
R1891 VTAIL.n43 VTAIL.n42 185
R1892 VTAIL.n28 VTAIL.n27 185
R1893 VTAIL.n49 VTAIL.n48 185
R1894 VTAIL.n51 VTAIL.n50 185
R1895 VTAIL.n24 VTAIL.n23 185
R1896 VTAIL.n57 VTAIL.n56 185
R1897 VTAIL.n59 VTAIL.n58 185
R1898 VTAIL.n20 VTAIL.n19 185
R1899 VTAIL.n65 VTAIL.n64 185
R1900 VTAIL.n67 VTAIL.n66 185
R1901 VTAIL.n16 VTAIL.n15 185
R1902 VTAIL.n73 VTAIL.n72 185
R1903 VTAIL.n76 VTAIL.n75 185
R1904 VTAIL.n74 VTAIL.n12 185
R1905 VTAIL.n81 VTAIL.n11 185
R1906 VTAIL.n83 VTAIL.n82 185
R1907 VTAIL.n85 VTAIL.n84 185
R1908 VTAIL.n8 VTAIL.n7 185
R1909 VTAIL.n91 VTAIL.n90 185
R1910 VTAIL.n93 VTAIL.n92 185
R1911 VTAIL.n4 VTAIL.n3 185
R1912 VTAIL.n99 VTAIL.n98 185
R1913 VTAIL.n101 VTAIL.n100 185
R1914 VTAIL.n141 VTAIL.n140 185
R1915 VTAIL.n138 VTAIL.n137 185
R1916 VTAIL.n147 VTAIL.n146 185
R1917 VTAIL.n149 VTAIL.n148 185
R1918 VTAIL.n134 VTAIL.n133 185
R1919 VTAIL.n155 VTAIL.n154 185
R1920 VTAIL.n157 VTAIL.n156 185
R1921 VTAIL.n130 VTAIL.n129 185
R1922 VTAIL.n163 VTAIL.n162 185
R1923 VTAIL.n165 VTAIL.n164 185
R1924 VTAIL.n126 VTAIL.n125 185
R1925 VTAIL.n171 VTAIL.n170 185
R1926 VTAIL.n173 VTAIL.n172 185
R1927 VTAIL.n122 VTAIL.n121 185
R1928 VTAIL.n179 VTAIL.n178 185
R1929 VTAIL.n182 VTAIL.n181 185
R1930 VTAIL.n180 VTAIL.n118 185
R1931 VTAIL.n187 VTAIL.n117 185
R1932 VTAIL.n189 VTAIL.n188 185
R1933 VTAIL.n191 VTAIL.n190 185
R1934 VTAIL.n114 VTAIL.n113 185
R1935 VTAIL.n197 VTAIL.n196 185
R1936 VTAIL.n199 VTAIL.n198 185
R1937 VTAIL.n110 VTAIL.n109 185
R1938 VTAIL.n205 VTAIL.n204 185
R1939 VTAIL.n207 VTAIL.n206 185
R1940 VTAIL.n247 VTAIL.n246 185
R1941 VTAIL.n244 VTAIL.n243 185
R1942 VTAIL.n253 VTAIL.n252 185
R1943 VTAIL.n255 VTAIL.n254 185
R1944 VTAIL.n240 VTAIL.n239 185
R1945 VTAIL.n261 VTAIL.n260 185
R1946 VTAIL.n263 VTAIL.n262 185
R1947 VTAIL.n236 VTAIL.n235 185
R1948 VTAIL.n269 VTAIL.n268 185
R1949 VTAIL.n271 VTAIL.n270 185
R1950 VTAIL.n232 VTAIL.n231 185
R1951 VTAIL.n277 VTAIL.n276 185
R1952 VTAIL.n279 VTAIL.n278 185
R1953 VTAIL.n228 VTAIL.n227 185
R1954 VTAIL.n285 VTAIL.n284 185
R1955 VTAIL.n288 VTAIL.n287 185
R1956 VTAIL.n286 VTAIL.n224 185
R1957 VTAIL.n293 VTAIL.n223 185
R1958 VTAIL.n295 VTAIL.n294 185
R1959 VTAIL.n297 VTAIL.n296 185
R1960 VTAIL.n220 VTAIL.n219 185
R1961 VTAIL.n303 VTAIL.n302 185
R1962 VTAIL.n305 VTAIL.n304 185
R1963 VTAIL.n216 VTAIL.n215 185
R1964 VTAIL.n311 VTAIL.n310 185
R1965 VTAIL.n313 VTAIL.n312 185
R1966 VTAIL.n737 VTAIL.n736 185
R1967 VTAIL.n735 VTAIL.n734 185
R1968 VTAIL.n640 VTAIL.n639 185
R1969 VTAIL.n729 VTAIL.n728 185
R1970 VTAIL.n727 VTAIL.n726 185
R1971 VTAIL.n644 VTAIL.n643 185
R1972 VTAIL.n721 VTAIL.n720 185
R1973 VTAIL.n719 VTAIL.n718 185
R1974 VTAIL.n717 VTAIL.n647 185
R1975 VTAIL.n651 VTAIL.n648 185
R1976 VTAIL.n712 VTAIL.n711 185
R1977 VTAIL.n710 VTAIL.n709 185
R1978 VTAIL.n653 VTAIL.n652 185
R1979 VTAIL.n704 VTAIL.n703 185
R1980 VTAIL.n702 VTAIL.n701 185
R1981 VTAIL.n657 VTAIL.n656 185
R1982 VTAIL.n696 VTAIL.n695 185
R1983 VTAIL.n694 VTAIL.n693 185
R1984 VTAIL.n661 VTAIL.n660 185
R1985 VTAIL.n688 VTAIL.n687 185
R1986 VTAIL.n686 VTAIL.n685 185
R1987 VTAIL.n665 VTAIL.n664 185
R1988 VTAIL.n680 VTAIL.n679 185
R1989 VTAIL.n678 VTAIL.n677 185
R1990 VTAIL.n669 VTAIL.n668 185
R1991 VTAIL.n672 VTAIL.n671 185
R1992 VTAIL.n631 VTAIL.n630 185
R1993 VTAIL.n629 VTAIL.n628 185
R1994 VTAIL.n534 VTAIL.n533 185
R1995 VTAIL.n623 VTAIL.n622 185
R1996 VTAIL.n621 VTAIL.n620 185
R1997 VTAIL.n538 VTAIL.n537 185
R1998 VTAIL.n615 VTAIL.n614 185
R1999 VTAIL.n613 VTAIL.n612 185
R2000 VTAIL.n611 VTAIL.n541 185
R2001 VTAIL.n545 VTAIL.n542 185
R2002 VTAIL.n606 VTAIL.n605 185
R2003 VTAIL.n604 VTAIL.n603 185
R2004 VTAIL.n547 VTAIL.n546 185
R2005 VTAIL.n598 VTAIL.n597 185
R2006 VTAIL.n596 VTAIL.n595 185
R2007 VTAIL.n551 VTAIL.n550 185
R2008 VTAIL.n590 VTAIL.n589 185
R2009 VTAIL.n588 VTAIL.n587 185
R2010 VTAIL.n555 VTAIL.n554 185
R2011 VTAIL.n582 VTAIL.n581 185
R2012 VTAIL.n580 VTAIL.n579 185
R2013 VTAIL.n559 VTAIL.n558 185
R2014 VTAIL.n574 VTAIL.n573 185
R2015 VTAIL.n572 VTAIL.n571 185
R2016 VTAIL.n563 VTAIL.n562 185
R2017 VTAIL.n566 VTAIL.n565 185
R2018 VTAIL.n525 VTAIL.n524 185
R2019 VTAIL.n523 VTAIL.n522 185
R2020 VTAIL.n428 VTAIL.n427 185
R2021 VTAIL.n517 VTAIL.n516 185
R2022 VTAIL.n515 VTAIL.n514 185
R2023 VTAIL.n432 VTAIL.n431 185
R2024 VTAIL.n509 VTAIL.n508 185
R2025 VTAIL.n507 VTAIL.n506 185
R2026 VTAIL.n505 VTAIL.n435 185
R2027 VTAIL.n439 VTAIL.n436 185
R2028 VTAIL.n500 VTAIL.n499 185
R2029 VTAIL.n498 VTAIL.n497 185
R2030 VTAIL.n441 VTAIL.n440 185
R2031 VTAIL.n492 VTAIL.n491 185
R2032 VTAIL.n490 VTAIL.n489 185
R2033 VTAIL.n445 VTAIL.n444 185
R2034 VTAIL.n484 VTAIL.n483 185
R2035 VTAIL.n482 VTAIL.n481 185
R2036 VTAIL.n449 VTAIL.n448 185
R2037 VTAIL.n476 VTAIL.n475 185
R2038 VTAIL.n474 VTAIL.n473 185
R2039 VTAIL.n453 VTAIL.n452 185
R2040 VTAIL.n468 VTAIL.n467 185
R2041 VTAIL.n466 VTAIL.n465 185
R2042 VTAIL.n457 VTAIL.n456 185
R2043 VTAIL.n460 VTAIL.n459 185
R2044 VTAIL.n419 VTAIL.n418 185
R2045 VTAIL.n417 VTAIL.n416 185
R2046 VTAIL.n322 VTAIL.n321 185
R2047 VTAIL.n411 VTAIL.n410 185
R2048 VTAIL.n409 VTAIL.n408 185
R2049 VTAIL.n326 VTAIL.n325 185
R2050 VTAIL.n403 VTAIL.n402 185
R2051 VTAIL.n401 VTAIL.n400 185
R2052 VTAIL.n399 VTAIL.n329 185
R2053 VTAIL.n333 VTAIL.n330 185
R2054 VTAIL.n394 VTAIL.n393 185
R2055 VTAIL.n392 VTAIL.n391 185
R2056 VTAIL.n335 VTAIL.n334 185
R2057 VTAIL.n386 VTAIL.n385 185
R2058 VTAIL.n384 VTAIL.n383 185
R2059 VTAIL.n339 VTAIL.n338 185
R2060 VTAIL.n378 VTAIL.n377 185
R2061 VTAIL.n376 VTAIL.n375 185
R2062 VTAIL.n343 VTAIL.n342 185
R2063 VTAIL.n370 VTAIL.n369 185
R2064 VTAIL.n368 VTAIL.n367 185
R2065 VTAIL.n347 VTAIL.n346 185
R2066 VTAIL.n362 VTAIL.n361 185
R2067 VTAIL.n360 VTAIL.n359 185
R2068 VTAIL.n351 VTAIL.n350 185
R2069 VTAIL.n354 VTAIL.n353 185
R2070 VTAIL.t3 VTAIL.n670 147.659
R2071 VTAIL.t1 VTAIL.n564 147.659
R2072 VTAIL.t6 VTAIL.n458 147.659
R2073 VTAIL.t7 VTAIL.n352 147.659
R2074 VTAIL.t5 VTAIL.n775 147.659
R2075 VTAIL.t4 VTAIL.n33 147.659
R2076 VTAIL.t2 VTAIL.n139 147.659
R2077 VTAIL.t0 VTAIL.n245 147.659
R2078 VTAIL.n776 VTAIL.n773 104.615
R2079 VTAIL.n783 VTAIL.n773 104.615
R2080 VTAIL.n784 VTAIL.n783 104.615
R2081 VTAIL.n784 VTAIL.n769 104.615
R2082 VTAIL.n791 VTAIL.n769 104.615
R2083 VTAIL.n792 VTAIL.n791 104.615
R2084 VTAIL.n792 VTAIL.n765 104.615
R2085 VTAIL.n799 VTAIL.n765 104.615
R2086 VTAIL.n800 VTAIL.n799 104.615
R2087 VTAIL.n800 VTAIL.n761 104.615
R2088 VTAIL.n807 VTAIL.n761 104.615
R2089 VTAIL.n808 VTAIL.n807 104.615
R2090 VTAIL.n808 VTAIL.n757 104.615
R2091 VTAIL.n815 VTAIL.n757 104.615
R2092 VTAIL.n817 VTAIL.n815 104.615
R2093 VTAIL.n817 VTAIL.n816 104.615
R2094 VTAIL.n816 VTAIL.n753 104.615
R2095 VTAIL.n825 VTAIL.n753 104.615
R2096 VTAIL.n826 VTAIL.n825 104.615
R2097 VTAIL.n826 VTAIL.n749 104.615
R2098 VTAIL.n833 VTAIL.n749 104.615
R2099 VTAIL.n834 VTAIL.n833 104.615
R2100 VTAIL.n834 VTAIL.n745 104.615
R2101 VTAIL.n841 VTAIL.n745 104.615
R2102 VTAIL.n842 VTAIL.n841 104.615
R2103 VTAIL.n34 VTAIL.n31 104.615
R2104 VTAIL.n41 VTAIL.n31 104.615
R2105 VTAIL.n42 VTAIL.n41 104.615
R2106 VTAIL.n42 VTAIL.n27 104.615
R2107 VTAIL.n49 VTAIL.n27 104.615
R2108 VTAIL.n50 VTAIL.n49 104.615
R2109 VTAIL.n50 VTAIL.n23 104.615
R2110 VTAIL.n57 VTAIL.n23 104.615
R2111 VTAIL.n58 VTAIL.n57 104.615
R2112 VTAIL.n58 VTAIL.n19 104.615
R2113 VTAIL.n65 VTAIL.n19 104.615
R2114 VTAIL.n66 VTAIL.n65 104.615
R2115 VTAIL.n66 VTAIL.n15 104.615
R2116 VTAIL.n73 VTAIL.n15 104.615
R2117 VTAIL.n75 VTAIL.n73 104.615
R2118 VTAIL.n75 VTAIL.n74 104.615
R2119 VTAIL.n74 VTAIL.n11 104.615
R2120 VTAIL.n83 VTAIL.n11 104.615
R2121 VTAIL.n84 VTAIL.n83 104.615
R2122 VTAIL.n84 VTAIL.n7 104.615
R2123 VTAIL.n91 VTAIL.n7 104.615
R2124 VTAIL.n92 VTAIL.n91 104.615
R2125 VTAIL.n92 VTAIL.n3 104.615
R2126 VTAIL.n99 VTAIL.n3 104.615
R2127 VTAIL.n100 VTAIL.n99 104.615
R2128 VTAIL.n140 VTAIL.n137 104.615
R2129 VTAIL.n147 VTAIL.n137 104.615
R2130 VTAIL.n148 VTAIL.n147 104.615
R2131 VTAIL.n148 VTAIL.n133 104.615
R2132 VTAIL.n155 VTAIL.n133 104.615
R2133 VTAIL.n156 VTAIL.n155 104.615
R2134 VTAIL.n156 VTAIL.n129 104.615
R2135 VTAIL.n163 VTAIL.n129 104.615
R2136 VTAIL.n164 VTAIL.n163 104.615
R2137 VTAIL.n164 VTAIL.n125 104.615
R2138 VTAIL.n171 VTAIL.n125 104.615
R2139 VTAIL.n172 VTAIL.n171 104.615
R2140 VTAIL.n172 VTAIL.n121 104.615
R2141 VTAIL.n179 VTAIL.n121 104.615
R2142 VTAIL.n181 VTAIL.n179 104.615
R2143 VTAIL.n181 VTAIL.n180 104.615
R2144 VTAIL.n180 VTAIL.n117 104.615
R2145 VTAIL.n189 VTAIL.n117 104.615
R2146 VTAIL.n190 VTAIL.n189 104.615
R2147 VTAIL.n190 VTAIL.n113 104.615
R2148 VTAIL.n197 VTAIL.n113 104.615
R2149 VTAIL.n198 VTAIL.n197 104.615
R2150 VTAIL.n198 VTAIL.n109 104.615
R2151 VTAIL.n205 VTAIL.n109 104.615
R2152 VTAIL.n206 VTAIL.n205 104.615
R2153 VTAIL.n246 VTAIL.n243 104.615
R2154 VTAIL.n253 VTAIL.n243 104.615
R2155 VTAIL.n254 VTAIL.n253 104.615
R2156 VTAIL.n254 VTAIL.n239 104.615
R2157 VTAIL.n261 VTAIL.n239 104.615
R2158 VTAIL.n262 VTAIL.n261 104.615
R2159 VTAIL.n262 VTAIL.n235 104.615
R2160 VTAIL.n269 VTAIL.n235 104.615
R2161 VTAIL.n270 VTAIL.n269 104.615
R2162 VTAIL.n270 VTAIL.n231 104.615
R2163 VTAIL.n277 VTAIL.n231 104.615
R2164 VTAIL.n278 VTAIL.n277 104.615
R2165 VTAIL.n278 VTAIL.n227 104.615
R2166 VTAIL.n285 VTAIL.n227 104.615
R2167 VTAIL.n287 VTAIL.n285 104.615
R2168 VTAIL.n287 VTAIL.n286 104.615
R2169 VTAIL.n286 VTAIL.n223 104.615
R2170 VTAIL.n295 VTAIL.n223 104.615
R2171 VTAIL.n296 VTAIL.n295 104.615
R2172 VTAIL.n296 VTAIL.n219 104.615
R2173 VTAIL.n303 VTAIL.n219 104.615
R2174 VTAIL.n304 VTAIL.n303 104.615
R2175 VTAIL.n304 VTAIL.n215 104.615
R2176 VTAIL.n311 VTAIL.n215 104.615
R2177 VTAIL.n312 VTAIL.n311 104.615
R2178 VTAIL.n736 VTAIL.n735 104.615
R2179 VTAIL.n735 VTAIL.n639 104.615
R2180 VTAIL.n728 VTAIL.n639 104.615
R2181 VTAIL.n728 VTAIL.n727 104.615
R2182 VTAIL.n727 VTAIL.n643 104.615
R2183 VTAIL.n720 VTAIL.n643 104.615
R2184 VTAIL.n720 VTAIL.n719 104.615
R2185 VTAIL.n719 VTAIL.n647 104.615
R2186 VTAIL.n651 VTAIL.n647 104.615
R2187 VTAIL.n711 VTAIL.n651 104.615
R2188 VTAIL.n711 VTAIL.n710 104.615
R2189 VTAIL.n710 VTAIL.n652 104.615
R2190 VTAIL.n703 VTAIL.n652 104.615
R2191 VTAIL.n703 VTAIL.n702 104.615
R2192 VTAIL.n702 VTAIL.n656 104.615
R2193 VTAIL.n695 VTAIL.n656 104.615
R2194 VTAIL.n695 VTAIL.n694 104.615
R2195 VTAIL.n694 VTAIL.n660 104.615
R2196 VTAIL.n687 VTAIL.n660 104.615
R2197 VTAIL.n687 VTAIL.n686 104.615
R2198 VTAIL.n686 VTAIL.n664 104.615
R2199 VTAIL.n679 VTAIL.n664 104.615
R2200 VTAIL.n679 VTAIL.n678 104.615
R2201 VTAIL.n678 VTAIL.n668 104.615
R2202 VTAIL.n671 VTAIL.n668 104.615
R2203 VTAIL.n630 VTAIL.n629 104.615
R2204 VTAIL.n629 VTAIL.n533 104.615
R2205 VTAIL.n622 VTAIL.n533 104.615
R2206 VTAIL.n622 VTAIL.n621 104.615
R2207 VTAIL.n621 VTAIL.n537 104.615
R2208 VTAIL.n614 VTAIL.n537 104.615
R2209 VTAIL.n614 VTAIL.n613 104.615
R2210 VTAIL.n613 VTAIL.n541 104.615
R2211 VTAIL.n545 VTAIL.n541 104.615
R2212 VTAIL.n605 VTAIL.n545 104.615
R2213 VTAIL.n605 VTAIL.n604 104.615
R2214 VTAIL.n604 VTAIL.n546 104.615
R2215 VTAIL.n597 VTAIL.n546 104.615
R2216 VTAIL.n597 VTAIL.n596 104.615
R2217 VTAIL.n596 VTAIL.n550 104.615
R2218 VTAIL.n589 VTAIL.n550 104.615
R2219 VTAIL.n589 VTAIL.n588 104.615
R2220 VTAIL.n588 VTAIL.n554 104.615
R2221 VTAIL.n581 VTAIL.n554 104.615
R2222 VTAIL.n581 VTAIL.n580 104.615
R2223 VTAIL.n580 VTAIL.n558 104.615
R2224 VTAIL.n573 VTAIL.n558 104.615
R2225 VTAIL.n573 VTAIL.n572 104.615
R2226 VTAIL.n572 VTAIL.n562 104.615
R2227 VTAIL.n565 VTAIL.n562 104.615
R2228 VTAIL.n524 VTAIL.n523 104.615
R2229 VTAIL.n523 VTAIL.n427 104.615
R2230 VTAIL.n516 VTAIL.n427 104.615
R2231 VTAIL.n516 VTAIL.n515 104.615
R2232 VTAIL.n515 VTAIL.n431 104.615
R2233 VTAIL.n508 VTAIL.n431 104.615
R2234 VTAIL.n508 VTAIL.n507 104.615
R2235 VTAIL.n507 VTAIL.n435 104.615
R2236 VTAIL.n439 VTAIL.n435 104.615
R2237 VTAIL.n499 VTAIL.n439 104.615
R2238 VTAIL.n499 VTAIL.n498 104.615
R2239 VTAIL.n498 VTAIL.n440 104.615
R2240 VTAIL.n491 VTAIL.n440 104.615
R2241 VTAIL.n491 VTAIL.n490 104.615
R2242 VTAIL.n490 VTAIL.n444 104.615
R2243 VTAIL.n483 VTAIL.n444 104.615
R2244 VTAIL.n483 VTAIL.n482 104.615
R2245 VTAIL.n482 VTAIL.n448 104.615
R2246 VTAIL.n475 VTAIL.n448 104.615
R2247 VTAIL.n475 VTAIL.n474 104.615
R2248 VTAIL.n474 VTAIL.n452 104.615
R2249 VTAIL.n467 VTAIL.n452 104.615
R2250 VTAIL.n467 VTAIL.n466 104.615
R2251 VTAIL.n466 VTAIL.n456 104.615
R2252 VTAIL.n459 VTAIL.n456 104.615
R2253 VTAIL.n418 VTAIL.n417 104.615
R2254 VTAIL.n417 VTAIL.n321 104.615
R2255 VTAIL.n410 VTAIL.n321 104.615
R2256 VTAIL.n410 VTAIL.n409 104.615
R2257 VTAIL.n409 VTAIL.n325 104.615
R2258 VTAIL.n402 VTAIL.n325 104.615
R2259 VTAIL.n402 VTAIL.n401 104.615
R2260 VTAIL.n401 VTAIL.n329 104.615
R2261 VTAIL.n333 VTAIL.n329 104.615
R2262 VTAIL.n393 VTAIL.n333 104.615
R2263 VTAIL.n393 VTAIL.n392 104.615
R2264 VTAIL.n392 VTAIL.n334 104.615
R2265 VTAIL.n385 VTAIL.n334 104.615
R2266 VTAIL.n385 VTAIL.n384 104.615
R2267 VTAIL.n384 VTAIL.n338 104.615
R2268 VTAIL.n377 VTAIL.n338 104.615
R2269 VTAIL.n377 VTAIL.n376 104.615
R2270 VTAIL.n376 VTAIL.n342 104.615
R2271 VTAIL.n369 VTAIL.n342 104.615
R2272 VTAIL.n369 VTAIL.n368 104.615
R2273 VTAIL.n368 VTAIL.n346 104.615
R2274 VTAIL.n361 VTAIL.n346 104.615
R2275 VTAIL.n361 VTAIL.n360 104.615
R2276 VTAIL.n360 VTAIL.n350 104.615
R2277 VTAIL.n353 VTAIL.n350 104.615
R2278 VTAIL.n776 VTAIL.t5 52.3082
R2279 VTAIL.n34 VTAIL.t4 52.3082
R2280 VTAIL.n140 VTAIL.t2 52.3082
R2281 VTAIL.n246 VTAIL.t0 52.3082
R2282 VTAIL.n671 VTAIL.t3 52.3082
R2283 VTAIL.n565 VTAIL.t1 52.3082
R2284 VTAIL.n459 VTAIL.t6 52.3082
R2285 VTAIL.n353 VTAIL.t7 52.3082
R2286 VTAIL.n847 VTAIL.n846 32.7672
R2287 VTAIL.n105 VTAIL.n104 32.7672
R2288 VTAIL.n211 VTAIL.n210 32.7672
R2289 VTAIL.n317 VTAIL.n316 32.7672
R2290 VTAIL.n741 VTAIL.n740 32.7672
R2291 VTAIL.n635 VTAIL.n634 32.7672
R2292 VTAIL.n529 VTAIL.n528 32.7672
R2293 VTAIL.n423 VTAIL.n422 32.7672
R2294 VTAIL.n847 VTAIL.n741 31.9186
R2295 VTAIL.n423 VTAIL.n317 31.9186
R2296 VTAIL.n777 VTAIL.n775 15.6677
R2297 VTAIL.n35 VTAIL.n33 15.6677
R2298 VTAIL.n141 VTAIL.n139 15.6677
R2299 VTAIL.n247 VTAIL.n245 15.6677
R2300 VTAIL.n672 VTAIL.n670 15.6677
R2301 VTAIL.n566 VTAIL.n564 15.6677
R2302 VTAIL.n460 VTAIL.n458 15.6677
R2303 VTAIL.n354 VTAIL.n352 15.6677
R2304 VTAIL.n824 VTAIL.n823 13.1884
R2305 VTAIL.n82 VTAIL.n81 13.1884
R2306 VTAIL.n188 VTAIL.n187 13.1884
R2307 VTAIL.n294 VTAIL.n293 13.1884
R2308 VTAIL.n718 VTAIL.n717 13.1884
R2309 VTAIL.n612 VTAIL.n611 13.1884
R2310 VTAIL.n506 VTAIL.n505 13.1884
R2311 VTAIL.n400 VTAIL.n399 13.1884
R2312 VTAIL.n778 VTAIL.n774 12.8005
R2313 VTAIL.n822 VTAIL.n754 12.8005
R2314 VTAIL.n827 VTAIL.n752 12.8005
R2315 VTAIL.n36 VTAIL.n32 12.8005
R2316 VTAIL.n80 VTAIL.n12 12.8005
R2317 VTAIL.n85 VTAIL.n10 12.8005
R2318 VTAIL.n142 VTAIL.n138 12.8005
R2319 VTAIL.n186 VTAIL.n118 12.8005
R2320 VTAIL.n191 VTAIL.n116 12.8005
R2321 VTAIL.n248 VTAIL.n244 12.8005
R2322 VTAIL.n292 VTAIL.n224 12.8005
R2323 VTAIL.n297 VTAIL.n222 12.8005
R2324 VTAIL.n721 VTAIL.n646 12.8005
R2325 VTAIL.n716 VTAIL.n648 12.8005
R2326 VTAIL.n673 VTAIL.n669 12.8005
R2327 VTAIL.n615 VTAIL.n540 12.8005
R2328 VTAIL.n610 VTAIL.n542 12.8005
R2329 VTAIL.n567 VTAIL.n563 12.8005
R2330 VTAIL.n509 VTAIL.n434 12.8005
R2331 VTAIL.n504 VTAIL.n436 12.8005
R2332 VTAIL.n461 VTAIL.n457 12.8005
R2333 VTAIL.n403 VTAIL.n328 12.8005
R2334 VTAIL.n398 VTAIL.n330 12.8005
R2335 VTAIL.n355 VTAIL.n351 12.8005
R2336 VTAIL.n782 VTAIL.n781 12.0247
R2337 VTAIL.n819 VTAIL.n818 12.0247
R2338 VTAIL.n828 VTAIL.n750 12.0247
R2339 VTAIL.n40 VTAIL.n39 12.0247
R2340 VTAIL.n77 VTAIL.n76 12.0247
R2341 VTAIL.n86 VTAIL.n8 12.0247
R2342 VTAIL.n146 VTAIL.n145 12.0247
R2343 VTAIL.n183 VTAIL.n182 12.0247
R2344 VTAIL.n192 VTAIL.n114 12.0247
R2345 VTAIL.n252 VTAIL.n251 12.0247
R2346 VTAIL.n289 VTAIL.n288 12.0247
R2347 VTAIL.n298 VTAIL.n220 12.0247
R2348 VTAIL.n722 VTAIL.n644 12.0247
R2349 VTAIL.n713 VTAIL.n712 12.0247
R2350 VTAIL.n677 VTAIL.n676 12.0247
R2351 VTAIL.n616 VTAIL.n538 12.0247
R2352 VTAIL.n607 VTAIL.n606 12.0247
R2353 VTAIL.n571 VTAIL.n570 12.0247
R2354 VTAIL.n510 VTAIL.n432 12.0247
R2355 VTAIL.n501 VTAIL.n500 12.0247
R2356 VTAIL.n465 VTAIL.n464 12.0247
R2357 VTAIL.n404 VTAIL.n326 12.0247
R2358 VTAIL.n395 VTAIL.n394 12.0247
R2359 VTAIL.n359 VTAIL.n358 12.0247
R2360 VTAIL.n785 VTAIL.n772 11.249
R2361 VTAIL.n814 VTAIL.n756 11.249
R2362 VTAIL.n832 VTAIL.n831 11.249
R2363 VTAIL.n43 VTAIL.n30 11.249
R2364 VTAIL.n72 VTAIL.n14 11.249
R2365 VTAIL.n90 VTAIL.n89 11.249
R2366 VTAIL.n149 VTAIL.n136 11.249
R2367 VTAIL.n178 VTAIL.n120 11.249
R2368 VTAIL.n196 VTAIL.n195 11.249
R2369 VTAIL.n255 VTAIL.n242 11.249
R2370 VTAIL.n284 VTAIL.n226 11.249
R2371 VTAIL.n302 VTAIL.n301 11.249
R2372 VTAIL.n726 VTAIL.n725 11.249
R2373 VTAIL.n709 VTAIL.n650 11.249
R2374 VTAIL.n680 VTAIL.n667 11.249
R2375 VTAIL.n620 VTAIL.n619 11.249
R2376 VTAIL.n603 VTAIL.n544 11.249
R2377 VTAIL.n574 VTAIL.n561 11.249
R2378 VTAIL.n514 VTAIL.n513 11.249
R2379 VTAIL.n497 VTAIL.n438 11.249
R2380 VTAIL.n468 VTAIL.n455 11.249
R2381 VTAIL.n408 VTAIL.n407 11.249
R2382 VTAIL.n391 VTAIL.n332 11.249
R2383 VTAIL.n362 VTAIL.n349 11.249
R2384 VTAIL.n786 VTAIL.n770 10.4732
R2385 VTAIL.n813 VTAIL.n758 10.4732
R2386 VTAIL.n835 VTAIL.n748 10.4732
R2387 VTAIL.n44 VTAIL.n28 10.4732
R2388 VTAIL.n71 VTAIL.n16 10.4732
R2389 VTAIL.n93 VTAIL.n6 10.4732
R2390 VTAIL.n150 VTAIL.n134 10.4732
R2391 VTAIL.n177 VTAIL.n122 10.4732
R2392 VTAIL.n199 VTAIL.n112 10.4732
R2393 VTAIL.n256 VTAIL.n240 10.4732
R2394 VTAIL.n283 VTAIL.n228 10.4732
R2395 VTAIL.n305 VTAIL.n218 10.4732
R2396 VTAIL.n729 VTAIL.n642 10.4732
R2397 VTAIL.n708 VTAIL.n653 10.4732
R2398 VTAIL.n681 VTAIL.n665 10.4732
R2399 VTAIL.n623 VTAIL.n536 10.4732
R2400 VTAIL.n602 VTAIL.n547 10.4732
R2401 VTAIL.n575 VTAIL.n559 10.4732
R2402 VTAIL.n517 VTAIL.n430 10.4732
R2403 VTAIL.n496 VTAIL.n441 10.4732
R2404 VTAIL.n469 VTAIL.n453 10.4732
R2405 VTAIL.n411 VTAIL.n324 10.4732
R2406 VTAIL.n390 VTAIL.n335 10.4732
R2407 VTAIL.n363 VTAIL.n347 10.4732
R2408 VTAIL.n790 VTAIL.n789 9.69747
R2409 VTAIL.n810 VTAIL.n809 9.69747
R2410 VTAIL.n836 VTAIL.n746 9.69747
R2411 VTAIL.n48 VTAIL.n47 9.69747
R2412 VTAIL.n68 VTAIL.n67 9.69747
R2413 VTAIL.n94 VTAIL.n4 9.69747
R2414 VTAIL.n154 VTAIL.n153 9.69747
R2415 VTAIL.n174 VTAIL.n173 9.69747
R2416 VTAIL.n200 VTAIL.n110 9.69747
R2417 VTAIL.n260 VTAIL.n259 9.69747
R2418 VTAIL.n280 VTAIL.n279 9.69747
R2419 VTAIL.n306 VTAIL.n216 9.69747
R2420 VTAIL.n730 VTAIL.n640 9.69747
R2421 VTAIL.n705 VTAIL.n704 9.69747
R2422 VTAIL.n685 VTAIL.n684 9.69747
R2423 VTAIL.n624 VTAIL.n534 9.69747
R2424 VTAIL.n599 VTAIL.n598 9.69747
R2425 VTAIL.n579 VTAIL.n578 9.69747
R2426 VTAIL.n518 VTAIL.n428 9.69747
R2427 VTAIL.n493 VTAIL.n492 9.69747
R2428 VTAIL.n473 VTAIL.n472 9.69747
R2429 VTAIL.n412 VTAIL.n322 9.69747
R2430 VTAIL.n387 VTAIL.n386 9.69747
R2431 VTAIL.n367 VTAIL.n366 9.69747
R2432 VTAIL.n846 VTAIL.n845 9.45567
R2433 VTAIL.n104 VTAIL.n103 9.45567
R2434 VTAIL.n210 VTAIL.n209 9.45567
R2435 VTAIL.n316 VTAIL.n315 9.45567
R2436 VTAIL.n740 VTAIL.n739 9.45567
R2437 VTAIL.n634 VTAIL.n633 9.45567
R2438 VTAIL.n528 VTAIL.n527 9.45567
R2439 VTAIL.n422 VTAIL.n421 9.45567
R2440 VTAIL.n744 VTAIL.n743 9.3005
R2441 VTAIL.n839 VTAIL.n838 9.3005
R2442 VTAIL.n837 VTAIL.n836 9.3005
R2443 VTAIL.n748 VTAIL.n747 9.3005
R2444 VTAIL.n831 VTAIL.n830 9.3005
R2445 VTAIL.n829 VTAIL.n828 9.3005
R2446 VTAIL.n752 VTAIL.n751 9.3005
R2447 VTAIL.n797 VTAIL.n796 9.3005
R2448 VTAIL.n795 VTAIL.n794 9.3005
R2449 VTAIL.n768 VTAIL.n767 9.3005
R2450 VTAIL.n789 VTAIL.n788 9.3005
R2451 VTAIL.n787 VTAIL.n786 9.3005
R2452 VTAIL.n772 VTAIL.n771 9.3005
R2453 VTAIL.n781 VTAIL.n780 9.3005
R2454 VTAIL.n779 VTAIL.n778 9.3005
R2455 VTAIL.n764 VTAIL.n763 9.3005
R2456 VTAIL.n803 VTAIL.n802 9.3005
R2457 VTAIL.n805 VTAIL.n804 9.3005
R2458 VTAIL.n760 VTAIL.n759 9.3005
R2459 VTAIL.n811 VTAIL.n810 9.3005
R2460 VTAIL.n813 VTAIL.n812 9.3005
R2461 VTAIL.n756 VTAIL.n755 9.3005
R2462 VTAIL.n820 VTAIL.n819 9.3005
R2463 VTAIL.n822 VTAIL.n821 9.3005
R2464 VTAIL.n845 VTAIL.n844 9.3005
R2465 VTAIL.n2 VTAIL.n1 9.3005
R2466 VTAIL.n97 VTAIL.n96 9.3005
R2467 VTAIL.n95 VTAIL.n94 9.3005
R2468 VTAIL.n6 VTAIL.n5 9.3005
R2469 VTAIL.n89 VTAIL.n88 9.3005
R2470 VTAIL.n87 VTAIL.n86 9.3005
R2471 VTAIL.n10 VTAIL.n9 9.3005
R2472 VTAIL.n55 VTAIL.n54 9.3005
R2473 VTAIL.n53 VTAIL.n52 9.3005
R2474 VTAIL.n26 VTAIL.n25 9.3005
R2475 VTAIL.n47 VTAIL.n46 9.3005
R2476 VTAIL.n45 VTAIL.n44 9.3005
R2477 VTAIL.n30 VTAIL.n29 9.3005
R2478 VTAIL.n39 VTAIL.n38 9.3005
R2479 VTAIL.n37 VTAIL.n36 9.3005
R2480 VTAIL.n22 VTAIL.n21 9.3005
R2481 VTAIL.n61 VTAIL.n60 9.3005
R2482 VTAIL.n63 VTAIL.n62 9.3005
R2483 VTAIL.n18 VTAIL.n17 9.3005
R2484 VTAIL.n69 VTAIL.n68 9.3005
R2485 VTAIL.n71 VTAIL.n70 9.3005
R2486 VTAIL.n14 VTAIL.n13 9.3005
R2487 VTAIL.n78 VTAIL.n77 9.3005
R2488 VTAIL.n80 VTAIL.n79 9.3005
R2489 VTAIL.n103 VTAIL.n102 9.3005
R2490 VTAIL.n108 VTAIL.n107 9.3005
R2491 VTAIL.n203 VTAIL.n202 9.3005
R2492 VTAIL.n201 VTAIL.n200 9.3005
R2493 VTAIL.n112 VTAIL.n111 9.3005
R2494 VTAIL.n195 VTAIL.n194 9.3005
R2495 VTAIL.n193 VTAIL.n192 9.3005
R2496 VTAIL.n116 VTAIL.n115 9.3005
R2497 VTAIL.n161 VTAIL.n160 9.3005
R2498 VTAIL.n159 VTAIL.n158 9.3005
R2499 VTAIL.n132 VTAIL.n131 9.3005
R2500 VTAIL.n153 VTAIL.n152 9.3005
R2501 VTAIL.n151 VTAIL.n150 9.3005
R2502 VTAIL.n136 VTAIL.n135 9.3005
R2503 VTAIL.n145 VTAIL.n144 9.3005
R2504 VTAIL.n143 VTAIL.n142 9.3005
R2505 VTAIL.n128 VTAIL.n127 9.3005
R2506 VTAIL.n167 VTAIL.n166 9.3005
R2507 VTAIL.n169 VTAIL.n168 9.3005
R2508 VTAIL.n124 VTAIL.n123 9.3005
R2509 VTAIL.n175 VTAIL.n174 9.3005
R2510 VTAIL.n177 VTAIL.n176 9.3005
R2511 VTAIL.n120 VTAIL.n119 9.3005
R2512 VTAIL.n184 VTAIL.n183 9.3005
R2513 VTAIL.n186 VTAIL.n185 9.3005
R2514 VTAIL.n209 VTAIL.n208 9.3005
R2515 VTAIL.n214 VTAIL.n213 9.3005
R2516 VTAIL.n309 VTAIL.n308 9.3005
R2517 VTAIL.n307 VTAIL.n306 9.3005
R2518 VTAIL.n218 VTAIL.n217 9.3005
R2519 VTAIL.n301 VTAIL.n300 9.3005
R2520 VTAIL.n299 VTAIL.n298 9.3005
R2521 VTAIL.n222 VTAIL.n221 9.3005
R2522 VTAIL.n267 VTAIL.n266 9.3005
R2523 VTAIL.n265 VTAIL.n264 9.3005
R2524 VTAIL.n238 VTAIL.n237 9.3005
R2525 VTAIL.n259 VTAIL.n258 9.3005
R2526 VTAIL.n257 VTAIL.n256 9.3005
R2527 VTAIL.n242 VTAIL.n241 9.3005
R2528 VTAIL.n251 VTAIL.n250 9.3005
R2529 VTAIL.n249 VTAIL.n248 9.3005
R2530 VTAIL.n234 VTAIL.n233 9.3005
R2531 VTAIL.n273 VTAIL.n272 9.3005
R2532 VTAIL.n275 VTAIL.n274 9.3005
R2533 VTAIL.n230 VTAIL.n229 9.3005
R2534 VTAIL.n281 VTAIL.n280 9.3005
R2535 VTAIL.n283 VTAIL.n282 9.3005
R2536 VTAIL.n226 VTAIL.n225 9.3005
R2537 VTAIL.n290 VTAIL.n289 9.3005
R2538 VTAIL.n292 VTAIL.n291 9.3005
R2539 VTAIL.n315 VTAIL.n314 9.3005
R2540 VTAIL.n698 VTAIL.n697 9.3005
R2541 VTAIL.n700 VTAIL.n699 9.3005
R2542 VTAIL.n655 VTAIL.n654 9.3005
R2543 VTAIL.n706 VTAIL.n705 9.3005
R2544 VTAIL.n708 VTAIL.n707 9.3005
R2545 VTAIL.n650 VTAIL.n649 9.3005
R2546 VTAIL.n714 VTAIL.n713 9.3005
R2547 VTAIL.n716 VTAIL.n715 9.3005
R2548 VTAIL.n739 VTAIL.n738 9.3005
R2549 VTAIL.n638 VTAIL.n637 9.3005
R2550 VTAIL.n733 VTAIL.n732 9.3005
R2551 VTAIL.n731 VTAIL.n730 9.3005
R2552 VTAIL.n642 VTAIL.n641 9.3005
R2553 VTAIL.n725 VTAIL.n724 9.3005
R2554 VTAIL.n723 VTAIL.n722 9.3005
R2555 VTAIL.n646 VTAIL.n645 9.3005
R2556 VTAIL.n659 VTAIL.n658 9.3005
R2557 VTAIL.n692 VTAIL.n691 9.3005
R2558 VTAIL.n690 VTAIL.n689 9.3005
R2559 VTAIL.n663 VTAIL.n662 9.3005
R2560 VTAIL.n684 VTAIL.n683 9.3005
R2561 VTAIL.n682 VTAIL.n681 9.3005
R2562 VTAIL.n667 VTAIL.n666 9.3005
R2563 VTAIL.n676 VTAIL.n675 9.3005
R2564 VTAIL.n674 VTAIL.n673 9.3005
R2565 VTAIL.n592 VTAIL.n591 9.3005
R2566 VTAIL.n594 VTAIL.n593 9.3005
R2567 VTAIL.n549 VTAIL.n548 9.3005
R2568 VTAIL.n600 VTAIL.n599 9.3005
R2569 VTAIL.n602 VTAIL.n601 9.3005
R2570 VTAIL.n544 VTAIL.n543 9.3005
R2571 VTAIL.n608 VTAIL.n607 9.3005
R2572 VTAIL.n610 VTAIL.n609 9.3005
R2573 VTAIL.n633 VTAIL.n632 9.3005
R2574 VTAIL.n532 VTAIL.n531 9.3005
R2575 VTAIL.n627 VTAIL.n626 9.3005
R2576 VTAIL.n625 VTAIL.n624 9.3005
R2577 VTAIL.n536 VTAIL.n535 9.3005
R2578 VTAIL.n619 VTAIL.n618 9.3005
R2579 VTAIL.n617 VTAIL.n616 9.3005
R2580 VTAIL.n540 VTAIL.n539 9.3005
R2581 VTAIL.n553 VTAIL.n552 9.3005
R2582 VTAIL.n586 VTAIL.n585 9.3005
R2583 VTAIL.n584 VTAIL.n583 9.3005
R2584 VTAIL.n557 VTAIL.n556 9.3005
R2585 VTAIL.n578 VTAIL.n577 9.3005
R2586 VTAIL.n576 VTAIL.n575 9.3005
R2587 VTAIL.n561 VTAIL.n560 9.3005
R2588 VTAIL.n570 VTAIL.n569 9.3005
R2589 VTAIL.n568 VTAIL.n567 9.3005
R2590 VTAIL.n486 VTAIL.n485 9.3005
R2591 VTAIL.n488 VTAIL.n487 9.3005
R2592 VTAIL.n443 VTAIL.n442 9.3005
R2593 VTAIL.n494 VTAIL.n493 9.3005
R2594 VTAIL.n496 VTAIL.n495 9.3005
R2595 VTAIL.n438 VTAIL.n437 9.3005
R2596 VTAIL.n502 VTAIL.n501 9.3005
R2597 VTAIL.n504 VTAIL.n503 9.3005
R2598 VTAIL.n527 VTAIL.n526 9.3005
R2599 VTAIL.n426 VTAIL.n425 9.3005
R2600 VTAIL.n521 VTAIL.n520 9.3005
R2601 VTAIL.n519 VTAIL.n518 9.3005
R2602 VTAIL.n430 VTAIL.n429 9.3005
R2603 VTAIL.n513 VTAIL.n512 9.3005
R2604 VTAIL.n511 VTAIL.n510 9.3005
R2605 VTAIL.n434 VTAIL.n433 9.3005
R2606 VTAIL.n447 VTAIL.n446 9.3005
R2607 VTAIL.n480 VTAIL.n479 9.3005
R2608 VTAIL.n478 VTAIL.n477 9.3005
R2609 VTAIL.n451 VTAIL.n450 9.3005
R2610 VTAIL.n472 VTAIL.n471 9.3005
R2611 VTAIL.n470 VTAIL.n469 9.3005
R2612 VTAIL.n455 VTAIL.n454 9.3005
R2613 VTAIL.n464 VTAIL.n463 9.3005
R2614 VTAIL.n462 VTAIL.n461 9.3005
R2615 VTAIL.n380 VTAIL.n379 9.3005
R2616 VTAIL.n382 VTAIL.n381 9.3005
R2617 VTAIL.n337 VTAIL.n336 9.3005
R2618 VTAIL.n388 VTAIL.n387 9.3005
R2619 VTAIL.n390 VTAIL.n389 9.3005
R2620 VTAIL.n332 VTAIL.n331 9.3005
R2621 VTAIL.n396 VTAIL.n395 9.3005
R2622 VTAIL.n398 VTAIL.n397 9.3005
R2623 VTAIL.n421 VTAIL.n420 9.3005
R2624 VTAIL.n320 VTAIL.n319 9.3005
R2625 VTAIL.n415 VTAIL.n414 9.3005
R2626 VTAIL.n413 VTAIL.n412 9.3005
R2627 VTAIL.n324 VTAIL.n323 9.3005
R2628 VTAIL.n407 VTAIL.n406 9.3005
R2629 VTAIL.n405 VTAIL.n404 9.3005
R2630 VTAIL.n328 VTAIL.n327 9.3005
R2631 VTAIL.n341 VTAIL.n340 9.3005
R2632 VTAIL.n374 VTAIL.n373 9.3005
R2633 VTAIL.n372 VTAIL.n371 9.3005
R2634 VTAIL.n345 VTAIL.n344 9.3005
R2635 VTAIL.n366 VTAIL.n365 9.3005
R2636 VTAIL.n364 VTAIL.n363 9.3005
R2637 VTAIL.n349 VTAIL.n348 9.3005
R2638 VTAIL.n358 VTAIL.n357 9.3005
R2639 VTAIL.n356 VTAIL.n355 9.3005
R2640 VTAIL.n793 VTAIL.n768 8.92171
R2641 VTAIL.n806 VTAIL.n760 8.92171
R2642 VTAIL.n840 VTAIL.n839 8.92171
R2643 VTAIL.n51 VTAIL.n26 8.92171
R2644 VTAIL.n64 VTAIL.n18 8.92171
R2645 VTAIL.n98 VTAIL.n97 8.92171
R2646 VTAIL.n157 VTAIL.n132 8.92171
R2647 VTAIL.n170 VTAIL.n124 8.92171
R2648 VTAIL.n204 VTAIL.n203 8.92171
R2649 VTAIL.n263 VTAIL.n238 8.92171
R2650 VTAIL.n276 VTAIL.n230 8.92171
R2651 VTAIL.n310 VTAIL.n309 8.92171
R2652 VTAIL.n734 VTAIL.n733 8.92171
R2653 VTAIL.n701 VTAIL.n655 8.92171
R2654 VTAIL.n688 VTAIL.n663 8.92171
R2655 VTAIL.n628 VTAIL.n627 8.92171
R2656 VTAIL.n595 VTAIL.n549 8.92171
R2657 VTAIL.n582 VTAIL.n557 8.92171
R2658 VTAIL.n522 VTAIL.n521 8.92171
R2659 VTAIL.n489 VTAIL.n443 8.92171
R2660 VTAIL.n476 VTAIL.n451 8.92171
R2661 VTAIL.n416 VTAIL.n415 8.92171
R2662 VTAIL.n383 VTAIL.n337 8.92171
R2663 VTAIL.n370 VTAIL.n345 8.92171
R2664 VTAIL.n794 VTAIL.n766 8.14595
R2665 VTAIL.n805 VTAIL.n762 8.14595
R2666 VTAIL.n843 VTAIL.n744 8.14595
R2667 VTAIL.n52 VTAIL.n24 8.14595
R2668 VTAIL.n63 VTAIL.n20 8.14595
R2669 VTAIL.n101 VTAIL.n2 8.14595
R2670 VTAIL.n158 VTAIL.n130 8.14595
R2671 VTAIL.n169 VTAIL.n126 8.14595
R2672 VTAIL.n207 VTAIL.n108 8.14595
R2673 VTAIL.n264 VTAIL.n236 8.14595
R2674 VTAIL.n275 VTAIL.n232 8.14595
R2675 VTAIL.n313 VTAIL.n214 8.14595
R2676 VTAIL.n737 VTAIL.n638 8.14595
R2677 VTAIL.n700 VTAIL.n657 8.14595
R2678 VTAIL.n689 VTAIL.n661 8.14595
R2679 VTAIL.n631 VTAIL.n532 8.14595
R2680 VTAIL.n594 VTAIL.n551 8.14595
R2681 VTAIL.n583 VTAIL.n555 8.14595
R2682 VTAIL.n525 VTAIL.n426 8.14595
R2683 VTAIL.n488 VTAIL.n445 8.14595
R2684 VTAIL.n477 VTAIL.n449 8.14595
R2685 VTAIL.n419 VTAIL.n320 8.14595
R2686 VTAIL.n382 VTAIL.n339 8.14595
R2687 VTAIL.n371 VTAIL.n343 8.14595
R2688 VTAIL.n798 VTAIL.n797 7.3702
R2689 VTAIL.n802 VTAIL.n801 7.3702
R2690 VTAIL.n844 VTAIL.n742 7.3702
R2691 VTAIL.n56 VTAIL.n55 7.3702
R2692 VTAIL.n60 VTAIL.n59 7.3702
R2693 VTAIL.n102 VTAIL.n0 7.3702
R2694 VTAIL.n162 VTAIL.n161 7.3702
R2695 VTAIL.n166 VTAIL.n165 7.3702
R2696 VTAIL.n208 VTAIL.n106 7.3702
R2697 VTAIL.n268 VTAIL.n267 7.3702
R2698 VTAIL.n272 VTAIL.n271 7.3702
R2699 VTAIL.n314 VTAIL.n212 7.3702
R2700 VTAIL.n738 VTAIL.n636 7.3702
R2701 VTAIL.n697 VTAIL.n696 7.3702
R2702 VTAIL.n693 VTAIL.n692 7.3702
R2703 VTAIL.n632 VTAIL.n530 7.3702
R2704 VTAIL.n591 VTAIL.n590 7.3702
R2705 VTAIL.n587 VTAIL.n586 7.3702
R2706 VTAIL.n526 VTAIL.n424 7.3702
R2707 VTAIL.n485 VTAIL.n484 7.3702
R2708 VTAIL.n481 VTAIL.n480 7.3702
R2709 VTAIL.n420 VTAIL.n318 7.3702
R2710 VTAIL.n379 VTAIL.n378 7.3702
R2711 VTAIL.n375 VTAIL.n374 7.3702
R2712 VTAIL.n798 VTAIL.n764 6.59444
R2713 VTAIL.n801 VTAIL.n764 6.59444
R2714 VTAIL.n846 VTAIL.n742 6.59444
R2715 VTAIL.n56 VTAIL.n22 6.59444
R2716 VTAIL.n59 VTAIL.n22 6.59444
R2717 VTAIL.n104 VTAIL.n0 6.59444
R2718 VTAIL.n162 VTAIL.n128 6.59444
R2719 VTAIL.n165 VTAIL.n128 6.59444
R2720 VTAIL.n210 VTAIL.n106 6.59444
R2721 VTAIL.n268 VTAIL.n234 6.59444
R2722 VTAIL.n271 VTAIL.n234 6.59444
R2723 VTAIL.n316 VTAIL.n212 6.59444
R2724 VTAIL.n740 VTAIL.n636 6.59444
R2725 VTAIL.n696 VTAIL.n659 6.59444
R2726 VTAIL.n693 VTAIL.n659 6.59444
R2727 VTAIL.n634 VTAIL.n530 6.59444
R2728 VTAIL.n590 VTAIL.n553 6.59444
R2729 VTAIL.n587 VTAIL.n553 6.59444
R2730 VTAIL.n528 VTAIL.n424 6.59444
R2731 VTAIL.n484 VTAIL.n447 6.59444
R2732 VTAIL.n481 VTAIL.n447 6.59444
R2733 VTAIL.n422 VTAIL.n318 6.59444
R2734 VTAIL.n378 VTAIL.n341 6.59444
R2735 VTAIL.n375 VTAIL.n341 6.59444
R2736 VTAIL.n797 VTAIL.n766 5.81868
R2737 VTAIL.n802 VTAIL.n762 5.81868
R2738 VTAIL.n844 VTAIL.n843 5.81868
R2739 VTAIL.n55 VTAIL.n24 5.81868
R2740 VTAIL.n60 VTAIL.n20 5.81868
R2741 VTAIL.n102 VTAIL.n101 5.81868
R2742 VTAIL.n161 VTAIL.n130 5.81868
R2743 VTAIL.n166 VTAIL.n126 5.81868
R2744 VTAIL.n208 VTAIL.n207 5.81868
R2745 VTAIL.n267 VTAIL.n236 5.81868
R2746 VTAIL.n272 VTAIL.n232 5.81868
R2747 VTAIL.n314 VTAIL.n313 5.81868
R2748 VTAIL.n738 VTAIL.n737 5.81868
R2749 VTAIL.n697 VTAIL.n657 5.81868
R2750 VTAIL.n692 VTAIL.n661 5.81868
R2751 VTAIL.n632 VTAIL.n631 5.81868
R2752 VTAIL.n591 VTAIL.n551 5.81868
R2753 VTAIL.n586 VTAIL.n555 5.81868
R2754 VTAIL.n526 VTAIL.n525 5.81868
R2755 VTAIL.n485 VTAIL.n445 5.81868
R2756 VTAIL.n480 VTAIL.n449 5.81868
R2757 VTAIL.n420 VTAIL.n419 5.81868
R2758 VTAIL.n379 VTAIL.n339 5.81868
R2759 VTAIL.n374 VTAIL.n343 5.81868
R2760 VTAIL.n794 VTAIL.n793 5.04292
R2761 VTAIL.n806 VTAIL.n805 5.04292
R2762 VTAIL.n840 VTAIL.n744 5.04292
R2763 VTAIL.n52 VTAIL.n51 5.04292
R2764 VTAIL.n64 VTAIL.n63 5.04292
R2765 VTAIL.n98 VTAIL.n2 5.04292
R2766 VTAIL.n158 VTAIL.n157 5.04292
R2767 VTAIL.n170 VTAIL.n169 5.04292
R2768 VTAIL.n204 VTAIL.n108 5.04292
R2769 VTAIL.n264 VTAIL.n263 5.04292
R2770 VTAIL.n276 VTAIL.n275 5.04292
R2771 VTAIL.n310 VTAIL.n214 5.04292
R2772 VTAIL.n734 VTAIL.n638 5.04292
R2773 VTAIL.n701 VTAIL.n700 5.04292
R2774 VTAIL.n689 VTAIL.n688 5.04292
R2775 VTAIL.n628 VTAIL.n532 5.04292
R2776 VTAIL.n595 VTAIL.n594 5.04292
R2777 VTAIL.n583 VTAIL.n582 5.04292
R2778 VTAIL.n522 VTAIL.n426 5.04292
R2779 VTAIL.n489 VTAIL.n488 5.04292
R2780 VTAIL.n477 VTAIL.n476 5.04292
R2781 VTAIL.n416 VTAIL.n320 5.04292
R2782 VTAIL.n383 VTAIL.n382 5.04292
R2783 VTAIL.n371 VTAIL.n370 5.04292
R2784 VTAIL.n674 VTAIL.n670 4.38563
R2785 VTAIL.n568 VTAIL.n564 4.38563
R2786 VTAIL.n462 VTAIL.n458 4.38563
R2787 VTAIL.n356 VTAIL.n352 4.38563
R2788 VTAIL.n779 VTAIL.n775 4.38563
R2789 VTAIL.n37 VTAIL.n33 4.38563
R2790 VTAIL.n143 VTAIL.n139 4.38563
R2791 VTAIL.n249 VTAIL.n245 4.38563
R2792 VTAIL.n790 VTAIL.n768 4.26717
R2793 VTAIL.n809 VTAIL.n760 4.26717
R2794 VTAIL.n839 VTAIL.n746 4.26717
R2795 VTAIL.n48 VTAIL.n26 4.26717
R2796 VTAIL.n67 VTAIL.n18 4.26717
R2797 VTAIL.n97 VTAIL.n4 4.26717
R2798 VTAIL.n154 VTAIL.n132 4.26717
R2799 VTAIL.n173 VTAIL.n124 4.26717
R2800 VTAIL.n203 VTAIL.n110 4.26717
R2801 VTAIL.n260 VTAIL.n238 4.26717
R2802 VTAIL.n279 VTAIL.n230 4.26717
R2803 VTAIL.n309 VTAIL.n216 4.26717
R2804 VTAIL.n733 VTAIL.n640 4.26717
R2805 VTAIL.n704 VTAIL.n655 4.26717
R2806 VTAIL.n685 VTAIL.n663 4.26717
R2807 VTAIL.n627 VTAIL.n534 4.26717
R2808 VTAIL.n598 VTAIL.n549 4.26717
R2809 VTAIL.n579 VTAIL.n557 4.26717
R2810 VTAIL.n521 VTAIL.n428 4.26717
R2811 VTAIL.n492 VTAIL.n443 4.26717
R2812 VTAIL.n473 VTAIL.n451 4.26717
R2813 VTAIL.n415 VTAIL.n322 4.26717
R2814 VTAIL.n386 VTAIL.n337 4.26717
R2815 VTAIL.n367 VTAIL.n345 4.26717
R2816 VTAIL.n789 VTAIL.n770 3.49141
R2817 VTAIL.n810 VTAIL.n758 3.49141
R2818 VTAIL.n836 VTAIL.n835 3.49141
R2819 VTAIL.n47 VTAIL.n28 3.49141
R2820 VTAIL.n68 VTAIL.n16 3.49141
R2821 VTAIL.n94 VTAIL.n93 3.49141
R2822 VTAIL.n153 VTAIL.n134 3.49141
R2823 VTAIL.n174 VTAIL.n122 3.49141
R2824 VTAIL.n200 VTAIL.n199 3.49141
R2825 VTAIL.n259 VTAIL.n240 3.49141
R2826 VTAIL.n280 VTAIL.n228 3.49141
R2827 VTAIL.n306 VTAIL.n305 3.49141
R2828 VTAIL.n730 VTAIL.n729 3.49141
R2829 VTAIL.n705 VTAIL.n653 3.49141
R2830 VTAIL.n684 VTAIL.n665 3.49141
R2831 VTAIL.n624 VTAIL.n623 3.49141
R2832 VTAIL.n599 VTAIL.n547 3.49141
R2833 VTAIL.n578 VTAIL.n559 3.49141
R2834 VTAIL.n518 VTAIL.n517 3.49141
R2835 VTAIL.n493 VTAIL.n441 3.49141
R2836 VTAIL.n472 VTAIL.n453 3.49141
R2837 VTAIL.n412 VTAIL.n411 3.49141
R2838 VTAIL.n387 VTAIL.n335 3.49141
R2839 VTAIL.n366 VTAIL.n347 3.49141
R2840 VTAIL.n529 VTAIL.n423 3.18153
R2841 VTAIL.n741 VTAIL.n635 3.18153
R2842 VTAIL.n317 VTAIL.n211 3.18153
R2843 VTAIL.n786 VTAIL.n785 2.71565
R2844 VTAIL.n814 VTAIL.n813 2.71565
R2845 VTAIL.n832 VTAIL.n748 2.71565
R2846 VTAIL.n44 VTAIL.n43 2.71565
R2847 VTAIL.n72 VTAIL.n71 2.71565
R2848 VTAIL.n90 VTAIL.n6 2.71565
R2849 VTAIL.n150 VTAIL.n149 2.71565
R2850 VTAIL.n178 VTAIL.n177 2.71565
R2851 VTAIL.n196 VTAIL.n112 2.71565
R2852 VTAIL.n256 VTAIL.n255 2.71565
R2853 VTAIL.n284 VTAIL.n283 2.71565
R2854 VTAIL.n302 VTAIL.n218 2.71565
R2855 VTAIL.n726 VTAIL.n642 2.71565
R2856 VTAIL.n709 VTAIL.n708 2.71565
R2857 VTAIL.n681 VTAIL.n680 2.71565
R2858 VTAIL.n620 VTAIL.n536 2.71565
R2859 VTAIL.n603 VTAIL.n602 2.71565
R2860 VTAIL.n575 VTAIL.n574 2.71565
R2861 VTAIL.n514 VTAIL.n430 2.71565
R2862 VTAIL.n497 VTAIL.n496 2.71565
R2863 VTAIL.n469 VTAIL.n468 2.71565
R2864 VTAIL.n408 VTAIL.n324 2.71565
R2865 VTAIL.n391 VTAIL.n390 2.71565
R2866 VTAIL.n363 VTAIL.n362 2.71565
R2867 VTAIL.n782 VTAIL.n772 1.93989
R2868 VTAIL.n818 VTAIL.n756 1.93989
R2869 VTAIL.n831 VTAIL.n750 1.93989
R2870 VTAIL.n40 VTAIL.n30 1.93989
R2871 VTAIL.n76 VTAIL.n14 1.93989
R2872 VTAIL.n89 VTAIL.n8 1.93989
R2873 VTAIL.n146 VTAIL.n136 1.93989
R2874 VTAIL.n182 VTAIL.n120 1.93989
R2875 VTAIL.n195 VTAIL.n114 1.93989
R2876 VTAIL.n252 VTAIL.n242 1.93989
R2877 VTAIL.n288 VTAIL.n226 1.93989
R2878 VTAIL.n301 VTAIL.n220 1.93989
R2879 VTAIL.n725 VTAIL.n644 1.93989
R2880 VTAIL.n712 VTAIL.n650 1.93989
R2881 VTAIL.n677 VTAIL.n667 1.93989
R2882 VTAIL.n619 VTAIL.n538 1.93989
R2883 VTAIL.n606 VTAIL.n544 1.93989
R2884 VTAIL.n571 VTAIL.n561 1.93989
R2885 VTAIL.n513 VTAIL.n432 1.93989
R2886 VTAIL.n500 VTAIL.n438 1.93989
R2887 VTAIL.n465 VTAIL.n455 1.93989
R2888 VTAIL.n407 VTAIL.n326 1.93989
R2889 VTAIL.n394 VTAIL.n332 1.93989
R2890 VTAIL.n359 VTAIL.n349 1.93989
R2891 VTAIL VTAIL.n105 1.64921
R2892 VTAIL VTAIL.n847 1.53283
R2893 VTAIL.n781 VTAIL.n774 1.16414
R2894 VTAIL.n819 VTAIL.n754 1.16414
R2895 VTAIL.n828 VTAIL.n827 1.16414
R2896 VTAIL.n39 VTAIL.n32 1.16414
R2897 VTAIL.n77 VTAIL.n12 1.16414
R2898 VTAIL.n86 VTAIL.n85 1.16414
R2899 VTAIL.n145 VTAIL.n138 1.16414
R2900 VTAIL.n183 VTAIL.n118 1.16414
R2901 VTAIL.n192 VTAIL.n191 1.16414
R2902 VTAIL.n251 VTAIL.n244 1.16414
R2903 VTAIL.n289 VTAIL.n224 1.16414
R2904 VTAIL.n298 VTAIL.n297 1.16414
R2905 VTAIL.n722 VTAIL.n721 1.16414
R2906 VTAIL.n713 VTAIL.n648 1.16414
R2907 VTAIL.n676 VTAIL.n669 1.16414
R2908 VTAIL.n616 VTAIL.n615 1.16414
R2909 VTAIL.n607 VTAIL.n542 1.16414
R2910 VTAIL.n570 VTAIL.n563 1.16414
R2911 VTAIL.n510 VTAIL.n509 1.16414
R2912 VTAIL.n501 VTAIL.n436 1.16414
R2913 VTAIL.n464 VTAIL.n457 1.16414
R2914 VTAIL.n404 VTAIL.n403 1.16414
R2915 VTAIL.n395 VTAIL.n330 1.16414
R2916 VTAIL.n358 VTAIL.n351 1.16414
R2917 VTAIL.n635 VTAIL.n529 0.470328
R2918 VTAIL.n211 VTAIL.n105 0.470328
R2919 VTAIL.n778 VTAIL.n777 0.388379
R2920 VTAIL.n823 VTAIL.n822 0.388379
R2921 VTAIL.n824 VTAIL.n752 0.388379
R2922 VTAIL.n36 VTAIL.n35 0.388379
R2923 VTAIL.n81 VTAIL.n80 0.388379
R2924 VTAIL.n82 VTAIL.n10 0.388379
R2925 VTAIL.n142 VTAIL.n141 0.388379
R2926 VTAIL.n187 VTAIL.n186 0.388379
R2927 VTAIL.n188 VTAIL.n116 0.388379
R2928 VTAIL.n248 VTAIL.n247 0.388379
R2929 VTAIL.n293 VTAIL.n292 0.388379
R2930 VTAIL.n294 VTAIL.n222 0.388379
R2931 VTAIL.n718 VTAIL.n646 0.388379
R2932 VTAIL.n717 VTAIL.n716 0.388379
R2933 VTAIL.n673 VTAIL.n672 0.388379
R2934 VTAIL.n612 VTAIL.n540 0.388379
R2935 VTAIL.n611 VTAIL.n610 0.388379
R2936 VTAIL.n567 VTAIL.n566 0.388379
R2937 VTAIL.n506 VTAIL.n434 0.388379
R2938 VTAIL.n505 VTAIL.n504 0.388379
R2939 VTAIL.n461 VTAIL.n460 0.388379
R2940 VTAIL.n400 VTAIL.n328 0.388379
R2941 VTAIL.n399 VTAIL.n398 0.388379
R2942 VTAIL.n355 VTAIL.n354 0.388379
R2943 VTAIL.n780 VTAIL.n779 0.155672
R2944 VTAIL.n780 VTAIL.n771 0.155672
R2945 VTAIL.n787 VTAIL.n771 0.155672
R2946 VTAIL.n788 VTAIL.n787 0.155672
R2947 VTAIL.n788 VTAIL.n767 0.155672
R2948 VTAIL.n795 VTAIL.n767 0.155672
R2949 VTAIL.n796 VTAIL.n795 0.155672
R2950 VTAIL.n796 VTAIL.n763 0.155672
R2951 VTAIL.n803 VTAIL.n763 0.155672
R2952 VTAIL.n804 VTAIL.n803 0.155672
R2953 VTAIL.n804 VTAIL.n759 0.155672
R2954 VTAIL.n811 VTAIL.n759 0.155672
R2955 VTAIL.n812 VTAIL.n811 0.155672
R2956 VTAIL.n812 VTAIL.n755 0.155672
R2957 VTAIL.n820 VTAIL.n755 0.155672
R2958 VTAIL.n821 VTAIL.n820 0.155672
R2959 VTAIL.n821 VTAIL.n751 0.155672
R2960 VTAIL.n829 VTAIL.n751 0.155672
R2961 VTAIL.n830 VTAIL.n829 0.155672
R2962 VTAIL.n830 VTAIL.n747 0.155672
R2963 VTAIL.n837 VTAIL.n747 0.155672
R2964 VTAIL.n838 VTAIL.n837 0.155672
R2965 VTAIL.n838 VTAIL.n743 0.155672
R2966 VTAIL.n845 VTAIL.n743 0.155672
R2967 VTAIL.n38 VTAIL.n37 0.155672
R2968 VTAIL.n38 VTAIL.n29 0.155672
R2969 VTAIL.n45 VTAIL.n29 0.155672
R2970 VTAIL.n46 VTAIL.n45 0.155672
R2971 VTAIL.n46 VTAIL.n25 0.155672
R2972 VTAIL.n53 VTAIL.n25 0.155672
R2973 VTAIL.n54 VTAIL.n53 0.155672
R2974 VTAIL.n54 VTAIL.n21 0.155672
R2975 VTAIL.n61 VTAIL.n21 0.155672
R2976 VTAIL.n62 VTAIL.n61 0.155672
R2977 VTAIL.n62 VTAIL.n17 0.155672
R2978 VTAIL.n69 VTAIL.n17 0.155672
R2979 VTAIL.n70 VTAIL.n69 0.155672
R2980 VTAIL.n70 VTAIL.n13 0.155672
R2981 VTAIL.n78 VTAIL.n13 0.155672
R2982 VTAIL.n79 VTAIL.n78 0.155672
R2983 VTAIL.n79 VTAIL.n9 0.155672
R2984 VTAIL.n87 VTAIL.n9 0.155672
R2985 VTAIL.n88 VTAIL.n87 0.155672
R2986 VTAIL.n88 VTAIL.n5 0.155672
R2987 VTAIL.n95 VTAIL.n5 0.155672
R2988 VTAIL.n96 VTAIL.n95 0.155672
R2989 VTAIL.n96 VTAIL.n1 0.155672
R2990 VTAIL.n103 VTAIL.n1 0.155672
R2991 VTAIL.n144 VTAIL.n143 0.155672
R2992 VTAIL.n144 VTAIL.n135 0.155672
R2993 VTAIL.n151 VTAIL.n135 0.155672
R2994 VTAIL.n152 VTAIL.n151 0.155672
R2995 VTAIL.n152 VTAIL.n131 0.155672
R2996 VTAIL.n159 VTAIL.n131 0.155672
R2997 VTAIL.n160 VTAIL.n159 0.155672
R2998 VTAIL.n160 VTAIL.n127 0.155672
R2999 VTAIL.n167 VTAIL.n127 0.155672
R3000 VTAIL.n168 VTAIL.n167 0.155672
R3001 VTAIL.n168 VTAIL.n123 0.155672
R3002 VTAIL.n175 VTAIL.n123 0.155672
R3003 VTAIL.n176 VTAIL.n175 0.155672
R3004 VTAIL.n176 VTAIL.n119 0.155672
R3005 VTAIL.n184 VTAIL.n119 0.155672
R3006 VTAIL.n185 VTAIL.n184 0.155672
R3007 VTAIL.n185 VTAIL.n115 0.155672
R3008 VTAIL.n193 VTAIL.n115 0.155672
R3009 VTAIL.n194 VTAIL.n193 0.155672
R3010 VTAIL.n194 VTAIL.n111 0.155672
R3011 VTAIL.n201 VTAIL.n111 0.155672
R3012 VTAIL.n202 VTAIL.n201 0.155672
R3013 VTAIL.n202 VTAIL.n107 0.155672
R3014 VTAIL.n209 VTAIL.n107 0.155672
R3015 VTAIL.n250 VTAIL.n249 0.155672
R3016 VTAIL.n250 VTAIL.n241 0.155672
R3017 VTAIL.n257 VTAIL.n241 0.155672
R3018 VTAIL.n258 VTAIL.n257 0.155672
R3019 VTAIL.n258 VTAIL.n237 0.155672
R3020 VTAIL.n265 VTAIL.n237 0.155672
R3021 VTAIL.n266 VTAIL.n265 0.155672
R3022 VTAIL.n266 VTAIL.n233 0.155672
R3023 VTAIL.n273 VTAIL.n233 0.155672
R3024 VTAIL.n274 VTAIL.n273 0.155672
R3025 VTAIL.n274 VTAIL.n229 0.155672
R3026 VTAIL.n281 VTAIL.n229 0.155672
R3027 VTAIL.n282 VTAIL.n281 0.155672
R3028 VTAIL.n282 VTAIL.n225 0.155672
R3029 VTAIL.n290 VTAIL.n225 0.155672
R3030 VTAIL.n291 VTAIL.n290 0.155672
R3031 VTAIL.n291 VTAIL.n221 0.155672
R3032 VTAIL.n299 VTAIL.n221 0.155672
R3033 VTAIL.n300 VTAIL.n299 0.155672
R3034 VTAIL.n300 VTAIL.n217 0.155672
R3035 VTAIL.n307 VTAIL.n217 0.155672
R3036 VTAIL.n308 VTAIL.n307 0.155672
R3037 VTAIL.n308 VTAIL.n213 0.155672
R3038 VTAIL.n315 VTAIL.n213 0.155672
R3039 VTAIL.n739 VTAIL.n637 0.155672
R3040 VTAIL.n732 VTAIL.n637 0.155672
R3041 VTAIL.n732 VTAIL.n731 0.155672
R3042 VTAIL.n731 VTAIL.n641 0.155672
R3043 VTAIL.n724 VTAIL.n641 0.155672
R3044 VTAIL.n724 VTAIL.n723 0.155672
R3045 VTAIL.n723 VTAIL.n645 0.155672
R3046 VTAIL.n715 VTAIL.n645 0.155672
R3047 VTAIL.n715 VTAIL.n714 0.155672
R3048 VTAIL.n714 VTAIL.n649 0.155672
R3049 VTAIL.n707 VTAIL.n649 0.155672
R3050 VTAIL.n707 VTAIL.n706 0.155672
R3051 VTAIL.n706 VTAIL.n654 0.155672
R3052 VTAIL.n699 VTAIL.n654 0.155672
R3053 VTAIL.n699 VTAIL.n698 0.155672
R3054 VTAIL.n698 VTAIL.n658 0.155672
R3055 VTAIL.n691 VTAIL.n658 0.155672
R3056 VTAIL.n691 VTAIL.n690 0.155672
R3057 VTAIL.n690 VTAIL.n662 0.155672
R3058 VTAIL.n683 VTAIL.n662 0.155672
R3059 VTAIL.n683 VTAIL.n682 0.155672
R3060 VTAIL.n682 VTAIL.n666 0.155672
R3061 VTAIL.n675 VTAIL.n666 0.155672
R3062 VTAIL.n675 VTAIL.n674 0.155672
R3063 VTAIL.n633 VTAIL.n531 0.155672
R3064 VTAIL.n626 VTAIL.n531 0.155672
R3065 VTAIL.n626 VTAIL.n625 0.155672
R3066 VTAIL.n625 VTAIL.n535 0.155672
R3067 VTAIL.n618 VTAIL.n535 0.155672
R3068 VTAIL.n618 VTAIL.n617 0.155672
R3069 VTAIL.n617 VTAIL.n539 0.155672
R3070 VTAIL.n609 VTAIL.n539 0.155672
R3071 VTAIL.n609 VTAIL.n608 0.155672
R3072 VTAIL.n608 VTAIL.n543 0.155672
R3073 VTAIL.n601 VTAIL.n543 0.155672
R3074 VTAIL.n601 VTAIL.n600 0.155672
R3075 VTAIL.n600 VTAIL.n548 0.155672
R3076 VTAIL.n593 VTAIL.n548 0.155672
R3077 VTAIL.n593 VTAIL.n592 0.155672
R3078 VTAIL.n592 VTAIL.n552 0.155672
R3079 VTAIL.n585 VTAIL.n552 0.155672
R3080 VTAIL.n585 VTAIL.n584 0.155672
R3081 VTAIL.n584 VTAIL.n556 0.155672
R3082 VTAIL.n577 VTAIL.n556 0.155672
R3083 VTAIL.n577 VTAIL.n576 0.155672
R3084 VTAIL.n576 VTAIL.n560 0.155672
R3085 VTAIL.n569 VTAIL.n560 0.155672
R3086 VTAIL.n569 VTAIL.n568 0.155672
R3087 VTAIL.n527 VTAIL.n425 0.155672
R3088 VTAIL.n520 VTAIL.n425 0.155672
R3089 VTAIL.n520 VTAIL.n519 0.155672
R3090 VTAIL.n519 VTAIL.n429 0.155672
R3091 VTAIL.n512 VTAIL.n429 0.155672
R3092 VTAIL.n512 VTAIL.n511 0.155672
R3093 VTAIL.n511 VTAIL.n433 0.155672
R3094 VTAIL.n503 VTAIL.n433 0.155672
R3095 VTAIL.n503 VTAIL.n502 0.155672
R3096 VTAIL.n502 VTAIL.n437 0.155672
R3097 VTAIL.n495 VTAIL.n437 0.155672
R3098 VTAIL.n495 VTAIL.n494 0.155672
R3099 VTAIL.n494 VTAIL.n442 0.155672
R3100 VTAIL.n487 VTAIL.n442 0.155672
R3101 VTAIL.n487 VTAIL.n486 0.155672
R3102 VTAIL.n486 VTAIL.n446 0.155672
R3103 VTAIL.n479 VTAIL.n446 0.155672
R3104 VTAIL.n479 VTAIL.n478 0.155672
R3105 VTAIL.n478 VTAIL.n450 0.155672
R3106 VTAIL.n471 VTAIL.n450 0.155672
R3107 VTAIL.n471 VTAIL.n470 0.155672
R3108 VTAIL.n470 VTAIL.n454 0.155672
R3109 VTAIL.n463 VTAIL.n454 0.155672
R3110 VTAIL.n463 VTAIL.n462 0.155672
R3111 VTAIL.n421 VTAIL.n319 0.155672
R3112 VTAIL.n414 VTAIL.n319 0.155672
R3113 VTAIL.n414 VTAIL.n413 0.155672
R3114 VTAIL.n413 VTAIL.n323 0.155672
R3115 VTAIL.n406 VTAIL.n323 0.155672
R3116 VTAIL.n406 VTAIL.n405 0.155672
R3117 VTAIL.n405 VTAIL.n327 0.155672
R3118 VTAIL.n397 VTAIL.n327 0.155672
R3119 VTAIL.n397 VTAIL.n396 0.155672
R3120 VTAIL.n396 VTAIL.n331 0.155672
R3121 VTAIL.n389 VTAIL.n331 0.155672
R3122 VTAIL.n389 VTAIL.n388 0.155672
R3123 VTAIL.n388 VTAIL.n336 0.155672
R3124 VTAIL.n381 VTAIL.n336 0.155672
R3125 VTAIL.n381 VTAIL.n380 0.155672
R3126 VTAIL.n380 VTAIL.n340 0.155672
R3127 VTAIL.n373 VTAIL.n340 0.155672
R3128 VTAIL.n373 VTAIL.n372 0.155672
R3129 VTAIL.n372 VTAIL.n344 0.155672
R3130 VTAIL.n365 VTAIL.n344 0.155672
R3131 VTAIL.n365 VTAIL.n364 0.155672
R3132 VTAIL.n364 VTAIL.n348 0.155672
R3133 VTAIL.n357 VTAIL.n348 0.155672
R3134 VTAIL.n357 VTAIL.n356 0.155672
R3135 VP.n5 VP.t0 171.273
R3136 VP.n5 VP.t3 170.139
R3137 VP.n17 VP.n16 161.3
R3138 VP.n15 VP.n1 161.3
R3139 VP.n14 VP.n13 161.3
R3140 VP.n12 VP.n2 161.3
R3141 VP.n11 VP.n10 161.3
R3142 VP.n9 VP.n3 161.3
R3143 VP.n8 VP.n7 161.3
R3144 VP.n4 VP.t2 136.208
R3145 VP.n0 VP.t1 136.208
R3146 VP.n6 VP.n4 73.1852
R3147 VP.n18 VP.n0 73.1852
R3148 VP.n6 VP.n5 56.4575
R3149 VP.n10 VP.n2 40.4934
R3150 VP.n14 VP.n2 40.4934
R3151 VP.n9 VP.n8 24.4675
R3152 VP.n10 VP.n9 24.4675
R3153 VP.n15 VP.n14 24.4675
R3154 VP.n16 VP.n15 24.4675
R3155 VP.n8 VP.n4 16.8827
R3156 VP.n16 VP.n0 16.8827
R3157 VP.n7 VP.n6 0.354971
R3158 VP.n18 VP.n17 0.354971
R3159 VP VP.n18 0.26696
R3160 VP.n7 VP.n3 0.189894
R3161 VP.n11 VP.n3 0.189894
R3162 VP.n12 VP.n11 0.189894
R3163 VP.n13 VP.n12 0.189894
R3164 VP.n13 VP.n1 0.189894
R3165 VP.n17 VP.n1 0.189894
R3166 VDD1 VDD1.n1 111.358
R3167 VDD1 VDD1.n0 61.2618
R3168 VDD1.n0 VDD1.t3 1.04315
R3169 VDD1.n0 VDD1.t0 1.04315
R3170 VDD1.n1 VDD1.t1 1.04315
R3171 VDD1.n1 VDD1.t2 1.04315
C0 VDD1 VDD2 1.20298f
C1 VDD1 VN 0.149534f
C2 VDD2 VN 7.64913f
C3 VDD1 VTAIL 7.1089f
C4 VDD2 VTAIL 7.1682f
C5 VN VTAIL 7.34273f
C6 VP VDD1 7.94117f
C7 VP VDD2 0.442513f
C8 VP VN 8.03145f
C9 VP VTAIL 7.35683f
C10 VDD2 B 4.744762f
C11 VDD1 B 9.83364f
C12 VTAIL B 14.737252f
C13 VN B 12.69946f
C14 VP B 11.026055f
C15 VDD1.t3 B 0.40139f
C16 VDD1.t0 B 0.40139f
C17 VDD1.n0 B 3.66508f
C18 VDD1.t1 B 0.40139f
C19 VDD1.t2 B 0.40139f
C20 VDD1.n1 B 4.67755f
C21 VP.t1 B 3.59437f
C22 VP.n0 B 1.3232f
C23 VP.n1 B 0.02046f
C24 VP.n2 B 0.01654f
C25 VP.n3 B 0.02046f
C26 VP.t2 B 3.59437f
C27 VP.n4 B 1.3232f
C28 VP.t0 B 3.88022f
C29 VP.t3 B 3.87134f
C30 VP.n5 B 3.83362f
C31 VP.n6 B 1.37959f
C32 VP.n7 B 0.033022f
C33 VP.n8 B 0.032295f
C34 VP.n9 B 0.038132f
C35 VP.n10 B 0.040664f
C36 VP.n11 B 0.02046f
C37 VP.n12 B 0.02046f
C38 VP.n13 B 0.02046f
C39 VP.n14 B 0.040664f
C40 VP.n15 B 0.038132f
C41 VP.n16 B 0.032295f
C42 VP.n17 B 0.033022f
C43 VP.n18 B 0.048072f
C44 VTAIL.n0 B 0.022487f
C45 VTAIL.n1 B 0.015478f
C46 VTAIL.n2 B 0.008317f
C47 VTAIL.n3 B 0.019659f
C48 VTAIL.n4 B 0.008807f
C49 VTAIL.n5 B 0.015478f
C50 VTAIL.n6 B 0.008317f
C51 VTAIL.n7 B 0.019659f
C52 VTAIL.n8 B 0.008807f
C53 VTAIL.n9 B 0.015478f
C54 VTAIL.n10 B 0.008317f
C55 VTAIL.n11 B 0.019659f
C56 VTAIL.n12 B 0.008807f
C57 VTAIL.n13 B 0.015478f
C58 VTAIL.n14 B 0.008317f
C59 VTAIL.n15 B 0.019659f
C60 VTAIL.n16 B 0.008807f
C61 VTAIL.n17 B 0.015478f
C62 VTAIL.n18 B 0.008317f
C63 VTAIL.n19 B 0.019659f
C64 VTAIL.n20 B 0.008807f
C65 VTAIL.n21 B 0.015478f
C66 VTAIL.n22 B 0.008317f
C67 VTAIL.n23 B 0.019659f
C68 VTAIL.n24 B 0.008807f
C69 VTAIL.n25 B 0.015478f
C70 VTAIL.n26 B 0.008317f
C71 VTAIL.n27 B 0.019659f
C72 VTAIL.n28 B 0.008807f
C73 VTAIL.n29 B 0.015478f
C74 VTAIL.n30 B 0.008317f
C75 VTAIL.n31 B 0.019659f
C76 VTAIL.n32 B 0.008807f
C77 VTAIL.n33 B 0.116437f
C78 VTAIL.t4 B 0.032627f
C79 VTAIL.n34 B 0.014744f
C80 VTAIL.n35 B 0.011613f
C81 VTAIL.n36 B 0.008317f
C82 VTAIL.n37 B 1.29007f
C83 VTAIL.n38 B 0.015478f
C84 VTAIL.n39 B 0.008317f
C85 VTAIL.n40 B 0.008807f
C86 VTAIL.n41 B 0.019659f
C87 VTAIL.n42 B 0.019659f
C88 VTAIL.n43 B 0.008807f
C89 VTAIL.n44 B 0.008317f
C90 VTAIL.n45 B 0.015478f
C91 VTAIL.n46 B 0.015478f
C92 VTAIL.n47 B 0.008317f
C93 VTAIL.n48 B 0.008807f
C94 VTAIL.n49 B 0.019659f
C95 VTAIL.n50 B 0.019659f
C96 VTAIL.n51 B 0.008807f
C97 VTAIL.n52 B 0.008317f
C98 VTAIL.n53 B 0.015478f
C99 VTAIL.n54 B 0.015478f
C100 VTAIL.n55 B 0.008317f
C101 VTAIL.n56 B 0.008807f
C102 VTAIL.n57 B 0.019659f
C103 VTAIL.n58 B 0.019659f
C104 VTAIL.n59 B 0.008807f
C105 VTAIL.n60 B 0.008317f
C106 VTAIL.n61 B 0.015478f
C107 VTAIL.n62 B 0.015478f
C108 VTAIL.n63 B 0.008317f
C109 VTAIL.n64 B 0.008807f
C110 VTAIL.n65 B 0.019659f
C111 VTAIL.n66 B 0.019659f
C112 VTAIL.n67 B 0.008807f
C113 VTAIL.n68 B 0.008317f
C114 VTAIL.n69 B 0.015478f
C115 VTAIL.n70 B 0.015478f
C116 VTAIL.n71 B 0.008317f
C117 VTAIL.n72 B 0.008807f
C118 VTAIL.n73 B 0.019659f
C119 VTAIL.n74 B 0.019659f
C120 VTAIL.n75 B 0.019659f
C121 VTAIL.n76 B 0.008807f
C122 VTAIL.n77 B 0.008317f
C123 VTAIL.n78 B 0.015478f
C124 VTAIL.n79 B 0.015478f
C125 VTAIL.n80 B 0.008317f
C126 VTAIL.n81 B 0.008562f
C127 VTAIL.n82 B 0.008562f
C128 VTAIL.n83 B 0.019659f
C129 VTAIL.n84 B 0.019659f
C130 VTAIL.n85 B 0.008807f
C131 VTAIL.n86 B 0.008317f
C132 VTAIL.n87 B 0.015478f
C133 VTAIL.n88 B 0.015478f
C134 VTAIL.n89 B 0.008317f
C135 VTAIL.n90 B 0.008807f
C136 VTAIL.n91 B 0.019659f
C137 VTAIL.n92 B 0.019659f
C138 VTAIL.n93 B 0.008807f
C139 VTAIL.n94 B 0.008317f
C140 VTAIL.n95 B 0.015478f
C141 VTAIL.n96 B 0.015478f
C142 VTAIL.n97 B 0.008317f
C143 VTAIL.n98 B 0.008807f
C144 VTAIL.n99 B 0.019659f
C145 VTAIL.n100 B 0.043851f
C146 VTAIL.n101 B 0.008807f
C147 VTAIL.n102 B 0.008317f
C148 VTAIL.n103 B 0.036411f
C149 VTAIL.n104 B 0.024689f
C150 VTAIL.n105 B 0.119238f
C151 VTAIL.n106 B 0.022487f
C152 VTAIL.n107 B 0.015478f
C153 VTAIL.n108 B 0.008317f
C154 VTAIL.n109 B 0.019659f
C155 VTAIL.n110 B 0.008807f
C156 VTAIL.n111 B 0.015478f
C157 VTAIL.n112 B 0.008317f
C158 VTAIL.n113 B 0.019659f
C159 VTAIL.n114 B 0.008807f
C160 VTAIL.n115 B 0.015478f
C161 VTAIL.n116 B 0.008317f
C162 VTAIL.n117 B 0.019659f
C163 VTAIL.n118 B 0.008807f
C164 VTAIL.n119 B 0.015478f
C165 VTAIL.n120 B 0.008317f
C166 VTAIL.n121 B 0.019659f
C167 VTAIL.n122 B 0.008807f
C168 VTAIL.n123 B 0.015478f
C169 VTAIL.n124 B 0.008317f
C170 VTAIL.n125 B 0.019659f
C171 VTAIL.n126 B 0.008807f
C172 VTAIL.n127 B 0.015478f
C173 VTAIL.n128 B 0.008317f
C174 VTAIL.n129 B 0.019659f
C175 VTAIL.n130 B 0.008807f
C176 VTAIL.n131 B 0.015478f
C177 VTAIL.n132 B 0.008317f
C178 VTAIL.n133 B 0.019659f
C179 VTAIL.n134 B 0.008807f
C180 VTAIL.n135 B 0.015478f
C181 VTAIL.n136 B 0.008317f
C182 VTAIL.n137 B 0.019659f
C183 VTAIL.n138 B 0.008807f
C184 VTAIL.n139 B 0.116437f
C185 VTAIL.t2 B 0.032627f
C186 VTAIL.n140 B 0.014744f
C187 VTAIL.n141 B 0.011613f
C188 VTAIL.n142 B 0.008317f
C189 VTAIL.n143 B 1.29007f
C190 VTAIL.n144 B 0.015478f
C191 VTAIL.n145 B 0.008317f
C192 VTAIL.n146 B 0.008807f
C193 VTAIL.n147 B 0.019659f
C194 VTAIL.n148 B 0.019659f
C195 VTAIL.n149 B 0.008807f
C196 VTAIL.n150 B 0.008317f
C197 VTAIL.n151 B 0.015478f
C198 VTAIL.n152 B 0.015478f
C199 VTAIL.n153 B 0.008317f
C200 VTAIL.n154 B 0.008807f
C201 VTAIL.n155 B 0.019659f
C202 VTAIL.n156 B 0.019659f
C203 VTAIL.n157 B 0.008807f
C204 VTAIL.n158 B 0.008317f
C205 VTAIL.n159 B 0.015478f
C206 VTAIL.n160 B 0.015478f
C207 VTAIL.n161 B 0.008317f
C208 VTAIL.n162 B 0.008807f
C209 VTAIL.n163 B 0.019659f
C210 VTAIL.n164 B 0.019659f
C211 VTAIL.n165 B 0.008807f
C212 VTAIL.n166 B 0.008317f
C213 VTAIL.n167 B 0.015478f
C214 VTAIL.n168 B 0.015478f
C215 VTAIL.n169 B 0.008317f
C216 VTAIL.n170 B 0.008807f
C217 VTAIL.n171 B 0.019659f
C218 VTAIL.n172 B 0.019659f
C219 VTAIL.n173 B 0.008807f
C220 VTAIL.n174 B 0.008317f
C221 VTAIL.n175 B 0.015478f
C222 VTAIL.n176 B 0.015478f
C223 VTAIL.n177 B 0.008317f
C224 VTAIL.n178 B 0.008807f
C225 VTAIL.n179 B 0.019659f
C226 VTAIL.n180 B 0.019659f
C227 VTAIL.n181 B 0.019659f
C228 VTAIL.n182 B 0.008807f
C229 VTAIL.n183 B 0.008317f
C230 VTAIL.n184 B 0.015478f
C231 VTAIL.n185 B 0.015478f
C232 VTAIL.n186 B 0.008317f
C233 VTAIL.n187 B 0.008562f
C234 VTAIL.n188 B 0.008562f
C235 VTAIL.n189 B 0.019659f
C236 VTAIL.n190 B 0.019659f
C237 VTAIL.n191 B 0.008807f
C238 VTAIL.n192 B 0.008317f
C239 VTAIL.n193 B 0.015478f
C240 VTAIL.n194 B 0.015478f
C241 VTAIL.n195 B 0.008317f
C242 VTAIL.n196 B 0.008807f
C243 VTAIL.n197 B 0.019659f
C244 VTAIL.n198 B 0.019659f
C245 VTAIL.n199 B 0.008807f
C246 VTAIL.n200 B 0.008317f
C247 VTAIL.n201 B 0.015478f
C248 VTAIL.n202 B 0.015478f
C249 VTAIL.n203 B 0.008317f
C250 VTAIL.n204 B 0.008807f
C251 VTAIL.n205 B 0.019659f
C252 VTAIL.n206 B 0.043851f
C253 VTAIL.n207 B 0.008807f
C254 VTAIL.n208 B 0.008317f
C255 VTAIL.n209 B 0.036411f
C256 VTAIL.n210 B 0.024689f
C257 VTAIL.n211 B 0.195662f
C258 VTAIL.n212 B 0.022487f
C259 VTAIL.n213 B 0.015478f
C260 VTAIL.n214 B 0.008317f
C261 VTAIL.n215 B 0.019659f
C262 VTAIL.n216 B 0.008807f
C263 VTAIL.n217 B 0.015478f
C264 VTAIL.n218 B 0.008317f
C265 VTAIL.n219 B 0.019659f
C266 VTAIL.n220 B 0.008807f
C267 VTAIL.n221 B 0.015478f
C268 VTAIL.n222 B 0.008317f
C269 VTAIL.n223 B 0.019659f
C270 VTAIL.n224 B 0.008807f
C271 VTAIL.n225 B 0.015478f
C272 VTAIL.n226 B 0.008317f
C273 VTAIL.n227 B 0.019659f
C274 VTAIL.n228 B 0.008807f
C275 VTAIL.n229 B 0.015478f
C276 VTAIL.n230 B 0.008317f
C277 VTAIL.n231 B 0.019659f
C278 VTAIL.n232 B 0.008807f
C279 VTAIL.n233 B 0.015478f
C280 VTAIL.n234 B 0.008317f
C281 VTAIL.n235 B 0.019659f
C282 VTAIL.n236 B 0.008807f
C283 VTAIL.n237 B 0.015478f
C284 VTAIL.n238 B 0.008317f
C285 VTAIL.n239 B 0.019659f
C286 VTAIL.n240 B 0.008807f
C287 VTAIL.n241 B 0.015478f
C288 VTAIL.n242 B 0.008317f
C289 VTAIL.n243 B 0.019659f
C290 VTAIL.n244 B 0.008807f
C291 VTAIL.n245 B 0.116437f
C292 VTAIL.t0 B 0.032627f
C293 VTAIL.n246 B 0.014744f
C294 VTAIL.n247 B 0.011613f
C295 VTAIL.n248 B 0.008317f
C296 VTAIL.n249 B 1.29007f
C297 VTAIL.n250 B 0.015478f
C298 VTAIL.n251 B 0.008317f
C299 VTAIL.n252 B 0.008807f
C300 VTAIL.n253 B 0.019659f
C301 VTAIL.n254 B 0.019659f
C302 VTAIL.n255 B 0.008807f
C303 VTAIL.n256 B 0.008317f
C304 VTAIL.n257 B 0.015478f
C305 VTAIL.n258 B 0.015478f
C306 VTAIL.n259 B 0.008317f
C307 VTAIL.n260 B 0.008807f
C308 VTAIL.n261 B 0.019659f
C309 VTAIL.n262 B 0.019659f
C310 VTAIL.n263 B 0.008807f
C311 VTAIL.n264 B 0.008317f
C312 VTAIL.n265 B 0.015478f
C313 VTAIL.n266 B 0.015478f
C314 VTAIL.n267 B 0.008317f
C315 VTAIL.n268 B 0.008807f
C316 VTAIL.n269 B 0.019659f
C317 VTAIL.n270 B 0.019659f
C318 VTAIL.n271 B 0.008807f
C319 VTAIL.n272 B 0.008317f
C320 VTAIL.n273 B 0.015478f
C321 VTAIL.n274 B 0.015478f
C322 VTAIL.n275 B 0.008317f
C323 VTAIL.n276 B 0.008807f
C324 VTAIL.n277 B 0.019659f
C325 VTAIL.n278 B 0.019659f
C326 VTAIL.n279 B 0.008807f
C327 VTAIL.n280 B 0.008317f
C328 VTAIL.n281 B 0.015478f
C329 VTAIL.n282 B 0.015478f
C330 VTAIL.n283 B 0.008317f
C331 VTAIL.n284 B 0.008807f
C332 VTAIL.n285 B 0.019659f
C333 VTAIL.n286 B 0.019659f
C334 VTAIL.n287 B 0.019659f
C335 VTAIL.n288 B 0.008807f
C336 VTAIL.n289 B 0.008317f
C337 VTAIL.n290 B 0.015478f
C338 VTAIL.n291 B 0.015478f
C339 VTAIL.n292 B 0.008317f
C340 VTAIL.n293 B 0.008562f
C341 VTAIL.n294 B 0.008562f
C342 VTAIL.n295 B 0.019659f
C343 VTAIL.n296 B 0.019659f
C344 VTAIL.n297 B 0.008807f
C345 VTAIL.n298 B 0.008317f
C346 VTAIL.n299 B 0.015478f
C347 VTAIL.n300 B 0.015478f
C348 VTAIL.n301 B 0.008317f
C349 VTAIL.n302 B 0.008807f
C350 VTAIL.n303 B 0.019659f
C351 VTAIL.n304 B 0.019659f
C352 VTAIL.n305 B 0.008807f
C353 VTAIL.n306 B 0.008317f
C354 VTAIL.n307 B 0.015478f
C355 VTAIL.n308 B 0.015478f
C356 VTAIL.n309 B 0.008317f
C357 VTAIL.n310 B 0.008807f
C358 VTAIL.n311 B 0.019659f
C359 VTAIL.n312 B 0.043851f
C360 VTAIL.n313 B 0.008807f
C361 VTAIL.n314 B 0.008317f
C362 VTAIL.n315 B 0.036411f
C363 VTAIL.n316 B 0.024689f
C364 VTAIL.n317 B 1.35761f
C365 VTAIL.n318 B 0.022487f
C366 VTAIL.n319 B 0.015478f
C367 VTAIL.n320 B 0.008317f
C368 VTAIL.n321 B 0.019659f
C369 VTAIL.n322 B 0.008807f
C370 VTAIL.n323 B 0.015478f
C371 VTAIL.n324 B 0.008317f
C372 VTAIL.n325 B 0.019659f
C373 VTAIL.n326 B 0.008807f
C374 VTAIL.n327 B 0.015478f
C375 VTAIL.n328 B 0.008317f
C376 VTAIL.n329 B 0.019659f
C377 VTAIL.n330 B 0.008807f
C378 VTAIL.n331 B 0.015478f
C379 VTAIL.n332 B 0.008317f
C380 VTAIL.n333 B 0.019659f
C381 VTAIL.n334 B 0.019659f
C382 VTAIL.n335 B 0.008807f
C383 VTAIL.n336 B 0.015478f
C384 VTAIL.n337 B 0.008317f
C385 VTAIL.n338 B 0.019659f
C386 VTAIL.n339 B 0.008807f
C387 VTAIL.n340 B 0.015478f
C388 VTAIL.n341 B 0.008317f
C389 VTAIL.n342 B 0.019659f
C390 VTAIL.n343 B 0.008807f
C391 VTAIL.n344 B 0.015478f
C392 VTAIL.n345 B 0.008317f
C393 VTAIL.n346 B 0.019659f
C394 VTAIL.n347 B 0.008807f
C395 VTAIL.n348 B 0.015478f
C396 VTAIL.n349 B 0.008317f
C397 VTAIL.n350 B 0.019659f
C398 VTAIL.n351 B 0.008807f
C399 VTAIL.n352 B 0.116437f
C400 VTAIL.t7 B 0.032627f
C401 VTAIL.n353 B 0.014744f
C402 VTAIL.n354 B 0.011613f
C403 VTAIL.n355 B 0.008317f
C404 VTAIL.n356 B 1.29007f
C405 VTAIL.n357 B 0.015478f
C406 VTAIL.n358 B 0.008317f
C407 VTAIL.n359 B 0.008807f
C408 VTAIL.n360 B 0.019659f
C409 VTAIL.n361 B 0.019659f
C410 VTAIL.n362 B 0.008807f
C411 VTAIL.n363 B 0.008317f
C412 VTAIL.n364 B 0.015478f
C413 VTAIL.n365 B 0.015478f
C414 VTAIL.n366 B 0.008317f
C415 VTAIL.n367 B 0.008807f
C416 VTAIL.n368 B 0.019659f
C417 VTAIL.n369 B 0.019659f
C418 VTAIL.n370 B 0.008807f
C419 VTAIL.n371 B 0.008317f
C420 VTAIL.n372 B 0.015478f
C421 VTAIL.n373 B 0.015478f
C422 VTAIL.n374 B 0.008317f
C423 VTAIL.n375 B 0.008807f
C424 VTAIL.n376 B 0.019659f
C425 VTAIL.n377 B 0.019659f
C426 VTAIL.n378 B 0.008807f
C427 VTAIL.n379 B 0.008317f
C428 VTAIL.n380 B 0.015478f
C429 VTAIL.n381 B 0.015478f
C430 VTAIL.n382 B 0.008317f
C431 VTAIL.n383 B 0.008807f
C432 VTAIL.n384 B 0.019659f
C433 VTAIL.n385 B 0.019659f
C434 VTAIL.n386 B 0.008807f
C435 VTAIL.n387 B 0.008317f
C436 VTAIL.n388 B 0.015478f
C437 VTAIL.n389 B 0.015478f
C438 VTAIL.n390 B 0.008317f
C439 VTAIL.n391 B 0.008807f
C440 VTAIL.n392 B 0.019659f
C441 VTAIL.n393 B 0.019659f
C442 VTAIL.n394 B 0.008807f
C443 VTAIL.n395 B 0.008317f
C444 VTAIL.n396 B 0.015478f
C445 VTAIL.n397 B 0.015478f
C446 VTAIL.n398 B 0.008317f
C447 VTAIL.n399 B 0.008562f
C448 VTAIL.n400 B 0.008562f
C449 VTAIL.n401 B 0.019659f
C450 VTAIL.n402 B 0.019659f
C451 VTAIL.n403 B 0.008807f
C452 VTAIL.n404 B 0.008317f
C453 VTAIL.n405 B 0.015478f
C454 VTAIL.n406 B 0.015478f
C455 VTAIL.n407 B 0.008317f
C456 VTAIL.n408 B 0.008807f
C457 VTAIL.n409 B 0.019659f
C458 VTAIL.n410 B 0.019659f
C459 VTAIL.n411 B 0.008807f
C460 VTAIL.n412 B 0.008317f
C461 VTAIL.n413 B 0.015478f
C462 VTAIL.n414 B 0.015478f
C463 VTAIL.n415 B 0.008317f
C464 VTAIL.n416 B 0.008807f
C465 VTAIL.n417 B 0.019659f
C466 VTAIL.n418 B 0.043851f
C467 VTAIL.n419 B 0.008807f
C468 VTAIL.n420 B 0.008317f
C469 VTAIL.n421 B 0.036411f
C470 VTAIL.n422 B 0.024689f
C471 VTAIL.n423 B 1.35761f
C472 VTAIL.n424 B 0.022487f
C473 VTAIL.n425 B 0.015478f
C474 VTAIL.n426 B 0.008317f
C475 VTAIL.n427 B 0.019659f
C476 VTAIL.n428 B 0.008807f
C477 VTAIL.n429 B 0.015478f
C478 VTAIL.n430 B 0.008317f
C479 VTAIL.n431 B 0.019659f
C480 VTAIL.n432 B 0.008807f
C481 VTAIL.n433 B 0.015478f
C482 VTAIL.n434 B 0.008317f
C483 VTAIL.n435 B 0.019659f
C484 VTAIL.n436 B 0.008807f
C485 VTAIL.n437 B 0.015478f
C486 VTAIL.n438 B 0.008317f
C487 VTAIL.n439 B 0.019659f
C488 VTAIL.n440 B 0.019659f
C489 VTAIL.n441 B 0.008807f
C490 VTAIL.n442 B 0.015478f
C491 VTAIL.n443 B 0.008317f
C492 VTAIL.n444 B 0.019659f
C493 VTAIL.n445 B 0.008807f
C494 VTAIL.n446 B 0.015478f
C495 VTAIL.n447 B 0.008317f
C496 VTAIL.n448 B 0.019659f
C497 VTAIL.n449 B 0.008807f
C498 VTAIL.n450 B 0.015478f
C499 VTAIL.n451 B 0.008317f
C500 VTAIL.n452 B 0.019659f
C501 VTAIL.n453 B 0.008807f
C502 VTAIL.n454 B 0.015478f
C503 VTAIL.n455 B 0.008317f
C504 VTAIL.n456 B 0.019659f
C505 VTAIL.n457 B 0.008807f
C506 VTAIL.n458 B 0.116437f
C507 VTAIL.t6 B 0.032627f
C508 VTAIL.n459 B 0.014744f
C509 VTAIL.n460 B 0.011613f
C510 VTAIL.n461 B 0.008317f
C511 VTAIL.n462 B 1.29007f
C512 VTAIL.n463 B 0.015478f
C513 VTAIL.n464 B 0.008317f
C514 VTAIL.n465 B 0.008807f
C515 VTAIL.n466 B 0.019659f
C516 VTAIL.n467 B 0.019659f
C517 VTAIL.n468 B 0.008807f
C518 VTAIL.n469 B 0.008317f
C519 VTAIL.n470 B 0.015478f
C520 VTAIL.n471 B 0.015478f
C521 VTAIL.n472 B 0.008317f
C522 VTAIL.n473 B 0.008807f
C523 VTAIL.n474 B 0.019659f
C524 VTAIL.n475 B 0.019659f
C525 VTAIL.n476 B 0.008807f
C526 VTAIL.n477 B 0.008317f
C527 VTAIL.n478 B 0.015478f
C528 VTAIL.n479 B 0.015478f
C529 VTAIL.n480 B 0.008317f
C530 VTAIL.n481 B 0.008807f
C531 VTAIL.n482 B 0.019659f
C532 VTAIL.n483 B 0.019659f
C533 VTAIL.n484 B 0.008807f
C534 VTAIL.n485 B 0.008317f
C535 VTAIL.n486 B 0.015478f
C536 VTAIL.n487 B 0.015478f
C537 VTAIL.n488 B 0.008317f
C538 VTAIL.n489 B 0.008807f
C539 VTAIL.n490 B 0.019659f
C540 VTAIL.n491 B 0.019659f
C541 VTAIL.n492 B 0.008807f
C542 VTAIL.n493 B 0.008317f
C543 VTAIL.n494 B 0.015478f
C544 VTAIL.n495 B 0.015478f
C545 VTAIL.n496 B 0.008317f
C546 VTAIL.n497 B 0.008807f
C547 VTAIL.n498 B 0.019659f
C548 VTAIL.n499 B 0.019659f
C549 VTAIL.n500 B 0.008807f
C550 VTAIL.n501 B 0.008317f
C551 VTAIL.n502 B 0.015478f
C552 VTAIL.n503 B 0.015478f
C553 VTAIL.n504 B 0.008317f
C554 VTAIL.n505 B 0.008562f
C555 VTAIL.n506 B 0.008562f
C556 VTAIL.n507 B 0.019659f
C557 VTAIL.n508 B 0.019659f
C558 VTAIL.n509 B 0.008807f
C559 VTAIL.n510 B 0.008317f
C560 VTAIL.n511 B 0.015478f
C561 VTAIL.n512 B 0.015478f
C562 VTAIL.n513 B 0.008317f
C563 VTAIL.n514 B 0.008807f
C564 VTAIL.n515 B 0.019659f
C565 VTAIL.n516 B 0.019659f
C566 VTAIL.n517 B 0.008807f
C567 VTAIL.n518 B 0.008317f
C568 VTAIL.n519 B 0.015478f
C569 VTAIL.n520 B 0.015478f
C570 VTAIL.n521 B 0.008317f
C571 VTAIL.n522 B 0.008807f
C572 VTAIL.n523 B 0.019659f
C573 VTAIL.n524 B 0.043851f
C574 VTAIL.n525 B 0.008807f
C575 VTAIL.n526 B 0.008317f
C576 VTAIL.n527 B 0.036411f
C577 VTAIL.n528 B 0.024689f
C578 VTAIL.n529 B 0.195662f
C579 VTAIL.n530 B 0.022487f
C580 VTAIL.n531 B 0.015478f
C581 VTAIL.n532 B 0.008317f
C582 VTAIL.n533 B 0.019659f
C583 VTAIL.n534 B 0.008807f
C584 VTAIL.n535 B 0.015478f
C585 VTAIL.n536 B 0.008317f
C586 VTAIL.n537 B 0.019659f
C587 VTAIL.n538 B 0.008807f
C588 VTAIL.n539 B 0.015478f
C589 VTAIL.n540 B 0.008317f
C590 VTAIL.n541 B 0.019659f
C591 VTAIL.n542 B 0.008807f
C592 VTAIL.n543 B 0.015478f
C593 VTAIL.n544 B 0.008317f
C594 VTAIL.n545 B 0.019659f
C595 VTAIL.n546 B 0.019659f
C596 VTAIL.n547 B 0.008807f
C597 VTAIL.n548 B 0.015478f
C598 VTAIL.n549 B 0.008317f
C599 VTAIL.n550 B 0.019659f
C600 VTAIL.n551 B 0.008807f
C601 VTAIL.n552 B 0.015478f
C602 VTAIL.n553 B 0.008317f
C603 VTAIL.n554 B 0.019659f
C604 VTAIL.n555 B 0.008807f
C605 VTAIL.n556 B 0.015478f
C606 VTAIL.n557 B 0.008317f
C607 VTAIL.n558 B 0.019659f
C608 VTAIL.n559 B 0.008807f
C609 VTAIL.n560 B 0.015478f
C610 VTAIL.n561 B 0.008317f
C611 VTAIL.n562 B 0.019659f
C612 VTAIL.n563 B 0.008807f
C613 VTAIL.n564 B 0.116437f
C614 VTAIL.t1 B 0.032627f
C615 VTAIL.n565 B 0.014744f
C616 VTAIL.n566 B 0.011613f
C617 VTAIL.n567 B 0.008317f
C618 VTAIL.n568 B 1.29007f
C619 VTAIL.n569 B 0.015478f
C620 VTAIL.n570 B 0.008317f
C621 VTAIL.n571 B 0.008807f
C622 VTAIL.n572 B 0.019659f
C623 VTAIL.n573 B 0.019659f
C624 VTAIL.n574 B 0.008807f
C625 VTAIL.n575 B 0.008317f
C626 VTAIL.n576 B 0.015478f
C627 VTAIL.n577 B 0.015478f
C628 VTAIL.n578 B 0.008317f
C629 VTAIL.n579 B 0.008807f
C630 VTAIL.n580 B 0.019659f
C631 VTAIL.n581 B 0.019659f
C632 VTAIL.n582 B 0.008807f
C633 VTAIL.n583 B 0.008317f
C634 VTAIL.n584 B 0.015478f
C635 VTAIL.n585 B 0.015478f
C636 VTAIL.n586 B 0.008317f
C637 VTAIL.n587 B 0.008807f
C638 VTAIL.n588 B 0.019659f
C639 VTAIL.n589 B 0.019659f
C640 VTAIL.n590 B 0.008807f
C641 VTAIL.n591 B 0.008317f
C642 VTAIL.n592 B 0.015478f
C643 VTAIL.n593 B 0.015478f
C644 VTAIL.n594 B 0.008317f
C645 VTAIL.n595 B 0.008807f
C646 VTAIL.n596 B 0.019659f
C647 VTAIL.n597 B 0.019659f
C648 VTAIL.n598 B 0.008807f
C649 VTAIL.n599 B 0.008317f
C650 VTAIL.n600 B 0.015478f
C651 VTAIL.n601 B 0.015478f
C652 VTAIL.n602 B 0.008317f
C653 VTAIL.n603 B 0.008807f
C654 VTAIL.n604 B 0.019659f
C655 VTAIL.n605 B 0.019659f
C656 VTAIL.n606 B 0.008807f
C657 VTAIL.n607 B 0.008317f
C658 VTAIL.n608 B 0.015478f
C659 VTAIL.n609 B 0.015478f
C660 VTAIL.n610 B 0.008317f
C661 VTAIL.n611 B 0.008562f
C662 VTAIL.n612 B 0.008562f
C663 VTAIL.n613 B 0.019659f
C664 VTAIL.n614 B 0.019659f
C665 VTAIL.n615 B 0.008807f
C666 VTAIL.n616 B 0.008317f
C667 VTAIL.n617 B 0.015478f
C668 VTAIL.n618 B 0.015478f
C669 VTAIL.n619 B 0.008317f
C670 VTAIL.n620 B 0.008807f
C671 VTAIL.n621 B 0.019659f
C672 VTAIL.n622 B 0.019659f
C673 VTAIL.n623 B 0.008807f
C674 VTAIL.n624 B 0.008317f
C675 VTAIL.n625 B 0.015478f
C676 VTAIL.n626 B 0.015478f
C677 VTAIL.n627 B 0.008317f
C678 VTAIL.n628 B 0.008807f
C679 VTAIL.n629 B 0.019659f
C680 VTAIL.n630 B 0.043851f
C681 VTAIL.n631 B 0.008807f
C682 VTAIL.n632 B 0.008317f
C683 VTAIL.n633 B 0.036411f
C684 VTAIL.n634 B 0.024689f
C685 VTAIL.n635 B 0.195662f
C686 VTAIL.n636 B 0.022487f
C687 VTAIL.n637 B 0.015478f
C688 VTAIL.n638 B 0.008317f
C689 VTAIL.n639 B 0.019659f
C690 VTAIL.n640 B 0.008807f
C691 VTAIL.n641 B 0.015478f
C692 VTAIL.n642 B 0.008317f
C693 VTAIL.n643 B 0.019659f
C694 VTAIL.n644 B 0.008807f
C695 VTAIL.n645 B 0.015478f
C696 VTAIL.n646 B 0.008317f
C697 VTAIL.n647 B 0.019659f
C698 VTAIL.n648 B 0.008807f
C699 VTAIL.n649 B 0.015478f
C700 VTAIL.n650 B 0.008317f
C701 VTAIL.n651 B 0.019659f
C702 VTAIL.n652 B 0.019659f
C703 VTAIL.n653 B 0.008807f
C704 VTAIL.n654 B 0.015478f
C705 VTAIL.n655 B 0.008317f
C706 VTAIL.n656 B 0.019659f
C707 VTAIL.n657 B 0.008807f
C708 VTAIL.n658 B 0.015478f
C709 VTAIL.n659 B 0.008317f
C710 VTAIL.n660 B 0.019659f
C711 VTAIL.n661 B 0.008807f
C712 VTAIL.n662 B 0.015478f
C713 VTAIL.n663 B 0.008317f
C714 VTAIL.n664 B 0.019659f
C715 VTAIL.n665 B 0.008807f
C716 VTAIL.n666 B 0.015478f
C717 VTAIL.n667 B 0.008317f
C718 VTAIL.n668 B 0.019659f
C719 VTAIL.n669 B 0.008807f
C720 VTAIL.n670 B 0.116437f
C721 VTAIL.t3 B 0.032627f
C722 VTAIL.n671 B 0.014744f
C723 VTAIL.n672 B 0.011613f
C724 VTAIL.n673 B 0.008317f
C725 VTAIL.n674 B 1.29007f
C726 VTAIL.n675 B 0.015478f
C727 VTAIL.n676 B 0.008317f
C728 VTAIL.n677 B 0.008807f
C729 VTAIL.n678 B 0.019659f
C730 VTAIL.n679 B 0.019659f
C731 VTAIL.n680 B 0.008807f
C732 VTAIL.n681 B 0.008317f
C733 VTAIL.n682 B 0.015478f
C734 VTAIL.n683 B 0.015478f
C735 VTAIL.n684 B 0.008317f
C736 VTAIL.n685 B 0.008807f
C737 VTAIL.n686 B 0.019659f
C738 VTAIL.n687 B 0.019659f
C739 VTAIL.n688 B 0.008807f
C740 VTAIL.n689 B 0.008317f
C741 VTAIL.n690 B 0.015478f
C742 VTAIL.n691 B 0.015478f
C743 VTAIL.n692 B 0.008317f
C744 VTAIL.n693 B 0.008807f
C745 VTAIL.n694 B 0.019659f
C746 VTAIL.n695 B 0.019659f
C747 VTAIL.n696 B 0.008807f
C748 VTAIL.n697 B 0.008317f
C749 VTAIL.n698 B 0.015478f
C750 VTAIL.n699 B 0.015478f
C751 VTAIL.n700 B 0.008317f
C752 VTAIL.n701 B 0.008807f
C753 VTAIL.n702 B 0.019659f
C754 VTAIL.n703 B 0.019659f
C755 VTAIL.n704 B 0.008807f
C756 VTAIL.n705 B 0.008317f
C757 VTAIL.n706 B 0.015478f
C758 VTAIL.n707 B 0.015478f
C759 VTAIL.n708 B 0.008317f
C760 VTAIL.n709 B 0.008807f
C761 VTAIL.n710 B 0.019659f
C762 VTAIL.n711 B 0.019659f
C763 VTAIL.n712 B 0.008807f
C764 VTAIL.n713 B 0.008317f
C765 VTAIL.n714 B 0.015478f
C766 VTAIL.n715 B 0.015478f
C767 VTAIL.n716 B 0.008317f
C768 VTAIL.n717 B 0.008562f
C769 VTAIL.n718 B 0.008562f
C770 VTAIL.n719 B 0.019659f
C771 VTAIL.n720 B 0.019659f
C772 VTAIL.n721 B 0.008807f
C773 VTAIL.n722 B 0.008317f
C774 VTAIL.n723 B 0.015478f
C775 VTAIL.n724 B 0.015478f
C776 VTAIL.n725 B 0.008317f
C777 VTAIL.n726 B 0.008807f
C778 VTAIL.n727 B 0.019659f
C779 VTAIL.n728 B 0.019659f
C780 VTAIL.n729 B 0.008807f
C781 VTAIL.n730 B 0.008317f
C782 VTAIL.n731 B 0.015478f
C783 VTAIL.n732 B 0.015478f
C784 VTAIL.n733 B 0.008317f
C785 VTAIL.n734 B 0.008807f
C786 VTAIL.n735 B 0.019659f
C787 VTAIL.n736 B 0.043851f
C788 VTAIL.n737 B 0.008807f
C789 VTAIL.n738 B 0.008317f
C790 VTAIL.n739 B 0.036411f
C791 VTAIL.n740 B 0.024689f
C792 VTAIL.n741 B 1.35761f
C793 VTAIL.n742 B 0.022487f
C794 VTAIL.n743 B 0.015478f
C795 VTAIL.n744 B 0.008317f
C796 VTAIL.n745 B 0.019659f
C797 VTAIL.n746 B 0.008807f
C798 VTAIL.n747 B 0.015478f
C799 VTAIL.n748 B 0.008317f
C800 VTAIL.n749 B 0.019659f
C801 VTAIL.n750 B 0.008807f
C802 VTAIL.n751 B 0.015478f
C803 VTAIL.n752 B 0.008317f
C804 VTAIL.n753 B 0.019659f
C805 VTAIL.n754 B 0.008807f
C806 VTAIL.n755 B 0.015478f
C807 VTAIL.n756 B 0.008317f
C808 VTAIL.n757 B 0.019659f
C809 VTAIL.n758 B 0.008807f
C810 VTAIL.n759 B 0.015478f
C811 VTAIL.n760 B 0.008317f
C812 VTAIL.n761 B 0.019659f
C813 VTAIL.n762 B 0.008807f
C814 VTAIL.n763 B 0.015478f
C815 VTAIL.n764 B 0.008317f
C816 VTAIL.n765 B 0.019659f
C817 VTAIL.n766 B 0.008807f
C818 VTAIL.n767 B 0.015478f
C819 VTAIL.n768 B 0.008317f
C820 VTAIL.n769 B 0.019659f
C821 VTAIL.n770 B 0.008807f
C822 VTAIL.n771 B 0.015478f
C823 VTAIL.n772 B 0.008317f
C824 VTAIL.n773 B 0.019659f
C825 VTAIL.n774 B 0.008807f
C826 VTAIL.n775 B 0.116437f
C827 VTAIL.t5 B 0.032627f
C828 VTAIL.n776 B 0.014744f
C829 VTAIL.n777 B 0.011613f
C830 VTAIL.n778 B 0.008317f
C831 VTAIL.n779 B 1.29007f
C832 VTAIL.n780 B 0.015478f
C833 VTAIL.n781 B 0.008317f
C834 VTAIL.n782 B 0.008807f
C835 VTAIL.n783 B 0.019659f
C836 VTAIL.n784 B 0.019659f
C837 VTAIL.n785 B 0.008807f
C838 VTAIL.n786 B 0.008317f
C839 VTAIL.n787 B 0.015478f
C840 VTAIL.n788 B 0.015478f
C841 VTAIL.n789 B 0.008317f
C842 VTAIL.n790 B 0.008807f
C843 VTAIL.n791 B 0.019659f
C844 VTAIL.n792 B 0.019659f
C845 VTAIL.n793 B 0.008807f
C846 VTAIL.n794 B 0.008317f
C847 VTAIL.n795 B 0.015478f
C848 VTAIL.n796 B 0.015478f
C849 VTAIL.n797 B 0.008317f
C850 VTAIL.n798 B 0.008807f
C851 VTAIL.n799 B 0.019659f
C852 VTAIL.n800 B 0.019659f
C853 VTAIL.n801 B 0.008807f
C854 VTAIL.n802 B 0.008317f
C855 VTAIL.n803 B 0.015478f
C856 VTAIL.n804 B 0.015478f
C857 VTAIL.n805 B 0.008317f
C858 VTAIL.n806 B 0.008807f
C859 VTAIL.n807 B 0.019659f
C860 VTAIL.n808 B 0.019659f
C861 VTAIL.n809 B 0.008807f
C862 VTAIL.n810 B 0.008317f
C863 VTAIL.n811 B 0.015478f
C864 VTAIL.n812 B 0.015478f
C865 VTAIL.n813 B 0.008317f
C866 VTAIL.n814 B 0.008807f
C867 VTAIL.n815 B 0.019659f
C868 VTAIL.n816 B 0.019659f
C869 VTAIL.n817 B 0.019659f
C870 VTAIL.n818 B 0.008807f
C871 VTAIL.n819 B 0.008317f
C872 VTAIL.n820 B 0.015478f
C873 VTAIL.n821 B 0.015478f
C874 VTAIL.n822 B 0.008317f
C875 VTAIL.n823 B 0.008562f
C876 VTAIL.n824 B 0.008562f
C877 VTAIL.n825 B 0.019659f
C878 VTAIL.n826 B 0.019659f
C879 VTAIL.n827 B 0.008807f
C880 VTAIL.n828 B 0.008317f
C881 VTAIL.n829 B 0.015478f
C882 VTAIL.n830 B 0.015478f
C883 VTAIL.n831 B 0.008317f
C884 VTAIL.n832 B 0.008807f
C885 VTAIL.n833 B 0.019659f
C886 VTAIL.n834 B 0.019659f
C887 VTAIL.n835 B 0.008807f
C888 VTAIL.n836 B 0.008317f
C889 VTAIL.n837 B 0.015478f
C890 VTAIL.n838 B 0.015478f
C891 VTAIL.n839 B 0.008317f
C892 VTAIL.n840 B 0.008807f
C893 VTAIL.n841 B 0.019659f
C894 VTAIL.n842 B 0.043851f
C895 VTAIL.n843 B 0.008807f
C896 VTAIL.n844 B 0.008317f
C897 VTAIL.n845 B 0.036411f
C898 VTAIL.n846 B 0.024689f
C899 VTAIL.n847 B 1.27538f
C900 VDD2.t2 B 0.398664f
C901 VDD2.t3 B 0.398664f
C902 VDD2.n0 B 4.61675f
C903 VDD2.t1 B 0.398664f
C904 VDD2.t0 B 0.398664f
C905 VDD2.n1 B 3.6397f
C906 VDD2.n2 B 4.67087f
C907 VN.t2 B 3.80019f
C908 VN.t3 B 3.80891f
C909 VN.n0 B 2.34633f
C910 VN.t0 B 3.80019f
C911 VN.t1 B 3.80891f
C912 VN.n1 B 3.77101f
.ends

