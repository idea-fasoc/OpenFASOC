* NGSPICE file created from diff_pair_sample_0051.ext - technology: sky130A

.subckt diff_pair_sample_0051 VTAIL VN VP B VDD2 VDD1
X0 B.t19 B.t17 B.t18 B.t11 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=2.65
X1 B.t16 B.t14 B.t15 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=2.65
X2 VDD2.t5 VN.t0 VTAIL.t9 B.t2 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=2.65
X3 VTAIL.t7 VN.t1 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=2.65
X4 VDD1.t5 VP.t0 VTAIL.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=2.65
X5 VDD1.t4 VP.t1 VTAIL.t5 B.t2 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=2.65
X6 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=2.65
X7 VDD1.t3 VP.t2 VTAIL.t2 B.t5 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=2.65
X8 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=0 ps=0 w=16.16 l=2.65
X9 VDD2.t3 VN.t2 VTAIL.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=2.65
X10 VDD2.t2 VN.t3 VTAIL.t8 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=2.65
X11 VTAIL.t0 VP.t3 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=2.65
X12 VDD2.t1 VN.t4 VTAIL.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=6.3024 pd=33.1 as=2.6664 ps=16.49 w=16.16 l=2.65
X13 VTAIL.t3 VP.t4 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=2.65
X14 VTAIL.t10 VN.t5 VDD2.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=2.6664 ps=16.49 w=16.16 l=2.65
X15 VDD1.t0 VP.t5 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.6664 pd=16.49 as=6.3024 ps=33.1 w=16.16 l=2.65
R0 B.n940 B.n939 585
R1 B.n941 B.n940 585
R2 B.n373 B.n139 585
R3 B.n372 B.n371 585
R4 B.n370 B.n369 585
R5 B.n368 B.n367 585
R6 B.n366 B.n365 585
R7 B.n364 B.n363 585
R8 B.n362 B.n361 585
R9 B.n360 B.n359 585
R10 B.n358 B.n357 585
R11 B.n356 B.n355 585
R12 B.n354 B.n353 585
R13 B.n352 B.n351 585
R14 B.n350 B.n349 585
R15 B.n348 B.n347 585
R16 B.n346 B.n345 585
R17 B.n344 B.n343 585
R18 B.n342 B.n341 585
R19 B.n340 B.n339 585
R20 B.n338 B.n337 585
R21 B.n336 B.n335 585
R22 B.n334 B.n333 585
R23 B.n332 B.n331 585
R24 B.n330 B.n329 585
R25 B.n328 B.n327 585
R26 B.n326 B.n325 585
R27 B.n324 B.n323 585
R28 B.n322 B.n321 585
R29 B.n320 B.n319 585
R30 B.n318 B.n317 585
R31 B.n316 B.n315 585
R32 B.n314 B.n313 585
R33 B.n312 B.n311 585
R34 B.n310 B.n309 585
R35 B.n308 B.n307 585
R36 B.n306 B.n305 585
R37 B.n304 B.n303 585
R38 B.n302 B.n301 585
R39 B.n300 B.n299 585
R40 B.n298 B.n297 585
R41 B.n296 B.n295 585
R42 B.n294 B.n293 585
R43 B.n292 B.n291 585
R44 B.n290 B.n289 585
R45 B.n288 B.n287 585
R46 B.n286 B.n285 585
R47 B.n284 B.n283 585
R48 B.n282 B.n281 585
R49 B.n280 B.n279 585
R50 B.n278 B.n277 585
R51 B.n276 B.n275 585
R52 B.n274 B.n273 585
R53 B.n272 B.n271 585
R54 B.n270 B.n269 585
R55 B.n267 B.n266 585
R56 B.n265 B.n264 585
R57 B.n263 B.n262 585
R58 B.n261 B.n260 585
R59 B.n259 B.n258 585
R60 B.n257 B.n256 585
R61 B.n255 B.n254 585
R62 B.n253 B.n252 585
R63 B.n251 B.n250 585
R64 B.n249 B.n248 585
R65 B.n247 B.n246 585
R66 B.n245 B.n244 585
R67 B.n243 B.n242 585
R68 B.n241 B.n240 585
R69 B.n239 B.n238 585
R70 B.n237 B.n236 585
R71 B.n235 B.n234 585
R72 B.n233 B.n232 585
R73 B.n231 B.n230 585
R74 B.n229 B.n228 585
R75 B.n227 B.n226 585
R76 B.n225 B.n224 585
R77 B.n223 B.n222 585
R78 B.n221 B.n220 585
R79 B.n219 B.n218 585
R80 B.n217 B.n216 585
R81 B.n215 B.n214 585
R82 B.n213 B.n212 585
R83 B.n211 B.n210 585
R84 B.n209 B.n208 585
R85 B.n207 B.n206 585
R86 B.n205 B.n204 585
R87 B.n203 B.n202 585
R88 B.n201 B.n200 585
R89 B.n199 B.n198 585
R90 B.n197 B.n196 585
R91 B.n195 B.n194 585
R92 B.n193 B.n192 585
R93 B.n191 B.n190 585
R94 B.n189 B.n188 585
R95 B.n187 B.n186 585
R96 B.n185 B.n184 585
R97 B.n183 B.n182 585
R98 B.n181 B.n180 585
R99 B.n179 B.n178 585
R100 B.n177 B.n176 585
R101 B.n175 B.n174 585
R102 B.n173 B.n172 585
R103 B.n171 B.n170 585
R104 B.n169 B.n168 585
R105 B.n167 B.n166 585
R106 B.n165 B.n164 585
R107 B.n163 B.n162 585
R108 B.n161 B.n160 585
R109 B.n159 B.n158 585
R110 B.n157 B.n156 585
R111 B.n155 B.n154 585
R112 B.n153 B.n152 585
R113 B.n151 B.n150 585
R114 B.n149 B.n148 585
R115 B.n147 B.n146 585
R116 B.n81 B.n80 585
R117 B.n944 B.n943 585
R118 B.n938 B.n140 585
R119 B.n140 B.n78 585
R120 B.n937 B.n77 585
R121 B.n948 B.n77 585
R122 B.n936 B.n76 585
R123 B.n949 B.n76 585
R124 B.n935 B.n75 585
R125 B.n950 B.n75 585
R126 B.n934 B.n933 585
R127 B.n933 B.n71 585
R128 B.n932 B.n70 585
R129 B.n956 B.n70 585
R130 B.n931 B.n69 585
R131 B.n957 B.n69 585
R132 B.n930 B.n68 585
R133 B.n958 B.n68 585
R134 B.n929 B.n928 585
R135 B.n928 B.n64 585
R136 B.n927 B.n63 585
R137 B.n964 B.n63 585
R138 B.n926 B.n62 585
R139 B.n965 B.n62 585
R140 B.n925 B.n61 585
R141 B.n966 B.n61 585
R142 B.n924 B.n923 585
R143 B.n923 B.n57 585
R144 B.n922 B.n56 585
R145 B.n972 B.n56 585
R146 B.n921 B.n55 585
R147 B.n973 B.n55 585
R148 B.n920 B.n54 585
R149 B.n974 B.n54 585
R150 B.n919 B.n918 585
R151 B.n918 B.n50 585
R152 B.n917 B.n49 585
R153 B.n980 B.n49 585
R154 B.n916 B.n48 585
R155 B.n981 B.n48 585
R156 B.n915 B.n47 585
R157 B.n982 B.n47 585
R158 B.n914 B.n913 585
R159 B.n913 B.n43 585
R160 B.n912 B.n42 585
R161 B.n988 B.n42 585
R162 B.n911 B.n41 585
R163 B.n989 B.n41 585
R164 B.n910 B.n40 585
R165 B.n990 B.n40 585
R166 B.n909 B.n908 585
R167 B.n908 B.n36 585
R168 B.n907 B.n35 585
R169 B.n996 B.n35 585
R170 B.n906 B.n34 585
R171 B.n997 B.n34 585
R172 B.n905 B.n33 585
R173 B.n998 B.n33 585
R174 B.n904 B.n903 585
R175 B.n903 B.n32 585
R176 B.n902 B.n28 585
R177 B.n1004 B.n28 585
R178 B.n901 B.n27 585
R179 B.n1005 B.n27 585
R180 B.n900 B.n26 585
R181 B.n1006 B.n26 585
R182 B.n899 B.n898 585
R183 B.n898 B.n22 585
R184 B.n897 B.n21 585
R185 B.n1012 B.n21 585
R186 B.n896 B.n20 585
R187 B.n1013 B.n20 585
R188 B.n895 B.n19 585
R189 B.n1014 B.n19 585
R190 B.n894 B.n893 585
R191 B.n893 B.n15 585
R192 B.n892 B.n14 585
R193 B.n1020 B.n14 585
R194 B.n891 B.n13 585
R195 B.n1021 B.n13 585
R196 B.n890 B.n12 585
R197 B.n1022 B.n12 585
R198 B.n889 B.n888 585
R199 B.n888 B.n8 585
R200 B.n887 B.n7 585
R201 B.n1028 B.n7 585
R202 B.n886 B.n6 585
R203 B.n1029 B.n6 585
R204 B.n885 B.n5 585
R205 B.n1030 B.n5 585
R206 B.n884 B.n883 585
R207 B.n883 B.n4 585
R208 B.n882 B.n374 585
R209 B.n882 B.n881 585
R210 B.n872 B.n375 585
R211 B.n376 B.n375 585
R212 B.n874 B.n873 585
R213 B.n875 B.n874 585
R214 B.n871 B.n381 585
R215 B.n381 B.n380 585
R216 B.n870 B.n869 585
R217 B.n869 B.n868 585
R218 B.n383 B.n382 585
R219 B.n384 B.n383 585
R220 B.n861 B.n860 585
R221 B.n862 B.n861 585
R222 B.n859 B.n389 585
R223 B.n389 B.n388 585
R224 B.n858 B.n857 585
R225 B.n857 B.n856 585
R226 B.n391 B.n390 585
R227 B.n392 B.n391 585
R228 B.n849 B.n848 585
R229 B.n850 B.n849 585
R230 B.n847 B.n397 585
R231 B.n397 B.n396 585
R232 B.n846 B.n845 585
R233 B.n845 B.n844 585
R234 B.n399 B.n398 585
R235 B.n837 B.n399 585
R236 B.n836 B.n835 585
R237 B.n838 B.n836 585
R238 B.n834 B.n404 585
R239 B.n404 B.n403 585
R240 B.n833 B.n832 585
R241 B.n832 B.n831 585
R242 B.n406 B.n405 585
R243 B.n407 B.n406 585
R244 B.n824 B.n823 585
R245 B.n825 B.n824 585
R246 B.n822 B.n412 585
R247 B.n412 B.n411 585
R248 B.n821 B.n820 585
R249 B.n820 B.n819 585
R250 B.n414 B.n413 585
R251 B.n415 B.n414 585
R252 B.n812 B.n811 585
R253 B.n813 B.n812 585
R254 B.n810 B.n420 585
R255 B.n420 B.n419 585
R256 B.n809 B.n808 585
R257 B.n808 B.n807 585
R258 B.n422 B.n421 585
R259 B.n423 B.n422 585
R260 B.n800 B.n799 585
R261 B.n801 B.n800 585
R262 B.n798 B.n428 585
R263 B.n428 B.n427 585
R264 B.n797 B.n796 585
R265 B.n796 B.n795 585
R266 B.n430 B.n429 585
R267 B.n431 B.n430 585
R268 B.n788 B.n787 585
R269 B.n789 B.n788 585
R270 B.n786 B.n436 585
R271 B.n436 B.n435 585
R272 B.n785 B.n784 585
R273 B.n784 B.n783 585
R274 B.n438 B.n437 585
R275 B.n439 B.n438 585
R276 B.n776 B.n775 585
R277 B.n777 B.n776 585
R278 B.n774 B.n444 585
R279 B.n444 B.n443 585
R280 B.n773 B.n772 585
R281 B.n772 B.n771 585
R282 B.n446 B.n445 585
R283 B.n447 B.n446 585
R284 B.n764 B.n763 585
R285 B.n765 B.n764 585
R286 B.n762 B.n452 585
R287 B.n452 B.n451 585
R288 B.n761 B.n760 585
R289 B.n760 B.n759 585
R290 B.n454 B.n453 585
R291 B.n455 B.n454 585
R292 B.n755 B.n754 585
R293 B.n458 B.n457 585
R294 B.n751 B.n750 585
R295 B.n752 B.n751 585
R296 B.n749 B.n516 585
R297 B.n748 B.n747 585
R298 B.n746 B.n745 585
R299 B.n744 B.n743 585
R300 B.n742 B.n741 585
R301 B.n740 B.n739 585
R302 B.n738 B.n737 585
R303 B.n736 B.n735 585
R304 B.n734 B.n733 585
R305 B.n732 B.n731 585
R306 B.n730 B.n729 585
R307 B.n728 B.n727 585
R308 B.n726 B.n725 585
R309 B.n724 B.n723 585
R310 B.n722 B.n721 585
R311 B.n720 B.n719 585
R312 B.n718 B.n717 585
R313 B.n716 B.n715 585
R314 B.n714 B.n713 585
R315 B.n712 B.n711 585
R316 B.n710 B.n709 585
R317 B.n708 B.n707 585
R318 B.n706 B.n705 585
R319 B.n704 B.n703 585
R320 B.n702 B.n701 585
R321 B.n700 B.n699 585
R322 B.n698 B.n697 585
R323 B.n696 B.n695 585
R324 B.n694 B.n693 585
R325 B.n692 B.n691 585
R326 B.n690 B.n689 585
R327 B.n688 B.n687 585
R328 B.n686 B.n685 585
R329 B.n684 B.n683 585
R330 B.n682 B.n681 585
R331 B.n680 B.n679 585
R332 B.n678 B.n677 585
R333 B.n676 B.n675 585
R334 B.n674 B.n673 585
R335 B.n672 B.n671 585
R336 B.n670 B.n669 585
R337 B.n668 B.n667 585
R338 B.n666 B.n665 585
R339 B.n664 B.n663 585
R340 B.n662 B.n661 585
R341 B.n660 B.n659 585
R342 B.n658 B.n657 585
R343 B.n656 B.n655 585
R344 B.n654 B.n653 585
R345 B.n652 B.n651 585
R346 B.n650 B.n649 585
R347 B.n647 B.n646 585
R348 B.n645 B.n644 585
R349 B.n643 B.n642 585
R350 B.n641 B.n640 585
R351 B.n639 B.n638 585
R352 B.n637 B.n636 585
R353 B.n635 B.n634 585
R354 B.n633 B.n632 585
R355 B.n631 B.n630 585
R356 B.n629 B.n628 585
R357 B.n627 B.n626 585
R358 B.n625 B.n624 585
R359 B.n623 B.n622 585
R360 B.n621 B.n620 585
R361 B.n619 B.n618 585
R362 B.n617 B.n616 585
R363 B.n615 B.n614 585
R364 B.n613 B.n612 585
R365 B.n611 B.n610 585
R366 B.n609 B.n608 585
R367 B.n607 B.n606 585
R368 B.n605 B.n604 585
R369 B.n603 B.n602 585
R370 B.n601 B.n600 585
R371 B.n599 B.n598 585
R372 B.n597 B.n596 585
R373 B.n595 B.n594 585
R374 B.n593 B.n592 585
R375 B.n591 B.n590 585
R376 B.n589 B.n588 585
R377 B.n587 B.n586 585
R378 B.n585 B.n584 585
R379 B.n583 B.n582 585
R380 B.n581 B.n580 585
R381 B.n579 B.n578 585
R382 B.n577 B.n576 585
R383 B.n575 B.n574 585
R384 B.n573 B.n572 585
R385 B.n571 B.n570 585
R386 B.n569 B.n568 585
R387 B.n567 B.n566 585
R388 B.n565 B.n564 585
R389 B.n563 B.n562 585
R390 B.n561 B.n560 585
R391 B.n559 B.n558 585
R392 B.n557 B.n556 585
R393 B.n555 B.n554 585
R394 B.n553 B.n552 585
R395 B.n551 B.n550 585
R396 B.n549 B.n548 585
R397 B.n547 B.n546 585
R398 B.n545 B.n544 585
R399 B.n543 B.n542 585
R400 B.n541 B.n540 585
R401 B.n539 B.n538 585
R402 B.n537 B.n536 585
R403 B.n535 B.n534 585
R404 B.n533 B.n532 585
R405 B.n531 B.n530 585
R406 B.n529 B.n528 585
R407 B.n527 B.n526 585
R408 B.n525 B.n524 585
R409 B.n523 B.n522 585
R410 B.n756 B.n456 585
R411 B.n456 B.n455 585
R412 B.n758 B.n757 585
R413 B.n759 B.n758 585
R414 B.n450 B.n449 585
R415 B.n451 B.n450 585
R416 B.n767 B.n766 585
R417 B.n766 B.n765 585
R418 B.n768 B.n448 585
R419 B.n448 B.n447 585
R420 B.n770 B.n769 585
R421 B.n771 B.n770 585
R422 B.n442 B.n441 585
R423 B.n443 B.n442 585
R424 B.n779 B.n778 585
R425 B.n778 B.n777 585
R426 B.n780 B.n440 585
R427 B.n440 B.n439 585
R428 B.n782 B.n781 585
R429 B.n783 B.n782 585
R430 B.n434 B.n433 585
R431 B.n435 B.n434 585
R432 B.n791 B.n790 585
R433 B.n790 B.n789 585
R434 B.n792 B.n432 585
R435 B.n432 B.n431 585
R436 B.n794 B.n793 585
R437 B.n795 B.n794 585
R438 B.n426 B.n425 585
R439 B.n427 B.n426 585
R440 B.n803 B.n802 585
R441 B.n802 B.n801 585
R442 B.n804 B.n424 585
R443 B.n424 B.n423 585
R444 B.n806 B.n805 585
R445 B.n807 B.n806 585
R446 B.n418 B.n417 585
R447 B.n419 B.n418 585
R448 B.n815 B.n814 585
R449 B.n814 B.n813 585
R450 B.n816 B.n416 585
R451 B.n416 B.n415 585
R452 B.n818 B.n817 585
R453 B.n819 B.n818 585
R454 B.n410 B.n409 585
R455 B.n411 B.n410 585
R456 B.n827 B.n826 585
R457 B.n826 B.n825 585
R458 B.n828 B.n408 585
R459 B.n408 B.n407 585
R460 B.n830 B.n829 585
R461 B.n831 B.n830 585
R462 B.n402 B.n401 585
R463 B.n403 B.n402 585
R464 B.n840 B.n839 585
R465 B.n839 B.n838 585
R466 B.n841 B.n400 585
R467 B.n837 B.n400 585
R468 B.n843 B.n842 585
R469 B.n844 B.n843 585
R470 B.n395 B.n394 585
R471 B.n396 B.n395 585
R472 B.n852 B.n851 585
R473 B.n851 B.n850 585
R474 B.n853 B.n393 585
R475 B.n393 B.n392 585
R476 B.n855 B.n854 585
R477 B.n856 B.n855 585
R478 B.n387 B.n386 585
R479 B.n388 B.n387 585
R480 B.n864 B.n863 585
R481 B.n863 B.n862 585
R482 B.n865 B.n385 585
R483 B.n385 B.n384 585
R484 B.n867 B.n866 585
R485 B.n868 B.n867 585
R486 B.n379 B.n378 585
R487 B.n380 B.n379 585
R488 B.n877 B.n876 585
R489 B.n876 B.n875 585
R490 B.n878 B.n377 585
R491 B.n377 B.n376 585
R492 B.n880 B.n879 585
R493 B.n881 B.n880 585
R494 B.n2 B.n0 585
R495 B.n4 B.n2 585
R496 B.n3 B.n1 585
R497 B.n1029 B.n3 585
R498 B.n1027 B.n1026 585
R499 B.n1028 B.n1027 585
R500 B.n1025 B.n9 585
R501 B.n9 B.n8 585
R502 B.n1024 B.n1023 585
R503 B.n1023 B.n1022 585
R504 B.n11 B.n10 585
R505 B.n1021 B.n11 585
R506 B.n1019 B.n1018 585
R507 B.n1020 B.n1019 585
R508 B.n1017 B.n16 585
R509 B.n16 B.n15 585
R510 B.n1016 B.n1015 585
R511 B.n1015 B.n1014 585
R512 B.n18 B.n17 585
R513 B.n1013 B.n18 585
R514 B.n1011 B.n1010 585
R515 B.n1012 B.n1011 585
R516 B.n1009 B.n23 585
R517 B.n23 B.n22 585
R518 B.n1008 B.n1007 585
R519 B.n1007 B.n1006 585
R520 B.n25 B.n24 585
R521 B.n1005 B.n25 585
R522 B.n1003 B.n1002 585
R523 B.n1004 B.n1003 585
R524 B.n1001 B.n29 585
R525 B.n32 B.n29 585
R526 B.n1000 B.n999 585
R527 B.n999 B.n998 585
R528 B.n31 B.n30 585
R529 B.n997 B.n31 585
R530 B.n995 B.n994 585
R531 B.n996 B.n995 585
R532 B.n993 B.n37 585
R533 B.n37 B.n36 585
R534 B.n992 B.n991 585
R535 B.n991 B.n990 585
R536 B.n39 B.n38 585
R537 B.n989 B.n39 585
R538 B.n987 B.n986 585
R539 B.n988 B.n987 585
R540 B.n985 B.n44 585
R541 B.n44 B.n43 585
R542 B.n984 B.n983 585
R543 B.n983 B.n982 585
R544 B.n46 B.n45 585
R545 B.n981 B.n46 585
R546 B.n979 B.n978 585
R547 B.n980 B.n979 585
R548 B.n977 B.n51 585
R549 B.n51 B.n50 585
R550 B.n976 B.n975 585
R551 B.n975 B.n974 585
R552 B.n53 B.n52 585
R553 B.n973 B.n53 585
R554 B.n971 B.n970 585
R555 B.n972 B.n971 585
R556 B.n969 B.n58 585
R557 B.n58 B.n57 585
R558 B.n968 B.n967 585
R559 B.n967 B.n966 585
R560 B.n60 B.n59 585
R561 B.n965 B.n60 585
R562 B.n963 B.n962 585
R563 B.n964 B.n963 585
R564 B.n961 B.n65 585
R565 B.n65 B.n64 585
R566 B.n960 B.n959 585
R567 B.n959 B.n958 585
R568 B.n67 B.n66 585
R569 B.n957 B.n67 585
R570 B.n955 B.n954 585
R571 B.n956 B.n955 585
R572 B.n953 B.n72 585
R573 B.n72 B.n71 585
R574 B.n952 B.n951 585
R575 B.n951 B.n950 585
R576 B.n74 B.n73 585
R577 B.n949 B.n74 585
R578 B.n947 B.n946 585
R579 B.n948 B.n947 585
R580 B.n945 B.n79 585
R581 B.n79 B.n78 585
R582 B.n1032 B.n1031 585
R583 B.n1031 B.n1030 585
R584 B.n754 B.n456 550.159
R585 B.n943 B.n79 550.159
R586 B.n522 B.n454 550.159
R587 B.n940 B.n140 550.159
R588 B.n519 B.t16 411.628
R589 B.n141 B.t12 411.628
R590 B.n517 B.t9 411.628
R591 B.n143 B.t18 411.628
R592 B.n519 B.t14 355.086
R593 B.n517 B.t6 355.086
R594 B.n143 B.t17 355.086
R595 B.n141 B.t10 355.086
R596 B.n520 B.t15 353.834
R597 B.n142 B.t13 353.834
R598 B.n518 B.t8 353.834
R599 B.n144 B.t19 353.834
R600 B.n941 B.n138 256.663
R601 B.n941 B.n137 256.663
R602 B.n941 B.n136 256.663
R603 B.n941 B.n135 256.663
R604 B.n941 B.n134 256.663
R605 B.n941 B.n133 256.663
R606 B.n941 B.n132 256.663
R607 B.n941 B.n131 256.663
R608 B.n941 B.n130 256.663
R609 B.n941 B.n129 256.663
R610 B.n941 B.n128 256.663
R611 B.n941 B.n127 256.663
R612 B.n941 B.n126 256.663
R613 B.n941 B.n125 256.663
R614 B.n941 B.n124 256.663
R615 B.n941 B.n123 256.663
R616 B.n941 B.n122 256.663
R617 B.n941 B.n121 256.663
R618 B.n941 B.n120 256.663
R619 B.n941 B.n119 256.663
R620 B.n941 B.n118 256.663
R621 B.n941 B.n117 256.663
R622 B.n941 B.n116 256.663
R623 B.n941 B.n115 256.663
R624 B.n941 B.n114 256.663
R625 B.n941 B.n113 256.663
R626 B.n941 B.n112 256.663
R627 B.n941 B.n111 256.663
R628 B.n941 B.n110 256.663
R629 B.n941 B.n109 256.663
R630 B.n941 B.n108 256.663
R631 B.n941 B.n107 256.663
R632 B.n941 B.n106 256.663
R633 B.n941 B.n105 256.663
R634 B.n941 B.n104 256.663
R635 B.n941 B.n103 256.663
R636 B.n941 B.n102 256.663
R637 B.n941 B.n101 256.663
R638 B.n941 B.n100 256.663
R639 B.n941 B.n99 256.663
R640 B.n941 B.n98 256.663
R641 B.n941 B.n97 256.663
R642 B.n941 B.n96 256.663
R643 B.n941 B.n95 256.663
R644 B.n941 B.n94 256.663
R645 B.n941 B.n93 256.663
R646 B.n941 B.n92 256.663
R647 B.n941 B.n91 256.663
R648 B.n941 B.n90 256.663
R649 B.n941 B.n89 256.663
R650 B.n941 B.n88 256.663
R651 B.n941 B.n87 256.663
R652 B.n941 B.n86 256.663
R653 B.n941 B.n85 256.663
R654 B.n941 B.n84 256.663
R655 B.n941 B.n83 256.663
R656 B.n941 B.n82 256.663
R657 B.n942 B.n941 256.663
R658 B.n753 B.n752 256.663
R659 B.n752 B.n459 256.663
R660 B.n752 B.n460 256.663
R661 B.n752 B.n461 256.663
R662 B.n752 B.n462 256.663
R663 B.n752 B.n463 256.663
R664 B.n752 B.n464 256.663
R665 B.n752 B.n465 256.663
R666 B.n752 B.n466 256.663
R667 B.n752 B.n467 256.663
R668 B.n752 B.n468 256.663
R669 B.n752 B.n469 256.663
R670 B.n752 B.n470 256.663
R671 B.n752 B.n471 256.663
R672 B.n752 B.n472 256.663
R673 B.n752 B.n473 256.663
R674 B.n752 B.n474 256.663
R675 B.n752 B.n475 256.663
R676 B.n752 B.n476 256.663
R677 B.n752 B.n477 256.663
R678 B.n752 B.n478 256.663
R679 B.n752 B.n479 256.663
R680 B.n752 B.n480 256.663
R681 B.n752 B.n481 256.663
R682 B.n752 B.n482 256.663
R683 B.n752 B.n483 256.663
R684 B.n752 B.n484 256.663
R685 B.n752 B.n485 256.663
R686 B.n752 B.n486 256.663
R687 B.n752 B.n487 256.663
R688 B.n752 B.n488 256.663
R689 B.n752 B.n489 256.663
R690 B.n752 B.n490 256.663
R691 B.n752 B.n491 256.663
R692 B.n752 B.n492 256.663
R693 B.n752 B.n493 256.663
R694 B.n752 B.n494 256.663
R695 B.n752 B.n495 256.663
R696 B.n752 B.n496 256.663
R697 B.n752 B.n497 256.663
R698 B.n752 B.n498 256.663
R699 B.n752 B.n499 256.663
R700 B.n752 B.n500 256.663
R701 B.n752 B.n501 256.663
R702 B.n752 B.n502 256.663
R703 B.n752 B.n503 256.663
R704 B.n752 B.n504 256.663
R705 B.n752 B.n505 256.663
R706 B.n752 B.n506 256.663
R707 B.n752 B.n507 256.663
R708 B.n752 B.n508 256.663
R709 B.n752 B.n509 256.663
R710 B.n752 B.n510 256.663
R711 B.n752 B.n511 256.663
R712 B.n752 B.n512 256.663
R713 B.n752 B.n513 256.663
R714 B.n752 B.n514 256.663
R715 B.n752 B.n515 256.663
R716 B.n758 B.n456 163.367
R717 B.n758 B.n450 163.367
R718 B.n766 B.n450 163.367
R719 B.n766 B.n448 163.367
R720 B.n770 B.n448 163.367
R721 B.n770 B.n442 163.367
R722 B.n778 B.n442 163.367
R723 B.n778 B.n440 163.367
R724 B.n782 B.n440 163.367
R725 B.n782 B.n434 163.367
R726 B.n790 B.n434 163.367
R727 B.n790 B.n432 163.367
R728 B.n794 B.n432 163.367
R729 B.n794 B.n426 163.367
R730 B.n802 B.n426 163.367
R731 B.n802 B.n424 163.367
R732 B.n806 B.n424 163.367
R733 B.n806 B.n418 163.367
R734 B.n814 B.n418 163.367
R735 B.n814 B.n416 163.367
R736 B.n818 B.n416 163.367
R737 B.n818 B.n410 163.367
R738 B.n826 B.n410 163.367
R739 B.n826 B.n408 163.367
R740 B.n830 B.n408 163.367
R741 B.n830 B.n402 163.367
R742 B.n839 B.n402 163.367
R743 B.n839 B.n400 163.367
R744 B.n843 B.n400 163.367
R745 B.n843 B.n395 163.367
R746 B.n851 B.n395 163.367
R747 B.n851 B.n393 163.367
R748 B.n855 B.n393 163.367
R749 B.n855 B.n387 163.367
R750 B.n863 B.n387 163.367
R751 B.n863 B.n385 163.367
R752 B.n867 B.n385 163.367
R753 B.n867 B.n379 163.367
R754 B.n876 B.n379 163.367
R755 B.n876 B.n377 163.367
R756 B.n880 B.n377 163.367
R757 B.n880 B.n2 163.367
R758 B.n1031 B.n2 163.367
R759 B.n1031 B.n3 163.367
R760 B.n1027 B.n3 163.367
R761 B.n1027 B.n9 163.367
R762 B.n1023 B.n9 163.367
R763 B.n1023 B.n11 163.367
R764 B.n1019 B.n11 163.367
R765 B.n1019 B.n16 163.367
R766 B.n1015 B.n16 163.367
R767 B.n1015 B.n18 163.367
R768 B.n1011 B.n18 163.367
R769 B.n1011 B.n23 163.367
R770 B.n1007 B.n23 163.367
R771 B.n1007 B.n25 163.367
R772 B.n1003 B.n25 163.367
R773 B.n1003 B.n29 163.367
R774 B.n999 B.n29 163.367
R775 B.n999 B.n31 163.367
R776 B.n995 B.n31 163.367
R777 B.n995 B.n37 163.367
R778 B.n991 B.n37 163.367
R779 B.n991 B.n39 163.367
R780 B.n987 B.n39 163.367
R781 B.n987 B.n44 163.367
R782 B.n983 B.n44 163.367
R783 B.n983 B.n46 163.367
R784 B.n979 B.n46 163.367
R785 B.n979 B.n51 163.367
R786 B.n975 B.n51 163.367
R787 B.n975 B.n53 163.367
R788 B.n971 B.n53 163.367
R789 B.n971 B.n58 163.367
R790 B.n967 B.n58 163.367
R791 B.n967 B.n60 163.367
R792 B.n963 B.n60 163.367
R793 B.n963 B.n65 163.367
R794 B.n959 B.n65 163.367
R795 B.n959 B.n67 163.367
R796 B.n955 B.n67 163.367
R797 B.n955 B.n72 163.367
R798 B.n951 B.n72 163.367
R799 B.n951 B.n74 163.367
R800 B.n947 B.n74 163.367
R801 B.n947 B.n79 163.367
R802 B.n751 B.n458 163.367
R803 B.n751 B.n516 163.367
R804 B.n747 B.n746 163.367
R805 B.n743 B.n742 163.367
R806 B.n739 B.n738 163.367
R807 B.n735 B.n734 163.367
R808 B.n731 B.n730 163.367
R809 B.n727 B.n726 163.367
R810 B.n723 B.n722 163.367
R811 B.n719 B.n718 163.367
R812 B.n715 B.n714 163.367
R813 B.n711 B.n710 163.367
R814 B.n707 B.n706 163.367
R815 B.n703 B.n702 163.367
R816 B.n699 B.n698 163.367
R817 B.n695 B.n694 163.367
R818 B.n691 B.n690 163.367
R819 B.n687 B.n686 163.367
R820 B.n683 B.n682 163.367
R821 B.n679 B.n678 163.367
R822 B.n675 B.n674 163.367
R823 B.n671 B.n670 163.367
R824 B.n667 B.n666 163.367
R825 B.n663 B.n662 163.367
R826 B.n659 B.n658 163.367
R827 B.n655 B.n654 163.367
R828 B.n651 B.n650 163.367
R829 B.n646 B.n645 163.367
R830 B.n642 B.n641 163.367
R831 B.n638 B.n637 163.367
R832 B.n634 B.n633 163.367
R833 B.n630 B.n629 163.367
R834 B.n626 B.n625 163.367
R835 B.n622 B.n621 163.367
R836 B.n618 B.n617 163.367
R837 B.n614 B.n613 163.367
R838 B.n610 B.n609 163.367
R839 B.n606 B.n605 163.367
R840 B.n602 B.n601 163.367
R841 B.n598 B.n597 163.367
R842 B.n594 B.n593 163.367
R843 B.n590 B.n589 163.367
R844 B.n586 B.n585 163.367
R845 B.n582 B.n581 163.367
R846 B.n578 B.n577 163.367
R847 B.n574 B.n573 163.367
R848 B.n570 B.n569 163.367
R849 B.n566 B.n565 163.367
R850 B.n562 B.n561 163.367
R851 B.n558 B.n557 163.367
R852 B.n554 B.n553 163.367
R853 B.n550 B.n549 163.367
R854 B.n546 B.n545 163.367
R855 B.n542 B.n541 163.367
R856 B.n538 B.n537 163.367
R857 B.n534 B.n533 163.367
R858 B.n530 B.n529 163.367
R859 B.n526 B.n525 163.367
R860 B.n760 B.n454 163.367
R861 B.n760 B.n452 163.367
R862 B.n764 B.n452 163.367
R863 B.n764 B.n446 163.367
R864 B.n772 B.n446 163.367
R865 B.n772 B.n444 163.367
R866 B.n776 B.n444 163.367
R867 B.n776 B.n438 163.367
R868 B.n784 B.n438 163.367
R869 B.n784 B.n436 163.367
R870 B.n788 B.n436 163.367
R871 B.n788 B.n430 163.367
R872 B.n796 B.n430 163.367
R873 B.n796 B.n428 163.367
R874 B.n800 B.n428 163.367
R875 B.n800 B.n422 163.367
R876 B.n808 B.n422 163.367
R877 B.n808 B.n420 163.367
R878 B.n812 B.n420 163.367
R879 B.n812 B.n414 163.367
R880 B.n820 B.n414 163.367
R881 B.n820 B.n412 163.367
R882 B.n824 B.n412 163.367
R883 B.n824 B.n406 163.367
R884 B.n832 B.n406 163.367
R885 B.n832 B.n404 163.367
R886 B.n836 B.n404 163.367
R887 B.n836 B.n399 163.367
R888 B.n845 B.n399 163.367
R889 B.n845 B.n397 163.367
R890 B.n849 B.n397 163.367
R891 B.n849 B.n391 163.367
R892 B.n857 B.n391 163.367
R893 B.n857 B.n389 163.367
R894 B.n861 B.n389 163.367
R895 B.n861 B.n383 163.367
R896 B.n869 B.n383 163.367
R897 B.n869 B.n381 163.367
R898 B.n874 B.n381 163.367
R899 B.n874 B.n375 163.367
R900 B.n882 B.n375 163.367
R901 B.n883 B.n882 163.367
R902 B.n883 B.n5 163.367
R903 B.n6 B.n5 163.367
R904 B.n7 B.n6 163.367
R905 B.n888 B.n7 163.367
R906 B.n888 B.n12 163.367
R907 B.n13 B.n12 163.367
R908 B.n14 B.n13 163.367
R909 B.n893 B.n14 163.367
R910 B.n893 B.n19 163.367
R911 B.n20 B.n19 163.367
R912 B.n21 B.n20 163.367
R913 B.n898 B.n21 163.367
R914 B.n898 B.n26 163.367
R915 B.n27 B.n26 163.367
R916 B.n28 B.n27 163.367
R917 B.n903 B.n28 163.367
R918 B.n903 B.n33 163.367
R919 B.n34 B.n33 163.367
R920 B.n35 B.n34 163.367
R921 B.n908 B.n35 163.367
R922 B.n908 B.n40 163.367
R923 B.n41 B.n40 163.367
R924 B.n42 B.n41 163.367
R925 B.n913 B.n42 163.367
R926 B.n913 B.n47 163.367
R927 B.n48 B.n47 163.367
R928 B.n49 B.n48 163.367
R929 B.n918 B.n49 163.367
R930 B.n918 B.n54 163.367
R931 B.n55 B.n54 163.367
R932 B.n56 B.n55 163.367
R933 B.n923 B.n56 163.367
R934 B.n923 B.n61 163.367
R935 B.n62 B.n61 163.367
R936 B.n63 B.n62 163.367
R937 B.n928 B.n63 163.367
R938 B.n928 B.n68 163.367
R939 B.n69 B.n68 163.367
R940 B.n70 B.n69 163.367
R941 B.n933 B.n70 163.367
R942 B.n933 B.n75 163.367
R943 B.n76 B.n75 163.367
R944 B.n77 B.n76 163.367
R945 B.n140 B.n77 163.367
R946 B.n146 B.n81 163.367
R947 B.n150 B.n149 163.367
R948 B.n154 B.n153 163.367
R949 B.n158 B.n157 163.367
R950 B.n162 B.n161 163.367
R951 B.n166 B.n165 163.367
R952 B.n170 B.n169 163.367
R953 B.n174 B.n173 163.367
R954 B.n178 B.n177 163.367
R955 B.n182 B.n181 163.367
R956 B.n186 B.n185 163.367
R957 B.n190 B.n189 163.367
R958 B.n194 B.n193 163.367
R959 B.n198 B.n197 163.367
R960 B.n202 B.n201 163.367
R961 B.n206 B.n205 163.367
R962 B.n210 B.n209 163.367
R963 B.n214 B.n213 163.367
R964 B.n218 B.n217 163.367
R965 B.n222 B.n221 163.367
R966 B.n226 B.n225 163.367
R967 B.n230 B.n229 163.367
R968 B.n234 B.n233 163.367
R969 B.n238 B.n237 163.367
R970 B.n242 B.n241 163.367
R971 B.n246 B.n245 163.367
R972 B.n250 B.n249 163.367
R973 B.n254 B.n253 163.367
R974 B.n258 B.n257 163.367
R975 B.n262 B.n261 163.367
R976 B.n266 B.n265 163.367
R977 B.n271 B.n270 163.367
R978 B.n275 B.n274 163.367
R979 B.n279 B.n278 163.367
R980 B.n283 B.n282 163.367
R981 B.n287 B.n286 163.367
R982 B.n291 B.n290 163.367
R983 B.n295 B.n294 163.367
R984 B.n299 B.n298 163.367
R985 B.n303 B.n302 163.367
R986 B.n307 B.n306 163.367
R987 B.n311 B.n310 163.367
R988 B.n315 B.n314 163.367
R989 B.n319 B.n318 163.367
R990 B.n323 B.n322 163.367
R991 B.n327 B.n326 163.367
R992 B.n331 B.n330 163.367
R993 B.n335 B.n334 163.367
R994 B.n339 B.n338 163.367
R995 B.n343 B.n342 163.367
R996 B.n347 B.n346 163.367
R997 B.n351 B.n350 163.367
R998 B.n355 B.n354 163.367
R999 B.n359 B.n358 163.367
R1000 B.n363 B.n362 163.367
R1001 B.n367 B.n366 163.367
R1002 B.n371 B.n370 163.367
R1003 B.n940 B.n139 163.367
R1004 B.n754 B.n753 71.676
R1005 B.n516 B.n459 71.676
R1006 B.n746 B.n460 71.676
R1007 B.n742 B.n461 71.676
R1008 B.n738 B.n462 71.676
R1009 B.n734 B.n463 71.676
R1010 B.n730 B.n464 71.676
R1011 B.n726 B.n465 71.676
R1012 B.n722 B.n466 71.676
R1013 B.n718 B.n467 71.676
R1014 B.n714 B.n468 71.676
R1015 B.n710 B.n469 71.676
R1016 B.n706 B.n470 71.676
R1017 B.n702 B.n471 71.676
R1018 B.n698 B.n472 71.676
R1019 B.n694 B.n473 71.676
R1020 B.n690 B.n474 71.676
R1021 B.n686 B.n475 71.676
R1022 B.n682 B.n476 71.676
R1023 B.n678 B.n477 71.676
R1024 B.n674 B.n478 71.676
R1025 B.n670 B.n479 71.676
R1026 B.n666 B.n480 71.676
R1027 B.n662 B.n481 71.676
R1028 B.n658 B.n482 71.676
R1029 B.n654 B.n483 71.676
R1030 B.n650 B.n484 71.676
R1031 B.n645 B.n485 71.676
R1032 B.n641 B.n486 71.676
R1033 B.n637 B.n487 71.676
R1034 B.n633 B.n488 71.676
R1035 B.n629 B.n489 71.676
R1036 B.n625 B.n490 71.676
R1037 B.n621 B.n491 71.676
R1038 B.n617 B.n492 71.676
R1039 B.n613 B.n493 71.676
R1040 B.n609 B.n494 71.676
R1041 B.n605 B.n495 71.676
R1042 B.n601 B.n496 71.676
R1043 B.n597 B.n497 71.676
R1044 B.n593 B.n498 71.676
R1045 B.n589 B.n499 71.676
R1046 B.n585 B.n500 71.676
R1047 B.n581 B.n501 71.676
R1048 B.n577 B.n502 71.676
R1049 B.n573 B.n503 71.676
R1050 B.n569 B.n504 71.676
R1051 B.n565 B.n505 71.676
R1052 B.n561 B.n506 71.676
R1053 B.n557 B.n507 71.676
R1054 B.n553 B.n508 71.676
R1055 B.n549 B.n509 71.676
R1056 B.n545 B.n510 71.676
R1057 B.n541 B.n511 71.676
R1058 B.n537 B.n512 71.676
R1059 B.n533 B.n513 71.676
R1060 B.n529 B.n514 71.676
R1061 B.n525 B.n515 71.676
R1062 B.n943 B.n942 71.676
R1063 B.n146 B.n82 71.676
R1064 B.n150 B.n83 71.676
R1065 B.n154 B.n84 71.676
R1066 B.n158 B.n85 71.676
R1067 B.n162 B.n86 71.676
R1068 B.n166 B.n87 71.676
R1069 B.n170 B.n88 71.676
R1070 B.n174 B.n89 71.676
R1071 B.n178 B.n90 71.676
R1072 B.n182 B.n91 71.676
R1073 B.n186 B.n92 71.676
R1074 B.n190 B.n93 71.676
R1075 B.n194 B.n94 71.676
R1076 B.n198 B.n95 71.676
R1077 B.n202 B.n96 71.676
R1078 B.n206 B.n97 71.676
R1079 B.n210 B.n98 71.676
R1080 B.n214 B.n99 71.676
R1081 B.n218 B.n100 71.676
R1082 B.n222 B.n101 71.676
R1083 B.n226 B.n102 71.676
R1084 B.n230 B.n103 71.676
R1085 B.n234 B.n104 71.676
R1086 B.n238 B.n105 71.676
R1087 B.n242 B.n106 71.676
R1088 B.n246 B.n107 71.676
R1089 B.n250 B.n108 71.676
R1090 B.n254 B.n109 71.676
R1091 B.n258 B.n110 71.676
R1092 B.n262 B.n111 71.676
R1093 B.n266 B.n112 71.676
R1094 B.n271 B.n113 71.676
R1095 B.n275 B.n114 71.676
R1096 B.n279 B.n115 71.676
R1097 B.n283 B.n116 71.676
R1098 B.n287 B.n117 71.676
R1099 B.n291 B.n118 71.676
R1100 B.n295 B.n119 71.676
R1101 B.n299 B.n120 71.676
R1102 B.n303 B.n121 71.676
R1103 B.n307 B.n122 71.676
R1104 B.n311 B.n123 71.676
R1105 B.n315 B.n124 71.676
R1106 B.n319 B.n125 71.676
R1107 B.n323 B.n126 71.676
R1108 B.n327 B.n127 71.676
R1109 B.n331 B.n128 71.676
R1110 B.n335 B.n129 71.676
R1111 B.n339 B.n130 71.676
R1112 B.n343 B.n131 71.676
R1113 B.n347 B.n132 71.676
R1114 B.n351 B.n133 71.676
R1115 B.n355 B.n134 71.676
R1116 B.n359 B.n135 71.676
R1117 B.n363 B.n136 71.676
R1118 B.n367 B.n137 71.676
R1119 B.n371 B.n138 71.676
R1120 B.n139 B.n138 71.676
R1121 B.n370 B.n137 71.676
R1122 B.n366 B.n136 71.676
R1123 B.n362 B.n135 71.676
R1124 B.n358 B.n134 71.676
R1125 B.n354 B.n133 71.676
R1126 B.n350 B.n132 71.676
R1127 B.n346 B.n131 71.676
R1128 B.n342 B.n130 71.676
R1129 B.n338 B.n129 71.676
R1130 B.n334 B.n128 71.676
R1131 B.n330 B.n127 71.676
R1132 B.n326 B.n126 71.676
R1133 B.n322 B.n125 71.676
R1134 B.n318 B.n124 71.676
R1135 B.n314 B.n123 71.676
R1136 B.n310 B.n122 71.676
R1137 B.n306 B.n121 71.676
R1138 B.n302 B.n120 71.676
R1139 B.n298 B.n119 71.676
R1140 B.n294 B.n118 71.676
R1141 B.n290 B.n117 71.676
R1142 B.n286 B.n116 71.676
R1143 B.n282 B.n115 71.676
R1144 B.n278 B.n114 71.676
R1145 B.n274 B.n113 71.676
R1146 B.n270 B.n112 71.676
R1147 B.n265 B.n111 71.676
R1148 B.n261 B.n110 71.676
R1149 B.n257 B.n109 71.676
R1150 B.n253 B.n108 71.676
R1151 B.n249 B.n107 71.676
R1152 B.n245 B.n106 71.676
R1153 B.n241 B.n105 71.676
R1154 B.n237 B.n104 71.676
R1155 B.n233 B.n103 71.676
R1156 B.n229 B.n102 71.676
R1157 B.n225 B.n101 71.676
R1158 B.n221 B.n100 71.676
R1159 B.n217 B.n99 71.676
R1160 B.n213 B.n98 71.676
R1161 B.n209 B.n97 71.676
R1162 B.n205 B.n96 71.676
R1163 B.n201 B.n95 71.676
R1164 B.n197 B.n94 71.676
R1165 B.n193 B.n93 71.676
R1166 B.n189 B.n92 71.676
R1167 B.n185 B.n91 71.676
R1168 B.n181 B.n90 71.676
R1169 B.n177 B.n89 71.676
R1170 B.n173 B.n88 71.676
R1171 B.n169 B.n87 71.676
R1172 B.n165 B.n86 71.676
R1173 B.n161 B.n85 71.676
R1174 B.n157 B.n84 71.676
R1175 B.n153 B.n83 71.676
R1176 B.n149 B.n82 71.676
R1177 B.n942 B.n81 71.676
R1178 B.n753 B.n458 71.676
R1179 B.n747 B.n459 71.676
R1180 B.n743 B.n460 71.676
R1181 B.n739 B.n461 71.676
R1182 B.n735 B.n462 71.676
R1183 B.n731 B.n463 71.676
R1184 B.n727 B.n464 71.676
R1185 B.n723 B.n465 71.676
R1186 B.n719 B.n466 71.676
R1187 B.n715 B.n467 71.676
R1188 B.n711 B.n468 71.676
R1189 B.n707 B.n469 71.676
R1190 B.n703 B.n470 71.676
R1191 B.n699 B.n471 71.676
R1192 B.n695 B.n472 71.676
R1193 B.n691 B.n473 71.676
R1194 B.n687 B.n474 71.676
R1195 B.n683 B.n475 71.676
R1196 B.n679 B.n476 71.676
R1197 B.n675 B.n477 71.676
R1198 B.n671 B.n478 71.676
R1199 B.n667 B.n479 71.676
R1200 B.n663 B.n480 71.676
R1201 B.n659 B.n481 71.676
R1202 B.n655 B.n482 71.676
R1203 B.n651 B.n483 71.676
R1204 B.n646 B.n484 71.676
R1205 B.n642 B.n485 71.676
R1206 B.n638 B.n486 71.676
R1207 B.n634 B.n487 71.676
R1208 B.n630 B.n488 71.676
R1209 B.n626 B.n489 71.676
R1210 B.n622 B.n490 71.676
R1211 B.n618 B.n491 71.676
R1212 B.n614 B.n492 71.676
R1213 B.n610 B.n493 71.676
R1214 B.n606 B.n494 71.676
R1215 B.n602 B.n495 71.676
R1216 B.n598 B.n496 71.676
R1217 B.n594 B.n497 71.676
R1218 B.n590 B.n498 71.676
R1219 B.n586 B.n499 71.676
R1220 B.n582 B.n500 71.676
R1221 B.n578 B.n501 71.676
R1222 B.n574 B.n502 71.676
R1223 B.n570 B.n503 71.676
R1224 B.n566 B.n504 71.676
R1225 B.n562 B.n505 71.676
R1226 B.n558 B.n506 71.676
R1227 B.n554 B.n507 71.676
R1228 B.n550 B.n508 71.676
R1229 B.n546 B.n509 71.676
R1230 B.n542 B.n510 71.676
R1231 B.n538 B.n511 71.676
R1232 B.n534 B.n512 71.676
R1233 B.n530 B.n513 71.676
R1234 B.n526 B.n514 71.676
R1235 B.n522 B.n515 71.676
R1236 B.n752 B.n455 69.2797
R1237 B.n941 B.n78 69.2797
R1238 B.n521 B.n520 59.5399
R1239 B.n648 B.n518 59.5399
R1240 B.n145 B.n144 59.5399
R1241 B.n268 B.n142 59.5399
R1242 B.n520 B.n519 57.7944
R1243 B.n518 B.n517 57.7944
R1244 B.n144 B.n143 57.7944
R1245 B.n142 B.n141 57.7944
R1246 B.n945 B.n944 35.7468
R1247 B.n939 B.n938 35.7468
R1248 B.n523 B.n453 35.7468
R1249 B.n756 B.n755 35.7468
R1250 B.n759 B.n455 34.8967
R1251 B.n759 B.n451 34.8967
R1252 B.n765 B.n451 34.8967
R1253 B.n765 B.n447 34.8967
R1254 B.n771 B.n447 34.8967
R1255 B.n771 B.n443 34.8967
R1256 B.n777 B.n443 34.8967
R1257 B.n783 B.n439 34.8967
R1258 B.n783 B.n435 34.8967
R1259 B.n789 B.n435 34.8967
R1260 B.n789 B.n431 34.8967
R1261 B.n795 B.n431 34.8967
R1262 B.n795 B.n427 34.8967
R1263 B.n801 B.n427 34.8967
R1264 B.n801 B.n423 34.8967
R1265 B.n807 B.n423 34.8967
R1266 B.n807 B.n419 34.8967
R1267 B.n813 B.n419 34.8967
R1268 B.n819 B.n415 34.8967
R1269 B.n819 B.n411 34.8967
R1270 B.n825 B.n411 34.8967
R1271 B.n825 B.n407 34.8967
R1272 B.n831 B.n407 34.8967
R1273 B.n831 B.n403 34.8967
R1274 B.n838 B.n403 34.8967
R1275 B.n838 B.n837 34.8967
R1276 B.n844 B.n396 34.8967
R1277 B.n850 B.n396 34.8967
R1278 B.n850 B.n392 34.8967
R1279 B.n856 B.n392 34.8967
R1280 B.n856 B.n388 34.8967
R1281 B.n862 B.n388 34.8967
R1282 B.n862 B.n384 34.8967
R1283 B.n868 B.n384 34.8967
R1284 B.n875 B.n380 34.8967
R1285 B.n875 B.n376 34.8967
R1286 B.n881 B.n376 34.8967
R1287 B.n881 B.n4 34.8967
R1288 B.n1030 B.n4 34.8967
R1289 B.n1030 B.n1029 34.8967
R1290 B.n1029 B.n1028 34.8967
R1291 B.n1028 B.n8 34.8967
R1292 B.n1022 B.n8 34.8967
R1293 B.n1022 B.n1021 34.8967
R1294 B.n1020 B.n15 34.8967
R1295 B.n1014 B.n15 34.8967
R1296 B.n1014 B.n1013 34.8967
R1297 B.n1013 B.n1012 34.8967
R1298 B.n1012 B.n22 34.8967
R1299 B.n1006 B.n22 34.8967
R1300 B.n1006 B.n1005 34.8967
R1301 B.n1005 B.n1004 34.8967
R1302 B.n998 B.n32 34.8967
R1303 B.n998 B.n997 34.8967
R1304 B.n997 B.n996 34.8967
R1305 B.n996 B.n36 34.8967
R1306 B.n990 B.n36 34.8967
R1307 B.n990 B.n989 34.8967
R1308 B.n989 B.n988 34.8967
R1309 B.n988 B.n43 34.8967
R1310 B.n982 B.n981 34.8967
R1311 B.n981 B.n980 34.8967
R1312 B.n980 B.n50 34.8967
R1313 B.n974 B.n50 34.8967
R1314 B.n974 B.n973 34.8967
R1315 B.n973 B.n972 34.8967
R1316 B.n972 B.n57 34.8967
R1317 B.n966 B.n57 34.8967
R1318 B.n966 B.n965 34.8967
R1319 B.n965 B.n964 34.8967
R1320 B.n964 B.n64 34.8967
R1321 B.n958 B.n957 34.8967
R1322 B.n957 B.n956 34.8967
R1323 B.n956 B.n71 34.8967
R1324 B.n950 B.n71 34.8967
R1325 B.n950 B.n949 34.8967
R1326 B.n949 B.n948 34.8967
R1327 B.n948 B.n78 34.8967
R1328 B.t1 B.n380 34.3835
R1329 B.n1021 B.t2 34.3835
R1330 B.n844 B.t4 26.1726
R1331 B.n1004 B.t0 26.1726
R1332 B B.n1032 18.0485
R1333 B.n777 B.t7 17.9618
R1334 B.t5 B.n415 17.9618
R1335 B.t3 B.n43 17.9618
R1336 B.n958 B.t11 17.9618
R1337 B.t7 B.n439 16.9354
R1338 B.n813 B.t5 16.9354
R1339 B.n982 B.t3 16.9354
R1340 B.t11 B.n64 16.9354
R1341 B.n944 B.n80 10.6151
R1342 B.n147 B.n80 10.6151
R1343 B.n148 B.n147 10.6151
R1344 B.n151 B.n148 10.6151
R1345 B.n152 B.n151 10.6151
R1346 B.n155 B.n152 10.6151
R1347 B.n156 B.n155 10.6151
R1348 B.n159 B.n156 10.6151
R1349 B.n160 B.n159 10.6151
R1350 B.n163 B.n160 10.6151
R1351 B.n164 B.n163 10.6151
R1352 B.n167 B.n164 10.6151
R1353 B.n168 B.n167 10.6151
R1354 B.n171 B.n168 10.6151
R1355 B.n172 B.n171 10.6151
R1356 B.n175 B.n172 10.6151
R1357 B.n176 B.n175 10.6151
R1358 B.n179 B.n176 10.6151
R1359 B.n180 B.n179 10.6151
R1360 B.n183 B.n180 10.6151
R1361 B.n184 B.n183 10.6151
R1362 B.n187 B.n184 10.6151
R1363 B.n188 B.n187 10.6151
R1364 B.n191 B.n188 10.6151
R1365 B.n192 B.n191 10.6151
R1366 B.n195 B.n192 10.6151
R1367 B.n196 B.n195 10.6151
R1368 B.n199 B.n196 10.6151
R1369 B.n200 B.n199 10.6151
R1370 B.n203 B.n200 10.6151
R1371 B.n204 B.n203 10.6151
R1372 B.n207 B.n204 10.6151
R1373 B.n208 B.n207 10.6151
R1374 B.n211 B.n208 10.6151
R1375 B.n212 B.n211 10.6151
R1376 B.n215 B.n212 10.6151
R1377 B.n216 B.n215 10.6151
R1378 B.n219 B.n216 10.6151
R1379 B.n220 B.n219 10.6151
R1380 B.n223 B.n220 10.6151
R1381 B.n224 B.n223 10.6151
R1382 B.n227 B.n224 10.6151
R1383 B.n228 B.n227 10.6151
R1384 B.n231 B.n228 10.6151
R1385 B.n232 B.n231 10.6151
R1386 B.n235 B.n232 10.6151
R1387 B.n236 B.n235 10.6151
R1388 B.n239 B.n236 10.6151
R1389 B.n240 B.n239 10.6151
R1390 B.n243 B.n240 10.6151
R1391 B.n244 B.n243 10.6151
R1392 B.n247 B.n244 10.6151
R1393 B.n248 B.n247 10.6151
R1394 B.n252 B.n251 10.6151
R1395 B.n255 B.n252 10.6151
R1396 B.n256 B.n255 10.6151
R1397 B.n259 B.n256 10.6151
R1398 B.n260 B.n259 10.6151
R1399 B.n263 B.n260 10.6151
R1400 B.n264 B.n263 10.6151
R1401 B.n267 B.n264 10.6151
R1402 B.n272 B.n269 10.6151
R1403 B.n273 B.n272 10.6151
R1404 B.n276 B.n273 10.6151
R1405 B.n277 B.n276 10.6151
R1406 B.n280 B.n277 10.6151
R1407 B.n281 B.n280 10.6151
R1408 B.n284 B.n281 10.6151
R1409 B.n285 B.n284 10.6151
R1410 B.n288 B.n285 10.6151
R1411 B.n289 B.n288 10.6151
R1412 B.n292 B.n289 10.6151
R1413 B.n293 B.n292 10.6151
R1414 B.n296 B.n293 10.6151
R1415 B.n297 B.n296 10.6151
R1416 B.n300 B.n297 10.6151
R1417 B.n301 B.n300 10.6151
R1418 B.n304 B.n301 10.6151
R1419 B.n305 B.n304 10.6151
R1420 B.n308 B.n305 10.6151
R1421 B.n309 B.n308 10.6151
R1422 B.n312 B.n309 10.6151
R1423 B.n313 B.n312 10.6151
R1424 B.n316 B.n313 10.6151
R1425 B.n317 B.n316 10.6151
R1426 B.n320 B.n317 10.6151
R1427 B.n321 B.n320 10.6151
R1428 B.n324 B.n321 10.6151
R1429 B.n325 B.n324 10.6151
R1430 B.n328 B.n325 10.6151
R1431 B.n329 B.n328 10.6151
R1432 B.n332 B.n329 10.6151
R1433 B.n333 B.n332 10.6151
R1434 B.n336 B.n333 10.6151
R1435 B.n337 B.n336 10.6151
R1436 B.n340 B.n337 10.6151
R1437 B.n341 B.n340 10.6151
R1438 B.n344 B.n341 10.6151
R1439 B.n345 B.n344 10.6151
R1440 B.n348 B.n345 10.6151
R1441 B.n349 B.n348 10.6151
R1442 B.n352 B.n349 10.6151
R1443 B.n353 B.n352 10.6151
R1444 B.n356 B.n353 10.6151
R1445 B.n357 B.n356 10.6151
R1446 B.n360 B.n357 10.6151
R1447 B.n361 B.n360 10.6151
R1448 B.n364 B.n361 10.6151
R1449 B.n365 B.n364 10.6151
R1450 B.n368 B.n365 10.6151
R1451 B.n369 B.n368 10.6151
R1452 B.n372 B.n369 10.6151
R1453 B.n373 B.n372 10.6151
R1454 B.n939 B.n373 10.6151
R1455 B.n761 B.n453 10.6151
R1456 B.n762 B.n761 10.6151
R1457 B.n763 B.n762 10.6151
R1458 B.n763 B.n445 10.6151
R1459 B.n773 B.n445 10.6151
R1460 B.n774 B.n773 10.6151
R1461 B.n775 B.n774 10.6151
R1462 B.n775 B.n437 10.6151
R1463 B.n785 B.n437 10.6151
R1464 B.n786 B.n785 10.6151
R1465 B.n787 B.n786 10.6151
R1466 B.n787 B.n429 10.6151
R1467 B.n797 B.n429 10.6151
R1468 B.n798 B.n797 10.6151
R1469 B.n799 B.n798 10.6151
R1470 B.n799 B.n421 10.6151
R1471 B.n809 B.n421 10.6151
R1472 B.n810 B.n809 10.6151
R1473 B.n811 B.n810 10.6151
R1474 B.n811 B.n413 10.6151
R1475 B.n821 B.n413 10.6151
R1476 B.n822 B.n821 10.6151
R1477 B.n823 B.n822 10.6151
R1478 B.n823 B.n405 10.6151
R1479 B.n833 B.n405 10.6151
R1480 B.n834 B.n833 10.6151
R1481 B.n835 B.n834 10.6151
R1482 B.n835 B.n398 10.6151
R1483 B.n846 B.n398 10.6151
R1484 B.n847 B.n846 10.6151
R1485 B.n848 B.n847 10.6151
R1486 B.n848 B.n390 10.6151
R1487 B.n858 B.n390 10.6151
R1488 B.n859 B.n858 10.6151
R1489 B.n860 B.n859 10.6151
R1490 B.n860 B.n382 10.6151
R1491 B.n870 B.n382 10.6151
R1492 B.n871 B.n870 10.6151
R1493 B.n873 B.n871 10.6151
R1494 B.n873 B.n872 10.6151
R1495 B.n872 B.n374 10.6151
R1496 B.n884 B.n374 10.6151
R1497 B.n885 B.n884 10.6151
R1498 B.n886 B.n885 10.6151
R1499 B.n887 B.n886 10.6151
R1500 B.n889 B.n887 10.6151
R1501 B.n890 B.n889 10.6151
R1502 B.n891 B.n890 10.6151
R1503 B.n892 B.n891 10.6151
R1504 B.n894 B.n892 10.6151
R1505 B.n895 B.n894 10.6151
R1506 B.n896 B.n895 10.6151
R1507 B.n897 B.n896 10.6151
R1508 B.n899 B.n897 10.6151
R1509 B.n900 B.n899 10.6151
R1510 B.n901 B.n900 10.6151
R1511 B.n902 B.n901 10.6151
R1512 B.n904 B.n902 10.6151
R1513 B.n905 B.n904 10.6151
R1514 B.n906 B.n905 10.6151
R1515 B.n907 B.n906 10.6151
R1516 B.n909 B.n907 10.6151
R1517 B.n910 B.n909 10.6151
R1518 B.n911 B.n910 10.6151
R1519 B.n912 B.n911 10.6151
R1520 B.n914 B.n912 10.6151
R1521 B.n915 B.n914 10.6151
R1522 B.n916 B.n915 10.6151
R1523 B.n917 B.n916 10.6151
R1524 B.n919 B.n917 10.6151
R1525 B.n920 B.n919 10.6151
R1526 B.n921 B.n920 10.6151
R1527 B.n922 B.n921 10.6151
R1528 B.n924 B.n922 10.6151
R1529 B.n925 B.n924 10.6151
R1530 B.n926 B.n925 10.6151
R1531 B.n927 B.n926 10.6151
R1532 B.n929 B.n927 10.6151
R1533 B.n930 B.n929 10.6151
R1534 B.n931 B.n930 10.6151
R1535 B.n932 B.n931 10.6151
R1536 B.n934 B.n932 10.6151
R1537 B.n935 B.n934 10.6151
R1538 B.n936 B.n935 10.6151
R1539 B.n937 B.n936 10.6151
R1540 B.n938 B.n937 10.6151
R1541 B.n755 B.n457 10.6151
R1542 B.n750 B.n457 10.6151
R1543 B.n750 B.n749 10.6151
R1544 B.n749 B.n748 10.6151
R1545 B.n748 B.n745 10.6151
R1546 B.n745 B.n744 10.6151
R1547 B.n744 B.n741 10.6151
R1548 B.n741 B.n740 10.6151
R1549 B.n740 B.n737 10.6151
R1550 B.n737 B.n736 10.6151
R1551 B.n736 B.n733 10.6151
R1552 B.n733 B.n732 10.6151
R1553 B.n732 B.n729 10.6151
R1554 B.n729 B.n728 10.6151
R1555 B.n728 B.n725 10.6151
R1556 B.n725 B.n724 10.6151
R1557 B.n724 B.n721 10.6151
R1558 B.n721 B.n720 10.6151
R1559 B.n720 B.n717 10.6151
R1560 B.n717 B.n716 10.6151
R1561 B.n716 B.n713 10.6151
R1562 B.n713 B.n712 10.6151
R1563 B.n712 B.n709 10.6151
R1564 B.n709 B.n708 10.6151
R1565 B.n708 B.n705 10.6151
R1566 B.n705 B.n704 10.6151
R1567 B.n704 B.n701 10.6151
R1568 B.n701 B.n700 10.6151
R1569 B.n700 B.n697 10.6151
R1570 B.n697 B.n696 10.6151
R1571 B.n696 B.n693 10.6151
R1572 B.n693 B.n692 10.6151
R1573 B.n692 B.n689 10.6151
R1574 B.n689 B.n688 10.6151
R1575 B.n688 B.n685 10.6151
R1576 B.n685 B.n684 10.6151
R1577 B.n684 B.n681 10.6151
R1578 B.n681 B.n680 10.6151
R1579 B.n680 B.n677 10.6151
R1580 B.n677 B.n676 10.6151
R1581 B.n676 B.n673 10.6151
R1582 B.n673 B.n672 10.6151
R1583 B.n672 B.n669 10.6151
R1584 B.n669 B.n668 10.6151
R1585 B.n668 B.n665 10.6151
R1586 B.n665 B.n664 10.6151
R1587 B.n664 B.n661 10.6151
R1588 B.n661 B.n660 10.6151
R1589 B.n660 B.n657 10.6151
R1590 B.n657 B.n656 10.6151
R1591 B.n656 B.n653 10.6151
R1592 B.n653 B.n652 10.6151
R1593 B.n652 B.n649 10.6151
R1594 B.n647 B.n644 10.6151
R1595 B.n644 B.n643 10.6151
R1596 B.n643 B.n640 10.6151
R1597 B.n640 B.n639 10.6151
R1598 B.n639 B.n636 10.6151
R1599 B.n636 B.n635 10.6151
R1600 B.n635 B.n632 10.6151
R1601 B.n632 B.n631 10.6151
R1602 B.n628 B.n627 10.6151
R1603 B.n627 B.n624 10.6151
R1604 B.n624 B.n623 10.6151
R1605 B.n623 B.n620 10.6151
R1606 B.n620 B.n619 10.6151
R1607 B.n619 B.n616 10.6151
R1608 B.n616 B.n615 10.6151
R1609 B.n615 B.n612 10.6151
R1610 B.n612 B.n611 10.6151
R1611 B.n611 B.n608 10.6151
R1612 B.n608 B.n607 10.6151
R1613 B.n607 B.n604 10.6151
R1614 B.n604 B.n603 10.6151
R1615 B.n603 B.n600 10.6151
R1616 B.n600 B.n599 10.6151
R1617 B.n599 B.n596 10.6151
R1618 B.n596 B.n595 10.6151
R1619 B.n595 B.n592 10.6151
R1620 B.n592 B.n591 10.6151
R1621 B.n591 B.n588 10.6151
R1622 B.n588 B.n587 10.6151
R1623 B.n587 B.n584 10.6151
R1624 B.n584 B.n583 10.6151
R1625 B.n583 B.n580 10.6151
R1626 B.n580 B.n579 10.6151
R1627 B.n579 B.n576 10.6151
R1628 B.n576 B.n575 10.6151
R1629 B.n575 B.n572 10.6151
R1630 B.n572 B.n571 10.6151
R1631 B.n571 B.n568 10.6151
R1632 B.n568 B.n567 10.6151
R1633 B.n567 B.n564 10.6151
R1634 B.n564 B.n563 10.6151
R1635 B.n563 B.n560 10.6151
R1636 B.n560 B.n559 10.6151
R1637 B.n559 B.n556 10.6151
R1638 B.n556 B.n555 10.6151
R1639 B.n555 B.n552 10.6151
R1640 B.n552 B.n551 10.6151
R1641 B.n551 B.n548 10.6151
R1642 B.n548 B.n547 10.6151
R1643 B.n547 B.n544 10.6151
R1644 B.n544 B.n543 10.6151
R1645 B.n543 B.n540 10.6151
R1646 B.n540 B.n539 10.6151
R1647 B.n539 B.n536 10.6151
R1648 B.n536 B.n535 10.6151
R1649 B.n535 B.n532 10.6151
R1650 B.n532 B.n531 10.6151
R1651 B.n531 B.n528 10.6151
R1652 B.n528 B.n527 10.6151
R1653 B.n527 B.n524 10.6151
R1654 B.n524 B.n523 10.6151
R1655 B.n757 B.n756 10.6151
R1656 B.n757 B.n449 10.6151
R1657 B.n767 B.n449 10.6151
R1658 B.n768 B.n767 10.6151
R1659 B.n769 B.n768 10.6151
R1660 B.n769 B.n441 10.6151
R1661 B.n779 B.n441 10.6151
R1662 B.n780 B.n779 10.6151
R1663 B.n781 B.n780 10.6151
R1664 B.n781 B.n433 10.6151
R1665 B.n791 B.n433 10.6151
R1666 B.n792 B.n791 10.6151
R1667 B.n793 B.n792 10.6151
R1668 B.n793 B.n425 10.6151
R1669 B.n803 B.n425 10.6151
R1670 B.n804 B.n803 10.6151
R1671 B.n805 B.n804 10.6151
R1672 B.n805 B.n417 10.6151
R1673 B.n815 B.n417 10.6151
R1674 B.n816 B.n815 10.6151
R1675 B.n817 B.n816 10.6151
R1676 B.n817 B.n409 10.6151
R1677 B.n827 B.n409 10.6151
R1678 B.n828 B.n827 10.6151
R1679 B.n829 B.n828 10.6151
R1680 B.n829 B.n401 10.6151
R1681 B.n840 B.n401 10.6151
R1682 B.n841 B.n840 10.6151
R1683 B.n842 B.n841 10.6151
R1684 B.n842 B.n394 10.6151
R1685 B.n852 B.n394 10.6151
R1686 B.n853 B.n852 10.6151
R1687 B.n854 B.n853 10.6151
R1688 B.n854 B.n386 10.6151
R1689 B.n864 B.n386 10.6151
R1690 B.n865 B.n864 10.6151
R1691 B.n866 B.n865 10.6151
R1692 B.n866 B.n378 10.6151
R1693 B.n877 B.n378 10.6151
R1694 B.n878 B.n877 10.6151
R1695 B.n879 B.n878 10.6151
R1696 B.n879 B.n0 10.6151
R1697 B.n1026 B.n1 10.6151
R1698 B.n1026 B.n1025 10.6151
R1699 B.n1025 B.n1024 10.6151
R1700 B.n1024 B.n10 10.6151
R1701 B.n1018 B.n10 10.6151
R1702 B.n1018 B.n1017 10.6151
R1703 B.n1017 B.n1016 10.6151
R1704 B.n1016 B.n17 10.6151
R1705 B.n1010 B.n17 10.6151
R1706 B.n1010 B.n1009 10.6151
R1707 B.n1009 B.n1008 10.6151
R1708 B.n1008 B.n24 10.6151
R1709 B.n1002 B.n24 10.6151
R1710 B.n1002 B.n1001 10.6151
R1711 B.n1001 B.n1000 10.6151
R1712 B.n1000 B.n30 10.6151
R1713 B.n994 B.n30 10.6151
R1714 B.n994 B.n993 10.6151
R1715 B.n993 B.n992 10.6151
R1716 B.n992 B.n38 10.6151
R1717 B.n986 B.n38 10.6151
R1718 B.n986 B.n985 10.6151
R1719 B.n985 B.n984 10.6151
R1720 B.n984 B.n45 10.6151
R1721 B.n978 B.n45 10.6151
R1722 B.n978 B.n977 10.6151
R1723 B.n977 B.n976 10.6151
R1724 B.n976 B.n52 10.6151
R1725 B.n970 B.n52 10.6151
R1726 B.n970 B.n969 10.6151
R1727 B.n969 B.n968 10.6151
R1728 B.n968 B.n59 10.6151
R1729 B.n962 B.n59 10.6151
R1730 B.n962 B.n961 10.6151
R1731 B.n961 B.n960 10.6151
R1732 B.n960 B.n66 10.6151
R1733 B.n954 B.n66 10.6151
R1734 B.n954 B.n953 10.6151
R1735 B.n953 B.n952 10.6151
R1736 B.n952 B.n73 10.6151
R1737 B.n946 B.n73 10.6151
R1738 B.n946 B.n945 10.6151
R1739 B.n837 B.t4 8.72455
R1740 B.n32 B.t0 8.72455
R1741 B.n251 B.n145 6.5566
R1742 B.n268 B.n267 6.5566
R1743 B.n648 B.n647 6.5566
R1744 B.n631 B.n521 6.5566
R1745 B.n248 B.n145 4.05904
R1746 B.n269 B.n268 4.05904
R1747 B.n649 B.n648 4.05904
R1748 B.n628 B.n521 4.05904
R1749 B.n1032 B.n0 2.81026
R1750 B.n1032 B.n1 2.81026
R1751 B.n868 B.t1 0.513679
R1752 B.t2 B.n1020 0.513679
R1753 VN.n4 VN.t0 181
R1754 VN.n20 VN.t3 181
R1755 VN.n29 VN.n16 161.3
R1756 VN.n28 VN.n27 161.3
R1757 VN.n26 VN.n17 161.3
R1758 VN.n25 VN.n24 161.3
R1759 VN.n23 VN.n18 161.3
R1760 VN.n22 VN.n21 161.3
R1761 VN.n13 VN.n0 161.3
R1762 VN.n12 VN.n11 161.3
R1763 VN.n10 VN.n1 161.3
R1764 VN.n9 VN.n8 161.3
R1765 VN.n7 VN.n2 161.3
R1766 VN.n6 VN.n5 161.3
R1767 VN.n3 VN.t5 146.965
R1768 VN.n14 VN.t2 146.965
R1769 VN.n19 VN.t1 146.965
R1770 VN.n30 VN.t4 146.965
R1771 VN.n15 VN.n14 99.596
R1772 VN.n31 VN.n30 99.596
R1773 VN.n4 VN.n3 60.4656
R1774 VN.n20 VN.n19 60.4656
R1775 VN.n8 VN.n1 56.5617
R1776 VN.n24 VN.n17 56.5617
R1777 VN VN.n31 52.3542
R1778 VN.n7 VN.n6 24.5923
R1779 VN.n8 VN.n7 24.5923
R1780 VN.n12 VN.n1 24.5923
R1781 VN.n13 VN.n12 24.5923
R1782 VN.n24 VN.n23 24.5923
R1783 VN.n23 VN.n22 24.5923
R1784 VN.n29 VN.n28 24.5923
R1785 VN.n28 VN.n17 24.5923
R1786 VN.n6 VN.n3 12.2964
R1787 VN.n22 VN.n19 12.2964
R1788 VN.n14 VN.n13 11.3127
R1789 VN.n30 VN.n29 11.3127
R1790 VN.n21 VN.n20 6.75133
R1791 VN.n5 VN.n4 6.75133
R1792 VN.n31 VN.n16 0.278335
R1793 VN.n15 VN.n0 0.278335
R1794 VN.n27 VN.n16 0.189894
R1795 VN.n27 VN.n26 0.189894
R1796 VN.n26 VN.n25 0.189894
R1797 VN.n25 VN.n18 0.189894
R1798 VN.n21 VN.n18 0.189894
R1799 VN.n5 VN.n2 0.189894
R1800 VN.n9 VN.n2 0.189894
R1801 VN.n10 VN.n9 0.189894
R1802 VN.n11 VN.n10 0.189894
R1803 VN.n11 VN.n0 0.189894
R1804 VN VN.n15 0.153485
R1805 VTAIL.n362 VTAIL.n278 289.615
R1806 VTAIL.n86 VTAIL.n2 289.615
R1807 VTAIL.n272 VTAIL.n188 289.615
R1808 VTAIL.n180 VTAIL.n96 289.615
R1809 VTAIL.n306 VTAIL.n305 185
R1810 VTAIL.n311 VTAIL.n310 185
R1811 VTAIL.n313 VTAIL.n312 185
R1812 VTAIL.n302 VTAIL.n301 185
R1813 VTAIL.n319 VTAIL.n318 185
R1814 VTAIL.n321 VTAIL.n320 185
R1815 VTAIL.n298 VTAIL.n297 185
R1816 VTAIL.n327 VTAIL.n326 185
R1817 VTAIL.n329 VTAIL.n328 185
R1818 VTAIL.n294 VTAIL.n293 185
R1819 VTAIL.n335 VTAIL.n334 185
R1820 VTAIL.n337 VTAIL.n336 185
R1821 VTAIL.n290 VTAIL.n289 185
R1822 VTAIL.n343 VTAIL.n342 185
R1823 VTAIL.n345 VTAIL.n344 185
R1824 VTAIL.n286 VTAIL.n285 185
R1825 VTAIL.n352 VTAIL.n351 185
R1826 VTAIL.n353 VTAIL.n284 185
R1827 VTAIL.n355 VTAIL.n354 185
R1828 VTAIL.n282 VTAIL.n281 185
R1829 VTAIL.n361 VTAIL.n360 185
R1830 VTAIL.n363 VTAIL.n362 185
R1831 VTAIL.n30 VTAIL.n29 185
R1832 VTAIL.n35 VTAIL.n34 185
R1833 VTAIL.n37 VTAIL.n36 185
R1834 VTAIL.n26 VTAIL.n25 185
R1835 VTAIL.n43 VTAIL.n42 185
R1836 VTAIL.n45 VTAIL.n44 185
R1837 VTAIL.n22 VTAIL.n21 185
R1838 VTAIL.n51 VTAIL.n50 185
R1839 VTAIL.n53 VTAIL.n52 185
R1840 VTAIL.n18 VTAIL.n17 185
R1841 VTAIL.n59 VTAIL.n58 185
R1842 VTAIL.n61 VTAIL.n60 185
R1843 VTAIL.n14 VTAIL.n13 185
R1844 VTAIL.n67 VTAIL.n66 185
R1845 VTAIL.n69 VTAIL.n68 185
R1846 VTAIL.n10 VTAIL.n9 185
R1847 VTAIL.n76 VTAIL.n75 185
R1848 VTAIL.n77 VTAIL.n8 185
R1849 VTAIL.n79 VTAIL.n78 185
R1850 VTAIL.n6 VTAIL.n5 185
R1851 VTAIL.n85 VTAIL.n84 185
R1852 VTAIL.n87 VTAIL.n86 185
R1853 VTAIL.n273 VTAIL.n272 185
R1854 VTAIL.n271 VTAIL.n270 185
R1855 VTAIL.n192 VTAIL.n191 185
R1856 VTAIL.n265 VTAIL.n264 185
R1857 VTAIL.n263 VTAIL.n194 185
R1858 VTAIL.n262 VTAIL.n261 185
R1859 VTAIL.n197 VTAIL.n195 185
R1860 VTAIL.n256 VTAIL.n255 185
R1861 VTAIL.n254 VTAIL.n253 185
R1862 VTAIL.n201 VTAIL.n200 185
R1863 VTAIL.n248 VTAIL.n247 185
R1864 VTAIL.n246 VTAIL.n245 185
R1865 VTAIL.n205 VTAIL.n204 185
R1866 VTAIL.n240 VTAIL.n239 185
R1867 VTAIL.n238 VTAIL.n237 185
R1868 VTAIL.n209 VTAIL.n208 185
R1869 VTAIL.n232 VTAIL.n231 185
R1870 VTAIL.n230 VTAIL.n229 185
R1871 VTAIL.n213 VTAIL.n212 185
R1872 VTAIL.n224 VTAIL.n223 185
R1873 VTAIL.n222 VTAIL.n221 185
R1874 VTAIL.n217 VTAIL.n216 185
R1875 VTAIL.n181 VTAIL.n180 185
R1876 VTAIL.n179 VTAIL.n178 185
R1877 VTAIL.n100 VTAIL.n99 185
R1878 VTAIL.n173 VTAIL.n172 185
R1879 VTAIL.n171 VTAIL.n102 185
R1880 VTAIL.n170 VTAIL.n169 185
R1881 VTAIL.n105 VTAIL.n103 185
R1882 VTAIL.n164 VTAIL.n163 185
R1883 VTAIL.n162 VTAIL.n161 185
R1884 VTAIL.n109 VTAIL.n108 185
R1885 VTAIL.n156 VTAIL.n155 185
R1886 VTAIL.n154 VTAIL.n153 185
R1887 VTAIL.n113 VTAIL.n112 185
R1888 VTAIL.n148 VTAIL.n147 185
R1889 VTAIL.n146 VTAIL.n145 185
R1890 VTAIL.n117 VTAIL.n116 185
R1891 VTAIL.n140 VTAIL.n139 185
R1892 VTAIL.n138 VTAIL.n137 185
R1893 VTAIL.n121 VTAIL.n120 185
R1894 VTAIL.n132 VTAIL.n131 185
R1895 VTAIL.n130 VTAIL.n129 185
R1896 VTAIL.n125 VTAIL.n124 185
R1897 VTAIL.n307 VTAIL.t11 147.659
R1898 VTAIL.n31 VTAIL.t1 147.659
R1899 VTAIL.n218 VTAIL.t4 147.659
R1900 VTAIL.n126 VTAIL.t8 147.659
R1901 VTAIL.n311 VTAIL.n305 104.615
R1902 VTAIL.n312 VTAIL.n311 104.615
R1903 VTAIL.n312 VTAIL.n301 104.615
R1904 VTAIL.n319 VTAIL.n301 104.615
R1905 VTAIL.n320 VTAIL.n319 104.615
R1906 VTAIL.n320 VTAIL.n297 104.615
R1907 VTAIL.n327 VTAIL.n297 104.615
R1908 VTAIL.n328 VTAIL.n327 104.615
R1909 VTAIL.n328 VTAIL.n293 104.615
R1910 VTAIL.n335 VTAIL.n293 104.615
R1911 VTAIL.n336 VTAIL.n335 104.615
R1912 VTAIL.n336 VTAIL.n289 104.615
R1913 VTAIL.n343 VTAIL.n289 104.615
R1914 VTAIL.n344 VTAIL.n343 104.615
R1915 VTAIL.n344 VTAIL.n285 104.615
R1916 VTAIL.n352 VTAIL.n285 104.615
R1917 VTAIL.n353 VTAIL.n352 104.615
R1918 VTAIL.n354 VTAIL.n353 104.615
R1919 VTAIL.n354 VTAIL.n281 104.615
R1920 VTAIL.n361 VTAIL.n281 104.615
R1921 VTAIL.n362 VTAIL.n361 104.615
R1922 VTAIL.n35 VTAIL.n29 104.615
R1923 VTAIL.n36 VTAIL.n35 104.615
R1924 VTAIL.n36 VTAIL.n25 104.615
R1925 VTAIL.n43 VTAIL.n25 104.615
R1926 VTAIL.n44 VTAIL.n43 104.615
R1927 VTAIL.n44 VTAIL.n21 104.615
R1928 VTAIL.n51 VTAIL.n21 104.615
R1929 VTAIL.n52 VTAIL.n51 104.615
R1930 VTAIL.n52 VTAIL.n17 104.615
R1931 VTAIL.n59 VTAIL.n17 104.615
R1932 VTAIL.n60 VTAIL.n59 104.615
R1933 VTAIL.n60 VTAIL.n13 104.615
R1934 VTAIL.n67 VTAIL.n13 104.615
R1935 VTAIL.n68 VTAIL.n67 104.615
R1936 VTAIL.n68 VTAIL.n9 104.615
R1937 VTAIL.n76 VTAIL.n9 104.615
R1938 VTAIL.n77 VTAIL.n76 104.615
R1939 VTAIL.n78 VTAIL.n77 104.615
R1940 VTAIL.n78 VTAIL.n5 104.615
R1941 VTAIL.n85 VTAIL.n5 104.615
R1942 VTAIL.n86 VTAIL.n85 104.615
R1943 VTAIL.n272 VTAIL.n271 104.615
R1944 VTAIL.n271 VTAIL.n191 104.615
R1945 VTAIL.n264 VTAIL.n191 104.615
R1946 VTAIL.n264 VTAIL.n263 104.615
R1947 VTAIL.n263 VTAIL.n262 104.615
R1948 VTAIL.n262 VTAIL.n195 104.615
R1949 VTAIL.n255 VTAIL.n195 104.615
R1950 VTAIL.n255 VTAIL.n254 104.615
R1951 VTAIL.n254 VTAIL.n200 104.615
R1952 VTAIL.n247 VTAIL.n200 104.615
R1953 VTAIL.n247 VTAIL.n246 104.615
R1954 VTAIL.n246 VTAIL.n204 104.615
R1955 VTAIL.n239 VTAIL.n204 104.615
R1956 VTAIL.n239 VTAIL.n238 104.615
R1957 VTAIL.n238 VTAIL.n208 104.615
R1958 VTAIL.n231 VTAIL.n208 104.615
R1959 VTAIL.n231 VTAIL.n230 104.615
R1960 VTAIL.n230 VTAIL.n212 104.615
R1961 VTAIL.n223 VTAIL.n212 104.615
R1962 VTAIL.n223 VTAIL.n222 104.615
R1963 VTAIL.n222 VTAIL.n216 104.615
R1964 VTAIL.n180 VTAIL.n179 104.615
R1965 VTAIL.n179 VTAIL.n99 104.615
R1966 VTAIL.n172 VTAIL.n99 104.615
R1967 VTAIL.n172 VTAIL.n171 104.615
R1968 VTAIL.n171 VTAIL.n170 104.615
R1969 VTAIL.n170 VTAIL.n103 104.615
R1970 VTAIL.n163 VTAIL.n103 104.615
R1971 VTAIL.n163 VTAIL.n162 104.615
R1972 VTAIL.n162 VTAIL.n108 104.615
R1973 VTAIL.n155 VTAIL.n108 104.615
R1974 VTAIL.n155 VTAIL.n154 104.615
R1975 VTAIL.n154 VTAIL.n112 104.615
R1976 VTAIL.n147 VTAIL.n112 104.615
R1977 VTAIL.n147 VTAIL.n146 104.615
R1978 VTAIL.n146 VTAIL.n116 104.615
R1979 VTAIL.n139 VTAIL.n116 104.615
R1980 VTAIL.n139 VTAIL.n138 104.615
R1981 VTAIL.n138 VTAIL.n120 104.615
R1982 VTAIL.n131 VTAIL.n120 104.615
R1983 VTAIL.n131 VTAIL.n130 104.615
R1984 VTAIL.n130 VTAIL.n124 104.615
R1985 VTAIL.t11 VTAIL.n305 52.3082
R1986 VTAIL.t1 VTAIL.n29 52.3082
R1987 VTAIL.t4 VTAIL.n216 52.3082
R1988 VTAIL.t8 VTAIL.n124 52.3082
R1989 VTAIL.n187 VTAIL.n186 45.6505
R1990 VTAIL.n95 VTAIL.n94 45.6505
R1991 VTAIL.n1 VTAIL.n0 45.6503
R1992 VTAIL.n93 VTAIL.n92 45.6503
R1993 VTAIL.n367 VTAIL.n366 33.7369
R1994 VTAIL.n91 VTAIL.n90 33.7369
R1995 VTAIL.n277 VTAIL.n276 33.7369
R1996 VTAIL.n185 VTAIL.n184 33.7369
R1997 VTAIL.n95 VTAIL.n93 31.4358
R1998 VTAIL.n367 VTAIL.n277 28.8669
R1999 VTAIL.n307 VTAIL.n306 15.6677
R2000 VTAIL.n31 VTAIL.n30 15.6677
R2001 VTAIL.n218 VTAIL.n217 15.6677
R2002 VTAIL.n126 VTAIL.n125 15.6677
R2003 VTAIL.n355 VTAIL.n284 13.1884
R2004 VTAIL.n79 VTAIL.n8 13.1884
R2005 VTAIL.n265 VTAIL.n194 13.1884
R2006 VTAIL.n173 VTAIL.n102 13.1884
R2007 VTAIL.n310 VTAIL.n309 12.8005
R2008 VTAIL.n351 VTAIL.n350 12.8005
R2009 VTAIL.n356 VTAIL.n282 12.8005
R2010 VTAIL.n34 VTAIL.n33 12.8005
R2011 VTAIL.n75 VTAIL.n74 12.8005
R2012 VTAIL.n80 VTAIL.n6 12.8005
R2013 VTAIL.n266 VTAIL.n192 12.8005
R2014 VTAIL.n261 VTAIL.n196 12.8005
R2015 VTAIL.n221 VTAIL.n220 12.8005
R2016 VTAIL.n174 VTAIL.n100 12.8005
R2017 VTAIL.n169 VTAIL.n104 12.8005
R2018 VTAIL.n129 VTAIL.n128 12.8005
R2019 VTAIL.n313 VTAIL.n304 12.0247
R2020 VTAIL.n349 VTAIL.n286 12.0247
R2021 VTAIL.n360 VTAIL.n359 12.0247
R2022 VTAIL.n37 VTAIL.n28 12.0247
R2023 VTAIL.n73 VTAIL.n10 12.0247
R2024 VTAIL.n84 VTAIL.n83 12.0247
R2025 VTAIL.n270 VTAIL.n269 12.0247
R2026 VTAIL.n260 VTAIL.n197 12.0247
R2027 VTAIL.n224 VTAIL.n215 12.0247
R2028 VTAIL.n178 VTAIL.n177 12.0247
R2029 VTAIL.n168 VTAIL.n105 12.0247
R2030 VTAIL.n132 VTAIL.n123 12.0247
R2031 VTAIL.n314 VTAIL.n302 11.249
R2032 VTAIL.n346 VTAIL.n345 11.249
R2033 VTAIL.n363 VTAIL.n280 11.249
R2034 VTAIL.n38 VTAIL.n26 11.249
R2035 VTAIL.n70 VTAIL.n69 11.249
R2036 VTAIL.n87 VTAIL.n4 11.249
R2037 VTAIL.n273 VTAIL.n190 11.249
R2038 VTAIL.n257 VTAIL.n256 11.249
R2039 VTAIL.n225 VTAIL.n213 11.249
R2040 VTAIL.n181 VTAIL.n98 11.249
R2041 VTAIL.n165 VTAIL.n164 11.249
R2042 VTAIL.n133 VTAIL.n121 11.249
R2043 VTAIL.n318 VTAIL.n317 10.4732
R2044 VTAIL.n342 VTAIL.n288 10.4732
R2045 VTAIL.n364 VTAIL.n278 10.4732
R2046 VTAIL.n42 VTAIL.n41 10.4732
R2047 VTAIL.n66 VTAIL.n12 10.4732
R2048 VTAIL.n88 VTAIL.n2 10.4732
R2049 VTAIL.n274 VTAIL.n188 10.4732
R2050 VTAIL.n253 VTAIL.n199 10.4732
R2051 VTAIL.n229 VTAIL.n228 10.4732
R2052 VTAIL.n182 VTAIL.n96 10.4732
R2053 VTAIL.n161 VTAIL.n107 10.4732
R2054 VTAIL.n137 VTAIL.n136 10.4732
R2055 VTAIL.n321 VTAIL.n300 9.69747
R2056 VTAIL.n341 VTAIL.n290 9.69747
R2057 VTAIL.n45 VTAIL.n24 9.69747
R2058 VTAIL.n65 VTAIL.n14 9.69747
R2059 VTAIL.n252 VTAIL.n201 9.69747
R2060 VTAIL.n232 VTAIL.n211 9.69747
R2061 VTAIL.n160 VTAIL.n109 9.69747
R2062 VTAIL.n140 VTAIL.n119 9.69747
R2063 VTAIL.n366 VTAIL.n365 9.45567
R2064 VTAIL.n90 VTAIL.n89 9.45567
R2065 VTAIL.n276 VTAIL.n275 9.45567
R2066 VTAIL.n184 VTAIL.n183 9.45567
R2067 VTAIL.n365 VTAIL.n364 9.3005
R2068 VTAIL.n280 VTAIL.n279 9.3005
R2069 VTAIL.n359 VTAIL.n358 9.3005
R2070 VTAIL.n357 VTAIL.n356 9.3005
R2071 VTAIL.n296 VTAIL.n295 9.3005
R2072 VTAIL.n325 VTAIL.n324 9.3005
R2073 VTAIL.n323 VTAIL.n322 9.3005
R2074 VTAIL.n300 VTAIL.n299 9.3005
R2075 VTAIL.n317 VTAIL.n316 9.3005
R2076 VTAIL.n315 VTAIL.n314 9.3005
R2077 VTAIL.n304 VTAIL.n303 9.3005
R2078 VTAIL.n309 VTAIL.n308 9.3005
R2079 VTAIL.n331 VTAIL.n330 9.3005
R2080 VTAIL.n333 VTAIL.n332 9.3005
R2081 VTAIL.n292 VTAIL.n291 9.3005
R2082 VTAIL.n339 VTAIL.n338 9.3005
R2083 VTAIL.n341 VTAIL.n340 9.3005
R2084 VTAIL.n288 VTAIL.n287 9.3005
R2085 VTAIL.n347 VTAIL.n346 9.3005
R2086 VTAIL.n349 VTAIL.n348 9.3005
R2087 VTAIL.n350 VTAIL.n283 9.3005
R2088 VTAIL.n89 VTAIL.n88 9.3005
R2089 VTAIL.n4 VTAIL.n3 9.3005
R2090 VTAIL.n83 VTAIL.n82 9.3005
R2091 VTAIL.n81 VTAIL.n80 9.3005
R2092 VTAIL.n20 VTAIL.n19 9.3005
R2093 VTAIL.n49 VTAIL.n48 9.3005
R2094 VTAIL.n47 VTAIL.n46 9.3005
R2095 VTAIL.n24 VTAIL.n23 9.3005
R2096 VTAIL.n41 VTAIL.n40 9.3005
R2097 VTAIL.n39 VTAIL.n38 9.3005
R2098 VTAIL.n28 VTAIL.n27 9.3005
R2099 VTAIL.n33 VTAIL.n32 9.3005
R2100 VTAIL.n55 VTAIL.n54 9.3005
R2101 VTAIL.n57 VTAIL.n56 9.3005
R2102 VTAIL.n16 VTAIL.n15 9.3005
R2103 VTAIL.n63 VTAIL.n62 9.3005
R2104 VTAIL.n65 VTAIL.n64 9.3005
R2105 VTAIL.n12 VTAIL.n11 9.3005
R2106 VTAIL.n71 VTAIL.n70 9.3005
R2107 VTAIL.n73 VTAIL.n72 9.3005
R2108 VTAIL.n74 VTAIL.n7 9.3005
R2109 VTAIL.n244 VTAIL.n243 9.3005
R2110 VTAIL.n203 VTAIL.n202 9.3005
R2111 VTAIL.n250 VTAIL.n249 9.3005
R2112 VTAIL.n252 VTAIL.n251 9.3005
R2113 VTAIL.n199 VTAIL.n198 9.3005
R2114 VTAIL.n258 VTAIL.n257 9.3005
R2115 VTAIL.n260 VTAIL.n259 9.3005
R2116 VTAIL.n196 VTAIL.n193 9.3005
R2117 VTAIL.n275 VTAIL.n274 9.3005
R2118 VTAIL.n190 VTAIL.n189 9.3005
R2119 VTAIL.n269 VTAIL.n268 9.3005
R2120 VTAIL.n267 VTAIL.n266 9.3005
R2121 VTAIL.n242 VTAIL.n241 9.3005
R2122 VTAIL.n207 VTAIL.n206 9.3005
R2123 VTAIL.n236 VTAIL.n235 9.3005
R2124 VTAIL.n234 VTAIL.n233 9.3005
R2125 VTAIL.n211 VTAIL.n210 9.3005
R2126 VTAIL.n228 VTAIL.n227 9.3005
R2127 VTAIL.n226 VTAIL.n225 9.3005
R2128 VTAIL.n215 VTAIL.n214 9.3005
R2129 VTAIL.n220 VTAIL.n219 9.3005
R2130 VTAIL.n152 VTAIL.n151 9.3005
R2131 VTAIL.n111 VTAIL.n110 9.3005
R2132 VTAIL.n158 VTAIL.n157 9.3005
R2133 VTAIL.n160 VTAIL.n159 9.3005
R2134 VTAIL.n107 VTAIL.n106 9.3005
R2135 VTAIL.n166 VTAIL.n165 9.3005
R2136 VTAIL.n168 VTAIL.n167 9.3005
R2137 VTAIL.n104 VTAIL.n101 9.3005
R2138 VTAIL.n183 VTAIL.n182 9.3005
R2139 VTAIL.n98 VTAIL.n97 9.3005
R2140 VTAIL.n177 VTAIL.n176 9.3005
R2141 VTAIL.n175 VTAIL.n174 9.3005
R2142 VTAIL.n150 VTAIL.n149 9.3005
R2143 VTAIL.n115 VTAIL.n114 9.3005
R2144 VTAIL.n144 VTAIL.n143 9.3005
R2145 VTAIL.n142 VTAIL.n141 9.3005
R2146 VTAIL.n119 VTAIL.n118 9.3005
R2147 VTAIL.n136 VTAIL.n135 9.3005
R2148 VTAIL.n134 VTAIL.n133 9.3005
R2149 VTAIL.n123 VTAIL.n122 9.3005
R2150 VTAIL.n128 VTAIL.n127 9.3005
R2151 VTAIL.n322 VTAIL.n298 8.92171
R2152 VTAIL.n338 VTAIL.n337 8.92171
R2153 VTAIL.n46 VTAIL.n22 8.92171
R2154 VTAIL.n62 VTAIL.n61 8.92171
R2155 VTAIL.n249 VTAIL.n248 8.92171
R2156 VTAIL.n233 VTAIL.n209 8.92171
R2157 VTAIL.n157 VTAIL.n156 8.92171
R2158 VTAIL.n141 VTAIL.n117 8.92171
R2159 VTAIL.n326 VTAIL.n325 8.14595
R2160 VTAIL.n334 VTAIL.n292 8.14595
R2161 VTAIL.n50 VTAIL.n49 8.14595
R2162 VTAIL.n58 VTAIL.n16 8.14595
R2163 VTAIL.n245 VTAIL.n203 8.14595
R2164 VTAIL.n237 VTAIL.n236 8.14595
R2165 VTAIL.n153 VTAIL.n111 8.14595
R2166 VTAIL.n145 VTAIL.n144 8.14595
R2167 VTAIL.n329 VTAIL.n296 7.3702
R2168 VTAIL.n333 VTAIL.n294 7.3702
R2169 VTAIL.n53 VTAIL.n20 7.3702
R2170 VTAIL.n57 VTAIL.n18 7.3702
R2171 VTAIL.n244 VTAIL.n205 7.3702
R2172 VTAIL.n240 VTAIL.n207 7.3702
R2173 VTAIL.n152 VTAIL.n113 7.3702
R2174 VTAIL.n148 VTAIL.n115 7.3702
R2175 VTAIL.n330 VTAIL.n329 6.59444
R2176 VTAIL.n330 VTAIL.n294 6.59444
R2177 VTAIL.n54 VTAIL.n53 6.59444
R2178 VTAIL.n54 VTAIL.n18 6.59444
R2179 VTAIL.n241 VTAIL.n205 6.59444
R2180 VTAIL.n241 VTAIL.n240 6.59444
R2181 VTAIL.n149 VTAIL.n113 6.59444
R2182 VTAIL.n149 VTAIL.n148 6.59444
R2183 VTAIL.n326 VTAIL.n296 5.81868
R2184 VTAIL.n334 VTAIL.n333 5.81868
R2185 VTAIL.n50 VTAIL.n20 5.81868
R2186 VTAIL.n58 VTAIL.n57 5.81868
R2187 VTAIL.n245 VTAIL.n244 5.81868
R2188 VTAIL.n237 VTAIL.n207 5.81868
R2189 VTAIL.n153 VTAIL.n152 5.81868
R2190 VTAIL.n145 VTAIL.n115 5.81868
R2191 VTAIL.n325 VTAIL.n298 5.04292
R2192 VTAIL.n337 VTAIL.n292 5.04292
R2193 VTAIL.n49 VTAIL.n22 5.04292
R2194 VTAIL.n61 VTAIL.n16 5.04292
R2195 VTAIL.n248 VTAIL.n203 5.04292
R2196 VTAIL.n236 VTAIL.n209 5.04292
R2197 VTAIL.n156 VTAIL.n111 5.04292
R2198 VTAIL.n144 VTAIL.n117 5.04292
R2199 VTAIL.n308 VTAIL.n307 4.38563
R2200 VTAIL.n32 VTAIL.n31 4.38563
R2201 VTAIL.n219 VTAIL.n218 4.38563
R2202 VTAIL.n127 VTAIL.n126 4.38563
R2203 VTAIL.n322 VTAIL.n321 4.26717
R2204 VTAIL.n338 VTAIL.n290 4.26717
R2205 VTAIL.n46 VTAIL.n45 4.26717
R2206 VTAIL.n62 VTAIL.n14 4.26717
R2207 VTAIL.n249 VTAIL.n201 4.26717
R2208 VTAIL.n233 VTAIL.n232 4.26717
R2209 VTAIL.n157 VTAIL.n109 4.26717
R2210 VTAIL.n141 VTAIL.n140 4.26717
R2211 VTAIL.n318 VTAIL.n300 3.49141
R2212 VTAIL.n342 VTAIL.n341 3.49141
R2213 VTAIL.n366 VTAIL.n278 3.49141
R2214 VTAIL.n42 VTAIL.n24 3.49141
R2215 VTAIL.n66 VTAIL.n65 3.49141
R2216 VTAIL.n90 VTAIL.n2 3.49141
R2217 VTAIL.n276 VTAIL.n188 3.49141
R2218 VTAIL.n253 VTAIL.n252 3.49141
R2219 VTAIL.n229 VTAIL.n211 3.49141
R2220 VTAIL.n184 VTAIL.n96 3.49141
R2221 VTAIL.n161 VTAIL.n160 3.49141
R2222 VTAIL.n137 VTAIL.n119 3.49141
R2223 VTAIL.n317 VTAIL.n302 2.71565
R2224 VTAIL.n345 VTAIL.n288 2.71565
R2225 VTAIL.n364 VTAIL.n363 2.71565
R2226 VTAIL.n41 VTAIL.n26 2.71565
R2227 VTAIL.n69 VTAIL.n12 2.71565
R2228 VTAIL.n88 VTAIL.n87 2.71565
R2229 VTAIL.n274 VTAIL.n273 2.71565
R2230 VTAIL.n256 VTAIL.n199 2.71565
R2231 VTAIL.n228 VTAIL.n213 2.71565
R2232 VTAIL.n182 VTAIL.n181 2.71565
R2233 VTAIL.n164 VTAIL.n107 2.71565
R2234 VTAIL.n136 VTAIL.n121 2.71565
R2235 VTAIL.n185 VTAIL.n95 2.56947
R2236 VTAIL.n277 VTAIL.n187 2.56947
R2237 VTAIL.n93 VTAIL.n91 2.56947
R2238 VTAIL.n314 VTAIL.n313 1.93989
R2239 VTAIL.n346 VTAIL.n286 1.93989
R2240 VTAIL.n360 VTAIL.n280 1.93989
R2241 VTAIL.n38 VTAIL.n37 1.93989
R2242 VTAIL.n70 VTAIL.n10 1.93989
R2243 VTAIL.n84 VTAIL.n4 1.93989
R2244 VTAIL.n270 VTAIL.n190 1.93989
R2245 VTAIL.n257 VTAIL.n197 1.93989
R2246 VTAIL.n225 VTAIL.n224 1.93989
R2247 VTAIL.n178 VTAIL.n98 1.93989
R2248 VTAIL.n165 VTAIL.n105 1.93989
R2249 VTAIL.n133 VTAIL.n132 1.93989
R2250 VTAIL VTAIL.n367 1.86903
R2251 VTAIL.n187 VTAIL.n185 1.75481
R2252 VTAIL.n91 VTAIL.n1 1.75481
R2253 VTAIL.n0 VTAIL.t9 1.22575
R2254 VTAIL.n0 VTAIL.t10 1.22575
R2255 VTAIL.n92 VTAIL.t2 1.22575
R2256 VTAIL.n92 VTAIL.t3 1.22575
R2257 VTAIL.n186 VTAIL.t5 1.22575
R2258 VTAIL.n186 VTAIL.t0 1.22575
R2259 VTAIL.n94 VTAIL.t6 1.22575
R2260 VTAIL.n94 VTAIL.t7 1.22575
R2261 VTAIL.n310 VTAIL.n304 1.16414
R2262 VTAIL.n351 VTAIL.n349 1.16414
R2263 VTAIL.n359 VTAIL.n282 1.16414
R2264 VTAIL.n34 VTAIL.n28 1.16414
R2265 VTAIL.n75 VTAIL.n73 1.16414
R2266 VTAIL.n83 VTAIL.n6 1.16414
R2267 VTAIL.n269 VTAIL.n192 1.16414
R2268 VTAIL.n261 VTAIL.n260 1.16414
R2269 VTAIL.n221 VTAIL.n215 1.16414
R2270 VTAIL.n177 VTAIL.n100 1.16414
R2271 VTAIL.n169 VTAIL.n168 1.16414
R2272 VTAIL.n129 VTAIL.n123 1.16414
R2273 VTAIL VTAIL.n1 0.700931
R2274 VTAIL.n309 VTAIL.n306 0.388379
R2275 VTAIL.n350 VTAIL.n284 0.388379
R2276 VTAIL.n356 VTAIL.n355 0.388379
R2277 VTAIL.n33 VTAIL.n30 0.388379
R2278 VTAIL.n74 VTAIL.n8 0.388379
R2279 VTAIL.n80 VTAIL.n79 0.388379
R2280 VTAIL.n266 VTAIL.n265 0.388379
R2281 VTAIL.n196 VTAIL.n194 0.388379
R2282 VTAIL.n220 VTAIL.n217 0.388379
R2283 VTAIL.n174 VTAIL.n173 0.388379
R2284 VTAIL.n104 VTAIL.n102 0.388379
R2285 VTAIL.n128 VTAIL.n125 0.388379
R2286 VTAIL.n308 VTAIL.n303 0.155672
R2287 VTAIL.n315 VTAIL.n303 0.155672
R2288 VTAIL.n316 VTAIL.n315 0.155672
R2289 VTAIL.n316 VTAIL.n299 0.155672
R2290 VTAIL.n323 VTAIL.n299 0.155672
R2291 VTAIL.n324 VTAIL.n323 0.155672
R2292 VTAIL.n324 VTAIL.n295 0.155672
R2293 VTAIL.n331 VTAIL.n295 0.155672
R2294 VTAIL.n332 VTAIL.n331 0.155672
R2295 VTAIL.n332 VTAIL.n291 0.155672
R2296 VTAIL.n339 VTAIL.n291 0.155672
R2297 VTAIL.n340 VTAIL.n339 0.155672
R2298 VTAIL.n340 VTAIL.n287 0.155672
R2299 VTAIL.n347 VTAIL.n287 0.155672
R2300 VTAIL.n348 VTAIL.n347 0.155672
R2301 VTAIL.n348 VTAIL.n283 0.155672
R2302 VTAIL.n357 VTAIL.n283 0.155672
R2303 VTAIL.n358 VTAIL.n357 0.155672
R2304 VTAIL.n358 VTAIL.n279 0.155672
R2305 VTAIL.n365 VTAIL.n279 0.155672
R2306 VTAIL.n32 VTAIL.n27 0.155672
R2307 VTAIL.n39 VTAIL.n27 0.155672
R2308 VTAIL.n40 VTAIL.n39 0.155672
R2309 VTAIL.n40 VTAIL.n23 0.155672
R2310 VTAIL.n47 VTAIL.n23 0.155672
R2311 VTAIL.n48 VTAIL.n47 0.155672
R2312 VTAIL.n48 VTAIL.n19 0.155672
R2313 VTAIL.n55 VTAIL.n19 0.155672
R2314 VTAIL.n56 VTAIL.n55 0.155672
R2315 VTAIL.n56 VTAIL.n15 0.155672
R2316 VTAIL.n63 VTAIL.n15 0.155672
R2317 VTAIL.n64 VTAIL.n63 0.155672
R2318 VTAIL.n64 VTAIL.n11 0.155672
R2319 VTAIL.n71 VTAIL.n11 0.155672
R2320 VTAIL.n72 VTAIL.n71 0.155672
R2321 VTAIL.n72 VTAIL.n7 0.155672
R2322 VTAIL.n81 VTAIL.n7 0.155672
R2323 VTAIL.n82 VTAIL.n81 0.155672
R2324 VTAIL.n82 VTAIL.n3 0.155672
R2325 VTAIL.n89 VTAIL.n3 0.155672
R2326 VTAIL.n275 VTAIL.n189 0.155672
R2327 VTAIL.n268 VTAIL.n189 0.155672
R2328 VTAIL.n268 VTAIL.n267 0.155672
R2329 VTAIL.n267 VTAIL.n193 0.155672
R2330 VTAIL.n259 VTAIL.n193 0.155672
R2331 VTAIL.n259 VTAIL.n258 0.155672
R2332 VTAIL.n258 VTAIL.n198 0.155672
R2333 VTAIL.n251 VTAIL.n198 0.155672
R2334 VTAIL.n251 VTAIL.n250 0.155672
R2335 VTAIL.n250 VTAIL.n202 0.155672
R2336 VTAIL.n243 VTAIL.n202 0.155672
R2337 VTAIL.n243 VTAIL.n242 0.155672
R2338 VTAIL.n242 VTAIL.n206 0.155672
R2339 VTAIL.n235 VTAIL.n206 0.155672
R2340 VTAIL.n235 VTAIL.n234 0.155672
R2341 VTAIL.n234 VTAIL.n210 0.155672
R2342 VTAIL.n227 VTAIL.n210 0.155672
R2343 VTAIL.n227 VTAIL.n226 0.155672
R2344 VTAIL.n226 VTAIL.n214 0.155672
R2345 VTAIL.n219 VTAIL.n214 0.155672
R2346 VTAIL.n183 VTAIL.n97 0.155672
R2347 VTAIL.n176 VTAIL.n97 0.155672
R2348 VTAIL.n176 VTAIL.n175 0.155672
R2349 VTAIL.n175 VTAIL.n101 0.155672
R2350 VTAIL.n167 VTAIL.n101 0.155672
R2351 VTAIL.n167 VTAIL.n166 0.155672
R2352 VTAIL.n166 VTAIL.n106 0.155672
R2353 VTAIL.n159 VTAIL.n106 0.155672
R2354 VTAIL.n159 VTAIL.n158 0.155672
R2355 VTAIL.n158 VTAIL.n110 0.155672
R2356 VTAIL.n151 VTAIL.n110 0.155672
R2357 VTAIL.n151 VTAIL.n150 0.155672
R2358 VTAIL.n150 VTAIL.n114 0.155672
R2359 VTAIL.n143 VTAIL.n114 0.155672
R2360 VTAIL.n143 VTAIL.n142 0.155672
R2361 VTAIL.n142 VTAIL.n118 0.155672
R2362 VTAIL.n135 VTAIL.n118 0.155672
R2363 VTAIL.n135 VTAIL.n134 0.155672
R2364 VTAIL.n134 VTAIL.n122 0.155672
R2365 VTAIL.n127 VTAIL.n122 0.155672
R2366 VDD2.n175 VDD2.n91 289.615
R2367 VDD2.n84 VDD2.n0 289.615
R2368 VDD2.n176 VDD2.n175 185
R2369 VDD2.n174 VDD2.n173 185
R2370 VDD2.n95 VDD2.n94 185
R2371 VDD2.n168 VDD2.n167 185
R2372 VDD2.n166 VDD2.n97 185
R2373 VDD2.n165 VDD2.n164 185
R2374 VDD2.n100 VDD2.n98 185
R2375 VDD2.n159 VDD2.n158 185
R2376 VDD2.n157 VDD2.n156 185
R2377 VDD2.n104 VDD2.n103 185
R2378 VDD2.n151 VDD2.n150 185
R2379 VDD2.n149 VDD2.n148 185
R2380 VDD2.n108 VDD2.n107 185
R2381 VDD2.n143 VDD2.n142 185
R2382 VDD2.n141 VDD2.n140 185
R2383 VDD2.n112 VDD2.n111 185
R2384 VDD2.n135 VDD2.n134 185
R2385 VDD2.n133 VDD2.n132 185
R2386 VDD2.n116 VDD2.n115 185
R2387 VDD2.n127 VDD2.n126 185
R2388 VDD2.n125 VDD2.n124 185
R2389 VDD2.n120 VDD2.n119 185
R2390 VDD2.n28 VDD2.n27 185
R2391 VDD2.n33 VDD2.n32 185
R2392 VDD2.n35 VDD2.n34 185
R2393 VDD2.n24 VDD2.n23 185
R2394 VDD2.n41 VDD2.n40 185
R2395 VDD2.n43 VDD2.n42 185
R2396 VDD2.n20 VDD2.n19 185
R2397 VDD2.n49 VDD2.n48 185
R2398 VDD2.n51 VDD2.n50 185
R2399 VDD2.n16 VDD2.n15 185
R2400 VDD2.n57 VDD2.n56 185
R2401 VDD2.n59 VDD2.n58 185
R2402 VDD2.n12 VDD2.n11 185
R2403 VDD2.n65 VDD2.n64 185
R2404 VDD2.n67 VDD2.n66 185
R2405 VDD2.n8 VDD2.n7 185
R2406 VDD2.n74 VDD2.n73 185
R2407 VDD2.n75 VDD2.n6 185
R2408 VDD2.n77 VDD2.n76 185
R2409 VDD2.n4 VDD2.n3 185
R2410 VDD2.n83 VDD2.n82 185
R2411 VDD2.n85 VDD2.n84 185
R2412 VDD2.n121 VDD2.t1 147.659
R2413 VDD2.n29 VDD2.t5 147.659
R2414 VDD2.n175 VDD2.n174 104.615
R2415 VDD2.n174 VDD2.n94 104.615
R2416 VDD2.n167 VDD2.n94 104.615
R2417 VDD2.n167 VDD2.n166 104.615
R2418 VDD2.n166 VDD2.n165 104.615
R2419 VDD2.n165 VDD2.n98 104.615
R2420 VDD2.n158 VDD2.n98 104.615
R2421 VDD2.n158 VDD2.n157 104.615
R2422 VDD2.n157 VDD2.n103 104.615
R2423 VDD2.n150 VDD2.n103 104.615
R2424 VDD2.n150 VDD2.n149 104.615
R2425 VDD2.n149 VDD2.n107 104.615
R2426 VDD2.n142 VDD2.n107 104.615
R2427 VDD2.n142 VDD2.n141 104.615
R2428 VDD2.n141 VDD2.n111 104.615
R2429 VDD2.n134 VDD2.n111 104.615
R2430 VDD2.n134 VDD2.n133 104.615
R2431 VDD2.n133 VDD2.n115 104.615
R2432 VDD2.n126 VDD2.n115 104.615
R2433 VDD2.n126 VDD2.n125 104.615
R2434 VDD2.n125 VDD2.n119 104.615
R2435 VDD2.n33 VDD2.n27 104.615
R2436 VDD2.n34 VDD2.n33 104.615
R2437 VDD2.n34 VDD2.n23 104.615
R2438 VDD2.n41 VDD2.n23 104.615
R2439 VDD2.n42 VDD2.n41 104.615
R2440 VDD2.n42 VDD2.n19 104.615
R2441 VDD2.n49 VDD2.n19 104.615
R2442 VDD2.n50 VDD2.n49 104.615
R2443 VDD2.n50 VDD2.n15 104.615
R2444 VDD2.n57 VDD2.n15 104.615
R2445 VDD2.n58 VDD2.n57 104.615
R2446 VDD2.n58 VDD2.n11 104.615
R2447 VDD2.n65 VDD2.n11 104.615
R2448 VDD2.n66 VDD2.n65 104.615
R2449 VDD2.n66 VDD2.n7 104.615
R2450 VDD2.n74 VDD2.n7 104.615
R2451 VDD2.n75 VDD2.n74 104.615
R2452 VDD2.n76 VDD2.n75 104.615
R2453 VDD2.n76 VDD2.n3 104.615
R2454 VDD2.n83 VDD2.n3 104.615
R2455 VDD2.n84 VDD2.n83 104.615
R2456 VDD2.n90 VDD2.n89 62.916
R2457 VDD2 VDD2.n181 62.9131
R2458 VDD2.t1 VDD2.n119 52.3082
R2459 VDD2.t5 VDD2.n27 52.3082
R2460 VDD2.n90 VDD2.n88 52.287
R2461 VDD2.n180 VDD2.n179 50.4157
R2462 VDD2.n180 VDD2.n90 45.9955
R2463 VDD2.n121 VDD2.n120 15.6677
R2464 VDD2.n29 VDD2.n28 15.6677
R2465 VDD2.n168 VDD2.n97 13.1884
R2466 VDD2.n77 VDD2.n6 13.1884
R2467 VDD2.n169 VDD2.n95 12.8005
R2468 VDD2.n164 VDD2.n99 12.8005
R2469 VDD2.n124 VDD2.n123 12.8005
R2470 VDD2.n32 VDD2.n31 12.8005
R2471 VDD2.n73 VDD2.n72 12.8005
R2472 VDD2.n78 VDD2.n4 12.8005
R2473 VDD2.n173 VDD2.n172 12.0247
R2474 VDD2.n163 VDD2.n100 12.0247
R2475 VDD2.n127 VDD2.n118 12.0247
R2476 VDD2.n35 VDD2.n26 12.0247
R2477 VDD2.n71 VDD2.n8 12.0247
R2478 VDD2.n82 VDD2.n81 12.0247
R2479 VDD2.n176 VDD2.n93 11.249
R2480 VDD2.n160 VDD2.n159 11.249
R2481 VDD2.n128 VDD2.n116 11.249
R2482 VDD2.n36 VDD2.n24 11.249
R2483 VDD2.n68 VDD2.n67 11.249
R2484 VDD2.n85 VDD2.n2 11.249
R2485 VDD2.n177 VDD2.n91 10.4732
R2486 VDD2.n156 VDD2.n102 10.4732
R2487 VDD2.n132 VDD2.n131 10.4732
R2488 VDD2.n40 VDD2.n39 10.4732
R2489 VDD2.n64 VDD2.n10 10.4732
R2490 VDD2.n86 VDD2.n0 10.4732
R2491 VDD2.n155 VDD2.n104 9.69747
R2492 VDD2.n135 VDD2.n114 9.69747
R2493 VDD2.n43 VDD2.n22 9.69747
R2494 VDD2.n63 VDD2.n12 9.69747
R2495 VDD2.n179 VDD2.n178 9.45567
R2496 VDD2.n88 VDD2.n87 9.45567
R2497 VDD2.n147 VDD2.n146 9.3005
R2498 VDD2.n106 VDD2.n105 9.3005
R2499 VDD2.n153 VDD2.n152 9.3005
R2500 VDD2.n155 VDD2.n154 9.3005
R2501 VDD2.n102 VDD2.n101 9.3005
R2502 VDD2.n161 VDD2.n160 9.3005
R2503 VDD2.n163 VDD2.n162 9.3005
R2504 VDD2.n99 VDD2.n96 9.3005
R2505 VDD2.n178 VDD2.n177 9.3005
R2506 VDD2.n93 VDD2.n92 9.3005
R2507 VDD2.n172 VDD2.n171 9.3005
R2508 VDD2.n170 VDD2.n169 9.3005
R2509 VDD2.n145 VDD2.n144 9.3005
R2510 VDD2.n110 VDD2.n109 9.3005
R2511 VDD2.n139 VDD2.n138 9.3005
R2512 VDD2.n137 VDD2.n136 9.3005
R2513 VDD2.n114 VDD2.n113 9.3005
R2514 VDD2.n131 VDD2.n130 9.3005
R2515 VDD2.n129 VDD2.n128 9.3005
R2516 VDD2.n118 VDD2.n117 9.3005
R2517 VDD2.n123 VDD2.n122 9.3005
R2518 VDD2.n87 VDD2.n86 9.3005
R2519 VDD2.n2 VDD2.n1 9.3005
R2520 VDD2.n81 VDD2.n80 9.3005
R2521 VDD2.n79 VDD2.n78 9.3005
R2522 VDD2.n18 VDD2.n17 9.3005
R2523 VDD2.n47 VDD2.n46 9.3005
R2524 VDD2.n45 VDD2.n44 9.3005
R2525 VDD2.n22 VDD2.n21 9.3005
R2526 VDD2.n39 VDD2.n38 9.3005
R2527 VDD2.n37 VDD2.n36 9.3005
R2528 VDD2.n26 VDD2.n25 9.3005
R2529 VDD2.n31 VDD2.n30 9.3005
R2530 VDD2.n53 VDD2.n52 9.3005
R2531 VDD2.n55 VDD2.n54 9.3005
R2532 VDD2.n14 VDD2.n13 9.3005
R2533 VDD2.n61 VDD2.n60 9.3005
R2534 VDD2.n63 VDD2.n62 9.3005
R2535 VDD2.n10 VDD2.n9 9.3005
R2536 VDD2.n69 VDD2.n68 9.3005
R2537 VDD2.n71 VDD2.n70 9.3005
R2538 VDD2.n72 VDD2.n5 9.3005
R2539 VDD2.n152 VDD2.n151 8.92171
R2540 VDD2.n136 VDD2.n112 8.92171
R2541 VDD2.n44 VDD2.n20 8.92171
R2542 VDD2.n60 VDD2.n59 8.92171
R2543 VDD2.n148 VDD2.n106 8.14595
R2544 VDD2.n140 VDD2.n139 8.14595
R2545 VDD2.n48 VDD2.n47 8.14595
R2546 VDD2.n56 VDD2.n14 8.14595
R2547 VDD2.n147 VDD2.n108 7.3702
R2548 VDD2.n143 VDD2.n110 7.3702
R2549 VDD2.n51 VDD2.n18 7.3702
R2550 VDD2.n55 VDD2.n16 7.3702
R2551 VDD2.n144 VDD2.n108 6.59444
R2552 VDD2.n144 VDD2.n143 6.59444
R2553 VDD2.n52 VDD2.n51 6.59444
R2554 VDD2.n52 VDD2.n16 6.59444
R2555 VDD2.n148 VDD2.n147 5.81868
R2556 VDD2.n140 VDD2.n110 5.81868
R2557 VDD2.n48 VDD2.n18 5.81868
R2558 VDD2.n56 VDD2.n55 5.81868
R2559 VDD2.n151 VDD2.n106 5.04292
R2560 VDD2.n139 VDD2.n112 5.04292
R2561 VDD2.n47 VDD2.n20 5.04292
R2562 VDD2.n59 VDD2.n14 5.04292
R2563 VDD2.n122 VDD2.n121 4.38563
R2564 VDD2.n30 VDD2.n29 4.38563
R2565 VDD2.n152 VDD2.n104 4.26717
R2566 VDD2.n136 VDD2.n135 4.26717
R2567 VDD2.n44 VDD2.n43 4.26717
R2568 VDD2.n60 VDD2.n12 4.26717
R2569 VDD2.n179 VDD2.n91 3.49141
R2570 VDD2.n156 VDD2.n155 3.49141
R2571 VDD2.n132 VDD2.n114 3.49141
R2572 VDD2.n40 VDD2.n22 3.49141
R2573 VDD2.n64 VDD2.n63 3.49141
R2574 VDD2.n88 VDD2.n0 3.49141
R2575 VDD2.n177 VDD2.n176 2.71565
R2576 VDD2.n159 VDD2.n102 2.71565
R2577 VDD2.n131 VDD2.n116 2.71565
R2578 VDD2.n39 VDD2.n24 2.71565
R2579 VDD2.n67 VDD2.n10 2.71565
R2580 VDD2.n86 VDD2.n85 2.71565
R2581 VDD2 VDD2.n180 1.98541
R2582 VDD2.n173 VDD2.n93 1.93989
R2583 VDD2.n160 VDD2.n100 1.93989
R2584 VDD2.n128 VDD2.n127 1.93989
R2585 VDD2.n36 VDD2.n35 1.93989
R2586 VDD2.n68 VDD2.n8 1.93989
R2587 VDD2.n82 VDD2.n2 1.93989
R2588 VDD2.n181 VDD2.t4 1.22575
R2589 VDD2.n181 VDD2.t2 1.22575
R2590 VDD2.n89 VDD2.t0 1.22575
R2591 VDD2.n89 VDD2.t3 1.22575
R2592 VDD2.n172 VDD2.n95 1.16414
R2593 VDD2.n164 VDD2.n163 1.16414
R2594 VDD2.n124 VDD2.n118 1.16414
R2595 VDD2.n32 VDD2.n26 1.16414
R2596 VDD2.n73 VDD2.n71 1.16414
R2597 VDD2.n81 VDD2.n4 1.16414
R2598 VDD2.n169 VDD2.n168 0.388379
R2599 VDD2.n99 VDD2.n97 0.388379
R2600 VDD2.n123 VDD2.n120 0.388379
R2601 VDD2.n31 VDD2.n28 0.388379
R2602 VDD2.n72 VDD2.n6 0.388379
R2603 VDD2.n78 VDD2.n77 0.388379
R2604 VDD2.n178 VDD2.n92 0.155672
R2605 VDD2.n171 VDD2.n92 0.155672
R2606 VDD2.n171 VDD2.n170 0.155672
R2607 VDD2.n170 VDD2.n96 0.155672
R2608 VDD2.n162 VDD2.n96 0.155672
R2609 VDD2.n162 VDD2.n161 0.155672
R2610 VDD2.n161 VDD2.n101 0.155672
R2611 VDD2.n154 VDD2.n101 0.155672
R2612 VDD2.n154 VDD2.n153 0.155672
R2613 VDD2.n153 VDD2.n105 0.155672
R2614 VDD2.n146 VDD2.n105 0.155672
R2615 VDD2.n146 VDD2.n145 0.155672
R2616 VDD2.n145 VDD2.n109 0.155672
R2617 VDD2.n138 VDD2.n109 0.155672
R2618 VDD2.n138 VDD2.n137 0.155672
R2619 VDD2.n137 VDD2.n113 0.155672
R2620 VDD2.n130 VDD2.n113 0.155672
R2621 VDD2.n130 VDD2.n129 0.155672
R2622 VDD2.n129 VDD2.n117 0.155672
R2623 VDD2.n122 VDD2.n117 0.155672
R2624 VDD2.n30 VDD2.n25 0.155672
R2625 VDD2.n37 VDD2.n25 0.155672
R2626 VDD2.n38 VDD2.n37 0.155672
R2627 VDD2.n38 VDD2.n21 0.155672
R2628 VDD2.n45 VDD2.n21 0.155672
R2629 VDD2.n46 VDD2.n45 0.155672
R2630 VDD2.n46 VDD2.n17 0.155672
R2631 VDD2.n53 VDD2.n17 0.155672
R2632 VDD2.n54 VDD2.n53 0.155672
R2633 VDD2.n54 VDD2.n13 0.155672
R2634 VDD2.n61 VDD2.n13 0.155672
R2635 VDD2.n62 VDD2.n61 0.155672
R2636 VDD2.n62 VDD2.n9 0.155672
R2637 VDD2.n69 VDD2.n9 0.155672
R2638 VDD2.n70 VDD2.n69 0.155672
R2639 VDD2.n70 VDD2.n5 0.155672
R2640 VDD2.n79 VDD2.n5 0.155672
R2641 VDD2.n80 VDD2.n79 0.155672
R2642 VDD2.n80 VDD2.n1 0.155672
R2643 VDD2.n87 VDD2.n1 0.155672
R2644 VP.n11 VP.t1 181
R2645 VP.n13 VP.n12 161.3
R2646 VP.n14 VP.n9 161.3
R2647 VP.n16 VP.n15 161.3
R2648 VP.n17 VP.n8 161.3
R2649 VP.n19 VP.n18 161.3
R2650 VP.n20 VP.n7 161.3
R2651 VP.n42 VP.n0 161.3
R2652 VP.n41 VP.n40 161.3
R2653 VP.n39 VP.n1 161.3
R2654 VP.n38 VP.n37 161.3
R2655 VP.n36 VP.n2 161.3
R2656 VP.n35 VP.n34 161.3
R2657 VP.n33 VP.n32 161.3
R2658 VP.n31 VP.n4 161.3
R2659 VP.n30 VP.n29 161.3
R2660 VP.n28 VP.n5 161.3
R2661 VP.n27 VP.n26 161.3
R2662 VP.n25 VP.n6 161.3
R2663 VP.n24 VP.t2 146.965
R2664 VP.n3 VP.t4 146.965
R2665 VP.n43 VP.t5 146.965
R2666 VP.n21 VP.t0 146.965
R2667 VP.n10 VP.t3 146.965
R2668 VP.n24 VP.n23 99.596
R2669 VP.n44 VP.n43 99.596
R2670 VP.n22 VP.n21 99.596
R2671 VP.n11 VP.n10 60.4656
R2672 VP.n37 VP.n1 56.5617
R2673 VP.n30 VP.n5 56.5617
R2674 VP.n15 VP.n8 56.5617
R2675 VP.n23 VP.n22 52.0754
R2676 VP.n26 VP.n25 24.5923
R2677 VP.n26 VP.n5 24.5923
R2678 VP.n31 VP.n30 24.5923
R2679 VP.n32 VP.n31 24.5923
R2680 VP.n36 VP.n35 24.5923
R2681 VP.n37 VP.n36 24.5923
R2682 VP.n41 VP.n1 24.5923
R2683 VP.n42 VP.n41 24.5923
R2684 VP.n19 VP.n8 24.5923
R2685 VP.n20 VP.n19 24.5923
R2686 VP.n14 VP.n13 24.5923
R2687 VP.n15 VP.n14 24.5923
R2688 VP.n32 VP.n3 12.2964
R2689 VP.n35 VP.n3 12.2964
R2690 VP.n13 VP.n10 12.2964
R2691 VP.n25 VP.n24 11.3127
R2692 VP.n43 VP.n42 11.3127
R2693 VP.n21 VP.n20 11.3127
R2694 VP.n12 VP.n11 6.75133
R2695 VP.n22 VP.n7 0.278335
R2696 VP.n23 VP.n6 0.278335
R2697 VP.n44 VP.n0 0.278335
R2698 VP.n12 VP.n9 0.189894
R2699 VP.n16 VP.n9 0.189894
R2700 VP.n17 VP.n16 0.189894
R2701 VP.n18 VP.n17 0.189894
R2702 VP.n18 VP.n7 0.189894
R2703 VP.n27 VP.n6 0.189894
R2704 VP.n28 VP.n27 0.189894
R2705 VP.n29 VP.n28 0.189894
R2706 VP.n29 VP.n4 0.189894
R2707 VP.n33 VP.n4 0.189894
R2708 VP.n34 VP.n33 0.189894
R2709 VP.n34 VP.n2 0.189894
R2710 VP.n38 VP.n2 0.189894
R2711 VP.n39 VP.n38 0.189894
R2712 VP.n40 VP.n39 0.189894
R2713 VP.n40 VP.n0 0.189894
R2714 VP VP.n44 0.153485
R2715 VDD1.n84 VDD1.n0 289.615
R2716 VDD1.n173 VDD1.n89 289.615
R2717 VDD1.n85 VDD1.n84 185
R2718 VDD1.n83 VDD1.n82 185
R2719 VDD1.n4 VDD1.n3 185
R2720 VDD1.n77 VDD1.n76 185
R2721 VDD1.n75 VDD1.n6 185
R2722 VDD1.n74 VDD1.n73 185
R2723 VDD1.n9 VDD1.n7 185
R2724 VDD1.n68 VDD1.n67 185
R2725 VDD1.n66 VDD1.n65 185
R2726 VDD1.n13 VDD1.n12 185
R2727 VDD1.n60 VDD1.n59 185
R2728 VDD1.n58 VDD1.n57 185
R2729 VDD1.n17 VDD1.n16 185
R2730 VDD1.n52 VDD1.n51 185
R2731 VDD1.n50 VDD1.n49 185
R2732 VDD1.n21 VDD1.n20 185
R2733 VDD1.n44 VDD1.n43 185
R2734 VDD1.n42 VDD1.n41 185
R2735 VDD1.n25 VDD1.n24 185
R2736 VDD1.n36 VDD1.n35 185
R2737 VDD1.n34 VDD1.n33 185
R2738 VDD1.n29 VDD1.n28 185
R2739 VDD1.n117 VDD1.n116 185
R2740 VDD1.n122 VDD1.n121 185
R2741 VDD1.n124 VDD1.n123 185
R2742 VDD1.n113 VDD1.n112 185
R2743 VDD1.n130 VDD1.n129 185
R2744 VDD1.n132 VDD1.n131 185
R2745 VDD1.n109 VDD1.n108 185
R2746 VDD1.n138 VDD1.n137 185
R2747 VDD1.n140 VDD1.n139 185
R2748 VDD1.n105 VDD1.n104 185
R2749 VDD1.n146 VDD1.n145 185
R2750 VDD1.n148 VDD1.n147 185
R2751 VDD1.n101 VDD1.n100 185
R2752 VDD1.n154 VDD1.n153 185
R2753 VDD1.n156 VDD1.n155 185
R2754 VDD1.n97 VDD1.n96 185
R2755 VDD1.n163 VDD1.n162 185
R2756 VDD1.n164 VDD1.n95 185
R2757 VDD1.n166 VDD1.n165 185
R2758 VDD1.n93 VDD1.n92 185
R2759 VDD1.n172 VDD1.n171 185
R2760 VDD1.n174 VDD1.n173 185
R2761 VDD1.n30 VDD1.t4 147.659
R2762 VDD1.n118 VDD1.t3 147.659
R2763 VDD1.n84 VDD1.n83 104.615
R2764 VDD1.n83 VDD1.n3 104.615
R2765 VDD1.n76 VDD1.n3 104.615
R2766 VDD1.n76 VDD1.n75 104.615
R2767 VDD1.n75 VDD1.n74 104.615
R2768 VDD1.n74 VDD1.n7 104.615
R2769 VDD1.n67 VDD1.n7 104.615
R2770 VDD1.n67 VDD1.n66 104.615
R2771 VDD1.n66 VDD1.n12 104.615
R2772 VDD1.n59 VDD1.n12 104.615
R2773 VDD1.n59 VDD1.n58 104.615
R2774 VDD1.n58 VDD1.n16 104.615
R2775 VDD1.n51 VDD1.n16 104.615
R2776 VDD1.n51 VDD1.n50 104.615
R2777 VDD1.n50 VDD1.n20 104.615
R2778 VDD1.n43 VDD1.n20 104.615
R2779 VDD1.n43 VDD1.n42 104.615
R2780 VDD1.n42 VDD1.n24 104.615
R2781 VDD1.n35 VDD1.n24 104.615
R2782 VDD1.n35 VDD1.n34 104.615
R2783 VDD1.n34 VDD1.n28 104.615
R2784 VDD1.n122 VDD1.n116 104.615
R2785 VDD1.n123 VDD1.n122 104.615
R2786 VDD1.n123 VDD1.n112 104.615
R2787 VDD1.n130 VDD1.n112 104.615
R2788 VDD1.n131 VDD1.n130 104.615
R2789 VDD1.n131 VDD1.n108 104.615
R2790 VDD1.n138 VDD1.n108 104.615
R2791 VDD1.n139 VDD1.n138 104.615
R2792 VDD1.n139 VDD1.n104 104.615
R2793 VDD1.n146 VDD1.n104 104.615
R2794 VDD1.n147 VDD1.n146 104.615
R2795 VDD1.n147 VDD1.n100 104.615
R2796 VDD1.n154 VDD1.n100 104.615
R2797 VDD1.n155 VDD1.n154 104.615
R2798 VDD1.n155 VDD1.n96 104.615
R2799 VDD1.n163 VDD1.n96 104.615
R2800 VDD1.n164 VDD1.n163 104.615
R2801 VDD1.n165 VDD1.n164 104.615
R2802 VDD1.n165 VDD1.n92 104.615
R2803 VDD1.n172 VDD1.n92 104.615
R2804 VDD1.n173 VDD1.n172 104.615
R2805 VDD1.n179 VDD1.n178 62.916
R2806 VDD1.n181 VDD1.n180 62.3291
R2807 VDD1 VDD1.n88 52.4006
R2808 VDD1.t4 VDD1.n28 52.3082
R2809 VDD1.t3 VDD1.n116 52.3082
R2810 VDD1.n179 VDD1.n177 52.287
R2811 VDD1.n181 VDD1.n179 47.863
R2812 VDD1.n30 VDD1.n29 15.6677
R2813 VDD1.n118 VDD1.n117 15.6677
R2814 VDD1.n77 VDD1.n6 13.1884
R2815 VDD1.n166 VDD1.n95 13.1884
R2816 VDD1.n78 VDD1.n4 12.8005
R2817 VDD1.n73 VDD1.n8 12.8005
R2818 VDD1.n33 VDD1.n32 12.8005
R2819 VDD1.n121 VDD1.n120 12.8005
R2820 VDD1.n162 VDD1.n161 12.8005
R2821 VDD1.n167 VDD1.n93 12.8005
R2822 VDD1.n82 VDD1.n81 12.0247
R2823 VDD1.n72 VDD1.n9 12.0247
R2824 VDD1.n36 VDD1.n27 12.0247
R2825 VDD1.n124 VDD1.n115 12.0247
R2826 VDD1.n160 VDD1.n97 12.0247
R2827 VDD1.n171 VDD1.n170 12.0247
R2828 VDD1.n85 VDD1.n2 11.249
R2829 VDD1.n69 VDD1.n68 11.249
R2830 VDD1.n37 VDD1.n25 11.249
R2831 VDD1.n125 VDD1.n113 11.249
R2832 VDD1.n157 VDD1.n156 11.249
R2833 VDD1.n174 VDD1.n91 11.249
R2834 VDD1.n86 VDD1.n0 10.4732
R2835 VDD1.n65 VDD1.n11 10.4732
R2836 VDD1.n41 VDD1.n40 10.4732
R2837 VDD1.n129 VDD1.n128 10.4732
R2838 VDD1.n153 VDD1.n99 10.4732
R2839 VDD1.n175 VDD1.n89 10.4732
R2840 VDD1.n64 VDD1.n13 9.69747
R2841 VDD1.n44 VDD1.n23 9.69747
R2842 VDD1.n132 VDD1.n111 9.69747
R2843 VDD1.n152 VDD1.n101 9.69747
R2844 VDD1.n88 VDD1.n87 9.45567
R2845 VDD1.n177 VDD1.n176 9.45567
R2846 VDD1.n56 VDD1.n55 9.3005
R2847 VDD1.n15 VDD1.n14 9.3005
R2848 VDD1.n62 VDD1.n61 9.3005
R2849 VDD1.n64 VDD1.n63 9.3005
R2850 VDD1.n11 VDD1.n10 9.3005
R2851 VDD1.n70 VDD1.n69 9.3005
R2852 VDD1.n72 VDD1.n71 9.3005
R2853 VDD1.n8 VDD1.n5 9.3005
R2854 VDD1.n87 VDD1.n86 9.3005
R2855 VDD1.n2 VDD1.n1 9.3005
R2856 VDD1.n81 VDD1.n80 9.3005
R2857 VDD1.n79 VDD1.n78 9.3005
R2858 VDD1.n54 VDD1.n53 9.3005
R2859 VDD1.n19 VDD1.n18 9.3005
R2860 VDD1.n48 VDD1.n47 9.3005
R2861 VDD1.n46 VDD1.n45 9.3005
R2862 VDD1.n23 VDD1.n22 9.3005
R2863 VDD1.n40 VDD1.n39 9.3005
R2864 VDD1.n38 VDD1.n37 9.3005
R2865 VDD1.n27 VDD1.n26 9.3005
R2866 VDD1.n32 VDD1.n31 9.3005
R2867 VDD1.n176 VDD1.n175 9.3005
R2868 VDD1.n91 VDD1.n90 9.3005
R2869 VDD1.n170 VDD1.n169 9.3005
R2870 VDD1.n168 VDD1.n167 9.3005
R2871 VDD1.n107 VDD1.n106 9.3005
R2872 VDD1.n136 VDD1.n135 9.3005
R2873 VDD1.n134 VDD1.n133 9.3005
R2874 VDD1.n111 VDD1.n110 9.3005
R2875 VDD1.n128 VDD1.n127 9.3005
R2876 VDD1.n126 VDD1.n125 9.3005
R2877 VDD1.n115 VDD1.n114 9.3005
R2878 VDD1.n120 VDD1.n119 9.3005
R2879 VDD1.n142 VDD1.n141 9.3005
R2880 VDD1.n144 VDD1.n143 9.3005
R2881 VDD1.n103 VDD1.n102 9.3005
R2882 VDD1.n150 VDD1.n149 9.3005
R2883 VDD1.n152 VDD1.n151 9.3005
R2884 VDD1.n99 VDD1.n98 9.3005
R2885 VDD1.n158 VDD1.n157 9.3005
R2886 VDD1.n160 VDD1.n159 9.3005
R2887 VDD1.n161 VDD1.n94 9.3005
R2888 VDD1.n61 VDD1.n60 8.92171
R2889 VDD1.n45 VDD1.n21 8.92171
R2890 VDD1.n133 VDD1.n109 8.92171
R2891 VDD1.n149 VDD1.n148 8.92171
R2892 VDD1.n57 VDD1.n15 8.14595
R2893 VDD1.n49 VDD1.n48 8.14595
R2894 VDD1.n137 VDD1.n136 8.14595
R2895 VDD1.n145 VDD1.n103 8.14595
R2896 VDD1.n56 VDD1.n17 7.3702
R2897 VDD1.n52 VDD1.n19 7.3702
R2898 VDD1.n140 VDD1.n107 7.3702
R2899 VDD1.n144 VDD1.n105 7.3702
R2900 VDD1.n53 VDD1.n17 6.59444
R2901 VDD1.n53 VDD1.n52 6.59444
R2902 VDD1.n141 VDD1.n140 6.59444
R2903 VDD1.n141 VDD1.n105 6.59444
R2904 VDD1.n57 VDD1.n56 5.81868
R2905 VDD1.n49 VDD1.n19 5.81868
R2906 VDD1.n137 VDD1.n107 5.81868
R2907 VDD1.n145 VDD1.n144 5.81868
R2908 VDD1.n60 VDD1.n15 5.04292
R2909 VDD1.n48 VDD1.n21 5.04292
R2910 VDD1.n136 VDD1.n109 5.04292
R2911 VDD1.n148 VDD1.n103 5.04292
R2912 VDD1.n31 VDD1.n30 4.38563
R2913 VDD1.n119 VDD1.n118 4.38563
R2914 VDD1.n61 VDD1.n13 4.26717
R2915 VDD1.n45 VDD1.n44 4.26717
R2916 VDD1.n133 VDD1.n132 4.26717
R2917 VDD1.n149 VDD1.n101 4.26717
R2918 VDD1.n88 VDD1.n0 3.49141
R2919 VDD1.n65 VDD1.n64 3.49141
R2920 VDD1.n41 VDD1.n23 3.49141
R2921 VDD1.n129 VDD1.n111 3.49141
R2922 VDD1.n153 VDD1.n152 3.49141
R2923 VDD1.n177 VDD1.n89 3.49141
R2924 VDD1.n86 VDD1.n85 2.71565
R2925 VDD1.n68 VDD1.n11 2.71565
R2926 VDD1.n40 VDD1.n25 2.71565
R2927 VDD1.n128 VDD1.n113 2.71565
R2928 VDD1.n156 VDD1.n99 2.71565
R2929 VDD1.n175 VDD1.n174 2.71565
R2930 VDD1.n82 VDD1.n2 1.93989
R2931 VDD1.n69 VDD1.n9 1.93989
R2932 VDD1.n37 VDD1.n36 1.93989
R2933 VDD1.n125 VDD1.n124 1.93989
R2934 VDD1.n157 VDD1.n97 1.93989
R2935 VDD1.n171 VDD1.n91 1.93989
R2936 VDD1.n180 VDD1.t2 1.22575
R2937 VDD1.n180 VDD1.t5 1.22575
R2938 VDD1.n178 VDD1.t1 1.22575
R2939 VDD1.n178 VDD1.t0 1.22575
R2940 VDD1.n81 VDD1.n4 1.16414
R2941 VDD1.n73 VDD1.n72 1.16414
R2942 VDD1.n33 VDD1.n27 1.16414
R2943 VDD1.n121 VDD1.n115 1.16414
R2944 VDD1.n162 VDD1.n160 1.16414
R2945 VDD1.n170 VDD1.n93 1.16414
R2946 VDD1 VDD1.n181 0.584552
R2947 VDD1.n78 VDD1.n77 0.388379
R2948 VDD1.n8 VDD1.n6 0.388379
R2949 VDD1.n32 VDD1.n29 0.388379
R2950 VDD1.n120 VDD1.n117 0.388379
R2951 VDD1.n161 VDD1.n95 0.388379
R2952 VDD1.n167 VDD1.n166 0.388379
R2953 VDD1.n87 VDD1.n1 0.155672
R2954 VDD1.n80 VDD1.n1 0.155672
R2955 VDD1.n80 VDD1.n79 0.155672
R2956 VDD1.n79 VDD1.n5 0.155672
R2957 VDD1.n71 VDD1.n5 0.155672
R2958 VDD1.n71 VDD1.n70 0.155672
R2959 VDD1.n70 VDD1.n10 0.155672
R2960 VDD1.n63 VDD1.n10 0.155672
R2961 VDD1.n63 VDD1.n62 0.155672
R2962 VDD1.n62 VDD1.n14 0.155672
R2963 VDD1.n55 VDD1.n14 0.155672
R2964 VDD1.n55 VDD1.n54 0.155672
R2965 VDD1.n54 VDD1.n18 0.155672
R2966 VDD1.n47 VDD1.n18 0.155672
R2967 VDD1.n47 VDD1.n46 0.155672
R2968 VDD1.n46 VDD1.n22 0.155672
R2969 VDD1.n39 VDD1.n22 0.155672
R2970 VDD1.n39 VDD1.n38 0.155672
R2971 VDD1.n38 VDD1.n26 0.155672
R2972 VDD1.n31 VDD1.n26 0.155672
R2973 VDD1.n119 VDD1.n114 0.155672
R2974 VDD1.n126 VDD1.n114 0.155672
R2975 VDD1.n127 VDD1.n126 0.155672
R2976 VDD1.n127 VDD1.n110 0.155672
R2977 VDD1.n134 VDD1.n110 0.155672
R2978 VDD1.n135 VDD1.n134 0.155672
R2979 VDD1.n135 VDD1.n106 0.155672
R2980 VDD1.n142 VDD1.n106 0.155672
R2981 VDD1.n143 VDD1.n142 0.155672
R2982 VDD1.n143 VDD1.n102 0.155672
R2983 VDD1.n150 VDD1.n102 0.155672
R2984 VDD1.n151 VDD1.n150 0.155672
R2985 VDD1.n151 VDD1.n98 0.155672
R2986 VDD1.n158 VDD1.n98 0.155672
R2987 VDD1.n159 VDD1.n158 0.155672
R2988 VDD1.n159 VDD1.n94 0.155672
R2989 VDD1.n168 VDD1.n94 0.155672
R2990 VDD1.n169 VDD1.n168 0.155672
R2991 VDD1.n169 VDD1.n90 0.155672
R2992 VDD1.n176 VDD1.n90 0.155672
C0 VTAIL VDD1 9.23654f
C1 VTAIL VP 8.94904f
C2 VDD1 VP 9.2611f
C3 VTAIL VDD2 9.28681f
C4 VTAIL VN 8.93469f
C5 VDD1 VDD2 1.42752f
C6 VDD1 VN 0.151223f
C7 VDD2 VP 0.463301f
C8 VP VN 7.73779f
C9 VDD2 VN 8.95292f
C10 VDD2 B 6.766913f
C11 VDD1 B 6.897519f
C12 VTAIL B 9.512801f
C13 VN B 13.368101f
C14 VP B 11.930395f
C15 VDD1.n0 B 0.029561f
C16 VDD1.n1 B 0.021442f
C17 VDD1.n2 B 0.011522f
C18 VDD1.n3 B 0.027234f
C19 VDD1.n4 B 0.0122f
C20 VDD1.n5 B 0.021442f
C21 VDD1.n6 B 0.011861f
C22 VDD1.n7 B 0.027234f
C23 VDD1.n8 B 0.011522f
C24 VDD1.n9 B 0.0122f
C25 VDD1.n10 B 0.021442f
C26 VDD1.n11 B 0.011522f
C27 VDD1.n12 B 0.027234f
C28 VDD1.n13 B 0.0122f
C29 VDD1.n14 B 0.021442f
C30 VDD1.n15 B 0.011522f
C31 VDD1.n16 B 0.027234f
C32 VDD1.n17 B 0.0122f
C33 VDD1.n18 B 0.021442f
C34 VDD1.n19 B 0.011522f
C35 VDD1.n20 B 0.027234f
C36 VDD1.n21 B 0.0122f
C37 VDD1.n22 B 0.021442f
C38 VDD1.n23 B 0.011522f
C39 VDD1.n24 B 0.027234f
C40 VDD1.n25 B 0.0122f
C41 VDD1.n26 B 0.021442f
C42 VDD1.n27 B 0.011522f
C43 VDD1.n28 B 0.020426f
C44 VDD1.n29 B 0.016088f
C45 VDD1.t4 B 0.044992f
C46 VDD1.n30 B 0.146088f
C47 VDD1.n31 B 1.50907f
C48 VDD1.n32 B 0.011522f
C49 VDD1.n33 B 0.0122f
C50 VDD1.n34 B 0.027234f
C51 VDD1.n35 B 0.027234f
C52 VDD1.n36 B 0.0122f
C53 VDD1.n37 B 0.011522f
C54 VDD1.n38 B 0.021442f
C55 VDD1.n39 B 0.021442f
C56 VDD1.n40 B 0.011522f
C57 VDD1.n41 B 0.0122f
C58 VDD1.n42 B 0.027234f
C59 VDD1.n43 B 0.027234f
C60 VDD1.n44 B 0.0122f
C61 VDD1.n45 B 0.011522f
C62 VDD1.n46 B 0.021442f
C63 VDD1.n47 B 0.021442f
C64 VDD1.n48 B 0.011522f
C65 VDD1.n49 B 0.0122f
C66 VDD1.n50 B 0.027234f
C67 VDD1.n51 B 0.027234f
C68 VDD1.n52 B 0.0122f
C69 VDD1.n53 B 0.011522f
C70 VDD1.n54 B 0.021442f
C71 VDD1.n55 B 0.021442f
C72 VDD1.n56 B 0.011522f
C73 VDD1.n57 B 0.0122f
C74 VDD1.n58 B 0.027234f
C75 VDD1.n59 B 0.027234f
C76 VDD1.n60 B 0.0122f
C77 VDD1.n61 B 0.011522f
C78 VDD1.n62 B 0.021442f
C79 VDD1.n63 B 0.021442f
C80 VDD1.n64 B 0.011522f
C81 VDD1.n65 B 0.0122f
C82 VDD1.n66 B 0.027234f
C83 VDD1.n67 B 0.027234f
C84 VDD1.n68 B 0.0122f
C85 VDD1.n69 B 0.011522f
C86 VDD1.n70 B 0.021442f
C87 VDD1.n71 B 0.021442f
C88 VDD1.n72 B 0.011522f
C89 VDD1.n73 B 0.0122f
C90 VDD1.n74 B 0.027234f
C91 VDD1.n75 B 0.027234f
C92 VDD1.n76 B 0.027234f
C93 VDD1.n77 B 0.011861f
C94 VDD1.n78 B 0.011522f
C95 VDD1.n79 B 0.021442f
C96 VDD1.n80 B 0.021442f
C97 VDD1.n81 B 0.011522f
C98 VDD1.n82 B 0.0122f
C99 VDD1.n83 B 0.027234f
C100 VDD1.n84 B 0.057935f
C101 VDD1.n85 B 0.0122f
C102 VDD1.n86 B 0.011522f
C103 VDD1.n87 B 0.051907f
C104 VDD1.n88 B 0.05398f
C105 VDD1.n89 B 0.029561f
C106 VDD1.n90 B 0.021442f
C107 VDD1.n91 B 0.011522f
C108 VDD1.n92 B 0.027234f
C109 VDD1.n93 B 0.0122f
C110 VDD1.n94 B 0.021442f
C111 VDD1.n95 B 0.011861f
C112 VDD1.n96 B 0.027234f
C113 VDD1.n97 B 0.0122f
C114 VDD1.n98 B 0.021442f
C115 VDD1.n99 B 0.011522f
C116 VDD1.n100 B 0.027234f
C117 VDD1.n101 B 0.0122f
C118 VDD1.n102 B 0.021442f
C119 VDD1.n103 B 0.011522f
C120 VDD1.n104 B 0.027234f
C121 VDD1.n105 B 0.0122f
C122 VDD1.n106 B 0.021442f
C123 VDD1.n107 B 0.011522f
C124 VDD1.n108 B 0.027234f
C125 VDD1.n109 B 0.0122f
C126 VDD1.n110 B 0.021442f
C127 VDD1.n111 B 0.011522f
C128 VDD1.n112 B 0.027234f
C129 VDD1.n113 B 0.0122f
C130 VDD1.n114 B 0.021442f
C131 VDD1.n115 B 0.011522f
C132 VDD1.n116 B 0.020426f
C133 VDD1.n117 B 0.016088f
C134 VDD1.t3 B 0.044992f
C135 VDD1.n118 B 0.146088f
C136 VDD1.n119 B 1.50907f
C137 VDD1.n120 B 0.011522f
C138 VDD1.n121 B 0.0122f
C139 VDD1.n122 B 0.027234f
C140 VDD1.n123 B 0.027234f
C141 VDD1.n124 B 0.0122f
C142 VDD1.n125 B 0.011522f
C143 VDD1.n126 B 0.021442f
C144 VDD1.n127 B 0.021442f
C145 VDD1.n128 B 0.011522f
C146 VDD1.n129 B 0.0122f
C147 VDD1.n130 B 0.027234f
C148 VDD1.n131 B 0.027234f
C149 VDD1.n132 B 0.0122f
C150 VDD1.n133 B 0.011522f
C151 VDD1.n134 B 0.021442f
C152 VDD1.n135 B 0.021442f
C153 VDD1.n136 B 0.011522f
C154 VDD1.n137 B 0.0122f
C155 VDD1.n138 B 0.027234f
C156 VDD1.n139 B 0.027234f
C157 VDD1.n140 B 0.0122f
C158 VDD1.n141 B 0.011522f
C159 VDD1.n142 B 0.021442f
C160 VDD1.n143 B 0.021442f
C161 VDD1.n144 B 0.011522f
C162 VDD1.n145 B 0.0122f
C163 VDD1.n146 B 0.027234f
C164 VDD1.n147 B 0.027234f
C165 VDD1.n148 B 0.0122f
C166 VDD1.n149 B 0.011522f
C167 VDD1.n150 B 0.021442f
C168 VDD1.n151 B 0.021442f
C169 VDD1.n152 B 0.011522f
C170 VDD1.n153 B 0.0122f
C171 VDD1.n154 B 0.027234f
C172 VDD1.n155 B 0.027234f
C173 VDD1.n156 B 0.0122f
C174 VDD1.n157 B 0.011522f
C175 VDD1.n158 B 0.021442f
C176 VDD1.n159 B 0.021442f
C177 VDD1.n160 B 0.011522f
C178 VDD1.n161 B 0.011522f
C179 VDD1.n162 B 0.0122f
C180 VDD1.n163 B 0.027234f
C181 VDD1.n164 B 0.027234f
C182 VDD1.n165 B 0.027234f
C183 VDD1.n166 B 0.011861f
C184 VDD1.n167 B 0.011522f
C185 VDD1.n168 B 0.021442f
C186 VDD1.n169 B 0.021442f
C187 VDD1.n170 B 0.011522f
C188 VDD1.n171 B 0.0122f
C189 VDD1.n172 B 0.027234f
C190 VDD1.n173 B 0.057935f
C191 VDD1.n174 B 0.0122f
C192 VDD1.n175 B 0.011522f
C193 VDD1.n176 B 0.051907f
C194 VDD1.n177 B 0.053333f
C195 VDD1.t1 B 0.273822f
C196 VDD1.t0 B 0.273822f
C197 VDD1.n178 B 2.48859f
C198 VDD1.n179 B 2.64789f
C199 VDD1.t2 B 0.273822f
C200 VDD1.t5 B 0.273822f
C201 VDD1.n180 B 2.48483f
C202 VDD1.n181 B 2.67434f
C203 VP.n0 B 0.029635f
C204 VP.t5 B 2.64221f
C205 VP.n1 B 0.0333f
C206 VP.n2 B 0.02248f
C207 VP.t4 B 2.64221f
C208 VP.n3 B 0.919864f
C209 VP.n4 B 0.02248f
C210 VP.n5 B 0.0333f
C211 VP.n6 B 0.029635f
C212 VP.t2 B 2.64221f
C213 VP.n7 B 0.029635f
C214 VP.t0 B 2.64221f
C215 VP.n8 B 0.0333f
C216 VP.n9 B 0.02248f
C217 VP.t3 B 2.64221f
C218 VP.n10 B 0.984996f
C219 VP.t1 B 2.84175f
C220 VP.n11 B 0.957326f
C221 VP.n12 B 0.218348f
C222 VP.n13 B 0.031397f
C223 VP.n14 B 0.041687f
C224 VP.n15 B 0.032056f
C225 VP.n16 B 0.02248f
C226 VP.n17 B 0.02248f
C227 VP.n18 B 0.02248f
C228 VP.n19 B 0.041687f
C229 VP.n20 B 0.030574f
C230 VP.n21 B 0.998018f
C231 VP.n22 B 1.32712f
C232 VP.n23 B 1.34268f
C233 VP.n24 B 0.998018f
C234 VP.n25 B 0.030574f
C235 VP.n26 B 0.041687f
C236 VP.n27 B 0.02248f
C237 VP.n28 B 0.02248f
C238 VP.n29 B 0.02248f
C239 VP.n30 B 0.032056f
C240 VP.n31 B 0.041687f
C241 VP.n32 B 0.031397f
C242 VP.n33 B 0.02248f
C243 VP.n34 B 0.02248f
C244 VP.n35 B 0.031397f
C245 VP.n36 B 0.041687f
C246 VP.n37 B 0.032056f
C247 VP.n38 B 0.02248f
C248 VP.n39 B 0.02248f
C249 VP.n40 B 0.02248f
C250 VP.n41 B 0.041687f
C251 VP.n42 B 0.030574f
C252 VP.n43 B 0.998018f
C253 VP.n44 B 0.036124f
C254 VDD2.n0 B 0.029367f
C255 VDD2.n1 B 0.021302f
C256 VDD2.n2 B 0.011447f
C257 VDD2.n3 B 0.027056f
C258 VDD2.n4 B 0.01212f
C259 VDD2.n5 B 0.021302f
C260 VDD2.n6 B 0.011783f
C261 VDD2.n7 B 0.027056f
C262 VDD2.n8 B 0.01212f
C263 VDD2.n9 B 0.021302f
C264 VDD2.n10 B 0.011447f
C265 VDD2.n11 B 0.027056f
C266 VDD2.n12 B 0.01212f
C267 VDD2.n13 B 0.021302f
C268 VDD2.n14 B 0.011447f
C269 VDD2.n15 B 0.027056f
C270 VDD2.n16 B 0.01212f
C271 VDD2.n17 B 0.021302f
C272 VDD2.n18 B 0.011447f
C273 VDD2.n19 B 0.027056f
C274 VDD2.n20 B 0.01212f
C275 VDD2.n21 B 0.021302f
C276 VDD2.n22 B 0.011447f
C277 VDD2.n23 B 0.027056f
C278 VDD2.n24 B 0.01212f
C279 VDD2.n25 B 0.021302f
C280 VDD2.n26 B 0.011447f
C281 VDD2.n27 B 0.020292f
C282 VDD2.n28 B 0.015983f
C283 VDD2.t5 B 0.044696f
C284 VDD2.n29 B 0.14513f
C285 VDD2.n30 B 1.49917f
C286 VDD2.n31 B 0.011447f
C287 VDD2.n32 B 0.01212f
C288 VDD2.n33 B 0.027056f
C289 VDD2.n34 B 0.027056f
C290 VDD2.n35 B 0.01212f
C291 VDD2.n36 B 0.011447f
C292 VDD2.n37 B 0.021302f
C293 VDD2.n38 B 0.021302f
C294 VDD2.n39 B 0.011447f
C295 VDD2.n40 B 0.01212f
C296 VDD2.n41 B 0.027056f
C297 VDD2.n42 B 0.027056f
C298 VDD2.n43 B 0.01212f
C299 VDD2.n44 B 0.011447f
C300 VDD2.n45 B 0.021302f
C301 VDD2.n46 B 0.021302f
C302 VDD2.n47 B 0.011447f
C303 VDD2.n48 B 0.01212f
C304 VDD2.n49 B 0.027056f
C305 VDD2.n50 B 0.027056f
C306 VDD2.n51 B 0.01212f
C307 VDD2.n52 B 0.011447f
C308 VDD2.n53 B 0.021302f
C309 VDD2.n54 B 0.021302f
C310 VDD2.n55 B 0.011447f
C311 VDD2.n56 B 0.01212f
C312 VDD2.n57 B 0.027056f
C313 VDD2.n58 B 0.027056f
C314 VDD2.n59 B 0.01212f
C315 VDD2.n60 B 0.011447f
C316 VDD2.n61 B 0.021302f
C317 VDD2.n62 B 0.021302f
C318 VDD2.n63 B 0.011447f
C319 VDD2.n64 B 0.01212f
C320 VDD2.n65 B 0.027056f
C321 VDD2.n66 B 0.027056f
C322 VDD2.n67 B 0.01212f
C323 VDD2.n68 B 0.011447f
C324 VDD2.n69 B 0.021302f
C325 VDD2.n70 B 0.021302f
C326 VDD2.n71 B 0.011447f
C327 VDD2.n72 B 0.011447f
C328 VDD2.n73 B 0.01212f
C329 VDD2.n74 B 0.027056f
C330 VDD2.n75 B 0.027056f
C331 VDD2.n76 B 0.027056f
C332 VDD2.n77 B 0.011783f
C333 VDD2.n78 B 0.011447f
C334 VDD2.n79 B 0.021302f
C335 VDD2.n80 B 0.021302f
C336 VDD2.n81 B 0.011447f
C337 VDD2.n82 B 0.01212f
C338 VDD2.n83 B 0.027056f
C339 VDD2.n84 B 0.057554f
C340 VDD2.n85 B 0.01212f
C341 VDD2.n86 B 0.011447f
C342 VDD2.n87 B 0.051566f
C343 VDD2.n88 B 0.052983f
C344 VDD2.t0 B 0.272027f
C345 VDD2.t3 B 0.272027f
C346 VDD2.n89 B 2.47227f
C347 VDD2.n90 B 2.52116f
C348 VDD2.n91 B 0.029367f
C349 VDD2.n92 B 0.021302f
C350 VDD2.n93 B 0.011447f
C351 VDD2.n94 B 0.027056f
C352 VDD2.n95 B 0.01212f
C353 VDD2.n96 B 0.021302f
C354 VDD2.n97 B 0.011783f
C355 VDD2.n98 B 0.027056f
C356 VDD2.n99 B 0.011447f
C357 VDD2.n100 B 0.01212f
C358 VDD2.n101 B 0.021302f
C359 VDD2.n102 B 0.011447f
C360 VDD2.n103 B 0.027056f
C361 VDD2.n104 B 0.01212f
C362 VDD2.n105 B 0.021302f
C363 VDD2.n106 B 0.011447f
C364 VDD2.n107 B 0.027056f
C365 VDD2.n108 B 0.01212f
C366 VDD2.n109 B 0.021302f
C367 VDD2.n110 B 0.011447f
C368 VDD2.n111 B 0.027056f
C369 VDD2.n112 B 0.01212f
C370 VDD2.n113 B 0.021302f
C371 VDD2.n114 B 0.011447f
C372 VDD2.n115 B 0.027056f
C373 VDD2.n116 B 0.01212f
C374 VDD2.n117 B 0.021302f
C375 VDD2.n118 B 0.011447f
C376 VDD2.n119 B 0.020292f
C377 VDD2.n120 B 0.015983f
C378 VDD2.t1 B 0.044696f
C379 VDD2.n121 B 0.14513f
C380 VDD2.n122 B 1.49917f
C381 VDD2.n123 B 0.011447f
C382 VDD2.n124 B 0.01212f
C383 VDD2.n125 B 0.027056f
C384 VDD2.n126 B 0.027056f
C385 VDD2.n127 B 0.01212f
C386 VDD2.n128 B 0.011447f
C387 VDD2.n129 B 0.021302f
C388 VDD2.n130 B 0.021302f
C389 VDD2.n131 B 0.011447f
C390 VDD2.n132 B 0.01212f
C391 VDD2.n133 B 0.027056f
C392 VDD2.n134 B 0.027056f
C393 VDD2.n135 B 0.01212f
C394 VDD2.n136 B 0.011447f
C395 VDD2.n137 B 0.021302f
C396 VDD2.n138 B 0.021302f
C397 VDD2.n139 B 0.011447f
C398 VDD2.n140 B 0.01212f
C399 VDD2.n141 B 0.027056f
C400 VDD2.n142 B 0.027056f
C401 VDD2.n143 B 0.01212f
C402 VDD2.n144 B 0.011447f
C403 VDD2.n145 B 0.021302f
C404 VDD2.n146 B 0.021302f
C405 VDD2.n147 B 0.011447f
C406 VDD2.n148 B 0.01212f
C407 VDD2.n149 B 0.027056f
C408 VDD2.n150 B 0.027056f
C409 VDD2.n151 B 0.01212f
C410 VDD2.n152 B 0.011447f
C411 VDD2.n153 B 0.021302f
C412 VDD2.n154 B 0.021302f
C413 VDD2.n155 B 0.011447f
C414 VDD2.n156 B 0.01212f
C415 VDD2.n157 B 0.027056f
C416 VDD2.n158 B 0.027056f
C417 VDD2.n159 B 0.01212f
C418 VDD2.n160 B 0.011447f
C419 VDD2.n161 B 0.021302f
C420 VDD2.n162 B 0.021302f
C421 VDD2.n163 B 0.011447f
C422 VDD2.n164 B 0.01212f
C423 VDD2.n165 B 0.027056f
C424 VDD2.n166 B 0.027056f
C425 VDD2.n167 B 0.027056f
C426 VDD2.n168 B 0.011783f
C427 VDD2.n169 B 0.011447f
C428 VDD2.n170 B 0.021302f
C429 VDD2.n171 B 0.021302f
C430 VDD2.n172 B 0.011447f
C431 VDD2.n173 B 0.01212f
C432 VDD2.n174 B 0.027056f
C433 VDD2.n175 B 0.057554f
C434 VDD2.n176 B 0.01212f
C435 VDD2.n177 B 0.011447f
C436 VDD2.n178 B 0.051566f
C437 VDD2.n179 B 0.046861f
C438 VDD2.n180 B 2.46703f
C439 VDD2.t4 B 0.272027f
C440 VDD2.t2 B 0.272027f
C441 VDD2.n181 B 2.47224f
C442 VTAIL.t9 B 0.290553f
C443 VTAIL.t10 B 0.290553f
C444 VTAIL.n0 B 2.57032f
C445 VTAIL.n1 B 0.401278f
C446 VTAIL.n2 B 0.031367f
C447 VTAIL.n3 B 0.022753f
C448 VTAIL.n4 B 0.012226f
C449 VTAIL.n5 B 0.028898f
C450 VTAIL.n6 B 0.012945f
C451 VTAIL.n7 B 0.022753f
C452 VTAIL.n8 B 0.012586f
C453 VTAIL.n9 B 0.028898f
C454 VTAIL.n10 B 0.012945f
C455 VTAIL.n11 B 0.022753f
C456 VTAIL.n12 B 0.012226f
C457 VTAIL.n13 B 0.028898f
C458 VTAIL.n14 B 0.012945f
C459 VTAIL.n15 B 0.022753f
C460 VTAIL.n16 B 0.012226f
C461 VTAIL.n17 B 0.028898f
C462 VTAIL.n18 B 0.012945f
C463 VTAIL.n19 B 0.022753f
C464 VTAIL.n20 B 0.012226f
C465 VTAIL.n21 B 0.028898f
C466 VTAIL.n22 B 0.012945f
C467 VTAIL.n23 B 0.022753f
C468 VTAIL.n24 B 0.012226f
C469 VTAIL.n25 B 0.028898f
C470 VTAIL.n26 B 0.012945f
C471 VTAIL.n27 B 0.022753f
C472 VTAIL.n28 B 0.012226f
C473 VTAIL.n29 B 0.021674f
C474 VTAIL.n30 B 0.017071f
C475 VTAIL.t1 B 0.047741f
C476 VTAIL.n31 B 0.155015f
C477 VTAIL.n32 B 1.60128f
C478 VTAIL.n33 B 0.012226f
C479 VTAIL.n34 B 0.012945f
C480 VTAIL.n35 B 0.028898f
C481 VTAIL.n36 B 0.028898f
C482 VTAIL.n37 B 0.012945f
C483 VTAIL.n38 B 0.012226f
C484 VTAIL.n39 B 0.022753f
C485 VTAIL.n40 B 0.022753f
C486 VTAIL.n41 B 0.012226f
C487 VTAIL.n42 B 0.012945f
C488 VTAIL.n43 B 0.028898f
C489 VTAIL.n44 B 0.028898f
C490 VTAIL.n45 B 0.012945f
C491 VTAIL.n46 B 0.012226f
C492 VTAIL.n47 B 0.022753f
C493 VTAIL.n48 B 0.022753f
C494 VTAIL.n49 B 0.012226f
C495 VTAIL.n50 B 0.012945f
C496 VTAIL.n51 B 0.028898f
C497 VTAIL.n52 B 0.028898f
C498 VTAIL.n53 B 0.012945f
C499 VTAIL.n54 B 0.012226f
C500 VTAIL.n55 B 0.022753f
C501 VTAIL.n56 B 0.022753f
C502 VTAIL.n57 B 0.012226f
C503 VTAIL.n58 B 0.012945f
C504 VTAIL.n59 B 0.028898f
C505 VTAIL.n60 B 0.028898f
C506 VTAIL.n61 B 0.012945f
C507 VTAIL.n62 B 0.012226f
C508 VTAIL.n63 B 0.022753f
C509 VTAIL.n64 B 0.022753f
C510 VTAIL.n65 B 0.012226f
C511 VTAIL.n66 B 0.012945f
C512 VTAIL.n67 B 0.028898f
C513 VTAIL.n68 B 0.028898f
C514 VTAIL.n69 B 0.012945f
C515 VTAIL.n70 B 0.012226f
C516 VTAIL.n71 B 0.022753f
C517 VTAIL.n72 B 0.022753f
C518 VTAIL.n73 B 0.012226f
C519 VTAIL.n74 B 0.012226f
C520 VTAIL.n75 B 0.012945f
C521 VTAIL.n76 B 0.028898f
C522 VTAIL.n77 B 0.028898f
C523 VTAIL.n78 B 0.028898f
C524 VTAIL.n79 B 0.012586f
C525 VTAIL.n80 B 0.012226f
C526 VTAIL.n81 B 0.022753f
C527 VTAIL.n82 B 0.022753f
C528 VTAIL.n83 B 0.012226f
C529 VTAIL.n84 B 0.012945f
C530 VTAIL.n85 B 0.028898f
C531 VTAIL.n86 B 0.061474f
C532 VTAIL.n87 B 0.012945f
C533 VTAIL.n88 B 0.012226f
C534 VTAIL.n89 B 0.055078f
C535 VTAIL.n90 B 0.034361f
C536 VTAIL.n91 B 0.337794f
C537 VTAIL.t2 B 0.290553f
C538 VTAIL.t3 B 0.290553f
C539 VTAIL.n92 B 2.57032f
C540 VTAIL.n93 B 2.11674f
C541 VTAIL.t6 B 0.290553f
C542 VTAIL.t7 B 0.290553f
C543 VTAIL.n94 B 2.57033f
C544 VTAIL.n95 B 2.11673f
C545 VTAIL.n96 B 0.031367f
C546 VTAIL.n97 B 0.022753f
C547 VTAIL.n98 B 0.012226f
C548 VTAIL.n99 B 0.028898f
C549 VTAIL.n100 B 0.012945f
C550 VTAIL.n101 B 0.022753f
C551 VTAIL.n102 B 0.012586f
C552 VTAIL.n103 B 0.028898f
C553 VTAIL.n104 B 0.012226f
C554 VTAIL.n105 B 0.012945f
C555 VTAIL.n106 B 0.022753f
C556 VTAIL.n107 B 0.012226f
C557 VTAIL.n108 B 0.028898f
C558 VTAIL.n109 B 0.012945f
C559 VTAIL.n110 B 0.022753f
C560 VTAIL.n111 B 0.012226f
C561 VTAIL.n112 B 0.028898f
C562 VTAIL.n113 B 0.012945f
C563 VTAIL.n114 B 0.022753f
C564 VTAIL.n115 B 0.012226f
C565 VTAIL.n116 B 0.028898f
C566 VTAIL.n117 B 0.012945f
C567 VTAIL.n118 B 0.022753f
C568 VTAIL.n119 B 0.012226f
C569 VTAIL.n120 B 0.028898f
C570 VTAIL.n121 B 0.012945f
C571 VTAIL.n122 B 0.022753f
C572 VTAIL.n123 B 0.012226f
C573 VTAIL.n124 B 0.021674f
C574 VTAIL.n125 B 0.017071f
C575 VTAIL.t8 B 0.047741f
C576 VTAIL.n126 B 0.155015f
C577 VTAIL.n127 B 1.60128f
C578 VTAIL.n128 B 0.012226f
C579 VTAIL.n129 B 0.012945f
C580 VTAIL.n130 B 0.028898f
C581 VTAIL.n131 B 0.028898f
C582 VTAIL.n132 B 0.012945f
C583 VTAIL.n133 B 0.012226f
C584 VTAIL.n134 B 0.022753f
C585 VTAIL.n135 B 0.022753f
C586 VTAIL.n136 B 0.012226f
C587 VTAIL.n137 B 0.012945f
C588 VTAIL.n138 B 0.028898f
C589 VTAIL.n139 B 0.028898f
C590 VTAIL.n140 B 0.012945f
C591 VTAIL.n141 B 0.012226f
C592 VTAIL.n142 B 0.022753f
C593 VTAIL.n143 B 0.022753f
C594 VTAIL.n144 B 0.012226f
C595 VTAIL.n145 B 0.012945f
C596 VTAIL.n146 B 0.028898f
C597 VTAIL.n147 B 0.028898f
C598 VTAIL.n148 B 0.012945f
C599 VTAIL.n149 B 0.012226f
C600 VTAIL.n150 B 0.022753f
C601 VTAIL.n151 B 0.022753f
C602 VTAIL.n152 B 0.012226f
C603 VTAIL.n153 B 0.012945f
C604 VTAIL.n154 B 0.028898f
C605 VTAIL.n155 B 0.028898f
C606 VTAIL.n156 B 0.012945f
C607 VTAIL.n157 B 0.012226f
C608 VTAIL.n158 B 0.022753f
C609 VTAIL.n159 B 0.022753f
C610 VTAIL.n160 B 0.012226f
C611 VTAIL.n161 B 0.012945f
C612 VTAIL.n162 B 0.028898f
C613 VTAIL.n163 B 0.028898f
C614 VTAIL.n164 B 0.012945f
C615 VTAIL.n165 B 0.012226f
C616 VTAIL.n166 B 0.022753f
C617 VTAIL.n167 B 0.022753f
C618 VTAIL.n168 B 0.012226f
C619 VTAIL.n169 B 0.012945f
C620 VTAIL.n170 B 0.028898f
C621 VTAIL.n171 B 0.028898f
C622 VTAIL.n172 B 0.028898f
C623 VTAIL.n173 B 0.012586f
C624 VTAIL.n174 B 0.012226f
C625 VTAIL.n175 B 0.022753f
C626 VTAIL.n176 B 0.022753f
C627 VTAIL.n177 B 0.012226f
C628 VTAIL.n178 B 0.012945f
C629 VTAIL.n179 B 0.028898f
C630 VTAIL.n180 B 0.061474f
C631 VTAIL.n181 B 0.012945f
C632 VTAIL.n182 B 0.012226f
C633 VTAIL.n183 B 0.055078f
C634 VTAIL.n184 B 0.034361f
C635 VTAIL.n185 B 0.337794f
C636 VTAIL.t5 B 0.290553f
C637 VTAIL.t0 B 0.290553f
C638 VTAIL.n186 B 2.57033f
C639 VTAIL.n187 B 0.538256f
C640 VTAIL.n188 B 0.031367f
C641 VTAIL.n189 B 0.022753f
C642 VTAIL.n190 B 0.012226f
C643 VTAIL.n191 B 0.028898f
C644 VTAIL.n192 B 0.012945f
C645 VTAIL.n193 B 0.022753f
C646 VTAIL.n194 B 0.012586f
C647 VTAIL.n195 B 0.028898f
C648 VTAIL.n196 B 0.012226f
C649 VTAIL.n197 B 0.012945f
C650 VTAIL.n198 B 0.022753f
C651 VTAIL.n199 B 0.012226f
C652 VTAIL.n200 B 0.028898f
C653 VTAIL.n201 B 0.012945f
C654 VTAIL.n202 B 0.022753f
C655 VTAIL.n203 B 0.012226f
C656 VTAIL.n204 B 0.028898f
C657 VTAIL.n205 B 0.012945f
C658 VTAIL.n206 B 0.022753f
C659 VTAIL.n207 B 0.012226f
C660 VTAIL.n208 B 0.028898f
C661 VTAIL.n209 B 0.012945f
C662 VTAIL.n210 B 0.022753f
C663 VTAIL.n211 B 0.012226f
C664 VTAIL.n212 B 0.028898f
C665 VTAIL.n213 B 0.012945f
C666 VTAIL.n214 B 0.022753f
C667 VTAIL.n215 B 0.012226f
C668 VTAIL.n216 B 0.021674f
C669 VTAIL.n217 B 0.017071f
C670 VTAIL.t4 B 0.047741f
C671 VTAIL.n218 B 0.155015f
C672 VTAIL.n219 B 1.60128f
C673 VTAIL.n220 B 0.012226f
C674 VTAIL.n221 B 0.012945f
C675 VTAIL.n222 B 0.028898f
C676 VTAIL.n223 B 0.028898f
C677 VTAIL.n224 B 0.012945f
C678 VTAIL.n225 B 0.012226f
C679 VTAIL.n226 B 0.022753f
C680 VTAIL.n227 B 0.022753f
C681 VTAIL.n228 B 0.012226f
C682 VTAIL.n229 B 0.012945f
C683 VTAIL.n230 B 0.028898f
C684 VTAIL.n231 B 0.028898f
C685 VTAIL.n232 B 0.012945f
C686 VTAIL.n233 B 0.012226f
C687 VTAIL.n234 B 0.022753f
C688 VTAIL.n235 B 0.022753f
C689 VTAIL.n236 B 0.012226f
C690 VTAIL.n237 B 0.012945f
C691 VTAIL.n238 B 0.028898f
C692 VTAIL.n239 B 0.028898f
C693 VTAIL.n240 B 0.012945f
C694 VTAIL.n241 B 0.012226f
C695 VTAIL.n242 B 0.022753f
C696 VTAIL.n243 B 0.022753f
C697 VTAIL.n244 B 0.012226f
C698 VTAIL.n245 B 0.012945f
C699 VTAIL.n246 B 0.028898f
C700 VTAIL.n247 B 0.028898f
C701 VTAIL.n248 B 0.012945f
C702 VTAIL.n249 B 0.012226f
C703 VTAIL.n250 B 0.022753f
C704 VTAIL.n251 B 0.022753f
C705 VTAIL.n252 B 0.012226f
C706 VTAIL.n253 B 0.012945f
C707 VTAIL.n254 B 0.028898f
C708 VTAIL.n255 B 0.028898f
C709 VTAIL.n256 B 0.012945f
C710 VTAIL.n257 B 0.012226f
C711 VTAIL.n258 B 0.022753f
C712 VTAIL.n259 B 0.022753f
C713 VTAIL.n260 B 0.012226f
C714 VTAIL.n261 B 0.012945f
C715 VTAIL.n262 B 0.028898f
C716 VTAIL.n263 B 0.028898f
C717 VTAIL.n264 B 0.028898f
C718 VTAIL.n265 B 0.012586f
C719 VTAIL.n266 B 0.012226f
C720 VTAIL.n267 B 0.022753f
C721 VTAIL.n268 B 0.022753f
C722 VTAIL.n269 B 0.012226f
C723 VTAIL.n270 B 0.012945f
C724 VTAIL.n271 B 0.028898f
C725 VTAIL.n272 B 0.061474f
C726 VTAIL.n273 B 0.012945f
C727 VTAIL.n274 B 0.012226f
C728 VTAIL.n275 B 0.055078f
C729 VTAIL.n276 B 0.034361f
C730 VTAIL.n277 B 1.72793f
C731 VTAIL.n278 B 0.031367f
C732 VTAIL.n279 B 0.022753f
C733 VTAIL.n280 B 0.012226f
C734 VTAIL.n281 B 0.028898f
C735 VTAIL.n282 B 0.012945f
C736 VTAIL.n283 B 0.022753f
C737 VTAIL.n284 B 0.012586f
C738 VTAIL.n285 B 0.028898f
C739 VTAIL.n286 B 0.012945f
C740 VTAIL.n287 B 0.022753f
C741 VTAIL.n288 B 0.012226f
C742 VTAIL.n289 B 0.028898f
C743 VTAIL.n290 B 0.012945f
C744 VTAIL.n291 B 0.022753f
C745 VTAIL.n292 B 0.012226f
C746 VTAIL.n293 B 0.028898f
C747 VTAIL.n294 B 0.012945f
C748 VTAIL.n295 B 0.022753f
C749 VTAIL.n296 B 0.012226f
C750 VTAIL.n297 B 0.028898f
C751 VTAIL.n298 B 0.012945f
C752 VTAIL.n299 B 0.022753f
C753 VTAIL.n300 B 0.012226f
C754 VTAIL.n301 B 0.028898f
C755 VTAIL.n302 B 0.012945f
C756 VTAIL.n303 B 0.022753f
C757 VTAIL.n304 B 0.012226f
C758 VTAIL.n305 B 0.021674f
C759 VTAIL.n306 B 0.017071f
C760 VTAIL.t11 B 0.047741f
C761 VTAIL.n307 B 0.155015f
C762 VTAIL.n308 B 1.60128f
C763 VTAIL.n309 B 0.012226f
C764 VTAIL.n310 B 0.012945f
C765 VTAIL.n311 B 0.028898f
C766 VTAIL.n312 B 0.028898f
C767 VTAIL.n313 B 0.012945f
C768 VTAIL.n314 B 0.012226f
C769 VTAIL.n315 B 0.022753f
C770 VTAIL.n316 B 0.022753f
C771 VTAIL.n317 B 0.012226f
C772 VTAIL.n318 B 0.012945f
C773 VTAIL.n319 B 0.028898f
C774 VTAIL.n320 B 0.028898f
C775 VTAIL.n321 B 0.012945f
C776 VTAIL.n322 B 0.012226f
C777 VTAIL.n323 B 0.022753f
C778 VTAIL.n324 B 0.022753f
C779 VTAIL.n325 B 0.012226f
C780 VTAIL.n326 B 0.012945f
C781 VTAIL.n327 B 0.028898f
C782 VTAIL.n328 B 0.028898f
C783 VTAIL.n329 B 0.012945f
C784 VTAIL.n330 B 0.012226f
C785 VTAIL.n331 B 0.022753f
C786 VTAIL.n332 B 0.022753f
C787 VTAIL.n333 B 0.012226f
C788 VTAIL.n334 B 0.012945f
C789 VTAIL.n335 B 0.028898f
C790 VTAIL.n336 B 0.028898f
C791 VTAIL.n337 B 0.012945f
C792 VTAIL.n338 B 0.012226f
C793 VTAIL.n339 B 0.022753f
C794 VTAIL.n340 B 0.022753f
C795 VTAIL.n341 B 0.012226f
C796 VTAIL.n342 B 0.012945f
C797 VTAIL.n343 B 0.028898f
C798 VTAIL.n344 B 0.028898f
C799 VTAIL.n345 B 0.012945f
C800 VTAIL.n346 B 0.012226f
C801 VTAIL.n347 B 0.022753f
C802 VTAIL.n348 B 0.022753f
C803 VTAIL.n349 B 0.012226f
C804 VTAIL.n350 B 0.012226f
C805 VTAIL.n351 B 0.012945f
C806 VTAIL.n352 B 0.028898f
C807 VTAIL.n353 B 0.028898f
C808 VTAIL.n354 B 0.028898f
C809 VTAIL.n355 B 0.012586f
C810 VTAIL.n356 B 0.012226f
C811 VTAIL.n357 B 0.022753f
C812 VTAIL.n358 B 0.022753f
C813 VTAIL.n359 B 0.012226f
C814 VTAIL.n360 B 0.012945f
C815 VTAIL.n361 B 0.028898f
C816 VTAIL.n362 B 0.061474f
C817 VTAIL.n363 B 0.012945f
C818 VTAIL.n364 B 0.012226f
C819 VTAIL.n365 B 0.055078f
C820 VTAIL.n366 B 0.034361f
C821 VTAIL.n367 B 1.67657f
C822 VN.n0 B 0.029257f
C823 VN.t2 B 2.60842f
C824 VN.n1 B 0.032874f
C825 VN.n2 B 0.022192f
C826 VN.t5 B 2.60842f
C827 VN.n3 B 0.972401f
C828 VN.t0 B 2.80541f
C829 VN.n4 B 0.945084f
C830 VN.n5 B 0.215555f
C831 VN.n6 B 0.030995f
C832 VN.n7 B 0.041153f
C833 VN.n8 B 0.031646f
C834 VN.n9 B 0.022192f
C835 VN.n10 B 0.022192f
C836 VN.n11 B 0.022192f
C837 VN.n12 B 0.041153f
C838 VN.n13 B 0.030183f
C839 VN.n14 B 0.985256f
C840 VN.n15 B 0.035662f
C841 VN.n16 B 0.029257f
C842 VN.t4 B 2.60842f
C843 VN.n17 B 0.032874f
C844 VN.n18 B 0.022192f
C845 VN.t1 B 2.60842f
C846 VN.n19 B 0.972401f
C847 VN.t3 B 2.80541f
C848 VN.n20 B 0.945084f
C849 VN.n21 B 0.215555f
C850 VN.n22 B 0.030995f
C851 VN.n23 B 0.041153f
C852 VN.n24 B 0.031646f
C853 VN.n25 B 0.022192f
C854 VN.n26 B 0.022192f
C855 VN.n27 B 0.022192f
C856 VN.n28 B 0.041153f
C857 VN.n29 B 0.030183f
C858 VN.n30 B 0.985256f
C859 VN.n31 B 1.32199f
.ends

