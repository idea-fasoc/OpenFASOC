* NGSPICE file created from diff_pair_sample_1745.ext - technology: sky130A

.subckt diff_pair_sample_1745 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t2 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0.6903 ps=4.32 w=1.77 l=3.53
X1 VDD2.t1 VN.t0 VTAIL.t0 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0.6903 ps=4.32 w=1.77 l=3.53
X2 B.t11 B.t9 B.t10 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=3.53
X3 B.t8 B.t6 B.t7 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=3.53
X4 B.t5 B.t3 B.t4 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=3.53
X5 B.t2 B.t0 B.t1 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0 ps=0 w=1.77 l=3.53
X6 VDD2.t0 VN.t1 VTAIL.t1 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0.6903 ps=4.32 w=1.77 l=3.53
X7 VDD1.t0 VP.t1 VTAIL.t3 w_n2514_n1322# sky130_fd_pr__pfet_01v8 ad=0.6903 pd=4.32 as=0.6903 ps=4.32 w=1.77 l=3.53
R0 VP.n0 VP.t0 90.2449
R1 VP.n0 VP.t1 50.8724
R2 VP VP.n0 0.52637
R3 VTAIL.n26 VTAIL.n24 756.745
R4 VTAIL.n2 VTAIL.n0 756.745
R5 VTAIL.n18 VTAIL.n16 756.745
R6 VTAIL.n10 VTAIL.n8 756.745
R7 VTAIL.n27 VTAIL.n26 585
R8 VTAIL.n3 VTAIL.n2 585
R9 VTAIL.n19 VTAIL.n18 585
R10 VTAIL.n11 VTAIL.n10 585
R11 VTAIL.t1 VTAIL.n25 415.613
R12 VTAIL.t3 VTAIL.n1 415.613
R13 VTAIL.t2 VTAIL.n17 415.613
R14 VTAIL.t0 VTAIL.n9 415.613
R15 VTAIL.n26 VTAIL.t1 85.8723
R16 VTAIL.n2 VTAIL.t3 85.8723
R17 VTAIL.n18 VTAIL.t2 85.8723
R18 VTAIL.n10 VTAIL.t0 85.8723
R19 VTAIL.n31 VTAIL.n30 33.9308
R20 VTAIL.n7 VTAIL.n6 33.9308
R21 VTAIL.n23 VTAIL.n22 33.9308
R22 VTAIL.n15 VTAIL.n14 33.9308
R23 VTAIL.n15 VTAIL.n7 20.5479
R24 VTAIL.n31 VTAIL.n23 17.2203
R25 VTAIL.n27 VTAIL.n25 14.9339
R26 VTAIL.n3 VTAIL.n1 14.9339
R27 VTAIL.n19 VTAIL.n17 14.9339
R28 VTAIL.n11 VTAIL.n9 14.9339
R29 VTAIL.n28 VTAIL.n24 12.8005
R30 VTAIL.n4 VTAIL.n0 12.8005
R31 VTAIL.n20 VTAIL.n16 12.8005
R32 VTAIL.n12 VTAIL.n8 12.8005
R33 VTAIL.n30 VTAIL.n29 9.45567
R34 VTAIL.n6 VTAIL.n5 9.45567
R35 VTAIL.n22 VTAIL.n21 9.45567
R36 VTAIL.n14 VTAIL.n13 9.45567
R37 VTAIL.n29 VTAIL.n28 9.3005
R38 VTAIL.n5 VTAIL.n4 9.3005
R39 VTAIL.n21 VTAIL.n20 9.3005
R40 VTAIL.n13 VTAIL.n12 9.3005
R41 VTAIL.n29 VTAIL.n25 5.44463
R42 VTAIL.n5 VTAIL.n1 5.44463
R43 VTAIL.n21 VTAIL.n17 5.44463
R44 VTAIL.n13 VTAIL.n9 5.44463
R45 VTAIL.n23 VTAIL.n15 2.13412
R46 VTAIL VTAIL.n7 1.36041
R47 VTAIL.n30 VTAIL.n24 1.16414
R48 VTAIL.n6 VTAIL.n0 1.16414
R49 VTAIL.n22 VTAIL.n16 1.16414
R50 VTAIL.n14 VTAIL.n8 1.16414
R51 VTAIL VTAIL.n31 0.774207
R52 VTAIL.n28 VTAIL.n27 0.388379
R53 VTAIL.n4 VTAIL.n3 0.388379
R54 VTAIL.n20 VTAIL.n19 0.388379
R55 VTAIL.n12 VTAIL.n11 0.388379
R56 VDD1.n2 VDD1.n0 756.745
R57 VDD1.n9 VDD1.n7 756.745
R58 VDD1.n3 VDD1.n2 585
R59 VDD1.n10 VDD1.n9 585
R60 VDD1.t0 VDD1.n8 415.613
R61 VDD1.t1 VDD1.n1 415.613
R62 VDD1.n2 VDD1.t1 85.8723
R63 VDD1.n9 VDD1.t0 85.8723
R64 VDD1 VDD1.n13 83.8068
R65 VDD1 VDD1.n6 51.4997
R66 VDD1.n3 VDD1.n1 14.9339
R67 VDD1.n10 VDD1.n8 14.9339
R68 VDD1.n4 VDD1.n0 12.8005
R69 VDD1.n11 VDD1.n7 12.8005
R70 VDD1.n6 VDD1.n5 9.45567
R71 VDD1.n13 VDD1.n12 9.45567
R72 VDD1.n5 VDD1.n4 9.3005
R73 VDD1.n12 VDD1.n11 9.3005
R74 VDD1.n5 VDD1.n1 5.44463
R75 VDD1.n12 VDD1.n8 5.44463
R76 VDD1.n6 VDD1.n0 1.16414
R77 VDD1.n13 VDD1.n7 1.16414
R78 VDD1.n4 VDD1.n3 0.388379
R79 VDD1.n11 VDD1.n10 0.388379
R80 VN VN.t0 90.152
R81 VN VN.t1 51.3983
R82 VDD2.n9 VDD2.n7 756.745
R83 VDD2.n2 VDD2.n0 756.745
R84 VDD2.n10 VDD2.n9 585
R85 VDD2.n3 VDD2.n2 585
R86 VDD2.t0 VDD2.n1 415.613
R87 VDD2.t1 VDD2.n8 415.613
R88 VDD2.n9 VDD2.t1 85.8723
R89 VDD2.n2 VDD2.t0 85.8723
R90 VDD2.n14 VDD2.n6 82.4501
R91 VDD2.n14 VDD2.n13 50.6096
R92 VDD2.n10 VDD2.n8 14.9339
R93 VDD2.n3 VDD2.n1 14.9339
R94 VDD2.n11 VDD2.n7 12.8005
R95 VDD2.n4 VDD2.n0 12.8005
R96 VDD2.n13 VDD2.n12 9.45567
R97 VDD2.n6 VDD2.n5 9.45567
R98 VDD2.n12 VDD2.n11 9.3005
R99 VDD2.n5 VDD2.n4 9.3005
R100 VDD2.n12 VDD2.n8 5.44463
R101 VDD2.n5 VDD2.n1 5.44463
R102 VDD2.n13 VDD2.n7 1.16414
R103 VDD2.n6 VDD2.n0 1.16414
R104 VDD2 VDD2.n14 0.890586
R105 VDD2.n11 VDD2.n10 0.388379
R106 VDD2.n4 VDD2.n3 0.388379
R107 B.n297 B.n38 585
R108 B.n299 B.n298 585
R109 B.n300 B.n37 585
R110 B.n302 B.n301 585
R111 B.n303 B.n36 585
R112 B.n305 B.n304 585
R113 B.n306 B.n35 585
R114 B.n308 B.n307 585
R115 B.n309 B.n34 585
R116 B.n311 B.n310 585
R117 B.n312 B.n33 585
R118 B.n314 B.n313 585
R119 B.n316 B.n315 585
R120 B.n317 B.n29 585
R121 B.n319 B.n318 585
R122 B.n320 B.n28 585
R123 B.n322 B.n321 585
R124 B.n323 B.n27 585
R125 B.n325 B.n324 585
R126 B.n326 B.n26 585
R127 B.n328 B.n327 585
R128 B.n330 B.n23 585
R129 B.n332 B.n331 585
R130 B.n333 B.n22 585
R131 B.n335 B.n334 585
R132 B.n336 B.n21 585
R133 B.n338 B.n337 585
R134 B.n339 B.n20 585
R135 B.n341 B.n340 585
R136 B.n342 B.n19 585
R137 B.n344 B.n343 585
R138 B.n345 B.n18 585
R139 B.n347 B.n346 585
R140 B.n296 B.n295 585
R141 B.n294 B.n39 585
R142 B.n293 B.n292 585
R143 B.n291 B.n40 585
R144 B.n290 B.n289 585
R145 B.n288 B.n41 585
R146 B.n287 B.n286 585
R147 B.n285 B.n42 585
R148 B.n284 B.n283 585
R149 B.n282 B.n43 585
R150 B.n281 B.n280 585
R151 B.n279 B.n44 585
R152 B.n278 B.n277 585
R153 B.n276 B.n45 585
R154 B.n275 B.n274 585
R155 B.n273 B.n46 585
R156 B.n272 B.n271 585
R157 B.n270 B.n47 585
R158 B.n269 B.n268 585
R159 B.n267 B.n48 585
R160 B.n266 B.n265 585
R161 B.n264 B.n49 585
R162 B.n263 B.n262 585
R163 B.n261 B.n50 585
R164 B.n260 B.n259 585
R165 B.n258 B.n51 585
R166 B.n257 B.n256 585
R167 B.n255 B.n52 585
R168 B.n254 B.n253 585
R169 B.n252 B.n53 585
R170 B.n251 B.n250 585
R171 B.n249 B.n54 585
R172 B.n248 B.n247 585
R173 B.n246 B.n55 585
R174 B.n245 B.n244 585
R175 B.n243 B.n56 585
R176 B.n242 B.n241 585
R177 B.n240 B.n57 585
R178 B.n239 B.n238 585
R179 B.n237 B.n58 585
R180 B.n236 B.n235 585
R181 B.n234 B.n59 585
R182 B.n233 B.n232 585
R183 B.n231 B.n60 585
R184 B.n230 B.n229 585
R185 B.n228 B.n61 585
R186 B.n227 B.n226 585
R187 B.n225 B.n62 585
R188 B.n224 B.n223 585
R189 B.n222 B.n63 585
R190 B.n221 B.n220 585
R191 B.n219 B.n64 585
R192 B.n218 B.n217 585
R193 B.n216 B.n65 585
R194 B.n215 B.n214 585
R195 B.n213 B.n66 585
R196 B.n212 B.n211 585
R197 B.n210 B.n67 585
R198 B.n209 B.n208 585
R199 B.n207 B.n68 585
R200 B.n206 B.n205 585
R201 B.n204 B.n69 585
R202 B.n203 B.n202 585
R203 B.n152 B.n151 585
R204 B.n153 B.n90 585
R205 B.n155 B.n154 585
R206 B.n156 B.n89 585
R207 B.n158 B.n157 585
R208 B.n159 B.n88 585
R209 B.n161 B.n160 585
R210 B.n162 B.n87 585
R211 B.n164 B.n163 585
R212 B.n165 B.n86 585
R213 B.n167 B.n166 585
R214 B.n168 B.n83 585
R215 B.n171 B.n170 585
R216 B.n172 B.n82 585
R217 B.n174 B.n173 585
R218 B.n175 B.n81 585
R219 B.n177 B.n176 585
R220 B.n178 B.n80 585
R221 B.n180 B.n179 585
R222 B.n181 B.n79 585
R223 B.n183 B.n182 585
R224 B.n185 B.n184 585
R225 B.n186 B.n75 585
R226 B.n188 B.n187 585
R227 B.n189 B.n74 585
R228 B.n191 B.n190 585
R229 B.n192 B.n73 585
R230 B.n194 B.n193 585
R231 B.n195 B.n72 585
R232 B.n197 B.n196 585
R233 B.n198 B.n71 585
R234 B.n200 B.n199 585
R235 B.n201 B.n70 585
R236 B.n150 B.n91 585
R237 B.n149 B.n148 585
R238 B.n147 B.n92 585
R239 B.n146 B.n145 585
R240 B.n144 B.n93 585
R241 B.n143 B.n142 585
R242 B.n141 B.n94 585
R243 B.n140 B.n139 585
R244 B.n138 B.n95 585
R245 B.n137 B.n136 585
R246 B.n135 B.n96 585
R247 B.n134 B.n133 585
R248 B.n132 B.n97 585
R249 B.n131 B.n130 585
R250 B.n129 B.n98 585
R251 B.n128 B.n127 585
R252 B.n126 B.n99 585
R253 B.n125 B.n124 585
R254 B.n123 B.n100 585
R255 B.n122 B.n121 585
R256 B.n120 B.n101 585
R257 B.n119 B.n118 585
R258 B.n117 B.n102 585
R259 B.n116 B.n115 585
R260 B.n114 B.n103 585
R261 B.n113 B.n112 585
R262 B.n111 B.n104 585
R263 B.n110 B.n109 585
R264 B.n108 B.n105 585
R265 B.n107 B.n106 585
R266 B.n2 B.n0 585
R267 B.n393 B.n1 585
R268 B.n392 B.n391 585
R269 B.n390 B.n3 585
R270 B.n389 B.n388 585
R271 B.n387 B.n4 585
R272 B.n386 B.n385 585
R273 B.n384 B.n5 585
R274 B.n383 B.n382 585
R275 B.n381 B.n6 585
R276 B.n380 B.n379 585
R277 B.n378 B.n7 585
R278 B.n377 B.n376 585
R279 B.n375 B.n8 585
R280 B.n374 B.n373 585
R281 B.n372 B.n9 585
R282 B.n371 B.n370 585
R283 B.n369 B.n10 585
R284 B.n368 B.n367 585
R285 B.n366 B.n11 585
R286 B.n365 B.n364 585
R287 B.n363 B.n12 585
R288 B.n362 B.n361 585
R289 B.n360 B.n13 585
R290 B.n359 B.n358 585
R291 B.n357 B.n14 585
R292 B.n356 B.n355 585
R293 B.n354 B.n15 585
R294 B.n353 B.n352 585
R295 B.n351 B.n16 585
R296 B.n350 B.n349 585
R297 B.n348 B.n17 585
R298 B.n395 B.n394 585
R299 B.n152 B.n91 439.647
R300 B.n346 B.n17 439.647
R301 B.n202 B.n201 439.647
R302 B.n297 B.n296 439.647
R303 B.n76 B.t5 318.738
R304 B.n30 B.t7 318.738
R305 B.n84 B.t2 318.738
R306 B.n24 B.t10 318.738
R307 B.n77 B.t4 243.876
R308 B.n31 B.t8 243.876
R309 B.n85 B.t1 243.876
R310 B.n25 B.t11 243.876
R311 B.n76 B.t3 209.543
R312 B.n84 B.t0 209.543
R313 B.n24 B.t9 209.543
R314 B.n30 B.t6 209.543
R315 B.n148 B.n91 163.367
R316 B.n148 B.n147 163.367
R317 B.n147 B.n146 163.367
R318 B.n146 B.n93 163.367
R319 B.n142 B.n93 163.367
R320 B.n142 B.n141 163.367
R321 B.n141 B.n140 163.367
R322 B.n140 B.n95 163.367
R323 B.n136 B.n95 163.367
R324 B.n136 B.n135 163.367
R325 B.n135 B.n134 163.367
R326 B.n134 B.n97 163.367
R327 B.n130 B.n97 163.367
R328 B.n130 B.n129 163.367
R329 B.n129 B.n128 163.367
R330 B.n128 B.n99 163.367
R331 B.n124 B.n99 163.367
R332 B.n124 B.n123 163.367
R333 B.n123 B.n122 163.367
R334 B.n122 B.n101 163.367
R335 B.n118 B.n101 163.367
R336 B.n118 B.n117 163.367
R337 B.n117 B.n116 163.367
R338 B.n116 B.n103 163.367
R339 B.n112 B.n103 163.367
R340 B.n112 B.n111 163.367
R341 B.n111 B.n110 163.367
R342 B.n110 B.n105 163.367
R343 B.n106 B.n105 163.367
R344 B.n106 B.n2 163.367
R345 B.n394 B.n2 163.367
R346 B.n394 B.n393 163.367
R347 B.n393 B.n392 163.367
R348 B.n392 B.n3 163.367
R349 B.n388 B.n3 163.367
R350 B.n388 B.n387 163.367
R351 B.n387 B.n386 163.367
R352 B.n386 B.n5 163.367
R353 B.n382 B.n5 163.367
R354 B.n382 B.n381 163.367
R355 B.n381 B.n380 163.367
R356 B.n380 B.n7 163.367
R357 B.n376 B.n7 163.367
R358 B.n376 B.n375 163.367
R359 B.n375 B.n374 163.367
R360 B.n374 B.n9 163.367
R361 B.n370 B.n9 163.367
R362 B.n370 B.n369 163.367
R363 B.n369 B.n368 163.367
R364 B.n368 B.n11 163.367
R365 B.n364 B.n11 163.367
R366 B.n364 B.n363 163.367
R367 B.n363 B.n362 163.367
R368 B.n362 B.n13 163.367
R369 B.n358 B.n13 163.367
R370 B.n358 B.n357 163.367
R371 B.n357 B.n356 163.367
R372 B.n356 B.n15 163.367
R373 B.n352 B.n15 163.367
R374 B.n352 B.n351 163.367
R375 B.n351 B.n350 163.367
R376 B.n350 B.n17 163.367
R377 B.n153 B.n152 163.367
R378 B.n154 B.n153 163.367
R379 B.n154 B.n89 163.367
R380 B.n158 B.n89 163.367
R381 B.n159 B.n158 163.367
R382 B.n160 B.n159 163.367
R383 B.n160 B.n87 163.367
R384 B.n164 B.n87 163.367
R385 B.n165 B.n164 163.367
R386 B.n166 B.n165 163.367
R387 B.n166 B.n83 163.367
R388 B.n171 B.n83 163.367
R389 B.n172 B.n171 163.367
R390 B.n173 B.n172 163.367
R391 B.n173 B.n81 163.367
R392 B.n177 B.n81 163.367
R393 B.n178 B.n177 163.367
R394 B.n179 B.n178 163.367
R395 B.n179 B.n79 163.367
R396 B.n183 B.n79 163.367
R397 B.n184 B.n183 163.367
R398 B.n184 B.n75 163.367
R399 B.n188 B.n75 163.367
R400 B.n189 B.n188 163.367
R401 B.n190 B.n189 163.367
R402 B.n190 B.n73 163.367
R403 B.n194 B.n73 163.367
R404 B.n195 B.n194 163.367
R405 B.n196 B.n195 163.367
R406 B.n196 B.n71 163.367
R407 B.n200 B.n71 163.367
R408 B.n201 B.n200 163.367
R409 B.n202 B.n69 163.367
R410 B.n206 B.n69 163.367
R411 B.n207 B.n206 163.367
R412 B.n208 B.n207 163.367
R413 B.n208 B.n67 163.367
R414 B.n212 B.n67 163.367
R415 B.n213 B.n212 163.367
R416 B.n214 B.n213 163.367
R417 B.n214 B.n65 163.367
R418 B.n218 B.n65 163.367
R419 B.n219 B.n218 163.367
R420 B.n220 B.n219 163.367
R421 B.n220 B.n63 163.367
R422 B.n224 B.n63 163.367
R423 B.n225 B.n224 163.367
R424 B.n226 B.n225 163.367
R425 B.n226 B.n61 163.367
R426 B.n230 B.n61 163.367
R427 B.n231 B.n230 163.367
R428 B.n232 B.n231 163.367
R429 B.n232 B.n59 163.367
R430 B.n236 B.n59 163.367
R431 B.n237 B.n236 163.367
R432 B.n238 B.n237 163.367
R433 B.n238 B.n57 163.367
R434 B.n242 B.n57 163.367
R435 B.n243 B.n242 163.367
R436 B.n244 B.n243 163.367
R437 B.n244 B.n55 163.367
R438 B.n248 B.n55 163.367
R439 B.n249 B.n248 163.367
R440 B.n250 B.n249 163.367
R441 B.n250 B.n53 163.367
R442 B.n254 B.n53 163.367
R443 B.n255 B.n254 163.367
R444 B.n256 B.n255 163.367
R445 B.n256 B.n51 163.367
R446 B.n260 B.n51 163.367
R447 B.n261 B.n260 163.367
R448 B.n262 B.n261 163.367
R449 B.n262 B.n49 163.367
R450 B.n266 B.n49 163.367
R451 B.n267 B.n266 163.367
R452 B.n268 B.n267 163.367
R453 B.n268 B.n47 163.367
R454 B.n272 B.n47 163.367
R455 B.n273 B.n272 163.367
R456 B.n274 B.n273 163.367
R457 B.n274 B.n45 163.367
R458 B.n278 B.n45 163.367
R459 B.n279 B.n278 163.367
R460 B.n280 B.n279 163.367
R461 B.n280 B.n43 163.367
R462 B.n284 B.n43 163.367
R463 B.n285 B.n284 163.367
R464 B.n286 B.n285 163.367
R465 B.n286 B.n41 163.367
R466 B.n290 B.n41 163.367
R467 B.n291 B.n290 163.367
R468 B.n292 B.n291 163.367
R469 B.n292 B.n39 163.367
R470 B.n296 B.n39 163.367
R471 B.n346 B.n345 163.367
R472 B.n345 B.n344 163.367
R473 B.n344 B.n19 163.367
R474 B.n340 B.n19 163.367
R475 B.n340 B.n339 163.367
R476 B.n339 B.n338 163.367
R477 B.n338 B.n21 163.367
R478 B.n334 B.n21 163.367
R479 B.n334 B.n333 163.367
R480 B.n333 B.n332 163.367
R481 B.n332 B.n23 163.367
R482 B.n327 B.n23 163.367
R483 B.n327 B.n326 163.367
R484 B.n326 B.n325 163.367
R485 B.n325 B.n27 163.367
R486 B.n321 B.n27 163.367
R487 B.n321 B.n320 163.367
R488 B.n320 B.n319 163.367
R489 B.n319 B.n29 163.367
R490 B.n315 B.n29 163.367
R491 B.n315 B.n314 163.367
R492 B.n314 B.n33 163.367
R493 B.n310 B.n33 163.367
R494 B.n310 B.n309 163.367
R495 B.n309 B.n308 163.367
R496 B.n308 B.n35 163.367
R497 B.n304 B.n35 163.367
R498 B.n304 B.n303 163.367
R499 B.n303 B.n302 163.367
R500 B.n302 B.n37 163.367
R501 B.n298 B.n37 163.367
R502 B.n298 B.n297 163.367
R503 B.n77 B.n76 74.8611
R504 B.n85 B.n84 74.8611
R505 B.n25 B.n24 74.8611
R506 B.n31 B.n30 74.8611
R507 B.n78 B.n77 59.5399
R508 B.n169 B.n85 59.5399
R509 B.n329 B.n25 59.5399
R510 B.n32 B.n31 59.5399
R511 B.n348 B.n347 28.5664
R512 B.n203 B.n70 28.5664
R513 B.n151 B.n150 28.5664
R514 B.n295 B.n38 28.5664
R515 B B.n395 18.0485
R516 B.n347 B.n18 10.6151
R517 B.n343 B.n18 10.6151
R518 B.n343 B.n342 10.6151
R519 B.n342 B.n341 10.6151
R520 B.n341 B.n20 10.6151
R521 B.n337 B.n20 10.6151
R522 B.n337 B.n336 10.6151
R523 B.n336 B.n335 10.6151
R524 B.n335 B.n22 10.6151
R525 B.n331 B.n22 10.6151
R526 B.n331 B.n330 10.6151
R527 B.n328 B.n26 10.6151
R528 B.n324 B.n26 10.6151
R529 B.n324 B.n323 10.6151
R530 B.n323 B.n322 10.6151
R531 B.n322 B.n28 10.6151
R532 B.n318 B.n28 10.6151
R533 B.n318 B.n317 10.6151
R534 B.n317 B.n316 10.6151
R535 B.n313 B.n312 10.6151
R536 B.n312 B.n311 10.6151
R537 B.n311 B.n34 10.6151
R538 B.n307 B.n34 10.6151
R539 B.n307 B.n306 10.6151
R540 B.n306 B.n305 10.6151
R541 B.n305 B.n36 10.6151
R542 B.n301 B.n36 10.6151
R543 B.n301 B.n300 10.6151
R544 B.n300 B.n299 10.6151
R545 B.n299 B.n38 10.6151
R546 B.n204 B.n203 10.6151
R547 B.n205 B.n204 10.6151
R548 B.n205 B.n68 10.6151
R549 B.n209 B.n68 10.6151
R550 B.n210 B.n209 10.6151
R551 B.n211 B.n210 10.6151
R552 B.n211 B.n66 10.6151
R553 B.n215 B.n66 10.6151
R554 B.n216 B.n215 10.6151
R555 B.n217 B.n216 10.6151
R556 B.n217 B.n64 10.6151
R557 B.n221 B.n64 10.6151
R558 B.n222 B.n221 10.6151
R559 B.n223 B.n222 10.6151
R560 B.n223 B.n62 10.6151
R561 B.n227 B.n62 10.6151
R562 B.n228 B.n227 10.6151
R563 B.n229 B.n228 10.6151
R564 B.n229 B.n60 10.6151
R565 B.n233 B.n60 10.6151
R566 B.n234 B.n233 10.6151
R567 B.n235 B.n234 10.6151
R568 B.n235 B.n58 10.6151
R569 B.n239 B.n58 10.6151
R570 B.n240 B.n239 10.6151
R571 B.n241 B.n240 10.6151
R572 B.n241 B.n56 10.6151
R573 B.n245 B.n56 10.6151
R574 B.n246 B.n245 10.6151
R575 B.n247 B.n246 10.6151
R576 B.n247 B.n54 10.6151
R577 B.n251 B.n54 10.6151
R578 B.n252 B.n251 10.6151
R579 B.n253 B.n252 10.6151
R580 B.n253 B.n52 10.6151
R581 B.n257 B.n52 10.6151
R582 B.n258 B.n257 10.6151
R583 B.n259 B.n258 10.6151
R584 B.n259 B.n50 10.6151
R585 B.n263 B.n50 10.6151
R586 B.n264 B.n263 10.6151
R587 B.n265 B.n264 10.6151
R588 B.n265 B.n48 10.6151
R589 B.n269 B.n48 10.6151
R590 B.n270 B.n269 10.6151
R591 B.n271 B.n270 10.6151
R592 B.n271 B.n46 10.6151
R593 B.n275 B.n46 10.6151
R594 B.n276 B.n275 10.6151
R595 B.n277 B.n276 10.6151
R596 B.n277 B.n44 10.6151
R597 B.n281 B.n44 10.6151
R598 B.n282 B.n281 10.6151
R599 B.n283 B.n282 10.6151
R600 B.n283 B.n42 10.6151
R601 B.n287 B.n42 10.6151
R602 B.n288 B.n287 10.6151
R603 B.n289 B.n288 10.6151
R604 B.n289 B.n40 10.6151
R605 B.n293 B.n40 10.6151
R606 B.n294 B.n293 10.6151
R607 B.n295 B.n294 10.6151
R608 B.n151 B.n90 10.6151
R609 B.n155 B.n90 10.6151
R610 B.n156 B.n155 10.6151
R611 B.n157 B.n156 10.6151
R612 B.n157 B.n88 10.6151
R613 B.n161 B.n88 10.6151
R614 B.n162 B.n161 10.6151
R615 B.n163 B.n162 10.6151
R616 B.n163 B.n86 10.6151
R617 B.n167 B.n86 10.6151
R618 B.n168 B.n167 10.6151
R619 B.n170 B.n82 10.6151
R620 B.n174 B.n82 10.6151
R621 B.n175 B.n174 10.6151
R622 B.n176 B.n175 10.6151
R623 B.n176 B.n80 10.6151
R624 B.n180 B.n80 10.6151
R625 B.n181 B.n180 10.6151
R626 B.n182 B.n181 10.6151
R627 B.n186 B.n185 10.6151
R628 B.n187 B.n186 10.6151
R629 B.n187 B.n74 10.6151
R630 B.n191 B.n74 10.6151
R631 B.n192 B.n191 10.6151
R632 B.n193 B.n192 10.6151
R633 B.n193 B.n72 10.6151
R634 B.n197 B.n72 10.6151
R635 B.n198 B.n197 10.6151
R636 B.n199 B.n198 10.6151
R637 B.n199 B.n70 10.6151
R638 B.n150 B.n149 10.6151
R639 B.n149 B.n92 10.6151
R640 B.n145 B.n92 10.6151
R641 B.n145 B.n144 10.6151
R642 B.n144 B.n143 10.6151
R643 B.n143 B.n94 10.6151
R644 B.n139 B.n94 10.6151
R645 B.n139 B.n138 10.6151
R646 B.n138 B.n137 10.6151
R647 B.n137 B.n96 10.6151
R648 B.n133 B.n96 10.6151
R649 B.n133 B.n132 10.6151
R650 B.n132 B.n131 10.6151
R651 B.n131 B.n98 10.6151
R652 B.n127 B.n98 10.6151
R653 B.n127 B.n126 10.6151
R654 B.n126 B.n125 10.6151
R655 B.n125 B.n100 10.6151
R656 B.n121 B.n100 10.6151
R657 B.n121 B.n120 10.6151
R658 B.n120 B.n119 10.6151
R659 B.n119 B.n102 10.6151
R660 B.n115 B.n102 10.6151
R661 B.n115 B.n114 10.6151
R662 B.n114 B.n113 10.6151
R663 B.n113 B.n104 10.6151
R664 B.n109 B.n104 10.6151
R665 B.n109 B.n108 10.6151
R666 B.n108 B.n107 10.6151
R667 B.n107 B.n0 10.6151
R668 B.n391 B.n1 10.6151
R669 B.n391 B.n390 10.6151
R670 B.n390 B.n389 10.6151
R671 B.n389 B.n4 10.6151
R672 B.n385 B.n4 10.6151
R673 B.n385 B.n384 10.6151
R674 B.n384 B.n383 10.6151
R675 B.n383 B.n6 10.6151
R676 B.n379 B.n6 10.6151
R677 B.n379 B.n378 10.6151
R678 B.n378 B.n377 10.6151
R679 B.n377 B.n8 10.6151
R680 B.n373 B.n8 10.6151
R681 B.n373 B.n372 10.6151
R682 B.n372 B.n371 10.6151
R683 B.n371 B.n10 10.6151
R684 B.n367 B.n10 10.6151
R685 B.n367 B.n366 10.6151
R686 B.n366 B.n365 10.6151
R687 B.n365 B.n12 10.6151
R688 B.n361 B.n12 10.6151
R689 B.n361 B.n360 10.6151
R690 B.n360 B.n359 10.6151
R691 B.n359 B.n14 10.6151
R692 B.n355 B.n14 10.6151
R693 B.n355 B.n354 10.6151
R694 B.n354 B.n353 10.6151
R695 B.n353 B.n16 10.6151
R696 B.n349 B.n16 10.6151
R697 B.n349 B.n348 10.6151
R698 B.n329 B.n328 6.5566
R699 B.n316 B.n32 6.5566
R700 B.n170 B.n169 6.5566
R701 B.n182 B.n78 6.5566
R702 B.n330 B.n329 4.05904
R703 B.n313 B.n32 4.05904
R704 B.n169 B.n168 4.05904
R705 B.n185 B.n78 4.05904
R706 B.n395 B.n0 2.81026
R707 B.n395 B.n1 2.81026
C0 VDD1 VP 0.872506f
C1 VDD1 w_n2514_n1322# 1.17911f
C2 VDD1 VN 0.155186f
C3 VP VDD2 0.379024f
C4 w_n2514_n1322# VDD2 1.21571f
C5 VN VDD2 0.650442f
C6 VTAIL VP 1.09935f
C7 VTAIL w_n2514_n1322# 1.32774f
C8 VTAIL VN 1.08522f
C9 VP w_n2514_n1322# 3.65552f
C10 VP VN 4.00358f
C11 VN w_n2514_n1322# 3.33866f
C12 VDD1 B 1.00444f
C13 B VDD2 1.04332f
C14 VTAIL B 1.44346f
C15 VDD1 VDD2 0.775511f
C16 VDD1 VTAIL 2.67169f
C17 B VP 1.56481f
C18 B w_n2514_n1322# 7.00033f
C19 B VN 1.03214f
C20 VTAIL VDD2 2.73106f
C21 VDD2 VSUBS 0.642639f
C22 VDD1 VSUBS 2.527258f
C23 VTAIL VSUBS 0.384639f
C24 VN VSUBS 6.08151f
C25 VP VSUBS 1.481802f
C26 B VSUBS 3.525302f
C27 w_n2514_n1322# VSUBS 42.5067f
C28 B.n0 VSUBS 0.006173f
C29 B.n1 VSUBS 0.006173f
C30 B.n2 VSUBS 0.009762f
C31 B.n3 VSUBS 0.009762f
C32 B.n4 VSUBS 0.009762f
C33 B.n5 VSUBS 0.009762f
C34 B.n6 VSUBS 0.009762f
C35 B.n7 VSUBS 0.009762f
C36 B.n8 VSUBS 0.009762f
C37 B.n9 VSUBS 0.009762f
C38 B.n10 VSUBS 0.009762f
C39 B.n11 VSUBS 0.009762f
C40 B.n12 VSUBS 0.009762f
C41 B.n13 VSUBS 0.009762f
C42 B.n14 VSUBS 0.009762f
C43 B.n15 VSUBS 0.009762f
C44 B.n16 VSUBS 0.009762f
C45 B.n17 VSUBS 0.020332f
C46 B.n18 VSUBS 0.009762f
C47 B.n19 VSUBS 0.009762f
C48 B.n20 VSUBS 0.009762f
C49 B.n21 VSUBS 0.009762f
C50 B.n22 VSUBS 0.009762f
C51 B.n23 VSUBS 0.009762f
C52 B.t11 VSUBS 0.041797f
C53 B.t10 VSUBS 0.060431f
C54 B.t9 VSUBS 0.438039f
C55 B.n24 VSUBS 0.112431f
C56 B.n25 VSUBS 0.09326f
C57 B.n26 VSUBS 0.009762f
C58 B.n27 VSUBS 0.009762f
C59 B.n28 VSUBS 0.009762f
C60 B.n29 VSUBS 0.009762f
C61 B.t8 VSUBS 0.041797f
C62 B.t7 VSUBS 0.060431f
C63 B.t6 VSUBS 0.438039f
C64 B.n30 VSUBS 0.112431f
C65 B.n31 VSUBS 0.09326f
C66 B.n32 VSUBS 0.022617f
C67 B.n33 VSUBS 0.009762f
C68 B.n34 VSUBS 0.009762f
C69 B.n35 VSUBS 0.009762f
C70 B.n36 VSUBS 0.009762f
C71 B.n37 VSUBS 0.009762f
C72 B.n38 VSUBS 0.020268f
C73 B.n39 VSUBS 0.009762f
C74 B.n40 VSUBS 0.009762f
C75 B.n41 VSUBS 0.009762f
C76 B.n42 VSUBS 0.009762f
C77 B.n43 VSUBS 0.009762f
C78 B.n44 VSUBS 0.009762f
C79 B.n45 VSUBS 0.009762f
C80 B.n46 VSUBS 0.009762f
C81 B.n47 VSUBS 0.009762f
C82 B.n48 VSUBS 0.009762f
C83 B.n49 VSUBS 0.009762f
C84 B.n50 VSUBS 0.009762f
C85 B.n51 VSUBS 0.009762f
C86 B.n52 VSUBS 0.009762f
C87 B.n53 VSUBS 0.009762f
C88 B.n54 VSUBS 0.009762f
C89 B.n55 VSUBS 0.009762f
C90 B.n56 VSUBS 0.009762f
C91 B.n57 VSUBS 0.009762f
C92 B.n58 VSUBS 0.009762f
C93 B.n59 VSUBS 0.009762f
C94 B.n60 VSUBS 0.009762f
C95 B.n61 VSUBS 0.009762f
C96 B.n62 VSUBS 0.009762f
C97 B.n63 VSUBS 0.009762f
C98 B.n64 VSUBS 0.009762f
C99 B.n65 VSUBS 0.009762f
C100 B.n66 VSUBS 0.009762f
C101 B.n67 VSUBS 0.009762f
C102 B.n68 VSUBS 0.009762f
C103 B.n69 VSUBS 0.009762f
C104 B.n70 VSUBS 0.021587f
C105 B.n71 VSUBS 0.009762f
C106 B.n72 VSUBS 0.009762f
C107 B.n73 VSUBS 0.009762f
C108 B.n74 VSUBS 0.009762f
C109 B.n75 VSUBS 0.009762f
C110 B.t4 VSUBS 0.041797f
C111 B.t5 VSUBS 0.060431f
C112 B.t3 VSUBS 0.438039f
C113 B.n76 VSUBS 0.112431f
C114 B.n77 VSUBS 0.09326f
C115 B.n78 VSUBS 0.022617f
C116 B.n79 VSUBS 0.009762f
C117 B.n80 VSUBS 0.009762f
C118 B.n81 VSUBS 0.009762f
C119 B.n82 VSUBS 0.009762f
C120 B.n83 VSUBS 0.009762f
C121 B.t1 VSUBS 0.041797f
C122 B.t2 VSUBS 0.060431f
C123 B.t0 VSUBS 0.438039f
C124 B.n84 VSUBS 0.112431f
C125 B.n85 VSUBS 0.09326f
C126 B.n86 VSUBS 0.009762f
C127 B.n87 VSUBS 0.009762f
C128 B.n88 VSUBS 0.009762f
C129 B.n89 VSUBS 0.009762f
C130 B.n90 VSUBS 0.009762f
C131 B.n91 VSUBS 0.020332f
C132 B.n92 VSUBS 0.009762f
C133 B.n93 VSUBS 0.009762f
C134 B.n94 VSUBS 0.009762f
C135 B.n95 VSUBS 0.009762f
C136 B.n96 VSUBS 0.009762f
C137 B.n97 VSUBS 0.009762f
C138 B.n98 VSUBS 0.009762f
C139 B.n99 VSUBS 0.009762f
C140 B.n100 VSUBS 0.009762f
C141 B.n101 VSUBS 0.009762f
C142 B.n102 VSUBS 0.009762f
C143 B.n103 VSUBS 0.009762f
C144 B.n104 VSUBS 0.009762f
C145 B.n105 VSUBS 0.009762f
C146 B.n106 VSUBS 0.009762f
C147 B.n107 VSUBS 0.009762f
C148 B.n108 VSUBS 0.009762f
C149 B.n109 VSUBS 0.009762f
C150 B.n110 VSUBS 0.009762f
C151 B.n111 VSUBS 0.009762f
C152 B.n112 VSUBS 0.009762f
C153 B.n113 VSUBS 0.009762f
C154 B.n114 VSUBS 0.009762f
C155 B.n115 VSUBS 0.009762f
C156 B.n116 VSUBS 0.009762f
C157 B.n117 VSUBS 0.009762f
C158 B.n118 VSUBS 0.009762f
C159 B.n119 VSUBS 0.009762f
C160 B.n120 VSUBS 0.009762f
C161 B.n121 VSUBS 0.009762f
C162 B.n122 VSUBS 0.009762f
C163 B.n123 VSUBS 0.009762f
C164 B.n124 VSUBS 0.009762f
C165 B.n125 VSUBS 0.009762f
C166 B.n126 VSUBS 0.009762f
C167 B.n127 VSUBS 0.009762f
C168 B.n128 VSUBS 0.009762f
C169 B.n129 VSUBS 0.009762f
C170 B.n130 VSUBS 0.009762f
C171 B.n131 VSUBS 0.009762f
C172 B.n132 VSUBS 0.009762f
C173 B.n133 VSUBS 0.009762f
C174 B.n134 VSUBS 0.009762f
C175 B.n135 VSUBS 0.009762f
C176 B.n136 VSUBS 0.009762f
C177 B.n137 VSUBS 0.009762f
C178 B.n138 VSUBS 0.009762f
C179 B.n139 VSUBS 0.009762f
C180 B.n140 VSUBS 0.009762f
C181 B.n141 VSUBS 0.009762f
C182 B.n142 VSUBS 0.009762f
C183 B.n143 VSUBS 0.009762f
C184 B.n144 VSUBS 0.009762f
C185 B.n145 VSUBS 0.009762f
C186 B.n146 VSUBS 0.009762f
C187 B.n147 VSUBS 0.009762f
C188 B.n148 VSUBS 0.009762f
C189 B.n149 VSUBS 0.009762f
C190 B.n150 VSUBS 0.020332f
C191 B.n151 VSUBS 0.021587f
C192 B.n152 VSUBS 0.021587f
C193 B.n153 VSUBS 0.009762f
C194 B.n154 VSUBS 0.009762f
C195 B.n155 VSUBS 0.009762f
C196 B.n156 VSUBS 0.009762f
C197 B.n157 VSUBS 0.009762f
C198 B.n158 VSUBS 0.009762f
C199 B.n159 VSUBS 0.009762f
C200 B.n160 VSUBS 0.009762f
C201 B.n161 VSUBS 0.009762f
C202 B.n162 VSUBS 0.009762f
C203 B.n163 VSUBS 0.009762f
C204 B.n164 VSUBS 0.009762f
C205 B.n165 VSUBS 0.009762f
C206 B.n166 VSUBS 0.009762f
C207 B.n167 VSUBS 0.009762f
C208 B.n168 VSUBS 0.006747f
C209 B.n169 VSUBS 0.022617f
C210 B.n170 VSUBS 0.007896f
C211 B.n171 VSUBS 0.009762f
C212 B.n172 VSUBS 0.009762f
C213 B.n173 VSUBS 0.009762f
C214 B.n174 VSUBS 0.009762f
C215 B.n175 VSUBS 0.009762f
C216 B.n176 VSUBS 0.009762f
C217 B.n177 VSUBS 0.009762f
C218 B.n178 VSUBS 0.009762f
C219 B.n179 VSUBS 0.009762f
C220 B.n180 VSUBS 0.009762f
C221 B.n181 VSUBS 0.009762f
C222 B.n182 VSUBS 0.007896f
C223 B.n183 VSUBS 0.009762f
C224 B.n184 VSUBS 0.009762f
C225 B.n185 VSUBS 0.006747f
C226 B.n186 VSUBS 0.009762f
C227 B.n187 VSUBS 0.009762f
C228 B.n188 VSUBS 0.009762f
C229 B.n189 VSUBS 0.009762f
C230 B.n190 VSUBS 0.009762f
C231 B.n191 VSUBS 0.009762f
C232 B.n192 VSUBS 0.009762f
C233 B.n193 VSUBS 0.009762f
C234 B.n194 VSUBS 0.009762f
C235 B.n195 VSUBS 0.009762f
C236 B.n196 VSUBS 0.009762f
C237 B.n197 VSUBS 0.009762f
C238 B.n198 VSUBS 0.009762f
C239 B.n199 VSUBS 0.009762f
C240 B.n200 VSUBS 0.009762f
C241 B.n201 VSUBS 0.021587f
C242 B.n202 VSUBS 0.020332f
C243 B.n203 VSUBS 0.020332f
C244 B.n204 VSUBS 0.009762f
C245 B.n205 VSUBS 0.009762f
C246 B.n206 VSUBS 0.009762f
C247 B.n207 VSUBS 0.009762f
C248 B.n208 VSUBS 0.009762f
C249 B.n209 VSUBS 0.009762f
C250 B.n210 VSUBS 0.009762f
C251 B.n211 VSUBS 0.009762f
C252 B.n212 VSUBS 0.009762f
C253 B.n213 VSUBS 0.009762f
C254 B.n214 VSUBS 0.009762f
C255 B.n215 VSUBS 0.009762f
C256 B.n216 VSUBS 0.009762f
C257 B.n217 VSUBS 0.009762f
C258 B.n218 VSUBS 0.009762f
C259 B.n219 VSUBS 0.009762f
C260 B.n220 VSUBS 0.009762f
C261 B.n221 VSUBS 0.009762f
C262 B.n222 VSUBS 0.009762f
C263 B.n223 VSUBS 0.009762f
C264 B.n224 VSUBS 0.009762f
C265 B.n225 VSUBS 0.009762f
C266 B.n226 VSUBS 0.009762f
C267 B.n227 VSUBS 0.009762f
C268 B.n228 VSUBS 0.009762f
C269 B.n229 VSUBS 0.009762f
C270 B.n230 VSUBS 0.009762f
C271 B.n231 VSUBS 0.009762f
C272 B.n232 VSUBS 0.009762f
C273 B.n233 VSUBS 0.009762f
C274 B.n234 VSUBS 0.009762f
C275 B.n235 VSUBS 0.009762f
C276 B.n236 VSUBS 0.009762f
C277 B.n237 VSUBS 0.009762f
C278 B.n238 VSUBS 0.009762f
C279 B.n239 VSUBS 0.009762f
C280 B.n240 VSUBS 0.009762f
C281 B.n241 VSUBS 0.009762f
C282 B.n242 VSUBS 0.009762f
C283 B.n243 VSUBS 0.009762f
C284 B.n244 VSUBS 0.009762f
C285 B.n245 VSUBS 0.009762f
C286 B.n246 VSUBS 0.009762f
C287 B.n247 VSUBS 0.009762f
C288 B.n248 VSUBS 0.009762f
C289 B.n249 VSUBS 0.009762f
C290 B.n250 VSUBS 0.009762f
C291 B.n251 VSUBS 0.009762f
C292 B.n252 VSUBS 0.009762f
C293 B.n253 VSUBS 0.009762f
C294 B.n254 VSUBS 0.009762f
C295 B.n255 VSUBS 0.009762f
C296 B.n256 VSUBS 0.009762f
C297 B.n257 VSUBS 0.009762f
C298 B.n258 VSUBS 0.009762f
C299 B.n259 VSUBS 0.009762f
C300 B.n260 VSUBS 0.009762f
C301 B.n261 VSUBS 0.009762f
C302 B.n262 VSUBS 0.009762f
C303 B.n263 VSUBS 0.009762f
C304 B.n264 VSUBS 0.009762f
C305 B.n265 VSUBS 0.009762f
C306 B.n266 VSUBS 0.009762f
C307 B.n267 VSUBS 0.009762f
C308 B.n268 VSUBS 0.009762f
C309 B.n269 VSUBS 0.009762f
C310 B.n270 VSUBS 0.009762f
C311 B.n271 VSUBS 0.009762f
C312 B.n272 VSUBS 0.009762f
C313 B.n273 VSUBS 0.009762f
C314 B.n274 VSUBS 0.009762f
C315 B.n275 VSUBS 0.009762f
C316 B.n276 VSUBS 0.009762f
C317 B.n277 VSUBS 0.009762f
C318 B.n278 VSUBS 0.009762f
C319 B.n279 VSUBS 0.009762f
C320 B.n280 VSUBS 0.009762f
C321 B.n281 VSUBS 0.009762f
C322 B.n282 VSUBS 0.009762f
C323 B.n283 VSUBS 0.009762f
C324 B.n284 VSUBS 0.009762f
C325 B.n285 VSUBS 0.009762f
C326 B.n286 VSUBS 0.009762f
C327 B.n287 VSUBS 0.009762f
C328 B.n288 VSUBS 0.009762f
C329 B.n289 VSUBS 0.009762f
C330 B.n290 VSUBS 0.009762f
C331 B.n291 VSUBS 0.009762f
C332 B.n292 VSUBS 0.009762f
C333 B.n293 VSUBS 0.009762f
C334 B.n294 VSUBS 0.009762f
C335 B.n295 VSUBS 0.021651f
C336 B.n296 VSUBS 0.020332f
C337 B.n297 VSUBS 0.021587f
C338 B.n298 VSUBS 0.009762f
C339 B.n299 VSUBS 0.009762f
C340 B.n300 VSUBS 0.009762f
C341 B.n301 VSUBS 0.009762f
C342 B.n302 VSUBS 0.009762f
C343 B.n303 VSUBS 0.009762f
C344 B.n304 VSUBS 0.009762f
C345 B.n305 VSUBS 0.009762f
C346 B.n306 VSUBS 0.009762f
C347 B.n307 VSUBS 0.009762f
C348 B.n308 VSUBS 0.009762f
C349 B.n309 VSUBS 0.009762f
C350 B.n310 VSUBS 0.009762f
C351 B.n311 VSUBS 0.009762f
C352 B.n312 VSUBS 0.009762f
C353 B.n313 VSUBS 0.006747f
C354 B.n314 VSUBS 0.009762f
C355 B.n315 VSUBS 0.009762f
C356 B.n316 VSUBS 0.007896f
C357 B.n317 VSUBS 0.009762f
C358 B.n318 VSUBS 0.009762f
C359 B.n319 VSUBS 0.009762f
C360 B.n320 VSUBS 0.009762f
C361 B.n321 VSUBS 0.009762f
C362 B.n322 VSUBS 0.009762f
C363 B.n323 VSUBS 0.009762f
C364 B.n324 VSUBS 0.009762f
C365 B.n325 VSUBS 0.009762f
C366 B.n326 VSUBS 0.009762f
C367 B.n327 VSUBS 0.009762f
C368 B.n328 VSUBS 0.007896f
C369 B.n329 VSUBS 0.022617f
C370 B.n330 VSUBS 0.006747f
C371 B.n331 VSUBS 0.009762f
C372 B.n332 VSUBS 0.009762f
C373 B.n333 VSUBS 0.009762f
C374 B.n334 VSUBS 0.009762f
C375 B.n335 VSUBS 0.009762f
C376 B.n336 VSUBS 0.009762f
C377 B.n337 VSUBS 0.009762f
C378 B.n338 VSUBS 0.009762f
C379 B.n339 VSUBS 0.009762f
C380 B.n340 VSUBS 0.009762f
C381 B.n341 VSUBS 0.009762f
C382 B.n342 VSUBS 0.009762f
C383 B.n343 VSUBS 0.009762f
C384 B.n344 VSUBS 0.009762f
C385 B.n345 VSUBS 0.009762f
C386 B.n346 VSUBS 0.021587f
C387 B.n347 VSUBS 0.021587f
C388 B.n348 VSUBS 0.020332f
C389 B.n349 VSUBS 0.009762f
C390 B.n350 VSUBS 0.009762f
C391 B.n351 VSUBS 0.009762f
C392 B.n352 VSUBS 0.009762f
C393 B.n353 VSUBS 0.009762f
C394 B.n354 VSUBS 0.009762f
C395 B.n355 VSUBS 0.009762f
C396 B.n356 VSUBS 0.009762f
C397 B.n357 VSUBS 0.009762f
C398 B.n358 VSUBS 0.009762f
C399 B.n359 VSUBS 0.009762f
C400 B.n360 VSUBS 0.009762f
C401 B.n361 VSUBS 0.009762f
C402 B.n362 VSUBS 0.009762f
C403 B.n363 VSUBS 0.009762f
C404 B.n364 VSUBS 0.009762f
C405 B.n365 VSUBS 0.009762f
C406 B.n366 VSUBS 0.009762f
C407 B.n367 VSUBS 0.009762f
C408 B.n368 VSUBS 0.009762f
C409 B.n369 VSUBS 0.009762f
C410 B.n370 VSUBS 0.009762f
C411 B.n371 VSUBS 0.009762f
C412 B.n372 VSUBS 0.009762f
C413 B.n373 VSUBS 0.009762f
C414 B.n374 VSUBS 0.009762f
C415 B.n375 VSUBS 0.009762f
C416 B.n376 VSUBS 0.009762f
C417 B.n377 VSUBS 0.009762f
C418 B.n378 VSUBS 0.009762f
C419 B.n379 VSUBS 0.009762f
C420 B.n380 VSUBS 0.009762f
C421 B.n381 VSUBS 0.009762f
C422 B.n382 VSUBS 0.009762f
C423 B.n383 VSUBS 0.009762f
C424 B.n384 VSUBS 0.009762f
C425 B.n385 VSUBS 0.009762f
C426 B.n386 VSUBS 0.009762f
C427 B.n387 VSUBS 0.009762f
C428 B.n388 VSUBS 0.009762f
C429 B.n389 VSUBS 0.009762f
C430 B.n390 VSUBS 0.009762f
C431 B.n391 VSUBS 0.009762f
C432 B.n392 VSUBS 0.009762f
C433 B.n393 VSUBS 0.009762f
C434 B.n394 VSUBS 0.009762f
C435 B.n395 VSUBS 0.022104f
C436 VDD2.n0 VSUBS 0.018977f
C437 VDD2.n1 VSUBS 0.05048f
C438 VDD2.t0 VSUBS 0.048749f
C439 VDD2.n2 VSUBS 0.046503f
C440 VDD2.n3 VSUBS 0.012417f
C441 VDD2.n4 VSUBS 0.009891f
C442 VDD2.n5 VSUBS 0.106782f
C443 VDD2.n6 VSUBS 0.331669f
C444 VDD2.n7 VSUBS 0.018977f
C445 VDD2.n8 VSUBS 0.05048f
C446 VDD2.t1 VSUBS 0.048749f
C447 VDD2.n9 VSUBS 0.046503f
C448 VDD2.n10 VSUBS 0.012417f
C449 VDD2.n11 VSUBS 0.009891f
C450 VDD2.n12 VSUBS 0.106782f
C451 VDD2.n13 VSUBS 0.038897f
C452 VDD2.n14 VSUBS 1.58986f
C453 VN.t1 VSUBS 1.24479f
C454 VN.t0 VSUBS 2.26904f
C455 VDD1.n0 VSUBS 0.018511f
C456 VDD1.n1 VSUBS 0.04924f
C457 VDD1.t1 VSUBS 0.047551f
C458 VDD1.n2 VSUBS 0.045361f
C459 VDD1.n3 VSUBS 0.012112f
C460 VDD1.n4 VSUBS 0.009648f
C461 VDD1.n5 VSUBS 0.104159f
C462 VDD1.n6 VSUBS 0.039451f
C463 VDD1.n7 VSUBS 0.018511f
C464 VDD1.n8 VSUBS 0.04924f
C465 VDD1.t0 VSUBS 0.047551f
C466 VDD1.n9 VSUBS 0.045361f
C467 VDD1.n10 VSUBS 0.012112f
C468 VDD1.n11 VSUBS 0.009648f
C469 VDD1.n12 VSUBS 0.104159f
C470 VDD1.n13 VSUBS 0.355905f
C471 VTAIL.n0 VSUBS 0.023288f
C472 VTAIL.n1 VSUBS 0.061947f
C473 VTAIL.t3 VSUBS 0.059822f
C474 VTAIL.n2 VSUBS 0.057066f
C475 VTAIL.n3 VSUBS 0.015237f
C476 VTAIL.n4 VSUBS 0.012137f
C477 VTAIL.n5 VSUBS 0.131037f
C478 VTAIL.n6 VSUBS 0.032157f
C479 VTAIL.n7 VSUBS 1.02209f
C480 VTAIL.n8 VSUBS 0.023288f
C481 VTAIL.n9 VSUBS 0.061947f
C482 VTAIL.t0 VSUBS 0.059822f
C483 VTAIL.n10 VSUBS 0.057066f
C484 VTAIL.n11 VSUBS 0.015237f
C485 VTAIL.n12 VSUBS 0.012137f
C486 VTAIL.n13 VSUBS 0.131037f
C487 VTAIL.n14 VSUBS 0.032157f
C488 VTAIL.n15 VSUBS 1.0784f
C489 VTAIL.n16 VSUBS 0.023288f
C490 VTAIL.n17 VSUBS 0.061947f
C491 VTAIL.t2 VSUBS 0.059822f
C492 VTAIL.n18 VSUBS 0.057066f
C493 VTAIL.n19 VSUBS 0.015237f
C494 VTAIL.n20 VSUBS 0.012137f
C495 VTAIL.n21 VSUBS 0.131037f
C496 VTAIL.n22 VSUBS 0.032157f
C497 VTAIL.n23 VSUBS 0.836216f
C498 VTAIL.n24 VSUBS 0.023288f
C499 VTAIL.n25 VSUBS 0.061947f
C500 VTAIL.t1 VSUBS 0.059822f
C501 VTAIL.n26 VSUBS 0.057066f
C502 VTAIL.n27 VSUBS 0.015237f
C503 VTAIL.n28 VSUBS 0.012137f
C504 VTAIL.n29 VSUBS 0.131037f
C505 VTAIL.n30 VSUBS 0.032157f
C506 VTAIL.n31 VSUBS 0.737239f
C507 VP.t0 VSUBS 2.41342f
C508 VP.t1 VSUBS 1.31981f
C509 VP.n0 VSUBS 3.77161f
.ends

