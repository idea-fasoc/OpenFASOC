* NGSPICE file created from diff_pair_sample_0292.ext - technology: sky130A

.subckt diff_pair_sample_0292 VTAIL VN VP B VDD2 VDD1
X0 VDD2.t9 VN.t0 VTAIL.t10 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=1.96845 ps=12.26 w=11.93 l=0.67
X1 B.t11 B.t9 B.t10 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=0 ps=0 w=11.93 l=0.67
X2 VTAIL.t2 VP.t0 VDD1.t9 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X3 VDD2.t8 VN.t1 VTAIL.t15 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=4.6527 ps=24.64 w=11.93 l=0.67
X4 VTAIL.t18 VP.t1 VDD1.t8 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X5 VDD2.t7 VN.t2 VTAIL.t16 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X6 VDD1.t7 VP.t2 VTAIL.t5 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X7 VTAIL.t0 VP.t3 VDD1.t6 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X8 VTAIL.t12 VN.t3 VDD2.t6 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X9 VDD2.t5 VN.t4 VTAIL.t9 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=4.6527 ps=24.64 w=11.93 l=0.67
X10 B.t8 B.t6 B.t7 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=0 ps=0 w=11.93 l=0.67
X11 VTAIL.t19 VP.t4 VDD1.t5 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X12 B.t5 B.t3 B.t4 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=0 ps=0 w=11.93 l=0.67
X13 VDD1.t4 VP.t5 VTAIL.t1 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=4.6527 ps=24.64 w=11.93 l=0.67
X14 VDD2.t4 VN.t5 VTAIL.t13 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X15 VDD1.t3 VP.t6 VTAIL.t3 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=4.6527 ps=24.64 w=11.93 l=0.67
X16 VTAIL.t17 VN.t6 VDD2.t3 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X17 VTAIL.t11 VN.t7 VDD2.t2 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X18 VDD1.t2 VP.t7 VTAIL.t7 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X19 VTAIL.t8 VN.t8 VDD2.t1 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=1.96845 pd=12.26 as=1.96845 ps=12.26 w=11.93 l=0.67
X20 B.t2 B.t0 B.t1 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=0 ps=0 w=11.93 l=0.67
X21 VDD2.t0 VN.t9 VTAIL.t14 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=1.96845 ps=12.26 w=11.93 l=0.67
X22 VDD1.t1 VP.t8 VTAIL.t6 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=1.96845 ps=12.26 w=11.93 l=0.67
X23 VDD1.t0 VP.t9 VTAIL.t4 w_n2170_n3354# sky130_fd_pr__pfet_01v8 ad=4.6527 pd=24.64 as=1.96845 ps=12.26 w=11.93 l=0.67
R0 VN.n3 VN.t9 509.111
R1 VN.n17 VN.t4 509.111
R2 VN.n4 VN.t7 488.115
R3 VN.n6 VN.t5 488.115
R4 VN.n10 VN.t3 488.115
R5 VN.n12 VN.t1 488.115
R6 VN.n18 VN.t8 488.115
R7 VN.n20 VN.t2 488.115
R8 VN.n24 VN.t6 488.115
R9 VN.n26 VN.t0 488.115
R10 VN.n13 VN.n12 161.3
R11 VN.n27 VN.n26 161.3
R12 VN.n25 VN.n14 161.3
R13 VN.n24 VN.n23 161.3
R14 VN.n22 VN.n15 161.3
R15 VN.n21 VN.n20 161.3
R16 VN.n19 VN.n16 161.3
R17 VN.n11 VN.n0 161.3
R18 VN.n10 VN.n9 161.3
R19 VN.n8 VN.n1 161.3
R20 VN.n7 VN.n6 161.3
R21 VN.n5 VN.n2 161.3
R22 VN.n17 VN.n16 44.8515
R23 VN.n3 VN.n2 44.8515
R24 VN VN.n27 42.8963
R25 VN.n5 VN.n4 24.1005
R26 VN.n6 VN.n5 24.1005
R27 VN.n6 VN.n1 24.1005
R28 VN.n10 VN.n1 24.1005
R29 VN.n11 VN.n10 24.1005
R30 VN.n12 VN.n11 24.1005
R31 VN.n20 VN.n19 24.1005
R32 VN.n19 VN.n18 24.1005
R33 VN.n24 VN.n15 24.1005
R34 VN.n20 VN.n15 24.1005
R35 VN.n26 VN.n25 24.1005
R36 VN.n25 VN.n24 24.1005
R37 VN.n4 VN.n3 20.9471
R38 VN.n18 VN.n17 20.9471
R39 VN.n27 VN.n14 0.189894
R40 VN.n23 VN.n14 0.189894
R41 VN.n23 VN.n22 0.189894
R42 VN.n22 VN.n21 0.189894
R43 VN.n21 VN.n16 0.189894
R44 VN.n7 VN.n2 0.189894
R45 VN.n8 VN.n7 0.189894
R46 VN.n9 VN.n8 0.189894
R47 VN.n9 VN.n0 0.189894
R48 VN.n13 VN.n0 0.189894
R49 VN VN.n13 0.0516364
R50 VTAIL.n276 VTAIL.n275 756.745
R51 VTAIL.n66 VTAIL.n65 756.745
R52 VTAIL.n210 VTAIL.n209 756.745
R53 VTAIL.n140 VTAIL.n139 756.745
R54 VTAIL.n235 VTAIL.n234 585
R55 VTAIL.n237 VTAIL.n236 585
R56 VTAIL.n230 VTAIL.n229 585
R57 VTAIL.n243 VTAIL.n242 585
R58 VTAIL.n245 VTAIL.n244 585
R59 VTAIL.n226 VTAIL.n225 585
R60 VTAIL.n251 VTAIL.n250 585
R61 VTAIL.n253 VTAIL.n252 585
R62 VTAIL.n222 VTAIL.n221 585
R63 VTAIL.n259 VTAIL.n258 585
R64 VTAIL.n261 VTAIL.n260 585
R65 VTAIL.n218 VTAIL.n217 585
R66 VTAIL.n267 VTAIL.n266 585
R67 VTAIL.n269 VTAIL.n268 585
R68 VTAIL.n214 VTAIL.n213 585
R69 VTAIL.n275 VTAIL.n274 585
R70 VTAIL.n25 VTAIL.n24 585
R71 VTAIL.n27 VTAIL.n26 585
R72 VTAIL.n20 VTAIL.n19 585
R73 VTAIL.n33 VTAIL.n32 585
R74 VTAIL.n35 VTAIL.n34 585
R75 VTAIL.n16 VTAIL.n15 585
R76 VTAIL.n41 VTAIL.n40 585
R77 VTAIL.n43 VTAIL.n42 585
R78 VTAIL.n12 VTAIL.n11 585
R79 VTAIL.n49 VTAIL.n48 585
R80 VTAIL.n51 VTAIL.n50 585
R81 VTAIL.n8 VTAIL.n7 585
R82 VTAIL.n57 VTAIL.n56 585
R83 VTAIL.n59 VTAIL.n58 585
R84 VTAIL.n4 VTAIL.n3 585
R85 VTAIL.n65 VTAIL.n64 585
R86 VTAIL.n209 VTAIL.n208 585
R87 VTAIL.n148 VTAIL.n147 585
R88 VTAIL.n203 VTAIL.n202 585
R89 VTAIL.n201 VTAIL.n200 585
R90 VTAIL.n152 VTAIL.n151 585
R91 VTAIL.n195 VTAIL.n194 585
R92 VTAIL.n193 VTAIL.n192 585
R93 VTAIL.n156 VTAIL.n155 585
R94 VTAIL.n187 VTAIL.n186 585
R95 VTAIL.n185 VTAIL.n184 585
R96 VTAIL.n160 VTAIL.n159 585
R97 VTAIL.n179 VTAIL.n178 585
R98 VTAIL.n177 VTAIL.n176 585
R99 VTAIL.n164 VTAIL.n163 585
R100 VTAIL.n171 VTAIL.n170 585
R101 VTAIL.n169 VTAIL.n168 585
R102 VTAIL.n139 VTAIL.n138 585
R103 VTAIL.n78 VTAIL.n77 585
R104 VTAIL.n133 VTAIL.n132 585
R105 VTAIL.n131 VTAIL.n130 585
R106 VTAIL.n82 VTAIL.n81 585
R107 VTAIL.n125 VTAIL.n124 585
R108 VTAIL.n123 VTAIL.n122 585
R109 VTAIL.n86 VTAIL.n85 585
R110 VTAIL.n117 VTAIL.n116 585
R111 VTAIL.n115 VTAIL.n114 585
R112 VTAIL.n90 VTAIL.n89 585
R113 VTAIL.n109 VTAIL.n108 585
R114 VTAIL.n107 VTAIL.n106 585
R115 VTAIL.n94 VTAIL.n93 585
R116 VTAIL.n101 VTAIL.n100 585
R117 VTAIL.n99 VTAIL.n98 585
R118 VTAIL.n167 VTAIL.t1 327.466
R119 VTAIL.n97 VTAIL.t9 327.466
R120 VTAIL.n233 VTAIL.t15 327.466
R121 VTAIL.n23 VTAIL.t3 327.466
R122 VTAIL.n236 VTAIL.n235 171.744
R123 VTAIL.n236 VTAIL.n229 171.744
R124 VTAIL.n243 VTAIL.n229 171.744
R125 VTAIL.n244 VTAIL.n243 171.744
R126 VTAIL.n244 VTAIL.n225 171.744
R127 VTAIL.n251 VTAIL.n225 171.744
R128 VTAIL.n252 VTAIL.n251 171.744
R129 VTAIL.n252 VTAIL.n221 171.744
R130 VTAIL.n259 VTAIL.n221 171.744
R131 VTAIL.n260 VTAIL.n259 171.744
R132 VTAIL.n260 VTAIL.n217 171.744
R133 VTAIL.n267 VTAIL.n217 171.744
R134 VTAIL.n268 VTAIL.n267 171.744
R135 VTAIL.n268 VTAIL.n213 171.744
R136 VTAIL.n275 VTAIL.n213 171.744
R137 VTAIL.n26 VTAIL.n25 171.744
R138 VTAIL.n26 VTAIL.n19 171.744
R139 VTAIL.n33 VTAIL.n19 171.744
R140 VTAIL.n34 VTAIL.n33 171.744
R141 VTAIL.n34 VTAIL.n15 171.744
R142 VTAIL.n41 VTAIL.n15 171.744
R143 VTAIL.n42 VTAIL.n41 171.744
R144 VTAIL.n42 VTAIL.n11 171.744
R145 VTAIL.n49 VTAIL.n11 171.744
R146 VTAIL.n50 VTAIL.n49 171.744
R147 VTAIL.n50 VTAIL.n7 171.744
R148 VTAIL.n57 VTAIL.n7 171.744
R149 VTAIL.n58 VTAIL.n57 171.744
R150 VTAIL.n58 VTAIL.n3 171.744
R151 VTAIL.n65 VTAIL.n3 171.744
R152 VTAIL.n209 VTAIL.n147 171.744
R153 VTAIL.n202 VTAIL.n147 171.744
R154 VTAIL.n202 VTAIL.n201 171.744
R155 VTAIL.n201 VTAIL.n151 171.744
R156 VTAIL.n194 VTAIL.n151 171.744
R157 VTAIL.n194 VTAIL.n193 171.744
R158 VTAIL.n193 VTAIL.n155 171.744
R159 VTAIL.n186 VTAIL.n155 171.744
R160 VTAIL.n186 VTAIL.n185 171.744
R161 VTAIL.n185 VTAIL.n159 171.744
R162 VTAIL.n178 VTAIL.n159 171.744
R163 VTAIL.n178 VTAIL.n177 171.744
R164 VTAIL.n177 VTAIL.n163 171.744
R165 VTAIL.n170 VTAIL.n163 171.744
R166 VTAIL.n170 VTAIL.n169 171.744
R167 VTAIL.n139 VTAIL.n77 171.744
R168 VTAIL.n132 VTAIL.n77 171.744
R169 VTAIL.n132 VTAIL.n131 171.744
R170 VTAIL.n131 VTAIL.n81 171.744
R171 VTAIL.n124 VTAIL.n81 171.744
R172 VTAIL.n124 VTAIL.n123 171.744
R173 VTAIL.n123 VTAIL.n85 171.744
R174 VTAIL.n116 VTAIL.n85 171.744
R175 VTAIL.n116 VTAIL.n115 171.744
R176 VTAIL.n115 VTAIL.n89 171.744
R177 VTAIL.n108 VTAIL.n89 171.744
R178 VTAIL.n108 VTAIL.n107 171.744
R179 VTAIL.n107 VTAIL.n93 171.744
R180 VTAIL.n100 VTAIL.n93 171.744
R181 VTAIL.n100 VTAIL.n99 171.744
R182 VTAIL.n235 VTAIL.t15 85.8723
R183 VTAIL.n25 VTAIL.t3 85.8723
R184 VTAIL.n169 VTAIL.t1 85.8723
R185 VTAIL.n99 VTAIL.t9 85.8723
R186 VTAIL.n145 VTAIL.n144 60.0341
R187 VTAIL.n143 VTAIL.n142 60.0341
R188 VTAIL.n75 VTAIL.n74 60.0341
R189 VTAIL.n73 VTAIL.n72 60.0341
R190 VTAIL.n279 VTAIL.n278 60.0339
R191 VTAIL.n1 VTAIL.n0 60.0339
R192 VTAIL.n69 VTAIL.n68 60.0339
R193 VTAIL.n71 VTAIL.n70 60.0339
R194 VTAIL.n277 VTAIL.n276 34.3187
R195 VTAIL.n67 VTAIL.n66 34.3187
R196 VTAIL.n211 VTAIL.n210 34.3187
R197 VTAIL.n141 VTAIL.n140 34.3187
R198 VTAIL.n73 VTAIL.n71 24.3755
R199 VTAIL.n277 VTAIL.n211 23.5134
R200 VTAIL.n234 VTAIL.n233 16.3895
R201 VTAIL.n24 VTAIL.n23 16.3895
R202 VTAIL.n168 VTAIL.n167 16.3895
R203 VTAIL.n98 VTAIL.n97 16.3895
R204 VTAIL.n237 VTAIL.n232 12.8005
R205 VTAIL.n27 VTAIL.n22 12.8005
R206 VTAIL.n171 VTAIL.n166 12.8005
R207 VTAIL.n101 VTAIL.n96 12.8005
R208 VTAIL.n238 VTAIL.n230 12.0247
R209 VTAIL.n274 VTAIL.n212 12.0247
R210 VTAIL.n28 VTAIL.n20 12.0247
R211 VTAIL.n64 VTAIL.n2 12.0247
R212 VTAIL.n208 VTAIL.n146 12.0247
R213 VTAIL.n172 VTAIL.n164 12.0247
R214 VTAIL.n138 VTAIL.n76 12.0247
R215 VTAIL.n102 VTAIL.n94 12.0247
R216 VTAIL.n242 VTAIL.n241 11.249
R217 VTAIL.n273 VTAIL.n214 11.249
R218 VTAIL.n32 VTAIL.n31 11.249
R219 VTAIL.n63 VTAIL.n4 11.249
R220 VTAIL.n207 VTAIL.n148 11.249
R221 VTAIL.n176 VTAIL.n175 11.249
R222 VTAIL.n137 VTAIL.n78 11.249
R223 VTAIL.n106 VTAIL.n105 11.249
R224 VTAIL.n245 VTAIL.n228 10.4732
R225 VTAIL.n270 VTAIL.n269 10.4732
R226 VTAIL.n35 VTAIL.n18 10.4732
R227 VTAIL.n60 VTAIL.n59 10.4732
R228 VTAIL.n204 VTAIL.n203 10.4732
R229 VTAIL.n179 VTAIL.n162 10.4732
R230 VTAIL.n134 VTAIL.n133 10.4732
R231 VTAIL.n109 VTAIL.n92 10.4732
R232 VTAIL.n246 VTAIL.n226 9.69747
R233 VTAIL.n266 VTAIL.n216 9.69747
R234 VTAIL.n36 VTAIL.n16 9.69747
R235 VTAIL.n56 VTAIL.n6 9.69747
R236 VTAIL.n200 VTAIL.n150 9.69747
R237 VTAIL.n180 VTAIL.n160 9.69747
R238 VTAIL.n130 VTAIL.n80 9.69747
R239 VTAIL.n110 VTAIL.n90 9.69747
R240 VTAIL.n272 VTAIL.n212 9.45567
R241 VTAIL.n62 VTAIL.n2 9.45567
R242 VTAIL.n206 VTAIL.n146 9.45567
R243 VTAIL.n136 VTAIL.n76 9.45567
R244 VTAIL.n257 VTAIL.n256 9.3005
R245 VTAIL.n220 VTAIL.n219 9.3005
R246 VTAIL.n263 VTAIL.n262 9.3005
R247 VTAIL.n265 VTAIL.n264 9.3005
R248 VTAIL.n216 VTAIL.n215 9.3005
R249 VTAIL.n271 VTAIL.n270 9.3005
R250 VTAIL.n273 VTAIL.n272 9.3005
R251 VTAIL.n224 VTAIL.n223 9.3005
R252 VTAIL.n249 VTAIL.n248 9.3005
R253 VTAIL.n247 VTAIL.n246 9.3005
R254 VTAIL.n228 VTAIL.n227 9.3005
R255 VTAIL.n241 VTAIL.n240 9.3005
R256 VTAIL.n239 VTAIL.n238 9.3005
R257 VTAIL.n232 VTAIL.n231 9.3005
R258 VTAIL.n255 VTAIL.n254 9.3005
R259 VTAIL.n47 VTAIL.n46 9.3005
R260 VTAIL.n10 VTAIL.n9 9.3005
R261 VTAIL.n53 VTAIL.n52 9.3005
R262 VTAIL.n55 VTAIL.n54 9.3005
R263 VTAIL.n6 VTAIL.n5 9.3005
R264 VTAIL.n61 VTAIL.n60 9.3005
R265 VTAIL.n63 VTAIL.n62 9.3005
R266 VTAIL.n14 VTAIL.n13 9.3005
R267 VTAIL.n39 VTAIL.n38 9.3005
R268 VTAIL.n37 VTAIL.n36 9.3005
R269 VTAIL.n18 VTAIL.n17 9.3005
R270 VTAIL.n31 VTAIL.n30 9.3005
R271 VTAIL.n29 VTAIL.n28 9.3005
R272 VTAIL.n22 VTAIL.n21 9.3005
R273 VTAIL.n45 VTAIL.n44 9.3005
R274 VTAIL.n207 VTAIL.n206 9.3005
R275 VTAIL.n205 VTAIL.n204 9.3005
R276 VTAIL.n150 VTAIL.n149 9.3005
R277 VTAIL.n199 VTAIL.n198 9.3005
R278 VTAIL.n197 VTAIL.n196 9.3005
R279 VTAIL.n154 VTAIL.n153 9.3005
R280 VTAIL.n191 VTAIL.n190 9.3005
R281 VTAIL.n189 VTAIL.n188 9.3005
R282 VTAIL.n158 VTAIL.n157 9.3005
R283 VTAIL.n183 VTAIL.n182 9.3005
R284 VTAIL.n181 VTAIL.n180 9.3005
R285 VTAIL.n162 VTAIL.n161 9.3005
R286 VTAIL.n175 VTAIL.n174 9.3005
R287 VTAIL.n173 VTAIL.n172 9.3005
R288 VTAIL.n166 VTAIL.n165 9.3005
R289 VTAIL.n84 VTAIL.n83 9.3005
R290 VTAIL.n127 VTAIL.n126 9.3005
R291 VTAIL.n129 VTAIL.n128 9.3005
R292 VTAIL.n80 VTAIL.n79 9.3005
R293 VTAIL.n135 VTAIL.n134 9.3005
R294 VTAIL.n137 VTAIL.n136 9.3005
R295 VTAIL.n121 VTAIL.n120 9.3005
R296 VTAIL.n119 VTAIL.n118 9.3005
R297 VTAIL.n88 VTAIL.n87 9.3005
R298 VTAIL.n113 VTAIL.n112 9.3005
R299 VTAIL.n111 VTAIL.n110 9.3005
R300 VTAIL.n92 VTAIL.n91 9.3005
R301 VTAIL.n105 VTAIL.n104 9.3005
R302 VTAIL.n103 VTAIL.n102 9.3005
R303 VTAIL.n96 VTAIL.n95 9.3005
R304 VTAIL.n250 VTAIL.n249 8.92171
R305 VTAIL.n265 VTAIL.n218 8.92171
R306 VTAIL.n40 VTAIL.n39 8.92171
R307 VTAIL.n55 VTAIL.n8 8.92171
R308 VTAIL.n199 VTAIL.n152 8.92171
R309 VTAIL.n184 VTAIL.n183 8.92171
R310 VTAIL.n129 VTAIL.n82 8.92171
R311 VTAIL.n114 VTAIL.n113 8.92171
R312 VTAIL.n253 VTAIL.n224 8.14595
R313 VTAIL.n262 VTAIL.n261 8.14595
R314 VTAIL.n43 VTAIL.n14 8.14595
R315 VTAIL.n52 VTAIL.n51 8.14595
R316 VTAIL.n196 VTAIL.n195 8.14595
R317 VTAIL.n187 VTAIL.n158 8.14595
R318 VTAIL.n126 VTAIL.n125 8.14595
R319 VTAIL.n117 VTAIL.n88 8.14595
R320 VTAIL.n254 VTAIL.n222 7.3702
R321 VTAIL.n258 VTAIL.n220 7.3702
R322 VTAIL.n44 VTAIL.n12 7.3702
R323 VTAIL.n48 VTAIL.n10 7.3702
R324 VTAIL.n192 VTAIL.n154 7.3702
R325 VTAIL.n188 VTAIL.n156 7.3702
R326 VTAIL.n122 VTAIL.n84 7.3702
R327 VTAIL.n118 VTAIL.n86 7.3702
R328 VTAIL.n257 VTAIL.n222 6.59444
R329 VTAIL.n258 VTAIL.n257 6.59444
R330 VTAIL.n47 VTAIL.n12 6.59444
R331 VTAIL.n48 VTAIL.n47 6.59444
R332 VTAIL.n192 VTAIL.n191 6.59444
R333 VTAIL.n191 VTAIL.n156 6.59444
R334 VTAIL.n122 VTAIL.n121 6.59444
R335 VTAIL.n121 VTAIL.n86 6.59444
R336 VTAIL.n254 VTAIL.n253 5.81868
R337 VTAIL.n261 VTAIL.n220 5.81868
R338 VTAIL.n44 VTAIL.n43 5.81868
R339 VTAIL.n51 VTAIL.n10 5.81868
R340 VTAIL.n195 VTAIL.n154 5.81868
R341 VTAIL.n188 VTAIL.n187 5.81868
R342 VTAIL.n125 VTAIL.n84 5.81868
R343 VTAIL.n118 VTAIL.n117 5.81868
R344 VTAIL.n250 VTAIL.n224 5.04292
R345 VTAIL.n262 VTAIL.n218 5.04292
R346 VTAIL.n40 VTAIL.n14 5.04292
R347 VTAIL.n52 VTAIL.n8 5.04292
R348 VTAIL.n196 VTAIL.n152 5.04292
R349 VTAIL.n184 VTAIL.n158 5.04292
R350 VTAIL.n126 VTAIL.n82 5.04292
R351 VTAIL.n114 VTAIL.n88 5.04292
R352 VTAIL.n249 VTAIL.n226 4.26717
R353 VTAIL.n266 VTAIL.n265 4.26717
R354 VTAIL.n39 VTAIL.n16 4.26717
R355 VTAIL.n56 VTAIL.n55 4.26717
R356 VTAIL.n200 VTAIL.n199 4.26717
R357 VTAIL.n183 VTAIL.n160 4.26717
R358 VTAIL.n130 VTAIL.n129 4.26717
R359 VTAIL.n113 VTAIL.n90 4.26717
R360 VTAIL.n167 VTAIL.n165 3.70982
R361 VTAIL.n97 VTAIL.n95 3.70982
R362 VTAIL.n233 VTAIL.n231 3.70982
R363 VTAIL.n23 VTAIL.n21 3.70982
R364 VTAIL.n246 VTAIL.n245 3.49141
R365 VTAIL.n269 VTAIL.n216 3.49141
R366 VTAIL.n36 VTAIL.n35 3.49141
R367 VTAIL.n59 VTAIL.n6 3.49141
R368 VTAIL.n203 VTAIL.n150 3.49141
R369 VTAIL.n180 VTAIL.n179 3.49141
R370 VTAIL.n133 VTAIL.n80 3.49141
R371 VTAIL.n110 VTAIL.n109 3.49141
R372 VTAIL.n278 VTAIL.t13 2.72514
R373 VTAIL.n278 VTAIL.t12 2.72514
R374 VTAIL.n0 VTAIL.t14 2.72514
R375 VTAIL.n0 VTAIL.t11 2.72514
R376 VTAIL.n68 VTAIL.t5 2.72514
R377 VTAIL.n68 VTAIL.t19 2.72514
R378 VTAIL.n70 VTAIL.t6 2.72514
R379 VTAIL.n70 VTAIL.t2 2.72514
R380 VTAIL.n144 VTAIL.t7 2.72514
R381 VTAIL.n144 VTAIL.t18 2.72514
R382 VTAIL.n142 VTAIL.t4 2.72514
R383 VTAIL.n142 VTAIL.t0 2.72514
R384 VTAIL.n74 VTAIL.t16 2.72514
R385 VTAIL.n74 VTAIL.t8 2.72514
R386 VTAIL.n72 VTAIL.t10 2.72514
R387 VTAIL.n72 VTAIL.t17 2.72514
R388 VTAIL.n242 VTAIL.n228 2.71565
R389 VTAIL.n270 VTAIL.n214 2.71565
R390 VTAIL.n32 VTAIL.n18 2.71565
R391 VTAIL.n60 VTAIL.n4 2.71565
R392 VTAIL.n204 VTAIL.n148 2.71565
R393 VTAIL.n176 VTAIL.n162 2.71565
R394 VTAIL.n134 VTAIL.n78 2.71565
R395 VTAIL.n106 VTAIL.n92 2.71565
R396 VTAIL.n241 VTAIL.n230 1.93989
R397 VTAIL.n274 VTAIL.n273 1.93989
R398 VTAIL.n31 VTAIL.n20 1.93989
R399 VTAIL.n64 VTAIL.n63 1.93989
R400 VTAIL.n208 VTAIL.n207 1.93989
R401 VTAIL.n175 VTAIL.n164 1.93989
R402 VTAIL.n138 VTAIL.n137 1.93989
R403 VTAIL.n105 VTAIL.n94 1.93989
R404 VTAIL.n238 VTAIL.n237 1.16414
R405 VTAIL.n276 VTAIL.n212 1.16414
R406 VTAIL.n28 VTAIL.n27 1.16414
R407 VTAIL.n66 VTAIL.n2 1.16414
R408 VTAIL.n210 VTAIL.n146 1.16414
R409 VTAIL.n172 VTAIL.n171 1.16414
R410 VTAIL.n140 VTAIL.n76 1.16414
R411 VTAIL.n102 VTAIL.n101 1.16414
R412 VTAIL.n143 VTAIL.n141 0.901362
R413 VTAIL.n67 VTAIL.n1 0.901362
R414 VTAIL.n75 VTAIL.n73 0.862569
R415 VTAIL.n141 VTAIL.n75 0.862569
R416 VTAIL.n145 VTAIL.n143 0.862569
R417 VTAIL.n211 VTAIL.n145 0.862569
R418 VTAIL.n71 VTAIL.n69 0.862569
R419 VTAIL.n69 VTAIL.n67 0.862569
R420 VTAIL.n279 VTAIL.n277 0.862569
R421 VTAIL VTAIL.n1 0.705241
R422 VTAIL.n234 VTAIL.n232 0.388379
R423 VTAIL.n24 VTAIL.n22 0.388379
R424 VTAIL.n168 VTAIL.n166 0.388379
R425 VTAIL.n98 VTAIL.n96 0.388379
R426 VTAIL VTAIL.n279 0.157828
R427 VTAIL.n239 VTAIL.n231 0.155672
R428 VTAIL.n240 VTAIL.n239 0.155672
R429 VTAIL.n240 VTAIL.n227 0.155672
R430 VTAIL.n247 VTAIL.n227 0.155672
R431 VTAIL.n248 VTAIL.n247 0.155672
R432 VTAIL.n248 VTAIL.n223 0.155672
R433 VTAIL.n255 VTAIL.n223 0.155672
R434 VTAIL.n256 VTAIL.n255 0.155672
R435 VTAIL.n256 VTAIL.n219 0.155672
R436 VTAIL.n263 VTAIL.n219 0.155672
R437 VTAIL.n264 VTAIL.n263 0.155672
R438 VTAIL.n264 VTAIL.n215 0.155672
R439 VTAIL.n271 VTAIL.n215 0.155672
R440 VTAIL.n272 VTAIL.n271 0.155672
R441 VTAIL.n29 VTAIL.n21 0.155672
R442 VTAIL.n30 VTAIL.n29 0.155672
R443 VTAIL.n30 VTAIL.n17 0.155672
R444 VTAIL.n37 VTAIL.n17 0.155672
R445 VTAIL.n38 VTAIL.n37 0.155672
R446 VTAIL.n38 VTAIL.n13 0.155672
R447 VTAIL.n45 VTAIL.n13 0.155672
R448 VTAIL.n46 VTAIL.n45 0.155672
R449 VTAIL.n46 VTAIL.n9 0.155672
R450 VTAIL.n53 VTAIL.n9 0.155672
R451 VTAIL.n54 VTAIL.n53 0.155672
R452 VTAIL.n54 VTAIL.n5 0.155672
R453 VTAIL.n61 VTAIL.n5 0.155672
R454 VTAIL.n62 VTAIL.n61 0.155672
R455 VTAIL.n206 VTAIL.n205 0.155672
R456 VTAIL.n205 VTAIL.n149 0.155672
R457 VTAIL.n198 VTAIL.n149 0.155672
R458 VTAIL.n198 VTAIL.n197 0.155672
R459 VTAIL.n197 VTAIL.n153 0.155672
R460 VTAIL.n190 VTAIL.n153 0.155672
R461 VTAIL.n190 VTAIL.n189 0.155672
R462 VTAIL.n189 VTAIL.n157 0.155672
R463 VTAIL.n182 VTAIL.n157 0.155672
R464 VTAIL.n182 VTAIL.n181 0.155672
R465 VTAIL.n181 VTAIL.n161 0.155672
R466 VTAIL.n174 VTAIL.n161 0.155672
R467 VTAIL.n174 VTAIL.n173 0.155672
R468 VTAIL.n173 VTAIL.n165 0.155672
R469 VTAIL.n136 VTAIL.n135 0.155672
R470 VTAIL.n135 VTAIL.n79 0.155672
R471 VTAIL.n128 VTAIL.n79 0.155672
R472 VTAIL.n128 VTAIL.n127 0.155672
R473 VTAIL.n127 VTAIL.n83 0.155672
R474 VTAIL.n120 VTAIL.n83 0.155672
R475 VTAIL.n120 VTAIL.n119 0.155672
R476 VTAIL.n119 VTAIL.n87 0.155672
R477 VTAIL.n112 VTAIL.n87 0.155672
R478 VTAIL.n112 VTAIL.n111 0.155672
R479 VTAIL.n111 VTAIL.n91 0.155672
R480 VTAIL.n104 VTAIL.n91 0.155672
R481 VTAIL.n104 VTAIL.n103 0.155672
R482 VTAIL.n103 VTAIL.n95 0.155672
R483 VDD2.n133 VDD2.n132 756.745
R484 VDD2.n64 VDD2.n63 756.745
R485 VDD2.n132 VDD2.n131 585
R486 VDD2.n71 VDD2.n70 585
R487 VDD2.n126 VDD2.n125 585
R488 VDD2.n124 VDD2.n123 585
R489 VDD2.n75 VDD2.n74 585
R490 VDD2.n118 VDD2.n117 585
R491 VDD2.n116 VDD2.n115 585
R492 VDD2.n79 VDD2.n78 585
R493 VDD2.n110 VDD2.n109 585
R494 VDD2.n108 VDD2.n107 585
R495 VDD2.n83 VDD2.n82 585
R496 VDD2.n102 VDD2.n101 585
R497 VDD2.n100 VDD2.n99 585
R498 VDD2.n87 VDD2.n86 585
R499 VDD2.n94 VDD2.n93 585
R500 VDD2.n92 VDD2.n91 585
R501 VDD2.n23 VDD2.n22 585
R502 VDD2.n25 VDD2.n24 585
R503 VDD2.n18 VDD2.n17 585
R504 VDD2.n31 VDD2.n30 585
R505 VDD2.n33 VDD2.n32 585
R506 VDD2.n14 VDD2.n13 585
R507 VDD2.n39 VDD2.n38 585
R508 VDD2.n41 VDD2.n40 585
R509 VDD2.n10 VDD2.n9 585
R510 VDD2.n47 VDD2.n46 585
R511 VDD2.n49 VDD2.n48 585
R512 VDD2.n6 VDD2.n5 585
R513 VDD2.n55 VDD2.n54 585
R514 VDD2.n57 VDD2.n56 585
R515 VDD2.n2 VDD2.n1 585
R516 VDD2.n63 VDD2.n62 585
R517 VDD2.n90 VDD2.t9 327.466
R518 VDD2.n21 VDD2.t0 327.466
R519 VDD2.n132 VDD2.n70 171.744
R520 VDD2.n125 VDD2.n70 171.744
R521 VDD2.n125 VDD2.n124 171.744
R522 VDD2.n124 VDD2.n74 171.744
R523 VDD2.n117 VDD2.n74 171.744
R524 VDD2.n117 VDD2.n116 171.744
R525 VDD2.n116 VDD2.n78 171.744
R526 VDD2.n109 VDD2.n78 171.744
R527 VDD2.n109 VDD2.n108 171.744
R528 VDD2.n108 VDD2.n82 171.744
R529 VDD2.n101 VDD2.n82 171.744
R530 VDD2.n101 VDD2.n100 171.744
R531 VDD2.n100 VDD2.n86 171.744
R532 VDD2.n93 VDD2.n86 171.744
R533 VDD2.n93 VDD2.n92 171.744
R534 VDD2.n24 VDD2.n23 171.744
R535 VDD2.n24 VDD2.n17 171.744
R536 VDD2.n31 VDD2.n17 171.744
R537 VDD2.n32 VDD2.n31 171.744
R538 VDD2.n32 VDD2.n13 171.744
R539 VDD2.n39 VDD2.n13 171.744
R540 VDD2.n40 VDD2.n39 171.744
R541 VDD2.n40 VDD2.n9 171.744
R542 VDD2.n47 VDD2.n9 171.744
R543 VDD2.n48 VDD2.n47 171.744
R544 VDD2.n48 VDD2.n5 171.744
R545 VDD2.n55 VDD2.n5 171.744
R546 VDD2.n56 VDD2.n55 171.744
R547 VDD2.n56 VDD2.n1 171.744
R548 VDD2.n63 VDD2.n1 171.744
R549 VDD2.n92 VDD2.t9 85.8723
R550 VDD2.n23 VDD2.t0 85.8723
R551 VDD2.n68 VDD2.n67 77.3039
R552 VDD2 VDD2.n137 77.3002
R553 VDD2.n136 VDD2.n135 76.7129
R554 VDD2.n66 VDD2.n65 76.7127
R555 VDD2.n66 VDD2.n64 51.8595
R556 VDD2.n134 VDD2.n133 50.9975
R557 VDD2.n134 VDD2.n68 38.0946
R558 VDD2.n91 VDD2.n90 16.3895
R559 VDD2.n22 VDD2.n21 16.3895
R560 VDD2.n94 VDD2.n89 12.8005
R561 VDD2.n25 VDD2.n20 12.8005
R562 VDD2.n131 VDD2.n69 12.0247
R563 VDD2.n95 VDD2.n87 12.0247
R564 VDD2.n26 VDD2.n18 12.0247
R565 VDD2.n62 VDD2.n0 12.0247
R566 VDD2.n130 VDD2.n71 11.249
R567 VDD2.n99 VDD2.n98 11.249
R568 VDD2.n30 VDD2.n29 11.249
R569 VDD2.n61 VDD2.n2 11.249
R570 VDD2.n127 VDD2.n126 10.4732
R571 VDD2.n102 VDD2.n85 10.4732
R572 VDD2.n33 VDD2.n16 10.4732
R573 VDD2.n58 VDD2.n57 10.4732
R574 VDD2.n123 VDD2.n73 9.69747
R575 VDD2.n103 VDD2.n83 9.69747
R576 VDD2.n34 VDD2.n14 9.69747
R577 VDD2.n54 VDD2.n4 9.69747
R578 VDD2.n129 VDD2.n69 9.45567
R579 VDD2.n60 VDD2.n0 9.45567
R580 VDD2.n77 VDD2.n76 9.3005
R581 VDD2.n120 VDD2.n119 9.3005
R582 VDD2.n122 VDD2.n121 9.3005
R583 VDD2.n73 VDD2.n72 9.3005
R584 VDD2.n128 VDD2.n127 9.3005
R585 VDD2.n130 VDD2.n129 9.3005
R586 VDD2.n114 VDD2.n113 9.3005
R587 VDD2.n112 VDD2.n111 9.3005
R588 VDD2.n81 VDD2.n80 9.3005
R589 VDD2.n106 VDD2.n105 9.3005
R590 VDD2.n104 VDD2.n103 9.3005
R591 VDD2.n85 VDD2.n84 9.3005
R592 VDD2.n98 VDD2.n97 9.3005
R593 VDD2.n96 VDD2.n95 9.3005
R594 VDD2.n89 VDD2.n88 9.3005
R595 VDD2.n45 VDD2.n44 9.3005
R596 VDD2.n8 VDD2.n7 9.3005
R597 VDD2.n51 VDD2.n50 9.3005
R598 VDD2.n53 VDD2.n52 9.3005
R599 VDD2.n4 VDD2.n3 9.3005
R600 VDD2.n59 VDD2.n58 9.3005
R601 VDD2.n61 VDD2.n60 9.3005
R602 VDD2.n12 VDD2.n11 9.3005
R603 VDD2.n37 VDD2.n36 9.3005
R604 VDD2.n35 VDD2.n34 9.3005
R605 VDD2.n16 VDD2.n15 9.3005
R606 VDD2.n29 VDD2.n28 9.3005
R607 VDD2.n27 VDD2.n26 9.3005
R608 VDD2.n20 VDD2.n19 9.3005
R609 VDD2.n43 VDD2.n42 9.3005
R610 VDD2.n122 VDD2.n75 8.92171
R611 VDD2.n107 VDD2.n106 8.92171
R612 VDD2.n38 VDD2.n37 8.92171
R613 VDD2.n53 VDD2.n6 8.92171
R614 VDD2.n119 VDD2.n118 8.14595
R615 VDD2.n110 VDD2.n81 8.14595
R616 VDD2.n41 VDD2.n12 8.14595
R617 VDD2.n50 VDD2.n49 8.14595
R618 VDD2.n115 VDD2.n77 7.3702
R619 VDD2.n111 VDD2.n79 7.3702
R620 VDD2.n42 VDD2.n10 7.3702
R621 VDD2.n46 VDD2.n8 7.3702
R622 VDD2.n115 VDD2.n114 6.59444
R623 VDD2.n114 VDD2.n79 6.59444
R624 VDD2.n45 VDD2.n10 6.59444
R625 VDD2.n46 VDD2.n45 6.59444
R626 VDD2.n118 VDD2.n77 5.81868
R627 VDD2.n111 VDD2.n110 5.81868
R628 VDD2.n42 VDD2.n41 5.81868
R629 VDD2.n49 VDD2.n8 5.81868
R630 VDD2.n119 VDD2.n75 5.04292
R631 VDD2.n107 VDD2.n81 5.04292
R632 VDD2.n38 VDD2.n12 5.04292
R633 VDD2.n50 VDD2.n6 5.04292
R634 VDD2.n123 VDD2.n122 4.26717
R635 VDD2.n106 VDD2.n83 4.26717
R636 VDD2.n37 VDD2.n14 4.26717
R637 VDD2.n54 VDD2.n53 4.26717
R638 VDD2.n90 VDD2.n88 3.70982
R639 VDD2.n21 VDD2.n19 3.70982
R640 VDD2.n126 VDD2.n73 3.49141
R641 VDD2.n103 VDD2.n102 3.49141
R642 VDD2.n34 VDD2.n33 3.49141
R643 VDD2.n57 VDD2.n4 3.49141
R644 VDD2.n137 VDD2.t1 2.72514
R645 VDD2.n137 VDD2.t5 2.72514
R646 VDD2.n135 VDD2.t3 2.72514
R647 VDD2.n135 VDD2.t7 2.72514
R648 VDD2.n67 VDD2.t6 2.72514
R649 VDD2.n67 VDD2.t8 2.72514
R650 VDD2.n65 VDD2.t2 2.72514
R651 VDD2.n65 VDD2.t4 2.72514
R652 VDD2.n127 VDD2.n71 2.71565
R653 VDD2.n99 VDD2.n85 2.71565
R654 VDD2.n30 VDD2.n16 2.71565
R655 VDD2.n58 VDD2.n2 2.71565
R656 VDD2.n131 VDD2.n130 1.93989
R657 VDD2.n98 VDD2.n87 1.93989
R658 VDD2.n29 VDD2.n18 1.93989
R659 VDD2.n62 VDD2.n61 1.93989
R660 VDD2.n133 VDD2.n69 1.16414
R661 VDD2.n95 VDD2.n94 1.16414
R662 VDD2.n26 VDD2.n25 1.16414
R663 VDD2.n64 VDD2.n0 1.16414
R664 VDD2.n136 VDD2.n134 0.862569
R665 VDD2.n91 VDD2.n89 0.388379
R666 VDD2.n22 VDD2.n20 0.388379
R667 VDD2 VDD2.n136 0.274207
R668 VDD2.n68 VDD2.n66 0.160671
R669 VDD2.n129 VDD2.n128 0.155672
R670 VDD2.n128 VDD2.n72 0.155672
R671 VDD2.n121 VDD2.n72 0.155672
R672 VDD2.n121 VDD2.n120 0.155672
R673 VDD2.n120 VDD2.n76 0.155672
R674 VDD2.n113 VDD2.n76 0.155672
R675 VDD2.n113 VDD2.n112 0.155672
R676 VDD2.n112 VDD2.n80 0.155672
R677 VDD2.n105 VDD2.n80 0.155672
R678 VDD2.n105 VDD2.n104 0.155672
R679 VDD2.n104 VDD2.n84 0.155672
R680 VDD2.n97 VDD2.n84 0.155672
R681 VDD2.n97 VDD2.n96 0.155672
R682 VDD2.n96 VDD2.n88 0.155672
R683 VDD2.n27 VDD2.n19 0.155672
R684 VDD2.n28 VDD2.n27 0.155672
R685 VDD2.n28 VDD2.n15 0.155672
R686 VDD2.n35 VDD2.n15 0.155672
R687 VDD2.n36 VDD2.n35 0.155672
R688 VDD2.n36 VDD2.n11 0.155672
R689 VDD2.n43 VDD2.n11 0.155672
R690 VDD2.n44 VDD2.n43 0.155672
R691 VDD2.n44 VDD2.n7 0.155672
R692 VDD2.n51 VDD2.n7 0.155672
R693 VDD2.n52 VDD2.n51 0.155672
R694 VDD2.n52 VDD2.n3 0.155672
R695 VDD2.n59 VDD2.n3 0.155672
R696 VDD2.n60 VDD2.n59 0.155672
R697 B.n247 B.t6 632.475
R698 B.n112 B.t0 632.475
R699 B.n42 B.t3 632.475
R700 B.n36 B.t9 632.475
R701 B.n328 B.n91 585
R702 B.n327 B.n326 585
R703 B.n325 B.n92 585
R704 B.n324 B.n323 585
R705 B.n322 B.n93 585
R706 B.n321 B.n320 585
R707 B.n319 B.n94 585
R708 B.n318 B.n317 585
R709 B.n316 B.n95 585
R710 B.n315 B.n314 585
R711 B.n313 B.n96 585
R712 B.n312 B.n311 585
R713 B.n310 B.n97 585
R714 B.n309 B.n308 585
R715 B.n307 B.n98 585
R716 B.n306 B.n305 585
R717 B.n304 B.n99 585
R718 B.n303 B.n302 585
R719 B.n301 B.n100 585
R720 B.n300 B.n299 585
R721 B.n298 B.n101 585
R722 B.n297 B.n296 585
R723 B.n295 B.n102 585
R724 B.n294 B.n293 585
R725 B.n292 B.n103 585
R726 B.n291 B.n290 585
R727 B.n289 B.n104 585
R728 B.n288 B.n287 585
R729 B.n286 B.n105 585
R730 B.n285 B.n284 585
R731 B.n283 B.n106 585
R732 B.n282 B.n281 585
R733 B.n280 B.n107 585
R734 B.n279 B.n278 585
R735 B.n277 B.n108 585
R736 B.n276 B.n275 585
R737 B.n274 B.n109 585
R738 B.n273 B.n272 585
R739 B.n271 B.n110 585
R740 B.n270 B.n269 585
R741 B.n268 B.n111 585
R742 B.n266 B.n265 585
R743 B.n264 B.n114 585
R744 B.n263 B.n262 585
R745 B.n261 B.n115 585
R746 B.n260 B.n259 585
R747 B.n258 B.n116 585
R748 B.n257 B.n256 585
R749 B.n255 B.n117 585
R750 B.n254 B.n253 585
R751 B.n252 B.n118 585
R752 B.n251 B.n250 585
R753 B.n246 B.n119 585
R754 B.n245 B.n244 585
R755 B.n243 B.n120 585
R756 B.n242 B.n241 585
R757 B.n240 B.n121 585
R758 B.n239 B.n238 585
R759 B.n237 B.n122 585
R760 B.n236 B.n235 585
R761 B.n234 B.n123 585
R762 B.n233 B.n232 585
R763 B.n231 B.n124 585
R764 B.n230 B.n229 585
R765 B.n228 B.n125 585
R766 B.n227 B.n226 585
R767 B.n225 B.n126 585
R768 B.n224 B.n223 585
R769 B.n222 B.n127 585
R770 B.n221 B.n220 585
R771 B.n219 B.n128 585
R772 B.n218 B.n217 585
R773 B.n216 B.n129 585
R774 B.n215 B.n214 585
R775 B.n213 B.n130 585
R776 B.n212 B.n211 585
R777 B.n210 B.n131 585
R778 B.n209 B.n208 585
R779 B.n207 B.n132 585
R780 B.n206 B.n205 585
R781 B.n204 B.n133 585
R782 B.n203 B.n202 585
R783 B.n201 B.n134 585
R784 B.n200 B.n199 585
R785 B.n198 B.n135 585
R786 B.n197 B.n196 585
R787 B.n195 B.n136 585
R788 B.n194 B.n193 585
R789 B.n192 B.n137 585
R790 B.n191 B.n190 585
R791 B.n189 B.n138 585
R792 B.n188 B.n187 585
R793 B.n330 B.n329 585
R794 B.n331 B.n90 585
R795 B.n333 B.n332 585
R796 B.n334 B.n89 585
R797 B.n336 B.n335 585
R798 B.n337 B.n88 585
R799 B.n339 B.n338 585
R800 B.n340 B.n87 585
R801 B.n342 B.n341 585
R802 B.n343 B.n86 585
R803 B.n345 B.n344 585
R804 B.n346 B.n85 585
R805 B.n348 B.n347 585
R806 B.n349 B.n84 585
R807 B.n351 B.n350 585
R808 B.n352 B.n83 585
R809 B.n354 B.n353 585
R810 B.n355 B.n82 585
R811 B.n357 B.n356 585
R812 B.n358 B.n81 585
R813 B.n360 B.n359 585
R814 B.n361 B.n80 585
R815 B.n363 B.n362 585
R816 B.n364 B.n79 585
R817 B.n366 B.n365 585
R818 B.n367 B.n78 585
R819 B.n369 B.n368 585
R820 B.n370 B.n77 585
R821 B.n372 B.n371 585
R822 B.n373 B.n76 585
R823 B.n375 B.n374 585
R824 B.n376 B.n75 585
R825 B.n378 B.n377 585
R826 B.n379 B.n74 585
R827 B.n381 B.n380 585
R828 B.n382 B.n73 585
R829 B.n384 B.n383 585
R830 B.n385 B.n72 585
R831 B.n387 B.n386 585
R832 B.n388 B.n71 585
R833 B.n390 B.n389 585
R834 B.n391 B.n70 585
R835 B.n393 B.n392 585
R836 B.n394 B.n69 585
R837 B.n396 B.n395 585
R838 B.n397 B.n68 585
R839 B.n399 B.n398 585
R840 B.n400 B.n67 585
R841 B.n402 B.n401 585
R842 B.n403 B.n66 585
R843 B.n405 B.n404 585
R844 B.n406 B.n65 585
R845 B.n546 B.n545 585
R846 B.n544 B.n15 585
R847 B.n543 B.n542 585
R848 B.n541 B.n16 585
R849 B.n540 B.n539 585
R850 B.n538 B.n17 585
R851 B.n537 B.n536 585
R852 B.n535 B.n18 585
R853 B.n534 B.n533 585
R854 B.n532 B.n19 585
R855 B.n531 B.n530 585
R856 B.n529 B.n20 585
R857 B.n528 B.n527 585
R858 B.n526 B.n21 585
R859 B.n525 B.n524 585
R860 B.n523 B.n22 585
R861 B.n522 B.n521 585
R862 B.n520 B.n23 585
R863 B.n519 B.n518 585
R864 B.n517 B.n24 585
R865 B.n516 B.n515 585
R866 B.n514 B.n25 585
R867 B.n513 B.n512 585
R868 B.n511 B.n26 585
R869 B.n510 B.n509 585
R870 B.n508 B.n27 585
R871 B.n507 B.n506 585
R872 B.n505 B.n28 585
R873 B.n504 B.n503 585
R874 B.n502 B.n29 585
R875 B.n501 B.n500 585
R876 B.n499 B.n30 585
R877 B.n498 B.n497 585
R878 B.n496 B.n31 585
R879 B.n495 B.n494 585
R880 B.n493 B.n32 585
R881 B.n492 B.n491 585
R882 B.n490 B.n33 585
R883 B.n489 B.n488 585
R884 B.n487 B.n34 585
R885 B.n486 B.n485 585
R886 B.n483 B.n35 585
R887 B.n482 B.n481 585
R888 B.n480 B.n38 585
R889 B.n479 B.n478 585
R890 B.n477 B.n39 585
R891 B.n476 B.n475 585
R892 B.n474 B.n40 585
R893 B.n473 B.n472 585
R894 B.n471 B.n41 585
R895 B.n470 B.n469 585
R896 B.n468 B.n467 585
R897 B.n466 B.n45 585
R898 B.n465 B.n464 585
R899 B.n463 B.n46 585
R900 B.n462 B.n461 585
R901 B.n460 B.n47 585
R902 B.n459 B.n458 585
R903 B.n457 B.n48 585
R904 B.n456 B.n455 585
R905 B.n454 B.n49 585
R906 B.n453 B.n452 585
R907 B.n451 B.n50 585
R908 B.n450 B.n449 585
R909 B.n448 B.n51 585
R910 B.n447 B.n446 585
R911 B.n445 B.n52 585
R912 B.n444 B.n443 585
R913 B.n442 B.n53 585
R914 B.n441 B.n440 585
R915 B.n439 B.n54 585
R916 B.n438 B.n437 585
R917 B.n436 B.n55 585
R918 B.n435 B.n434 585
R919 B.n433 B.n56 585
R920 B.n432 B.n431 585
R921 B.n430 B.n57 585
R922 B.n429 B.n428 585
R923 B.n427 B.n58 585
R924 B.n426 B.n425 585
R925 B.n424 B.n59 585
R926 B.n423 B.n422 585
R927 B.n421 B.n60 585
R928 B.n420 B.n419 585
R929 B.n418 B.n61 585
R930 B.n417 B.n416 585
R931 B.n415 B.n62 585
R932 B.n414 B.n413 585
R933 B.n412 B.n63 585
R934 B.n411 B.n410 585
R935 B.n409 B.n64 585
R936 B.n408 B.n407 585
R937 B.n547 B.n14 585
R938 B.n549 B.n548 585
R939 B.n550 B.n13 585
R940 B.n552 B.n551 585
R941 B.n553 B.n12 585
R942 B.n555 B.n554 585
R943 B.n556 B.n11 585
R944 B.n558 B.n557 585
R945 B.n559 B.n10 585
R946 B.n561 B.n560 585
R947 B.n562 B.n9 585
R948 B.n564 B.n563 585
R949 B.n565 B.n8 585
R950 B.n567 B.n566 585
R951 B.n568 B.n7 585
R952 B.n570 B.n569 585
R953 B.n571 B.n6 585
R954 B.n573 B.n572 585
R955 B.n574 B.n5 585
R956 B.n576 B.n575 585
R957 B.n577 B.n4 585
R958 B.n579 B.n578 585
R959 B.n580 B.n3 585
R960 B.n582 B.n581 585
R961 B.n583 B.n0 585
R962 B.n2 B.n1 585
R963 B.n152 B.n151 585
R964 B.n153 B.n150 585
R965 B.n155 B.n154 585
R966 B.n156 B.n149 585
R967 B.n158 B.n157 585
R968 B.n159 B.n148 585
R969 B.n161 B.n160 585
R970 B.n162 B.n147 585
R971 B.n164 B.n163 585
R972 B.n165 B.n146 585
R973 B.n167 B.n166 585
R974 B.n168 B.n145 585
R975 B.n170 B.n169 585
R976 B.n171 B.n144 585
R977 B.n173 B.n172 585
R978 B.n174 B.n143 585
R979 B.n176 B.n175 585
R980 B.n177 B.n142 585
R981 B.n179 B.n178 585
R982 B.n180 B.n141 585
R983 B.n182 B.n181 585
R984 B.n183 B.n140 585
R985 B.n185 B.n184 585
R986 B.n186 B.n139 585
R987 B.n188 B.n139 574.183
R988 B.n330 B.n91 574.183
R989 B.n408 B.n65 574.183
R990 B.n547 B.n546 574.183
R991 B.n112 B.t1 393.567
R992 B.n42 B.t5 393.567
R993 B.n247 B.t7 393.567
R994 B.n36 B.t11 393.567
R995 B.n113 B.t2 374.173
R996 B.n43 B.t4 374.173
R997 B.n248 B.t8 374.173
R998 B.n37 B.t10 374.173
R999 B.n585 B.n584 256.663
R1000 B.n584 B.n583 235.042
R1001 B.n584 B.n2 235.042
R1002 B.n189 B.n188 163.367
R1003 B.n190 B.n189 163.367
R1004 B.n190 B.n137 163.367
R1005 B.n194 B.n137 163.367
R1006 B.n195 B.n194 163.367
R1007 B.n196 B.n195 163.367
R1008 B.n196 B.n135 163.367
R1009 B.n200 B.n135 163.367
R1010 B.n201 B.n200 163.367
R1011 B.n202 B.n201 163.367
R1012 B.n202 B.n133 163.367
R1013 B.n206 B.n133 163.367
R1014 B.n207 B.n206 163.367
R1015 B.n208 B.n207 163.367
R1016 B.n208 B.n131 163.367
R1017 B.n212 B.n131 163.367
R1018 B.n213 B.n212 163.367
R1019 B.n214 B.n213 163.367
R1020 B.n214 B.n129 163.367
R1021 B.n218 B.n129 163.367
R1022 B.n219 B.n218 163.367
R1023 B.n220 B.n219 163.367
R1024 B.n220 B.n127 163.367
R1025 B.n224 B.n127 163.367
R1026 B.n225 B.n224 163.367
R1027 B.n226 B.n225 163.367
R1028 B.n226 B.n125 163.367
R1029 B.n230 B.n125 163.367
R1030 B.n231 B.n230 163.367
R1031 B.n232 B.n231 163.367
R1032 B.n232 B.n123 163.367
R1033 B.n236 B.n123 163.367
R1034 B.n237 B.n236 163.367
R1035 B.n238 B.n237 163.367
R1036 B.n238 B.n121 163.367
R1037 B.n242 B.n121 163.367
R1038 B.n243 B.n242 163.367
R1039 B.n244 B.n243 163.367
R1040 B.n244 B.n119 163.367
R1041 B.n251 B.n119 163.367
R1042 B.n252 B.n251 163.367
R1043 B.n253 B.n252 163.367
R1044 B.n253 B.n117 163.367
R1045 B.n257 B.n117 163.367
R1046 B.n258 B.n257 163.367
R1047 B.n259 B.n258 163.367
R1048 B.n259 B.n115 163.367
R1049 B.n263 B.n115 163.367
R1050 B.n264 B.n263 163.367
R1051 B.n265 B.n264 163.367
R1052 B.n265 B.n111 163.367
R1053 B.n270 B.n111 163.367
R1054 B.n271 B.n270 163.367
R1055 B.n272 B.n271 163.367
R1056 B.n272 B.n109 163.367
R1057 B.n276 B.n109 163.367
R1058 B.n277 B.n276 163.367
R1059 B.n278 B.n277 163.367
R1060 B.n278 B.n107 163.367
R1061 B.n282 B.n107 163.367
R1062 B.n283 B.n282 163.367
R1063 B.n284 B.n283 163.367
R1064 B.n284 B.n105 163.367
R1065 B.n288 B.n105 163.367
R1066 B.n289 B.n288 163.367
R1067 B.n290 B.n289 163.367
R1068 B.n290 B.n103 163.367
R1069 B.n294 B.n103 163.367
R1070 B.n295 B.n294 163.367
R1071 B.n296 B.n295 163.367
R1072 B.n296 B.n101 163.367
R1073 B.n300 B.n101 163.367
R1074 B.n301 B.n300 163.367
R1075 B.n302 B.n301 163.367
R1076 B.n302 B.n99 163.367
R1077 B.n306 B.n99 163.367
R1078 B.n307 B.n306 163.367
R1079 B.n308 B.n307 163.367
R1080 B.n308 B.n97 163.367
R1081 B.n312 B.n97 163.367
R1082 B.n313 B.n312 163.367
R1083 B.n314 B.n313 163.367
R1084 B.n314 B.n95 163.367
R1085 B.n318 B.n95 163.367
R1086 B.n319 B.n318 163.367
R1087 B.n320 B.n319 163.367
R1088 B.n320 B.n93 163.367
R1089 B.n324 B.n93 163.367
R1090 B.n325 B.n324 163.367
R1091 B.n326 B.n325 163.367
R1092 B.n326 B.n91 163.367
R1093 B.n404 B.n65 163.367
R1094 B.n404 B.n403 163.367
R1095 B.n403 B.n402 163.367
R1096 B.n402 B.n67 163.367
R1097 B.n398 B.n67 163.367
R1098 B.n398 B.n397 163.367
R1099 B.n397 B.n396 163.367
R1100 B.n396 B.n69 163.367
R1101 B.n392 B.n69 163.367
R1102 B.n392 B.n391 163.367
R1103 B.n391 B.n390 163.367
R1104 B.n390 B.n71 163.367
R1105 B.n386 B.n71 163.367
R1106 B.n386 B.n385 163.367
R1107 B.n385 B.n384 163.367
R1108 B.n384 B.n73 163.367
R1109 B.n380 B.n73 163.367
R1110 B.n380 B.n379 163.367
R1111 B.n379 B.n378 163.367
R1112 B.n378 B.n75 163.367
R1113 B.n374 B.n75 163.367
R1114 B.n374 B.n373 163.367
R1115 B.n373 B.n372 163.367
R1116 B.n372 B.n77 163.367
R1117 B.n368 B.n77 163.367
R1118 B.n368 B.n367 163.367
R1119 B.n367 B.n366 163.367
R1120 B.n366 B.n79 163.367
R1121 B.n362 B.n79 163.367
R1122 B.n362 B.n361 163.367
R1123 B.n361 B.n360 163.367
R1124 B.n360 B.n81 163.367
R1125 B.n356 B.n81 163.367
R1126 B.n356 B.n355 163.367
R1127 B.n355 B.n354 163.367
R1128 B.n354 B.n83 163.367
R1129 B.n350 B.n83 163.367
R1130 B.n350 B.n349 163.367
R1131 B.n349 B.n348 163.367
R1132 B.n348 B.n85 163.367
R1133 B.n344 B.n85 163.367
R1134 B.n344 B.n343 163.367
R1135 B.n343 B.n342 163.367
R1136 B.n342 B.n87 163.367
R1137 B.n338 B.n87 163.367
R1138 B.n338 B.n337 163.367
R1139 B.n337 B.n336 163.367
R1140 B.n336 B.n89 163.367
R1141 B.n332 B.n89 163.367
R1142 B.n332 B.n331 163.367
R1143 B.n331 B.n330 163.367
R1144 B.n546 B.n15 163.367
R1145 B.n542 B.n15 163.367
R1146 B.n542 B.n541 163.367
R1147 B.n541 B.n540 163.367
R1148 B.n540 B.n17 163.367
R1149 B.n536 B.n17 163.367
R1150 B.n536 B.n535 163.367
R1151 B.n535 B.n534 163.367
R1152 B.n534 B.n19 163.367
R1153 B.n530 B.n19 163.367
R1154 B.n530 B.n529 163.367
R1155 B.n529 B.n528 163.367
R1156 B.n528 B.n21 163.367
R1157 B.n524 B.n21 163.367
R1158 B.n524 B.n523 163.367
R1159 B.n523 B.n522 163.367
R1160 B.n522 B.n23 163.367
R1161 B.n518 B.n23 163.367
R1162 B.n518 B.n517 163.367
R1163 B.n517 B.n516 163.367
R1164 B.n516 B.n25 163.367
R1165 B.n512 B.n25 163.367
R1166 B.n512 B.n511 163.367
R1167 B.n511 B.n510 163.367
R1168 B.n510 B.n27 163.367
R1169 B.n506 B.n27 163.367
R1170 B.n506 B.n505 163.367
R1171 B.n505 B.n504 163.367
R1172 B.n504 B.n29 163.367
R1173 B.n500 B.n29 163.367
R1174 B.n500 B.n499 163.367
R1175 B.n499 B.n498 163.367
R1176 B.n498 B.n31 163.367
R1177 B.n494 B.n31 163.367
R1178 B.n494 B.n493 163.367
R1179 B.n493 B.n492 163.367
R1180 B.n492 B.n33 163.367
R1181 B.n488 B.n33 163.367
R1182 B.n488 B.n487 163.367
R1183 B.n487 B.n486 163.367
R1184 B.n486 B.n35 163.367
R1185 B.n481 B.n35 163.367
R1186 B.n481 B.n480 163.367
R1187 B.n480 B.n479 163.367
R1188 B.n479 B.n39 163.367
R1189 B.n475 B.n39 163.367
R1190 B.n475 B.n474 163.367
R1191 B.n474 B.n473 163.367
R1192 B.n473 B.n41 163.367
R1193 B.n469 B.n41 163.367
R1194 B.n469 B.n468 163.367
R1195 B.n468 B.n45 163.367
R1196 B.n464 B.n45 163.367
R1197 B.n464 B.n463 163.367
R1198 B.n463 B.n462 163.367
R1199 B.n462 B.n47 163.367
R1200 B.n458 B.n47 163.367
R1201 B.n458 B.n457 163.367
R1202 B.n457 B.n456 163.367
R1203 B.n456 B.n49 163.367
R1204 B.n452 B.n49 163.367
R1205 B.n452 B.n451 163.367
R1206 B.n451 B.n450 163.367
R1207 B.n450 B.n51 163.367
R1208 B.n446 B.n51 163.367
R1209 B.n446 B.n445 163.367
R1210 B.n445 B.n444 163.367
R1211 B.n444 B.n53 163.367
R1212 B.n440 B.n53 163.367
R1213 B.n440 B.n439 163.367
R1214 B.n439 B.n438 163.367
R1215 B.n438 B.n55 163.367
R1216 B.n434 B.n55 163.367
R1217 B.n434 B.n433 163.367
R1218 B.n433 B.n432 163.367
R1219 B.n432 B.n57 163.367
R1220 B.n428 B.n57 163.367
R1221 B.n428 B.n427 163.367
R1222 B.n427 B.n426 163.367
R1223 B.n426 B.n59 163.367
R1224 B.n422 B.n59 163.367
R1225 B.n422 B.n421 163.367
R1226 B.n421 B.n420 163.367
R1227 B.n420 B.n61 163.367
R1228 B.n416 B.n61 163.367
R1229 B.n416 B.n415 163.367
R1230 B.n415 B.n414 163.367
R1231 B.n414 B.n63 163.367
R1232 B.n410 B.n63 163.367
R1233 B.n410 B.n409 163.367
R1234 B.n409 B.n408 163.367
R1235 B.n548 B.n547 163.367
R1236 B.n548 B.n13 163.367
R1237 B.n552 B.n13 163.367
R1238 B.n553 B.n552 163.367
R1239 B.n554 B.n553 163.367
R1240 B.n554 B.n11 163.367
R1241 B.n558 B.n11 163.367
R1242 B.n559 B.n558 163.367
R1243 B.n560 B.n559 163.367
R1244 B.n560 B.n9 163.367
R1245 B.n564 B.n9 163.367
R1246 B.n565 B.n564 163.367
R1247 B.n566 B.n565 163.367
R1248 B.n566 B.n7 163.367
R1249 B.n570 B.n7 163.367
R1250 B.n571 B.n570 163.367
R1251 B.n572 B.n571 163.367
R1252 B.n572 B.n5 163.367
R1253 B.n576 B.n5 163.367
R1254 B.n577 B.n576 163.367
R1255 B.n578 B.n577 163.367
R1256 B.n578 B.n3 163.367
R1257 B.n582 B.n3 163.367
R1258 B.n583 B.n582 163.367
R1259 B.n152 B.n2 163.367
R1260 B.n153 B.n152 163.367
R1261 B.n154 B.n153 163.367
R1262 B.n154 B.n149 163.367
R1263 B.n158 B.n149 163.367
R1264 B.n159 B.n158 163.367
R1265 B.n160 B.n159 163.367
R1266 B.n160 B.n147 163.367
R1267 B.n164 B.n147 163.367
R1268 B.n165 B.n164 163.367
R1269 B.n166 B.n165 163.367
R1270 B.n166 B.n145 163.367
R1271 B.n170 B.n145 163.367
R1272 B.n171 B.n170 163.367
R1273 B.n172 B.n171 163.367
R1274 B.n172 B.n143 163.367
R1275 B.n176 B.n143 163.367
R1276 B.n177 B.n176 163.367
R1277 B.n178 B.n177 163.367
R1278 B.n178 B.n141 163.367
R1279 B.n182 B.n141 163.367
R1280 B.n183 B.n182 163.367
R1281 B.n184 B.n183 163.367
R1282 B.n184 B.n139 163.367
R1283 B.n249 B.n248 59.5399
R1284 B.n267 B.n113 59.5399
R1285 B.n44 B.n43 59.5399
R1286 B.n484 B.n37 59.5399
R1287 B.n545 B.n14 37.3078
R1288 B.n407 B.n406 37.3078
R1289 B.n329 B.n328 37.3078
R1290 B.n187 B.n186 37.3078
R1291 B.n248 B.n247 19.3944
R1292 B.n113 B.n112 19.3944
R1293 B.n43 B.n42 19.3944
R1294 B.n37 B.n36 19.3944
R1295 B B.n585 18.0485
R1296 B.n549 B.n14 10.6151
R1297 B.n550 B.n549 10.6151
R1298 B.n551 B.n550 10.6151
R1299 B.n551 B.n12 10.6151
R1300 B.n555 B.n12 10.6151
R1301 B.n556 B.n555 10.6151
R1302 B.n557 B.n556 10.6151
R1303 B.n557 B.n10 10.6151
R1304 B.n561 B.n10 10.6151
R1305 B.n562 B.n561 10.6151
R1306 B.n563 B.n562 10.6151
R1307 B.n563 B.n8 10.6151
R1308 B.n567 B.n8 10.6151
R1309 B.n568 B.n567 10.6151
R1310 B.n569 B.n568 10.6151
R1311 B.n569 B.n6 10.6151
R1312 B.n573 B.n6 10.6151
R1313 B.n574 B.n573 10.6151
R1314 B.n575 B.n574 10.6151
R1315 B.n575 B.n4 10.6151
R1316 B.n579 B.n4 10.6151
R1317 B.n580 B.n579 10.6151
R1318 B.n581 B.n580 10.6151
R1319 B.n581 B.n0 10.6151
R1320 B.n545 B.n544 10.6151
R1321 B.n544 B.n543 10.6151
R1322 B.n543 B.n16 10.6151
R1323 B.n539 B.n16 10.6151
R1324 B.n539 B.n538 10.6151
R1325 B.n538 B.n537 10.6151
R1326 B.n537 B.n18 10.6151
R1327 B.n533 B.n18 10.6151
R1328 B.n533 B.n532 10.6151
R1329 B.n532 B.n531 10.6151
R1330 B.n531 B.n20 10.6151
R1331 B.n527 B.n20 10.6151
R1332 B.n527 B.n526 10.6151
R1333 B.n526 B.n525 10.6151
R1334 B.n525 B.n22 10.6151
R1335 B.n521 B.n22 10.6151
R1336 B.n521 B.n520 10.6151
R1337 B.n520 B.n519 10.6151
R1338 B.n519 B.n24 10.6151
R1339 B.n515 B.n24 10.6151
R1340 B.n515 B.n514 10.6151
R1341 B.n514 B.n513 10.6151
R1342 B.n513 B.n26 10.6151
R1343 B.n509 B.n26 10.6151
R1344 B.n509 B.n508 10.6151
R1345 B.n508 B.n507 10.6151
R1346 B.n507 B.n28 10.6151
R1347 B.n503 B.n28 10.6151
R1348 B.n503 B.n502 10.6151
R1349 B.n502 B.n501 10.6151
R1350 B.n501 B.n30 10.6151
R1351 B.n497 B.n30 10.6151
R1352 B.n497 B.n496 10.6151
R1353 B.n496 B.n495 10.6151
R1354 B.n495 B.n32 10.6151
R1355 B.n491 B.n32 10.6151
R1356 B.n491 B.n490 10.6151
R1357 B.n490 B.n489 10.6151
R1358 B.n489 B.n34 10.6151
R1359 B.n485 B.n34 10.6151
R1360 B.n483 B.n482 10.6151
R1361 B.n482 B.n38 10.6151
R1362 B.n478 B.n38 10.6151
R1363 B.n478 B.n477 10.6151
R1364 B.n477 B.n476 10.6151
R1365 B.n476 B.n40 10.6151
R1366 B.n472 B.n40 10.6151
R1367 B.n472 B.n471 10.6151
R1368 B.n471 B.n470 10.6151
R1369 B.n467 B.n466 10.6151
R1370 B.n466 B.n465 10.6151
R1371 B.n465 B.n46 10.6151
R1372 B.n461 B.n46 10.6151
R1373 B.n461 B.n460 10.6151
R1374 B.n460 B.n459 10.6151
R1375 B.n459 B.n48 10.6151
R1376 B.n455 B.n48 10.6151
R1377 B.n455 B.n454 10.6151
R1378 B.n454 B.n453 10.6151
R1379 B.n453 B.n50 10.6151
R1380 B.n449 B.n50 10.6151
R1381 B.n449 B.n448 10.6151
R1382 B.n448 B.n447 10.6151
R1383 B.n447 B.n52 10.6151
R1384 B.n443 B.n52 10.6151
R1385 B.n443 B.n442 10.6151
R1386 B.n442 B.n441 10.6151
R1387 B.n441 B.n54 10.6151
R1388 B.n437 B.n54 10.6151
R1389 B.n437 B.n436 10.6151
R1390 B.n436 B.n435 10.6151
R1391 B.n435 B.n56 10.6151
R1392 B.n431 B.n56 10.6151
R1393 B.n431 B.n430 10.6151
R1394 B.n430 B.n429 10.6151
R1395 B.n429 B.n58 10.6151
R1396 B.n425 B.n58 10.6151
R1397 B.n425 B.n424 10.6151
R1398 B.n424 B.n423 10.6151
R1399 B.n423 B.n60 10.6151
R1400 B.n419 B.n60 10.6151
R1401 B.n419 B.n418 10.6151
R1402 B.n418 B.n417 10.6151
R1403 B.n417 B.n62 10.6151
R1404 B.n413 B.n62 10.6151
R1405 B.n413 B.n412 10.6151
R1406 B.n412 B.n411 10.6151
R1407 B.n411 B.n64 10.6151
R1408 B.n407 B.n64 10.6151
R1409 B.n406 B.n405 10.6151
R1410 B.n405 B.n66 10.6151
R1411 B.n401 B.n66 10.6151
R1412 B.n401 B.n400 10.6151
R1413 B.n400 B.n399 10.6151
R1414 B.n399 B.n68 10.6151
R1415 B.n395 B.n68 10.6151
R1416 B.n395 B.n394 10.6151
R1417 B.n394 B.n393 10.6151
R1418 B.n393 B.n70 10.6151
R1419 B.n389 B.n70 10.6151
R1420 B.n389 B.n388 10.6151
R1421 B.n388 B.n387 10.6151
R1422 B.n387 B.n72 10.6151
R1423 B.n383 B.n72 10.6151
R1424 B.n383 B.n382 10.6151
R1425 B.n382 B.n381 10.6151
R1426 B.n381 B.n74 10.6151
R1427 B.n377 B.n74 10.6151
R1428 B.n377 B.n376 10.6151
R1429 B.n376 B.n375 10.6151
R1430 B.n375 B.n76 10.6151
R1431 B.n371 B.n76 10.6151
R1432 B.n371 B.n370 10.6151
R1433 B.n370 B.n369 10.6151
R1434 B.n369 B.n78 10.6151
R1435 B.n365 B.n78 10.6151
R1436 B.n365 B.n364 10.6151
R1437 B.n364 B.n363 10.6151
R1438 B.n363 B.n80 10.6151
R1439 B.n359 B.n80 10.6151
R1440 B.n359 B.n358 10.6151
R1441 B.n358 B.n357 10.6151
R1442 B.n357 B.n82 10.6151
R1443 B.n353 B.n82 10.6151
R1444 B.n353 B.n352 10.6151
R1445 B.n352 B.n351 10.6151
R1446 B.n351 B.n84 10.6151
R1447 B.n347 B.n84 10.6151
R1448 B.n347 B.n346 10.6151
R1449 B.n346 B.n345 10.6151
R1450 B.n345 B.n86 10.6151
R1451 B.n341 B.n86 10.6151
R1452 B.n341 B.n340 10.6151
R1453 B.n340 B.n339 10.6151
R1454 B.n339 B.n88 10.6151
R1455 B.n335 B.n88 10.6151
R1456 B.n335 B.n334 10.6151
R1457 B.n334 B.n333 10.6151
R1458 B.n333 B.n90 10.6151
R1459 B.n329 B.n90 10.6151
R1460 B.n151 B.n1 10.6151
R1461 B.n151 B.n150 10.6151
R1462 B.n155 B.n150 10.6151
R1463 B.n156 B.n155 10.6151
R1464 B.n157 B.n156 10.6151
R1465 B.n157 B.n148 10.6151
R1466 B.n161 B.n148 10.6151
R1467 B.n162 B.n161 10.6151
R1468 B.n163 B.n162 10.6151
R1469 B.n163 B.n146 10.6151
R1470 B.n167 B.n146 10.6151
R1471 B.n168 B.n167 10.6151
R1472 B.n169 B.n168 10.6151
R1473 B.n169 B.n144 10.6151
R1474 B.n173 B.n144 10.6151
R1475 B.n174 B.n173 10.6151
R1476 B.n175 B.n174 10.6151
R1477 B.n175 B.n142 10.6151
R1478 B.n179 B.n142 10.6151
R1479 B.n180 B.n179 10.6151
R1480 B.n181 B.n180 10.6151
R1481 B.n181 B.n140 10.6151
R1482 B.n185 B.n140 10.6151
R1483 B.n186 B.n185 10.6151
R1484 B.n187 B.n138 10.6151
R1485 B.n191 B.n138 10.6151
R1486 B.n192 B.n191 10.6151
R1487 B.n193 B.n192 10.6151
R1488 B.n193 B.n136 10.6151
R1489 B.n197 B.n136 10.6151
R1490 B.n198 B.n197 10.6151
R1491 B.n199 B.n198 10.6151
R1492 B.n199 B.n134 10.6151
R1493 B.n203 B.n134 10.6151
R1494 B.n204 B.n203 10.6151
R1495 B.n205 B.n204 10.6151
R1496 B.n205 B.n132 10.6151
R1497 B.n209 B.n132 10.6151
R1498 B.n210 B.n209 10.6151
R1499 B.n211 B.n210 10.6151
R1500 B.n211 B.n130 10.6151
R1501 B.n215 B.n130 10.6151
R1502 B.n216 B.n215 10.6151
R1503 B.n217 B.n216 10.6151
R1504 B.n217 B.n128 10.6151
R1505 B.n221 B.n128 10.6151
R1506 B.n222 B.n221 10.6151
R1507 B.n223 B.n222 10.6151
R1508 B.n223 B.n126 10.6151
R1509 B.n227 B.n126 10.6151
R1510 B.n228 B.n227 10.6151
R1511 B.n229 B.n228 10.6151
R1512 B.n229 B.n124 10.6151
R1513 B.n233 B.n124 10.6151
R1514 B.n234 B.n233 10.6151
R1515 B.n235 B.n234 10.6151
R1516 B.n235 B.n122 10.6151
R1517 B.n239 B.n122 10.6151
R1518 B.n240 B.n239 10.6151
R1519 B.n241 B.n240 10.6151
R1520 B.n241 B.n120 10.6151
R1521 B.n245 B.n120 10.6151
R1522 B.n246 B.n245 10.6151
R1523 B.n250 B.n246 10.6151
R1524 B.n254 B.n118 10.6151
R1525 B.n255 B.n254 10.6151
R1526 B.n256 B.n255 10.6151
R1527 B.n256 B.n116 10.6151
R1528 B.n260 B.n116 10.6151
R1529 B.n261 B.n260 10.6151
R1530 B.n262 B.n261 10.6151
R1531 B.n262 B.n114 10.6151
R1532 B.n266 B.n114 10.6151
R1533 B.n269 B.n268 10.6151
R1534 B.n269 B.n110 10.6151
R1535 B.n273 B.n110 10.6151
R1536 B.n274 B.n273 10.6151
R1537 B.n275 B.n274 10.6151
R1538 B.n275 B.n108 10.6151
R1539 B.n279 B.n108 10.6151
R1540 B.n280 B.n279 10.6151
R1541 B.n281 B.n280 10.6151
R1542 B.n281 B.n106 10.6151
R1543 B.n285 B.n106 10.6151
R1544 B.n286 B.n285 10.6151
R1545 B.n287 B.n286 10.6151
R1546 B.n287 B.n104 10.6151
R1547 B.n291 B.n104 10.6151
R1548 B.n292 B.n291 10.6151
R1549 B.n293 B.n292 10.6151
R1550 B.n293 B.n102 10.6151
R1551 B.n297 B.n102 10.6151
R1552 B.n298 B.n297 10.6151
R1553 B.n299 B.n298 10.6151
R1554 B.n299 B.n100 10.6151
R1555 B.n303 B.n100 10.6151
R1556 B.n304 B.n303 10.6151
R1557 B.n305 B.n304 10.6151
R1558 B.n305 B.n98 10.6151
R1559 B.n309 B.n98 10.6151
R1560 B.n310 B.n309 10.6151
R1561 B.n311 B.n310 10.6151
R1562 B.n311 B.n96 10.6151
R1563 B.n315 B.n96 10.6151
R1564 B.n316 B.n315 10.6151
R1565 B.n317 B.n316 10.6151
R1566 B.n317 B.n94 10.6151
R1567 B.n321 B.n94 10.6151
R1568 B.n322 B.n321 10.6151
R1569 B.n323 B.n322 10.6151
R1570 B.n323 B.n92 10.6151
R1571 B.n327 B.n92 10.6151
R1572 B.n328 B.n327 10.6151
R1573 B.n485 B.n484 9.36635
R1574 B.n467 B.n44 9.36635
R1575 B.n250 B.n249 9.36635
R1576 B.n268 B.n267 9.36635
R1577 B.n585 B.n0 8.11757
R1578 B.n585 B.n1 8.11757
R1579 B.n484 B.n483 1.24928
R1580 B.n470 B.n44 1.24928
R1581 B.n249 B.n118 1.24928
R1582 B.n267 B.n266 1.24928
R1583 VP.n7 VP.t9 509.111
R1584 VP.n18 VP.t8 488.115
R1585 VP.n22 VP.t0 488.115
R1586 VP.n24 VP.t2 488.115
R1587 VP.n28 VP.t4 488.115
R1588 VP.n30 VP.t6 488.115
R1589 VP.n16 VP.t5 488.115
R1590 VP.n14 VP.t1 488.115
R1591 VP.n6 VP.t7 488.115
R1592 VP.n8 VP.t3 488.115
R1593 VP.n31 VP.n30 161.3
R1594 VP.n10 VP.n9 161.3
R1595 VP.n11 VP.n6 161.3
R1596 VP.n13 VP.n12 161.3
R1597 VP.n14 VP.n5 161.3
R1598 VP.n15 VP.n4 161.3
R1599 VP.n17 VP.n16 161.3
R1600 VP.n29 VP.n0 161.3
R1601 VP.n28 VP.n27 161.3
R1602 VP.n26 VP.n1 161.3
R1603 VP.n25 VP.n24 161.3
R1604 VP.n23 VP.n2 161.3
R1605 VP.n22 VP.n21 161.3
R1606 VP.n20 VP.n3 161.3
R1607 VP.n19 VP.n18 161.3
R1608 VP.n10 VP.n7 44.8515
R1609 VP.n19 VP.n17 42.5156
R1610 VP.n18 VP.n3 24.1005
R1611 VP.n22 VP.n3 24.1005
R1612 VP.n23 VP.n22 24.1005
R1613 VP.n24 VP.n23 24.1005
R1614 VP.n24 VP.n1 24.1005
R1615 VP.n28 VP.n1 24.1005
R1616 VP.n29 VP.n28 24.1005
R1617 VP.n30 VP.n29 24.1005
R1618 VP.n15 VP.n14 24.1005
R1619 VP.n16 VP.n15 24.1005
R1620 VP.n13 VP.n6 24.1005
R1621 VP.n14 VP.n13 24.1005
R1622 VP.n9 VP.n8 24.1005
R1623 VP.n9 VP.n6 24.1005
R1624 VP.n8 VP.n7 20.9471
R1625 VP.n11 VP.n10 0.189894
R1626 VP.n12 VP.n11 0.189894
R1627 VP.n12 VP.n5 0.189894
R1628 VP.n5 VP.n4 0.189894
R1629 VP.n17 VP.n4 0.189894
R1630 VP.n20 VP.n19 0.189894
R1631 VP.n21 VP.n20 0.189894
R1632 VP.n21 VP.n2 0.189894
R1633 VP.n25 VP.n2 0.189894
R1634 VP.n26 VP.n25 0.189894
R1635 VP.n27 VP.n26 0.189894
R1636 VP.n27 VP.n0 0.189894
R1637 VP.n31 VP.n0 0.189894
R1638 VP VP.n31 0.0516364
R1639 VDD1.n64 VDD1.n63 756.745
R1640 VDD1.n131 VDD1.n130 756.745
R1641 VDD1.n63 VDD1.n62 585
R1642 VDD1.n2 VDD1.n1 585
R1643 VDD1.n57 VDD1.n56 585
R1644 VDD1.n55 VDD1.n54 585
R1645 VDD1.n6 VDD1.n5 585
R1646 VDD1.n49 VDD1.n48 585
R1647 VDD1.n47 VDD1.n46 585
R1648 VDD1.n10 VDD1.n9 585
R1649 VDD1.n41 VDD1.n40 585
R1650 VDD1.n39 VDD1.n38 585
R1651 VDD1.n14 VDD1.n13 585
R1652 VDD1.n33 VDD1.n32 585
R1653 VDD1.n31 VDD1.n30 585
R1654 VDD1.n18 VDD1.n17 585
R1655 VDD1.n25 VDD1.n24 585
R1656 VDD1.n23 VDD1.n22 585
R1657 VDD1.n90 VDD1.n89 585
R1658 VDD1.n92 VDD1.n91 585
R1659 VDD1.n85 VDD1.n84 585
R1660 VDD1.n98 VDD1.n97 585
R1661 VDD1.n100 VDD1.n99 585
R1662 VDD1.n81 VDD1.n80 585
R1663 VDD1.n106 VDD1.n105 585
R1664 VDD1.n108 VDD1.n107 585
R1665 VDD1.n77 VDD1.n76 585
R1666 VDD1.n114 VDD1.n113 585
R1667 VDD1.n116 VDD1.n115 585
R1668 VDD1.n73 VDD1.n72 585
R1669 VDD1.n122 VDD1.n121 585
R1670 VDD1.n124 VDD1.n123 585
R1671 VDD1.n69 VDD1.n68 585
R1672 VDD1.n130 VDD1.n129 585
R1673 VDD1.n21 VDD1.t0 327.466
R1674 VDD1.n88 VDD1.t1 327.466
R1675 VDD1.n63 VDD1.n1 171.744
R1676 VDD1.n56 VDD1.n1 171.744
R1677 VDD1.n56 VDD1.n55 171.744
R1678 VDD1.n55 VDD1.n5 171.744
R1679 VDD1.n48 VDD1.n5 171.744
R1680 VDD1.n48 VDD1.n47 171.744
R1681 VDD1.n47 VDD1.n9 171.744
R1682 VDD1.n40 VDD1.n9 171.744
R1683 VDD1.n40 VDD1.n39 171.744
R1684 VDD1.n39 VDD1.n13 171.744
R1685 VDD1.n32 VDD1.n13 171.744
R1686 VDD1.n32 VDD1.n31 171.744
R1687 VDD1.n31 VDD1.n17 171.744
R1688 VDD1.n24 VDD1.n17 171.744
R1689 VDD1.n24 VDD1.n23 171.744
R1690 VDD1.n91 VDD1.n90 171.744
R1691 VDD1.n91 VDD1.n84 171.744
R1692 VDD1.n98 VDD1.n84 171.744
R1693 VDD1.n99 VDD1.n98 171.744
R1694 VDD1.n99 VDD1.n80 171.744
R1695 VDD1.n106 VDD1.n80 171.744
R1696 VDD1.n107 VDD1.n106 171.744
R1697 VDD1.n107 VDD1.n76 171.744
R1698 VDD1.n114 VDD1.n76 171.744
R1699 VDD1.n115 VDD1.n114 171.744
R1700 VDD1.n115 VDD1.n72 171.744
R1701 VDD1.n122 VDD1.n72 171.744
R1702 VDD1.n123 VDD1.n122 171.744
R1703 VDD1.n123 VDD1.n68 171.744
R1704 VDD1.n130 VDD1.n68 171.744
R1705 VDD1.n23 VDD1.t0 85.8723
R1706 VDD1.n90 VDD1.t1 85.8723
R1707 VDD1.n135 VDD1.n134 77.3039
R1708 VDD1.n66 VDD1.n65 76.7129
R1709 VDD1.n133 VDD1.n132 76.7127
R1710 VDD1.n137 VDD1.n136 76.7118
R1711 VDD1.n66 VDD1.n64 51.8595
R1712 VDD1.n133 VDD1.n131 51.8595
R1713 VDD1.n137 VDD1.n135 39.1087
R1714 VDD1.n22 VDD1.n21 16.3895
R1715 VDD1.n89 VDD1.n88 16.3895
R1716 VDD1.n25 VDD1.n20 12.8005
R1717 VDD1.n92 VDD1.n87 12.8005
R1718 VDD1.n62 VDD1.n0 12.0247
R1719 VDD1.n26 VDD1.n18 12.0247
R1720 VDD1.n93 VDD1.n85 12.0247
R1721 VDD1.n129 VDD1.n67 12.0247
R1722 VDD1.n61 VDD1.n2 11.249
R1723 VDD1.n30 VDD1.n29 11.249
R1724 VDD1.n97 VDD1.n96 11.249
R1725 VDD1.n128 VDD1.n69 11.249
R1726 VDD1.n58 VDD1.n57 10.4732
R1727 VDD1.n33 VDD1.n16 10.4732
R1728 VDD1.n100 VDD1.n83 10.4732
R1729 VDD1.n125 VDD1.n124 10.4732
R1730 VDD1.n54 VDD1.n4 9.69747
R1731 VDD1.n34 VDD1.n14 9.69747
R1732 VDD1.n101 VDD1.n81 9.69747
R1733 VDD1.n121 VDD1.n71 9.69747
R1734 VDD1.n60 VDD1.n0 9.45567
R1735 VDD1.n127 VDD1.n67 9.45567
R1736 VDD1.n8 VDD1.n7 9.3005
R1737 VDD1.n51 VDD1.n50 9.3005
R1738 VDD1.n53 VDD1.n52 9.3005
R1739 VDD1.n4 VDD1.n3 9.3005
R1740 VDD1.n59 VDD1.n58 9.3005
R1741 VDD1.n61 VDD1.n60 9.3005
R1742 VDD1.n45 VDD1.n44 9.3005
R1743 VDD1.n43 VDD1.n42 9.3005
R1744 VDD1.n12 VDD1.n11 9.3005
R1745 VDD1.n37 VDD1.n36 9.3005
R1746 VDD1.n35 VDD1.n34 9.3005
R1747 VDD1.n16 VDD1.n15 9.3005
R1748 VDD1.n29 VDD1.n28 9.3005
R1749 VDD1.n27 VDD1.n26 9.3005
R1750 VDD1.n20 VDD1.n19 9.3005
R1751 VDD1.n112 VDD1.n111 9.3005
R1752 VDD1.n75 VDD1.n74 9.3005
R1753 VDD1.n118 VDD1.n117 9.3005
R1754 VDD1.n120 VDD1.n119 9.3005
R1755 VDD1.n71 VDD1.n70 9.3005
R1756 VDD1.n126 VDD1.n125 9.3005
R1757 VDD1.n128 VDD1.n127 9.3005
R1758 VDD1.n79 VDD1.n78 9.3005
R1759 VDD1.n104 VDD1.n103 9.3005
R1760 VDD1.n102 VDD1.n101 9.3005
R1761 VDD1.n83 VDD1.n82 9.3005
R1762 VDD1.n96 VDD1.n95 9.3005
R1763 VDD1.n94 VDD1.n93 9.3005
R1764 VDD1.n87 VDD1.n86 9.3005
R1765 VDD1.n110 VDD1.n109 9.3005
R1766 VDD1.n53 VDD1.n6 8.92171
R1767 VDD1.n38 VDD1.n37 8.92171
R1768 VDD1.n105 VDD1.n104 8.92171
R1769 VDD1.n120 VDD1.n73 8.92171
R1770 VDD1.n50 VDD1.n49 8.14595
R1771 VDD1.n41 VDD1.n12 8.14595
R1772 VDD1.n108 VDD1.n79 8.14595
R1773 VDD1.n117 VDD1.n116 8.14595
R1774 VDD1.n46 VDD1.n8 7.3702
R1775 VDD1.n42 VDD1.n10 7.3702
R1776 VDD1.n109 VDD1.n77 7.3702
R1777 VDD1.n113 VDD1.n75 7.3702
R1778 VDD1.n46 VDD1.n45 6.59444
R1779 VDD1.n45 VDD1.n10 6.59444
R1780 VDD1.n112 VDD1.n77 6.59444
R1781 VDD1.n113 VDD1.n112 6.59444
R1782 VDD1.n49 VDD1.n8 5.81868
R1783 VDD1.n42 VDD1.n41 5.81868
R1784 VDD1.n109 VDD1.n108 5.81868
R1785 VDD1.n116 VDD1.n75 5.81868
R1786 VDD1.n50 VDD1.n6 5.04292
R1787 VDD1.n38 VDD1.n12 5.04292
R1788 VDD1.n105 VDD1.n79 5.04292
R1789 VDD1.n117 VDD1.n73 5.04292
R1790 VDD1.n54 VDD1.n53 4.26717
R1791 VDD1.n37 VDD1.n14 4.26717
R1792 VDD1.n104 VDD1.n81 4.26717
R1793 VDD1.n121 VDD1.n120 4.26717
R1794 VDD1.n21 VDD1.n19 3.70982
R1795 VDD1.n88 VDD1.n86 3.70982
R1796 VDD1.n57 VDD1.n4 3.49141
R1797 VDD1.n34 VDD1.n33 3.49141
R1798 VDD1.n101 VDD1.n100 3.49141
R1799 VDD1.n124 VDD1.n71 3.49141
R1800 VDD1.n136 VDD1.t8 2.72514
R1801 VDD1.n136 VDD1.t4 2.72514
R1802 VDD1.n65 VDD1.t6 2.72514
R1803 VDD1.n65 VDD1.t2 2.72514
R1804 VDD1.n134 VDD1.t5 2.72514
R1805 VDD1.n134 VDD1.t3 2.72514
R1806 VDD1.n132 VDD1.t9 2.72514
R1807 VDD1.n132 VDD1.t7 2.72514
R1808 VDD1.n58 VDD1.n2 2.71565
R1809 VDD1.n30 VDD1.n16 2.71565
R1810 VDD1.n97 VDD1.n83 2.71565
R1811 VDD1.n125 VDD1.n69 2.71565
R1812 VDD1.n62 VDD1.n61 1.93989
R1813 VDD1.n29 VDD1.n18 1.93989
R1814 VDD1.n96 VDD1.n85 1.93989
R1815 VDD1.n129 VDD1.n128 1.93989
R1816 VDD1.n64 VDD1.n0 1.16414
R1817 VDD1.n26 VDD1.n25 1.16414
R1818 VDD1.n93 VDD1.n92 1.16414
R1819 VDD1.n131 VDD1.n67 1.16414
R1820 VDD1 VDD1.n137 0.588862
R1821 VDD1.n22 VDD1.n20 0.388379
R1822 VDD1.n89 VDD1.n87 0.388379
R1823 VDD1 VDD1.n66 0.274207
R1824 VDD1.n135 VDD1.n133 0.160671
R1825 VDD1.n60 VDD1.n59 0.155672
R1826 VDD1.n59 VDD1.n3 0.155672
R1827 VDD1.n52 VDD1.n3 0.155672
R1828 VDD1.n52 VDD1.n51 0.155672
R1829 VDD1.n51 VDD1.n7 0.155672
R1830 VDD1.n44 VDD1.n7 0.155672
R1831 VDD1.n44 VDD1.n43 0.155672
R1832 VDD1.n43 VDD1.n11 0.155672
R1833 VDD1.n36 VDD1.n11 0.155672
R1834 VDD1.n36 VDD1.n35 0.155672
R1835 VDD1.n35 VDD1.n15 0.155672
R1836 VDD1.n28 VDD1.n15 0.155672
R1837 VDD1.n28 VDD1.n27 0.155672
R1838 VDD1.n27 VDD1.n19 0.155672
R1839 VDD1.n94 VDD1.n86 0.155672
R1840 VDD1.n95 VDD1.n94 0.155672
R1841 VDD1.n95 VDD1.n82 0.155672
R1842 VDD1.n102 VDD1.n82 0.155672
R1843 VDD1.n103 VDD1.n102 0.155672
R1844 VDD1.n103 VDD1.n78 0.155672
R1845 VDD1.n110 VDD1.n78 0.155672
R1846 VDD1.n111 VDD1.n110 0.155672
R1847 VDD1.n111 VDD1.n74 0.155672
R1848 VDD1.n118 VDD1.n74 0.155672
R1849 VDD1.n119 VDD1.n118 0.155672
R1850 VDD1.n119 VDD1.n70 0.155672
R1851 VDD1.n126 VDD1.n70 0.155672
R1852 VDD1.n127 VDD1.n126 0.155672
C0 VDD2 VDD1 0.950406f
C1 VN w_n2170_n3354# 4.07137f
C2 w_n2170_n3354# VP 4.34794f
C3 VN B 0.789855f
C4 B VP 1.24427f
C5 w_n2170_n3354# VDD2 2.0582f
C6 VTAIL VDD1 14.4186f
C7 VDD2 B 1.72836f
C8 VTAIL w_n2170_n3354# 2.9876f
C9 VTAIL B 2.69914f
C10 VN VP 5.5433f
C11 VN VDD2 6.5078f
C12 VDD2 VP 0.33728f
C13 w_n2170_n3354# VDD1 2.01514f
C14 B VDD1 1.68523f
C15 VTAIL VN 6.3313f
C16 VTAIL VP 6.34591f
C17 VTAIL VDD2 14.452499f
C18 w_n2170_n3354# B 7.28441f
C19 VN VDD1 0.148475f
C20 VDD1 VP 6.69189f
C21 VDD2 VSUBS 1.437567f
C22 VDD1 VSUBS 1.150134f
C23 VTAIL VSUBS 0.755948f
C24 VN VSUBS 4.87902f
C25 VP VSUBS 1.772159f
C26 B VSUBS 2.967307f
C27 w_n2170_n3354# VSUBS 89.60361f
C28 VDD1.n0 VSUBS 0.015243f
C29 VDD1.n1 VSUBS 0.034382f
C30 VDD1.n2 VSUBS 0.015402f
C31 VDD1.n3 VSUBS 0.02707f
C32 VDD1.n4 VSUBS 0.014546f
C33 VDD1.n5 VSUBS 0.034382f
C34 VDD1.n6 VSUBS 0.015402f
C35 VDD1.n7 VSUBS 0.02707f
C36 VDD1.n8 VSUBS 0.014546f
C37 VDD1.n9 VSUBS 0.034382f
C38 VDD1.n10 VSUBS 0.015402f
C39 VDD1.n11 VSUBS 0.02707f
C40 VDD1.n12 VSUBS 0.014546f
C41 VDD1.n13 VSUBS 0.034382f
C42 VDD1.n14 VSUBS 0.015402f
C43 VDD1.n15 VSUBS 0.02707f
C44 VDD1.n16 VSUBS 0.014546f
C45 VDD1.n17 VSUBS 0.034382f
C46 VDD1.n18 VSUBS 0.015402f
C47 VDD1.n19 VSUBS 1.35119f
C48 VDD1.n20 VSUBS 0.014546f
C49 VDD1.t0 VSUBS 0.073402f
C50 VDD1.n21 VSUBS 0.166311f
C51 VDD1.n22 VSUBS 0.021872f
C52 VDD1.n23 VSUBS 0.025786f
C53 VDD1.n24 VSUBS 0.034382f
C54 VDD1.n25 VSUBS 0.015402f
C55 VDD1.n26 VSUBS 0.014546f
C56 VDD1.n27 VSUBS 0.02707f
C57 VDD1.n28 VSUBS 0.02707f
C58 VDD1.n29 VSUBS 0.014546f
C59 VDD1.n30 VSUBS 0.015402f
C60 VDD1.n31 VSUBS 0.034382f
C61 VDD1.n32 VSUBS 0.034382f
C62 VDD1.n33 VSUBS 0.015402f
C63 VDD1.n34 VSUBS 0.014546f
C64 VDD1.n35 VSUBS 0.02707f
C65 VDD1.n36 VSUBS 0.02707f
C66 VDD1.n37 VSUBS 0.014546f
C67 VDD1.n38 VSUBS 0.015402f
C68 VDD1.n39 VSUBS 0.034382f
C69 VDD1.n40 VSUBS 0.034382f
C70 VDD1.n41 VSUBS 0.015402f
C71 VDD1.n42 VSUBS 0.014546f
C72 VDD1.n43 VSUBS 0.02707f
C73 VDD1.n44 VSUBS 0.02707f
C74 VDD1.n45 VSUBS 0.014546f
C75 VDD1.n46 VSUBS 0.015402f
C76 VDD1.n47 VSUBS 0.034382f
C77 VDD1.n48 VSUBS 0.034382f
C78 VDD1.n49 VSUBS 0.015402f
C79 VDD1.n50 VSUBS 0.014546f
C80 VDD1.n51 VSUBS 0.02707f
C81 VDD1.n52 VSUBS 0.02707f
C82 VDD1.n53 VSUBS 0.014546f
C83 VDD1.n54 VSUBS 0.015402f
C84 VDD1.n55 VSUBS 0.034382f
C85 VDD1.n56 VSUBS 0.034382f
C86 VDD1.n57 VSUBS 0.015402f
C87 VDD1.n58 VSUBS 0.014546f
C88 VDD1.n59 VSUBS 0.02707f
C89 VDD1.n60 VSUBS 0.068857f
C90 VDD1.n61 VSUBS 0.014546f
C91 VDD1.n62 VSUBS 0.015402f
C92 VDD1.n63 VSUBS 0.075423f
C93 VDD1.n64 VSUBS 0.071192f
C94 VDD1.t6 VSUBS 0.2552f
C95 VDD1.t2 VSUBS 0.2552f
C96 VDD1.n65 VSUBS 2.01243f
C97 VDD1.n66 VSUBS 0.711276f
C98 VDD1.n67 VSUBS 0.015243f
C99 VDD1.n68 VSUBS 0.034382f
C100 VDD1.n69 VSUBS 0.015402f
C101 VDD1.n70 VSUBS 0.02707f
C102 VDD1.n71 VSUBS 0.014546f
C103 VDD1.n72 VSUBS 0.034382f
C104 VDD1.n73 VSUBS 0.015402f
C105 VDD1.n74 VSUBS 0.02707f
C106 VDD1.n75 VSUBS 0.014546f
C107 VDD1.n76 VSUBS 0.034382f
C108 VDD1.n77 VSUBS 0.015402f
C109 VDD1.n78 VSUBS 0.02707f
C110 VDD1.n79 VSUBS 0.014546f
C111 VDD1.n80 VSUBS 0.034382f
C112 VDD1.n81 VSUBS 0.015402f
C113 VDD1.n82 VSUBS 0.02707f
C114 VDD1.n83 VSUBS 0.014546f
C115 VDD1.n84 VSUBS 0.034382f
C116 VDD1.n85 VSUBS 0.015402f
C117 VDD1.n86 VSUBS 1.35119f
C118 VDD1.n87 VSUBS 0.014546f
C119 VDD1.t1 VSUBS 0.073402f
C120 VDD1.n88 VSUBS 0.166311f
C121 VDD1.n89 VSUBS 0.021872f
C122 VDD1.n90 VSUBS 0.025786f
C123 VDD1.n91 VSUBS 0.034382f
C124 VDD1.n92 VSUBS 0.015402f
C125 VDD1.n93 VSUBS 0.014546f
C126 VDD1.n94 VSUBS 0.02707f
C127 VDD1.n95 VSUBS 0.02707f
C128 VDD1.n96 VSUBS 0.014546f
C129 VDD1.n97 VSUBS 0.015402f
C130 VDD1.n98 VSUBS 0.034382f
C131 VDD1.n99 VSUBS 0.034382f
C132 VDD1.n100 VSUBS 0.015402f
C133 VDD1.n101 VSUBS 0.014546f
C134 VDD1.n102 VSUBS 0.02707f
C135 VDD1.n103 VSUBS 0.02707f
C136 VDD1.n104 VSUBS 0.014546f
C137 VDD1.n105 VSUBS 0.015402f
C138 VDD1.n106 VSUBS 0.034382f
C139 VDD1.n107 VSUBS 0.034382f
C140 VDD1.n108 VSUBS 0.015402f
C141 VDD1.n109 VSUBS 0.014546f
C142 VDD1.n110 VSUBS 0.02707f
C143 VDD1.n111 VSUBS 0.02707f
C144 VDD1.n112 VSUBS 0.014546f
C145 VDD1.n113 VSUBS 0.015402f
C146 VDD1.n114 VSUBS 0.034382f
C147 VDD1.n115 VSUBS 0.034382f
C148 VDD1.n116 VSUBS 0.015402f
C149 VDD1.n117 VSUBS 0.014546f
C150 VDD1.n118 VSUBS 0.02707f
C151 VDD1.n119 VSUBS 0.02707f
C152 VDD1.n120 VSUBS 0.014546f
C153 VDD1.n121 VSUBS 0.015402f
C154 VDD1.n122 VSUBS 0.034382f
C155 VDD1.n123 VSUBS 0.034382f
C156 VDD1.n124 VSUBS 0.015402f
C157 VDD1.n125 VSUBS 0.014546f
C158 VDD1.n126 VSUBS 0.02707f
C159 VDD1.n127 VSUBS 0.068857f
C160 VDD1.n128 VSUBS 0.014546f
C161 VDD1.n129 VSUBS 0.015402f
C162 VDD1.n130 VSUBS 0.075423f
C163 VDD1.n131 VSUBS 0.071192f
C164 VDD1.t9 VSUBS 0.2552f
C165 VDD1.t7 VSUBS 0.2552f
C166 VDD1.n132 VSUBS 2.01242f
C167 VDD1.n133 VSUBS 0.705298f
C168 VDD1.t5 VSUBS 0.2552f
C169 VDD1.t3 VSUBS 0.2552f
C170 VDD1.n134 VSUBS 2.01719f
C171 VDD1.n135 VSUBS 2.3819f
C172 VDD1.t8 VSUBS 0.2552f
C173 VDD1.t4 VSUBS 0.2552f
C174 VDD1.n136 VSUBS 2.01242f
C175 VDD1.n137 VSUBS 2.82679f
C176 VP.n0 VSUBS 0.054022f
C177 VP.n1 VSUBS 0.012259f
C178 VP.n2 VSUBS 0.054022f
C179 VP.n3 VSUBS 0.012259f
C180 VP.n4 VSUBS 0.054022f
C181 VP.t5 VSUBS 1.23176f
C182 VP.t1 VSUBS 1.23176f
C183 VP.n5 VSUBS 0.054022f
C184 VP.t7 VSUBS 1.23176f
C185 VP.n6 VSUBS 0.493399f
C186 VP.t9 VSUBS 1.25205f
C187 VP.n7 VSUBS 0.477043f
C188 VP.t3 VSUBS 1.23176f
C189 VP.n8 VSUBS 0.49729f
C190 VP.n9 VSUBS 0.012259f
C191 VP.n10 VSUBS 0.220688f
C192 VP.n11 VSUBS 0.054022f
C193 VP.n12 VSUBS 0.054022f
C194 VP.n13 VSUBS 0.012259f
C195 VP.n14 VSUBS 0.493399f
C196 VP.n15 VSUBS 0.012259f
C197 VP.n16 VSUBS 0.487903f
C198 VP.n17 VSUBS 2.27549f
C199 VP.t8 VSUBS 1.23176f
C200 VP.n18 VSUBS 0.487903f
C201 VP.n19 VSUBS 2.32117f
C202 VP.n20 VSUBS 0.054022f
C203 VP.n21 VSUBS 0.054022f
C204 VP.t0 VSUBS 1.23176f
C205 VP.n22 VSUBS 0.493399f
C206 VP.n23 VSUBS 0.012259f
C207 VP.t2 VSUBS 1.23176f
C208 VP.n24 VSUBS 0.493399f
C209 VP.n25 VSUBS 0.054022f
C210 VP.n26 VSUBS 0.054022f
C211 VP.n27 VSUBS 0.054022f
C212 VP.t4 VSUBS 1.23176f
C213 VP.n28 VSUBS 0.493399f
C214 VP.n29 VSUBS 0.012259f
C215 VP.t6 VSUBS 1.23176f
C216 VP.n30 VSUBS 0.487903f
C217 VP.n31 VSUBS 0.041865f
C218 B.n0 VSUBS 0.006495f
C219 B.n1 VSUBS 0.006495f
C220 B.n2 VSUBS 0.009606f
C221 B.n3 VSUBS 0.007361f
C222 B.n4 VSUBS 0.007361f
C223 B.n5 VSUBS 0.007361f
C224 B.n6 VSUBS 0.007361f
C225 B.n7 VSUBS 0.007361f
C226 B.n8 VSUBS 0.007361f
C227 B.n9 VSUBS 0.007361f
C228 B.n10 VSUBS 0.007361f
C229 B.n11 VSUBS 0.007361f
C230 B.n12 VSUBS 0.007361f
C231 B.n13 VSUBS 0.007361f
C232 B.n14 VSUBS 0.018437f
C233 B.n15 VSUBS 0.007361f
C234 B.n16 VSUBS 0.007361f
C235 B.n17 VSUBS 0.007361f
C236 B.n18 VSUBS 0.007361f
C237 B.n19 VSUBS 0.007361f
C238 B.n20 VSUBS 0.007361f
C239 B.n21 VSUBS 0.007361f
C240 B.n22 VSUBS 0.007361f
C241 B.n23 VSUBS 0.007361f
C242 B.n24 VSUBS 0.007361f
C243 B.n25 VSUBS 0.007361f
C244 B.n26 VSUBS 0.007361f
C245 B.n27 VSUBS 0.007361f
C246 B.n28 VSUBS 0.007361f
C247 B.n29 VSUBS 0.007361f
C248 B.n30 VSUBS 0.007361f
C249 B.n31 VSUBS 0.007361f
C250 B.n32 VSUBS 0.007361f
C251 B.n33 VSUBS 0.007361f
C252 B.n34 VSUBS 0.007361f
C253 B.n35 VSUBS 0.007361f
C254 B.t10 VSUBS 0.220037f
C255 B.t11 VSUBS 0.232117f
C256 B.t9 VSUBS 0.345804f
C257 B.n36 VSUBS 0.323809f
C258 B.n37 VSUBS 0.255639f
C259 B.n38 VSUBS 0.007361f
C260 B.n39 VSUBS 0.007361f
C261 B.n40 VSUBS 0.007361f
C262 B.n41 VSUBS 0.007361f
C263 B.t4 VSUBS 0.220041f
C264 B.t5 VSUBS 0.23212f
C265 B.t3 VSUBS 0.345804f
C266 B.n42 VSUBS 0.323806f
C267 B.n43 VSUBS 0.255635f
C268 B.n44 VSUBS 0.017055f
C269 B.n45 VSUBS 0.007361f
C270 B.n46 VSUBS 0.007361f
C271 B.n47 VSUBS 0.007361f
C272 B.n48 VSUBS 0.007361f
C273 B.n49 VSUBS 0.007361f
C274 B.n50 VSUBS 0.007361f
C275 B.n51 VSUBS 0.007361f
C276 B.n52 VSUBS 0.007361f
C277 B.n53 VSUBS 0.007361f
C278 B.n54 VSUBS 0.007361f
C279 B.n55 VSUBS 0.007361f
C280 B.n56 VSUBS 0.007361f
C281 B.n57 VSUBS 0.007361f
C282 B.n58 VSUBS 0.007361f
C283 B.n59 VSUBS 0.007361f
C284 B.n60 VSUBS 0.007361f
C285 B.n61 VSUBS 0.007361f
C286 B.n62 VSUBS 0.007361f
C287 B.n63 VSUBS 0.007361f
C288 B.n64 VSUBS 0.007361f
C289 B.n65 VSUBS 0.018437f
C290 B.n66 VSUBS 0.007361f
C291 B.n67 VSUBS 0.007361f
C292 B.n68 VSUBS 0.007361f
C293 B.n69 VSUBS 0.007361f
C294 B.n70 VSUBS 0.007361f
C295 B.n71 VSUBS 0.007361f
C296 B.n72 VSUBS 0.007361f
C297 B.n73 VSUBS 0.007361f
C298 B.n74 VSUBS 0.007361f
C299 B.n75 VSUBS 0.007361f
C300 B.n76 VSUBS 0.007361f
C301 B.n77 VSUBS 0.007361f
C302 B.n78 VSUBS 0.007361f
C303 B.n79 VSUBS 0.007361f
C304 B.n80 VSUBS 0.007361f
C305 B.n81 VSUBS 0.007361f
C306 B.n82 VSUBS 0.007361f
C307 B.n83 VSUBS 0.007361f
C308 B.n84 VSUBS 0.007361f
C309 B.n85 VSUBS 0.007361f
C310 B.n86 VSUBS 0.007361f
C311 B.n87 VSUBS 0.007361f
C312 B.n88 VSUBS 0.007361f
C313 B.n89 VSUBS 0.007361f
C314 B.n90 VSUBS 0.007361f
C315 B.n91 VSUBS 0.019235f
C316 B.n92 VSUBS 0.007361f
C317 B.n93 VSUBS 0.007361f
C318 B.n94 VSUBS 0.007361f
C319 B.n95 VSUBS 0.007361f
C320 B.n96 VSUBS 0.007361f
C321 B.n97 VSUBS 0.007361f
C322 B.n98 VSUBS 0.007361f
C323 B.n99 VSUBS 0.007361f
C324 B.n100 VSUBS 0.007361f
C325 B.n101 VSUBS 0.007361f
C326 B.n102 VSUBS 0.007361f
C327 B.n103 VSUBS 0.007361f
C328 B.n104 VSUBS 0.007361f
C329 B.n105 VSUBS 0.007361f
C330 B.n106 VSUBS 0.007361f
C331 B.n107 VSUBS 0.007361f
C332 B.n108 VSUBS 0.007361f
C333 B.n109 VSUBS 0.007361f
C334 B.n110 VSUBS 0.007361f
C335 B.n111 VSUBS 0.007361f
C336 B.t2 VSUBS 0.220041f
C337 B.t1 VSUBS 0.23212f
C338 B.t0 VSUBS 0.345804f
C339 B.n112 VSUBS 0.323806f
C340 B.n113 VSUBS 0.255635f
C341 B.n114 VSUBS 0.007361f
C342 B.n115 VSUBS 0.007361f
C343 B.n116 VSUBS 0.007361f
C344 B.n117 VSUBS 0.007361f
C345 B.n118 VSUBS 0.004114f
C346 B.n119 VSUBS 0.007361f
C347 B.n120 VSUBS 0.007361f
C348 B.n121 VSUBS 0.007361f
C349 B.n122 VSUBS 0.007361f
C350 B.n123 VSUBS 0.007361f
C351 B.n124 VSUBS 0.007361f
C352 B.n125 VSUBS 0.007361f
C353 B.n126 VSUBS 0.007361f
C354 B.n127 VSUBS 0.007361f
C355 B.n128 VSUBS 0.007361f
C356 B.n129 VSUBS 0.007361f
C357 B.n130 VSUBS 0.007361f
C358 B.n131 VSUBS 0.007361f
C359 B.n132 VSUBS 0.007361f
C360 B.n133 VSUBS 0.007361f
C361 B.n134 VSUBS 0.007361f
C362 B.n135 VSUBS 0.007361f
C363 B.n136 VSUBS 0.007361f
C364 B.n137 VSUBS 0.007361f
C365 B.n138 VSUBS 0.007361f
C366 B.n139 VSUBS 0.018437f
C367 B.n140 VSUBS 0.007361f
C368 B.n141 VSUBS 0.007361f
C369 B.n142 VSUBS 0.007361f
C370 B.n143 VSUBS 0.007361f
C371 B.n144 VSUBS 0.007361f
C372 B.n145 VSUBS 0.007361f
C373 B.n146 VSUBS 0.007361f
C374 B.n147 VSUBS 0.007361f
C375 B.n148 VSUBS 0.007361f
C376 B.n149 VSUBS 0.007361f
C377 B.n150 VSUBS 0.007361f
C378 B.n151 VSUBS 0.007361f
C379 B.n152 VSUBS 0.007361f
C380 B.n153 VSUBS 0.007361f
C381 B.n154 VSUBS 0.007361f
C382 B.n155 VSUBS 0.007361f
C383 B.n156 VSUBS 0.007361f
C384 B.n157 VSUBS 0.007361f
C385 B.n158 VSUBS 0.007361f
C386 B.n159 VSUBS 0.007361f
C387 B.n160 VSUBS 0.007361f
C388 B.n161 VSUBS 0.007361f
C389 B.n162 VSUBS 0.007361f
C390 B.n163 VSUBS 0.007361f
C391 B.n164 VSUBS 0.007361f
C392 B.n165 VSUBS 0.007361f
C393 B.n166 VSUBS 0.007361f
C394 B.n167 VSUBS 0.007361f
C395 B.n168 VSUBS 0.007361f
C396 B.n169 VSUBS 0.007361f
C397 B.n170 VSUBS 0.007361f
C398 B.n171 VSUBS 0.007361f
C399 B.n172 VSUBS 0.007361f
C400 B.n173 VSUBS 0.007361f
C401 B.n174 VSUBS 0.007361f
C402 B.n175 VSUBS 0.007361f
C403 B.n176 VSUBS 0.007361f
C404 B.n177 VSUBS 0.007361f
C405 B.n178 VSUBS 0.007361f
C406 B.n179 VSUBS 0.007361f
C407 B.n180 VSUBS 0.007361f
C408 B.n181 VSUBS 0.007361f
C409 B.n182 VSUBS 0.007361f
C410 B.n183 VSUBS 0.007361f
C411 B.n184 VSUBS 0.007361f
C412 B.n185 VSUBS 0.007361f
C413 B.n186 VSUBS 0.018437f
C414 B.n187 VSUBS 0.019235f
C415 B.n188 VSUBS 0.019235f
C416 B.n189 VSUBS 0.007361f
C417 B.n190 VSUBS 0.007361f
C418 B.n191 VSUBS 0.007361f
C419 B.n192 VSUBS 0.007361f
C420 B.n193 VSUBS 0.007361f
C421 B.n194 VSUBS 0.007361f
C422 B.n195 VSUBS 0.007361f
C423 B.n196 VSUBS 0.007361f
C424 B.n197 VSUBS 0.007361f
C425 B.n198 VSUBS 0.007361f
C426 B.n199 VSUBS 0.007361f
C427 B.n200 VSUBS 0.007361f
C428 B.n201 VSUBS 0.007361f
C429 B.n202 VSUBS 0.007361f
C430 B.n203 VSUBS 0.007361f
C431 B.n204 VSUBS 0.007361f
C432 B.n205 VSUBS 0.007361f
C433 B.n206 VSUBS 0.007361f
C434 B.n207 VSUBS 0.007361f
C435 B.n208 VSUBS 0.007361f
C436 B.n209 VSUBS 0.007361f
C437 B.n210 VSUBS 0.007361f
C438 B.n211 VSUBS 0.007361f
C439 B.n212 VSUBS 0.007361f
C440 B.n213 VSUBS 0.007361f
C441 B.n214 VSUBS 0.007361f
C442 B.n215 VSUBS 0.007361f
C443 B.n216 VSUBS 0.007361f
C444 B.n217 VSUBS 0.007361f
C445 B.n218 VSUBS 0.007361f
C446 B.n219 VSUBS 0.007361f
C447 B.n220 VSUBS 0.007361f
C448 B.n221 VSUBS 0.007361f
C449 B.n222 VSUBS 0.007361f
C450 B.n223 VSUBS 0.007361f
C451 B.n224 VSUBS 0.007361f
C452 B.n225 VSUBS 0.007361f
C453 B.n226 VSUBS 0.007361f
C454 B.n227 VSUBS 0.007361f
C455 B.n228 VSUBS 0.007361f
C456 B.n229 VSUBS 0.007361f
C457 B.n230 VSUBS 0.007361f
C458 B.n231 VSUBS 0.007361f
C459 B.n232 VSUBS 0.007361f
C460 B.n233 VSUBS 0.007361f
C461 B.n234 VSUBS 0.007361f
C462 B.n235 VSUBS 0.007361f
C463 B.n236 VSUBS 0.007361f
C464 B.n237 VSUBS 0.007361f
C465 B.n238 VSUBS 0.007361f
C466 B.n239 VSUBS 0.007361f
C467 B.n240 VSUBS 0.007361f
C468 B.n241 VSUBS 0.007361f
C469 B.n242 VSUBS 0.007361f
C470 B.n243 VSUBS 0.007361f
C471 B.n244 VSUBS 0.007361f
C472 B.n245 VSUBS 0.007361f
C473 B.n246 VSUBS 0.007361f
C474 B.t8 VSUBS 0.220037f
C475 B.t7 VSUBS 0.232117f
C476 B.t6 VSUBS 0.345804f
C477 B.n247 VSUBS 0.323809f
C478 B.n248 VSUBS 0.255639f
C479 B.n249 VSUBS 0.017055f
C480 B.n250 VSUBS 0.006928f
C481 B.n251 VSUBS 0.007361f
C482 B.n252 VSUBS 0.007361f
C483 B.n253 VSUBS 0.007361f
C484 B.n254 VSUBS 0.007361f
C485 B.n255 VSUBS 0.007361f
C486 B.n256 VSUBS 0.007361f
C487 B.n257 VSUBS 0.007361f
C488 B.n258 VSUBS 0.007361f
C489 B.n259 VSUBS 0.007361f
C490 B.n260 VSUBS 0.007361f
C491 B.n261 VSUBS 0.007361f
C492 B.n262 VSUBS 0.007361f
C493 B.n263 VSUBS 0.007361f
C494 B.n264 VSUBS 0.007361f
C495 B.n265 VSUBS 0.007361f
C496 B.n266 VSUBS 0.004114f
C497 B.n267 VSUBS 0.017055f
C498 B.n268 VSUBS 0.006928f
C499 B.n269 VSUBS 0.007361f
C500 B.n270 VSUBS 0.007361f
C501 B.n271 VSUBS 0.007361f
C502 B.n272 VSUBS 0.007361f
C503 B.n273 VSUBS 0.007361f
C504 B.n274 VSUBS 0.007361f
C505 B.n275 VSUBS 0.007361f
C506 B.n276 VSUBS 0.007361f
C507 B.n277 VSUBS 0.007361f
C508 B.n278 VSUBS 0.007361f
C509 B.n279 VSUBS 0.007361f
C510 B.n280 VSUBS 0.007361f
C511 B.n281 VSUBS 0.007361f
C512 B.n282 VSUBS 0.007361f
C513 B.n283 VSUBS 0.007361f
C514 B.n284 VSUBS 0.007361f
C515 B.n285 VSUBS 0.007361f
C516 B.n286 VSUBS 0.007361f
C517 B.n287 VSUBS 0.007361f
C518 B.n288 VSUBS 0.007361f
C519 B.n289 VSUBS 0.007361f
C520 B.n290 VSUBS 0.007361f
C521 B.n291 VSUBS 0.007361f
C522 B.n292 VSUBS 0.007361f
C523 B.n293 VSUBS 0.007361f
C524 B.n294 VSUBS 0.007361f
C525 B.n295 VSUBS 0.007361f
C526 B.n296 VSUBS 0.007361f
C527 B.n297 VSUBS 0.007361f
C528 B.n298 VSUBS 0.007361f
C529 B.n299 VSUBS 0.007361f
C530 B.n300 VSUBS 0.007361f
C531 B.n301 VSUBS 0.007361f
C532 B.n302 VSUBS 0.007361f
C533 B.n303 VSUBS 0.007361f
C534 B.n304 VSUBS 0.007361f
C535 B.n305 VSUBS 0.007361f
C536 B.n306 VSUBS 0.007361f
C537 B.n307 VSUBS 0.007361f
C538 B.n308 VSUBS 0.007361f
C539 B.n309 VSUBS 0.007361f
C540 B.n310 VSUBS 0.007361f
C541 B.n311 VSUBS 0.007361f
C542 B.n312 VSUBS 0.007361f
C543 B.n313 VSUBS 0.007361f
C544 B.n314 VSUBS 0.007361f
C545 B.n315 VSUBS 0.007361f
C546 B.n316 VSUBS 0.007361f
C547 B.n317 VSUBS 0.007361f
C548 B.n318 VSUBS 0.007361f
C549 B.n319 VSUBS 0.007361f
C550 B.n320 VSUBS 0.007361f
C551 B.n321 VSUBS 0.007361f
C552 B.n322 VSUBS 0.007361f
C553 B.n323 VSUBS 0.007361f
C554 B.n324 VSUBS 0.007361f
C555 B.n325 VSUBS 0.007361f
C556 B.n326 VSUBS 0.007361f
C557 B.n327 VSUBS 0.007361f
C558 B.n328 VSUBS 0.018474f
C559 B.n329 VSUBS 0.019198f
C560 B.n330 VSUBS 0.018437f
C561 B.n331 VSUBS 0.007361f
C562 B.n332 VSUBS 0.007361f
C563 B.n333 VSUBS 0.007361f
C564 B.n334 VSUBS 0.007361f
C565 B.n335 VSUBS 0.007361f
C566 B.n336 VSUBS 0.007361f
C567 B.n337 VSUBS 0.007361f
C568 B.n338 VSUBS 0.007361f
C569 B.n339 VSUBS 0.007361f
C570 B.n340 VSUBS 0.007361f
C571 B.n341 VSUBS 0.007361f
C572 B.n342 VSUBS 0.007361f
C573 B.n343 VSUBS 0.007361f
C574 B.n344 VSUBS 0.007361f
C575 B.n345 VSUBS 0.007361f
C576 B.n346 VSUBS 0.007361f
C577 B.n347 VSUBS 0.007361f
C578 B.n348 VSUBS 0.007361f
C579 B.n349 VSUBS 0.007361f
C580 B.n350 VSUBS 0.007361f
C581 B.n351 VSUBS 0.007361f
C582 B.n352 VSUBS 0.007361f
C583 B.n353 VSUBS 0.007361f
C584 B.n354 VSUBS 0.007361f
C585 B.n355 VSUBS 0.007361f
C586 B.n356 VSUBS 0.007361f
C587 B.n357 VSUBS 0.007361f
C588 B.n358 VSUBS 0.007361f
C589 B.n359 VSUBS 0.007361f
C590 B.n360 VSUBS 0.007361f
C591 B.n361 VSUBS 0.007361f
C592 B.n362 VSUBS 0.007361f
C593 B.n363 VSUBS 0.007361f
C594 B.n364 VSUBS 0.007361f
C595 B.n365 VSUBS 0.007361f
C596 B.n366 VSUBS 0.007361f
C597 B.n367 VSUBS 0.007361f
C598 B.n368 VSUBS 0.007361f
C599 B.n369 VSUBS 0.007361f
C600 B.n370 VSUBS 0.007361f
C601 B.n371 VSUBS 0.007361f
C602 B.n372 VSUBS 0.007361f
C603 B.n373 VSUBS 0.007361f
C604 B.n374 VSUBS 0.007361f
C605 B.n375 VSUBS 0.007361f
C606 B.n376 VSUBS 0.007361f
C607 B.n377 VSUBS 0.007361f
C608 B.n378 VSUBS 0.007361f
C609 B.n379 VSUBS 0.007361f
C610 B.n380 VSUBS 0.007361f
C611 B.n381 VSUBS 0.007361f
C612 B.n382 VSUBS 0.007361f
C613 B.n383 VSUBS 0.007361f
C614 B.n384 VSUBS 0.007361f
C615 B.n385 VSUBS 0.007361f
C616 B.n386 VSUBS 0.007361f
C617 B.n387 VSUBS 0.007361f
C618 B.n388 VSUBS 0.007361f
C619 B.n389 VSUBS 0.007361f
C620 B.n390 VSUBS 0.007361f
C621 B.n391 VSUBS 0.007361f
C622 B.n392 VSUBS 0.007361f
C623 B.n393 VSUBS 0.007361f
C624 B.n394 VSUBS 0.007361f
C625 B.n395 VSUBS 0.007361f
C626 B.n396 VSUBS 0.007361f
C627 B.n397 VSUBS 0.007361f
C628 B.n398 VSUBS 0.007361f
C629 B.n399 VSUBS 0.007361f
C630 B.n400 VSUBS 0.007361f
C631 B.n401 VSUBS 0.007361f
C632 B.n402 VSUBS 0.007361f
C633 B.n403 VSUBS 0.007361f
C634 B.n404 VSUBS 0.007361f
C635 B.n405 VSUBS 0.007361f
C636 B.n406 VSUBS 0.018437f
C637 B.n407 VSUBS 0.019235f
C638 B.n408 VSUBS 0.019235f
C639 B.n409 VSUBS 0.007361f
C640 B.n410 VSUBS 0.007361f
C641 B.n411 VSUBS 0.007361f
C642 B.n412 VSUBS 0.007361f
C643 B.n413 VSUBS 0.007361f
C644 B.n414 VSUBS 0.007361f
C645 B.n415 VSUBS 0.007361f
C646 B.n416 VSUBS 0.007361f
C647 B.n417 VSUBS 0.007361f
C648 B.n418 VSUBS 0.007361f
C649 B.n419 VSUBS 0.007361f
C650 B.n420 VSUBS 0.007361f
C651 B.n421 VSUBS 0.007361f
C652 B.n422 VSUBS 0.007361f
C653 B.n423 VSUBS 0.007361f
C654 B.n424 VSUBS 0.007361f
C655 B.n425 VSUBS 0.007361f
C656 B.n426 VSUBS 0.007361f
C657 B.n427 VSUBS 0.007361f
C658 B.n428 VSUBS 0.007361f
C659 B.n429 VSUBS 0.007361f
C660 B.n430 VSUBS 0.007361f
C661 B.n431 VSUBS 0.007361f
C662 B.n432 VSUBS 0.007361f
C663 B.n433 VSUBS 0.007361f
C664 B.n434 VSUBS 0.007361f
C665 B.n435 VSUBS 0.007361f
C666 B.n436 VSUBS 0.007361f
C667 B.n437 VSUBS 0.007361f
C668 B.n438 VSUBS 0.007361f
C669 B.n439 VSUBS 0.007361f
C670 B.n440 VSUBS 0.007361f
C671 B.n441 VSUBS 0.007361f
C672 B.n442 VSUBS 0.007361f
C673 B.n443 VSUBS 0.007361f
C674 B.n444 VSUBS 0.007361f
C675 B.n445 VSUBS 0.007361f
C676 B.n446 VSUBS 0.007361f
C677 B.n447 VSUBS 0.007361f
C678 B.n448 VSUBS 0.007361f
C679 B.n449 VSUBS 0.007361f
C680 B.n450 VSUBS 0.007361f
C681 B.n451 VSUBS 0.007361f
C682 B.n452 VSUBS 0.007361f
C683 B.n453 VSUBS 0.007361f
C684 B.n454 VSUBS 0.007361f
C685 B.n455 VSUBS 0.007361f
C686 B.n456 VSUBS 0.007361f
C687 B.n457 VSUBS 0.007361f
C688 B.n458 VSUBS 0.007361f
C689 B.n459 VSUBS 0.007361f
C690 B.n460 VSUBS 0.007361f
C691 B.n461 VSUBS 0.007361f
C692 B.n462 VSUBS 0.007361f
C693 B.n463 VSUBS 0.007361f
C694 B.n464 VSUBS 0.007361f
C695 B.n465 VSUBS 0.007361f
C696 B.n466 VSUBS 0.007361f
C697 B.n467 VSUBS 0.006928f
C698 B.n468 VSUBS 0.007361f
C699 B.n469 VSUBS 0.007361f
C700 B.n470 VSUBS 0.004114f
C701 B.n471 VSUBS 0.007361f
C702 B.n472 VSUBS 0.007361f
C703 B.n473 VSUBS 0.007361f
C704 B.n474 VSUBS 0.007361f
C705 B.n475 VSUBS 0.007361f
C706 B.n476 VSUBS 0.007361f
C707 B.n477 VSUBS 0.007361f
C708 B.n478 VSUBS 0.007361f
C709 B.n479 VSUBS 0.007361f
C710 B.n480 VSUBS 0.007361f
C711 B.n481 VSUBS 0.007361f
C712 B.n482 VSUBS 0.007361f
C713 B.n483 VSUBS 0.004114f
C714 B.n484 VSUBS 0.017055f
C715 B.n485 VSUBS 0.006928f
C716 B.n486 VSUBS 0.007361f
C717 B.n487 VSUBS 0.007361f
C718 B.n488 VSUBS 0.007361f
C719 B.n489 VSUBS 0.007361f
C720 B.n490 VSUBS 0.007361f
C721 B.n491 VSUBS 0.007361f
C722 B.n492 VSUBS 0.007361f
C723 B.n493 VSUBS 0.007361f
C724 B.n494 VSUBS 0.007361f
C725 B.n495 VSUBS 0.007361f
C726 B.n496 VSUBS 0.007361f
C727 B.n497 VSUBS 0.007361f
C728 B.n498 VSUBS 0.007361f
C729 B.n499 VSUBS 0.007361f
C730 B.n500 VSUBS 0.007361f
C731 B.n501 VSUBS 0.007361f
C732 B.n502 VSUBS 0.007361f
C733 B.n503 VSUBS 0.007361f
C734 B.n504 VSUBS 0.007361f
C735 B.n505 VSUBS 0.007361f
C736 B.n506 VSUBS 0.007361f
C737 B.n507 VSUBS 0.007361f
C738 B.n508 VSUBS 0.007361f
C739 B.n509 VSUBS 0.007361f
C740 B.n510 VSUBS 0.007361f
C741 B.n511 VSUBS 0.007361f
C742 B.n512 VSUBS 0.007361f
C743 B.n513 VSUBS 0.007361f
C744 B.n514 VSUBS 0.007361f
C745 B.n515 VSUBS 0.007361f
C746 B.n516 VSUBS 0.007361f
C747 B.n517 VSUBS 0.007361f
C748 B.n518 VSUBS 0.007361f
C749 B.n519 VSUBS 0.007361f
C750 B.n520 VSUBS 0.007361f
C751 B.n521 VSUBS 0.007361f
C752 B.n522 VSUBS 0.007361f
C753 B.n523 VSUBS 0.007361f
C754 B.n524 VSUBS 0.007361f
C755 B.n525 VSUBS 0.007361f
C756 B.n526 VSUBS 0.007361f
C757 B.n527 VSUBS 0.007361f
C758 B.n528 VSUBS 0.007361f
C759 B.n529 VSUBS 0.007361f
C760 B.n530 VSUBS 0.007361f
C761 B.n531 VSUBS 0.007361f
C762 B.n532 VSUBS 0.007361f
C763 B.n533 VSUBS 0.007361f
C764 B.n534 VSUBS 0.007361f
C765 B.n535 VSUBS 0.007361f
C766 B.n536 VSUBS 0.007361f
C767 B.n537 VSUBS 0.007361f
C768 B.n538 VSUBS 0.007361f
C769 B.n539 VSUBS 0.007361f
C770 B.n540 VSUBS 0.007361f
C771 B.n541 VSUBS 0.007361f
C772 B.n542 VSUBS 0.007361f
C773 B.n543 VSUBS 0.007361f
C774 B.n544 VSUBS 0.007361f
C775 B.n545 VSUBS 0.019235f
C776 B.n546 VSUBS 0.019235f
C777 B.n547 VSUBS 0.018437f
C778 B.n548 VSUBS 0.007361f
C779 B.n549 VSUBS 0.007361f
C780 B.n550 VSUBS 0.007361f
C781 B.n551 VSUBS 0.007361f
C782 B.n552 VSUBS 0.007361f
C783 B.n553 VSUBS 0.007361f
C784 B.n554 VSUBS 0.007361f
C785 B.n555 VSUBS 0.007361f
C786 B.n556 VSUBS 0.007361f
C787 B.n557 VSUBS 0.007361f
C788 B.n558 VSUBS 0.007361f
C789 B.n559 VSUBS 0.007361f
C790 B.n560 VSUBS 0.007361f
C791 B.n561 VSUBS 0.007361f
C792 B.n562 VSUBS 0.007361f
C793 B.n563 VSUBS 0.007361f
C794 B.n564 VSUBS 0.007361f
C795 B.n565 VSUBS 0.007361f
C796 B.n566 VSUBS 0.007361f
C797 B.n567 VSUBS 0.007361f
C798 B.n568 VSUBS 0.007361f
C799 B.n569 VSUBS 0.007361f
C800 B.n570 VSUBS 0.007361f
C801 B.n571 VSUBS 0.007361f
C802 B.n572 VSUBS 0.007361f
C803 B.n573 VSUBS 0.007361f
C804 B.n574 VSUBS 0.007361f
C805 B.n575 VSUBS 0.007361f
C806 B.n576 VSUBS 0.007361f
C807 B.n577 VSUBS 0.007361f
C808 B.n578 VSUBS 0.007361f
C809 B.n579 VSUBS 0.007361f
C810 B.n580 VSUBS 0.007361f
C811 B.n581 VSUBS 0.007361f
C812 B.n582 VSUBS 0.007361f
C813 B.n583 VSUBS 0.009606f
C814 B.n584 VSUBS 0.010233f
C815 B.n585 VSUBS 0.020349f
C816 VDD2.n0 VSUBS 0.01531f
C817 VDD2.n1 VSUBS 0.034531f
C818 VDD2.n2 VSUBS 0.015469f
C819 VDD2.n3 VSUBS 0.027188f
C820 VDD2.n4 VSUBS 0.014609f
C821 VDD2.n5 VSUBS 0.034531f
C822 VDD2.n6 VSUBS 0.015469f
C823 VDD2.n7 VSUBS 0.027188f
C824 VDD2.n8 VSUBS 0.014609f
C825 VDD2.n9 VSUBS 0.034531f
C826 VDD2.n10 VSUBS 0.015469f
C827 VDD2.n11 VSUBS 0.027188f
C828 VDD2.n12 VSUBS 0.014609f
C829 VDD2.n13 VSUBS 0.034531f
C830 VDD2.n14 VSUBS 0.015469f
C831 VDD2.n15 VSUBS 0.027188f
C832 VDD2.n16 VSUBS 0.014609f
C833 VDD2.n17 VSUBS 0.034531f
C834 VDD2.n18 VSUBS 0.015469f
C835 VDD2.n19 VSUBS 1.35706f
C836 VDD2.n20 VSUBS 0.014609f
C837 VDD2.t0 VSUBS 0.073721f
C838 VDD2.n21 VSUBS 0.167034f
C839 VDD2.n22 VSUBS 0.021967f
C840 VDD2.n23 VSUBS 0.025899f
C841 VDD2.n24 VSUBS 0.034531f
C842 VDD2.n25 VSUBS 0.015469f
C843 VDD2.n26 VSUBS 0.014609f
C844 VDD2.n27 VSUBS 0.027188f
C845 VDD2.n28 VSUBS 0.027188f
C846 VDD2.n29 VSUBS 0.014609f
C847 VDD2.n30 VSUBS 0.015469f
C848 VDD2.n31 VSUBS 0.034531f
C849 VDD2.n32 VSUBS 0.034531f
C850 VDD2.n33 VSUBS 0.015469f
C851 VDD2.n34 VSUBS 0.014609f
C852 VDD2.n35 VSUBS 0.027188f
C853 VDD2.n36 VSUBS 0.027188f
C854 VDD2.n37 VSUBS 0.014609f
C855 VDD2.n38 VSUBS 0.015469f
C856 VDD2.n39 VSUBS 0.034531f
C857 VDD2.n40 VSUBS 0.034531f
C858 VDD2.n41 VSUBS 0.015469f
C859 VDD2.n42 VSUBS 0.014609f
C860 VDD2.n43 VSUBS 0.027188f
C861 VDD2.n44 VSUBS 0.027188f
C862 VDD2.n45 VSUBS 0.014609f
C863 VDD2.n46 VSUBS 0.015469f
C864 VDD2.n47 VSUBS 0.034531f
C865 VDD2.n48 VSUBS 0.034531f
C866 VDD2.n49 VSUBS 0.015469f
C867 VDD2.n50 VSUBS 0.014609f
C868 VDD2.n51 VSUBS 0.027188f
C869 VDD2.n52 VSUBS 0.027188f
C870 VDD2.n53 VSUBS 0.014609f
C871 VDD2.n54 VSUBS 0.015469f
C872 VDD2.n55 VSUBS 0.034531f
C873 VDD2.n56 VSUBS 0.034531f
C874 VDD2.n57 VSUBS 0.015469f
C875 VDD2.n58 VSUBS 0.014609f
C876 VDD2.n59 VSUBS 0.027188f
C877 VDD2.n60 VSUBS 0.069157f
C878 VDD2.n61 VSUBS 0.014609f
C879 VDD2.n62 VSUBS 0.015469f
C880 VDD2.n63 VSUBS 0.075751f
C881 VDD2.n64 VSUBS 0.071502f
C882 VDD2.t2 VSUBS 0.256309f
C883 VDD2.t4 VSUBS 0.256309f
C884 VDD2.n65 VSUBS 2.02117f
C885 VDD2.n66 VSUBS 0.708364f
C886 VDD2.t6 VSUBS 0.256309f
C887 VDD2.t8 VSUBS 0.256309f
C888 VDD2.n67 VSUBS 2.02596f
C889 VDD2.n68 VSUBS 2.3093f
C890 VDD2.n69 VSUBS 0.01531f
C891 VDD2.n70 VSUBS 0.034531f
C892 VDD2.n71 VSUBS 0.015469f
C893 VDD2.n72 VSUBS 0.027188f
C894 VDD2.n73 VSUBS 0.014609f
C895 VDD2.n74 VSUBS 0.034531f
C896 VDD2.n75 VSUBS 0.015469f
C897 VDD2.n76 VSUBS 0.027188f
C898 VDD2.n77 VSUBS 0.014609f
C899 VDD2.n78 VSUBS 0.034531f
C900 VDD2.n79 VSUBS 0.015469f
C901 VDD2.n80 VSUBS 0.027188f
C902 VDD2.n81 VSUBS 0.014609f
C903 VDD2.n82 VSUBS 0.034531f
C904 VDD2.n83 VSUBS 0.015469f
C905 VDD2.n84 VSUBS 0.027188f
C906 VDD2.n85 VSUBS 0.014609f
C907 VDD2.n86 VSUBS 0.034531f
C908 VDD2.n87 VSUBS 0.015469f
C909 VDD2.n88 VSUBS 1.35706f
C910 VDD2.n89 VSUBS 0.014609f
C911 VDD2.t9 VSUBS 0.073721f
C912 VDD2.n90 VSUBS 0.167034f
C913 VDD2.n91 VSUBS 0.021967f
C914 VDD2.n92 VSUBS 0.025899f
C915 VDD2.n93 VSUBS 0.034531f
C916 VDD2.n94 VSUBS 0.015469f
C917 VDD2.n95 VSUBS 0.014609f
C918 VDD2.n96 VSUBS 0.027188f
C919 VDD2.n97 VSUBS 0.027188f
C920 VDD2.n98 VSUBS 0.014609f
C921 VDD2.n99 VSUBS 0.015469f
C922 VDD2.n100 VSUBS 0.034531f
C923 VDD2.n101 VSUBS 0.034531f
C924 VDD2.n102 VSUBS 0.015469f
C925 VDD2.n103 VSUBS 0.014609f
C926 VDD2.n104 VSUBS 0.027188f
C927 VDD2.n105 VSUBS 0.027188f
C928 VDD2.n106 VSUBS 0.014609f
C929 VDD2.n107 VSUBS 0.015469f
C930 VDD2.n108 VSUBS 0.034531f
C931 VDD2.n109 VSUBS 0.034531f
C932 VDD2.n110 VSUBS 0.015469f
C933 VDD2.n111 VSUBS 0.014609f
C934 VDD2.n112 VSUBS 0.027188f
C935 VDD2.n113 VSUBS 0.027188f
C936 VDD2.n114 VSUBS 0.014609f
C937 VDD2.n115 VSUBS 0.015469f
C938 VDD2.n116 VSUBS 0.034531f
C939 VDD2.n117 VSUBS 0.034531f
C940 VDD2.n118 VSUBS 0.015469f
C941 VDD2.n119 VSUBS 0.014609f
C942 VDD2.n120 VSUBS 0.027188f
C943 VDD2.n121 VSUBS 0.027188f
C944 VDD2.n122 VSUBS 0.014609f
C945 VDD2.n123 VSUBS 0.015469f
C946 VDD2.n124 VSUBS 0.034531f
C947 VDD2.n125 VSUBS 0.034531f
C948 VDD2.n126 VSUBS 0.015469f
C949 VDD2.n127 VSUBS 0.014609f
C950 VDD2.n128 VSUBS 0.027188f
C951 VDD2.n129 VSUBS 0.069157f
C952 VDD2.n130 VSUBS 0.014609f
C953 VDD2.n131 VSUBS 0.015469f
C954 VDD2.n132 VSUBS 0.075751f
C955 VDD2.n133 VSUBS 0.069337f
C956 VDD2.n134 VSUBS 2.32698f
C957 VDD2.t3 VSUBS 0.256309f
C958 VDD2.t7 VSUBS 0.256309f
C959 VDD2.n135 VSUBS 2.02118f
C960 VDD2.n136 VSUBS 0.58632f
C961 VDD2.t1 VSUBS 0.256309f
C962 VDD2.t5 VSUBS 0.256309f
C963 VDD2.n137 VSUBS 2.02592f
C964 VTAIL.t14 VSUBS 0.277422f
C965 VTAIL.t11 VSUBS 0.277422f
C966 VTAIL.n0 VSUBS 2.04282f
C967 VTAIL.n1 VSUBS 0.784017f
C968 VTAIL.n2 VSUBS 0.016571f
C969 VTAIL.n3 VSUBS 0.037376f
C970 VTAIL.n4 VSUBS 0.016743f
C971 VTAIL.n5 VSUBS 0.029427f
C972 VTAIL.n6 VSUBS 0.015813f
C973 VTAIL.n7 VSUBS 0.037376f
C974 VTAIL.n8 VSUBS 0.016743f
C975 VTAIL.n9 VSUBS 0.029427f
C976 VTAIL.n10 VSUBS 0.015813f
C977 VTAIL.n11 VSUBS 0.037376f
C978 VTAIL.n12 VSUBS 0.016743f
C979 VTAIL.n13 VSUBS 0.029427f
C980 VTAIL.n14 VSUBS 0.015813f
C981 VTAIL.n15 VSUBS 0.037376f
C982 VTAIL.n16 VSUBS 0.016743f
C983 VTAIL.n17 VSUBS 0.029427f
C984 VTAIL.n18 VSUBS 0.015813f
C985 VTAIL.n19 VSUBS 0.037376f
C986 VTAIL.n20 VSUBS 0.016743f
C987 VTAIL.n21 VSUBS 1.46885f
C988 VTAIL.n22 VSUBS 0.015813f
C989 VTAIL.t3 VSUBS 0.079794f
C990 VTAIL.n23 VSUBS 0.180793f
C991 VTAIL.n24 VSUBS 0.023777f
C992 VTAIL.n25 VSUBS 0.028032f
C993 VTAIL.n26 VSUBS 0.037376f
C994 VTAIL.n27 VSUBS 0.016743f
C995 VTAIL.n28 VSUBS 0.015813f
C996 VTAIL.n29 VSUBS 0.029427f
C997 VTAIL.n30 VSUBS 0.029427f
C998 VTAIL.n31 VSUBS 0.015813f
C999 VTAIL.n32 VSUBS 0.016743f
C1000 VTAIL.n33 VSUBS 0.037376f
C1001 VTAIL.n34 VSUBS 0.037376f
C1002 VTAIL.n35 VSUBS 0.016743f
C1003 VTAIL.n36 VSUBS 0.015813f
C1004 VTAIL.n37 VSUBS 0.029427f
C1005 VTAIL.n38 VSUBS 0.029427f
C1006 VTAIL.n39 VSUBS 0.015813f
C1007 VTAIL.n40 VSUBS 0.016743f
C1008 VTAIL.n41 VSUBS 0.037376f
C1009 VTAIL.n42 VSUBS 0.037376f
C1010 VTAIL.n43 VSUBS 0.016743f
C1011 VTAIL.n44 VSUBS 0.015813f
C1012 VTAIL.n45 VSUBS 0.029427f
C1013 VTAIL.n46 VSUBS 0.029427f
C1014 VTAIL.n47 VSUBS 0.015813f
C1015 VTAIL.n48 VSUBS 0.016743f
C1016 VTAIL.n49 VSUBS 0.037376f
C1017 VTAIL.n50 VSUBS 0.037376f
C1018 VTAIL.n51 VSUBS 0.016743f
C1019 VTAIL.n52 VSUBS 0.015813f
C1020 VTAIL.n53 VSUBS 0.029427f
C1021 VTAIL.n54 VSUBS 0.029427f
C1022 VTAIL.n55 VSUBS 0.015813f
C1023 VTAIL.n56 VSUBS 0.016743f
C1024 VTAIL.n57 VSUBS 0.037376f
C1025 VTAIL.n58 VSUBS 0.037376f
C1026 VTAIL.n59 VSUBS 0.016743f
C1027 VTAIL.n60 VSUBS 0.015813f
C1028 VTAIL.n61 VSUBS 0.029427f
C1029 VTAIL.n62 VSUBS 0.074853f
C1030 VTAIL.n63 VSUBS 0.015813f
C1031 VTAIL.n64 VSUBS 0.016743f
C1032 VTAIL.n65 VSUBS 0.081991f
C1033 VTAIL.n66 VSUBS 0.054763f
C1034 VTAIL.n67 VSUBS 0.194795f
C1035 VTAIL.t5 VSUBS 0.277422f
C1036 VTAIL.t19 VSUBS 0.277422f
C1037 VTAIL.n68 VSUBS 2.04282f
C1038 VTAIL.n69 VSUBS 0.795256f
C1039 VTAIL.t6 VSUBS 0.277422f
C1040 VTAIL.t2 VSUBS 0.277422f
C1041 VTAIL.n70 VSUBS 2.04282f
C1042 VTAIL.n71 VSUBS 2.25191f
C1043 VTAIL.t10 VSUBS 0.277422f
C1044 VTAIL.t17 VSUBS 0.277422f
C1045 VTAIL.n72 VSUBS 2.04283f
C1046 VTAIL.n73 VSUBS 2.2519f
C1047 VTAIL.t16 VSUBS 0.277422f
C1048 VTAIL.t8 VSUBS 0.277422f
C1049 VTAIL.n74 VSUBS 2.04283f
C1050 VTAIL.n75 VSUBS 0.795246f
C1051 VTAIL.n76 VSUBS 0.016571f
C1052 VTAIL.n77 VSUBS 0.037376f
C1053 VTAIL.n78 VSUBS 0.016743f
C1054 VTAIL.n79 VSUBS 0.029427f
C1055 VTAIL.n80 VSUBS 0.015813f
C1056 VTAIL.n81 VSUBS 0.037376f
C1057 VTAIL.n82 VSUBS 0.016743f
C1058 VTAIL.n83 VSUBS 0.029427f
C1059 VTAIL.n84 VSUBS 0.015813f
C1060 VTAIL.n85 VSUBS 0.037376f
C1061 VTAIL.n86 VSUBS 0.016743f
C1062 VTAIL.n87 VSUBS 0.029427f
C1063 VTAIL.n88 VSUBS 0.015813f
C1064 VTAIL.n89 VSUBS 0.037376f
C1065 VTAIL.n90 VSUBS 0.016743f
C1066 VTAIL.n91 VSUBS 0.029427f
C1067 VTAIL.n92 VSUBS 0.015813f
C1068 VTAIL.n93 VSUBS 0.037376f
C1069 VTAIL.n94 VSUBS 0.016743f
C1070 VTAIL.n95 VSUBS 1.46885f
C1071 VTAIL.n96 VSUBS 0.015813f
C1072 VTAIL.t9 VSUBS 0.079794f
C1073 VTAIL.n97 VSUBS 0.180793f
C1074 VTAIL.n98 VSUBS 0.023777f
C1075 VTAIL.n99 VSUBS 0.028032f
C1076 VTAIL.n100 VSUBS 0.037376f
C1077 VTAIL.n101 VSUBS 0.016743f
C1078 VTAIL.n102 VSUBS 0.015813f
C1079 VTAIL.n103 VSUBS 0.029427f
C1080 VTAIL.n104 VSUBS 0.029427f
C1081 VTAIL.n105 VSUBS 0.015813f
C1082 VTAIL.n106 VSUBS 0.016743f
C1083 VTAIL.n107 VSUBS 0.037376f
C1084 VTAIL.n108 VSUBS 0.037376f
C1085 VTAIL.n109 VSUBS 0.016743f
C1086 VTAIL.n110 VSUBS 0.015813f
C1087 VTAIL.n111 VSUBS 0.029427f
C1088 VTAIL.n112 VSUBS 0.029427f
C1089 VTAIL.n113 VSUBS 0.015813f
C1090 VTAIL.n114 VSUBS 0.016743f
C1091 VTAIL.n115 VSUBS 0.037376f
C1092 VTAIL.n116 VSUBS 0.037376f
C1093 VTAIL.n117 VSUBS 0.016743f
C1094 VTAIL.n118 VSUBS 0.015813f
C1095 VTAIL.n119 VSUBS 0.029427f
C1096 VTAIL.n120 VSUBS 0.029427f
C1097 VTAIL.n121 VSUBS 0.015813f
C1098 VTAIL.n122 VSUBS 0.016743f
C1099 VTAIL.n123 VSUBS 0.037376f
C1100 VTAIL.n124 VSUBS 0.037376f
C1101 VTAIL.n125 VSUBS 0.016743f
C1102 VTAIL.n126 VSUBS 0.015813f
C1103 VTAIL.n127 VSUBS 0.029427f
C1104 VTAIL.n128 VSUBS 0.029427f
C1105 VTAIL.n129 VSUBS 0.015813f
C1106 VTAIL.n130 VSUBS 0.016743f
C1107 VTAIL.n131 VSUBS 0.037376f
C1108 VTAIL.n132 VSUBS 0.037376f
C1109 VTAIL.n133 VSUBS 0.016743f
C1110 VTAIL.n134 VSUBS 0.015813f
C1111 VTAIL.n135 VSUBS 0.029427f
C1112 VTAIL.n136 VSUBS 0.074853f
C1113 VTAIL.n137 VSUBS 0.015813f
C1114 VTAIL.n138 VSUBS 0.016743f
C1115 VTAIL.n139 VSUBS 0.081991f
C1116 VTAIL.n140 VSUBS 0.054763f
C1117 VTAIL.n141 VSUBS 0.194795f
C1118 VTAIL.t4 VSUBS 0.277422f
C1119 VTAIL.t0 VSUBS 0.277422f
C1120 VTAIL.n142 VSUBS 2.04283f
C1121 VTAIL.n143 VSUBS 0.798924f
C1122 VTAIL.t7 VSUBS 0.277422f
C1123 VTAIL.t18 VSUBS 0.277422f
C1124 VTAIL.n144 VSUBS 2.04283f
C1125 VTAIL.n145 VSUBS 0.795246f
C1126 VTAIL.n146 VSUBS 0.016571f
C1127 VTAIL.n147 VSUBS 0.037376f
C1128 VTAIL.n148 VSUBS 0.016743f
C1129 VTAIL.n149 VSUBS 0.029427f
C1130 VTAIL.n150 VSUBS 0.015813f
C1131 VTAIL.n151 VSUBS 0.037376f
C1132 VTAIL.n152 VSUBS 0.016743f
C1133 VTAIL.n153 VSUBS 0.029427f
C1134 VTAIL.n154 VSUBS 0.015813f
C1135 VTAIL.n155 VSUBS 0.037376f
C1136 VTAIL.n156 VSUBS 0.016743f
C1137 VTAIL.n157 VSUBS 0.029427f
C1138 VTAIL.n158 VSUBS 0.015813f
C1139 VTAIL.n159 VSUBS 0.037376f
C1140 VTAIL.n160 VSUBS 0.016743f
C1141 VTAIL.n161 VSUBS 0.029427f
C1142 VTAIL.n162 VSUBS 0.015813f
C1143 VTAIL.n163 VSUBS 0.037376f
C1144 VTAIL.n164 VSUBS 0.016743f
C1145 VTAIL.n165 VSUBS 1.46885f
C1146 VTAIL.n166 VSUBS 0.015813f
C1147 VTAIL.t1 VSUBS 0.079794f
C1148 VTAIL.n167 VSUBS 0.180793f
C1149 VTAIL.n168 VSUBS 0.023777f
C1150 VTAIL.n169 VSUBS 0.028032f
C1151 VTAIL.n170 VSUBS 0.037376f
C1152 VTAIL.n171 VSUBS 0.016743f
C1153 VTAIL.n172 VSUBS 0.015813f
C1154 VTAIL.n173 VSUBS 0.029427f
C1155 VTAIL.n174 VSUBS 0.029427f
C1156 VTAIL.n175 VSUBS 0.015813f
C1157 VTAIL.n176 VSUBS 0.016743f
C1158 VTAIL.n177 VSUBS 0.037376f
C1159 VTAIL.n178 VSUBS 0.037376f
C1160 VTAIL.n179 VSUBS 0.016743f
C1161 VTAIL.n180 VSUBS 0.015813f
C1162 VTAIL.n181 VSUBS 0.029427f
C1163 VTAIL.n182 VSUBS 0.029427f
C1164 VTAIL.n183 VSUBS 0.015813f
C1165 VTAIL.n184 VSUBS 0.016743f
C1166 VTAIL.n185 VSUBS 0.037376f
C1167 VTAIL.n186 VSUBS 0.037376f
C1168 VTAIL.n187 VSUBS 0.016743f
C1169 VTAIL.n188 VSUBS 0.015813f
C1170 VTAIL.n189 VSUBS 0.029427f
C1171 VTAIL.n190 VSUBS 0.029427f
C1172 VTAIL.n191 VSUBS 0.015813f
C1173 VTAIL.n192 VSUBS 0.016743f
C1174 VTAIL.n193 VSUBS 0.037376f
C1175 VTAIL.n194 VSUBS 0.037376f
C1176 VTAIL.n195 VSUBS 0.016743f
C1177 VTAIL.n196 VSUBS 0.015813f
C1178 VTAIL.n197 VSUBS 0.029427f
C1179 VTAIL.n198 VSUBS 0.029427f
C1180 VTAIL.n199 VSUBS 0.015813f
C1181 VTAIL.n200 VSUBS 0.016743f
C1182 VTAIL.n201 VSUBS 0.037376f
C1183 VTAIL.n202 VSUBS 0.037376f
C1184 VTAIL.n203 VSUBS 0.016743f
C1185 VTAIL.n204 VSUBS 0.015813f
C1186 VTAIL.n205 VSUBS 0.029427f
C1187 VTAIL.n206 VSUBS 0.074853f
C1188 VTAIL.n207 VSUBS 0.015813f
C1189 VTAIL.n208 VSUBS 0.016743f
C1190 VTAIL.n209 VSUBS 0.081991f
C1191 VTAIL.n210 VSUBS 0.054763f
C1192 VTAIL.n211 VSUBS 1.56603f
C1193 VTAIL.n212 VSUBS 0.016571f
C1194 VTAIL.n213 VSUBS 0.037376f
C1195 VTAIL.n214 VSUBS 0.016743f
C1196 VTAIL.n215 VSUBS 0.029427f
C1197 VTAIL.n216 VSUBS 0.015813f
C1198 VTAIL.n217 VSUBS 0.037376f
C1199 VTAIL.n218 VSUBS 0.016743f
C1200 VTAIL.n219 VSUBS 0.029427f
C1201 VTAIL.n220 VSUBS 0.015813f
C1202 VTAIL.n221 VSUBS 0.037376f
C1203 VTAIL.n222 VSUBS 0.016743f
C1204 VTAIL.n223 VSUBS 0.029427f
C1205 VTAIL.n224 VSUBS 0.015813f
C1206 VTAIL.n225 VSUBS 0.037376f
C1207 VTAIL.n226 VSUBS 0.016743f
C1208 VTAIL.n227 VSUBS 0.029427f
C1209 VTAIL.n228 VSUBS 0.015813f
C1210 VTAIL.n229 VSUBS 0.037376f
C1211 VTAIL.n230 VSUBS 0.016743f
C1212 VTAIL.n231 VSUBS 1.46885f
C1213 VTAIL.n232 VSUBS 0.015813f
C1214 VTAIL.t15 VSUBS 0.079794f
C1215 VTAIL.n233 VSUBS 0.180793f
C1216 VTAIL.n234 VSUBS 0.023777f
C1217 VTAIL.n235 VSUBS 0.028032f
C1218 VTAIL.n236 VSUBS 0.037376f
C1219 VTAIL.n237 VSUBS 0.016743f
C1220 VTAIL.n238 VSUBS 0.015813f
C1221 VTAIL.n239 VSUBS 0.029427f
C1222 VTAIL.n240 VSUBS 0.029427f
C1223 VTAIL.n241 VSUBS 0.015813f
C1224 VTAIL.n242 VSUBS 0.016743f
C1225 VTAIL.n243 VSUBS 0.037376f
C1226 VTAIL.n244 VSUBS 0.037376f
C1227 VTAIL.n245 VSUBS 0.016743f
C1228 VTAIL.n246 VSUBS 0.015813f
C1229 VTAIL.n247 VSUBS 0.029427f
C1230 VTAIL.n248 VSUBS 0.029427f
C1231 VTAIL.n249 VSUBS 0.015813f
C1232 VTAIL.n250 VSUBS 0.016743f
C1233 VTAIL.n251 VSUBS 0.037376f
C1234 VTAIL.n252 VSUBS 0.037376f
C1235 VTAIL.n253 VSUBS 0.016743f
C1236 VTAIL.n254 VSUBS 0.015813f
C1237 VTAIL.n255 VSUBS 0.029427f
C1238 VTAIL.n256 VSUBS 0.029427f
C1239 VTAIL.n257 VSUBS 0.015813f
C1240 VTAIL.n258 VSUBS 0.016743f
C1241 VTAIL.n259 VSUBS 0.037376f
C1242 VTAIL.n260 VSUBS 0.037376f
C1243 VTAIL.n261 VSUBS 0.016743f
C1244 VTAIL.n262 VSUBS 0.015813f
C1245 VTAIL.n263 VSUBS 0.029427f
C1246 VTAIL.n264 VSUBS 0.029427f
C1247 VTAIL.n265 VSUBS 0.015813f
C1248 VTAIL.n266 VSUBS 0.016743f
C1249 VTAIL.n267 VSUBS 0.037376f
C1250 VTAIL.n268 VSUBS 0.037376f
C1251 VTAIL.n269 VSUBS 0.016743f
C1252 VTAIL.n270 VSUBS 0.015813f
C1253 VTAIL.n271 VSUBS 0.029427f
C1254 VTAIL.n272 VSUBS 0.074853f
C1255 VTAIL.n273 VSUBS 0.015813f
C1256 VTAIL.n274 VSUBS 0.016743f
C1257 VTAIL.n275 VSUBS 0.081991f
C1258 VTAIL.n276 VSUBS 0.054763f
C1259 VTAIL.n277 VSUBS 1.56603f
C1260 VTAIL.t13 VSUBS 0.277422f
C1261 VTAIL.t12 VSUBS 0.277422f
C1262 VTAIL.n278 VSUBS 2.04282f
C1263 VTAIL.n279 VSUBS 0.728432f
C1264 VN.n0 VSUBS 0.052898f
C1265 VN.n1 VSUBS 0.012004f
C1266 VN.n2 VSUBS 0.216097f
C1267 VN.t9 VSUBS 1.226f
C1268 VN.n3 VSUBS 0.467118f
C1269 VN.t7 VSUBS 1.20613f
C1270 VN.n4 VSUBS 0.486944f
C1271 VN.n5 VSUBS 0.012004f
C1272 VN.t5 VSUBS 1.20613f
C1273 VN.n6 VSUBS 0.483133f
C1274 VN.n7 VSUBS 0.052898f
C1275 VN.n8 VSUBS 0.052898f
C1276 VN.n9 VSUBS 0.052898f
C1277 VN.t3 VSUBS 1.20613f
C1278 VN.n10 VSUBS 0.483133f
C1279 VN.n11 VSUBS 0.012004f
C1280 VN.t1 VSUBS 1.20613f
C1281 VN.n12 VSUBS 0.477752f
C1282 VN.n13 VSUBS 0.040994f
C1283 VN.n14 VSUBS 0.052898f
C1284 VN.n15 VSUBS 0.012004f
C1285 VN.t6 VSUBS 1.20613f
C1286 VN.n16 VSUBS 0.216097f
C1287 VN.t4 VSUBS 1.226f
C1288 VN.n17 VSUBS 0.467118f
C1289 VN.t8 VSUBS 1.20613f
C1290 VN.n18 VSUBS 0.486944f
C1291 VN.n19 VSUBS 0.012004f
C1292 VN.t2 VSUBS 1.20613f
C1293 VN.n20 VSUBS 0.483133f
C1294 VN.n21 VSUBS 0.052898f
C1295 VN.n22 VSUBS 0.052898f
C1296 VN.n23 VSUBS 0.052898f
C1297 VN.n24 VSUBS 0.483133f
C1298 VN.n25 VSUBS 0.012004f
C1299 VN.t0 VSUBS 1.20613f
C1300 VN.n26 VSUBS 0.477752f
C1301 VN.n27 VSUBS 2.26285f
.ends

