* NGSPICE file created from diff_pair_sample_0107.ext - technology: sky130A

.subckt diff_pair_sample_0107 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=0.69
X1 VDD1.t5 VP.t0 VTAIL.t7 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=1.8447 ps=10.24 w=4.73 l=0.69
X2 VDD1.t4 VP.t1 VTAIL.t11 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0.78045 ps=5.06 w=4.73 l=0.69
X3 VDD2.t5 VN.t0 VTAIL.t4 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=1.8447 ps=10.24 w=4.73 l=0.69
X4 VDD2.t4 VN.t1 VTAIL.t5 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0.78045 ps=5.06 w=4.73 l=0.69
X5 B.t8 B.t6 B.t7 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=0.69
X6 VDD2.t3 VN.t2 VTAIL.t0 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=1.8447 ps=10.24 w=4.73 l=0.69
X7 VTAIL.t1 VN.t3 VDD2.t2 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=0.78045 ps=5.06 w=4.73 l=0.69
X8 VTAIL.t3 VN.t4 VDD2.t1 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=0.78045 ps=5.06 w=4.73 l=0.69
X9 VDD2.t0 VN.t5 VTAIL.t2 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0.78045 ps=5.06 w=4.73 l=0.69
X10 VDD1.t3 VP.t2 VTAIL.t6 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0.78045 ps=5.06 w=4.73 l=0.69
X11 B.t5 B.t3 B.t4 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=0.69
X12 B.t2 B.t0 B.t1 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=1.8447 pd=10.24 as=0 ps=0 w=4.73 l=0.69
X13 VTAIL.t10 VP.t3 VDD1.t2 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=0.78045 ps=5.06 w=4.73 l=0.69
X14 VTAIL.t9 VP.t4 VDD1.t1 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=0.78045 ps=5.06 w=4.73 l=0.69
X15 VDD1.t0 VP.t5 VTAIL.t8 w_n1786_n1914# sky130_fd_pr__pfet_01v8 ad=0.78045 pd=5.06 as=1.8447 ps=10.24 w=4.73 l=0.69
R0 B.n268 B.n41 585
R1 B.n270 B.n269 585
R2 B.n271 B.n40 585
R3 B.n273 B.n272 585
R4 B.n274 B.n39 585
R5 B.n276 B.n275 585
R6 B.n277 B.n38 585
R7 B.n279 B.n278 585
R8 B.n280 B.n37 585
R9 B.n282 B.n281 585
R10 B.n283 B.n36 585
R11 B.n285 B.n284 585
R12 B.n286 B.n35 585
R13 B.n288 B.n287 585
R14 B.n289 B.n34 585
R15 B.n291 B.n290 585
R16 B.n292 B.n33 585
R17 B.n294 B.n293 585
R18 B.n295 B.n32 585
R19 B.n297 B.n296 585
R20 B.n299 B.n29 585
R21 B.n301 B.n300 585
R22 B.n302 B.n28 585
R23 B.n304 B.n303 585
R24 B.n305 B.n27 585
R25 B.n307 B.n306 585
R26 B.n308 B.n26 585
R27 B.n310 B.n309 585
R28 B.n311 B.n25 585
R29 B.n313 B.n312 585
R30 B.n315 B.n314 585
R31 B.n316 B.n21 585
R32 B.n318 B.n317 585
R33 B.n319 B.n20 585
R34 B.n321 B.n320 585
R35 B.n322 B.n19 585
R36 B.n324 B.n323 585
R37 B.n325 B.n18 585
R38 B.n327 B.n326 585
R39 B.n328 B.n17 585
R40 B.n330 B.n329 585
R41 B.n331 B.n16 585
R42 B.n333 B.n332 585
R43 B.n334 B.n15 585
R44 B.n336 B.n335 585
R45 B.n337 B.n14 585
R46 B.n339 B.n338 585
R47 B.n340 B.n13 585
R48 B.n342 B.n341 585
R49 B.n343 B.n12 585
R50 B.n267 B.n266 585
R51 B.n265 B.n42 585
R52 B.n264 B.n263 585
R53 B.n262 B.n43 585
R54 B.n261 B.n260 585
R55 B.n259 B.n44 585
R56 B.n258 B.n257 585
R57 B.n256 B.n45 585
R58 B.n255 B.n254 585
R59 B.n253 B.n46 585
R60 B.n252 B.n251 585
R61 B.n250 B.n47 585
R62 B.n249 B.n248 585
R63 B.n247 B.n48 585
R64 B.n246 B.n245 585
R65 B.n244 B.n49 585
R66 B.n243 B.n242 585
R67 B.n241 B.n50 585
R68 B.n240 B.n239 585
R69 B.n238 B.n51 585
R70 B.n237 B.n236 585
R71 B.n235 B.n52 585
R72 B.n234 B.n233 585
R73 B.n232 B.n53 585
R74 B.n231 B.n230 585
R75 B.n229 B.n54 585
R76 B.n228 B.n227 585
R77 B.n226 B.n55 585
R78 B.n225 B.n224 585
R79 B.n223 B.n56 585
R80 B.n222 B.n221 585
R81 B.n220 B.n57 585
R82 B.n219 B.n218 585
R83 B.n217 B.n58 585
R84 B.n216 B.n215 585
R85 B.n214 B.n59 585
R86 B.n213 B.n212 585
R87 B.n211 B.n60 585
R88 B.n210 B.n209 585
R89 B.n208 B.n61 585
R90 B.n207 B.n206 585
R91 B.n130 B.n91 585
R92 B.n132 B.n131 585
R93 B.n133 B.n90 585
R94 B.n135 B.n134 585
R95 B.n136 B.n89 585
R96 B.n138 B.n137 585
R97 B.n139 B.n88 585
R98 B.n141 B.n140 585
R99 B.n142 B.n87 585
R100 B.n144 B.n143 585
R101 B.n145 B.n86 585
R102 B.n147 B.n146 585
R103 B.n148 B.n85 585
R104 B.n150 B.n149 585
R105 B.n151 B.n84 585
R106 B.n153 B.n152 585
R107 B.n154 B.n83 585
R108 B.n156 B.n155 585
R109 B.n157 B.n82 585
R110 B.n159 B.n158 585
R111 B.n161 B.n79 585
R112 B.n163 B.n162 585
R113 B.n164 B.n78 585
R114 B.n166 B.n165 585
R115 B.n167 B.n77 585
R116 B.n169 B.n168 585
R117 B.n170 B.n76 585
R118 B.n172 B.n171 585
R119 B.n173 B.n75 585
R120 B.n175 B.n174 585
R121 B.n177 B.n176 585
R122 B.n178 B.n71 585
R123 B.n180 B.n179 585
R124 B.n181 B.n70 585
R125 B.n183 B.n182 585
R126 B.n184 B.n69 585
R127 B.n186 B.n185 585
R128 B.n187 B.n68 585
R129 B.n189 B.n188 585
R130 B.n190 B.n67 585
R131 B.n192 B.n191 585
R132 B.n193 B.n66 585
R133 B.n195 B.n194 585
R134 B.n196 B.n65 585
R135 B.n198 B.n197 585
R136 B.n199 B.n64 585
R137 B.n201 B.n200 585
R138 B.n202 B.n63 585
R139 B.n204 B.n203 585
R140 B.n205 B.n62 585
R141 B.n129 B.n128 585
R142 B.n127 B.n92 585
R143 B.n126 B.n125 585
R144 B.n124 B.n93 585
R145 B.n123 B.n122 585
R146 B.n121 B.n94 585
R147 B.n120 B.n119 585
R148 B.n118 B.n95 585
R149 B.n117 B.n116 585
R150 B.n115 B.n96 585
R151 B.n114 B.n113 585
R152 B.n112 B.n97 585
R153 B.n111 B.n110 585
R154 B.n109 B.n98 585
R155 B.n108 B.n107 585
R156 B.n106 B.n99 585
R157 B.n105 B.n104 585
R158 B.n103 B.n100 585
R159 B.n102 B.n101 585
R160 B.n2 B.n0 585
R161 B.n373 B.n1 585
R162 B.n372 B.n371 585
R163 B.n370 B.n3 585
R164 B.n369 B.n368 585
R165 B.n367 B.n4 585
R166 B.n366 B.n365 585
R167 B.n364 B.n5 585
R168 B.n363 B.n362 585
R169 B.n361 B.n6 585
R170 B.n360 B.n359 585
R171 B.n358 B.n7 585
R172 B.n357 B.n356 585
R173 B.n355 B.n8 585
R174 B.n354 B.n353 585
R175 B.n352 B.n9 585
R176 B.n351 B.n350 585
R177 B.n349 B.n10 585
R178 B.n348 B.n347 585
R179 B.n346 B.n11 585
R180 B.n345 B.n344 585
R181 B.n375 B.n374 585
R182 B.n128 B.n91 521.33
R183 B.n344 B.n343 521.33
R184 B.n206 B.n205 521.33
R185 B.n266 B.n41 521.33
R186 B.n72 B.t3 368.298
R187 B.n80 B.t6 368.298
R188 B.n22 B.t0 368.298
R189 B.n30 B.t9 368.298
R190 B.n72 B.t5 266.647
R191 B.n30 B.t10 266.647
R192 B.n80 B.t8 266.647
R193 B.n22 B.t1 266.647
R194 B.n73 B.t4 246.865
R195 B.n31 B.t11 246.865
R196 B.n81 B.t7 246.865
R197 B.n23 B.t2 246.865
R198 B.n128 B.n127 163.367
R199 B.n127 B.n126 163.367
R200 B.n126 B.n93 163.367
R201 B.n122 B.n93 163.367
R202 B.n122 B.n121 163.367
R203 B.n121 B.n120 163.367
R204 B.n120 B.n95 163.367
R205 B.n116 B.n95 163.367
R206 B.n116 B.n115 163.367
R207 B.n115 B.n114 163.367
R208 B.n114 B.n97 163.367
R209 B.n110 B.n97 163.367
R210 B.n110 B.n109 163.367
R211 B.n109 B.n108 163.367
R212 B.n108 B.n99 163.367
R213 B.n104 B.n99 163.367
R214 B.n104 B.n103 163.367
R215 B.n103 B.n102 163.367
R216 B.n102 B.n2 163.367
R217 B.n374 B.n2 163.367
R218 B.n374 B.n373 163.367
R219 B.n373 B.n372 163.367
R220 B.n372 B.n3 163.367
R221 B.n368 B.n3 163.367
R222 B.n368 B.n367 163.367
R223 B.n367 B.n366 163.367
R224 B.n366 B.n5 163.367
R225 B.n362 B.n5 163.367
R226 B.n362 B.n361 163.367
R227 B.n361 B.n360 163.367
R228 B.n360 B.n7 163.367
R229 B.n356 B.n7 163.367
R230 B.n356 B.n355 163.367
R231 B.n355 B.n354 163.367
R232 B.n354 B.n9 163.367
R233 B.n350 B.n9 163.367
R234 B.n350 B.n349 163.367
R235 B.n349 B.n348 163.367
R236 B.n348 B.n11 163.367
R237 B.n344 B.n11 163.367
R238 B.n132 B.n91 163.367
R239 B.n133 B.n132 163.367
R240 B.n134 B.n133 163.367
R241 B.n134 B.n89 163.367
R242 B.n138 B.n89 163.367
R243 B.n139 B.n138 163.367
R244 B.n140 B.n139 163.367
R245 B.n140 B.n87 163.367
R246 B.n144 B.n87 163.367
R247 B.n145 B.n144 163.367
R248 B.n146 B.n145 163.367
R249 B.n146 B.n85 163.367
R250 B.n150 B.n85 163.367
R251 B.n151 B.n150 163.367
R252 B.n152 B.n151 163.367
R253 B.n152 B.n83 163.367
R254 B.n156 B.n83 163.367
R255 B.n157 B.n156 163.367
R256 B.n158 B.n157 163.367
R257 B.n158 B.n79 163.367
R258 B.n163 B.n79 163.367
R259 B.n164 B.n163 163.367
R260 B.n165 B.n164 163.367
R261 B.n165 B.n77 163.367
R262 B.n169 B.n77 163.367
R263 B.n170 B.n169 163.367
R264 B.n171 B.n170 163.367
R265 B.n171 B.n75 163.367
R266 B.n175 B.n75 163.367
R267 B.n176 B.n175 163.367
R268 B.n176 B.n71 163.367
R269 B.n180 B.n71 163.367
R270 B.n181 B.n180 163.367
R271 B.n182 B.n181 163.367
R272 B.n182 B.n69 163.367
R273 B.n186 B.n69 163.367
R274 B.n187 B.n186 163.367
R275 B.n188 B.n187 163.367
R276 B.n188 B.n67 163.367
R277 B.n192 B.n67 163.367
R278 B.n193 B.n192 163.367
R279 B.n194 B.n193 163.367
R280 B.n194 B.n65 163.367
R281 B.n198 B.n65 163.367
R282 B.n199 B.n198 163.367
R283 B.n200 B.n199 163.367
R284 B.n200 B.n63 163.367
R285 B.n204 B.n63 163.367
R286 B.n205 B.n204 163.367
R287 B.n206 B.n61 163.367
R288 B.n210 B.n61 163.367
R289 B.n211 B.n210 163.367
R290 B.n212 B.n211 163.367
R291 B.n212 B.n59 163.367
R292 B.n216 B.n59 163.367
R293 B.n217 B.n216 163.367
R294 B.n218 B.n217 163.367
R295 B.n218 B.n57 163.367
R296 B.n222 B.n57 163.367
R297 B.n223 B.n222 163.367
R298 B.n224 B.n223 163.367
R299 B.n224 B.n55 163.367
R300 B.n228 B.n55 163.367
R301 B.n229 B.n228 163.367
R302 B.n230 B.n229 163.367
R303 B.n230 B.n53 163.367
R304 B.n234 B.n53 163.367
R305 B.n235 B.n234 163.367
R306 B.n236 B.n235 163.367
R307 B.n236 B.n51 163.367
R308 B.n240 B.n51 163.367
R309 B.n241 B.n240 163.367
R310 B.n242 B.n241 163.367
R311 B.n242 B.n49 163.367
R312 B.n246 B.n49 163.367
R313 B.n247 B.n246 163.367
R314 B.n248 B.n247 163.367
R315 B.n248 B.n47 163.367
R316 B.n252 B.n47 163.367
R317 B.n253 B.n252 163.367
R318 B.n254 B.n253 163.367
R319 B.n254 B.n45 163.367
R320 B.n258 B.n45 163.367
R321 B.n259 B.n258 163.367
R322 B.n260 B.n259 163.367
R323 B.n260 B.n43 163.367
R324 B.n264 B.n43 163.367
R325 B.n265 B.n264 163.367
R326 B.n266 B.n265 163.367
R327 B.n343 B.n342 163.367
R328 B.n342 B.n13 163.367
R329 B.n338 B.n13 163.367
R330 B.n338 B.n337 163.367
R331 B.n337 B.n336 163.367
R332 B.n336 B.n15 163.367
R333 B.n332 B.n15 163.367
R334 B.n332 B.n331 163.367
R335 B.n331 B.n330 163.367
R336 B.n330 B.n17 163.367
R337 B.n326 B.n17 163.367
R338 B.n326 B.n325 163.367
R339 B.n325 B.n324 163.367
R340 B.n324 B.n19 163.367
R341 B.n320 B.n19 163.367
R342 B.n320 B.n319 163.367
R343 B.n319 B.n318 163.367
R344 B.n318 B.n21 163.367
R345 B.n314 B.n21 163.367
R346 B.n314 B.n313 163.367
R347 B.n313 B.n25 163.367
R348 B.n309 B.n25 163.367
R349 B.n309 B.n308 163.367
R350 B.n308 B.n307 163.367
R351 B.n307 B.n27 163.367
R352 B.n303 B.n27 163.367
R353 B.n303 B.n302 163.367
R354 B.n302 B.n301 163.367
R355 B.n301 B.n29 163.367
R356 B.n296 B.n29 163.367
R357 B.n296 B.n295 163.367
R358 B.n295 B.n294 163.367
R359 B.n294 B.n33 163.367
R360 B.n290 B.n33 163.367
R361 B.n290 B.n289 163.367
R362 B.n289 B.n288 163.367
R363 B.n288 B.n35 163.367
R364 B.n284 B.n35 163.367
R365 B.n284 B.n283 163.367
R366 B.n283 B.n282 163.367
R367 B.n282 B.n37 163.367
R368 B.n278 B.n37 163.367
R369 B.n278 B.n277 163.367
R370 B.n277 B.n276 163.367
R371 B.n276 B.n39 163.367
R372 B.n272 B.n39 163.367
R373 B.n272 B.n271 163.367
R374 B.n271 B.n270 163.367
R375 B.n270 B.n41 163.367
R376 B.n74 B.n73 59.5399
R377 B.n160 B.n81 59.5399
R378 B.n24 B.n23 59.5399
R379 B.n298 B.n31 59.5399
R380 B.n345 B.n12 33.8737
R381 B.n268 B.n267 33.8737
R382 B.n207 B.n62 33.8737
R383 B.n130 B.n129 33.8737
R384 B.n73 B.n72 19.7823
R385 B.n81 B.n80 19.7823
R386 B.n23 B.n22 19.7823
R387 B.n31 B.n30 19.7823
R388 B B.n375 18.0485
R389 B.n341 B.n12 10.6151
R390 B.n341 B.n340 10.6151
R391 B.n340 B.n339 10.6151
R392 B.n339 B.n14 10.6151
R393 B.n335 B.n14 10.6151
R394 B.n335 B.n334 10.6151
R395 B.n334 B.n333 10.6151
R396 B.n333 B.n16 10.6151
R397 B.n329 B.n16 10.6151
R398 B.n329 B.n328 10.6151
R399 B.n328 B.n327 10.6151
R400 B.n327 B.n18 10.6151
R401 B.n323 B.n18 10.6151
R402 B.n323 B.n322 10.6151
R403 B.n322 B.n321 10.6151
R404 B.n321 B.n20 10.6151
R405 B.n317 B.n20 10.6151
R406 B.n317 B.n316 10.6151
R407 B.n316 B.n315 10.6151
R408 B.n312 B.n311 10.6151
R409 B.n311 B.n310 10.6151
R410 B.n310 B.n26 10.6151
R411 B.n306 B.n26 10.6151
R412 B.n306 B.n305 10.6151
R413 B.n305 B.n304 10.6151
R414 B.n304 B.n28 10.6151
R415 B.n300 B.n28 10.6151
R416 B.n300 B.n299 10.6151
R417 B.n297 B.n32 10.6151
R418 B.n293 B.n32 10.6151
R419 B.n293 B.n292 10.6151
R420 B.n292 B.n291 10.6151
R421 B.n291 B.n34 10.6151
R422 B.n287 B.n34 10.6151
R423 B.n287 B.n286 10.6151
R424 B.n286 B.n285 10.6151
R425 B.n285 B.n36 10.6151
R426 B.n281 B.n36 10.6151
R427 B.n281 B.n280 10.6151
R428 B.n280 B.n279 10.6151
R429 B.n279 B.n38 10.6151
R430 B.n275 B.n38 10.6151
R431 B.n275 B.n274 10.6151
R432 B.n274 B.n273 10.6151
R433 B.n273 B.n40 10.6151
R434 B.n269 B.n40 10.6151
R435 B.n269 B.n268 10.6151
R436 B.n208 B.n207 10.6151
R437 B.n209 B.n208 10.6151
R438 B.n209 B.n60 10.6151
R439 B.n213 B.n60 10.6151
R440 B.n214 B.n213 10.6151
R441 B.n215 B.n214 10.6151
R442 B.n215 B.n58 10.6151
R443 B.n219 B.n58 10.6151
R444 B.n220 B.n219 10.6151
R445 B.n221 B.n220 10.6151
R446 B.n221 B.n56 10.6151
R447 B.n225 B.n56 10.6151
R448 B.n226 B.n225 10.6151
R449 B.n227 B.n226 10.6151
R450 B.n227 B.n54 10.6151
R451 B.n231 B.n54 10.6151
R452 B.n232 B.n231 10.6151
R453 B.n233 B.n232 10.6151
R454 B.n233 B.n52 10.6151
R455 B.n237 B.n52 10.6151
R456 B.n238 B.n237 10.6151
R457 B.n239 B.n238 10.6151
R458 B.n239 B.n50 10.6151
R459 B.n243 B.n50 10.6151
R460 B.n244 B.n243 10.6151
R461 B.n245 B.n244 10.6151
R462 B.n245 B.n48 10.6151
R463 B.n249 B.n48 10.6151
R464 B.n250 B.n249 10.6151
R465 B.n251 B.n250 10.6151
R466 B.n251 B.n46 10.6151
R467 B.n255 B.n46 10.6151
R468 B.n256 B.n255 10.6151
R469 B.n257 B.n256 10.6151
R470 B.n257 B.n44 10.6151
R471 B.n261 B.n44 10.6151
R472 B.n262 B.n261 10.6151
R473 B.n263 B.n262 10.6151
R474 B.n263 B.n42 10.6151
R475 B.n267 B.n42 10.6151
R476 B.n131 B.n130 10.6151
R477 B.n131 B.n90 10.6151
R478 B.n135 B.n90 10.6151
R479 B.n136 B.n135 10.6151
R480 B.n137 B.n136 10.6151
R481 B.n137 B.n88 10.6151
R482 B.n141 B.n88 10.6151
R483 B.n142 B.n141 10.6151
R484 B.n143 B.n142 10.6151
R485 B.n143 B.n86 10.6151
R486 B.n147 B.n86 10.6151
R487 B.n148 B.n147 10.6151
R488 B.n149 B.n148 10.6151
R489 B.n149 B.n84 10.6151
R490 B.n153 B.n84 10.6151
R491 B.n154 B.n153 10.6151
R492 B.n155 B.n154 10.6151
R493 B.n155 B.n82 10.6151
R494 B.n159 B.n82 10.6151
R495 B.n162 B.n161 10.6151
R496 B.n162 B.n78 10.6151
R497 B.n166 B.n78 10.6151
R498 B.n167 B.n166 10.6151
R499 B.n168 B.n167 10.6151
R500 B.n168 B.n76 10.6151
R501 B.n172 B.n76 10.6151
R502 B.n173 B.n172 10.6151
R503 B.n174 B.n173 10.6151
R504 B.n178 B.n177 10.6151
R505 B.n179 B.n178 10.6151
R506 B.n179 B.n70 10.6151
R507 B.n183 B.n70 10.6151
R508 B.n184 B.n183 10.6151
R509 B.n185 B.n184 10.6151
R510 B.n185 B.n68 10.6151
R511 B.n189 B.n68 10.6151
R512 B.n190 B.n189 10.6151
R513 B.n191 B.n190 10.6151
R514 B.n191 B.n66 10.6151
R515 B.n195 B.n66 10.6151
R516 B.n196 B.n195 10.6151
R517 B.n197 B.n196 10.6151
R518 B.n197 B.n64 10.6151
R519 B.n201 B.n64 10.6151
R520 B.n202 B.n201 10.6151
R521 B.n203 B.n202 10.6151
R522 B.n203 B.n62 10.6151
R523 B.n129 B.n92 10.6151
R524 B.n125 B.n92 10.6151
R525 B.n125 B.n124 10.6151
R526 B.n124 B.n123 10.6151
R527 B.n123 B.n94 10.6151
R528 B.n119 B.n94 10.6151
R529 B.n119 B.n118 10.6151
R530 B.n118 B.n117 10.6151
R531 B.n117 B.n96 10.6151
R532 B.n113 B.n96 10.6151
R533 B.n113 B.n112 10.6151
R534 B.n112 B.n111 10.6151
R535 B.n111 B.n98 10.6151
R536 B.n107 B.n98 10.6151
R537 B.n107 B.n106 10.6151
R538 B.n106 B.n105 10.6151
R539 B.n105 B.n100 10.6151
R540 B.n101 B.n100 10.6151
R541 B.n101 B.n0 10.6151
R542 B.n371 B.n1 10.6151
R543 B.n371 B.n370 10.6151
R544 B.n370 B.n369 10.6151
R545 B.n369 B.n4 10.6151
R546 B.n365 B.n4 10.6151
R547 B.n365 B.n364 10.6151
R548 B.n364 B.n363 10.6151
R549 B.n363 B.n6 10.6151
R550 B.n359 B.n6 10.6151
R551 B.n359 B.n358 10.6151
R552 B.n358 B.n357 10.6151
R553 B.n357 B.n8 10.6151
R554 B.n353 B.n8 10.6151
R555 B.n353 B.n352 10.6151
R556 B.n352 B.n351 10.6151
R557 B.n351 B.n10 10.6151
R558 B.n347 B.n10 10.6151
R559 B.n347 B.n346 10.6151
R560 B.n346 B.n345 10.6151
R561 B.n315 B.n24 9.36635
R562 B.n298 B.n297 9.36635
R563 B.n160 B.n159 9.36635
R564 B.n177 B.n74 9.36635
R565 B.n375 B.n0 2.81026
R566 B.n375 B.n1 2.81026
R567 B.n312 B.n24 1.24928
R568 B.n299 B.n298 1.24928
R569 B.n161 B.n160 1.24928
R570 B.n174 B.n74 1.24928
R571 VP.n3 VP.t2 243.886
R572 VP.n8 VP.t1 222.488
R573 VP.n12 VP.t3 222.488
R574 VP.n14 VP.t0 222.488
R575 VP.n6 VP.t5 222.488
R576 VP.n4 VP.t4 222.488
R577 VP.n15 VP.n14 161.3
R578 VP.n5 VP.n2 161.3
R579 VP.n7 VP.n6 161.3
R580 VP.n13 VP.n0 161.3
R581 VP.n12 VP.n11 161.3
R582 VP.n10 VP.n1 161.3
R583 VP.n9 VP.n8 161.3
R584 VP.n3 VP.n2 44.853
R585 VP.n9 VP.n7 35.6444
R586 VP.n8 VP.n1 25.5611
R587 VP.n14 VP.n13 25.5611
R588 VP.n6 VP.n5 25.5611
R589 VP.n12 VP.n1 22.6399
R590 VP.n13 VP.n12 22.6399
R591 VP.n5 VP.n4 22.6399
R592 VP.n4 VP.n3 20.5405
R593 VP.n7 VP.n2 0.189894
R594 VP.n10 VP.n9 0.189894
R595 VP.n11 VP.n10 0.189894
R596 VP.n11 VP.n0 0.189894
R597 VP.n15 VP.n0 0.189894
R598 VP VP.n15 0.0516364
R599 VTAIL.n98 VTAIL.n80 756.745
R600 VTAIL.n20 VTAIL.n2 756.745
R601 VTAIL.n74 VTAIL.n56 756.745
R602 VTAIL.n48 VTAIL.n30 756.745
R603 VTAIL.n89 VTAIL.n88 585
R604 VTAIL.n91 VTAIL.n90 585
R605 VTAIL.n84 VTAIL.n83 585
R606 VTAIL.n97 VTAIL.n96 585
R607 VTAIL.n99 VTAIL.n98 585
R608 VTAIL.n11 VTAIL.n10 585
R609 VTAIL.n13 VTAIL.n12 585
R610 VTAIL.n6 VTAIL.n5 585
R611 VTAIL.n19 VTAIL.n18 585
R612 VTAIL.n21 VTAIL.n20 585
R613 VTAIL.n75 VTAIL.n74 585
R614 VTAIL.n73 VTAIL.n72 585
R615 VTAIL.n60 VTAIL.n59 585
R616 VTAIL.n67 VTAIL.n66 585
R617 VTAIL.n65 VTAIL.n64 585
R618 VTAIL.n49 VTAIL.n48 585
R619 VTAIL.n47 VTAIL.n46 585
R620 VTAIL.n34 VTAIL.n33 585
R621 VTAIL.n41 VTAIL.n40 585
R622 VTAIL.n39 VTAIL.n38 585
R623 VTAIL.n87 VTAIL.t4 328.587
R624 VTAIL.n9 VTAIL.t7 328.587
R625 VTAIL.n63 VTAIL.t8 328.587
R626 VTAIL.n37 VTAIL.t0 328.587
R627 VTAIL.n90 VTAIL.n89 171.744
R628 VTAIL.n90 VTAIL.n83 171.744
R629 VTAIL.n97 VTAIL.n83 171.744
R630 VTAIL.n98 VTAIL.n97 171.744
R631 VTAIL.n12 VTAIL.n11 171.744
R632 VTAIL.n12 VTAIL.n5 171.744
R633 VTAIL.n19 VTAIL.n5 171.744
R634 VTAIL.n20 VTAIL.n19 171.744
R635 VTAIL.n74 VTAIL.n73 171.744
R636 VTAIL.n73 VTAIL.n59 171.744
R637 VTAIL.n66 VTAIL.n59 171.744
R638 VTAIL.n66 VTAIL.n65 171.744
R639 VTAIL.n48 VTAIL.n47 171.744
R640 VTAIL.n47 VTAIL.n33 171.744
R641 VTAIL.n40 VTAIL.n33 171.744
R642 VTAIL.n40 VTAIL.n39 171.744
R643 VTAIL.n55 VTAIL.n54 90.698
R644 VTAIL.n29 VTAIL.n28 90.698
R645 VTAIL.n1 VTAIL.n0 90.6978
R646 VTAIL.n27 VTAIL.n26 90.6978
R647 VTAIL.n89 VTAIL.t4 85.8723
R648 VTAIL.n11 VTAIL.t7 85.8723
R649 VTAIL.n65 VTAIL.t8 85.8723
R650 VTAIL.n39 VTAIL.t0 85.8723
R651 VTAIL.n103 VTAIL.n102 35.4823
R652 VTAIL.n25 VTAIL.n24 35.4823
R653 VTAIL.n79 VTAIL.n78 35.4823
R654 VTAIL.n53 VTAIL.n52 35.4823
R655 VTAIL.n29 VTAIL.n27 18.2031
R656 VTAIL.n103 VTAIL.n79 17.3238
R657 VTAIL.n88 VTAIL.n87 16.3651
R658 VTAIL.n10 VTAIL.n9 16.3651
R659 VTAIL.n64 VTAIL.n63 16.3651
R660 VTAIL.n38 VTAIL.n37 16.3651
R661 VTAIL.n91 VTAIL.n86 12.8005
R662 VTAIL.n13 VTAIL.n8 12.8005
R663 VTAIL.n67 VTAIL.n62 12.8005
R664 VTAIL.n41 VTAIL.n36 12.8005
R665 VTAIL.n92 VTAIL.n84 12.0247
R666 VTAIL.n14 VTAIL.n6 12.0247
R667 VTAIL.n68 VTAIL.n60 12.0247
R668 VTAIL.n42 VTAIL.n34 12.0247
R669 VTAIL.n96 VTAIL.n95 11.249
R670 VTAIL.n18 VTAIL.n17 11.249
R671 VTAIL.n72 VTAIL.n71 11.249
R672 VTAIL.n46 VTAIL.n45 11.249
R673 VTAIL.n99 VTAIL.n82 10.4732
R674 VTAIL.n21 VTAIL.n4 10.4732
R675 VTAIL.n75 VTAIL.n58 10.4732
R676 VTAIL.n49 VTAIL.n32 10.4732
R677 VTAIL.n100 VTAIL.n80 9.69747
R678 VTAIL.n22 VTAIL.n2 9.69747
R679 VTAIL.n76 VTAIL.n56 9.69747
R680 VTAIL.n50 VTAIL.n30 9.69747
R681 VTAIL.n102 VTAIL.n101 9.45567
R682 VTAIL.n24 VTAIL.n23 9.45567
R683 VTAIL.n78 VTAIL.n77 9.45567
R684 VTAIL.n52 VTAIL.n51 9.45567
R685 VTAIL.n101 VTAIL.n100 9.3005
R686 VTAIL.n82 VTAIL.n81 9.3005
R687 VTAIL.n95 VTAIL.n94 9.3005
R688 VTAIL.n93 VTAIL.n92 9.3005
R689 VTAIL.n86 VTAIL.n85 9.3005
R690 VTAIL.n23 VTAIL.n22 9.3005
R691 VTAIL.n4 VTAIL.n3 9.3005
R692 VTAIL.n17 VTAIL.n16 9.3005
R693 VTAIL.n15 VTAIL.n14 9.3005
R694 VTAIL.n8 VTAIL.n7 9.3005
R695 VTAIL.n77 VTAIL.n76 9.3005
R696 VTAIL.n58 VTAIL.n57 9.3005
R697 VTAIL.n71 VTAIL.n70 9.3005
R698 VTAIL.n69 VTAIL.n68 9.3005
R699 VTAIL.n62 VTAIL.n61 9.3005
R700 VTAIL.n51 VTAIL.n50 9.3005
R701 VTAIL.n32 VTAIL.n31 9.3005
R702 VTAIL.n45 VTAIL.n44 9.3005
R703 VTAIL.n43 VTAIL.n42 9.3005
R704 VTAIL.n36 VTAIL.n35 9.3005
R705 VTAIL.n0 VTAIL.t5 6.87259
R706 VTAIL.n0 VTAIL.t3 6.87259
R707 VTAIL.n26 VTAIL.t11 6.87259
R708 VTAIL.n26 VTAIL.t10 6.87259
R709 VTAIL.n54 VTAIL.t6 6.87259
R710 VTAIL.n54 VTAIL.t9 6.87259
R711 VTAIL.n28 VTAIL.t2 6.87259
R712 VTAIL.n28 VTAIL.t1 6.87259
R713 VTAIL.n102 VTAIL.n80 4.26717
R714 VTAIL.n24 VTAIL.n2 4.26717
R715 VTAIL.n78 VTAIL.n56 4.26717
R716 VTAIL.n52 VTAIL.n30 4.26717
R717 VTAIL.n87 VTAIL.n85 3.73474
R718 VTAIL.n9 VTAIL.n7 3.73474
R719 VTAIL.n63 VTAIL.n61 3.73474
R720 VTAIL.n37 VTAIL.n35 3.73474
R721 VTAIL.n100 VTAIL.n99 3.49141
R722 VTAIL.n22 VTAIL.n21 3.49141
R723 VTAIL.n76 VTAIL.n75 3.49141
R724 VTAIL.n50 VTAIL.n49 3.49141
R725 VTAIL.n96 VTAIL.n82 2.71565
R726 VTAIL.n18 VTAIL.n4 2.71565
R727 VTAIL.n72 VTAIL.n58 2.71565
R728 VTAIL.n46 VTAIL.n32 2.71565
R729 VTAIL.n95 VTAIL.n84 1.93989
R730 VTAIL.n17 VTAIL.n6 1.93989
R731 VTAIL.n71 VTAIL.n60 1.93989
R732 VTAIL.n45 VTAIL.n34 1.93989
R733 VTAIL.n92 VTAIL.n91 1.16414
R734 VTAIL.n14 VTAIL.n13 1.16414
R735 VTAIL.n68 VTAIL.n67 1.16414
R736 VTAIL.n42 VTAIL.n41 1.16414
R737 VTAIL.n55 VTAIL.n53 0.909983
R738 VTAIL.n25 VTAIL.n1 0.909983
R739 VTAIL.n53 VTAIL.n29 0.87981
R740 VTAIL.n79 VTAIL.n55 0.87981
R741 VTAIL.n27 VTAIL.n25 0.87981
R742 VTAIL VTAIL.n103 0.601793
R743 VTAIL.n88 VTAIL.n86 0.388379
R744 VTAIL.n10 VTAIL.n8 0.388379
R745 VTAIL.n64 VTAIL.n62 0.388379
R746 VTAIL.n38 VTAIL.n36 0.388379
R747 VTAIL VTAIL.n1 0.278517
R748 VTAIL.n93 VTAIL.n85 0.155672
R749 VTAIL.n94 VTAIL.n93 0.155672
R750 VTAIL.n94 VTAIL.n81 0.155672
R751 VTAIL.n101 VTAIL.n81 0.155672
R752 VTAIL.n15 VTAIL.n7 0.155672
R753 VTAIL.n16 VTAIL.n15 0.155672
R754 VTAIL.n16 VTAIL.n3 0.155672
R755 VTAIL.n23 VTAIL.n3 0.155672
R756 VTAIL.n77 VTAIL.n57 0.155672
R757 VTAIL.n70 VTAIL.n57 0.155672
R758 VTAIL.n70 VTAIL.n69 0.155672
R759 VTAIL.n69 VTAIL.n61 0.155672
R760 VTAIL.n51 VTAIL.n31 0.155672
R761 VTAIL.n44 VTAIL.n31 0.155672
R762 VTAIL.n44 VTAIL.n43 0.155672
R763 VTAIL.n43 VTAIL.n35 0.155672
R764 VDD1.n18 VDD1.n0 756.745
R765 VDD1.n41 VDD1.n23 756.745
R766 VDD1.n19 VDD1.n18 585
R767 VDD1.n17 VDD1.n16 585
R768 VDD1.n4 VDD1.n3 585
R769 VDD1.n11 VDD1.n10 585
R770 VDD1.n9 VDD1.n8 585
R771 VDD1.n32 VDD1.n31 585
R772 VDD1.n34 VDD1.n33 585
R773 VDD1.n27 VDD1.n26 585
R774 VDD1.n40 VDD1.n39 585
R775 VDD1.n42 VDD1.n41 585
R776 VDD1.n7 VDD1.t3 328.587
R777 VDD1.n30 VDD1.t4 328.587
R778 VDD1.n18 VDD1.n17 171.744
R779 VDD1.n17 VDD1.n3 171.744
R780 VDD1.n10 VDD1.n3 171.744
R781 VDD1.n10 VDD1.n9 171.744
R782 VDD1.n33 VDD1.n32 171.744
R783 VDD1.n33 VDD1.n26 171.744
R784 VDD1.n40 VDD1.n26 171.744
R785 VDD1.n41 VDD1.n40 171.744
R786 VDD1.n47 VDD1.n46 107.541
R787 VDD1.n49 VDD1.n48 107.376
R788 VDD1.n9 VDD1.t3 85.8723
R789 VDD1.n32 VDD1.t4 85.8723
R790 VDD1 VDD1.n22 52.8788
R791 VDD1.n47 VDD1.n45 52.7652
R792 VDD1.n49 VDD1.n47 31.6733
R793 VDD1.n8 VDD1.n7 16.3651
R794 VDD1.n31 VDD1.n30 16.3651
R795 VDD1.n11 VDD1.n6 12.8005
R796 VDD1.n34 VDD1.n29 12.8005
R797 VDD1.n12 VDD1.n4 12.0247
R798 VDD1.n35 VDD1.n27 12.0247
R799 VDD1.n16 VDD1.n15 11.249
R800 VDD1.n39 VDD1.n38 11.249
R801 VDD1.n19 VDD1.n2 10.4732
R802 VDD1.n42 VDD1.n25 10.4732
R803 VDD1.n20 VDD1.n0 9.69747
R804 VDD1.n43 VDD1.n23 9.69747
R805 VDD1.n22 VDD1.n21 9.45567
R806 VDD1.n45 VDD1.n44 9.45567
R807 VDD1.n21 VDD1.n20 9.3005
R808 VDD1.n2 VDD1.n1 9.3005
R809 VDD1.n15 VDD1.n14 9.3005
R810 VDD1.n13 VDD1.n12 9.3005
R811 VDD1.n6 VDD1.n5 9.3005
R812 VDD1.n44 VDD1.n43 9.3005
R813 VDD1.n25 VDD1.n24 9.3005
R814 VDD1.n38 VDD1.n37 9.3005
R815 VDD1.n36 VDD1.n35 9.3005
R816 VDD1.n29 VDD1.n28 9.3005
R817 VDD1.n48 VDD1.t1 6.87259
R818 VDD1.n48 VDD1.t0 6.87259
R819 VDD1.n46 VDD1.t2 6.87259
R820 VDD1.n46 VDD1.t5 6.87259
R821 VDD1.n22 VDD1.n0 4.26717
R822 VDD1.n45 VDD1.n23 4.26717
R823 VDD1.n7 VDD1.n5 3.73474
R824 VDD1.n30 VDD1.n28 3.73474
R825 VDD1.n20 VDD1.n19 3.49141
R826 VDD1.n43 VDD1.n42 3.49141
R827 VDD1.n16 VDD1.n2 2.71565
R828 VDD1.n39 VDD1.n25 2.71565
R829 VDD1.n15 VDD1.n4 1.93989
R830 VDD1.n38 VDD1.n27 1.93989
R831 VDD1.n12 VDD1.n11 1.16414
R832 VDD1.n35 VDD1.n34 1.16414
R833 VDD1.n8 VDD1.n6 0.388379
R834 VDD1.n31 VDD1.n29 0.388379
R835 VDD1 VDD1.n49 0.162138
R836 VDD1.n21 VDD1.n1 0.155672
R837 VDD1.n14 VDD1.n1 0.155672
R838 VDD1.n14 VDD1.n13 0.155672
R839 VDD1.n13 VDD1.n5 0.155672
R840 VDD1.n36 VDD1.n28 0.155672
R841 VDD1.n37 VDD1.n36 0.155672
R842 VDD1.n37 VDD1.n24 0.155672
R843 VDD1.n44 VDD1.n24 0.155672
R844 VN.n1 VN.t1 243.886
R845 VN.n7 VN.t2 243.886
R846 VN.n2 VN.t4 222.488
R847 VN.n4 VN.t0 222.488
R848 VN.n8 VN.t3 222.488
R849 VN.n10 VN.t5 222.488
R850 VN.n5 VN.n4 161.3
R851 VN.n11 VN.n10 161.3
R852 VN.n9 VN.n6 161.3
R853 VN.n3 VN.n0 161.3
R854 VN.n7 VN.n6 44.853
R855 VN.n1 VN.n0 44.853
R856 VN VN.n11 36.0251
R857 VN.n4 VN.n3 25.5611
R858 VN.n10 VN.n9 25.5611
R859 VN.n3 VN.n2 22.6399
R860 VN.n9 VN.n8 22.6399
R861 VN.n2 VN.n1 20.5405
R862 VN.n8 VN.n7 20.5405
R863 VN.n11 VN.n6 0.189894
R864 VN.n5 VN.n0 0.189894
R865 VN VN.n5 0.0516364
R866 VDD2.n43 VDD2.n25 756.745
R867 VDD2.n18 VDD2.n0 756.745
R868 VDD2.n44 VDD2.n43 585
R869 VDD2.n42 VDD2.n41 585
R870 VDD2.n29 VDD2.n28 585
R871 VDD2.n36 VDD2.n35 585
R872 VDD2.n34 VDD2.n33 585
R873 VDD2.n9 VDD2.n8 585
R874 VDD2.n11 VDD2.n10 585
R875 VDD2.n4 VDD2.n3 585
R876 VDD2.n17 VDD2.n16 585
R877 VDD2.n19 VDD2.n18 585
R878 VDD2.n32 VDD2.t0 328.587
R879 VDD2.n7 VDD2.t4 328.587
R880 VDD2.n43 VDD2.n42 171.744
R881 VDD2.n42 VDD2.n28 171.744
R882 VDD2.n35 VDD2.n28 171.744
R883 VDD2.n35 VDD2.n34 171.744
R884 VDD2.n10 VDD2.n9 171.744
R885 VDD2.n10 VDD2.n3 171.744
R886 VDD2.n17 VDD2.n3 171.744
R887 VDD2.n18 VDD2.n17 171.744
R888 VDD2.n24 VDD2.n23 107.541
R889 VDD2 VDD2.n49 107.538
R890 VDD2.n34 VDD2.t0 85.8723
R891 VDD2.n9 VDD2.t4 85.8723
R892 VDD2.n24 VDD2.n22 52.7652
R893 VDD2.n48 VDD2.n47 52.1611
R894 VDD2.n48 VDD2.n24 30.6506
R895 VDD2.n33 VDD2.n32 16.3651
R896 VDD2.n8 VDD2.n7 16.3651
R897 VDD2.n36 VDD2.n31 12.8005
R898 VDD2.n11 VDD2.n6 12.8005
R899 VDD2.n37 VDD2.n29 12.0247
R900 VDD2.n12 VDD2.n4 12.0247
R901 VDD2.n41 VDD2.n40 11.249
R902 VDD2.n16 VDD2.n15 11.249
R903 VDD2.n44 VDD2.n27 10.4732
R904 VDD2.n19 VDD2.n2 10.4732
R905 VDD2.n45 VDD2.n25 9.69747
R906 VDD2.n20 VDD2.n0 9.69747
R907 VDD2.n47 VDD2.n46 9.45567
R908 VDD2.n22 VDD2.n21 9.45567
R909 VDD2.n46 VDD2.n45 9.3005
R910 VDD2.n27 VDD2.n26 9.3005
R911 VDD2.n40 VDD2.n39 9.3005
R912 VDD2.n38 VDD2.n37 9.3005
R913 VDD2.n31 VDD2.n30 9.3005
R914 VDD2.n21 VDD2.n20 9.3005
R915 VDD2.n2 VDD2.n1 9.3005
R916 VDD2.n15 VDD2.n14 9.3005
R917 VDD2.n13 VDD2.n12 9.3005
R918 VDD2.n6 VDD2.n5 9.3005
R919 VDD2.n49 VDD2.t2 6.87259
R920 VDD2.n49 VDD2.t3 6.87259
R921 VDD2.n23 VDD2.t1 6.87259
R922 VDD2.n23 VDD2.t5 6.87259
R923 VDD2.n47 VDD2.n25 4.26717
R924 VDD2.n22 VDD2.n0 4.26717
R925 VDD2.n32 VDD2.n30 3.73474
R926 VDD2.n7 VDD2.n5 3.73474
R927 VDD2.n45 VDD2.n44 3.49141
R928 VDD2.n20 VDD2.n19 3.49141
R929 VDD2.n41 VDD2.n27 2.71565
R930 VDD2.n16 VDD2.n2 2.71565
R931 VDD2.n40 VDD2.n29 1.93989
R932 VDD2.n15 VDD2.n4 1.93989
R933 VDD2.n37 VDD2.n36 1.16414
R934 VDD2.n12 VDD2.n11 1.16414
R935 VDD2 VDD2.n48 0.718172
R936 VDD2.n33 VDD2.n31 0.388379
R937 VDD2.n8 VDD2.n6 0.388379
R938 VDD2.n46 VDD2.n26 0.155672
R939 VDD2.n39 VDD2.n26 0.155672
R940 VDD2.n39 VDD2.n38 0.155672
R941 VDD2.n38 VDD2.n30 0.155672
R942 VDD2.n13 VDD2.n5 0.155672
R943 VDD2.n14 VDD2.n13 0.155672
R944 VDD2.n14 VDD2.n1 0.155672
R945 VDD2.n21 VDD2.n1 0.155672
C0 VP VN 3.72649f
C1 B VDD2 1.0565f
C2 VP B 1.0458f
C3 VP VDD2 0.29965f
C4 w_n1786_n1914# VN 2.79025f
C5 w_n1786_n1914# B 5.00108f
C6 VDD1 VN 0.151794f
C7 w_n1786_n1914# VDD2 1.29041f
C8 B VDD1 1.02772f
C9 VP w_n1786_n1914# 3.01574f
C10 VDD1 VDD2 0.703623f
C11 VP VDD1 2.05128f
C12 w_n1786_n1914# VDD1 1.26694f
C13 VTAIL VN 1.94357f
C14 B VTAIL 1.39832f
C15 VDD2 VTAIL 5.10521f
C16 VP VTAIL 1.95787f
C17 w_n1786_n1914# VTAIL 1.76942f
C18 VDD1 VTAIL 5.06717f
C19 B VN 0.678871f
C20 VDD2 VN 1.90575f
C21 VDD2 VSUBS 0.845228f
C22 VDD1 VSUBS 0.898919f
C23 VTAIL VSUBS 0.375744f
C24 VN VSUBS 3.08873f
C25 VP VSUBS 1.103979f
C26 B VSUBS 2.038693f
C27 w_n1786_n1914# VSUBS 42.8854f
C28 VDD2.n0 VSUBS 0.019363f
C29 VDD2.n1 VSUBS 0.017094f
C30 VDD2.n2 VSUBS 0.009185f
C31 VDD2.n3 VSUBS 0.021711f
C32 VDD2.n4 VSUBS 0.009726f
C33 VDD2.n5 VSUBS 0.291647f
C34 VDD2.n6 VSUBS 0.009185f
C35 VDD2.t4 VSUBS 0.047603f
C36 VDD2.n7 VSUBS 0.070076f
C37 VDD2.n8 VSUBS 0.013754f
C38 VDD2.n9 VSUBS 0.016283f
C39 VDD2.n10 VSUBS 0.021711f
C40 VDD2.n11 VSUBS 0.009726f
C41 VDD2.n12 VSUBS 0.009185f
C42 VDD2.n13 VSUBS 0.017094f
C43 VDD2.n14 VSUBS 0.017094f
C44 VDD2.n15 VSUBS 0.009185f
C45 VDD2.n16 VSUBS 0.009726f
C46 VDD2.n17 VSUBS 0.021711f
C47 VDD2.n18 VSUBS 0.054538f
C48 VDD2.n19 VSUBS 0.009726f
C49 VDD2.n20 VSUBS 0.009185f
C50 VDD2.n21 VSUBS 0.043481f
C51 VDD2.n22 VSUBS 0.040198f
C52 VDD2.t1 VSUBS 0.063893f
C53 VDD2.t5 VSUBS 0.063893f
C54 VDD2.n23 VSUBS 0.395996f
C55 VDD2.n24 VSUBS 1.08792f
C56 VDD2.n25 VSUBS 0.019363f
C57 VDD2.n26 VSUBS 0.017094f
C58 VDD2.n27 VSUBS 0.009185f
C59 VDD2.n28 VSUBS 0.021711f
C60 VDD2.n29 VSUBS 0.009726f
C61 VDD2.n30 VSUBS 0.291647f
C62 VDD2.n31 VSUBS 0.009185f
C63 VDD2.t0 VSUBS 0.047603f
C64 VDD2.n32 VSUBS 0.070076f
C65 VDD2.n33 VSUBS 0.013754f
C66 VDD2.n34 VSUBS 0.016283f
C67 VDD2.n35 VSUBS 0.021711f
C68 VDD2.n36 VSUBS 0.009726f
C69 VDD2.n37 VSUBS 0.009185f
C70 VDD2.n38 VSUBS 0.017094f
C71 VDD2.n39 VSUBS 0.017094f
C72 VDD2.n40 VSUBS 0.009185f
C73 VDD2.n41 VSUBS 0.009726f
C74 VDD2.n42 VSUBS 0.021711f
C75 VDD2.n43 VSUBS 0.054538f
C76 VDD2.n44 VSUBS 0.009726f
C77 VDD2.n45 VSUBS 0.009185f
C78 VDD2.n46 VSUBS 0.043481f
C79 VDD2.n47 VSUBS 0.039406f
C80 VDD2.n48 VSUBS 1.00083f
C81 VDD2.t2 VSUBS 0.063893f
C82 VDD2.t3 VSUBS 0.063893f
C83 VDD2.n49 VSUBS 0.395984f
C84 VN.n0 VSUBS 0.1687f
C85 VN.t1 VSUBS 0.408228f
C86 VN.n1 VSUBS 0.180759f
C87 VN.t4 VSUBS 0.391234f
C88 VN.n2 VSUBS 0.197432f
C89 VN.n3 VSUBS 0.009288f
C90 VN.t0 VSUBS 0.391234f
C91 VN.n4 VSUBS 0.190836f
C92 VN.n5 VSUBS 0.031718f
C93 VN.n6 VSUBS 0.1687f
C94 VN.t2 VSUBS 0.408228f
C95 VN.n7 VSUBS 0.180759f
C96 VN.t3 VSUBS 0.391234f
C97 VN.n8 VSUBS 0.197432f
C98 VN.n9 VSUBS 0.009288f
C99 VN.t5 VSUBS 0.391234f
C100 VN.n10 VSUBS 0.190836f
C101 VN.n11 VSUBS 1.29005f
C102 VDD1.n0 VSUBS 0.027002f
C103 VDD1.n1 VSUBS 0.023837f
C104 VDD1.n2 VSUBS 0.012809f
C105 VDD1.n3 VSUBS 0.030276f
C106 VDD1.n4 VSUBS 0.013563f
C107 VDD1.n5 VSUBS 0.406702f
C108 VDD1.n6 VSUBS 0.012809f
C109 VDD1.t3 VSUBS 0.066382f
C110 VDD1.n7 VSUBS 0.097721f
C111 VDD1.n8 VSUBS 0.01918f
C112 VDD1.n9 VSUBS 0.022707f
C113 VDD1.n10 VSUBS 0.030276f
C114 VDD1.n11 VSUBS 0.013563f
C115 VDD1.n12 VSUBS 0.012809f
C116 VDD1.n13 VSUBS 0.023837f
C117 VDD1.n14 VSUBS 0.023837f
C118 VDD1.n15 VSUBS 0.012809f
C119 VDD1.n16 VSUBS 0.013563f
C120 VDD1.n17 VSUBS 0.030276f
C121 VDD1.n18 VSUBS 0.076054f
C122 VDD1.n19 VSUBS 0.013563f
C123 VDD1.n20 VSUBS 0.012809f
C124 VDD1.n21 VSUBS 0.060635f
C125 VDD1.n22 VSUBS 0.056366f
C126 VDD1.n23 VSUBS 0.027002f
C127 VDD1.n24 VSUBS 0.023837f
C128 VDD1.n25 VSUBS 0.012809f
C129 VDD1.n26 VSUBS 0.030276f
C130 VDD1.n27 VSUBS 0.013563f
C131 VDD1.n28 VSUBS 0.406702f
C132 VDD1.n29 VSUBS 0.012809f
C133 VDD1.t4 VSUBS 0.066382f
C134 VDD1.n30 VSUBS 0.097721f
C135 VDD1.n31 VSUBS 0.01918f
C136 VDD1.n32 VSUBS 0.022707f
C137 VDD1.n33 VSUBS 0.030276f
C138 VDD1.n34 VSUBS 0.013563f
C139 VDD1.n35 VSUBS 0.012809f
C140 VDD1.n36 VSUBS 0.023837f
C141 VDD1.n37 VSUBS 0.023837f
C142 VDD1.n38 VSUBS 0.012809f
C143 VDD1.n39 VSUBS 0.013563f
C144 VDD1.n40 VSUBS 0.030276f
C145 VDD1.n41 VSUBS 0.076054f
C146 VDD1.n42 VSUBS 0.013563f
C147 VDD1.n43 VSUBS 0.012809f
C148 VDD1.n44 VSUBS 0.060635f
C149 VDD1.n45 VSUBS 0.056056f
C150 VDD1.t2 VSUBS 0.089099f
C151 VDD1.t5 VSUBS 0.089099f
C152 VDD1.n46 VSUBS 0.552218f
C153 VDD1.n47 VSUBS 1.58733f
C154 VDD1.t1 VSUBS 0.089099f
C155 VDD1.t0 VSUBS 0.089099f
C156 VDD1.n48 VSUBS 0.551529f
C157 VDD1.n49 VSUBS 1.75574f
C158 VTAIL.t5 VSUBS 0.072902f
C159 VTAIL.t3 VSUBS 0.072902f
C160 VTAIL.n0 VSUBS 0.39825f
C161 VTAIL.n1 VSUBS 0.393176f
C162 VTAIL.n2 VSUBS 0.022093f
C163 VTAIL.n3 VSUBS 0.019504f
C164 VTAIL.n4 VSUBS 0.010481f
C165 VTAIL.n5 VSUBS 0.024772f
C166 VTAIL.n6 VSUBS 0.011097f
C167 VTAIL.n7 VSUBS 0.332771f
C168 VTAIL.n8 VSUBS 0.010481f
C169 VTAIL.t7 VSUBS 0.054315f
C170 VTAIL.n9 VSUBS 0.079957f
C171 VTAIL.n10 VSUBS 0.015694f
C172 VTAIL.n11 VSUBS 0.018579f
C173 VTAIL.n12 VSUBS 0.024772f
C174 VTAIL.n13 VSUBS 0.011097f
C175 VTAIL.n14 VSUBS 0.010481f
C176 VTAIL.n15 VSUBS 0.019504f
C177 VTAIL.n16 VSUBS 0.019504f
C178 VTAIL.n17 VSUBS 0.010481f
C179 VTAIL.n18 VSUBS 0.011097f
C180 VTAIL.n19 VSUBS 0.024772f
C181 VTAIL.n20 VSUBS 0.062228f
C182 VTAIL.n21 VSUBS 0.011097f
C183 VTAIL.n22 VSUBS 0.010481f
C184 VTAIL.n23 VSUBS 0.049612f
C185 VTAIL.n24 VSUBS 0.031528f
C186 VTAIL.n25 VSUBS 0.13164f
C187 VTAIL.t11 VSUBS 0.072902f
C188 VTAIL.t10 VSUBS 0.072902f
C189 VTAIL.n26 VSUBS 0.39825f
C190 VTAIL.n27 VSUBS 1.00553f
C191 VTAIL.t2 VSUBS 0.072902f
C192 VTAIL.t1 VSUBS 0.072902f
C193 VTAIL.n28 VSUBS 0.398253f
C194 VTAIL.n29 VSUBS 1.00553f
C195 VTAIL.n30 VSUBS 0.022093f
C196 VTAIL.n31 VSUBS 0.019504f
C197 VTAIL.n32 VSUBS 0.010481f
C198 VTAIL.n33 VSUBS 0.024772f
C199 VTAIL.n34 VSUBS 0.011097f
C200 VTAIL.n35 VSUBS 0.332771f
C201 VTAIL.n36 VSUBS 0.010481f
C202 VTAIL.t0 VSUBS 0.054315f
C203 VTAIL.n37 VSUBS 0.079957f
C204 VTAIL.n38 VSUBS 0.015694f
C205 VTAIL.n39 VSUBS 0.018579f
C206 VTAIL.n40 VSUBS 0.024772f
C207 VTAIL.n41 VSUBS 0.011097f
C208 VTAIL.n42 VSUBS 0.010481f
C209 VTAIL.n43 VSUBS 0.019504f
C210 VTAIL.n44 VSUBS 0.019504f
C211 VTAIL.n45 VSUBS 0.010481f
C212 VTAIL.n46 VSUBS 0.011097f
C213 VTAIL.n47 VSUBS 0.024772f
C214 VTAIL.n48 VSUBS 0.062228f
C215 VTAIL.n49 VSUBS 0.011097f
C216 VTAIL.n50 VSUBS 0.010481f
C217 VTAIL.n51 VSUBS 0.049612f
C218 VTAIL.n52 VSUBS 0.031528f
C219 VTAIL.n53 VSUBS 0.13164f
C220 VTAIL.t6 VSUBS 0.072902f
C221 VTAIL.t9 VSUBS 0.072902f
C222 VTAIL.n54 VSUBS 0.398253f
C223 VTAIL.n55 VSUBS 0.430963f
C224 VTAIL.n56 VSUBS 0.022093f
C225 VTAIL.n57 VSUBS 0.019504f
C226 VTAIL.n58 VSUBS 0.010481f
C227 VTAIL.n59 VSUBS 0.024772f
C228 VTAIL.n60 VSUBS 0.011097f
C229 VTAIL.n61 VSUBS 0.332771f
C230 VTAIL.n62 VSUBS 0.010481f
C231 VTAIL.t8 VSUBS 0.054315f
C232 VTAIL.n63 VSUBS 0.079957f
C233 VTAIL.n64 VSUBS 0.015694f
C234 VTAIL.n65 VSUBS 0.018579f
C235 VTAIL.n66 VSUBS 0.024772f
C236 VTAIL.n67 VSUBS 0.011097f
C237 VTAIL.n68 VSUBS 0.010481f
C238 VTAIL.n69 VSUBS 0.019504f
C239 VTAIL.n70 VSUBS 0.019504f
C240 VTAIL.n71 VSUBS 0.010481f
C241 VTAIL.n72 VSUBS 0.011097f
C242 VTAIL.n73 VSUBS 0.024772f
C243 VTAIL.n74 VSUBS 0.062228f
C244 VTAIL.n75 VSUBS 0.011097f
C245 VTAIL.n76 VSUBS 0.010481f
C246 VTAIL.n77 VSUBS 0.049612f
C247 VTAIL.n78 VSUBS 0.031528f
C248 VTAIL.n79 VSUBS 0.650947f
C249 VTAIL.n80 VSUBS 0.022093f
C250 VTAIL.n81 VSUBS 0.019504f
C251 VTAIL.n82 VSUBS 0.010481f
C252 VTAIL.n83 VSUBS 0.024772f
C253 VTAIL.n84 VSUBS 0.011097f
C254 VTAIL.n85 VSUBS 0.332771f
C255 VTAIL.n86 VSUBS 0.010481f
C256 VTAIL.t4 VSUBS 0.054315f
C257 VTAIL.n87 VSUBS 0.079957f
C258 VTAIL.n88 VSUBS 0.015694f
C259 VTAIL.n89 VSUBS 0.018579f
C260 VTAIL.n90 VSUBS 0.024772f
C261 VTAIL.n91 VSUBS 0.011097f
C262 VTAIL.n92 VSUBS 0.010481f
C263 VTAIL.n93 VSUBS 0.019504f
C264 VTAIL.n94 VSUBS 0.019504f
C265 VTAIL.n95 VSUBS 0.010481f
C266 VTAIL.n96 VSUBS 0.011097f
C267 VTAIL.n97 VSUBS 0.024772f
C268 VTAIL.n98 VSUBS 0.062228f
C269 VTAIL.n99 VSUBS 0.011097f
C270 VTAIL.n100 VSUBS 0.010481f
C271 VTAIL.n101 VSUBS 0.049612f
C272 VTAIL.n102 VSUBS 0.031528f
C273 VTAIL.n103 VSUBS 0.633475f
C274 VP.n0 VSUBS 0.055906f
C275 VP.n1 VSUBS 0.012686f
C276 VP.n2 VSUBS 0.230434f
C277 VP.t5 VSUBS 0.5344f
C278 VP.t4 VSUBS 0.5344f
C279 VP.t2 VSUBS 0.557614f
C280 VP.n3 VSUBS 0.246905f
C281 VP.n4 VSUBS 0.269679f
C282 VP.n5 VSUBS 0.012686f
C283 VP.n6 VSUBS 0.26067f
C284 VP.n7 VSUBS 1.72502f
C285 VP.t1 VSUBS 0.5344f
C286 VP.n8 VSUBS 0.26067f
C287 VP.n9 VSUBS 1.7814f
C288 VP.n10 VSUBS 0.055906f
C289 VP.n11 VSUBS 0.055906f
C290 VP.t3 VSUBS 0.5344f
C291 VP.n12 VSUBS 0.265324f
C292 VP.n13 VSUBS 0.012686f
C293 VP.t0 VSUBS 0.5344f
C294 VP.n14 VSUBS 0.26067f
C295 VP.n15 VSUBS 0.043325f
C296 B.n0 VSUBS 0.004448f
C297 B.n1 VSUBS 0.004448f
C298 B.n2 VSUBS 0.007034f
C299 B.n3 VSUBS 0.007034f
C300 B.n4 VSUBS 0.007034f
C301 B.n5 VSUBS 0.007034f
C302 B.n6 VSUBS 0.007034f
C303 B.n7 VSUBS 0.007034f
C304 B.n8 VSUBS 0.007034f
C305 B.n9 VSUBS 0.007034f
C306 B.n10 VSUBS 0.007034f
C307 B.n11 VSUBS 0.007034f
C308 B.n12 VSUBS 0.0173f
C309 B.n13 VSUBS 0.007034f
C310 B.n14 VSUBS 0.007034f
C311 B.n15 VSUBS 0.007034f
C312 B.n16 VSUBS 0.007034f
C313 B.n17 VSUBS 0.007034f
C314 B.n18 VSUBS 0.007034f
C315 B.n19 VSUBS 0.007034f
C316 B.n20 VSUBS 0.007034f
C317 B.n21 VSUBS 0.007034f
C318 B.t2 VSUBS 0.069222f
C319 B.t1 VSUBS 0.077662f
C320 B.t0 VSUBS 0.144458f
C321 B.n22 VSUBS 0.139539f
C322 B.n23 VSUBS 0.123805f
C323 B.n24 VSUBS 0.016296f
C324 B.n25 VSUBS 0.007034f
C325 B.n26 VSUBS 0.007034f
C326 B.n27 VSUBS 0.007034f
C327 B.n28 VSUBS 0.007034f
C328 B.n29 VSUBS 0.007034f
C329 B.t11 VSUBS 0.069223f
C330 B.t10 VSUBS 0.077663f
C331 B.t9 VSUBS 0.144458f
C332 B.n30 VSUBS 0.139538f
C333 B.n31 VSUBS 0.123803f
C334 B.n32 VSUBS 0.007034f
C335 B.n33 VSUBS 0.007034f
C336 B.n34 VSUBS 0.007034f
C337 B.n35 VSUBS 0.007034f
C338 B.n36 VSUBS 0.007034f
C339 B.n37 VSUBS 0.007034f
C340 B.n38 VSUBS 0.007034f
C341 B.n39 VSUBS 0.007034f
C342 B.n40 VSUBS 0.007034f
C343 B.n41 VSUBS 0.0173f
C344 B.n42 VSUBS 0.007034f
C345 B.n43 VSUBS 0.007034f
C346 B.n44 VSUBS 0.007034f
C347 B.n45 VSUBS 0.007034f
C348 B.n46 VSUBS 0.007034f
C349 B.n47 VSUBS 0.007034f
C350 B.n48 VSUBS 0.007034f
C351 B.n49 VSUBS 0.007034f
C352 B.n50 VSUBS 0.007034f
C353 B.n51 VSUBS 0.007034f
C354 B.n52 VSUBS 0.007034f
C355 B.n53 VSUBS 0.007034f
C356 B.n54 VSUBS 0.007034f
C357 B.n55 VSUBS 0.007034f
C358 B.n56 VSUBS 0.007034f
C359 B.n57 VSUBS 0.007034f
C360 B.n58 VSUBS 0.007034f
C361 B.n59 VSUBS 0.007034f
C362 B.n60 VSUBS 0.007034f
C363 B.n61 VSUBS 0.007034f
C364 B.n62 VSUBS 0.0173f
C365 B.n63 VSUBS 0.007034f
C366 B.n64 VSUBS 0.007034f
C367 B.n65 VSUBS 0.007034f
C368 B.n66 VSUBS 0.007034f
C369 B.n67 VSUBS 0.007034f
C370 B.n68 VSUBS 0.007034f
C371 B.n69 VSUBS 0.007034f
C372 B.n70 VSUBS 0.007034f
C373 B.n71 VSUBS 0.007034f
C374 B.t4 VSUBS 0.069223f
C375 B.t5 VSUBS 0.077663f
C376 B.t3 VSUBS 0.144458f
C377 B.n72 VSUBS 0.139538f
C378 B.n73 VSUBS 0.123803f
C379 B.n74 VSUBS 0.016296f
C380 B.n75 VSUBS 0.007034f
C381 B.n76 VSUBS 0.007034f
C382 B.n77 VSUBS 0.007034f
C383 B.n78 VSUBS 0.007034f
C384 B.n79 VSUBS 0.007034f
C385 B.t7 VSUBS 0.069222f
C386 B.t8 VSUBS 0.077662f
C387 B.t6 VSUBS 0.144458f
C388 B.n80 VSUBS 0.139539f
C389 B.n81 VSUBS 0.123805f
C390 B.n82 VSUBS 0.007034f
C391 B.n83 VSUBS 0.007034f
C392 B.n84 VSUBS 0.007034f
C393 B.n85 VSUBS 0.007034f
C394 B.n86 VSUBS 0.007034f
C395 B.n87 VSUBS 0.007034f
C396 B.n88 VSUBS 0.007034f
C397 B.n89 VSUBS 0.007034f
C398 B.n90 VSUBS 0.007034f
C399 B.n91 VSUBS 0.0173f
C400 B.n92 VSUBS 0.007034f
C401 B.n93 VSUBS 0.007034f
C402 B.n94 VSUBS 0.007034f
C403 B.n95 VSUBS 0.007034f
C404 B.n96 VSUBS 0.007034f
C405 B.n97 VSUBS 0.007034f
C406 B.n98 VSUBS 0.007034f
C407 B.n99 VSUBS 0.007034f
C408 B.n100 VSUBS 0.007034f
C409 B.n101 VSUBS 0.007034f
C410 B.n102 VSUBS 0.007034f
C411 B.n103 VSUBS 0.007034f
C412 B.n104 VSUBS 0.007034f
C413 B.n105 VSUBS 0.007034f
C414 B.n106 VSUBS 0.007034f
C415 B.n107 VSUBS 0.007034f
C416 B.n108 VSUBS 0.007034f
C417 B.n109 VSUBS 0.007034f
C418 B.n110 VSUBS 0.007034f
C419 B.n111 VSUBS 0.007034f
C420 B.n112 VSUBS 0.007034f
C421 B.n113 VSUBS 0.007034f
C422 B.n114 VSUBS 0.007034f
C423 B.n115 VSUBS 0.007034f
C424 B.n116 VSUBS 0.007034f
C425 B.n117 VSUBS 0.007034f
C426 B.n118 VSUBS 0.007034f
C427 B.n119 VSUBS 0.007034f
C428 B.n120 VSUBS 0.007034f
C429 B.n121 VSUBS 0.007034f
C430 B.n122 VSUBS 0.007034f
C431 B.n123 VSUBS 0.007034f
C432 B.n124 VSUBS 0.007034f
C433 B.n125 VSUBS 0.007034f
C434 B.n126 VSUBS 0.007034f
C435 B.n127 VSUBS 0.007034f
C436 B.n128 VSUBS 0.016421f
C437 B.n129 VSUBS 0.016421f
C438 B.n130 VSUBS 0.0173f
C439 B.n131 VSUBS 0.007034f
C440 B.n132 VSUBS 0.007034f
C441 B.n133 VSUBS 0.007034f
C442 B.n134 VSUBS 0.007034f
C443 B.n135 VSUBS 0.007034f
C444 B.n136 VSUBS 0.007034f
C445 B.n137 VSUBS 0.007034f
C446 B.n138 VSUBS 0.007034f
C447 B.n139 VSUBS 0.007034f
C448 B.n140 VSUBS 0.007034f
C449 B.n141 VSUBS 0.007034f
C450 B.n142 VSUBS 0.007034f
C451 B.n143 VSUBS 0.007034f
C452 B.n144 VSUBS 0.007034f
C453 B.n145 VSUBS 0.007034f
C454 B.n146 VSUBS 0.007034f
C455 B.n147 VSUBS 0.007034f
C456 B.n148 VSUBS 0.007034f
C457 B.n149 VSUBS 0.007034f
C458 B.n150 VSUBS 0.007034f
C459 B.n151 VSUBS 0.007034f
C460 B.n152 VSUBS 0.007034f
C461 B.n153 VSUBS 0.007034f
C462 B.n154 VSUBS 0.007034f
C463 B.n155 VSUBS 0.007034f
C464 B.n156 VSUBS 0.007034f
C465 B.n157 VSUBS 0.007034f
C466 B.n158 VSUBS 0.007034f
C467 B.n159 VSUBS 0.00662f
C468 B.n160 VSUBS 0.016296f
C469 B.n161 VSUBS 0.003931f
C470 B.n162 VSUBS 0.007034f
C471 B.n163 VSUBS 0.007034f
C472 B.n164 VSUBS 0.007034f
C473 B.n165 VSUBS 0.007034f
C474 B.n166 VSUBS 0.007034f
C475 B.n167 VSUBS 0.007034f
C476 B.n168 VSUBS 0.007034f
C477 B.n169 VSUBS 0.007034f
C478 B.n170 VSUBS 0.007034f
C479 B.n171 VSUBS 0.007034f
C480 B.n172 VSUBS 0.007034f
C481 B.n173 VSUBS 0.007034f
C482 B.n174 VSUBS 0.003931f
C483 B.n175 VSUBS 0.007034f
C484 B.n176 VSUBS 0.007034f
C485 B.n177 VSUBS 0.00662f
C486 B.n178 VSUBS 0.007034f
C487 B.n179 VSUBS 0.007034f
C488 B.n180 VSUBS 0.007034f
C489 B.n181 VSUBS 0.007034f
C490 B.n182 VSUBS 0.007034f
C491 B.n183 VSUBS 0.007034f
C492 B.n184 VSUBS 0.007034f
C493 B.n185 VSUBS 0.007034f
C494 B.n186 VSUBS 0.007034f
C495 B.n187 VSUBS 0.007034f
C496 B.n188 VSUBS 0.007034f
C497 B.n189 VSUBS 0.007034f
C498 B.n190 VSUBS 0.007034f
C499 B.n191 VSUBS 0.007034f
C500 B.n192 VSUBS 0.007034f
C501 B.n193 VSUBS 0.007034f
C502 B.n194 VSUBS 0.007034f
C503 B.n195 VSUBS 0.007034f
C504 B.n196 VSUBS 0.007034f
C505 B.n197 VSUBS 0.007034f
C506 B.n198 VSUBS 0.007034f
C507 B.n199 VSUBS 0.007034f
C508 B.n200 VSUBS 0.007034f
C509 B.n201 VSUBS 0.007034f
C510 B.n202 VSUBS 0.007034f
C511 B.n203 VSUBS 0.007034f
C512 B.n204 VSUBS 0.007034f
C513 B.n205 VSUBS 0.0173f
C514 B.n206 VSUBS 0.016421f
C515 B.n207 VSUBS 0.016421f
C516 B.n208 VSUBS 0.007034f
C517 B.n209 VSUBS 0.007034f
C518 B.n210 VSUBS 0.007034f
C519 B.n211 VSUBS 0.007034f
C520 B.n212 VSUBS 0.007034f
C521 B.n213 VSUBS 0.007034f
C522 B.n214 VSUBS 0.007034f
C523 B.n215 VSUBS 0.007034f
C524 B.n216 VSUBS 0.007034f
C525 B.n217 VSUBS 0.007034f
C526 B.n218 VSUBS 0.007034f
C527 B.n219 VSUBS 0.007034f
C528 B.n220 VSUBS 0.007034f
C529 B.n221 VSUBS 0.007034f
C530 B.n222 VSUBS 0.007034f
C531 B.n223 VSUBS 0.007034f
C532 B.n224 VSUBS 0.007034f
C533 B.n225 VSUBS 0.007034f
C534 B.n226 VSUBS 0.007034f
C535 B.n227 VSUBS 0.007034f
C536 B.n228 VSUBS 0.007034f
C537 B.n229 VSUBS 0.007034f
C538 B.n230 VSUBS 0.007034f
C539 B.n231 VSUBS 0.007034f
C540 B.n232 VSUBS 0.007034f
C541 B.n233 VSUBS 0.007034f
C542 B.n234 VSUBS 0.007034f
C543 B.n235 VSUBS 0.007034f
C544 B.n236 VSUBS 0.007034f
C545 B.n237 VSUBS 0.007034f
C546 B.n238 VSUBS 0.007034f
C547 B.n239 VSUBS 0.007034f
C548 B.n240 VSUBS 0.007034f
C549 B.n241 VSUBS 0.007034f
C550 B.n242 VSUBS 0.007034f
C551 B.n243 VSUBS 0.007034f
C552 B.n244 VSUBS 0.007034f
C553 B.n245 VSUBS 0.007034f
C554 B.n246 VSUBS 0.007034f
C555 B.n247 VSUBS 0.007034f
C556 B.n248 VSUBS 0.007034f
C557 B.n249 VSUBS 0.007034f
C558 B.n250 VSUBS 0.007034f
C559 B.n251 VSUBS 0.007034f
C560 B.n252 VSUBS 0.007034f
C561 B.n253 VSUBS 0.007034f
C562 B.n254 VSUBS 0.007034f
C563 B.n255 VSUBS 0.007034f
C564 B.n256 VSUBS 0.007034f
C565 B.n257 VSUBS 0.007034f
C566 B.n258 VSUBS 0.007034f
C567 B.n259 VSUBS 0.007034f
C568 B.n260 VSUBS 0.007034f
C569 B.n261 VSUBS 0.007034f
C570 B.n262 VSUBS 0.007034f
C571 B.n263 VSUBS 0.007034f
C572 B.n264 VSUBS 0.007034f
C573 B.n265 VSUBS 0.007034f
C574 B.n266 VSUBS 0.016421f
C575 B.n267 VSUBS 0.017222f
C576 B.n268 VSUBS 0.016499f
C577 B.n269 VSUBS 0.007034f
C578 B.n270 VSUBS 0.007034f
C579 B.n271 VSUBS 0.007034f
C580 B.n272 VSUBS 0.007034f
C581 B.n273 VSUBS 0.007034f
C582 B.n274 VSUBS 0.007034f
C583 B.n275 VSUBS 0.007034f
C584 B.n276 VSUBS 0.007034f
C585 B.n277 VSUBS 0.007034f
C586 B.n278 VSUBS 0.007034f
C587 B.n279 VSUBS 0.007034f
C588 B.n280 VSUBS 0.007034f
C589 B.n281 VSUBS 0.007034f
C590 B.n282 VSUBS 0.007034f
C591 B.n283 VSUBS 0.007034f
C592 B.n284 VSUBS 0.007034f
C593 B.n285 VSUBS 0.007034f
C594 B.n286 VSUBS 0.007034f
C595 B.n287 VSUBS 0.007034f
C596 B.n288 VSUBS 0.007034f
C597 B.n289 VSUBS 0.007034f
C598 B.n290 VSUBS 0.007034f
C599 B.n291 VSUBS 0.007034f
C600 B.n292 VSUBS 0.007034f
C601 B.n293 VSUBS 0.007034f
C602 B.n294 VSUBS 0.007034f
C603 B.n295 VSUBS 0.007034f
C604 B.n296 VSUBS 0.007034f
C605 B.n297 VSUBS 0.00662f
C606 B.n298 VSUBS 0.016296f
C607 B.n299 VSUBS 0.003931f
C608 B.n300 VSUBS 0.007034f
C609 B.n301 VSUBS 0.007034f
C610 B.n302 VSUBS 0.007034f
C611 B.n303 VSUBS 0.007034f
C612 B.n304 VSUBS 0.007034f
C613 B.n305 VSUBS 0.007034f
C614 B.n306 VSUBS 0.007034f
C615 B.n307 VSUBS 0.007034f
C616 B.n308 VSUBS 0.007034f
C617 B.n309 VSUBS 0.007034f
C618 B.n310 VSUBS 0.007034f
C619 B.n311 VSUBS 0.007034f
C620 B.n312 VSUBS 0.003931f
C621 B.n313 VSUBS 0.007034f
C622 B.n314 VSUBS 0.007034f
C623 B.n315 VSUBS 0.00662f
C624 B.n316 VSUBS 0.007034f
C625 B.n317 VSUBS 0.007034f
C626 B.n318 VSUBS 0.007034f
C627 B.n319 VSUBS 0.007034f
C628 B.n320 VSUBS 0.007034f
C629 B.n321 VSUBS 0.007034f
C630 B.n322 VSUBS 0.007034f
C631 B.n323 VSUBS 0.007034f
C632 B.n324 VSUBS 0.007034f
C633 B.n325 VSUBS 0.007034f
C634 B.n326 VSUBS 0.007034f
C635 B.n327 VSUBS 0.007034f
C636 B.n328 VSUBS 0.007034f
C637 B.n329 VSUBS 0.007034f
C638 B.n330 VSUBS 0.007034f
C639 B.n331 VSUBS 0.007034f
C640 B.n332 VSUBS 0.007034f
C641 B.n333 VSUBS 0.007034f
C642 B.n334 VSUBS 0.007034f
C643 B.n335 VSUBS 0.007034f
C644 B.n336 VSUBS 0.007034f
C645 B.n337 VSUBS 0.007034f
C646 B.n338 VSUBS 0.007034f
C647 B.n339 VSUBS 0.007034f
C648 B.n340 VSUBS 0.007034f
C649 B.n341 VSUBS 0.007034f
C650 B.n342 VSUBS 0.007034f
C651 B.n343 VSUBS 0.0173f
C652 B.n344 VSUBS 0.016421f
C653 B.n345 VSUBS 0.016421f
C654 B.n346 VSUBS 0.007034f
C655 B.n347 VSUBS 0.007034f
C656 B.n348 VSUBS 0.007034f
C657 B.n349 VSUBS 0.007034f
C658 B.n350 VSUBS 0.007034f
C659 B.n351 VSUBS 0.007034f
C660 B.n352 VSUBS 0.007034f
C661 B.n353 VSUBS 0.007034f
C662 B.n354 VSUBS 0.007034f
C663 B.n355 VSUBS 0.007034f
C664 B.n356 VSUBS 0.007034f
C665 B.n357 VSUBS 0.007034f
C666 B.n358 VSUBS 0.007034f
C667 B.n359 VSUBS 0.007034f
C668 B.n360 VSUBS 0.007034f
C669 B.n361 VSUBS 0.007034f
C670 B.n362 VSUBS 0.007034f
C671 B.n363 VSUBS 0.007034f
C672 B.n364 VSUBS 0.007034f
C673 B.n365 VSUBS 0.007034f
C674 B.n366 VSUBS 0.007034f
C675 B.n367 VSUBS 0.007034f
C676 B.n368 VSUBS 0.007034f
C677 B.n369 VSUBS 0.007034f
C678 B.n370 VSUBS 0.007034f
C679 B.n371 VSUBS 0.007034f
C680 B.n372 VSUBS 0.007034f
C681 B.n373 VSUBS 0.007034f
C682 B.n374 VSUBS 0.007034f
C683 B.n375 VSUBS 0.015927f
.ends

