* NGSPICE file created from diff_pair_sample_0193.ext - technology: sky130A

.subckt diff_pair_sample_0193 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t9 VP.t0 VTAIL.t13 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=3.6504 ps=19.5 w=9.36 l=3.81
X1 B.t23 B.t21 B.t22 B.t18 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=0 ps=0 w=9.36 l=3.81
X2 VTAIL.t5 VN.t0 VDD2.t9 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X3 VTAIL.t6 VN.t1 VDD2.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X4 VTAIL.t12 VP.t1 VDD1.t8 B.t6 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X5 VDD1.t7 VP.t2 VTAIL.t14 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X6 VTAIL.t2 VN.t2 VDD2.t7 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X7 VTAIL.t3 VN.t3 VDD2.t6 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X8 VDD2.t5 VN.t4 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X9 VDD1.t6 VP.t3 VTAIL.t18 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X10 VTAIL.t15 VP.t4 VDD1.t5 B.t3 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X11 VDD2.t4 VN.t5 VTAIL.t8 B.t8 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=1.5444 ps=9.69 w=9.36 l=3.81
X12 B.t20 B.t17 B.t19 B.t18 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=0 ps=0 w=9.36 l=3.81
X13 VDD1.t4 VP.t5 VTAIL.t17 B.t4 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=1.5444 ps=9.69 w=9.36 l=3.81
X14 VDD2.t3 VN.t6 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=3.6504 ps=19.5 w=9.36 l=3.81
X15 B.t16 B.t14 B.t15 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=0 ps=0 w=9.36 l=3.81
X16 B.t13 B.t10 B.t12 B.t11 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=0 ps=0 w=9.36 l=3.81
X17 VDD2.t2 VN.t7 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X18 VDD2.t1 VN.t8 VTAIL.t9 B.t9 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=3.6504 ps=19.5 w=9.36 l=3.81
X19 VTAIL.t19 VP.t6 VDD1.t3 B.t2 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X20 VDD1.t2 VP.t7 VTAIL.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=1.5444 ps=9.69 w=9.36 l=3.81
X21 VDD1.t1 VP.t8 VTAIL.t11 B.t9 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=3.6504 ps=19.5 w=9.36 l=3.81
X22 VTAIL.t10 VP.t9 VDD1.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.5444 pd=9.69 as=1.5444 ps=9.69 w=9.36 l=3.81
X23 VDD2.t0 VN.t9 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.6504 pd=19.5 as=1.5444 ps=9.69 w=9.36 l=3.81
R0 VP.n34 VP.n33 161.3
R1 VP.n35 VP.n30 161.3
R2 VP.n37 VP.n36 161.3
R3 VP.n38 VP.n29 161.3
R4 VP.n40 VP.n39 161.3
R5 VP.n41 VP.n28 161.3
R6 VP.n43 VP.n42 161.3
R7 VP.n44 VP.n27 161.3
R8 VP.n47 VP.n46 161.3
R9 VP.n48 VP.n26 161.3
R10 VP.n50 VP.n49 161.3
R11 VP.n51 VP.n25 161.3
R12 VP.n53 VP.n52 161.3
R13 VP.n54 VP.n24 161.3
R14 VP.n56 VP.n55 161.3
R15 VP.n57 VP.n23 161.3
R16 VP.n60 VP.n59 161.3
R17 VP.n61 VP.n22 161.3
R18 VP.n63 VP.n62 161.3
R19 VP.n64 VP.n21 161.3
R20 VP.n66 VP.n65 161.3
R21 VP.n67 VP.n20 161.3
R22 VP.n69 VP.n68 161.3
R23 VP.n70 VP.n19 161.3
R24 VP.n72 VP.n71 161.3
R25 VP.n129 VP.n128 161.3
R26 VP.n127 VP.n1 161.3
R27 VP.n126 VP.n125 161.3
R28 VP.n124 VP.n2 161.3
R29 VP.n123 VP.n122 161.3
R30 VP.n121 VP.n3 161.3
R31 VP.n120 VP.n119 161.3
R32 VP.n118 VP.n4 161.3
R33 VP.n117 VP.n116 161.3
R34 VP.n114 VP.n5 161.3
R35 VP.n113 VP.n112 161.3
R36 VP.n111 VP.n6 161.3
R37 VP.n110 VP.n109 161.3
R38 VP.n108 VP.n7 161.3
R39 VP.n107 VP.n106 161.3
R40 VP.n105 VP.n8 161.3
R41 VP.n104 VP.n103 161.3
R42 VP.n101 VP.n9 161.3
R43 VP.n100 VP.n99 161.3
R44 VP.n98 VP.n10 161.3
R45 VP.n97 VP.n96 161.3
R46 VP.n95 VP.n11 161.3
R47 VP.n94 VP.n93 161.3
R48 VP.n92 VP.n12 161.3
R49 VP.n91 VP.n90 161.3
R50 VP.n88 VP.n13 161.3
R51 VP.n87 VP.n86 161.3
R52 VP.n85 VP.n14 161.3
R53 VP.n84 VP.n83 161.3
R54 VP.n82 VP.n15 161.3
R55 VP.n81 VP.n80 161.3
R56 VP.n79 VP.n16 161.3
R57 VP.n78 VP.n77 161.3
R58 VP.n76 VP.n17 161.3
R59 VP.n31 VP.t5 91.7699
R60 VP.n75 VP.n74 88.77
R61 VP.n130 VP.n0 88.77
R62 VP.n73 VP.n18 88.77
R63 VP.n75 VP.t7 59.2068
R64 VP.n89 VP.t6 59.2068
R65 VP.n102 VP.t3 59.2068
R66 VP.n115 VP.t1 59.2068
R67 VP.n0 VP.t0 59.2068
R68 VP.n18 VP.t8 59.2068
R69 VP.n58 VP.t4 59.2068
R70 VP.n45 VP.t2 59.2068
R71 VP.n32 VP.t9 59.2068
R72 VP.n74 VP.n73 57.7268
R73 VP.n96 VP.n95 56.5617
R74 VP.n109 VP.n108 56.5617
R75 VP.n52 VP.n51 56.5617
R76 VP.n39 VP.n38 56.5617
R77 VP.n32 VP.n31 56.1007
R78 VP.n83 VP.n82 44.4521
R79 VP.n122 VP.n121 44.4521
R80 VP.n65 VP.n64 44.4521
R81 VP.n82 VP.n81 36.702
R82 VP.n122 VP.n2 36.702
R83 VP.n65 VP.n20 36.702
R84 VP.n77 VP.n76 24.5923
R85 VP.n77 VP.n16 24.5923
R86 VP.n81 VP.n16 24.5923
R87 VP.n83 VP.n14 24.5923
R88 VP.n87 VP.n14 24.5923
R89 VP.n88 VP.n87 24.5923
R90 VP.n90 VP.n12 24.5923
R91 VP.n94 VP.n12 24.5923
R92 VP.n95 VP.n94 24.5923
R93 VP.n96 VP.n10 24.5923
R94 VP.n100 VP.n10 24.5923
R95 VP.n101 VP.n100 24.5923
R96 VP.n103 VP.n8 24.5923
R97 VP.n107 VP.n8 24.5923
R98 VP.n108 VP.n107 24.5923
R99 VP.n109 VP.n6 24.5923
R100 VP.n113 VP.n6 24.5923
R101 VP.n114 VP.n113 24.5923
R102 VP.n116 VP.n4 24.5923
R103 VP.n120 VP.n4 24.5923
R104 VP.n121 VP.n120 24.5923
R105 VP.n126 VP.n2 24.5923
R106 VP.n127 VP.n126 24.5923
R107 VP.n128 VP.n127 24.5923
R108 VP.n69 VP.n20 24.5923
R109 VP.n70 VP.n69 24.5923
R110 VP.n71 VP.n70 24.5923
R111 VP.n52 VP.n24 24.5923
R112 VP.n56 VP.n24 24.5923
R113 VP.n57 VP.n56 24.5923
R114 VP.n59 VP.n22 24.5923
R115 VP.n63 VP.n22 24.5923
R116 VP.n64 VP.n63 24.5923
R117 VP.n39 VP.n28 24.5923
R118 VP.n43 VP.n28 24.5923
R119 VP.n44 VP.n43 24.5923
R120 VP.n46 VP.n26 24.5923
R121 VP.n50 VP.n26 24.5923
R122 VP.n51 VP.n50 24.5923
R123 VP.n33 VP.n30 24.5923
R124 VP.n37 VP.n30 24.5923
R125 VP.n38 VP.n37 24.5923
R126 VP.n90 VP.n89 19.1821
R127 VP.n115 VP.n114 19.1821
R128 VP.n58 VP.n57 19.1821
R129 VP.n33 VP.n32 19.1821
R130 VP.n102 VP.n101 12.2964
R131 VP.n103 VP.n102 12.2964
R132 VP.n45 VP.n44 12.2964
R133 VP.n46 VP.n45 12.2964
R134 VP.n89 VP.n88 5.4107
R135 VP.n116 VP.n115 5.4107
R136 VP.n59 VP.n58 5.4107
R137 VP.n34 VP.n31 2.48416
R138 VP.n76 VP.n75 1.47601
R139 VP.n128 VP.n0 1.47601
R140 VP.n71 VP.n18 1.47601
R141 VP.n73 VP.n72 0.354861
R142 VP.n74 VP.n17 0.354861
R143 VP.n130 VP.n129 0.354861
R144 VP VP.n130 0.267071
R145 VP.n35 VP.n34 0.189894
R146 VP.n36 VP.n35 0.189894
R147 VP.n36 VP.n29 0.189894
R148 VP.n40 VP.n29 0.189894
R149 VP.n41 VP.n40 0.189894
R150 VP.n42 VP.n41 0.189894
R151 VP.n42 VP.n27 0.189894
R152 VP.n47 VP.n27 0.189894
R153 VP.n48 VP.n47 0.189894
R154 VP.n49 VP.n48 0.189894
R155 VP.n49 VP.n25 0.189894
R156 VP.n53 VP.n25 0.189894
R157 VP.n54 VP.n53 0.189894
R158 VP.n55 VP.n54 0.189894
R159 VP.n55 VP.n23 0.189894
R160 VP.n60 VP.n23 0.189894
R161 VP.n61 VP.n60 0.189894
R162 VP.n62 VP.n61 0.189894
R163 VP.n62 VP.n21 0.189894
R164 VP.n66 VP.n21 0.189894
R165 VP.n67 VP.n66 0.189894
R166 VP.n68 VP.n67 0.189894
R167 VP.n68 VP.n19 0.189894
R168 VP.n72 VP.n19 0.189894
R169 VP.n78 VP.n17 0.189894
R170 VP.n79 VP.n78 0.189894
R171 VP.n80 VP.n79 0.189894
R172 VP.n80 VP.n15 0.189894
R173 VP.n84 VP.n15 0.189894
R174 VP.n85 VP.n84 0.189894
R175 VP.n86 VP.n85 0.189894
R176 VP.n86 VP.n13 0.189894
R177 VP.n91 VP.n13 0.189894
R178 VP.n92 VP.n91 0.189894
R179 VP.n93 VP.n92 0.189894
R180 VP.n93 VP.n11 0.189894
R181 VP.n97 VP.n11 0.189894
R182 VP.n98 VP.n97 0.189894
R183 VP.n99 VP.n98 0.189894
R184 VP.n99 VP.n9 0.189894
R185 VP.n104 VP.n9 0.189894
R186 VP.n105 VP.n104 0.189894
R187 VP.n106 VP.n105 0.189894
R188 VP.n106 VP.n7 0.189894
R189 VP.n110 VP.n7 0.189894
R190 VP.n111 VP.n110 0.189894
R191 VP.n112 VP.n111 0.189894
R192 VP.n112 VP.n5 0.189894
R193 VP.n117 VP.n5 0.189894
R194 VP.n118 VP.n117 0.189894
R195 VP.n119 VP.n118 0.189894
R196 VP.n119 VP.n3 0.189894
R197 VP.n123 VP.n3 0.189894
R198 VP.n124 VP.n123 0.189894
R199 VP.n125 VP.n124 0.189894
R200 VP.n125 VP.n1 0.189894
R201 VP.n129 VP.n1 0.189894
R202 VTAIL.n208 VTAIL.n164 289.615
R203 VTAIL.n46 VTAIL.n2 289.615
R204 VTAIL.n158 VTAIL.n114 289.615
R205 VTAIL.n104 VTAIL.n60 289.615
R206 VTAIL.n181 VTAIL.n180 185
R207 VTAIL.n183 VTAIL.n182 185
R208 VTAIL.n176 VTAIL.n175 185
R209 VTAIL.n189 VTAIL.n188 185
R210 VTAIL.n191 VTAIL.n190 185
R211 VTAIL.n172 VTAIL.n171 185
R212 VTAIL.n198 VTAIL.n197 185
R213 VTAIL.n199 VTAIL.n170 185
R214 VTAIL.n201 VTAIL.n200 185
R215 VTAIL.n168 VTAIL.n167 185
R216 VTAIL.n207 VTAIL.n206 185
R217 VTAIL.n209 VTAIL.n208 185
R218 VTAIL.n19 VTAIL.n18 185
R219 VTAIL.n21 VTAIL.n20 185
R220 VTAIL.n14 VTAIL.n13 185
R221 VTAIL.n27 VTAIL.n26 185
R222 VTAIL.n29 VTAIL.n28 185
R223 VTAIL.n10 VTAIL.n9 185
R224 VTAIL.n36 VTAIL.n35 185
R225 VTAIL.n37 VTAIL.n8 185
R226 VTAIL.n39 VTAIL.n38 185
R227 VTAIL.n6 VTAIL.n5 185
R228 VTAIL.n45 VTAIL.n44 185
R229 VTAIL.n47 VTAIL.n46 185
R230 VTAIL.n159 VTAIL.n158 185
R231 VTAIL.n157 VTAIL.n156 185
R232 VTAIL.n118 VTAIL.n117 185
R233 VTAIL.n122 VTAIL.n120 185
R234 VTAIL.n151 VTAIL.n150 185
R235 VTAIL.n149 VTAIL.n148 185
R236 VTAIL.n124 VTAIL.n123 185
R237 VTAIL.n143 VTAIL.n142 185
R238 VTAIL.n141 VTAIL.n140 185
R239 VTAIL.n128 VTAIL.n127 185
R240 VTAIL.n135 VTAIL.n134 185
R241 VTAIL.n133 VTAIL.n132 185
R242 VTAIL.n105 VTAIL.n104 185
R243 VTAIL.n103 VTAIL.n102 185
R244 VTAIL.n64 VTAIL.n63 185
R245 VTAIL.n68 VTAIL.n66 185
R246 VTAIL.n97 VTAIL.n96 185
R247 VTAIL.n95 VTAIL.n94 185
R248 VTAIL.n70 VTAIL.n69 185
R249 VTAIL.n89 VTAIL.n88 185
R250 VTAIL.n87 VTAIL.n86 185
R251 VTAIL.n74 VTAIL.n73 185
R252 VTAIL.n81 VTAIL.n80 185
R253 VTAIL.n79 VTAIL.n78 185
R254 VTAIL.n179 VTAIL.t9 149.524
R255 VTAIL.n17 VTAIL.t13 149.524
R256 VTAIL.n131 VTAIL.t11 149.524
R257 VTAIL.n77 VTAIL.t0 149.524
R258 VTAIL.n182 VTAIL.n181 104.615
R259 VTAIL.n182 VTAIL.n175 104.615
R260 VTAIL.n189 VTAIL.n175 104.615
R261 VTAIL.n190 VTAIL.n189 104.615
R262 VTAIL.n190 VTAIL.n171 104.615
R263 VTAIL.n198 VTAIL.n171 104.615
R264 VTAIL.n199 VTAIL.n198 104.615
R265 VTAIL.n200 VTAIL.n199 104.615
R266 VTAIL.n200 VTAIL.n167 104.615
R267 VTAIL.n207 VTAIL.n167 104.615
R268 VTAIL.n208 VTAIL.n207 104.615
R269 VTAIL.n20 VTAIL.n19 104.615
R270 VTAIL.n20 VTAIL.n13 104.615
R271 VTAIL.n27 VTAIL.n13 104.615
R272 VTAIL.n28 VTAIL.n27 104.615
R273 VTAIL.n28 VTAIL.n9 104.615
R274 VTAIL.n36 VTAIL.n9 104.615
R275 VTAIL.n37 VTAIL.n36 104.615
R276 VTAIL.n38 VTAIL.n37 104.615
R277 VTAIL.n38 VTAIL.n5 104.615
R278 VTAIL.n45 VTAIL.n5 104.615
R279 VTAIL.n46 VTAIL.n45 104.615
R280 VTAIL.n158 VTAIL.n157 104.615
R281 VTAIL.n157 VTAIL.n117 104.615
R282 VTAIL.n122 VTAIL.n117 104.615
R283 VTAIL.n150 VTAIL.n122 104.615
R284 VTAIL.n150 VTAIL.n149 104.615
R285 VTAIL.n149 VTAIL.n123 104.615
R286 VTAIL.n142 VTAIL.n123 104.615
R287 VTAIL.n142 VTAIL.n141 104.615
R288 VTAIL.n141 VTAIL.n127 104.615
R289 VTAIL.n134 VTAIL.n127 104.615
R290 VTAIL.n134 VTAIL.n133 104.615
R291 VTAIL.n104 VTAIL.n103 104.615
R292 VTAIL.n103 VTAIL.n63 104.615
R293 VTAIL.n68 VTAIL.n63 104.615
R294 VTAIL.n96 VTAIL.n68 104.615
R295 VTAIL.n96 VTAIL.n95 104.615
R296 VTAIL.n95 VTAIL.n69 104.615
R297 VTAIL.n88 VTAIL.n69 104.615
R298 VTAIL.n88 VTAIL.n87 104.615
R299 VTAIL.n87 VTAIL.n73 104.615
R300 VTAIL.n80 VTAIL.n73 104.615
R301 VTAIL.n80 VTAIL.n79 104.615
R302 VTAIL.n181 VTAIL.t9 52.3082
R303 VTAIL.n19 VTAIL.t13 52.3082
R304 VTAIL.n133 VTAIL.t11 52.3082
R305 VTAIL.n79 VTAIL.t0 52.3082
R306 VTAIL.n113 VTAIL.n112 48.6505
R307 VTAIL.n111 VTAIL.n110 48.6505
R308 VTAIL.n59 VTAIL.n58 48.6505
R309 VTAIL.n57 VTAIL.n56 48.6505
R310 VTAIL.n215 VTAIL.n214 48.6504
R311 VTAIL.n1 VTAIL.n0 48.6504
R312 VTAIL.n53 VTAIL.n52 48.6504
R313 VTAIL.n55 VTAIL.n54 48.6504
R314 VTAIL.n213 VTAIL.n212 34.5126
R315 VTAIL.n51 VTAIL.n50 34.5126
R316 VTAIL.n163 VTAIL.n162 34.5126
R317 VTAIL.n109 VTAIL.n108 34.5126
R318 VTAIL.n57 VTAIL.n55 27.5738
R319 VTAIL.n213 VTAIL.n163 24.0048
R320 VTAIL.n201 VTAIL.n168 13.1884
R321 VTAIL.n39 VTAIL.n6 13.1884
R322 VTAIL.n120 VTAIL.n118 13.1884
R323 VTAIL.n66 VTAIL.n64 13.1884
R324 VTAIL.n202 VTAIL.n170 12.8005
R325 VTAIL.n206 VTAIL.n205 12.8005
R326 VTAIL.n40 VTAIL.n8 12.8005
R327 VTAIL.n44 VTAIL.n43 12.8005
R328 VTAIL.n156 VTAIL.n155 12.8005
R329 VTAIL.n152 VTAIL.n151 12.8005
R330 VTAIL.n102 VTAIL.n101 12.8005
R331 VTAIL.n98 VTAIL.n97 12.8005
R332 VTAIL.n197 VTAIL.n196 12.0247
R333 VTAIL.n209 VTAIL.n166 12.0247
R334 VTAIL.n35 VTAIL.n34 12.0247
R335 VTAIL.n47 VTAIL.n4 12.0247
R336 VTAIL.n159 VTAIL.n116 12.0247
R337 VTAIL.n148 VTAIL.n121 12.0247
R338 VTAIL.n105 VTAIL.n62 12.0247
R339 VTAIL.n94 VTAIL.n67 12.0247
R340 VTAIL.n195 VTAIL.n172 11.249
R341 VTAIL.n210 VTAIL.n164 11.249
R342 VTAIL.n33 VTAIL.n10 11.249
R343 VTAIL.n48 VTAIL.n2 11.249
R344 VTAIL.n160 VTAIL.n114 11.249
R345 VTAIL.n147 VTAIL.n124 11.249
R346 VTAIL.n106 VTAIL.n60 11.249
R347 VTAIL.n93 VTAIL.n70 11.249
R348 VTAIL.n192 VTAIL.n191 10.4732
R349 VTAIL.n30 VTAIL.n29 10.4732
R350 VTAIL.n144 VTAIL.n143 10.4732
R351 VTAIL.n90 VTAIL.n89 10.4732
R352 VTAIL.n180 VTAIL.n179 10.2747
R353 VTAIL.n18 VTAIL.n17 10.2747
R354 VTAIL.n132 VTAIL.n131 10.2747
R355 VTAIL.n78 VTAIL.n77 10.2747
R356 VTAIL.n188 VTAIL.n174 9.69747
R357 VTAIL.n26 VTAIL.n12 9.69747
R358 VTAIL.n140 VTAIL.n126 9.69747
R359 VTAIL.n86 VTAIL.n72 9.69747
R360 VTAIL.n212 VTAIL.n211 9.45567
R361 VTAIL.n50 VTAIL.n49 9.45567
R362 VTAIL.n162 VTAIL.n161 9.45567
R363 VTAIL.n108 VTAIL.n107 9.45567
R364 VTAIL.n211 VTAIL.n210 9.3005
R365 VTAIL.n166 VTAIL.n165 9.3005
R366 VTAIL.n205 VTAIL.n204 9.3005
R367 VTAIL.n178 VTAIL.n177 9.3005
R368 VTAIL.n185 VTAIL.n184 9.3005
R369 VTAIL.n187 VTAIL.n186 9.3005
R370 VTAIL.n174 VTAIL.n173 9.3005
R371 VTAIL.n193 VTAIL.n192 9.3005
R372 VTAIL.n195 VTAIL.n194 9.3005
R373 VTAIL.n196 VTAIL.n169 9.3005
R374 VTAIL.n203 VTAIL.n202 9.3005
R375 VTAIL.n49 VTAIL.n48 9.3005
R376 VTAIL.n4 VTAIL.n3 9.3005
R377 VTAIL.n43 VTAIL.n42 9.3005
R378 VTAIL.n16 VTAIL.n15 9.3005
R379 VTAIL.n23 VTAIL.n22 9.3005
R380 VTAIL.n25 VTAIL.n24 9.3005
R381 VTAIL.n12 VTAIL.n11 9.3005
R382 VTAIL.n31 VTAIL.n30 9.3005
R383 VTAIL.n33 VTAIL.n32 9.3005
R384 VTAIL.n34 VTAIL.n7 9.3005
R385 VTAIL.n41 VTAIL.n40 9.3005
R386 VTAIL.n130 VTAIL.n129 9.3005
R387 VTAIL.n137 VTAIL.n136 9.3005
R388 VTAIL.n139 VTAIL.n138 9.3005
R389 VTAIL.n126 VTAIL.n125 9.3005
R390 VTAIL.n145 VTAIL.n144 9.3005
R391 VTAIL.n147 VTAIL.n146 9.3005
R392 VTAIL.n121 VTAIL.n119 9.3005
R393 VTAIL.n153 VTAIL.n152 9.3005
R394 VTAIL.n161 VTAIL.n160 9.3005
R395 VTAIL.n116 VTAIL.n115 9.3005
R396 VTAIL.n155 VTAIL.n154 9.3005
R397 VTAIL.n76 VTAIL.n75 9.3005
R398 VTAIL.n83 VTAIL.n82 9.3005
R399 VTAIL.n85 VTAIL.n84 9.3005
R400 VTAIL.n72 VTAIL.n71 9.3005
R401 VTAIL.n91 VTAIL.n90 9.3005
R402 VTAIL.n93 VTAIL.n92 9.3005
R403 VTAIL.n67 VTAIL.n65 9.3005
R404 VTAIL.n99 VTAIL.n98 9.3005
R405 VTAIL.n107 VTAIL.n106 9.3005
R406 VTAIL.n62 VTAIL.n61 9.3005
R407 VTAIL.n101 VTAIL.n100 9.3005
R408 VTAIL.n187 VTAIL.n176 8.92171
R409 VTAIL.n25 VTAIL.n14 8.92171
R410 VTAIL.n139 VTAIL.n128 8.92171
R411 VTAIL.n85 VTAIL.n74 8.92171
R412 VTAIL.n184 VTAIL.n183 8.14595
R413 VTAIL.n22 VTAIL.n21 8.14595
R414 VTAIL.n136 VTAIL.n135 8.14595
R415 VTAIL.n82 VTAIL.n81 8.14595
R416 VTAIL.n180 VTAIL.n178 7.3702
R417 VTAIL.n18 VTAIL.n16 7.3702
R418 VTAIL.n132 VTAIL.n130 7.3702
R419 VTAIL.n78 VTAIL.n76 7.3702
R420 VTAIL.n183 VTAIL.n178 5.81868
R421 VTAIL.n21 VTAIL.n16 5.81868
R422 VTAIL.n135 VTAIL.n130 5.81868
R423 VTAIL.n81 VTAIL.n76 5.81868
R424 VTAIL.n184 VTAIL.n176 5.04292
R425 VTAIL.n22 VTAIL.n14 5.04292
R426 VTAIL.n136 VTAIL.n128 5.04292
R427 VTAIL.n82 VTAIL.n74 5.04292
R428 VTAIL.n188 VTAIL.n187 4.26717
R429 VTAIL.n26 VTAIL.n25 4.26717
R430 VTAIL.n140 VTAIL.n139 4.26717
R431 VTAIL.n86 VTAIL.n85 4.26717
R432 VTAIL.n59 VTAIL.n57 3.56947
R433 VTAIL.n109 VTAIL.n59 3.56947
R434 VTAIL.n113 VTAIL.n111 3.56947
R435 VTAIL.n163 VTAIL.n113 3.56947
R436 VTAIL.n55 VTAIL.n53 3.56947
R437 VTAIL.n53 VTAIL.n51 3.56947
R438 VTAIL.n215 VTAIL.n213 3.56947
R439 VTAIL.n191 VTAIL.n174 3.49141
R440 VTAIL.n29 VTAIL.n12 3.49141
R441 VTAIL.n143 VTAIL.n126 3.49141
R442 VTAIL.n89 VTAIL.n72 3.49141
R443 VTAIL.n179 VTAIL.n177 2.84303
R444 VTAIL.n17 VTAIL.n15 2.84303
R445 VTAIL.n131 VTAIL.n129 2.84303
R446 VTAIL.n77 VTAIL.n75 2.84303
R447 VTAIL VTAIL.n1 2.73541
R448 VTAIL.n192 VTAIL.n172 2.71565
R449 VTAIL.n212 VTAIL.n164 2.71565
R450 VTAIL.n30 VTAIL.n10 2.71565
R451 VTAIL.n50 VTAIL.n2 2.71565
R452 VTAIL.n162 VTAIL.n114 2.71565
R453 VTAIL.n144 VTAIL.n124 2.71565
R454 VTAIL.n108 VTAIL.n60 2.71565
R455 VTAIL.n90 VTAIL.n70 2.71565
R456 VTAIL.n111 VTAIL.n109 2.25481
R457 VTAIL.n51 VTAIL.n1 2.25481
R458 VTAIL.n214 VTAIL.t1 2.11588
R459 VTAIL.n214 VTAIL.t3 2.11588
R460 VTAIL.n0 VTAIL.t4 2.11588
R461 VTAIL.n0 VTAIL.t5 2.11588
R462 VTAIL.n52 VTAIL.t18 2.11588
R463 VTAIL.n52 VTAIL.t12 2.11588
R464 VTAIL.n54 VTAIL.t16 2.11588
R465 VTAIL.n54 VTAIL.t19 2.11588
R466 VTAIL.n112 VTAIL.t14 2.11588
R467 VTAIL.n112 VTAIL.t15 2.11588
R468 VTAIL.n110 VTAIL.t17 2.11588
R469 VTAIL.n110 VTAIL.t10 2.11588
R470 VTAIL.n58 VTAIL.t7 2.11588
R471 VTAIL.n58 VTAIL.t6 2.11588
R472 VTAIL.n56 VTAIL.t8 2.11588
R473 VTAIL.n56 VTAIL.t2 2.11588
R474 VTAIL.n197 VTAIL.n195 1.93989
R475 VTAIL.n210 VTAIL.n209 1.93989
R476 VTAIL.n35 VTAIL.n33 1.93989
R477 VTAIL.n48 VTAIL.n47 1.93989
R478 VTAIL.n160 VTAIL.n159 1.93989
R479 VTAIL.n148 VTAIL.n147 1.93989
R480 VTAIL.n106 VTAIL.n105 1.93989
R481 VTAIL.n94 VTAIL.n93 1.93989
R482 VTAIL.n196 VTAIL.n170 1.16414
R483 VTAIL.n206 VTAIL.n166 1.16414
R484 VTAIL.n34 VTAIL.n8 1.16414
R485 VTAIL.n44 VTAIL.n4 1.16414
R486 VTAIL.n156 VTAIL.n116 1.16414
R487 VTAIL.n151 VTAIL.n121 1.16414
R488 VTAIL.n102 VTAIL.n62 1.16414
R489 VTAIL.n97 VTAIL.n67 1.16414
R490 VTAIL VTAIL.n215 0.834552
R491 VTAIL.n202 VTAIL.n201 0.388379
R492 VTAIL.n205 VTAIL.n168 0.388379
R493 VTAIL.n40 VTAIL.n39 0.388379
R494 VTAIL.n43 VTAIL.n6 0.388379
R495 VTAIL.n155 VTAIL.n118 0.388379
R496 VTAIL.n152 VTAIL.n120 0.388379
R497 VTAIL.n101 VTAIL.n64 0.388379
R498 VTAIL.n98 VTAIL.n66 0.388379
R499 VTAIL.n185 VTAIL.n177 0.155672
R500 VTAIL.n186 VTAIL.n185 0.155672
R501 VTAIL.n186 VTAIL.n173 0.155672
R502 VTAIL.n193 VTAIL.n173 0.155672
R503 VTAIL.n194 VTAIL.n193 0.155672
R504 VTAIL.n194 VTAIL.n169 0.155672
R505 VTAIL.n203 VTAIL.n169 0.155672
R506 VTAIL.n204 VTAIL.n203 0.155672
R507 VTAIL.n204 VTAIL.n165 0.155672
R508 VTAIL.n211 VTAIL.n165 0.155672
R509 VTAIL.n23 VTAIL.n15 0.155672
R510 VTAIL.n24 VTAIL.n23 0.155672
R511 VTAIL.n24 VTAIL.n11 0.155672
R512 VTAIL.n31 VTAIL.n11 0.155672
R513 VTAIL.n32 VTAIL.n31 0.155672
R514 VTAIL.n32 VTAIL.n7 0.155672
R515 VTAIL.n41 VTAIL.n7 0.155672
R516 VTAIL.n42 VTAIL.n41 0.155672
R517 VTAIL.n42 VTAIL.n3 0.155672
R518 VTAIL.n49 VTAIL.n3 0.155672
R519 VTAIL.n161 VTAIL.n115 0.155672
R520 VTAIL.n154 VTAIL.n115 0.155672
R521 VTAIL.n154 VTAIL.n153 0.155672
R522 VTAIL.n153 VTAIL.n119 0.155672
R523 VTAIL.n146 VTAIL.n119 0.155672
R524 VTAIL.n146 VTAIL.n145 0.155672
R525 VTAIL.n145 VTAIL.n125 0.155672
R526 VTAIL.n138 VTAIL.n125 0.155672
R527 VTAIL.n138 VTAIL.n137 0.155672
R528 VTAIL.n137 VTAIL.n129 0.155672
R529 VTAIL.n107 VTAIL.n61 0.155672
R530 VTAIL.n100 VTAIL.n61 0.155672
R531 VTAIL.n100 VTAIL.n99 0.155672
R532 VTAIL.n99 VTAIL.n65 0.155672
R533 VTAIL.n92 VTAIL.n65 0.155672
R534 VTAIL.n92 VTAIL.n91 0.155672
R535 VTAIL.n91 VTAIL.n71 0.155672
R536 VTAIL.n84 VTAIL.n71 0.155672
R537 VTAIL.n84 VTAIL.n83 0.155672
R538 VTAIL.n83 VTAIL.n75 0.155672
R539 VDD1.n44 VDD1.n0 289.615
R540 VDD1.n95 VDD1.n51 289.615
R541 VDD1.n45 VDD1.n44 185
R542 VDD1.n43 VDD1.n42 185
R543 VDD1.n4 VDD1.n3 185
R544 VDD1.n8 VDD1.n6 185
R545 VDD1.n37 VDD1.n36 185
R546 VDD1.n35 VDD1.n34 185
R547 VDD1.n10 VDD1.n9 185
R548 VDD1.n29 VDD1.n28 185
R549 VDD1.n27 VDD1.n26 185
R550 VDD1.n14 VDD1.n13 185
R551 VDD1.n21 VDD1.n20 185
R552 VDD1.n19 VDD1.n18 185
R553 VDD1.n68 VDD1.n67 185
R554 VDD1.n70 VDD1.n69 185
R555 VDD1.n63 VDD1.n62 185
R556 VDD1.n76 VDD1.n75 185
R557 VDD1.n78 VDD1.n77 185
R558 VDD1.n59 VDD1.n58 185
R559 VDD1.n85 VDD1.n84 185
R560 VDD1.n86 VDD1.n57 185
R561 VDD1.n88 VDD1.n87 185
R562 VDD1.n55 VDD1.n54 185
R563 VDD1.n94 VDD1.n93 185
R564 VDD1.n96 VDD1.n95 185
R565 VDD1.n17 VDD1.t4 149.524
R566 VDD1.n66 VDD1.t2 149.524
R567 VDD1.n44 VDD1.n43 104.615
R568 VDD1.n43 VDD1.n3 104.615
R569 VDD1.n8 VDD1.n3 104.615
R570 VDD1.n36 VDD1.n8 104.615
R571 VDD1.n36 VDD1.n35 104.615
R572 VDD1.n35 VDD1.n9 104.615
R573 VDD1.n28 VDD1.n9 104.615
R574 VDD1.n28 VDD1.n27 104.615
R575 VDD1.n27 VDD1.n13 104.615
R576 VDD1.n20 VDD1.n13 104.615
R577 VDD1.n20 VDD1.n19 104.615
R578 VDD1.n69 VDD1.n68 104.615
R579 VDD1.n69 VDD1.n62 104.615
R580 VDD1.n76 VDD1.n62 104.615
R581 VDD1.n77 VDD1.n76 104.615
R582 VDD1.n77 VDD1.n58 104.615
R583 VDD1.n85 VDD1.n58 104.615
R584 VDD1.n86 VDD1.n85 104.615
R585 VDD1.n87 VDD1.n86 104.615
R586 VDD1.n87 VDD1.n54 104.615
R587 VDD1.n94 VDD1.n54 104.615
R588 VDD1.n95 VDD1.n94 104.615
R589 VDD1.n103 VDD1.n102 67.9505
R590 VDD1.n50 VDD1.n49 65.3293
R591 VDD1.n105 VDD1.n104 65.3292
R592 VDD1.n101 VDD1.n100 65.3292
R593 VDD1.n50 VDD1.n48 54.7604
R594 VDD1.n101 VDD1.n99 54.7604
R595 VDD1.n19 VDD1.t4 52.3082
R596 VDD1.n68 VDD1.t2 52.3082
R597 VDD1.n105 VDD1.n103 51.1043
R598 VDD1.n6 VDD1.n4 13.1884
R599 VDD1.n88 VDD1.n55 13.1884
R600 VDD1.n42 VDD1.n41 12.8005
R601 VDD1.n38 VDD1.n37 12.8005
R602 VDD1.n89 VDD1.n57 12.8005
R603 VDD1.n93 VDD1.n92 12.8005
R604 VDD1.n45 VDD1.n2 12.0247
R605 VDD1.n34 VDD1.n7 12.0247
R606 VDD1.n84 VDD1.n83 12.0247
R607 VDD1.n96 VDD1.n53 12.0247
R608 VDD1.n46 VDD1.n0 11.249
R609 VDD1.n33 VDD1.n10 11.249
R610 VDD1.n82 VDD1.n59 11.249
R611 VDD1.n97 VDD1.n51 11.249
R612 VDD1.n30 VDD1.n29 10.4732
R613 VDD1.n79 VDD1.n78 10.4732
R614 VDD1.n18 VDD1.n17 10.2747
R615 VDD1.n67 VDD1.n66 10.2747
R616 VDD1.n26 VDD1.n12 9.69747
R617 VDD1.n75 VDD1.n61 9.69747
R618 VDD1.n48 VDD1.n47 9.45567
R619 VDD1.n99 VDD1.n98 9.45567
R620 VDD1.n16 VDD1.n15 9.3005
R621 VDD1.n23 VDD1.n22 9.3005
R622 VDD1.n25 VDD1.n24 9.3005
R623 VDD1.n12 VDD1.n11 9.3005
R624 VDD1.n31 VDD1.n30 9.3005
R625 VDD1.n33 VDD1.n32 9.3005
R626 VDD1.n7 VDD1.n5 9.3005
R627 VDD1.n39 VDD1.n38 9.3005
R628 VDD1.n47 VDD1.n46 9.3005
R629 VDD1.n2 VDD1.n1 9.3005
R630 VDD1.n41 VDD1.n40 9.3005
R631 VDD1.n98 VDD1.n97 9.3005
R632 VDD1.n53 VDD1.n52 9.3005
R633 VDD1.n92 VDD1.n91 9.3005
R634 VDD1.n65 VDD1.n64 9.3005
R635 VDD1.n72 VDD1.n71 9.3005
R636 VDD1.n74 VDD1.n73 9.3005
R637 VDD1.n61 VDD1.n60 9.3005
R638 VDD1.n80 VDD1.n79 9.3005
R639 VDD1.n82 VDD1.n81 9.3005
R640 VDD1.n83 VDD1.n56 9.3005
R641 VDD1.n90 VDD1.n89 9.3005
R642 VDD1.n25 VDD1.n14 8.92171
R643 VDD1.n74 VDD1.n63 8.92171
R644 VDD1.n22 VDD1.n21 8.14595
R645 VDD1.n71 VDD1.n70 8.14595
R646 VDD1.n18 VDD1.n16 7.3702
R647 VDD1.n67 VDD1.n65 7.3702
R648 VDD1.n21 VDD1.n16 5.81868
R649 VDD1.n70 VDD1.n65 5.81868
R650 VDD1.n22 VDD1.n14 5.04292
R651 VDD1.n71 VDD1.n63 5.04292
R652 VDD1.n26 VDD1.n25 4.26717
R653 VDD1.n75 VDD1.n74 4.26717
R654 VDD1.n29 VDD1.n12 3.49141
R655 VDD1.n78 VDD1.n61 3.49141
R656 VDD1.n17 VDD1.n15 2.84303
R657 VDD1.n66 VDD1.n64 2.84303
R658 VDD1.n48 VDD1.n0 2.71565
R659 VDD1.n30 VDD1.n10 2.71565
R660 VDD1.n79 VDD1.n59 2.71565
R661 VDD1.n99 VDD1.n51 2.71565
R662 VDD1 VDD1.n105 2.61903
R663 VDD1.n104 VDD1.t5 2.11588
R664 VDD1.n104 VDD1.t1 2.11588
R665 VDD1.n49 VDD1.t0 2.11588
R666 VDD1.n49 VDD1.t7 2.11588
R667 VDD1.n102 VDD1.t8 2.11588
R668 VDD1.n102 VDD1.t9 2.11588
R669 VDD1.n100 VDD1.t3 2.11588
R670 VDD1.n100 VDD1.t6 2.11588
R671 VDD1.n46 VDD1.n45 1.93989
R672 VDD1.n34 VDD1.n33 1.93989
R673 VDD1.n84 VDD1.n82 1.93989
R674 VDD1.n97 VDD1.n96 1.93989
R675 VDD1.n42 VDD1.n2 1.16414
R676 VDD1.n37 VDD1.n7 1.16414
R677 VDD1.n83 VDD1.n57 1.16414
R678 VDD1.n93 VDD1.n53 1.16414
R679 VDD1 VDD1.n50 0.950931
R680 VDD1.n103 VDD1.n101 0.837395
R681 VDD1.n41 VDD1.n4 0.388379
R682 VDD1.n38 VDD1.n6 0.388379
R683 VDD1.n89 VDD1.n88 0.388379
R684 VDD1.n92 VDD1.n55 0.388379
R685 VDD1.n47 VDD1.n1 0.155672
R686 VDD1.n40 VDD1.n1 0.155672
R687 VDD1.n40 VDD1.n39 0.155672
R688 VDD1.n39 VDD1.n5 0.155672
R689 VDD1.n32 VDD1.n5 0.155672
R690 VDD1.n32 VDD1.n31 0.155672
R691 VDD1.n31 VDD1.n11 0.155672
R692 VDD1.n24 VDD1.n11 0.155672
R693 VDD1.n24 VDD1.n23 0.155672
R694 VDD1.n23 VDD1.n15 0.155672
R695 VDD1.n72 VDD1.n64 0.155672
R696 VDD1.n73 VDD1.n72 0.155672
R697 VDD1.n73 VDD1.n60 0.155672
R698 VDD1.n80 VDD1.n60 0.155672
R699 VDD1.n81 VDD1.n80 0.155672
R700 VDD1.n81 VDD1.n56 0.155672
R701 VDD1.n90 VDD1.n56 0.155672
R702 VDD1.n91 VDD1.n90 0.155672
R703 VDD1.n91 VDD1.n52 0.155672
R704 VDD1.n98 VDD1.n52 0.155672
R705 B.n1047 B.n1046 585
R706 B.n1048 B.n1047 585
R707 B.n342 B.n185 585
R708 B.n341 B.n340 585
R709 B.n339 B.n338 585
R710 B.n337 B.n336 585
R711 B.n335 B.n334 585
R712 B.n333 B.n332 585
R713 B.n331 B.n330 585
R714 B.n329 B.n328 585
R715 B.n327 B.n326 585
R716 B.n325 B.n324 585
R717 B.n323 B.n322 585
R718 B.n321 B.n320 585
R719 B.n319 B.n318 585
R720 B.n317 B.n316 585
R721 B.n315 B.n314 585
R722 B.n313 B.n312 585
R723 B.n311 B.n310 585
R724 B.n309 B.n308 585
R725 B.n307 B.n306 585
R726 B.n305 B.n304 585
R727 B.n303 B.n302 585
R728 B.n301 B.n300 585
R729 B.n299 B.n298 585
R730 B.n297 B.n296 585
R731 B.n295 B.n294 585
R732 B.n293 B.n292 585
R733 B.n291 B.n290 585
R734 B.n289 B.n288 585
R735 B.n287 B.n286 585
R736 B.n285 B.n284 585
R737 B.n283 B.n282 585
R738 B.n281 B.n280 585
R739 B.n279 B.n278 585
R740 B.n276 B.n275 585
R741 B.n274 B.n273 585
R742 B.n272 B.n271 585
R743 B.n270 B.n269 585
R744 B.n268 B.n267 585
R745 B.n266 B.n265 585
R746 B.n264 B.n263 585
R747 B.n262 B.n261 585
R748 B.n260 B.n259 585
R749 B.n258 B.n257 585
R750 B.n256 B.n255 585
R751 B.n254 B.n253 585
R752 B.n252 B.n251 585
R753 B.n250 B.n249 585
R754 B.n248 B.n247 585
R755 B.n246 B.n245 585
R756 B.n244 B.n243 585
R757 B.n242 B.n241 585
R758 B.n240 B.n239 585
R759 B.n238 B.n237 585
R760 B.n236 B.n235 585
R761 B.n234 B.n233 585
R762 B.n232 B.n231 585
R763 B.n230 B.n229 585
R764 B.n228 B.n227 585
R765 B.n226 B.n225 585
R766 B.n224 B.n223 585
R767 B.n222 B.n221 585
R768 B.n220 B.n219 585
R769 B.n218 B.n217 585
R770 B.n216 B.n215 585
R771 B.n214 B.n213 585
R772 B.n212 B.n211 585
R773 B.n210 B.n209 585
R774 B.n208 B.n207 585
R775 B.n206 B.n205 585
R776 B.n204 B.n203 585
R777 B.n202 B.n201 585
R778 B.n200 B.n199 585
R779 B.n198 B.n197 585
R780 B.n196 B.n195 585
R781 B.n194 B.n193 585
R782 B.n192 B.n191 585
R783 B.n1045 B.n146 585
R784 B.n1049 B.n146 585
R785 B.n1044 B.n145 585
R786 B.n1050 B.n145 585
R787 B.n1043 B.n1042 585
R788 B.n1042 B.n141 585
R789 B.n1041 B.n140 585
R790 B.n1056 B.n140 585
R791 B.n1040 B.n139 585
R792 B.n1057 B.n139 585
R793 B.n1039 B.n138 585
R794 B.n1058 B.n138 585
R795 B.n1038 B.n1037 585
R796 B.n1037 B.n134 585
R797 B.n1036 B.n133 585
R798 B.n1064 B.n133 585
R799 B.n1035 B.n132 585
R800 B.n1065 B.n132 585
R801 B.n1034 B.n131 585
R802 B.n1066 B.n131 585
R803 B.n1033 B.n1032 585
R804 B.n1032 B.n127 585
R805 B.n1031 B.n126 585
R806 B.n1072 B.n126 585
R807 B.n1030 B.n125 585
R808 B.n1073 B.n125 585
R809 B.n1029 B.n124 585
R810 B.n1074 B.n124 585
R811 B.n1028 B.n1027 585
R812 B.n1027 B.n120 585
R813 B.n1026 B.n119 585
R814 B.n1080 B.n119 585
R815 B.n1025 B.n118 585
R816 B.n1081 B.n118 585
R817 B.n1024 B.n117 585
R818 B.n1082 B.n117 585
R819 B.n1023 B.n1022 585
R820 B.n1022 B.n113 585
R821 B.n1021 B.n112 585
R822 B.n1088 B.n112 585
R823 B.n1020 B.n111 585
R824 B.n1089 B.n111 585
R825 B.n1019 B.n110 585
R826 B.n1090 B.n110 585
R827 B.n1018 B.n1017 585
R828 B.n1017 B.n106 585
R829 B.n1016 B.n105 585
R830 B.n1096 B.n105 585
R831 B.n1015 B.n104 585
R832 B.n1097 B.n104 585
R833 B.n1014 B.n103 585
R834 B.n1098 B.n103 585
R835 B.n1013 B.n1012 585
R836 B.n1012 B.n99 585
R837 B.n1011 B.n98 585
R838 B.n1104 B.n98 585
R839 B.n1010 B.n97 585
R840 B.n1105 B.n97 585
R841 B.n1009 B.n96 585
R842 B.n1106 B.n96 585
R843 B.n1008 B.n1007 585
R844 B.n1007 B.n92 585
R845 B.n1006 B.n91 585
R846 B.n1112 B.n91 585
R847 B.n1005 B.n90 585
R848 B.n1113 B.n90 585
R849 B.n1004 B.n89 585
R850 B.n1114 B.n89 585
R851 B.n1003 B.n1002 585
R852 B.n1002 B.n85 585
R853 B.n1001 B.n84 585
R854 B.n1120 B.n84 585
R855 B.n1000 B.n83 585
R856 B.n1121 B.n83 585
R857 B.n999 B.n82 585
R858 B.n1122 B.n82 585
R859 B.n998 B.n997 585
R860 B.n997 B.n78 585
R861 B.n996 B.n77 585
R862 B.n1128 B.n77 585
R863 B.n995 B.n76 585
R864 B.n1129 B.n76 585
R865 B.n994 B.n75 585
R866 B.n1130 B.n75 585
R867 B.n993 B.n992 585
R868 B.n992 B.n71 585
R869 B.n991 B.n70 585
R870 B.n1136 B.n70 585
R871 B.n990 B.n69 585
R872 B.n1137 B.n69 585
R873 B.n989 B.n68 585
R874 B.n1138 B.n68 585
R875 B.n988 B.n987 585
R876 B.n987 B.n64 585
R877 B.n986 B.n63 585
R878 B.n1144 B.n63 585
R879 B.n985 B.n62 585
R880 B.n1145 B.n62 585
R881 B.n984 B.n61 585
R882 B.n1146 B.n61 585
R883 B.n983 B.n982 585
R884 B.n982 B.n57 585
R885 B.n981 B.n56 585
R886 B.n1152 B.n56 585
R887 B.n980 B.n55 585
R888 B.n1153 B.n55 585
R889 B.n979 B.n54 585
R890 B.n1154 B.n54 585
R891 B.n978 B.n977 585
R892 B.n977 B.n50 585
R893 B.n976 B.n49 585
R894 B.n1160 B.n49 585
R895 B.n975 B.n48 585
R896 B.n1161 B.n48 585
R897 B.n974 B.n47 585
R898 B.n1162 B.n47 585
R899 B.n973 B.n972 585
R900 B.n972 B.n43 585
R901 B.n971 B.n42 585
R902 B.n1168 B.n42 585
R903 B.n970 B.n41 585
R904 B.n1169 B.n41 585
R905 B.n969 B.n40 585
R906 B.n1170 B.n40 585
R907 B.n968 B.n967 585
R908 B.n967 B.n36 585
R909 B.n966 B.n35 585
R910 B.n1176 B.n35 585
R911 B.n965 B.n34 585
R912 B.n1177 B.n34 585
R913 B.n964 B.n33 585
R914 B.n1178 B.n33 585
R915 B.n963 B.n962 585
R916 B.n962 B.n29 585
R917 B.n961 B.n28 585
R918 B.n1184 B.n28 585
R919 B.n960 B.n27 585
R920 B.n1185 B.n27 585
R921 B.n959 B.n26 585
R922 B.n1186 B.n26 585
R923 B.n958 B.n957 585
R924 B.n957 B.n22 585
R925 B.n956 B.n21 585
R926 B.n1192 B.n21 585
R927 B.n955 B.n20 585
R928 B.n1193 B.n20 585
R929 B.n954 B.n19 585
R930 B.n1194 B.n19 585
R931 B.n953 B.n952 585
R932 B.n952 B.n15 585
R933 B.n951 B.n14 585
R934 B.n1200 B.n14 585
R935 B.n950 B.n13 585
R936 B.n1201 B.n13 585
R937 B.n949 B.n12 585
R938 B.n1202 B.n12 585
R939 B.n948 B.n947 585
R940 B.n947 B.n8 585
R941 B.n946 B.n7 585
R942 B.n1208 B.n7 585
R943 B.n945 B.n6 585
R944 B.n1209 B.n6 585
R945 B.n944 B.n5 585
R946 B.n1210 B.n5 585
R947 B.n943 B.n942 585
R948 B.n942 B.n4 585
R949 B.n941 B.n343 585
R950 B.n941 B.n940 585
R951 B.n931 B.n344 585
R952 B.n345 B.n344 585
R953 B.n933 B.n932 585
R954 B.n934 B.n933 585
R955 B.n930 B.n350 585
R956 B.n350 B.n349 585
R957 B.n929 B.n928 585
R958 B.n928 B.n927 585
R959 B.n352 B.n351 585
R960 B.n353 B.n352 585
R961 B.n920 B.n919 585
R962 B.n921 B.n920 585
R963 B.n918 B.n358 585
R964 B.n358 B.n357 585
R965 B.n917 B.n916 585
R966 B.n916 B.n915 585
R967 B.n360 B.n359 585
R968 B.n361 B.n360 585
R969 B.n908 B.n907 585
R970 B.n909 B.n908 585
R971 B.n906 B.n366 585
R972 B.n366 B.n365 585
R973 B.n905 B.n904 585
R974 B.n904 B.n903 585
R975 B.n368 B.n367 585
R976 B.n369 B.n368 585
R977 B.n896 B.n895 585
R978 B.n897 B.n896 585
R979 B.n894 B.n374 585
R980 B.n374 B.n373 585
R981 B.n893 B.n892 585
R982 B.n892 B.n891 585
R983 B.n376 B.n375 585
R984 B.n377 B.n376 585
R985 B.n884 B.n883 585
R986 B.n885 B.n884 585
R987 B.n882 B.n382 585
R988 B.n382 B.n381 585
R989 B.n881 B.n880 585
R990 B.n880 B.n879 585
R991 B.n384 B.n383 585
R992 B.n385 B.n384 585
R993 B.n872 B.n871 585
R994 B.n873 B.n872 585
R995 B.n870 B.n390 585
R996 B.n390 B.n389 585
R997 B.n869 B.n868 585
R998 B.n868 B.n867 585
R999 B.n392 B.n391 585
R1000 B.n393 B.n392 585
R1001 B.n860 B.n859 585
R1002 B.n861 B.n860 585
R1003 B.n858 B.n398 585
R1004 B.n398 B.n397 585
R1005 B.n857 B.n856 585
R1006 B.n856 B.n855 585
R1007 B.n400 B.n399 585
R1008 B.n401 B.n400 585
R1009 B.n848 B.n847 585
R1010 B.n849 B.n848 585
R1011 B.n846 B.n405 585
R1012 B.n409 B.n405 585
R1013 B.n845 B.n844 585
R1014 B.n844 B.n843 585
R1015 B.n407 B.n406 585
R1016 B.n408 B.n407 585
R1017 B.n836 B.n835 585
R1018 B.n837 B.n836 585
R1019 B.n834 B.n414 585
R1020 B.n414 B.n413 585
R1021 B.n833 B.n832 585
R1022 B.n832 B.n831 585
R1023 B.n416 B.n415 585
R1024 B.n417 B.n416 585
R1025 B.n824 B.n823 585
R1026 B.n825 B.n824 585
R1027 B.n822 B.n422 585
R1028 B.n422 B.n421 585
R1029 B.n821 B.n820 585
R1030 B.n820 B.n819 585
R1031 B.n424 B.n423 585
R1032 B.n425 B.n424 585
R1033 B.n812 B.n811 585
R1034 B.n813 B.n812 585
R1035 B.n810 B.n429 585
R1036 B.n433 B.n429 585
R1037 B.n809 B.n808 585
R1038 B.n808 B.n807 585
R1039 B.n431 B.n430 585
R1040 B.n432 B.n431 585
R1041 B.n800 B.n799 585
R1042 B.n801 B.n800 585
R1043 B.n798 B.n438 585
R1044 B.n438 B.n437 585
R1045 B.n797 B.n796 585
R1046 B.n796 B.n795 585
R1047 B.n440 B.n439 585
R1048 B.n441 B.n440 585
R1049 B.n788 B.n787 585
R1050 B.n789 B.n788 585
R1051 B.n786 B.n446 585
R1052 B.n446 B.n445 585
R1053 B.n785 B.n784 585
R1054 B.n784 B.n783 585
R1055 B.n448 B.n447 585
R1056 B.n449 B.n448 585
R1057 B.n776 B.n775 585
R1058 B.n777 B.n776 585
R1059 B.n774 B.n453 585
R1060 B.n457 B.n453 585
R1061 B.n773 B.n772 585
R1062 B.n772 B.n771 585
R1063 B.n455 B.n454 585
R1064 B.n456 B.n455 585
R1065 B.n764 B.n763 585
R1066 B.n765 B.n764 585
R1067 B.n762 B.n462 585
R1068 B.n462 B.n461 585
R1069 B.n761 B.n760 585
R1070 B.n760 B.n759 585
R1071 B.n464 B.n463 585
R1072 B.n465 B.n464 585
R1073 B.n752 B.n751 585
R1074 B.n753 B.n752 585
R1075 B.n750 B.n470 585
R1076 B.n470 B.n469 585
R1077 B.n749 B.n748 585
R1078 B.n748 B.n747 585
R1079 B.n472 B.n471 585
R1080 B.n473 B.n472 585
R1081 B.n740 B.n739 585
R1082 B.n741 B.n740 585
R1083 B.n738 B.n478 585
R1084 B.n478 B.n477 585
R1085 B.n737 B.n736 585
R1086 B.n736 B.n735 585
R1087 B.n480 B.n479 585
R1088 B.n481 B.n480 585
R1089 B.n728 B.n727 585
R1090 B.n729 B.n728 585
R1091 B.n726 B.n486 585
R1092 B.n486 B.n485 585
R1093 B.n725 B.n724 585
R1094 B.n724 B.n723 585
R1095 B.n488 B.n487 585
R1096 B.n489 B.n488 585
R1097 B.n716 B.n715 585
R1098 B.n717 B.n716 585
R1099 B.n714 B.n494 585
R1100 B.n494 B.n493 585
R1101 B.n713 B.n712 585
R1102 B.n712 B.n711 585
R1103 B.n496 B.n495 585
R1104 B.n497 B.n496 585
R1105 B.n704 B.n703 585
R1106 B.n705 B.n704 585
R1107 B.n702 B.n502 585
R1108 B.n502 B.n501 585
R1109 B.n696 B.n695 585
R1110 B.n694 B.n542 585
R1111 B.n693 B.n541 585
R1112 B.n698 B.n541 585
R1113 B.n692 B.n691 585
R1114 B.n690 B.n689 585
R1115 B.n688 B.n687 585
R1116 B.n686 B.n685 585
R1117 B.n684 B.n683 585
R1118 B.n682 B.n681 585
R1119 B.n680 B.n679 585
R1120 B.n678 B.n677 585
R1121 B.n676 B.n675 585
R1122 B.n674 B.n673 585
R1123 B.n672 B.n671 585
R1124 B.n670 B.n669 585
R1125 B.n668 B.n667 585
R1126 B.n666 B.n665 585
R1127 B.n664 B.n663 585
R1128 B.n662 B.n661 585
R1129 B.n660 B.n659 585
R1130 B.n658 B.n657 585
R1131 B.n656 B.n655 585
R1132 B.n654 B.n653 585
R1133 B.n652 B.n651 585
R1134 B.n650 B.n649 585
R1135 B.n648 B.n647 585
R1136 B.n646 B.n645 585
R1137 B.n644 B.n643 585
R1138 B.n642 B.n641 585
R1139 B.n640 B.n639 585
R1140 B.n638 B.n637 585
R1141 B.n636 B.n635 585
R1142 B.n634 B.n633 585
R1143 B.n632 B.n631 585
R1144 B.n629 B.n628 585
R1145 B.n627 B.n626 585
R1146 B.n625 B.n624 585
R1147 B.n623 B.n622 585
R1148 B.n621 B.n620 585
R1149 B.n619 B.n618 585
R1150 B.n617 B.n616 585
R1151 B.n615 B.n614 585
R1152 B.n613 B.n612 585
R1153 B.n611 B.n610 585
R1154 B.n609 B.n608 585
R1155 B.n607 B.n606 585
R1156 B.n605 B.n604 585
R1157 B.n603 B.n602 585
R1158 B.n601 B.n600 585
R1159 B.n599 B.n598 585
R1160 B.n597 B.n596 585
R1161 B.n595 B.n594 585
R1162 B.n593 B.n592 585
R1163 B.n591 B.n590 585
R1164 B.n589 B.n588 585
R1165 B.n587 B.n586 585
R1166 B.n585 B.n584 585
R1167 B.n583 B.n582 585
R1168 B.n581 B.n580 585
R1169 B.n579 B.n578 585
R1170 B.n577 B.n576 585
R1171 B.n575 B.n574 585
R1172 B.n573 B.n572 585
R1173 B.n571 B.n570 585
R1174 B.n569 B.n568 585
R1175 B.n567 B.n566 585
R1176 B.n565 B.n564 585
R1177 B.n563 B.n562 585
R1178 B.n561 B.n560 585
R1179 B.n559 B.n558 585
R1180 B.n557 B.n556 585
R1181 B.n555 B.n554 585
R1182 B.n553 B.n552 585
R1183 B.n551 B.n550 585
R1184 B.n549 B.n548 585
R1185 B.n504 B.n503 585
R1186 B.n701 B.n700 585
R1187 B.n500 B.n499 585
R1188 B.n501 B.n500 585
R1189 B.n707 B.n706 585
R1190 B.n706 B.n705 585
R1191 B.n708 B.n498 585
R1192 B.n498 B.n497 585
R1193 B.n710 B.n709 585
R1194 B.n711 B.n710 585
R1195 B.n492 B.n491 585
R1196 B.n493 B.n492 585
R1197 B.n719 B.n718 585
R1198 B.n718 B.n717 585
R1199 B.n720 B.n490 585
R1200 B.n490 B.n489 585
R1201 B.n722 B.n721 585
R1202 B.n723 B.n722 585
R1203 B.n484 B.n483 585
R1204 B.n485 B.n484 585
R1205 B.n731 B.n730 585
R1206 B.n730 B.n729 585
R1207 B.n732 B.n482 585
R1208 B.n482 B.n481 585
R1209 B.n734 B.n733 585
R1210 B.n735 B.n734 585
R1211 B.n476 B.n475 585
R1212 B.n477 B.n476 585
R1213 B.n743 B.n742 585
R1214 B.n742 B.n741 585
R1215 B.n744 B.n474 585
R1216 B.n474 B.n473 585
R1217 B.n746 B.n745 585
R1218 B.n747 B.n746 585
R1219 B.n468 B.n467 585
R1220 B.n469 B.n468 585
R1221 B.n755 B.n754 585
R1222 B.n754 B.n753 585
R1223 B.n756 B.n466 585
R1224 B.n466 B.n465 585
R1225 B.n758 B.n757 585
R1226 B.n759 B.n758 585
R1227 B.n460 B.n459 585
R1228 B.n461 B.n460 585
R1229 B.n767 B.n766 585
R1230 B.n766 B.n765 585
R1231 B.n768 B.n458 585
R1232 B.n458 B.n456 585
R1233 B.n770 B.n769 585
R1234 B.n771 B.n770 585
R1235 B.n452 B.n451 585
R1236 B.n457 B.n452 585
R1237 B.n779 B.n778 585
R1238 B.n778 B.n777 585
R1239 B.n780 B.n450 585
R1240 B.n450 B.n449 585
R1241 B.n782 B.n781 585
R1242 B.n783 B.n782 585
R1243 B.n444 B.n443 585
R1244 B.n445 B.n444 585
R1245 B.n791 B.n790 585
R1246 B.n790 B.n789 585
R1247 B.n792 B.n442 585
R1248 B.n442 B.n441 585
R1249 B.n794 B.n793 585
R1250 B.n795 B.n794 585
R1251 B.n436 B.n435 585
R1252 B.n437 B.n436 585
R1253 B.n803 B.n802 585
R1254 B.n802 B.n801 585
R1255 B.n804 B.n434 585
R1256 B.n434 B.n432 585
R1257 B.n806 B.n805 585
R1258 B.n807 B.n806 585
R1259 B.n428 B.n427 585
R1260 B.n433 B.n428 585
R1261 B.n815 B.n814 585
R1262 B.n814 B.n813 585
R1263 B.n816 B.n426 585
R1264 B.n426 B.n425 585
R1265 B.n818 B.n817 585
R1266 B.n819 B.n818 585
R1267 B.n420 B.n419 585
R1268 B.n421 B.n420 585
R1269 B.n827 B.n826 585
R1270 B.n826 B.n825 585
R1271 B.n828 B.n418 585
R1272 B.n418 B.n417 585
R1273 B.n830 B.n829 585
R1274 B.n831 B.n830 585
R1275 B.n412 B.n411 585
R1276 B.n413 B.n412 585
R1277 B.n839 B.n838 585
R1278 B.n838 B.n837 585
R1279 B.n840 B.n410 585
R1280 B.n410 B.n408 585
R1281 B.n842 B.n841 585
R1282 B.n843 B.n842 585
R1283 B.n404 B.n403 585
R1284 B.n409 B.n404 585
R1285 B.n851 B.n850 585
R1286 B.n850 B.n849 585
R1287 B.n852 B.n402 585
R1288 B.n402 B.n401 585
R1289 B.n854 B.n853 585
R1290 B.n855 B.n854 585
R1291 B.n396 B.n395 585
R1292 B.n397 B.n396 585
R1293 B.n863 B.n862 585
R1294 B.n862 B.n861 585
R1295 B.n864 B.n394 585
R1296 B.n394 B.n393 585
R1297 B.n866 B.n865 585
R1298 B.n867 B.n866 585
R1299 B.n388 B.n387 585
R1300 B.n389 B.n388 585
R1301 B.n875 B.n874 585
R1302 B.n874 B.n873 585
R1303 B.n876 B.n386 585
R1304 B.n386 B.n385 585
R1305 B.n878 B.n877 585
R1306 B.n879 B.n878 585
R1307 B.n380 B.n379 585
R1308 B.n381 B.n380 585
R1309 B.n887 B.n886 585
R1310 B.n886 B.n885 585
R1311 B.n888 B.n378 585
R1312 B.n378 B.n377 585
R1313 B.n890 B.n889 585
R1314 B.n891 B.n890 585
R1315 B.n372 B.n371 585
R1316 B.n373 B.n372 585
R1317 B.n899 B.n898 585
R1318 B.n898 B.n897 585
R1319 B.n900 B.n370 585
R1320 B.n370 B.n369 585
R1321 B.n902 B.n901 585
R1322 B.n903 B.n902 585
R1323 B.n364 B.n363 585
R1324 B.n365 B.n364 585
R1325 B.n911 B.n910 585
R1326 B.n910 B.n909 585
R1327 B.n912 B.n362 585
R1328 B.n362 B.n361 585
R1329 B.n914 B.n913 585
R1330 B.n915 B.n914 585
R1331 B.n356 B.n355 585
R1332 B.n357 B.n356 585
R1333 B.n923 B.n922 585
R1334 B.n922 B.n921 585
R1335 B.n924 B.n354 585
R1336 B.n354 B.n353 585
R1337 B.n926 B.n925 585
R1338 B.n927 B.n926 585
R1339 B.n348 B.n347 585
R1340 B.n349 B.n348 585
R1341 B.n936 B.n935 585
R1342 B.n935 B.n934 585
R1343 B.n937 B.n346 585
R1344 B.n346 B.n345 585
R1345 B.n939 B.n938 585
R1346 B.n940 B.n939 585
R1347 B.n2 B.n0 585
R1348 B.n4 B.n2 585
R1349 B.n3 B.n1 585
R1350 B.n1209 B.n3 585
R1351 B.n1207 B.n1206 585
R1352 B.n1208 B.n1207 585
R1353 B.n1205 B.n9 585
R1354 B.n9 B.n8 585
R1355 B.n1204 B.n1203 585
R1356 B.n1203 B.n1202 585
R1357 B.n11 B.n10 585
R1358 B.n1201 B.n11 585
R1359 B.n1199 B.n1198 585
R1360 B.n1200 B.n1199 585
R1361 B.n1197 B.n16 585
R1362 B.n16 B.n15 585
R1363 B.n1196 B.n1195 585
R1364 B.n1195 B.n1194 585
R1365 B.n18 B.n17 585
R1366 B.n1193 B.n18 585
R1367 B.n1191 B.n1190 585
R1368 B.n1192 B.n1191 585
R1369 B.n1189 B.n23 585
R1370 B.n23 B.n22 585
R1371 B.n1188 B.n1187 585
R1372 B.n1187 B.n1186 585
R1373 B.n25 B.n24 585
R1374 B.n1185 B.n25 585
R1375 B.n1183 B.n1182 585
R1376 B.n1184 B.n1183 585
R1377 B.n1181 B.n30 585
R1378 B.n30 B.n29 585
R1379 B.n1180 B.n1179 585
R1380 B.n1179 B.n1178 585
R1381 B.n32 B.n31 585
R1382 B.n1177 B.n32 585
R1383 B.n1175 B.n1174 585
R1384 B.n1176 B.n1175 585
R1385 B.n1173 B.n37 585
R1386 B.n37 B.n36 585
R1387 B.n1172 B.n1171 585
R1388 B.n1171 B.n1170 585
R1389 B.n39 B.n38 585
R1390 B.n1169 B.n39 585
R1391 B.n1167 B.n1166 585
R1392 B.n1168 B.n1167 585
R1393 B.n1165 B.n44 585
R1394 B.n44 B.n43 585
R1395 B.n1164 B.n1163 585
R1396 B.n1163 B.n1162 585
R1397 B.n46 B.n45 585
R1398 B.n1161 B.n46 585
R1399 B.n1159 B.n1158 585
R1400 B.n1160 B.n1159 585
R1401 B.n1157 B.n51 585
R1402 B.n51 B.n50 585
R1403 B.n1156 B.n1155 585
R1404 B.n1155 B.n1154 585
R1405 B.n53 B.n52 585
R1406 B.n1153 B.n53 585
R1407 B.n1151 B.n1150 585
R1408 B.n1152 B.n1151 585
R1409 B.n1149 B.n58 585
R1410 B.n58 B.n57 585
R1411 B.n1148 B.n1147 585
R1412 B.n1147 B.n1146 585
R1413 B.n60 B.n59 585
R1414 B.n1145 B.n60 585
R1415 B.n1143 B.n1142 585
R1416 B.n1144 B.n1143 585
R1417 B.n1141 B.n65 585
R1418 B.n65 B.n64 585
R1419 B.n1140 B.n1139 585
R1420 B.n1139 B.n1138 585
R1421 B.n67 B.n66 585
R1422 B.n1137 B.n67 585
R1423 B.n1135 B.n1134 585
R1424 B.n1136 B.n1135 585
R1425 B.n1133 B.n72 585
R1426 B.n72 B.n71 585
R1427 B.n1132 B.n1131 585
R1428 B.n1131 B.n1130 585
R1429 B.n74 B.n73 585
R1430 B.n1129 B.n74 585
R1431 B.n1127 B.n1126 585
R1432 B.n1128 B.n1127 585
R1433 B.n1125 B.n79 585
R1434 B.n79 B.n78 585
R1435 B.n1124 B.n1123 585
R1436 B.n1123 B.n1122 585
R1437 B.n81 B.n80 585
R1438 B.n1121 B.n81 585
R1439 B.n1119 B.n1118 585
R1440 B.n1120 B.n1119 585
R1441 B.n1117 B.n86 585
R1442 B.n86 B.n85 585
R1443 B.n1116 B.n1115 585
R1444 B.n1115 B.n1114 585
R1445 B.n88 B.n87 585
R1446 B.n1113 B.n88 585
R1447 B.n1111 B.n1110 585
R1448 B.n1112 B.n1111 585
R1449 B.n1109 B.n93 585
R1450 B.n93 B.n92 585
R1451 B.n1108 B.n1107 585
R1452 B.n1107 B.n1106 585
R1453 B.n95 B.n94 585
R1454 B.n1105 B.n95 585
R1455 B.n1103 B.n1102 585
R1456 B.n1104 B.n1103 585
R1457 B.n1101 B.n100 585
R1458 B.n100 B.n99 585
R1459 B.n1100 B.n1099 585
R1460 B.n1099 B.n1098 585
R1461 B.n102 B.n101 585
R1462 B.n1097 B.n102 585
R1463 B.n1095 B.n1094 585
R1464 B.n1096 B.n1095 585
R1465 B.n1093 B.n107 585
R1466 B.n107 B.n106 585
R1467 B.n1092 B.n1091 585
R1468 B.n1091 B.n1090 585
R1469 B.n109 B.n108 585
R1470 B.n1089 B.n109 585
R1471 B.n1087 B.n1086 585
R1472 B.n1088 B.n1087 585
R1473 B.n1085 B.n114 585
R1474 B.n114 B.n113 585
R1475 B.n1084 B.n1083 585
R1476 B.n1083 B.n1082 585
R1477 B.n116 B.n115 585
R1478 B.n1081 B.n116 585
R1479 B.n1079 B.n1078 585
R1480 B.n1080 B.n1079 585
R1481 B.n1077 B.n121 585
R1482 B.n121 B.n120 585
R1483 B.n1076 B.n1075 585
R1484 B.n1075 B.n1074 585
R1485 B.n123 B.n122 585
R1486 B.n1073 B.n123 585
R1487 B.n1071 B.n1070 585
R1488 B.n1072 B.n1071 585
R1489 B.n1069 B.n128 585
R1490 B.n128 B.n127 585
R1491 B.n1068 B.n1067 585
R1492 B.n1067 B.n1066 585
R1493 B.n130 B.n129 585
R1494 B.n1065 B.n130 585
R1495 B.n1063 B.n1062 585
R1496 B.n1064 B.n1063 585
R1497 B.n1061 B.n135 585
R1498 B.n135 B.n134 585
R1499 B.n1060 B.n1059 585
R1500 B.n1059 B.n1058 585
R1501 B.n137 B.n136 585
R1502 B.n1057 B.n137 585
R1503 B.n1055 B.n1054 585
R1504 B.n1056 B.n1055 585
R1505 B.n1053 B.n142 585
R1506 B.n142 B.n141 585
R1507 B.n1052 B.n1051 585
R1508 B.n1051 B.n1050 585
R1509 B.n144 B.n143 585
R1510 B.n1049 B.n144 585
R1511 B.n1212 B.n1211 585
R1512 B.n1211 B.n1210 585
R1513 B.n696 B.n500 550.159
R1514 B.n191 B.n144 550.159
R1515 B.n700 B.n502 550.159
R1516 B.n1047 B.n146 550.159
R1517 B.n545 B.t23 317.002
R1518 B.n186 B.t12 317.002
R1519 B.n543 B.t20 317.002
R1520 B.n188 B.t15 317.002
R1521 B.n545 B.t21 268.558
R1522 B.n543 B.t17 268.558
R1523 B.n188 B.t14 268.558
R1524 B.n186 B.t10 268.558
R1525 B.n1048 B.n184 256.663
R1526 B.n1048 B.n183 256.663
R1527 B.n1048 B.n182 256.663
R1528 B.n1048 B.n181 256.663
R1529 B.n1048 B.n180 256.663
R1530 B.n1048 B.n179 256.663
R1531 B.n1048 B.n178 256.663
R1532 B.n1048 B.n177 256.663
R1533 B.n1048 B.n176 256.663
R1534 B.n1048 B.n175 256.663
R1535 B.n1048 B.n174 256.663
R1536 B.n1048 B.n173 256.663
R1537 B.n1048 B.n172 256.663
R1538 B.n1048 B.n171 256.663
R1539 B.n1048 B.n170 256.663
R1540 B.n1048 B.n169 256.663
R1541 B.n1048 B.n168 256.663
R1542 B.n1048 B.n167 256.663
R1543 B.n1048 B.n166 256.663
R1544 B.n1048 B.n165 256.663
R1545 B.n1048 B.n164 256.663
R1546 B.n1048 B.n163 256.663
R1547 B.n1048 B.n162 256.663
R1548 B.n1048 B.n161 256.663
R1549 B.n1048 B.n160 256.663
R1550 B.n1048 B.n159 256.663
R1551 B.n1048 B.n158 256.663
R1552 B.n1048 B.n157 256.663
R1553 B.n1048 B.n156 256.663
R1554 B.n1048 B.n155 256.663
R1555 B.n1048 B.n154 256.663
R1556 B.n1048 B.n153 256.663
R1557 B.n1048 B.n152 256.663
R1558 B.n1048 B.n151 256.663
R1559 B.n1048 B.n150 256.663
R1560 B.n1048 B.n149 256.663
R1561 B.n1048 B.n148 256.663
R1562 B.n1048 B.n147 256.663
R1563 B.n698 B.n697 256.663
R1564 B.n698 B.n505 256.663
R1565 B.n698 B.n506 256.663
R1566 B.n698 B.n507 256.663
R1567 B.n698 B.n508 256.663
R1568 B.n698 B.n509 256.663
R1569 B.n698 B.n510 256.663
R1570 B.n698 B.n511 256.663
R1571 B.n698 B.n512 256.663
R1572 B.n698 B.n513 256.663
R1573 B.n698 B.n514 256.663
R1574 B.n698 B.n515 256.663
R1575 B.n698 B.n516 256.663
R1576 B.n698 B.n517 256.663
R1577 B.n698 B.n518 256.663
R1578 B.n698 B.n519 256.663
R1579 B.n698 B.n520 256.663
R1580 B.n698 B.n521 256.663
R1581 B.n698 B.n522 256.663
R1582 B.n698 B.n523 256.663
R1583 B.n698 B.n524 256.663
R1584 B.n698 B.n525 256.663
R1585 B.n698 B.n526 256.663
R1586 B.n698 B.n527 256.663
R1587 B.n698 B.n528 256.663
R1588 B.n698 B.n529 256.663
R1589 B.n698 B.n530 256.663
R1590 B.n698 B.n531 256.663
R1591 B.n698 B.n532 256.663
R1592 B.n698 B.n533 256.663
R1593 B.n698 B.n534 256.663
R1594 B.n698 B.n535 256.663
R1595 B.n698 B.n536 256.663
R1596 B.n698 B.n537 256.663
R1597 B.n698 B.n538 256.663
R1598 B.n698 B.n539 256.663
R1599 B.n698 B.n540 256.663
R1600 B.n699 B.n698 256.663
R1601 B.n546 B.t22 236.712
R1602 B.n187 B.t13 236.712
R1603 B.n544 B.t19 236.712
R1604 B.n189 B.t16 236.712
R1605 B.n706 B.n500 163.367
R1606 B.n706 B.n498 163.367
R1607 B.n710 B.n498 163.367
R1608 B.n710 B.n492 163.367
R1609 B.n718 B.n492 163.367
R1610 B.n718 B.n490 163.367
R1611 B.n722 B.n490 163.367
R1612 B.n722 B.n484 163.367
R1613 B.n730 B.n484 163.367
R1614 B.n730 B.n482 163.367
R1615 B.n734 B.n482 163.367
R1616 B.n734 B.n476 163.367
R1617 B.n742 B.n476 163.367
R1618 B.n742 B.n474 163.367
R1619 B.n746 B.n474 163.367
R1620 B.n746 B.n468 163.367
R1621 B.n754 B.n468 163.367
R1622 B.n754 B.n466 163.367
R1623 B.n758 B.n466 163.367
R1624 B.n758 B.n460 163.367
R1625 B.n766 B.n460 163.367
R1626 B.n766 B.n458 163.367
R1627 B.n770 B.n458 163.367
R1628 B.n770 B.n452 163.367
R1629 B.n778 B.n452 163.367
R1630 B.n778 B.n450 163.367
R1631 B.n782 B.n450 163.367
R1632 B.n782 B.n444 163.367
R1633 B.n790 B.n444 163.367
R1634 B.n790 B.n442 163.367
R1635 B.n794 B.n442 163.367
R1636 B.n794 B.n436 163.367
R1637 B.n802 B.n436 163.367
R1638 B.n802 B.n434 163.367
R1639 B.n806 B.n434 163.367
R1640 B.n806 B.n428 163.367
R1641 B.n814 B.n428 163.367
R1642 B.n814 B.n426 163.367
R1643 B.n818 B.n426 163.367
R1644 B.n818 B.n420 163.367
R1645 B.n826 B.n420 163.367
R1646 B.n826 B.n418 163.367
R1647 B.n830 B.n418 163.367
R1648 B.n830 B.n412 163.367
R1649 B.n838 B.n412 163.367
R1650 B.n838 B.n410 163.367
R1651 B.n842 B.n410 163.367
R1652 B.n842 B.n404 163.367
R1653 B.n850 B.n404 163.367
R1654 B.n850 B.n402 163.367
R1655 B.n854 B.n402 163.367
R1656 B.n854 B.n396 163.367
R1657 B.n862 B.n396 163.367
R1658 B.n862 B.n394 163.367
R1659 B.n866 B.n394 163.367
R1660 B.n866 B.n388 163.367
R1661 B.n874 B.n388 163.367
R1662 B.n874 B.n386 163.367
R1663 B.n878 B.n386 163.367
R1664 B.n878 B.n380 163.367
R1665 B.n886 B.n380 163.367
R1666 B.n886 B.n378 163.367
R1667 B.n890 B.n378 163.367
R1668 B.n890 B.n372 163.367
R1669 B.n898 B.n372 163.367
R1670 B.n898 B.n370 163.367
R1671 B.n902 B.n370 163.367
R1672 B.n902 B.n364 163.367
R1673 B.n910 B.n364 163.367
R1674 B.n910 B.n362 163.367
R1675 B.n914 B.n362 163.367
R1676 B.n914 B.n356 163.367
R1677 B.n922 B.n356 163.367
R1678 B.n922 B.n354 163.367
R1679 B.n926 B.n354 163.367
R1680 B.n926 B.n348 163.367
R1681 B.n935 B.n348 163.367
R1682 B.n935 B.n346 163.367
R1683 B.n939 B.n346 163.367
R1684 B.n939 B.n2 163.367
R1685 B.n1211 B.n2 163.367
R1686 B.n1211 B.n3 163.367
R1687 B.n1207 B.n3 163.367
R1688 B.n1207 B.n9 163.367
R1689 B.n1203 B.n9 163.367
R1690 B.n1203 B.n11 163.367
R1691 B.n1199 B.n11 163.367
R1692 B.n1199 B.n16 163.367
R1693 B.n1195 B.n16 163.367
R1694 B.n1195 B.n18 163.367
R1695 B.n1191 B.n18 163.367
R1696 B.n1191 B.n23 163.367
R1697 B.n1187 B.n23 163.367
R1698 B.n1187 B.n25 163.367
R1699 B.n1183 B.n25 163.367
R1700 B.n1183 B.n30 163.367
R1701 B.n1179 B.n30 163.367
R1702 B.n1179 B.n32 163.367
R1703 B.n1175 B.n32 163.367
R1704 B.n1175 B.n37 163.367
R1705 B.n1171 B.n37 163.367
R1706 B.n1171 B.n39 163.367
R1707 B.n1167 B.n39 163.367
R1708 B.n1167 B.n44 163.367
R1709 B.n1163 B.n44 163.367
R1710 B.n1163 B.n46 163.367
R1711 B.n1159 B.n46 163.367
R1712 B.n1159 B.n51 163.367
R1713 B.n1155 B.n51 163.367
R1714 B.n1155 B.n53 163.367
R1715 B.n1151 B.n53 163.367
R1716 B.n1151 B.n58 163.367
R1717 B.n1147 B.n58 163.367
R1718 B.n1147 B.n60 163.367
R1719 B.n1143 B.n60 163.367
R1720 B.n1143 B.n65 163.367
R1721 B.n1139 B.n65 163.367
R1722 B.n1139 B.n67 163.367
R1723 B.n1135 B.n67 163.367
R1724 B.n1135 B.n72 163.367
R1725 B.n1131 B.n72 163.367
R1726 B.n1131 B.n74 163.367
R1727 B.n1127 B.n74 163.367
R1728 B.n1127 B.n79 163.367
R1729 B.n1123 B.n79 163.367
R1730 B.n1123 B.n81 163.367
R1731 B.n1119 B.n81 163.367
R1732 B.n1119 B.n86 163.367
R1733 B.n1115 B.n86 163.367
R1734 B.n1115 B.n88 163.367
R1735 B.n1111 B.n88 163.367
R1736 B.n1111 B.n93 163.367
R1737 B.n1107 B.n93 163.367
R1738 B.n1107 B.n95 163.367
R1739 B.n1103 B.n95 163.367
R1740 B.n1103 B.n100 163.367
R1741 B.n1099 B.n100 163.367
R1742 B.n1099 B.n102 163.367
R1743 B.n1095 B.n102 163.367
R1744 B.n1095 B.n107 163.367
R1745 B.n1091 B.n107 163.367
R1746 B.n1091 B.n109 163.367
R1747 B.n1087 B.n109 163.367
R1748 B.n1087 B.n114 163.367
R1749 B.n1083 B.n114 163.367
R1750 B.n1083 B.n116 163.367
R1751 B.n1079 B.n116 163.367
R1752 B.n1079 B.n121 163.367
R1753 B.n1075 B.n121 163.367
R1754 B.n1075 B.n123 163.367
R1755 B.n1071 B.n123 163.367
R1756 B.n1071 B.n128 163.367
R1757 B.n1067 B.n128 163.367
R1758 B.n1067 B.n130 163.367
R1759 B.n1063 B.n130 163.367
R1760 B.n1063 B.n135 163.367
R1761 B.n1059 B.n135 163.367
R1762 B.n1059 B.n137 163.367
R1763 B.n1055 B.n137 163.367
R1764 B.n1055 B.n142 163.367
R1765 B.n1051 B.n142 163.367
R1766 B.n1051 B.n144 163.367
R1767 B.n542 B.n541 163.367
R1768 B.n691 B.n541 163.367
R1769 B.n689 B.n688 163.367
R1770 B.n685 B.n684 163.367
R1771 B.n681 B.n680 163.367
R1772 B.n677 B.n676 163.367
R1773 B.n673 B.n672 163.367
R1774 B.n669 B.n668 163.367
R1775 B.n665 B.n664 163.367
R1776 B.n661 B.n660 163.367
R1777 B.n657 B.n656 163.367
R1778 B.n653 B.n652 163.367
R1779 B.n649 B.n648 163.367
R1780 B.n645 B.n644 163.367
R1781 B.n641 B.n640 163.367
R1782 B.n637 B.n636 163.367
R1783 B.n633 B.n632 163.367
R1784 B.n628 B.n627 163.367
R1785 B.n624 B.n623 163.367
R1786 B.n620 B.n619 163.367
R1787 B.n616 B.n615 163.367
R1788 B.n612 B.n611 163.367
R1789 B.n608 B.n607 163.367
R1790 B.n604 B.n603 163.367
R1791 B.n600 B.n599 163.367
R1792 B.n596 B.n595 163.367
R1793 B.n592 B.n591 163.367
R1794 B.n588 B.n587 163.367
R1795 B.n584 B.n583 163.367
R1796 B.n580 B.n579 163.367
R1797 B.n576 B.n575 163.367
R1798 B.n572 B.n571 163.367
R1799 B.n568 B.n567 163.367
R1800 B.n564 B.n563 163.367
R1801 B.n560 B.n559 163.367
R1802 B.n556 B.n555 163.367
R1803 B.n552 B.n551 163.367
R1804 B.n548 B.n504 163.367
R1805 B.n704 B.n502 163.367
R1806 B.n704 B.n496 163.367
R1807 B.n712 B.n496 163.367
R1808 B.n712 B.n494 163.367
R1809 B.n716 B.n494 163.367
R1810 B.n716 B.n488 163.367
R1811 B.n724 B.n488 163.367
R1812 B.n724 B.n486 163.367
R1813 B.n728 B.n486 163.367
R1814 B.n728 B.n480 163.367
R1815 B.n736 B.n480 163.367
R1816 B.n736 B.n478 163.367
R1817 B.n740 B.n478 163.367
R1818 B.n740 B.n472 163.367
R1819 B.n748 B.n472 163.367
R1820 B.n748 B.n470 163.367
R1821 B.n752 B.n470 163.367
R1822 B.n752 B.n464 163.367
R1823 B.n760 B.n464 163.367
R1824 B.n760 B.n462 163.367
R1825 B.n764 B.n462 163.367
R1826 B.n764 B.n455 163.367
R1827 B.n772 B.n455 163.367
R1828 B.n772 B.n453 163.367
R1829 B.n776 B.n453 163.367
R1830 B.n776 B.n448 163.367
R1831 B.n784 B.n448 163.367
R1832 B.n784 B.n446 163.367
R1833 B.n788 B.n446 163.367
R1834 B.n788 B.n440 163.367
R1835 B.n796 B.n440 163.367
R1836 B.n796 B.n438 163.367
R1837 B.n800 B.n438 163.367
R1838 B.n800 B.n431 163.367
R1839 B.n808 B.n431 163.367
R1840 B.n808 B.n429 163.367
R1841 B.n812 B.n429 163.367
R1842 B.n812 B.n424 163.367
R1843 B.n820 B.n424 163.367
R1844 B.n820 B.n422 163.367
R1845 B.n824 B.n422 163.367
R1846 B.n824 B.n416 163.367
R1847 B.n832 B.n416 163.367
R1848 B.n832 B.n414 163.367
R1849 B.n836 B.n414 163.367
R1850 B.n836 B.n407 163.367
R1851 B.n844 B.n407 163.367
R1852 B.n844 B.n405 163.367
R1853 B.n848 B.n405 163.367
R1854 B.n848 B.n400 163.367
R1855 B.n856 B.n400 163.367
R1856 B.n856 B.n398 163.367
R1857 B.n860 B.n398 163.367
R1858 B.n860 B.n392 163.367
R1859 B.n868 B.n392 163.367
R1860 B.n868 B.n390 163.367
R1861 B.n872 B.n390 163.367
R1862 B.n872 B.n384 163.367
R1863 B.n880 B.n384 163.367
R1864 B.n880 B.n382 163.367
R1865 B.n884 B.n382 163.367
R1866 B.n884 B.n376 163.367
R1867 B.n892 B.n376 163.367
R1868 B.n892 B.n374 163.367
R1869 B.n896 B.n374 163.367
R1870 B.n896 B.n368 163.367
R1871 B.n904 B.n368 163.367
R1872 B.n904 B.n366 163.367
R1873 B.n908 B.n366 163.367
R1874 B.n908 B.n360 163.367
R1875 B.n916 B.n360 163.367
R1876 B.n916 B.n358 163.367
R1877 B.n920 B.n358 163.367
R1878 B.n920 B.n352 163.367
R1879 B.n928 B.n352 163.367
R1880 B.n928 B.n350 163.367
R1881 B.n933 B.n350 163.367
R1882 B.n933 B.n344 163.367
R1883 B.n941 B.n344 163.367
R1884 B.n942 B.n941 163.367
R1885 B.n942 B.n5 163.367
R1886 B.n6 B.n5 163.367
R1887 B.n7 B.n6 163.367
R1888 B.n947 B.n7 163.367
R1889 B.n947 B.n12 163.367
R1890 B.n13 B.n12 163.367
R1891 B.n14 B.n13 163.367
R1892 B.n952 B.n14 163.367
R1893 B.n952 B.n19 163.367
R1894 B.n20 B.n19 163.367
R1895 B.n21 B.n20 163.367
R1896 B.n957 B.n21 163.367
R1897 B.n957 B.n26 163.367
R1898 B.n27 B.n26 163.367
R1899 B.n28 B.n27 163.367
R1900 B.n962 B.n28 163.367
R1901 B.n962 B.n33 163.367
R1902 B.n34 B.n33 163.367
R1903 B.n35 B.n34 163.367
R1904 B.n967 B.n35 163.367
R1905 B.n967 B.n40 163.367
R1906 B.n41 B.n40 163.367
R1907 B.n42 B.n41 163.367
R1908 B.n972 B.n42 163.367
R1909 B.n972 B.n47 163.367
R1910 B.n48 B.n47 163.367
R1911 B.n49 B.n48 163.367
R1912 B.n977 B.n49 163.367
R1913 B.n977 B.n54 163.367
R1914 B.n55 B.n54 163.367
R1915 B.n56 B.n55 163.367
R1916 B.n982 B.n56 163.367
R1917 B.n982 B.n61 163.367
R1918 B.n62 B.n61 163.367
R1919 B.n63 B.n62 163.367
R1920 B.n987 B.n63 163.367
R1921 B.n987 B.n68 163.367
R1922 B.n69 B.n68 163.367
R1923 B.n70 B.n69 163.367
R1924 B.n992 B.n70 163.367
R1925 B.n992 B.n75 163.367
R1926 B.n76 B.n75 163.367
R1927 B.n77 B.n76 163.367
R1928 B.n997 B.n77 163.367
R1929 B.n997 B.n82 163.367
R1930 B.n83 B.n82 163.367
R1931 B.n84 B.n83 163.367
R1932 B.n1002 B.n84 163.367
R1933 B.n1002 B.n89 163.367
R1934 B.n90 B.n89 163.367
R1935 B.n91 B.n90 163.367
R1936 B.n1007 B.n91 163.367
R1937 B.n1007 B.n96 163.367
R1938 B.n97 B.n96 163.367
R1939 B.n98 B.n97 163.367
R1940 B.n1012 B.n98 163.367
R1941 B.n1012 B.n103 163.367
R1942 B.n104 B.n103 163.367
R1943 B.n105 B.n104 163.367
R1944 B.n1017 B.n105 163.367
R1945 B.n1017 B.n110 163.367
R1946 B.n111 B.n110 163.367
R1947 B.n112 B.n111 163.367
R1948 B.n1022 B.n112 163.367
R1949 B.n1022 B.n117 163.367
R1950 B.n118 B.n117 163.367
R1951 B.n119 B.n118 163.367
R1952 B.n1027 B.n119 163.367
R1953 B.n1027 B.n124 163.367
R1954 B.n125 B.n124 163.367
R1955 B.n126 B.n125 163.367
R1956 B.n1032 B.n126 163.367
R1957 B.n1032 B.n131 163.367
R1958 B.n132 B.n131 163.367
R1959 B.n133 B.n132 163.367
R1960 B.n1037 B.n133 163.367
R1961 B.n1037 B.n138 163.367
R1962 B.n139 B.n138 163.367
R1963 B.n140 B.n139 163.367
R1964 B.n1042 B.n140 163.367
R1965 B.n1042 B.n145 163.367
R1966 B.n146 B.n145 163.367
R1967 B.n195 B.n194 163.367
R1968 B.n199 B.n198 163.367
R1969 B.n203 B.n202 163.367
R1970 B.n207 B.n206 163.367
R1971 B.n211 B.n210 163.367
R1972 B.n215 B.n214 163.367
R1973 B.n219 B.n218 163.367
R1974 B.n223 B.n222 163.367
R1975 B.n227 B.n226 163.367
R1976 B.n231 B.n230 163.367
R1977 B.n235 B.n234 163.367
R1978 B.n239 B.n238 163.367
R1979 B.n243 B.n242 163.367
R1980 B.n247 B.n246 163.367
R1981 B.n251 B.n250 163.367
R1982 B.n255 B.n254 163.367
R1983 B.n259 B.n258 163.367
R1984 B.n263 B.n262 163.367
R1985 B.n267 B.n266 163.367
R1986 B.n271 B.n270 163.367
R1987 B.n275 B.n274 163.367
R1988 B.n280 B.n279 163.367
R1989 B.n284 B.n283 163.367
R1990 B.n288 B.n287 163.367
R1991 B.n292 B.n291 163.367
R1992 B.n296 B.n295 163.367
R1993 B.n300 B.n299 163.367
R1994 B.n304 B.n303 163.367
R1995 B.n308 B.n307 163.367
R1996 B.n312 B.n311 163.367
R1997 B.n316 B.n315 163.367
R1998 B.n320 B.n319 163.367
R1999 B.n324 B.n323 163.367
R2000 B.n328 B.n327 163.367
R2001 B.n332 B.n331 163.367
R2002 B.n336 B.n335 163.367
R2003 B.n340 B.n339 163.367
R2004 B.n1047 B.n185 163.367
R2005 B.n698 B.n501 101.469
R2006 B.n1049 B.n1048 101.469
R2007 B.n546 B.n545 80.2914
R2008 B.n544 B.n543 80.2914
R2009 B.n189 B.n188 80.2914
R2010 B.n187 B.n186 80.2914
R2011 B.n697 B.n696 71.676
R2012 B.n691 B.n505 71.676
R2013 B.n688 B.n506 71.676
R2014 B.n684 B.n507 71.676
R2015 B.n680 B.n508 71.676
R2016 B.n676 B.n509 71.676
R2017 B.n672 B.n510 71.676
R2018 B.n668 B.n511 71.676
R2019 B.n664 B.n512 71.676
R2020 B.n660 B.n513 71.676
R2021 B.n656 B.n514 71.676
R2022 B.n652 B.n515 71.676
R2023 B.n648 B.n516 71.676
R2024 B.n644 B.n517 71.676
R2025 B.n640 B.n518 71.676
R2026 B.n636 B.n519 71.676
R2027 B.n632 B.n520 71.676
R2028 B.n627 B.n521 71.676
R2029 B.n623 B.n522 71.676
R2030 B.n619 B.n523 71.676
R2031 B.n615 B.n524 71.676
R2032 B.n611 B.n525 71.676
R2033 B.n607 B.n526 71.676
R2034 B.n603 B.n527 71.676
R2035 B.n599 B.n528 71.676
R2036 B.n595 B.n529 71.676
R2037 B.n591 B.n530 71.676
R2038 B.n587 B.n531 71.676
R2039 B.n583 B.n532 71.676
R2040 B.n579 B.n533 71.676
R2041 B.n575 B.n534 71.676
R2042 B.n571 B.n535 71.676
R2043 B.n567 B.n536 71.676
R2044 B.n563 B.n537 71.676
R2045 B.n559 B.n538 71.676
R2046 B.n555 B.n539 71.676
R2047 B.n551 B.n540 71.676
R2048 B.n699 B.n504 71.676
R2049 B.n191 B.n147 71.676
R2050 B.n195 B.n148 71.676
R2051 B.n199 B.n149 71.676
R2052 B.n203 B.n150 71.676
R2053 B.n207 B.n151 71.676
R2054 B.n211 B.n152 71.676
R2055 B.n215 B.n153 71.676
R2056 B.n219 B.n154 71.676
R2057 B.n223 B.n155 71.676
R2058 B.n227 B.n156 71.676
R2059 B.n231 B.n157 71.676
R2060 B.n235 B.n158 71.676
R2061 B.n239 B.n159 71.676
R2062 B.n243 B.n160 71.676
R2063 B.n247 B.n161 71.676
R2064 B.n251 B.n162 71.676
R2065 B.n255 B.n163 71.676
R2066 B.n259 B.n164 71.676
R2067 B.n263 B.n165 71.676
R2068 B.n267 B.n166 71.676
R2069 B.n271 B.n167 71.676
R2070 B.n275 B.n168 71.676
R2071 B.n280 B.n169 71.676
R2072 B.n284 B.n170 71.676
R2073 B.n288 B.n171 71.676
R2074 B.n292 B.n172 71.676
R2075 B.n296 B.n173 71.676
R2076 B.n300 B.n174 71.676
R2077 B.n304 B.n175 71.676
R2078 B.n308 B.n176 71.676
R2079 B.n312 B.n177 71.676
R2080 B.n316 B.n178 71.676
R2081 B.n320 B.n179 71.676
R2082 B.n324 B.n180 71.676
R2083 B.n328 B.n181 71.676
R2084 B.n332 B.n182 71.676
R2085 B.n336 B.n183 71.676
R2086 B.n340 B.n184 71.676
R2087 B.n185 B.n184 71.676
R2088 B.n339 B.n183 71.676
R2089 B.n335 B.n182 71.676
R2090 B.n331 B.n181 71.676
R2091 B.n327 B.n180 71.676
R2092 B.n323 B.n179 71.676
R2093 B.n319 B.n178 71.676
R2094 B.n315 B.n177 71.676
R2095 B.n311 B.n176 71.676
R2096 B.n307 B.n175 71.676
R2097 B.n303 B.n174 71.676
R2098 B.n299 B.n173 71.676
R2099 B.n295 B.n172 71.676
R2100 B.n291 B.n171 71.676
R2101 B.n287 B.n170 71.676
R2102 B.n283 B.n169 71.676
R2103 B.n279 B.n168 71.676
R2104 B.n274 B.n167 71.676
R2105 B.n270 B.n166 71.676
R2106 B.n266 B.n165 71.676
R2107 B.n262 B.n164 71.676
R2108 B.n258 B.n163 71.676
R2109 B.n254 B.n162 71.676
R2110 B.n250 B.n161 71.676
R2111 B.n246 B.n160 71.676
R2112 B.n242 B.n159 71.676
R2113 B.n238 B.n158 71.676
R2114 B.n234 B.n157 71.676
R2115 B.n230 B.n156 71.676
R2116 B.n226 B.n155 71.676
R2117 B.n222 B.n154 71.676
R2118 B.n218 B.n153 71.676
R2119 B.n214 B.n152 71.676
R2120 B.n210 B.n151 71.676
R2121 B.n206 B.n150 71.676
R2122 B.n202 B.n149 71.676
R2123 B.n198 B.n148 71.676
R2124 B.n194 B.n147 71.676
R2125 B.n697 B.n542 71.676
R2126 B.n689 B.n505 71.676
R2127 B.n685 B.n506 71.676
R2128 B.n681 B.n507 71.676
R2129 B.n677 B.n508 71.676
R2130 B.n673 B.n509 71.676
R2131 B.n669 B.n510 71.676
R2132 B.n665 B.n511 71.676
R2133 B.n661 B.n512 71.676
R2134 B.n657 B.n513 71.676
R2135 B.n653 B.n514 71.676
R2136 B.n649 B.n515 71.676
R2137 B.n645 B.n516 71.676
R2138 B.n641 B.n517 71.676
R2139 B.n637 B.n518 71.676
R2140 B.n633 B.n519 71.676
R2141 B.n628 B.n520 71.676
R2142 B.n624 B.n521 71.676
R2143 B.n620 B.n522 71.676
R2144 B.n616 B.n523 71.676
R2145 B.n612 B.n524 71.676
R2146 B.n608 B.n525 71.676
R2147 B.n604 B.n526 71.676
R2148 B.n600 B.n527 71.676
R2149 B.n596 B.n528 71.676
R2150 B.n592 B.n529 71.676
R2151 B.n588 B.n530 71.676
R2152 B.n584 B.n531 71.676
R2153 B.n580 B.n532 71.676
R2154 B.n576 B.n533 71.676
R2155 B.n572 B.n534 71.676
R2156 B.n568 B.n535 71.676
R2157 B.n564 B.n536 71.676
R2158 B.n560 B.n537 71.676
R2159 B.n556 B.n538 71.676
R2160 B.n552 B.n539 71.676
R2161 B.n548 B.n540 71.676
R2162 B.n700 B.n699 71.676
R2163 B.n547 B.n546 59.5399
R2164 B.n630 B.n544 59.5399
R2165 B.n190 B.n189 59.5399
R2166 B.n277 B.n187 59.5399
R2167 B.n705 B.n501 51.1109
R2168 B.n705 B.n497 51.1109
R2169 B.n711 B.n497 51.1109
R2170 B.n711 B.n493 51.1109
R2171 B.n717 B.n493 51.1109
R2172 B.n717 B.n489 51.1109
R2173 B.n723 B.n489 51.1109
R2174 B.n723 B.n485 51.1109
R2175 B.n729 B.n485 51.1109
R2176 B.n735 B.n481 51.1109
R2177 B.n735 B.n477 51.1109
R2178 B.n741 B.n477 51.1109
R2179 B.n741 B.n473 51.1109
R2180 B.n747 B.n473 51.1109
R2181 B.n747 B.n469 51.1109
R2182 B.n753 B.n469 51.1109
R2183 B.n753 B.n465 51.1109
R2184 B.n759 B.n465 51.1109
R2185 B.n759 B.n461 51.1109
R2186 B.n765 B.n461 51.1109
R2187 B.n765 B.n456 51.1109
R2188 B.n771 B.n456 51.1109
R2189 B.n771 B.n457 51.1109
R2190 B.n777 B.n449 51.1109
R2191 B.n783 B.n449 51.1109
R2192 B.n783 B.n445 51.1109
R2193 B.n789 B.n445 51.1109
R2194 B.n789 B.n441 51.1109
R2195 B.n795 B.n441 51.1109
R2196 B.n795 B.n437 51.1109
R2197 B.n801 B.n437 51.1109
R2198 B.n801 B.n432 51.1109
R2199 B.n807 B.n432 51.1109
R2200 B.n807 B.n433 51.1109
R2201 B.n813 B.n425 51.1109
R2202 B.n819 B.n425 51.1109
R2203 B.n819 B.n421 51.1109
R2204 B.n825 B.n421 51.1109
R2205 B.n825 B.n417 51.1109
R2206 B.n831 B.n417 51.1109
R2207 B.n831 B.n413 51.1109
R2208 B.n837 B.n413 51.1109
R2209 B.n837 B.n408 51.1109
R2210 B.n843 B.n408 51.1109
R2211 B.n843 B.n409 51.1109
R2212 B.n849 B.n401 51.1109
R2213 B.n855 B.n401 51.1109
R2214 B.n855 B.n397 51.1109
R2215 B.n861 B.n397 51.1109
R2216 B.n861 B.n393 51.1109
R2217 B.n867 B.n393 51.1109
R2218 B.n867 B.n389 51.1109
R2219 B.n873 B.n389 51.1109
R2220 B.n873 B.n385 51.1109
R2221 B.n879 B.n385 51.1109
R2222 B.n879 B.n381 51.1109
R2223 B.n885 B.n381 51.1109
R2224 B.n891 B.n377 51.1109
R2225 B.n891 B.n373 51.1109
R2226 B.n897 B.n373 51.1109
R2227 B.n897 B.n369 51.1109
R2228 B.n903 B.n369 51.1109
R2229 B.n903 B.n365 51.1109
R2230 B.n909 B.n365 51.1109
R2231 B.n909 B.n361 51.1109
R2232 B.n915 B.n361 51.1109
R2233 B.n915 B.n357 51.1109
R2234 B.n921 B.n357 51.1109
R2235 B.n927 B.n353 51.1109
R2236 B.n927 B.n349 51.1109
R2237 B.n934 B.n349 51.1109
R2238 B.n934 B.n345 51.1109
R2239 B.n940 B.n345 51.1109
R2240 B.n940 B.n4 51.1109
R2241 B.n1210 B.n4 51.1109
R2242 B.n1210 B.n1209 51.1109
R2243 B.n1209 B.n1208 51.1109
R2244 B.n1208 B.n8 51.1109
R2245 B.n1202 B.n8 51.1109
R2246 B.n1202 B.n1201 51.1109
R2247 B.n1201 B.n1200 51.1109
R2248 B.n1200 B.n15 51.1109
R2249 B.n1194 B.n1193 51.1109
R2250 B.n1193 B.n1192 51.1109
R2251 B.n1192 B.n22 51.1109
R2252 B.n1186 B.n22 51.1109
R2253 B.n1186 B.n1185 51.1109
R2254 B.n1185 B.n1184 51.1109
R2255 B.n1184 B.n29 51.1109
R2256 B.n1178 B.n29 51.1109
R2257 B.n1178 B.n1177 51.1109
R2258 B.n1177 B.n1176 51.1109
R2259 B.n1176 B.n36 51.1109
R2260 B.n1170 B.n1169 51.1109
R2261 B.n1169 B.n1168 51.1109
R2262 B.n1168 B.n43 51.1109
R2263 B.n1162 B.n43 51.1109
R2264 B.n1162 B.n1161 51.1109
R2265 B.n1161 B.n1160 51.1109
R2266 B.n1160 B.n50 51.1109
R2267 B.n1154 B.n50 51.1109
R2268 B.n1154 B.n1153 51.1109
R2269 B.n1153 B.n1152 51.1109
R2270 B.n1152 B.n57 51.1109
R2271 B.n1146 B.n57 51.1109
R2272 B.n1145 B.n1144 51.1109
R2273 B.n1144 B.n64 51.1109
R2274 B.n1138 B.n64 51.1109
R2275 B.n1138 B.n1137 51.1109
R2276 B.n1137 B.n1136 51.1109
R2277 B.n1136 B.n71 51.1109
R2278 B.n1130 B.n71 51.1109
R2279 B.n1130 B.n1129 51.1109
R2280 B.n1129 B.n1128 51.1109
R2281 B.n1128 B.n78 51.1109
R2282 B.n1122 B.n78 51.1109
R2283 B.n1121 B.n1120 51.1109
R2284 B.n1120 B.n85 51.1109
R2285 B.n1114 B.n85 51.1109
R2286 B.n1114 B.n1113 51.1109
R2287 B.n1113 B.n1112 51.1109
R2288 B.n1112 B.n92 51.1109
R2289 B.n1106 B.n92 51.1109
R2290 B.n1106 B.n1105 51.1109
R2291 B.n1105 B.n1104 51.1109
R2292 B.n1104 B.n99 51.1109
R2293 B.n1098 B.n99 51.1109
R2294 B.n1097 B.n1096 51.1109
R2295 B.n1096 B.n106 51.1109
R2296 B.n1090 B.n106 51.1109
R2297 B.n1090 B.n1089 51.1109
R2298 B.n1089 B.n1088 51.1109
R2299 B.n1088 B.n113 51.1109
R2300 B.n1082 B.n113 51.1109
R2301 B.n1082 B.n1081 51.1109
R2302 B.n1081 B.n1080 51.1109
R2303 B.n1080 B.n120 51.1109
R2304 B.n1074 B.n120 51.1109
R2305 B.n1074 B.n1073 51.1109
R2306 B.n1073 B.n1072 51.1109
R2307 B.n1072 B.n127 51.1109
R2308 B.n1066 B.n1065 51.1109
R2309 B.n1065 B.n1064 51.1109
R2310 B.n1064 B.n134 51.1109
R2311 B.n1058 B.n134 51.1109
R2312 B.n1058 B.n1057 51.1109
R2313 B.n1057 B.n1056 51.1109
R2314 B.n1056 B.n141 51.1109
R2315 B.n1050 B.n141 51.1109
R2316 B.n1050 B.n1049 51.1109
R2317 B.n409 B.t7 48.856
R2318 B.t1 B.n1145 48.856
R2319 B.t6 B.n377 44.3462
R2320 B.t5 B.n36 44.3462
R2321 B.t18 B.n481 39.8365
R2322 B.n433 B.t2 39.8365
R2323 B.t3 B.n1121 39.8365
R2324 B.t11 B.n127 39.8365
R2325 B.n192 B.n143 35.7468
R2326 B.n1046 B.n1045 35.7468
R2327 B.n702 B.n701 35.7468
R2328 B.n695 B.n499 35.7468
R2329 B.t0 B.n353 35.3268
R2330 B.t4 B.n15 35.3268
R2331 B.n457 B.t8 30.817
R2332 B.t9 B.n1097 30.817
R2333 B.n777 B.t8 20.2943
R2334 B.n1098 B.t9 20.2943
R2335 B B.n1212 18.0485
R2336 B.n921 B.t0 15.7846
R2337 B.n1194 B.t4 15.7846
R2338 B.n729 B.t18 11.2748
R2339 B.n813 B.t2 11.2748
R2340 B.n1122 B.t3 11.2748
R2341 B.n1066 B.t11 11.2748
R2342 B.n193 B.n192 10.6151
R2343 B.n196 B.n193 10.6151
R2344 B.n197 B.n196 10.6151
R2345 B.n200 B.n197 10.6151
R2346 B.n201 B.n200 10.6151
R2347 B.n204 B.n201 10.6151
R2348 B.n205 B.n204 10.6151
R2349 B.n208 B.n205 10.6151
R2350 B.n209 B.n208 10.6151
R2351 B.n212 B.n209 10.6151
R2352 B.n213 B.n212 10.6151
R2353 B.n216 B.n213 10.6151
R2354 B.n217 B.n216 10.6151
R2355 B.n220 B.n217 10.6151
R2356 B.n221 B.n220 10.6151
R2357 B.n224 B.n221 10.6151
R2358 B.n225 B.n224 10.6151
R2359 B.n228 B.n225 10.6151
R2360 B.n229 B.n228 10.6151
R2361 B.n232 B.n229 10.6151
R2362 B.n233 B.n232 10.6151
R2363 B.n236 B.n233 10.6151
R2364 B.n237 B.n236 10.6151
R2365 B.n240 B.n237 10.6151
R2366 B.n241 B.n240 10.6151
R2367 B.n244 B.n241 10.6151
R2368 B.n245 B.n244 10.6151
R2369 B.n248 B.n245 10.6151
R2370 B.n249 B.n248 10.6151
R2371 B.n252 B.n249 10.6151
R2372 B.n253 B.n252 10.6151
R2373 B.n256 B.n253 10.6151
R2374 B.n257 B.n256 10.6151
R2375 B.n261 B.n260 10.6151
R2376 B.n264 B.n261 10.6151
R2377 B.n265 B.n264 10.6151
R2378 B.n268 B.n265 10.6151
R2379 B.n269 B.n268 10.6151
R2380 B.n272 B.n269 10.6151
R2381 B.n273 B.n272 10.6151
R2382 B.n276 B.n273 10.6151
R2383 B.n281 B.n278 10.6151
R2384 B.n282 B.n281 10.6151
R2385 B.n285 B.n282 10.6151
R2386 B.n286 B.n285 10.6151
R2387 B.n289 B.n286 10.6151
R2388 B.n290 B.n289 10.6151
R2389 B.n293 B.n290 10.6151
R2390 B.n294 B.n293 10.6151
R2391 B.n297 B.n294 10.6151
R2392 B.n298 B.n297 10.6151
R2393 B.n301 B.n298 10.6151
R2394 B.n302 B.n301 10.6151
R2395 B.n305 B.n302 10.6151
R2396 B.n306 B.n305 10.6151
R2397 B.n309 B.n306 10.6151
R2398 B.n310 B.n309 10.6151
R2399 B.n313 B.n310 10.6151
R2400 B.n314 B.n313 10.6151
R2401 B.n317 B.n314 10.6151
R2402 B.n318 B.n317 10.6151
R2403 B.n321 B.n318 10.6151
R2404 B.n322 B.n321 10.6151
R2405 B.n325 B.n322 10.6151
R2406 B.n326 B.n325 10.6151
R2407 B.n329 B.n326 10.6151
R2408 B.n330 B.n329 10.6151
R2409 B.n333 B.n330 10.6151
R2410 B.n334 B.n333 10.6151
R2411 B.n337 B.n334 10.6151
R2412 B.n338 B.n337 10.6151
R2413 B.n341 B.n338 10.6151
R2414 B.n342 B.n341 10.6151
R2415 B.n1046 B.n342 10.6151
R2416 B.n703 B.n702 10.6151
R2417 B.n703 B.n495 10.6151
R2418 B.n713 B.n495 10.6151
R2419 B.n714 B.n713 10.6151
R2420 B.n715 B.n714 10.6151
R2421 B.n715 B.n487 10.6151
R2422 B.n725 B.n487 10.6151
R2423 B.n726 B.n725 10.6151
R2424 B.n727 B.n726 10.6151
R2425 B.n727 B.n479 10.6151
R2426 B.n737 B.n479 10.6151
R2427 B.n738 B.n737 10.6151
R2428 B.n739 B.n738 10.6151
R2429 B.n739 B.n471 10.6151
R2430 B.n749 B.n471 10.6151
R2431 B.n750 B.n749 10.6151
R2432 B.n751 B.n750 10.6151
R2433 B.n751 B.n463 10.6151
R2434 B.n761 B.n463 10.6151
R2435 B.n762 B.n761 10.6151
R2436 B.n763 B.n762 10.6151
R2437 B.n763 B.n454 10.6151
R2438 B.n773 B.n454 10.6151
R2439 B.n774 B.n773 10.6151
R2440 B.n775 B.n774 10.6151
R2441 B.n775 B.n447 10.6151
R2442 B.n785 B.n447 10.6151
R2443 B.n786 B.n785 10.6151
R2444 B.n787 B.n786 10.6151
R2445 B.n787 B.n439 10.6151
R2446 B.n797 B.n439 10.6151
R2447 B.n798 B.n797 10.6151
R2448 B.n799 B.n798 10.6151
R2449 B.n799 B.n430 10.6151
R2450 B.n809 B.n430 10.6151
R2451 B.n810 B.n809 10.6151
R2452 B.n811 B.n810 10.6151
R2453 B.n811 B.n423 10.6151
R2454 B.n821 B.n423 10.6151
R2455 B.n822 B.n821 10.6151
R2456 B.n823 B.n822 10.6151
R2457 B.n823 B.n415 10.6151
R2458 B.n833 B.n415 10.6151
R2459 B.n834 B.n833 10.6151
R2460 B.n835 B.n834 10.6151
R2461 B.n835 B.n406 10.6151
R2462 B.n845 B.n406 10.6151
R2463 B.n846 B.n845 10.6151
R2464 B.n847 B.n846 10.6151
R2465 B.n847 B.n399 10.6151
R2466 B.n857 B.n399 10.6151
R2467 B.n858 B.n857 10.6151
R2468 B.n859 B.n858 10.6151
R2469 B.n859 B.n391 10.6151
R2470 B.n869 B.n391 10.6151
R2471 B.n870 B.n869 10.6151
R2472 B.n871 B.n870 10.6151
R2473 B.n871 B.n383 10.6151
R2474 B.n881 B.n383 10.6151
R2475 B.n882 B.n881 10.6151
R2476 B.n883 B.n882 10.6151
R2477 B.n883 B.n375 10.6151
R2478 B.n893 B.n375 10.6151
R2479 B.n894 B.n893 10.6151
R2480 B.n895 B.n894 10.6151
R2481 B.n895 B.n367 10.6151
R2482 B.n905 B.n367 10.6151
R2483 B.n906 B.n905 10.6151
R2484 B.n907 B.n906 10.6151
R2485 B.n907 B.n359 10.6151
R2486 B.n917 B.n359 10.6151
R2487 B.n918 B.n917 10.6151
R2488 B.n919 B.n918 10.6151
R2489 B.n919 B.n351 10.6151
R2490 B.n929 B.n351 10.6151
R2491 B.n930 B.n929 10.6151
R2492 B.n932 B.n930 10.6151
R2493 B.n932 B.n931 10.6151
R2494 B.n931 B.n343 10.6151
R2495 B.n943 B.n343 10.6151
R2496 B.n944 B.n943 10.6151
R2497 B.n945 B.n944 10.6151
R2498 B.n946 B.n945 10.6151
R2499 B.n948 B.n946 10.6151
R2500 B.n949 B.n948 10.6151
R2501 B.n950 B.n949 10.6151
R2502 B.n951 B.n950 10.6151
R2503 B.n953 B.n951 10.6151
R2504 B.n954 B.n953 10.6151
R2505 B.n955 B.n954 10.6151
R2506 B.n956 B.n955 10.6151
R2507 B.n958 B.n956 10.6151
R2508 B.n959 B.n958 10.6151
R2509 B.n960 B.n959 10.6151
R2510 B.n961 B.n960 10.6151
R2511 B.n963 B.n961 10.6151
R2512 B.n964 B.n963 10.6151
R2513 B.n965 B.n964 10.6151
R2514 B.n966 B.n965 10.6151
R2515 B.n968 B.n966 10.6151
R2516 B.n969 B.n968 10.6151
R2517 B.n970 B.n969 10.6151
R2518 B.n971 B.n970 10.6151
R2519 B.n973 B.n971 10.6151
R2520 B.n974 B.n973 10.6151
R2521 B.n975 B.n974 10.6151
R2522 B.n976 B.n975 10.6151
R2523 B.n978 B.n976 10.6151
R2524 B.n979 B.n978 10.6151
R2525 B.n980 B.n979 10.6151
R2526 B.n981 B.n980 10.6151
R2527 B.n983 B.n981 10.6151
R2528 B.n984 B.n983 10.6151
R2529 B.n985 B.n984 10.6151
R2530 B.n986 B.n985 10.6151
R2531 B.n988 B.n986 10.6151
R2532 B.n989 B.n988 10.6151
R2533 B.n990 B.n989 10.6151
R2534 B.n991 B.n990 10.6151
R2535 B.n993 B.n991 10.6151
R2536 B.n994 B.n993 10.6151
R2537 B.n995 B.n994 10.6151
R2538 B.n996 B.n995 10.6151
R2539 B.n998 B.n996 10.6151
R2540 B.n999 B.n998 10.6151
R2541 B.n1000 B.n999 10.6151
R2542 B.n1001 B.n1000 10.6151
R2543 B.n1003 B.n1001 10.6151
R2544 B.n1004 B.n1003 10.6151
R2545 B.n1005 B.n1004 10.6151
R2546 B.n1006 B.n1005 10.6151
R2547 B.n1008 B.n1006 10.6151
R2548 B.n1009 B.n1008 10.6151
R2549 B.n1010 B.n1009 10.6151
R2550 B.n1011 B.n1010 10.6151
R2551 B.n1013 B.n1011 10.6151
R2552 B.n1014 B.n1013 10.6151
R2553 B.n1015 B.n1014 10.6151
R2554 B.n1016 B.n1015 10.6151
R2555 B.n1018 B.n1016 10.6151
R2556 B.n1019 B.n1018 10.6151
R2557 B.n1020 B.n1019 10.6151
R2558 B.n1021 B.n1020 10.6151
R2559 B.n1023 B.n1021 10.6151
R2560 B.n1024 B.n1023 10.6151
R2561 B.n1025 B.n1024 10.6151
R2562 B.n1026 B.n1025 10.6151
R2563 B.n1028 B.n1026 10.6151
R2564 B.n1029 B.n1028 10.6151
R2565 B.n1030 B.n1029 10.6151
R2566 B.n1031 B.n1030 10.6151
R2567 B.n1033 B.n1031 10.6151
R2568 B.n1034 B.n1033 10.6151
R2569 B.n1035 B.n1034 10.6151
R2570 B.n1036 B.n1035 10.6151
R2571 B.n1038 B.n1036 10.6151
R2572 B.n1039 B.n1038 10.6151
R2573 B.n1040 B.n1039 10.6151
R2574 B.n1041 B.n1040 10.6151
R2575 B.n1043 B.n1041 10.6151
R2576 B.n1044 B.n1043 10.6151
R2577 B.n1045 B.n1044 10.6151
R2578 B.n695 B.n694 10.6151
R2579 B.n694 B.n693 10.6151
R2580 B.n693 B.n692 10.6151
R2581 B.n692 B.n690 10.6151
R2582 B.n690 B.n687 10.6151
R2583 B.n687 B.n686 10.6151
R2584 B.n686 B.n683 10.6151
R2585 B.n683 B.n682 10.6151
R2586 B.n682 B.n679 10.6151
R2587 B.n679 B.n678 10.6151
R2588 B.n678 B.n675 10.6151
R2589 B.n675 B.n674 10.6151
R2590 B.n674 B.n671 10.6151
R2591 B.n671 B.n670 10.6151
R2592 B.n670 B.n667 10.6151
R2593 B.n667 B.n666 10.6151
R2594 B.n666 B.n663 10.6151
R2595 B.n663 B.n662 10.6151
R2596 B.n662 B.n659 10.6151
R2597 B.n659 B.n658 10.6151
R2598 B.n658 B.n655 10.6151
R2599 B.n655 B.n654 10.6151
R2600 B.n654 B.n651 10.6151
R2601 B.n651 B.n650 10.6151
R2602 B.n650 B.n647 10.6151
R2603 B.n647 B.n646 10.6151
R2604 B.n646 B.n643 10.6151
R2605 B.n643 B.n642 10.6151
R2606 B.n642 B.n639 10.6151
R2607 B.n639 B.n638 10.6151
R2608 B.n638 B.n635 10.6151
R2609 B.n635 B.n634 10.6151
R2610 B.n634 B.n631 10.6151
R2611 B.n629 B.n626 10.6151
R2612 B.n626 B.n625 10.6151
R2613 B.n625 B.n622 10.6151
R2614 B.n622 B.n621 10.6151
R2615 B.n621 B.n618 10.6151
R2616 B.n618 B.n617 10.6151
R2617 B.n617 B.n614 10.6151
R2618 B.n614 B.n613 10.6151
R2619 B.n610 B.n609 10.6151
R2620 B.n609 B.n606 10.6151
R2621 B.n606 B.n605 10.6151
R2622 B.n605 B.n602 10.6151
R2623 B.n602 B.n601 10.6151
R2624 B.n601 B.n598 10.6151
R2625 B.n598 B.n597 10.6151
R2626 B.n597 B.n594 10.6151
R2627 B.n594 B.n593 10.6151
R2628 B.n593 B.n590 10.6151
R2629 B.n590 B.n589 10.6151
R2630 B.n589 B.n586 10.6151
R2631 B.n586 B.n585 10.6151
R2632 B.n585 B.n582 10.6151
R2633 B.n582 B.n581 10.6151
R2634 B.n581 B.n578 10.6151
R2635 B.n578 B.n577 10.6151
R2636 B.n577 B.n574 10.6151
R2637 B.n574 B.n573 10.6151
R2638 B.n573 B.n570 10.6151
R2639 B.n570 B.n569 10.6151
R2640 B.n569 B.n566 10.6151
R2641 B.n566 B.n565 10.6151
R2642 B.n565 B.n562 10.6151
R2643 B.n562 B.n561 10.6151
R2644 B.n561 B.n558 10.6151
R2645 B.n558 B.n557 10.6151
R2646 B.n557 B.n554 10.6151
R2647 B.n554 B.n553 10.6151
R2648 B.n553 B.n550 10.6151
R2649 B.n550 B.n549 10.6151
R2650 B.n549 B.n503 10.6151
R2651 B.n701 B.n503 10.6151
R2652 B.n707 B.n499 10.6151
R2653 B.n708 B.n707 10.6151
R2654 B.n709 B.n708 10.6151
R2655 B.n709 B.n491 10.6151
R2656 B.n719 B.n491 10.6151
R2657 B.n720 B.n719 10.6151
R2658 B.n721 B.n720 10.6151
R2659 B.n721 B.n483 10.6151
R2660 B.n731 B.n483 10.6151
R2661 B.n732 B.n731 10.6151
R2662 B.n733 B.n732 10.6151
R2663 B.n733 B.n475 10.6151
R2664 B.n743 B.n475 10.6151
R2665 B.n744 B.n743 10.6151
R2666 B.n745 B.n744 10.6151
R2667 B.n745 B.n467 10.6151
R2668 B.n755 B.n467 10.6151
R2669 B.n756 B.n755 10.6151
R2670 B.n757 B.n756 10.6151
R2671 B.n757 B.n459 10.6151
R2672 B.n767 B.n459 10.6151
R2673 B.n768 B.n767 10.6151
R2674 B.n769 B.n768 10.6151
R2675 B.n769 B.n451 10.6151
R2676 B.n779 B.n451 10.6151
R2677 B.n780 B.n779 10.6151
R2678 B.n781 B.n780 10.6151
R2679 B.n781 B.n443 10.6151
R2680 B.n791 B.n443 10.6151
R2681 B.n792 B.n791 10.6151
R2682 B.n793 B.n792 10.6151
R2683 B.n793 B.n435 10.6151
R2684 B.n803 B.n435 10.6151
R2685 B.n804 B.n803 10.6151
R2686 B.n805 B.n804 10.6151
R2687 B.n805 B.n427 10.6151
R2688 B.n815 B.n427 10.6151
R2689 B.n816 B.n815 10.6151
R2690 B.n817 B.n816 10.6151
R2691 B.n817 B.n419 10.6151
R2692 B.n827 B.n419 10.6151
R2693 B.n828 B.n827 10.6151
R2694 B.n829 B.n828 10.6151
R2695 B.n829 B.n411 10.6151
R2696 B.n839 B.n411 10.6151
R2697 B.n840 B.n839 10.6151
R2698 B.n841 B.n840 10.6151
R2699 B.n841 B.n403 10.6151
R2700 B.n851 B.n403 10.6151
R2701 B.n852 B.n851 10.6151
R2702 B.n853 B.n852 10.6151
R2703 B.n853 B.n395 10.6151
R2704 B.n863 B.n395 10.6151
R2705 B.n864 B.n863 10.6151
R2706 B.n865 B.n864 10.6151
R2707 B.n865 B.n387 10.6151
R2708 B.n875 B.n387 10.6151
R2709 B.n876 B.n875 10.6151
R2710 B.n877 B.n876 10.6151
R2711 B.n877 B.n379 10.6151
R2712 B.n887 B.n379 10.6151
R2713 B.n888 B.n887 10.6151
R2714 B.n889 B.n888 10.6151
R2715 B.n889 B.n371 10.6151
R2716 B.n899 B.n371 10.6151
R2717 B.n900 B.n899 10.6151
R2718 B.n901 B.n900 10.6151
R2719 B.n901 B.n363 10.6151
R2720 B.n911 B.n363 10.6151
R2721 B.n912 B.n911 10.6151
R2722 B.n913 B.n912 10.6151
R2723 B.n913 B.n355 10.6151
R2724 B.n923 B.n355 10.6151
R2725 B.n924 B.n923 10.6151
R2726 B.n925 B.n924 10.6151
R2727 B.n925 B.n347 10.6151
R2728 B.n936 B.n347 10.6151
R2729 B.n937 B.n936 10.6151
R2730 B.n938 B.n937 10.6151
R2731 B.n938 B.n0 10.6151
R2732 B.n1206 B.n1 10.6151
R2733 B.n1206 B.n1205 10.6151
R2734 B.n1205 B.n1204 10.6151
R2735 B.n1204 B.n10 10.6151
R2736 B.n1198 B.n10 10.6151
R2737 B.n1198 B.n1197 10.6151
R2738 B.n1197 B.n1196 10.6151
R2739 B.n1196 B.n17 10.6151
R2740 B.n1190 B.n17 10.6151
R2741 B.n1190 B.n1189 10.6151
R2742 B.n1189 B.n1188 10.6151
R2743 B.n1188 B.n24 10.6151
R2744 B.n1182 B.n24 10.6151
R2745 B.n1182 B.n1181 10.6151
R2746 B.n1181 B.n1180 10.6151
R2747 B.n1180 B.n31 10.6151
R2748 B.n1174 B.n31 10.6151
R2749 B.n1174 B.n1173 10.6151
R2750 B.n1173 B.n1172 10.6151
R2751 B.n1172 B.n38 10.6151
R2752 B.n1166 B.n38 10.6151
R2753 B.n1166 B.n1165 10.6151
R2754 B.n1165 B.n1164 10.6151
R2755 B.n1164 B.n45 10.6151
R2756 B.n1158 B.n45 10.6151
R2757 B.n1158 B.n1157 10.6151
R2758 B.n1157 B.n1156 10.6151
R2759 B.n1156 B.n52 10.6151
R2760 B.n1150 B.n52 10.6151
R2761 B.n1150 B.n1149 10.6151
R2762 B.n1149 B.n1148 10.6151
R2763 B.n1148 B.n59 10.6151
R2764 B.n1142 B.n59 10.6151
R2765 B.n1142 B.n1141 10.6151
R2766 B.n1141 B.n1140 10.6151
R2767 B.n1140 B.n66 10.6151
R2768 B.n1134 B.n66 10.6151
R2769 B.n1134 B.n1133 10.6151
R2770 B.n1133 B.n1132 10.6151
R2771 B.n1132 B.n73 10.6151
R2772 B.n1126 B.n73 10.6151
R2773 B.n1126 B.n1125 10.6151
R2774 B.n1125 B.n1124 10.6151
R2775 B.n1124 B.n80 10.6151
R2776 B.n1118 B.n80 10.6151
R2777 B.n1118 B.n1117 10.6151
R2778 B.n1117 B.n1116 10.6151
R2779 B.n1116 B.n87 10.6151
R2780 B.n1110 B.n87 10.6151
R2781 B.n1110 B.n1109 10.6151
R2782 B.n1109 B.n1108 10.6151
R2783 B.n1108 B.n94 10.6151
R2784 B.n1102 B.n94 10.6151
R2785 B.n1102 B.n1101 10.6151
R2786 B.n1101 B.n1100 10.6151
R2787 B.n1100 B.n101 10.6151
R2788 B.n1094 B.n101 10.6151
R2789 B.n1094 B.n1093 10.6151
R2790 B.n1093 B.n1092 10.6151
R2791 B.n1092 B.n108 10.6151
R2792 B.n1086 B.n108 10.6151
R2793 B.n1086 B.n1085 10.6151
R2794 B.n1085 B.n1084 10.6151
R2795 B.n1084 B.n115 10.6151
R2796 B.n1078 B.n115 10.6151
R2797 B.n1078 B.n1077 10.6151
R2798 B.n1077 B.n1076 10.6151
R2799 B.n1076 B.n122 10.6151
R2800 B.n1070 B.n122 10.6151
R2801 B.n1070 B.n1069 10.6151
R2802 B.n1069 B.n1068 10.6151
R2803 B.n1068 B.n129 10.6151
R2804 B.n1062 B.n129 10.6151
R2805 B.n1062 B.n1061 10.6151
R2806 B.n1061 B.n1060 10.6151
R2807 B.n1060 B.n136 10.6151
R2808 B.n1054 B.n136 10.6151
R2809 B.n1054 B.n1053 10.6151
R2810 B.n1053 B.n1052 10.6151
R2811 B.n1052 B.n143 10.6151
R2812 B.n885 B.t6 6.76511
R2813 B.n1170 B.t5 6.76511
R2814 B.n260 B.n190 6.5566
R2815 B.n277 B.n276 6.5566
R2816 B.n630 B.n629 6.5566
R2817 B.n613 B.n547 6.5566
R2818 B.n257 B.n190 4.05904
R2819 B.n278 B.n277 4.05904
R2820 B.n631 B.n630 4.05904
R2821 B.n610 B.n547 4.05904
R2822 B.n1212 B.n0 2.81026
R2823 B.n1212 B.n1 2.81026
R2824 B.n849 B.t7 2.25537
R2825 B.n1146 B.t1 2.25537
R2826 VN.n110 VN.n109 161.3
R2827 VN.n108 VN.n57 161.3
R2828 VN.n107 VN.n106 161.3
R2829 VN.n105 VN.n58 161.3
R2830 VN.n104 VN.n103 161.3
R2831 VN.n102 VN.n59 161.3
R2832 VN.n101 VN.n100 161.3
R2833 VN.n99 VN.n60 161.3
R2834 VN.n98 VN.n97 161.3
R2835 VN.n95 VN.n61 161.3
R2836 VN.n94 VN.n93 161.3
R2837 VN.n92 VN.n62 161.3
R2838 VN.n91 VN.n90 161.3
R2839 VN.n89 VN.n63 161.3
R2840 VN.n88 VN.n87 161.3
R2841 VN.n86 VN.n64 161.3
R2842 VN.n85 VN.n84 161.3
R2843 VN.n82 VN.n65 161.3
R2844 VN.n81 VN.n80 161.3
R2845 VN.n79 VN.n66 161.3
R2846 VN.n78 VN.n77 161.3
R2847 VN.n76 VN.n67 161.3
R2848 VN.n75 VN.n74 161.3
R2849 VN.n73 VN.n68 161.3
R2850 VN.n72 VN.n71 161.3
R2851 VN.n54 VN.n53 161.3
R2852 VN.n52 VN.n1 161.3
R2853 VN.n51 VN.n50 161.3
R2854 VN.n49 VN.n2 161.3
R2855 VN.n48 VN.n47 161.3
R2856 VN.n46 VN.n3 161.3
R2857 VN.n45 VN.n44 161.3
R2858 VN.n43 VN.n4 161.3
R2859 VN.n42 VN.n41 161.3
R2860 VN.n39 VN.n5 161.3
R2861 VN.n38 VN.n37 161.3
R2862 VN.n36 VN.n6 161.3
R2863 VN.n35 VN.n34 161.3
R2864 VN.n33 VN.n7 161.3
R2865 VN.n32 VN.n31 161.3
R2866 VN.n30 VN.n8 161.3
R2867 VN.n29 VN.n28 161.3
R2868 VN.n26 VN.n9 161.3
R2869 VN.n25 VN.n24 161.3
R2870 VN.n23 VN.n10 161.3
R2871 VN.n22 VN.n21 161.3
R2872 VN.n20 VN.n11 161.3
R2873 VN.n19 VN.n18 161.3
R2874 VN.n17 VN.n12 161.3
R2875 VN.n16 VN.n15 161.3
R2876 VN.n69 VN.t6 91.7701
R2877 VN.n13 VN.t9 91.7701
R2878 VN.n55 VN.n0 88.77
R2879 VN.n111 VN.n56 88.77
R2880 VN.n14 VN.t0 59.2068
R2881 VN.n27 VN.t4 59.2068
R2882 VN.n40 VN.t3 59.2068
R2883 VN.n0 VN.t8 59.2068
R2884 VN.n70 VN.t1 59.2068
R2885 VN.n83 VN.t7 59.2068
R2886 VN.n96 VN.t2 59.2068
R2887 VN.n56 VN.t5 59.2068
R2888 VN VN.n111 57.8921
R2889 VN.n21 VN.n20 56.5617
R2890 VN.n34 VN.n33 56.5617
R2891 VN.n77 VN.n76 56.5617
R2892 VN.n90 VN.n89 56.5617
R2893 VN.n14 VN.n13 56.1007
R2894 VN.n70 VN.n69 56.1007
R2895 VN.n47 VN.n46 44.4521
R2896 VN.n103 VN.n102 44.4521
R2897 VN.n47 VN.n2 36.702
R2898 VN.n103 VN.n58 36.702
R2899 VN.n15 VN.n12 24.5923
R2900 VN.n19 VN.n12 24.5923
R2901 VN.n20 VN.n19 24.5923
R2902 VN.n21 VN.n10 24.5923
R2903 VN.n25 VN.n10 24.5923
R2904 VN.n26 VN.n25 24.5923
R2905 VN.n28 VN.n8 24.5923
R2906 VN.n32 VN.n8 24.5923
R2907 VN.n33 VN.n32 24.5923
R2908 VN.n34 VN.n6 24.5923
R2909 VN.n38 VN.n6 24.5923
R2910 VN.n39 VN.n38 24.5923
R2911 VN.n41 VN.n4 24.5923
R2912 VN.n45 VN.n4 24.5923
R2913 VN.n46 VN.n45 24.5923
R2914 VN.n51 VN.n2 24.5923
R2915 VN.n52 VN.n51 24.5923
R2916 VN.n53 VN.n52 24.5923
R2917 VN.n76 VN.n75 24.5923
R2918 VN.n75 VN.n68 24.5923
R2919 VN.n71 VN.n68 24.5923
R2920 VN.n89 VN.n88 24.5923
R2921 VN.n88 VN.n64 24.5923
R2922 VN.n84 VN.n64 24.5923
R2923 VN.n82 VN.n81 24.5923
R2924 VN.n81 VN.n66 24.5923
R2925 VN.n77 VN.n66 24.5923
R2926 VN.n102 VN.n101 24.5923
R2927 VN.n101 VN.n60 24.5923
R2928 VN.n97 VN.n60 24.5923
R2929 VN.n95 VN.n94 24.5923
R2930 VN.n94 VN.n62 24.5923
R2931 VN.n90 VN.n62 24.5923
R2932 VN.n109 VN.n108 24.5923
R2933 VN.n108 VN.n107 24.5923
R2934 VN.n107 VN.n58 24.5923
R2935 VN.n15 VN.n14 19.1821
R2936 VN.n40 VN.n39 19.1821
R2937 VN.n71 VN.n70 19.1821
R2938 VN.n96 VN.n95 19.1821
R2939 VN.n27 VN.n26 12.2964
R2940 VN.n28 VN.n27 12.2964
R2941 VN.n84 VN.n83 12.2964
R2942 VN.n83 VN.n82 12.2964
R2943 VN.n41 VN.n40 5.4107
R2944 VN.n97 VN.n96 5.4107
R2945 VN.n16 VN.n13 2.48417
R2946 VN.n72 VN.n69 2.48417
R2947 VN.n53 VN.n0 1.47601
R2948 VN.n109 VN.n56 1.47601
R2949 VN.n111 VN.n110 0.354861
R2950 VN.n55 VN.n54 0.354861
R2951 VN VN.n55 0.267071
R2952 VN.n110 VN.n57 0.189894
R2953 VN.n106 VN.n57 0.189894
R2954 VN.n106 VN.n105 0.189894
R2955 VN.n105 VN.n104 0.189894
R2956 VN.n104 VN.n59 0.189894
R2957 VN.n100 VN.n59 0.189894
R2958 VN.n100 VN.n99 0.189894
R2959 VN.n99 VN.n98 0.189894
R2960 VN.n98 VN.n61 0.189894
R2961 VN.n93 VN.n61 0.189894
R2962 VN.n93 VN.n92 0.189894
R2963 VN.n92 VN.n91 0.189894
R2964 VN.n91 VN.n63 0.189894
R2965 VN.n87 VN.n63 0.189894
R2966 VN.n87 VN.n86 0.189894
R2967 VN.n86 VN.n85 0.189894
R2968 VN.n85 VN.n65 0.189894
R2969 VN.n80 VN.n65 0.189894
R2970 VN.n80 VN.n79 0.189894
R2971 VN.n79 VN.n78 0.189894
R2972 VN.n78 VN.n67 0.189894
R2973 VN.n74 VN.n67 0.189894
R2974 VN.n74 VN.n73 0.189894
R2975 VN.n73 VN.n72 0.189894
R2976 VN.n17 VN.n16 0.189894
R2977 VN.n18 VN.n17 0.189894
R2978 VN.n18 VN.n11 0.189894
R2979 VN.n22 VN.n11 0.189894
R2980 VN.n23 VN.n22 0.189894
R2981 VN.n24 VN.n23 0.189894
R2982 VN.n24 VN.n9 0.189894
R2983 VN.n29 VN.n9 0.189894
R2984 VN.n30 VN.n29 0.189894
R2985 VN.n31 VN.n30 0.189894
R2986 VN.n31 VN.n7 0.189894
R2987 VN.n35 VN.n7 0.189894
R2988 VN.n36 VN.n35 0.189894
R2989 VN.n37 VN.n36 0.189894
R2990 VN.n37 VN.n5 0.189894
R2991 VN.n42 VN.n5 0.189894
R2992 VN.n43 VN.n42 0.189894
R2993 VN.n44 VN.n43 0.189894
R2994 VN.n44 VN.n3 0.189894
R2995 VN.n48 VN.n3 0.189894
R2996 VN.n49 VN.n48 0.189894
R2997 VN.n50 VN.n49 0.189894
R2998 VN.n50 VN.n1 0.189894
R2999 VN.n54 VN.n1 0.189894
R3000 VDD2.n97 VDD2.n53 289.615
R3001 VDD2.n44 VDD2.n0 289.615
R3002 VDD2.n98 VDD2.n97 185
R3003 VDD2.n96 VDD2.n95 185
R3004 VDD2.n57 VDD2.n56 185
R3005 VDD2.n61 VDD2.n59 185
R3006 VDD2.n90 VDD2.n89 185
R3007 VDD2.n88 VDD2.n87 185
R3008 VDD2.n63 VDD2.n62 185
R3009 VDD2.n82 VDD2.n81 185
R3010 VDD2.n80 VDD2.n79 185
R3011 VDD2.n67 VDD2.n66 185
R3012 VDD2.n74 VDD2.n73 185
R3013 VDD2.n72 VDD2.n71 185
R3014 VDD2.n17 VDD2.n16 185
R3015 VDD2.n19 VDD2.n18 185
R3016 VDD2.n12 VDD2.n11 185
R3017 VDD2.n25 VDD2.n24 185
R3018 VDD2.n27 VDD2.n26 185
R3019 VDD2.n8 VDD2.n7 185
R3020 VDD2.n34 VDD2.n33 185
R3021 VDD2.n35 VDD2.n6 185
R3022 VDD2.n37 VDD2.n36 185
R3023 VDD2.n4 VDD2.n3 185
R3024 VDD2.n43 VDD2.n42 185
R3025 VDD2.n45 VDD2.n44 185
R3026 VDD2.n70 VDD2.t4 149.524
R3027 VDD2.n15 VDD2.t0 149.524
R3028 VDD2.n97 VDD2.n96 104.615
R3029 VDD2.n96 VDD2.n56 104.615
R3030 VDD2.n61 VDD2.n56 104.615
R3031 VDD2.n89 VDD2.n61 104.615
R3032 VDD2.n89 VDD2.n88 104.615
R3033 VDD2.n88 VDD2.n62 104.615
R3034 VDD2.n81 VDD2.n62 104.615
R3035 VDD2.n81 VDD2.n80 104.615
R3036 VDD2.n80 VDD2.n66 104.615
R3037 VDD2.n73 VDD2.n66 104.615
R3038 VDD2.n73 VDD2.n72 104.615
R3039 VDD2.n18 VDD2.n17 104.615
R3040 VDD2.n18 VDD2.n11 104.615
R3041 VDD2.n25 VDD2.n11 104.615
R3042 VDD2.n26 VDD2.n25 104.615
R3043 VDD2.n26 VDD2.n7 104.615
R3044 VDD2.n34 VDD2.n7 104.615
R3045 VDD2.n35 VDD2.n34 104.615
R3046 VDD2.n36 VDD2.n35 104.615
R3047 VDD2.n36 VDD2.n3 104.615
R3048 VDD2.n43 VDD2.n3 104.615
R3049 VDD2.n44 VDD2.n43 104.615
R3050 VDD2.n52 VDD2.n51 67.9505
R3051 VDD2 VDD2.n105 67.9477
R3052 VDD2.n104 VDD2.n103 65.3293
R3053 VDD2.n50 VDD2.n49 65.3292
R3054 VDD2.n50 VDD2.n48 54.7604
R3055 VDD2.n72 VDD2.t4 52.3082
R3056 VDD2.n17 VDD2.t0 52.3082
R3057 VDD2.n102 VDD2.n101 51.1914
R3058 VDD2.n102 VDD2.n52 48.7368
R3059 VDD2.n59 VDD2.n57 13.1884
R3060 VDD2.n37 VDD2.n4 13.1884
R3061 VDD2.n95 VDD2.n94 12.8005
R3062 VDD2.n91 VDD2.n90 12.8005
R3063 VDD2.n38 VDD2.n6 12.8005
R3064 VDD2.n42 VDD2.n41 12.8005
R3065 VDD2.n98 VDD2.n55 12.0247
R3066 VDD2.n87 VDD2.n60 12.0247
R3067 VDD2.n33 VDD2.n32 12.0247
R3068 VDD2.n45 VDD2.n2 12.0247
R3069 VDD2.n99 VDD2.n53 11.249
R3070 VDD2.n86 VDD2.n63 11.249
R3071 VDD2.n31 VDD2.n8 11.249
R3072 VDD2.n46 VDD2.n0 11.249
R3073 VDD2.n83 VDD2.n82 10.4732
R3074 VDD2.n28 VDD2.n27 10.4732
R3075 VDD2.n71 VDD2.n70 10.2747
R3076 VDD2.n16 VDD2.n15 10.2747
R3077 VDD2.n79 VDD2.n65 9.69747
R3078 VDD2.n24 VDD2.n10 9.69747
R3079 VDD2.n101 VDD2.n100 9.45567
R3080 VDD2.n48 VDD2.n47 9.45567
R3081 VDD2.n69 VDD2.n68 9.3005
R3082 VDD2.n76 VDD2.n75 9.3005
R3083 VDD2.n78 VDD2.n77 9.3005
R3084 VDD2.n65 VDD2.n64 9.3005
R3085 VDD2.n84 VDD2.n83 9.3005
R3086 VDD2.n86 VDD2.n85 9.3005
R3087 VDD2.n60 VDD2.n58 9.3005
R3088 VDD2.n92 VDD2.n91 9.3005
R3089 VDD2.n100 VDD2.n99 9.3005
R3090 VDD2.n55 VDD2.n54 9.3005
R3091 VDD2.n94 VDD2.n93 9.3005
R3092 VDD2.n47 VDD2.n46 9.3005
R3093 VDD2.n2 VDD2.n1 9.3005
R3094 VDD2.n41 VDD2.n40 9.3005
R3095 VDD2.n14 VDD2.n13 9.3005
R3096 VDD2.n21 VDD2.n20 9.3005
R3097 VDD2.n23 VDD2.n22 9.3005
R3098 VDD2.n10 VDD2.n9 9.3005
R3099 VDD2.n29 VDD2.n28 9.3005
R3100 VDD2.n31 VDD2.n30 9.3005
R3101 VDD2.n32 VDD2.n5 9.3005
R3102 VDD2.n39 VDD2.n38 9.3005
R3103 VDD2.n78 VDD2.n67 8.92171
R3104 VDD2.n23 VDD2.n12 8.92171
R3105 VDD2.n75 VDD2.n74 8.14595
R3106 VDD2.n20 VDD2.n19 8.14595
R3107 VDD2.n71 VDD2.n69 7.3702
R3108 VDD2.n16 VDD2.n14 7.3702
R3109 VDD2.n74 VDD2.n69 5.81868
R3110 VDD2.n19 VDD2.n14 5.81868
R3111 VDD2.n75 VDD2.n67 5.04292
R3112 VDD2.n20 VDD2.n12 5.04292
R3113 VDD2.n79 VDD2.n78 4.26717
R3114 VDD2.n24 VDD2.n23 4.26717
R3115 VDD2.n104 VDD2.n102 3.56947
R3116 VDD2.n82 VDD2.n65 3.49141
R3117 VDD2.n27 VDD2.n10 3.49141
R3118 VDD2.n70 VDD2.n68 2.84303
R3119 VDD2.n15 VDD2.n13 2.84303
R3120 VDD2.n101 VDD2.n53 2.71565
R3121 VDD2.n83 VDD2.n63 2.71565
R3122 VDD2.n28 VDD2.n8 2.71565
R3123 VDD2.n48 VDD2.n0 2.71565
R3124 VDD2.n105 VDD2.t8 2.11588
R3125 VDD2.n105 VDD2.t3 2.11588
R3126 VDD2.n103 VDD2.t7 2.11588
R3127 VDD2.n103 VDD2.t2 2.11588
R3128 VDD2.n51 VDD2.t6 2.11588
R3129 VDD2.n51 VDD2.t1 2.11588
R3130 VDD2.n49 VDD2.t9 2.11588
R3131 VDD2.n49 VDD2.t5 2.11588
R3132 VDD2.n99 VDD2.n98 1.93989
R3133 VDD2.n87 VDD2.n86 1.93989
R3134 VDD2.n33 VDD2.n31 1.93989
R3135 VDD2.n46 VDD2.n45 1.93989
R3136 VDD2.n95 VDD2.n55 1.16414
R3137 VDD2.n90 VDD2.n60 1.16414
R3138 VDD2.n32 VDD2.n6 1.16414
R3139 VDD2.n42 VDD2.n2 1.16414
R3140 VDD2 VDD2.n104 0.950931
R3141 VDD2.n52 VDD2.n50 0.837395
R3142 VDD2.n94 VDD2.n57 0.388379
R3143 VDD2.n91 VDD2.n59 0.388379
R3144 VDD2.n38 VDD2.n37 0.388379
R3145 VDD2.n41 VDD2.n4 0.388379
R3146 VDD2.n100 VDD2.n54 0.155672
R3147 VDD2.n93 VDD2.n54 0.155672
R3148 VDD2.n93 VDD2.n92 0.155672
R3149 VDD2.n92 VDD2.n58 0.155672
R3150 VDD2.n85 VDD2.n58 0.155672
R3151 VDD2.n85 VDD2.n84 0.155672
R3152 VDD2.n84 VDD2.n64 0.155672
R3153 VDD2.n77 VDD2.n64 0.155672
R3154 VDD2.n77 VDD2.n76 0.155672
R3155 VDD2.n76 VDD2.n68 0.155672
R3156 VDD2.n21 VDD2.n13 0.155672
R3157 VDD2.n22 VDD2.n21 0.155672
R3158 VDD2.n22 VDD2.n9 0.155672
R3159 VDD2.n29 VDD2.n9 0.155672
R3160 VDD2.n30 VDD2.n29 0.155672
R3161 VDD2.n30 VDD2.n5 0.155672
R3162 VDD2.n39 VDD2.n5 0.155672
R3163 VDD2.n40 VDD2.n39 0.155672
R3164 VDD2.n40 VDD2.n1 0.155672
R3165 VDD2.n47 VDD2.n1 0.155672
C0 VDD1 VDD2 2.96221f
C1 VDD2 VP 0.73771f
C2 VN VDD1 0.15641f
C3 VN VP 9.686259f
C4 VTAIL VDD1 9.997691f
C5 VN VDD2 8.99606f
C6 VTAIL VP 10.2983f
C7 VTAIL VDD2 10.0581f
C8 VN VTAIL 10.2837f
C9 VDD1 VP 9.57408f
C10 VDD2 B 8.176821f
C11 VDD1 B 8.131026f
C12 VTAIL B 8.045068f
C13 VN B 23.73278f
C14 VP B 22.322727f
C15 VDD2.n0 B 0.035337f
C16 VDD2.n1 B 0.025632f
C17 VDD2.n2 B 0.013774f
C18 VDD2.n3 B 0.032556f
C19 VDD2.n4 B 0.014179f
C20 VDD2.n5 B 0.025632f
C21 VDD2.n6 B 0.014584f
C22 VDD2.n7 B 0.032556f
C23 VDD2.n8 B 0.014584f
C24 VDD2.n9 B 0.025632f
C25 VDD2.n10 B 0.013774f
C26 VDD2.n11 B 0.032556f
C27 VDD2.n12 B 0.014584f
C28 VDD2.n13 B 0.992113f
C29 VDD2.n14 B 0.013774f
C30 VDD2.t0 B 0.054625f
C31 VDD2.n15 B 0.158835f
C32 VDD2.n16 B 0.023015f
C33 VDD2.n17 B 0.024417f
C34 VDD2.n18 B 0.032556f
C35 VDD2.n19 B 0.014584f
C36 VDD2.n20 B 0.013774f
C37 VDD2.n21 B 0.025632f
C38 VDD2.n22 B 0.025632f
C39 VDD2.n23 B 0.013774f
C40 VDD2.n24 B 0.014584f
C41 VDD2.n25 B 0.032556f
C42 VDD2.n26 B 0.032556f
C43 VDD2.n27 B 0.014584f
C44 VDD2.n28 B 0.013774f
C45 VDD2.n29 B 0.025632f
C46 VDD2.n30 B 0.025632f
C47 VDD2.n31 B 0.013774f
C48 VDD2.n32 B 0.013774f
C49 VDD2.n33 B 0.014584f
C50 VDD2.n34 B 0.032556f
C51 VDD2.n35 B 0.032556f
C52 VDD2.n36 B 0.032556f
C53 VDD2.n37 B 0.014179f
C54 VDD2.n38 B 0.013774f
C55 VDD2.n39 B 0.025632f
C56 VDD2.n40 B 0.025632f
C57 VDD2.n41 B 0.013774f
C58 VDD2.n42 B 0.014584f
C59 VDD2.n43 B 0.032556f
C60 VDD2.n44 B 0.069255f
C61 VDD2.n45 B 0.014584f
C62 VDD2.n46 B 0.013774f
C63 VDD2.n47 B 0.06345f
C64 VDD2.n48 B 0.079004f
C65 VDD2.t9 B 0.189591f
C66 VDD2.t5 B 0.189591f
C67 VDD2.n49 B 1.66323f
C68 VDD2.n50 B 0.894543f
C69 VDD2.t6 B 0.189591f
C70 VDD2.t1 B 0.189591f
C71 VDD2.n51 B 1.6913f
C72 VDD2.n52 B 3.45214f
C73 VDD2.n53 B 0.035337f
C74 VDD2.n54 B 0.025632f
C75 VDD2.n55 B 0.013774f
C76 VDD2.n56 B 0.032556f
C77 VDD2.n57 B 0.014179f
C78 VDD2.n58 B 0.025632f
C79 VDD2.n59 B 0.014179f
C80 VDD2.n60 B 0.013774f
C81 VDD2.n61 B 0.032556f
C82 VDD2.n62 B 0.032556f
C83 VDD2.n63 B 0.014584f
C84 VDD2.n64 B 0.025632f
C85 VDD2.n65 B 0.013774f
C86 VDD2.n66 B 0.032556f
C87 VDD2.n67 B 0.014584f
C88 VDD2.n68 B 0.992113f
C89 VDD2.n69 B 0.013774f
C90 VDD2.t4 B 0.054625f
C91 VDD2.n70 B 0.158835f
C92 VDD2.n71 B 0.023015f
C93 VDD2.n72 B 0.024417f
C94 VDD2.n73 B 0.032556f
C95 VDD2.n74 B 0.014584f
C96 VDD2.n75 B 0.013774f
C97 VDD2.n76 B 0.025632f
C98 VDD2.n77 B 0.025632f
C99 VDD2.n78 B 0.013774f
C100 VDD2.n79 B 0.014584f
C101 VDD2.n80 B 0.032556f
C102 VDD2.n81 B 0.032556f
C103 VDD2.n82 B 0.014584f
C104 VDD2.n83 B 0.013774f
C105 VDD2.n84 B 0.025632f
C106 VDD2.n85 B 0.025632f
C107 VDD2.n86 B 0.013774f
C108 VDD2.n87 B 0.014584f
C109 VDD2.n88 B 0.032556f
C110 VDD2.n89 B 0.032556f
C111 VDD2.n90 B 0.014584f
C112 VDD2.n91 B 0.013774f
C113 VDD2.n92 B 0.025632f
C114 VDD2.n93 B 0.025632f
C115 VDD2.n94 B 0.013774f
C116 VDD2.n95 B 0.014584f
C117 VDD2.n96 B 0.032556f
C118 VDD2.n97 B 0.069255f
C119 VDD2.n98 B 0.014584f
C120 VDD2.n99 B 0.013774f
C121 VDD2.n100 B 0.06345f
C122 VDD2.n101 B 0.056418f
C123 VDD2.n102 B 3.24194f
C124 VDD2.t7 B 0.189591f
C125 VDD2.t2 B 0.189591f
C126 VDD2.n103 B 1.66323f
C127 VDD2.n104 B 0.579252f
C128 VDD2.t8 B 0.189591f
C129 VDD2.t3 B 0.189591f
C130 VDD2.n105 B 1.69126f
C131 VN.t8 B 1.6892f
C132 VN.n0 B 0.6641f
C133 VN.n1 B 0.017526f
C134 VN.n2 B 0.035148f
C135 VN.n3 B 0.017526f
C136 VN.n4 B 0.032501f
C137 VN.n5 B 0.017526f
C138 VN.t3 B 1.6892f
C139 VN.n6 B 0.032501f
C140 VN.n7 B 0.017526f
C141 VN.n8 B 0.032501f
C142 VN.n9 B 0.017526f
C143 VN.t4 B 1.6892f
C144 VN.n10 B 0.032501f
C145 VN.n11 B 0.017526f
C146 VN.n12 B 0.032501f
C147 VN.t9 B 1.95134f
C148 VN.n13 B 0.635713f
C149 VN.t0 B 1.6892f
C150 VN.n14 B 0.667285f
C151 VN.n15 B 0.028971f
C152 VN.n16 B 0.22579f
C153 VN.n17 B 0.017526f
C154 VN.n18 B 0.017526f
C155 VN.n19 B 0.032501f
C156 VN.n20 B 0.022083f
C157 VN.n21 B 0.028871f
C158 VN.n22 B 0.017526f
C159 VN.n23 B 0.017526f
C160 VN.n24 B 0.017526f
C161 VN.n25 B 0.032501f
C162 VN.n26 B 0.024478f
C163 VN.n27 B 0.599904f
C164 VN.n28 B 0.024478f
C165 VN.n29 B 0.017526f
C166 VN.n30 B 0.017526f
C167 VN.n31 B 0.017526f
C168 VN.n32 B 0.032501f
C169 VN.n33 B 0.028871f
C170 VN.n34 B 0.022083f
C171 VN.n35 B 0.017526f
C172 VN.n36 B 0.017526f
C173 VN.n37 B 0.017526f
C174 VN.n38 B 0.032501f
C175 VN.n39 B 0.028971f
C176 VN.n40 B 0.599904f
C177 VN.n41 B 0.019986f
C178 VN.n42 B 0.017526f
C179 VN.n43 B 0.017526f
C180 VN.n44 B 0.017526f
C181 VN.n45 B 0.032501f
C182 VN.n46 B 0.033791f
C183 VN.n47 B 0.014516f
C184 VN.n48 B 0.017526f
C185 VN.n49 B 0.017526f
C186 VN.n50 B 0.017526f
C187 VN.n51 B 0.032501f
C188 VN.n52 B 0.032501f
C189 VN.n53 B 0.017419f
C190 VN.n54 B 0.028282f
C191 VN.n55 B 0.054576f
C192 VN.t5 B 1.6892f
C193 VN.n56 B 0.6641f
C194 VN.n57 B 0.017526f
C195 VN.n58 B 0.035148f
C196 VN.n59 B 0.017526f
C197 VN.n60 B 0.032501f
C198 VN.n61 B 0.017526f
C199 VN.t2 B 1.6892f
C200 VN.n62 B 0.032501f
C201 VN.n63 B 0.017526f
C202 VN.n64 B 0.032501f
C203 VN.n65 B 0.017526f
C204 VN.t7 B 1.6892f
C205 VN.n66 B 0.032501f
C206 VN.n67 B 0.017526f
C207 VN.n68 B 0.032501f
C208 VN.t6 B 1.95134f
C209 VN.n69 B 0.635713f
C210 VN.t1 B 1.6892f
C211 VN.n70 B 0.667285f
C212 VN.n71 B 0.028971f
C213 VN.n72 B 0.225789f
C214 VN.n73 B 0.017526f
C215 VN.n74 B 0.017526f
C216 VN.n75 B 0.032501f
C217 VN.n76 B 0.022083f
C218 VN.n77 B 0.028871f
C219 VN.n78 B 0.017526f
C220 VN.n79 B 0.017526f
C221 VN.n80 B 0.017526f
C222 VN.n81 B 0.032501f
C223 VN.n82 B 0.024478f
C224 VN.n83 B 0.599904f
C225 VN.n84 B 0.024478f
C226 VN.n85 B 0.017526f
C227 VN.n86 B 0.017526f
C228 VN.n87 B 0.017526f
C229 VN.n88 B 0.032501f
C230 VN.n89 B 0.028871f
C231 VN.n90 B 0.022083f
C232 VN.n91 B 0.017526f
C233 VN.n92 B 0.017526f
C234 VN.n93 B 0.017526f
C235 VN.n94 B 0.032501f
C236 VN.n95 B 0.028971f
C237 VN.n96 B 0.599904f
C238 VN.n97 B 0.019986f
C239 VN.n98 B 0.017526f
C240 VN.n99 B 0.017526f
C241 VN.n100 B 0.017526f
C242 VN.n101 B 0.032501f
C243 VN.n102 B 0.033791f
C244 VN.n103 B 0.014516f
C245 VN.n104 B 0.017526f
C246 VN.n105 B 0.017526f
C247 VN.n106 B 0.017526f
C248 VN.n107 B 0.032501f
C249 VN.n108 B 0.032501f
C250 VN.n109 B 0.017419f
C251 VN.n110 B 0.028282f
C252 VN.n111 B 1.23715f
C253 VDD1.n0 B 0.035982f
C254 VDD1.n1 B 0.0261f
C255 VDD1.n2 B 0.014025f
C256 VDD1.n3 B 0.033151f
C257 VDD1.n4 B 0.014438f
C258 VDD1.n5 B 0.0261f
C259 VDD1.n6 B 0.014438f
C260 VDD1.n7 B 0.014025f
C261 VDD1.n8 B 0.033151f
C262 VDD1.n9 B 0.033151f
C263 VDD1.n10 B 0.01485f
C264 VDD1.n11 B 0.0261f
C265 VDD1.n12 B 0.014025f
C266 VDD1.n13 B 0.033151f
C267 VDD1.n14 B 0.01485f
C268 VDD1.n15 B 1.01023f
C269 VDD1.n16 B 0.014025f
C270 VDD1.t4 B 0.055623f
C271 VDD1.n17 B 0.161736f
C272 VDD1.n18 B 0.023435f
C273 VDD1.n19 B 0.024863f
C274 VDD1.n20 B 0.033151f
C275 VDD1.n21 B 0.01485f
C276 VDD1.n22 B 0.014025f
C277 VDD1.n23 B 0.0261f
C278 VDD1.n24 B 0.0261f
C279 VDD1.n25 B 0.014025f
C280 VDD1.n26 B 0.01485f
C281 VDD1.n27 B 0.033151f
C282 VDD1.n28 B 0.033151f
C283 VDD1.n29 B 0.01485f
C284 VDD1.n30 B 0.014025f
C285 VDD1.n31 B 0.0261f
C286 VDD1.n32 B 0.0261f
C287 VDD1.n33 B 0.014025f
C288 VDD1.n34 B 0.01485f
C289 VDD1.n35 B 0.033151f
C290 VDD1.n36 B 0.033151f
C291 VDD1.n37 B 0.01485f
C292 VDD1.n38 B 0.014025f
C293 VDD1.n39 B 0.0261f
C294 VDD1.n40 B 0.0261f
C295 VDD1.n41 B 0.014025f
C296 VDD1.n42 B 0.01485f
C297 VDD1.n43 B 0.033151f
C298 VDD1.n44 B 0.07052f
C299 VDD1.n45 B 0.01485f
C300 VDD1.n46 B 0.014025f
C301 VDD1.n47 B 0.064609f
C302 VDD1.n48 B 0.080447f
C303 VDD1.t0 B 0.193054f
C304 VDD1.t7 B 0.193054f
C305 VDD1.n49 B 1.69361f
C306 VDD1.n50 B 0.919697f
C307 VDD1.n51 B 0.035982f
C308 VDD1.n52 B 0.0261f
C309 VDD1.n53 B 0.014025f
C310 VDD1.n54 B 0.033151f
C311 VDD1.n55 B 0.014438f
C312 VDD1.n56 B 0.0261f
C313 VDD1.n57 B 0.01485f
C314 VDD1.n58 B 0.033151f
C315 VDD1.n59 B 0.01485f
C316 VDD1.n60 B 0.0261f
C317 VDD1.n61 B 0.014025f
C318 VDD1.n62 B 0.033151f
C319 VDD1.n63 B 0.01485f
C320 VDD1.n64 B 1.01023f
C321 VDD1.n65 B 0.014025f
C322 VDD1.t2 B 0.055623f
C323 VDD1.n66 B 0.161736f
C324 VDD1.n67 B 0.023435f
C325 VDD1.n68 B 0.024863f
C326 VDD1.n69 B 0.033151f
C327 VDD1.n70 B 0.01485f
C328 VDD1.n71 B 0.014025f
C329 VDD1.n72 B 0.0261f
C330 VDD1.n73 B 0.0261f
C331 VDD1.n74 B 0.014025f
C332 VDD1.n75 B 0.01485f
C333 VDD1.n76 B 0.033151f
C334 VDD1.n77 B 0.033151f
C335 VDD1.n78 B 0.01485f
C336 VDD1.n79 B 0.014025f
C337 VDD1.n80 B 0.0261f
C338 VDD1.n81 B 0.0261f
C339 VDD1.n82 B 0.014025f
C340 VDD1.n83 B 0.014025f
C341 VDD1.n84 B 0.01485f
C342 VDD1.n85 B 0.033151f
C343 VDD1.n86 B 0.033151f
C344 VDD1.n87 B 0.033151f
C345 VDD1.n88 B 0.014438f
C346 VDD1.n89 B 0.014025f
C347 VDD1.n90 B 0.0261f
C348 VDD1.n91 B 0.0261f
C349 VDD1.n92 B 0.014025f
C350 VDD1.n93 B 0.01485f
C351 VDD1.n94 B 0.033151f
C352 VDD1.n95 B 0.07052f
C353 VDD1.n96 B 0.01485f
C354 VDD1.n97 B 0.014025f
C355 VDD1.n98 B 0.064609f
C356 VDD1.n99 B 0.080447f
C357 VDD1.t3 B 0.193054f
C358 VDD1.t6 B 0.193054f
C359 VDD1.n100 B 1.6936f
C360 VDD1.n101 B 0.910879f
C361 VDD1.t8 B 0.193054f
C362 VDD1.t9 B 0.193054f
C363 VDD1.n102 B 1.72219f
C364 VDD1.n103 B 3.67828f
C365 VDD1.t5 B 0.193054f
C366 VDD1.t1 B 0.193054f
C367 VDD1.n104 B 1.6936f
C368 VDD1.n105 B 3.62223f
C369 VTAIL.t4 B 0.200934f
C370 VTAIL.t5 B 0.200934f
C371 VTAIL.n0 B 1.68966f
C372 VTAIL.n1 B 0.691188f
C373 VTAIL.n2 B 0.037451f
C374 VTAIL.n3 B 0.027166f
C375 VTAIL.n4 B 0.014598f
C376 VTAIL.n5 B 0.034504f
C377 VTAIL.n6 B 0.015027f
C378 VTAIL.n7 B 0.027166f
C379 VTAIL.n8 B 0.015457f
C380 VTAIL.n9 B 0.034504f
C381 VTAIL.n10 B 0.015457f
C382 VTAIL.n11 B 0.027166f
C383 VTAIL.n12 B 0.014598f
C384 VTAIL.n13 B 0.034504f
C385 VTAIL.n14 B 0.015457f
C386 VTAIL.n15 B 1.05147f
C387 VTAIL.n16 B 0.014598f
C388 VTAIL.t13 B 0.057893f
C389 VTAIL.n17 B 0.168338f
C390 VTAIL.n18 B 0.024392f
C391 VTAIL.n19 B 0.025878f
C392 VTAIL.n20 B 0.034504f
C393 VTAIL.n21 B 0.015457f
C394 VTAIL.n22 B 0.014598f
C395 VTAIL.n23 B 0.027166f
C396 VTAIL.n24 B 0.027166f
C397 VTAIL.n25 B 0.014598f
C398 VTAIL.n26 B 0.015457f
C399 VTAIL.n27 B 0.034504f
C400 VTAIL.n28 B 0.034504f
C401 VTAIL.n29 B 0.015457f
C402 VTAIL.n30 B 0.014598f
C403 VTAIL.n31 B 0.027166f
C404 VTAIL.n32 B 0.027166f
C405 VTAIL.n33 B 0.014598f
C406 VTAIL.n34 B 0.014598f
C407 VTAIL.n35 B 0.015457f
C408 VTAIL.n36 B 0.034504f
C409 VTAIL.n37 B 0.034504f
C410 VTAIL.n38 B 0.034504f
C411 VTAIL.n39 B 0.015027f
C412 VTAIL.n40 B 0.014598f
C413 VTAIL.n41 B 0.027166f
C414 VTAIL.n42 B 0.027166f
C415 VTAIL.n43 B 0.014598f
C416 VTAIL.n44 B 0.015457f
C417 VTAIL.n45 B 0.034504f
C418 VTAIL.n46 B 0.073399f
C419 VTAIL.n47 B 0.015457f
C420 VTAIL.n48 B 0.014598f
C421 VTAIL.n49 B 0.067246f
C422 VTAIL.n50 B 0.041069f
C423 VTAIL.n51 B 0.535458f
C424 VTAIL.t18 B 0.200934f
C425 VTAIL.t12 B 0.200934f
C426 VTAIL.n52 B 1.68966f
C427 VTAIL.n53 B 0.879274f
C428 VTAIL.t16 B 0.200934f
C429 VTAIL.t19 B 0.200934f
C430 VTAIL.n54 B 1.68966f
C431 VTAIL.n55 B 2.26701f
C432 VTAIL.t8 B 0.200934f
C433 VTAIL.t2 B 0.200934f
C434 VTAIL.n56 B 1.68967f
C435 VTAIL.n57 B 2.267f
C436 VTAIL.t7 B 0.200934f
C437 VTAIL.t6 B 0.200934f
C438 VTAIL.n58 B 1.68967f
C439 VTAIL.n59 B 0.879264f
C440 VTAIL.n60 B 0.037451f
C441 VTAIL.n61 B 0.027166f
C442 VTAIL.n62 B 0.014598f
C443 VTAIL.n63 B 0.034504f
C444 VTAIL.n64 B 0.015027f
C445 VTAIL.n65 B 0.027166f
C446 VTAIL.n66 B 0.015027f
C447 VTAIL.n67 B 0.014598f
C448 VTAIL.n68 B 0.034504f
C449 VTAIL.n69 B 0.034504f
C450 VTAIL.n70 B 0.015457f
C451 VTAIL.n71 B 0.027166f
C452 VTAIL.n72 B 0.014598f
C453 VTAIL.n73 B 0.034504f
C454 VTAIL.n74 B 0.015457f
C455 VTAIL.n75 B 1.05147f
C456 VTAIL.n76 B 0.014598f
C457 VTAIL.t0 B 0.057893f
C458 VTAIL.n77 B 0.168338f
C459 VTAIL.n78 B 0.024392f
C460 VTAIL.n79 B 0.025878f
C461 VTAIL.n80 B 0.034504f
C462 VTAIL.n81 B 0.015457f
C463 VTAIL.n82 B 0.014598f
C464 VTAIL.n83 B 0.027166f
C465 VTAIL.n84 B 0.027166f
C466 VTAIL.n85 B 0.014598f
C467 VTAIL.n86 B 0.015457f
C468 VTAIL.n87 B 0.034504f
C469 VTAIL.n88 B 0.034504f
C470 VTAIL.n89 B 0.015457f
C471 VTAIL.n90 B 0.014598f
C472 VTAIL.n91 B 0.027166f
C473 VTAIL.n92 B 0.027166f
C474 VTAIL.n93 B 0.014598f
C475 VTAIL.n94 B 0.015457f
C476 VTAIL.n95 B 0.034504f
C477 VTAIL.n96 B 0.034504f
C478 VTAIL.n97 B 0.015457f
C479 VTAIL.n98 B 0.014598f
C480 VTAIL.n99 B 0.027166f
C481 VTAIL.n100 B 0.027166f
C482 VTAIL.n101 B 0.014598f
C483 VTAIL.n102 B 0.015457f
C484 VTAIL.n103 B 0.034504f
C485 VTAIL.n104 B 0.073399f
C486 VTAIL.n105 B 0.015457f
C487 VTAIL.n106 B 0.014598f
C488 VTAIL.n107 B 0.067246f
C489 VTAIL.n108 B 0.041069f
C490 VTAIL.n109 B 0.535458f
C491 VTAIL.t17 B 0.200934f
C492 VTAIL.t10 B 0.200934f
C493 VTAIL.n110 B 1.68967f
C494 VTAIL.n111 B 0.764186f
C495 VTAIL.t14 B 0.200934f
C496 VTAIL.t15 B 0.200934f
C497 VTAIL.n112 B 1.68967f
C498 VTAIL.n113 B 0.879264f
C499 VTAIL.n114 B 0.037451f
C500 VTAIL.n115 B 0.027166f
C501 VTAIL.n116 B 0.014598f
C502 VTAIL.n117 B 0.034504f
C503 VTAIL.n118 B 0.015027f
C504 VTAIL.n119 B 0.027166f
C505 VTAIL.n120 B 0.015027f
C506 VTAIL.n121 B 0.014598f
C507 VTAIL.n122 B 0.034504f
C508 VTAIL.n123 B 0.034504f
C509 VTAIL.n124 B 0.015457f
C510 VTAIL.n125 B 0.027166f
C511 VTAIL.n126 B 0.014598f
C512 VTAIL.n127 B 0.034504f
C513 VTAIL.n128 B 0.015457f
C514 VTAIL.n129 B 1.05147f
C515 VTAIL.n130 B 0.014598f
C516 VTAIL.t11 B 0.057893f
C517 VTAIL.n131 B 0.168338f
C518 VTAIL.n132 B 0.024392f
C519 VTAIL.n133 B 0.025878f
C520 VTAIL.n134 B 0.034504f
C521 VTAIL.n135 B 0.015457f
C522 VTAIL.n136 B 0.014598f
C523 VTAIL.n137 B 0.027166f
C524 VTAIL.n138 B 0.027166f
C525 VTAIL.n139 B 0.014598f
C526 VTAIL.n140 B 0.015457f
C527 VTAIL.n141 B 0.034504f
C528 VTAIL.n142 B 0.034504f
C529 VTAIL.n143 B 0.015457f
C530 VTAIL.n144 B 0.014598f
C531 VTAIL.n145 B 0.027166f
C532 VTAIL.n146 B 0.027166f
C533 VTAIL.n147 B 0.014598f
C534 VTAIL.n148 B 0.015457f
C535 VTAIL.n149 B 0.034504f
C536 VTAIL.n150 B 0.034504f
C537 VTAIL.n151 B 0.015457f
C538 VTAIL.n152 B 0.014598f
C539 VTAIL.n153 B 0.027166f
C540 VTAIL.n154 B 0.027166f
C541 VTAIL.n155 B 0.014598f
C542 VTAIL.n156 B 0.015457f
C543 VTAIL.n157 B 0.034504f
C544 VTAIL.n158 B 0.073399f
C545 VTAIL.n159 B 0.015457f
C546 VTAIL.n160 B 0.014598f
C547 VTAIL.n161 B 0.067246f
C548 VTAIL.n162 B 0.041069f
C549 VTAIL.n163 B 1.72587f
C550 VTAIL.n164 B 0.037451f
C551 VTAIL.n165 B 0.027166f
C552 VTAIL.n166 B 0.014598f
C553 VTAIL.n167 B 0.034504f
C554 VTAIL.n168 B 0.015027f
C555 VTAIL.n169 B 0.027166f
C556 VTAIL.n170 B 0.015457f
C557 VTAIL.n171 B 0.034504f
C558 VTAIL.n172 B 0.015457f
C559 VTAIL.n173 B 0.027166f
C560 VTAIL.n174 B 0.014598f
C561 VTAIL.n175 B 0.034504f
C562 VTAIL.n176 B 0.015457f
C563 VTAIL.n177 B 1.05147f
C564 VTAIL.n178 B 0.014598f
C565 VTAIL.t9 B 0.057893f
C566 VTAIL.n179 B 0.168338f
C567 VTAIL.n180 B 0.024392f
C568 VTAIL.n181 B 0.025878f
C569 VTAIL.n182 B 0.034504f
C570 VTAIL.n183 B 0.015457f
C571 VTAIL.n184 B 0.014598f
C572 VTAIL.n185 B 0.027166f
C573 VTAIL.n186 B 0.027166f
C574 VTAIL.n187 B 0.014598f
C575 VTAIL.n188 B 0.015457f
C576 VTAIL.n189 B 0.034504f
C577 VTAIL.n190 B 0.034504f
C578 VTAIL.n191 B 0.015457f
C579 VTAIL.n192 B 0.014598f
C580 VTAIL.n193 B 0.027166f
C581 VTAIL.n194 B 0.027166f
C582 VTAIL.n195 B 0.014598f
C583 VTAIL.n196 B 0.014598f
C584 VTAIL.n197 B 0.015457f
C585 VTAIL.n198 B 0.034504f
C586 VTAIL.n199 B 0.034504f
C587 VTAIL.n200 B 0.034504f
C588 VTAIL.n201 B 0.015027f
C589 VTAIL.n202 B 0.014598f
C590 VTAIL.n203 B 0.027166f
C591 VTAIL.n204 B 0.027166f
C592 VTAIL.n205 B 0.014598f
C593 VTAIL.n206 B 0.015457f
C594 VTAIL.n207 B 0.034504f
C595 VTAIL.n208 B 0.073399f
C596 VTAIL.n209 B 0.015457f
C597 VTAIL.n210 B 0.014598f
C598 VTAIL.n211 B 0.067246f
C599 VTAIL.n212 B 0.041069f
C600 VTAIL.n213 B 1.72587f
C601 VTAIL.t1 B 0.200934f
C602 VTAIL.t3 B 0.200934f
C603 VTAIL.n214 B 1.68966f
C604 VTAIL.n215 B 0.639874f
C605 VP.t0 B 1.72562f
C606 VP.n0 B 0.678416f
C607 VP.n1 B 0.017904f
C608 VP.n2 B 0.035905f
C609 VP.n3 B 0.017904f
C610 VP.n4 B 0.033201f
C611 VP.n5 B 0.017904f
C612 VP.t1 B 1.72562f
C613 VP.n6 B 0.033201f
C614 VP.n7 B 0.017904f
C615 VP.n8 B 0.033201f
C616 VP.n9 B 0.017904f
C617 VP.t3 B 1.72562f
C618 VP.n10 B 0.033201f
C619 VP.n11 B 0.017904f
C620 VP.n12 B 0.033201f
C621 VP.n13 B 0.017904f
C622 VP.t6 B 1.72562f
C623 VP.n14 B 0.033201f
C624 VP.n15 B 0.017904f
C625 VP.n16 B 0.033201f
C626 VP.n17 B 0.028892f
C627 VP.t7 B 1.72562f
C628 VP.t8 B 1.72562f
C629 VP.n18 B 0.678416f
C630 VP.n19 B 0.017904f
C631 VP.n20 B 0.035905f
C632 VP.n21 B 0.017904f
C633 VP.n22 B 0.033201f
C634 VP.n23 B 0.017904f
C635 VP.t4 B 1.72562f
C636 VP.n24 B 0.033201f
C637 VP.n25 B 0.017904f
C638 VP.n26 B 0.033201f
C639 VP.n27 B 0.017904f
C640 VP.t2 B 1.72562f
C641 VP.n28 B 0.033201f
C642 VP.n29 B 0.017904f
C643 VP.n30 B 0.033201f
C644 VP.t5 B 1.9934f
C645 VP.n31 B 0.649418f
C646 VP.t9 B 1.72562f
C647 VP.n32 B 0.68167f
C648 VP.n33 B 0.029595f
C649 VP.n34 B 0.230657f
C650 VP.n35 B 0.017904f
C651 VP.n36 B 0.017904f
C652 VP.n37 B 0.033201f
C653 VP.n38 B 0.022559f
C654 VP.n39 B 0.029494f
C655 VP.n40 B 0.017904f
C656 VP.n41 B 0.017904f
C657 VP.n42 B 0.017904f
C658 VP.n43 B 0.033201f
C659 VP.n44 B 0.025006f
C660 VP.n45 B 0.612837f
C661 VP.n46 B 0.025006f
C662 VP.n47 B 0.017904f
C663 VP.n48 B 0.017904f
C664 VP.n49 B 0.017904f
C665 VP.n50 B 0.033201f
C666 VP.n51 B 0.029494f
C667 VP.n52 B 0.022559f
C668 VP.n53 B 0.017904f
C669 VP.n54 B 0.017904f
C670 VP.n55 B 0.017904f
C671 VP.n56 B 0.033201f
C672 VP.n57 B 0.029595f
C673 VP.n58 B 0.612837f
C674 VP.n59 B 0.020417f
C675 VP.n60 B 0.017904f
C676 VP.n61 B 0.017904f
C677 VP.n62 B 0.017904f
C678 VP.n63 B 0.033201f
C679 VP.n64 B 0.03452f
C680 VP.n65 B 0.014829f
C681 VP.n66 B 0.017904f
C682 VP.n67 B 0.017904f
C683 VP.n68 B 0.017904f
C684 VP.n69 B 0.033201f
C685 VP.n70 B 0.033201f
C686 VP.n71 B 0.017794f
C687 VP.n72 B 0.028892f
C688 VP.n73 B 1.25684f
C689 VP.n74 B 1.26802f
C690 VP.n75 B 0.678416f
C691 VP.n76 B 0.017794f
C692 VP.n77 B 0.033201f
C693 VP.n78 B 0.017904f
C694 VP.n79 B 0.017904f
C695 VP.n80 B 0.017904f
C696 VP.n81 B 0.035905f
C697 VP.n82 B 0.014829f
C698 VP.n83 B 0.03452f
C699 VP.n84 B 0.017904f
C700 VP.n85 B 0.017904f
C701 VP.n86 B 0.017904f
C702 VP.n87 B 0.033201f
C703 VP.n88 B 0.020417f
C704 VP.n89 B 0.612837f
C705 VP.n90 B 0.029595f
C706 VP.n91 B 0.017904f
C707 VP.n92 B 0.017904f
C708 VP.n93 B 0.017904f
C709 VP.n94 B 0.033201f
C710 VP.n95 B 0.022559f
C711 VP.n96 B 0.029494f
C712 VP.n97 B 0.017904f
C713 VP.n98 B 0.017904f
C714 VP.n99 B 0.017904f
C715 VP.n100 B 0.033201f
C716 VP.n101 B 0.025006f
C717 VP.n102 B 0.612837f
C718 VP.n103 B 0.025006f
C719 VP.n104 B 0.017904f
C720 VP.n105 B 0.017904f
C721 VP.n106 B 0.017904f
C722 VP.n107 B 0.033201f
C723 VP.n108 B 0.029494f
C724 VP.n109 B 0.022559f
C725 VP.n110 B 0.017904f
C726 VP.n111 B 0.017904f
C727 VP.n112 B 0.017904f
C728 VP.n113 B 0.033201f
C729 VP.n114 B 0.029595f
C730 VP.n115 B 0.612837f
C731 VP.n116 B 0.020417f
C732 VP.n117 B 0.017904f
C733 VP.n118 B 0.017904f
C734 VP.n119 B 0.017904f
C735 VP.n120 B 0.033201f
C736 VP.n121 B 0.03452f
C737 VP.n122 B 0.014829f
C738 VP.n123 B 0.017904f
C739 VP.n124 B 0.017904f
C740 VP.n125 B 0.017904f
C741 VP.n126 B 0.033201f
C742 VP.n127 B 0.033201f
C743 VP.n128 B 0.017794f
C744 VP.n129 B 0.028892f
C745 VP.n130 B 0.055752f
.ends

