* NGSPICE file created from diff_pair_sample_1740.ext - technology: sky130A

.subckt diff_pair_sample_1740 VTAIL VN VP B VDD2 VDD1
X0 B.t11 B.t9 B.t10 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=0 ps=0 w=14.99 l=2.46
X1 VDD2.t5 VN.t0 VTAIL.t6 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=2.47335 ps=15.32 w=14.99 l=2.46
X2 B.t8 B.t6 B.t7 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=0 ps=0 w=14.99 l=2.46
X3 VDD1.t5 VP.t0 VTAIL.t5 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=5.8461 ps=30.76 w=14.99 l=2.46
X4 VTAIL.t4 VP.t1 VDD1.t4 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=2.47335 ps=15.32 w=14.99 l=2.46
X5 VTAIL.t7 VN.t1 VDD2.t4 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=2.47335 ps=15.32 w=14.99 l=2.46
X6 VTAIL.t8 VN.t2 VDD2.t3 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=2.47335 ps=15.32 w=14.99 l=2.46
X7 VDD2.t2 VN.t3 VTAIL.t9 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=5.8461 ps=30.76 w=14.99 l=2.46
X8 VDD1.t3 VP.t2 VTAIL.t2 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=2.47335 ps=15.32 w=14.99 l=2.46
X9 B.t5 B.t3 B.t4 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=0 ps=0 w=14.99 l=2.46
X10 VDD2.t1 VN.t4 VTAIL.t10 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=5.8461 ps=30.76 w=14.99 l=2.46
X11 VDD2.t0 VN.t5 VTAIL.t11 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=2.47335 ps=15.32 w=14.99 l=2.46
X12 B.t2 B.t0 B.t1 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=0 ps=0 w=14.99 l=2.46
X13 VDD1.t2 VP.t3 VTAIL.t3 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=5.8461 ps=30.76 w=14.99 l=2.46
X14 VDD1.t1 VP.t4 VTAIL.t1 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=5.8461 pd=30.76 as=2.47335 ps=15.32 w=14.99 l=2.46
X15 VTAIL.t0 VP.t5 VDD1.t0 w_n3202_n3966# sky130_fd_pr__pfet_01v8 ad=2.47335 pd=15.32 as=2.47335 ps=15.32 w=14.99 l=2.46
R0 B.n555 B.n82 585
R1 B.n557 B.n556 585
R2 B.n558 B.n81 585
R3 B.n560 B.n559 585
R4 B.n561 B.n80 585
R5 B.n563 B.n562 585
R6 B.n564 B.n79 585
R7 B.n566 B.n565 585
R8 B.n567 B.n78 585
R9 B.n569 B.n568 585
R10 B.n570 B.n77 585
R11 B.n572 B.n571 585
R12 B.n573 B.n76 585
R13 B.n575 B.n574 585
R14 B.n576 B.n75 585
R15 B.n578 B.n577 585
R16 B.n579 B.n74 585
R17 B.n581 B.n580 585
R18 B.n582 B.n73 585
R19 B.n584 B.n583 585
R20 B.n585 B.n72 585
R21 B.n587 B.n586 585
R22 B.n588 B.n71 585
R23 B.n590 B.n589 585
R24 B.n591 B.n70 585
R25 B.n593 B.n592 585
R26 B.n594 B.n69 585
R27 B.n596 B.n595 585
R28 B.n597 B.n68 585
R29 B.n599 B.n598 585
R30 B.n600 B.n67 585
R31 B.n602 B.n601 585
R32 B.n603 B.n66 585
R33 B.n605 B.n604 585
R34 B.n606 B.n65 585
R35 B.n608 B.n607 585
R36 B.n609 B.n64 585
R37 B.n611 B.n610 585
R38 B.n612 B.n63 585
R39 B.n614 B.n613 585
R40 B.n615 B.n62 585
R41 B.n617 B.n616 585
R42 B.n618 B.n61 585
R43 B.n620 B.n619 585
R44 B.n621 B.n60 585
R45 B.n623 B.n622 585
R46 B.n624 B.n59 585
R47 B.n626 B.n625 585
R48 B.n627 B.n55 585
R49 B.n629 B.n628 585
R50 B.n630 B.n54 585
R51 B.n632 B.n631 585
R52 B.n633 B.n53 585
R53 B.n635 B.n634 585
R54 B.n636 B.n52 585
R55 B.n638 B.n637 585
R56 B.n639 B.n51 585
R57 B.n641 B.n640 585
R58 B.n642 B.n50 585
R59 B.n644 B.n643 585
R60 B.n646 B.n47 585
R61 B.n648 B.n647 585
R62 B.n649 B.n46 585
R63 B.n651 B.n650 585
R64 B.n652 B.n45 585
R65 B.n654 B.n653 585
R66 B.n655 B.n44 585
R67 B.n657 B.n656 585
R68 B.n658 B.n43 585
R69 B.n660 B.n659 585
R70 B.n661 B.n42 585
R71 B.n663 B.n662 585
R72 B.n664 B.n41 585
R73 B.n666 B.n665 585
R74 B.n667 B.n40 585
R75 B.n669 B.n668 585
R76 B.n670 B.n39 585
R77 B.n672 B.n671 585
R78 B.n673 B.n38 585
R79 B.n675 B.n674 585
R80 B.n676 B.n37 585
R81 B.n678 B.n677 585
R82 B.n679 B.n36 585
R83 B.n681 B.n680 585
R84 B.n682 B.n35 585
R85 B.n684 B.n683 585
R86 B.n685 B.n34 585
R87 B.n687 B.n686 585
R88 B.n688 B.n33 585
R89 B.n690 B.n689 585
R90 B.n691 B.n32 585
R91 B.n693 B.n692 585
R92 B.n694 B.n31 585
R93 B.n696 B.n695 585
R94 B.n697 B.n30 585
R95 B.n699 B.n698 585
R96 B.n700 B.n29 585
R97 B.n702 B.n701 585
R98 B.n703 B.n28 585
R99 B.n705 B.n704 585
R100 B.n706 B.n27 585
R101 B.n708 B.n707 585
R102 B.n709 B.n26 585
R103 B.n711 B.n710 585
R104 B.n712 B.n25 585
R105 B.n714 B.n713 585
R106 B.n715 B.n24 585
R107 B.n717 B.n716 585
R108 B.n718 B.n23 585
R109 B.n720 B.n719 585
R110 B.n554 B.n553 585
R111 B.n552 B.n83 585
R112 B.n551 B.n550 585
R113 B.n549 B.n84 585
R114 B.n548 B.n547 585
R115 B.n546 B.n85 585
R116 B.n545 B.n544 585
R117 B.n543 B.n86 585
R118 B.n542 B.n541 585
R119 B.n540 B.n87 585
R120 B.n539 B.n538 585
R121 B.n537 B.n88 585
R122 B.n536 B.n535 585
R123 B.n534 B.n89 585
R124 B.n533 B.n532 585
R125 B.n531 B.n90 585
R126 B.n530 B.n529 585
R127 B.n528 B.n91 585
R128 B.n527 B.n526 585
R129 B.n525 B.n92 585
R130 B.n524 B.n523 585
R131 B.n522 B.n93 585
R132 B.n521 B.n520 585
R133 B.n519 B.n94 585
R134 B.n518 B.n517 585
R135 B.n516 B.n95 585
R136 B.n515 B.n514 585
R137 B.n513 B.n96 585
R138 B.n512 B.n511 585
R139 B.n510 B.n97 585
R140 B.n509 B.n508 585
R141 B.n507 B.n98 585
R142 B.n506 B.n505 585
R143 B.n504 B.n99 585
R144 B.n503 B.n502 585
R145 B.n501 B.n100 585
R146 B.n500 B.n499 585
R147 B.n498 B.n101 585
R148 B.n497 B.n496 585
R149 B.n495 B.n102 585
R150 B.n494 B.n493 585
R151 B.n492 B.n103 585
R152 B.n491 B.n490 585
R153 B.n489 B.n104 585
R154 B.n488 B.n487 585
R155 B.n486 B.n105 585
R156 B.n485 B.n484 585
R157 B.n483 B.n106 585
R158 B.n482 B.n481 585
R159 B.n480 B.n107 585
R160 B.n479 B.n478 585
R161 B.n477 B.n108 585
R162 B.n476 B.n475 585
R163 B.n474 B.n109 585
R164 B.n473 B.n472 585
R165 B.n471 B.n110 585
R166 B.n470 B.n469 585
R167 B.n468 B.n111 585
R168 B.n467 B.n466 585
R169 B.n465 B.n112 585
R170 B.n464 B.n463 585
R171 B.n462 B.n113 585
R172 B.n461 B.n460 585
R173 B.n459 B.n114 585
R174 B.n458 B.n457 585
R175 B.n456 B.n115 585
R176 B.n455 B.n454 585
R177 B.n453 B.n116 585
R178 B.n452 B.n451 585
R179 B.n450 B.n117 585
R180 B.n449 B.n448 585
R181 B.n447 B.n118 585
R182 B.n446 B.n445 585
R183 B.n444 B.n119 585
R184 B.n443 B.n442 585
R185 B.n441 B.n120 585
R186 B.n440 B.n439 585
R187 B.n438 B.n121 585
R188 B.n437 B.n436 585
R189 B.n435 B.n122 585
R190 B.n434 B.n433 585
R191 B.n432 B.n123 585
R192 B.n431 B.n430 585
R193 B.n264 B.n183 585
R194 B.n266 B.n265 585
R195 B.n267 B.n182 585
R196 B.n269 B.n268 585
R197 B.n270 B.n181 585
R198 B.n272 B.n271 585
R199 B.n273 B.n180 585
R200 B.n275 B.n274 585
R201 B.n276 B.n179 585
R202 B.n278 B.n277 585
R203 B.n279 B.n178 585
R204 B.n281 B.n280 585
R205 B.n282 B.n177 585
R206 B.n284 B.n283 585
R207 B.n285 B.n176 585
R208 B.n287 B.n286 585
R209 B.n288 B.n175 585
R210 B.n290 B.n289 585
R211 B.n291 B.n174 585
R212 B.n293 B.n292 585
R213 B.n294 B.n173 585
R214 B.n296 B.n295 585
R215 B.n297 B.n172 585
R216 B.n299 B.n298 585
R217 B.n300 B.n171 585
R218 B.n302 B.n301 585
R219 B.n303 B.n170 585
R220 B.n305 B.n304 585
R221 B.n306 B.n169 585
R222 B.n308 B.n307 585
R223 B.n309 B.n168 585
R224 B.n311 B.n310 585
R225 B.n312 B.n167 585
R226 B.n314 B.n313 585
R227 B.n315 B.n166 585
R228 B.n317 B.n316 585
R229 B.n318 B.n165 585
R230 B.n320 B.n319 585
R231 B.n321 B.n164 585
R232 B.n323 B.n322 585
R233 B.n324 B.n163 585
R234 B.n326 B.n325 585
R235 B.n327 B.n162 585
R236 B.n329 B.n328 585
R237 B.n330 B.n161 585
R238 B.n332 B.n331 585
R239 B.n333 B.n160 585
R240 B.n335 B.n334 585
R241 B.n336 B.n159 585
R242 B.n338 B.n337 585
R243 B.n340 B.n156 585
R244 B.n342 B.n341 585
R245 B.n343 B.n155 585
R246 B.n345 B.n344 585
R247 B.n346 B.n154 585
R248 B.n348 B.n347 585
R249 B.n349 B.n153 585
R250 B.n351 B.n350 585
R251 B.n352 B.n152 585
R252 B.n354 B.n353 585
R253 B.n356 B.n355 585
R254 B.n357 B.n148 585
R255 B.n359 B.n358 585
R256 B.n360 B.n147 585
R257 B.n362 B.n361 585
R258 B.n363 B.n146 585
R259 B.n365 B.n364 585
R260 B.n366 B.n145 585
R261 B.n368 B.n367 585
R262 B.n369 B.n144 585
R263 B.n371 B.n370 585
R264 B.n372 B.n143 585
R265 B.n374 B.n373 585
R266 B.n375 B.n142 585
R267 B.n377 B.n376 585
R268 B.n378 B.n141 585
R269 B.n380 B.n379 585
R270 B.n381 B.n140 585
R271 B.n383 B.n382 585
R272 B.n384 B.n139 585
R273 B.n386 B.n385 585
R274 B.n387 B.n138 585
R275 B.n389 B.n388 585
R276 B.n390 B.n137 585
R277 B.n392 B.n391 585
R278 B.n393 B.n136 585
R279 B.n395 B.n394 585
R280 B.n396 B.n135 585
R281 B.n398 B.n397 585
R282 B.n399 B.n134 585
R283 B.n401 B.n400 585
R284 B.n402 B.n133 585
R285 B.n404 B.n403 585
R286 B.n405 B.n132 585
R287 B.n407 B.n406 585
R288 B.n408 B.n131 585
R289 B.n410 B.n409 585
R290 B.n411 B.n130 585
R291 B.n413 B.n412 585
R292 B.n414 B.n129 585
R293 B.n416 B.n415 585
R294 B.n417 B.n128 585
R295 B.n419 B.n418 585
R296 B.n420 B.n127 585
R297 B.n422 B.n421 585
R298 B.n423 B.n126 585
R299 B.n425 B.n424 585
R300 B.n426 B.n125 585
R301 B.n428 B.n427 585
R302 B.n429 B.n124 585
R303 B.n263 B.n262 585
R304 B.n261 B.n184 585
R305 B.n260 B.n259 585
R306 B.n258 B.n185 585
R307 B.n257 B.n256 585
R308 B.n255 B.n186 585
R309 B.n254 B.n253 585
R310 B.n252 B.n187 585
R311 B.n251 B.n250 585
R312 B.n249 B.n188 585
R313 B.n248 B.n247 585
R314 B.n246 B.n189 585
R315 B.n245 B.n244 585
R316 B.n243 B.n190 585
R317 B.n242 B.n241 585
R318 B.n240 B.n191 585
R319 B.n239 B.n238 585
R320 B.n237 B.n192 585
R321 B.n236 B.n235 585
R322 B.n234 B.n193 585
R323 B.n233 B.n232 585
R324 B.n231 B.n194 585
R325 B.n230 B.n229 585
R326 B.n228 B.n195 585
R327 B.n227 B.n226 585
R328 B.n225 B.n196 585
R329 B.n224 B.n223 585
R330 B.n222 B.n197 585
R331 B.n221 B.n220 585
R332 B.n219 B.n198 585
R333 B.n218 B.n217 585
R334 B.n216 B.n199 585
R335 B.n215 B.n214 585
R336 B.n213 B.n200 585
R337 B.n212 B.n211 585
R338 B.n210 B.n201 585
R339 B.n209 B.n208 585
R340 B.n207 B.n202 585
R341 B.n206 B.n205 585
R342 B.n204 B.n203 585
R343 B.n2 B.n0 585
R344 B.n781 B.n1 585
R345 B.n780 B.n779 585
R346 B.n778 B.n3 585
R347 B.n777 B.n776 585
R348 B.n775 B.n4 585
R349 B.n774 B.n773 585
R350 B.n772 B.n5 585
R351 B.n771 B.n770 585
R352 B.n769 B.n6 585
R353 B.n768 B.n767 585
R354 B.n766 B.n7 585
R355 B.n765 B.n764 585
R356 B.n763 B.n8 585
R357 B.n762 B.n761 585
R358 B.n760 B.n9 585
R359 B.n759 B.n758 585
R360 B.n757 B.n10 585
R361 B.n756 B.n755 585
R362 B.n754 B.n11 585
R363 B.n753 B.n752 585
R364 B.n751 B.n12 585
R365 B.n750 B.n749 585
R366 B.n748 B.n13 585
R367 B.n747 B.n746 585
R368 B.n745 B.n14 585
R369 B.n744 B.n743 585
R370 B.n742 B.n15 585
R371 B.n741 B.n740 585
R372 B.n739 B.n16 585
R373 B.n738 B.n737 585
R374 B.n736 B.n17 585
R375 B.n735 B.n734 585
R376 B.n733 B.n18 585
R377 B.n732 B.n731 585
R378 B.n730 B.n19 585
R379 B.n729 B.n728 585
R380 B.n727 B.n20 585
R381 B.n726 B.n725 585
R382 B.n724 B.n21 585
R383 B.n723 B.n722 585
R384 B.n721 B.n22 585
R385 B.n783 B.n782 585
R386 B.n264 B.n263 521.33
R387 B.n721 B.n720 521.33
R388 B.n431 B.n124 521.33
R389 B.n553 B.n82 521.33
R390 B.n149 B.t0 354.678
R391 B.n157 B.t6 354.678
R392 B.n48 B.t9 354.678
R393 B.n56 B.t3 354.678
R394 B.n263 B.n184 163.367
R395 B.n259 B.n184 163.367
R396 B.n259 B.n258 163.367
R397 B.n258 B.n257 163.367
R398 B.n257 B.n186 163.367
R399 B.n253 B.n186 163.367
R400 B.n253 B.n252 163.367
R401 B.n252 B.n251 163.367
R402 B.n251 B.n188 163.367
R403 B.n247 B.n188 163.367
R404 B.n247 B.n246 163.367
R405 B.n246 B.n245 163.367
R406 B.n245 B.n190 163.367
R407 B.n241 B.n190 163.367
R408 B.n241 B.n240 163.367
R409 B.n240 B.n239 163.367
R410 B.n239 B.n192 163.367
R411 B.n235 B.n192 163.367
R412 B.n235 B.n234 163.367
R413 B.n234 B.n233 163.367
R414 B.n233 B.n194 163.367
R415 B.n229 B.n194 163.367
R416 B.n229 B.n228 163.367
R417 B.n228 B.n227 163.367
R418 B.n227 B.n196 163.367
R419 B.n223 B.n196 163.367
R420 B.n223 B.n222 163.367
R421 B.n222 B.n221 163.367
R422 B.n221 B.n198 163.367
R423 B.n217 B.n198 163.367
R424 B.n217 B.n216 163.367
R425 B.n216 B.n215 163.367
R426 B.n215 B.n200 163.367
R427 B.n211 B.n200 163.367
R428 B.n211 B.n210 163.367
R429 B.n210 B.n209 163.367
R430 B.n209 B.n202 163.367
R431 B.n205 B.n202 163.367
R432 B.n205 B.n204 163.367
R433 B.n204 B.n2 163.367
R434 B.n782 B.n2 163.367
R435 B.n782 B.n781 163.367
R436 B.n781 B.n780 163.367
R437 B.n780 B.n3 163.367
R438 B.n776 B.n3 163.367
R439 B.n776 B.n775 163.367
R440 B.n775 B.n774 163.367
R441 B.n774 B.n5 163.367
R442 B.n770 B.n5 163.367
R443 B.n770 B.n769 163.367
R444 B.n769 B.n768 163.367
R445 B.n768 B.n7 163.367
R446 B.n764 B.n7 163.367
R447 B.n764 B.n763 163.367
R448 B.n763 B.n762 163.367
R449 B.n762 B.n9 163.367
R450 B.n758 B.n9 163.367
R451 B.n758 B.n757 163.367
R452 B.n757 B.n756 163.367
R453 B.n756 B.n11 163.367
R454 B.n752 B.n11 163.367
R455 B.n752 B.n751 163.367
R456 B.n751 B.n750 163.367
R457 B.n750 B.n13 163.367
R458 B.n746 B.n13 163.367
R459 B.n746 B.n745 163.367
R460 B.n745 B.n744 163.367
R461 B.n744 B.n15 163.367
R462 B.n740 B.n15 163.367
R463 B.n740 B.n739 163.367
R464 B.n739 B.n738 163.367
R465 B.n738 B.n17 163.367
R466 B.n734 B.n17 163.367
R467 B.n734 B.n733 163.367
R468 B.n733 B.n732 163.367
R469 B.n732 B.n19 163.367
R470 B.n728 B.n19 163.367
R471 B.n728 B.n727 163.367
R472 B.n727 B.n726 163.367
R473 B.n726 B.n21 163.367
R474 B.n722 B.n21 163.367
R475 B.n722 B.n721 163.367
R476 B.n265 B.n264 163.367
R477 B.n265 B.n182 163.367
R478 B.n269 B.n182 163.367
R479 B.n270 B.n269 163.367
R480 B.n271 B.n270 163.367
R481 B.n271 B.n180 163.367
R482 B.n275 B.n180 163.367
R483 B.n276 B.n275 163.367
R484 B.n277 B.n276 163.367
R485 B.n277 B.n178 163.367
R486 B.n281 B.n178 163.367
R487 B.n282 B.n281 163.367
R488 B.n283 B.n282 163.367
R489 B.n283 B.n176 163.367
R490 B.n287 B.n176 163.367
R491 B.n288 B.n287 163.367
R492 B.n289 B.n288 163.367
R493 B.n289 B.n174 163.367
R494 B.n293 B.n174 163.367
R495 B.n294 B.n293 163.367
R496 B.n295 B.n294 163.367
R497 B.n295 B.n172 163.367
R498 B.n299 B.n172 163.367
R499 B.n300 B.n299 163.367
R500 B.n301 B.n300 163.367
R501 B.n301 B.n170 163.367
R502 B.n305 B.n170 163.367
R503 B.n306 B.n305 163.367
R504 B.n307 B.n306 163.367
R505 B.n307 B.n168 163.367
R506 B.n311 B.n168 163.367
R507 B.n312 B.n311 163.367
R508 B.n313 B.n312 163.367
R509 B.n313 B.n166 163.367
R510 B.n317 B.n166 163.367
R511 B.n318 B.n317 163.367
R512 B.n319 B.n318 163.367
R513 B.n319 B.n164 163.367
R514 B.n323 B.n164 163.367
R515 B.n324 B.n323 163.367
R516 B.n325 B.n324 163.367
R517 B.n325 B.n162 163.367
R518 B.n329 B.n162 163.367
R519 B.n330 B.n329 163.367
R520 B.n331 B.n330 163.367
R521 B.n331 B.n160 163.367
R522 B.n335 B.n160 163.367
R523 B.n336 B.n335 163.367
R524 B.n337 B.n336 163.367
R525 B.n337 B.n156 163.367
R526 B.n342 B.n156 163.367
R527 B.n343 B.n342 163.367
R528 B.n344 B.n343 163.367
R529 B.n344 B.n154 163.367
R530 B.n348 B.n154 163.367
R531 B.n349 B.n348 163.367
R532 B.n350 B.n349 163.367
R533 B.n350 B.n152 163.367
R534 B.n354 B.n152 163.367
R535 B.n355 B.n354 163.367
R536 B.n355 B.n148 163.367
R537 B.n359 B.n148 163.367
R538 B.n360 B.n359 163.367
R539 B.n361 B.n360 163.367
R540 B.n361 B.n146 163.367
R541 B.n365 B.n146 163.367
R542 B.n366 B.n365 163.367
R543 B.n367 B.n366 163.367
R544 B.n367 B.n144 163.367
R545 B.n371 B.n144 163.367
R546 B.n372 B.n371 163.367
R547 B.n373 B.n372 163.367
R548 B.n373 B.n142 163.367
R549 B.n377 B.n142 163.367
R550 B.n378 B.n377 163.367
R551 B.n379 B.n378 163.367
R552 B.n379 B.n140 163.367
R553 B.n383 B.n140 163.367
R554 B.n384 B.n383 163.367
R555 B.n385 B.n384 163.367
R556 B.n385 B.n138 163.367
R557 B.n389 B.n138 163.367
R558 B.n390 B.n389 163.367
R559 B.n391 B.n390 163.367
R560 B.n391 B.n136 163.367
R561 B.n395 B.n136 163.367
R562 B.n396 B.n395 163.367
R563 B.n397 B.n396 163.367
R564 B.n397 B.n134 163.367
R565 B.n401 B.n134 163.367
R566 B.n402 B.n401 163.367
R567 B.n403 B.n402 163.367
R568 B.n403 B.n132 163.367
R569 B.n407 B.n132 163.367
R570 B.n408 B.n407 163.367
R571 B.n409 B.n408 163.367
R572 B.n409 B.n130 163.367
R573 B.n413 B.n130 163.367
R574 B.n414 B.n413 163.367
R575 B.n415 B.n414 163.367
R576 B.n415 B.n128 163.367
R577 B.n419 B.n128 163.367
R578 B.n420 B.n419 163.367
R579 B.n421 B.n420 163.367
R580 B.n421 B.n126 163.367
R581 B.n425 B.n126 163.367
R582 B.n426 B.n425 163.367
R583 B.n427 B.n426 163.367
R584 B.n427 B.n124 163.367
R585 B.n432 B.n431 163.367
R586 B.n433 B.n432 163.367
R587 B.n433 B.n122 163.367
R588 B.n437 B.n122 163.367
R589 B.n438 B.n437 163.367
R590 B.n439 B.n438 163.367
R591 B.n439 B.n120 163.367
R592 B.n443 B.n120 163.367
R593 B.n444 B.n443 163.367
R594 B.n445 B.n444 163.367
R595 B.n445 B.n118 163.367
R596 B.n449 B.n118 163.367
R597 B.n450 B.n449 163.367
R598 B.n451 B.n450 163.367
R599 B.n451 B.n116 163.367
R600 B.n455 B.n116 163.367
R601 B.n456 B.n455 163.367
R602 B.n457 B.n456 163.367
R603 B.n457 B.n114 163.367
R604 B.n461 B.n114 163.367
R605 B.n462 B.n461 163.367
R606 B.n463 B.n462 163.367
R607 B.n463 B.n112 163.367
R608 B.n467 B.n112 163.367
R609 B.n468 B.n467 163.367
R610 B.n469 B.n468 163.367
R611 B.n469 B.n110 163.367
R612 B.n473 B.n110 163.367
R613 B.n474 B.n473 163.367
R614 B.n475 B.n474 163.367
R615 B.n475 B.n108 163.367
R616 B.n479 B.n108 163.367
R617 B.n480 B.n479 163.367
R618 B.n481 B.n480 163.367
R619 B.n481 B.n106 163.367
R620 B.n485 B.n106 163.367
R621 B.n486 B.n485 163.367
R622 B.n487 B.n486 163.367
R623 B.n487 B.n104 163.367
R624 B.n491 B.n104 163.367
R625 B.n492 B.n491 163.367
R626 B.n493 B.n492 163.367
R627 B.n493 B.n102 163.367
R628 B.n497 B.n102 163.367
R629 B.n498 B.n497 163.367
R630 B.n499 B.n498 163.367
R631 B.n499 B.n100 163.367
R632 B.n503 B.n100 163.367
R633 B.n504 B.n503 163.367
R634 B.n505 B.n504 163.367
R635 B.n505 B.n98 163.367
R636 B.n509 B.n98 163.367
R637 B.n510 B.n509 163.367
R638 B.n511 B.n510 163.367
R639 B.n511 B.n96 163.367
R640 B.n515 B.n96 163.367
R641 B.n516 B.n515 163.367
R642 B.n517 B.n516 163.367
R643 B.n517 B.n94 163.367
R644 B.n521 B.n94 163.367
R645 B.n522 B.n521 163.367
R646 B.n523 B.n522 163.367
R647 B.n523 B.n92 163.367
R648 B.n527 B.n92 163.367
R649 B.n528 B.n527 163.367
R650 B.n529 B.n528 163.367
R651 B.n529 B.n90 163.367
R652 B.n533 B.n90 163.367
R653 B.n534 B.n533 163.367
R654 B.n535 B.n534 163.367
R655 B.n535 B.n88 163.367
R656 B.n539 B.n88 163.367
R657 B.n540 B.n539 163.367
R658 B.n541 B.n540 163.367
R659 B.n541 B.n86 163.367
R660 B.n545 B.n86 163.367
R661 B.n546 B.n545 163.367
R662 B.n547 B.n546 163.367
R663 B.n547 B.n84 163.367
R664 B.n551 B.n84 163.367
R665 B.n552 B.n551 163.367
R666 B.n553 B.n552 163.367
R667 B.n720 B.n23 163.367
R668 B.n716 B.n23 163.367
R669 B.n716 B.n715 163.367
R670 B.n715 B.n714 163.367
R671 B.n714 B.n25 163.367
R672 B.n710 B.n25 163.367
R673 B.n710 B.n709 163.367
R674 B.n709 B.n708 163.367
R675 B.n708 B.n27 163.367
R676 B.n704 B.n27 163.367
R677 B.n704 B.n703 163.367
R678 B.n703 B.n702 163.367
R679 B.n702 B.n29 163.367
R680 B.n698 B.n29 163.367
R681 B.n698 B.n697 163.367
R682 B.n697 B.n696 163.367
R683 B.n696 B.n31 163.367
R684 B.n692 B.n31 163.367
R685 B.n692 B.n691 163.367
R686 B.n691 B.n690 163.367
R687 B.n690 B.n33 163.367
R688 B.n686 B.n33 163.367
R689 B.n686 B.n685 163.367
R690 B.n685 B.n684 163.367
R691 B.n684 B.n35 163.367
R692 B.n680 B.n35 163.367
R693 B.n680 B.n679 163.367
R694 B.n679 B.n678 163.367
R695 B.n678 B.n37 163.367
R696 B.n674 B.n37 163.367
R697 B.n674 B.n673 163.367
R698 B.n673 B.n672 163.367
R699 B.n672 B.n39 163.367
R700 B.n668 B.n39 163.367
R701 B.n668 B.n667 163.367
R702 B.n667 B.n666 163.367
R703 B.n666 B.n41 163.367
R704 B.n662 B.n41 163.367
R705 B.n662 B.n661 163.367
R706 B.n661 B.n660 163.367
R707 B.n660 B.n43 163.367
R708 B.n656 B.n43 163.367
R709 B.n656 B.n655 163.367
R710 B.n655 B.n654 163.367
R711 B.n654 B.n45 163.367
R712 B.n650 B.n45 163.367
R713 B.n650 B.n649 163.367
R714 B.n649 B.n648 163.367
R715 B.n648 B.n47 163.367
R716 B.n643 B.n47 163.367
R717 B.n643 B.n642 163.367
R718 B.n642 B.n641 163.367
R719 B.n641 B.n51 163.367
R720 B.n637 B.n51 163.367
R721 B.n637 B.n636 163.367
R722 B.n636 B.n635 163.367
R723 B.n635 B.n53 163.367
R724 B.n631 B.n53 163.367
R725 B.n631 B.n630 163.367
R726 B.n630 B.n629 163.367
R727 B.n629 B.n55 163.367
R728 B.n625 B.n55 163.367
R729 B.n625 B.n624 163.367
R730 B.n624 B.n623 163.367
R731 B.n623 B.n60 163.367
R732 B.n619 B.n60 163.367
R733 B.n619 B.n618 163.367
R734 B.n618 B.n617 163.367
R735 B.n617 B.n62 163.367
R736 B.n613 B.n62 163.367
R737 B.n613 B.n612 163.367
R738 B.n612 B.n611 163.367
R739 B.n611 B.n64 163.367
R740 B.n607 B.n64 163.367
R741 B.n607 B.n606 163.367
R742 B.n606 B.n605 163.367
R743 B.n605 B.n66 163.367
R744 B.n601 B.n66 163.367
R745 B.n601 B.n600 163.367
R746 B.n600 B.n599 163.367
R747 B.n599 B.n68 163.367
R748 B.n595 B.n68 163.367
R749 B.n595 B.n594 163.367
R750 B.n594 B.n593 163.367
R751 B.n593 B.n70 163.367
R752 B.n589 B.n70 163.367
R753 B.n589 B.n588 163.367
R754 B.n588 B.n587 163.367
R755 B.n587 B.n72 163.367
R756 B.n583 B.n72 163.367
R757 B.n583 B.n582 163.367
R758 B.n582 B.n581 163.367
R759 B.n581 B.n74 163.367
R760 B.n577 B.n74 163.367
R761 B.n577 B.n576 163.367
R762 B.n576 B.n575 163.367
R763 B.n575 B.n76 163.367
R764 B.n571 B.n76 163.367
R765 B.n571 B.n570 163.367
R766 B.n570 B.n569 163.367
R767 B.n569 B.n78 163.367
R768 B.n565 B.n78 163.367
R769 B.n565 B.n564 163.367
R770 B.n564 B.n563 163.367
R771 B.n563 B.n80 163.367
R772 B.n559 B.n80 163.367
R773 B.n559 B.n558 163.367
R774 B.n558 B.n557 163.367
R775 B.n557 B.n82 163.367
R776 B.n149 B.t2 161.254
R777 B.n56 B.t4 161.254
R778 B.n157 B.t8 161.234
R779 B.n48 B.t10 161.234
R780 B.n150 B.t1 107.144
R781 B.n57 B.t5 107.144
R782 B.n158 B.t7 107.126
R783 B.n49 B.t11 107.126
R784 B.n151 B.n150 59.5399
R785 B.n339 B.n158 59.5399
R786 B.n645 B.n49 59.5399
R787 B.n58 B.n57 59.5399
R788 B.n150 B.n149 54.1096
R789 B.n158 B.n157 54.1096
R790 B.n49 B.n48 54.1096
R791 B.n57 B.n56 54.1096
R792 B.n719 B.n22 33.8737
R793 B.n555 B.n554 33.8737
R794 B.n430 B.n429 33.8737
R795 B.n262 B.n183 33.8737
R796 B B.n783 18.0485
R797 B.n719 B.n718 10.6151
R798 B.n718 B.n717 10.6151
R799 B.n717 B.n24 10.6151
R800 B.n713 B.n24 10.6151
R801 B.n713 B.n712 10.6151
R802 B.n712 B.n711 10.6151
R803 B.n711 B.n26 10.6151
R804 B.n707 B.n26 10.6151
R805 B.n707 B.n706 10.6151
R806 B.n706 B.n705 10.6151
R807 B.n705 B.n28 10.6151
R808 B.n701 B.n28 10.6151
R809 B.n701 B.n700 10.6151
R810 B.n700 B.n699 10.6151
R811 B.n699 B.n30 10.6151
R812 B.n695 B.n30 10.6151
R813 B.n695 B.n694 10.6151
R814 B.n694 B.n693 10.6151
R815 B.n693 B.n32 10.6151
R816 B.n689 B.n32 10.6151
R817 B.n689 B.n688 10.6151
R818 B.n688 B.n687 10.6151
R819 B.n687 B.n34 10.6151
R820 B.n683 B.n34 10.6151
R821 B.n683 B.n682 10.6151
R822 B.n682 B.n681 10.6151
R823 B.n681 B.n36 10.6151
R824 B.n677 B.n36 10.6151
R825 B.n677 B.n676 10.6151
R826 B.n676 B.n675 10.6151
R827 B.n675 B.n38 10.6151
R828 B.n671 B.n38 10.6151
R829 B.n671 B.n670 10.6151
R830 B.n670 B.n669 10.6151
R831 B.n669 B.n40 10.6151
R832 B.n665 B.n40 10.6151
R833 B.n665 B.n664 10.6151
R834 B.n664 B.n663 10.6151
R835 B.n663 B.n42 10.6151
R836 B.n659 B.n42 10.6151
R837 B.n659 B.n658 10.6151
R838 B.n658 B.n657 10.6151
R839 B.n657 B.n44 10.6151
R840 B.n653 B.n44 10.6151
R841 B.n653 B.n652 10.6151
R842 B.n652 B.n651 10.6151
R843 B.n651 B.n46 10.6151
R844 B.n647 B.n46 10.6151
R845 B.n647 B.n646 10.6151
R846 B.n644 B.n50 10.6151
R847 B.n640 B.n50 10.6151
R848 B.n640 B.n639 10.6151
R849 B.n639 B.n638 10.6151
R850 B.n638 B.n52 10.6151
R851 B.n634 B.n52 10.6151
R852 B.n634 B.n633 10.6151
R853 B.n633 B.n632 10.6151
R854 B.n632 B.n54 10.6151
R855 B.n628 B.n627 10.6151
R856 B.n627 B.n626 10.6151
R857 B.n626 B.n59 10.6151
R858 B.n622 B.n59 10.6151
R859 B.n622 B.n621 10.6151
R860 B.n621 B.n620 10.6151
R861 B.n620 B.n61 10.6151
R862 B.n616 B.n61 10.6151
R863 B.n616 B.n615 10.6151
R864 B.n615 B.n614 10.6151
R865 B.n614 B.n63 10.6151
R866 B.n610 B.n63 10.6151
R867 B.n610 B.n609 10.6151
R868 B.n609 B.n608 10.6151
R869 B.n608 B.n65 10.6151
R870 B.n604 B.n65 10.6151
R871 B.n604 B.n603 10.6151
R872 B.n603 B.n602 10.6151
R873 B.n602 B.n67 10.6151
R874 B.n598 B.n67 10.6151
R875 B.n598 B.n597 10.6151
R876 B.n597 B.n596 10.6151
R877 B.n596 B.n69 10.6151
R878 B.n592 B.n69 10.6151
R879 B.n592 B.n591 10.6151
R880 B.n591 B.n590 10.6151
R881 B.n590 B.n71 10.6151
R882 B.n586 B.n71 10.6151
R883 B.n586 B.n585 10.6151
R884 B.n585 B.n584 10.6151
R885 B.n584 B.n73 10.6151
R886 B.n580 B.n73 10.6151
R887 B.n580 B.n579 10.6151
R888 B.n579 B.n578 10.6151
R889 B.n578 B.n75 10.6151
R890 B.n574 B.n75 10.6151
R891 B.n574 B.n573 10.6151
R892 B.n573 B.n572 10.6151
R893 B.n572 B.n77 10.6151
R894 B.n568 B.n77 10.6151
R895 B.n568 B.n567 10.6151
R896 B.n567 B.n566 10.6151
R897 B.n566 B.n79 10.6151
R898 B.n562 B.n79 10.6151
R899 B.n562 B.n561 10.6151
R900 B.n561 B.n560 10.6151
R901 B.n560 B.n81 10.6151
R902 B.n556 B.n81 10.6151
R903 B.n556 B.n555 10.6151
R904 B.n430 B.n123 10.6151
R905 B.n434 B.n123 10.6151
R906 B.n435 B.n434 10.6151
R907 B.n436 B.n435 10.6151
R908 B.n436 B.n121 10.6151
R909 B.n440 B.n121 10.6151
R910 B.n441 B.n440 10.6151
R911 B.n442 B.n441 10.6151
R912 B.n442 B.n119 10.6151
R913 B.n446 B.n119 10.6151
R914 B.n447 B.n446 10.6151
R915 B.n448 B.n447 10.6151
R916 B.n448 B.n117 10.6151
R917 B.n452 B.n117 10.6151
R918 B.n453 B.n452 10.6151
R919 B.n454 B.n453 10.6151
R920 B.n454 B.n115 10.6151
R921 B.n458 B.n115 10.6151
R922 B.n459 B.n458 10.6151
R923 B.n460 B.n459 10.6151
R924 B.n460 B.n113 10.6151
R925 B.n464 B.n113 10.6151
R926 B.n465 B.n464 10.6151
R927 B.n466 B.n465 10.6151
R928 B.n466 B.n111 10.6151
R929 B.n470 B.n111 10.6151
R930 B.n471 B.n470 10.6151
R931 B.n472 B.n471 10.6151
R932 B.n472 B.n109 10.6151
R933 B.n476 B.n109 10.6151
R934 B.n477 B.n476 10.6151
R935 B.n478 B.n477 10.6151
R936 B.n478 B.n107 10.6151
R937 B.n482 B.n107 10.6151
R938 B.n483 B.n482 10.6151
R939 B.n484 B.n483 10.6151
R940 B.n484 B.n105 10.6151
R941 B.n488 B.n105 10.6151
R942 B.n489 B.n488 10.6151
R943 B.n490 B.n489 10.6151
R944 B.n490 B.n103 10.6151
R945 B.n494 B.n103 10.6151
R946 B.n495 B.n494 10.6151
R947 B.n496 B.n495 10.6151
R948 B.n496 B.n101 10.6151
R949 B.n500 B.n101 10.6151
R950 B.n501 B.n500 10.6151
R951 B.n502 B.n501 10.6151
R952 B.n502 B.n99 10.6151
R953 B.n506 B.n99 10.6151
R954 B.n507 B.n506 10.6151
R955 B.n508 B.n507 10.6151
R956 B.n508 B.n97 10.6151
R957 B.n512 B.n97 10.6151
R958 B.n513 B.n512 10.6151
R959 B.n514 B.n513 10.6151
R960 B.n514 B.n95 10.6151
R961 B.n518 B.n95 10.6151
R962 B.n519 B.n518 10.6151
R963 B.n520 B.n519 10.6151
R964 B.n520 B.n93 10.6151
R965 B.n524 B.n93 10.6151
R966 B.n525 B.n524 10.6151
R967 B.n526 B.n525 10.6151
R968 B.n526 B.n91 10.6151
R969 B.n530 B.n91 10.6151
R970 B.n531 B.n530 10.6151
R971 B.n532 B.n531 10.6151
R972 B.n532 B.n89 10.6151
R973 B.n536 B.n89 10.6151
R974 B.n537 B.n536 10.6151
R975 B.n538 B.n537 10.6151
R976 B.n538 B.n87 10.6151
R977 B.n542 B.n87 10.6151
R978 B.n543 B.n542 10.6151
R979 B.n544 B.n543 10.6151
R980 B.n544 B.n85 10.6151
R981 B.n548 B.n85 10.6151
R982 B.n549 B.n548 10.6151
R983 B.n550 B.n549 10.6151
R984 B.n550 B.n83 10.6151
R985 B.n554 B.n83 10.6151
R986 B.n266 B.n183 10.6151
R987 B.n267 B.n266 10.6151
R988 B.n268 B.n267 10.6151
R989 B.n268 B.n181 10.6151
R990 B.n272 B.n181 10.6151
R991 B.n273 B.n272 10.6151
R992 B.n274 B.n273 10.6151
R993 B.n274 B.n179 10.6151
R994 B.n278 B.n179 10.6151
R995 B.n279 B.n278 10.6151
R996 B.n280 B.n279 10.6151
R997 B.n280 B.n177 10.6151
R998 B.n284 B.n177 10.6151
R999 B.n285 B.n284 10.6151
R1000 B.n286 B.n285 10.6151
R1001 B.n286 B.n175 10.6151
R1002 B.n290 B.n175 10.6151
R1003 B.n291 B.n290 10.6151
R1004 B.n292 B.n291 10.6151
R1005 B.n292 B.n173 10.6151
R1006 B.n296 B.n173 10.6151
R1007 B.n297 B.n296 10.6151
R1008 B.n298 B.n297 10.6151
R1009 B.n298 B.n171 10.6151
R1010 B.n302 B.n171 10.6151
R1011 B.n303 B.n302 10.6151
R1012 B.n304 B.n303 10.6151
R1013 B.n304 B.n169 10.6151
R1014 B.n308 B.n169 10.6151
R1015 B.n309 B.n308 10.6151
R1016 B.n310 B.n309 10.6151
R1017 B.n310 B.n167 10.6151
R1018 B.n314 B.n167 10.6151
R1019 B.n315 B.n314 10.6151
R1020 B.n316 B.n315 10.6151
R1021 B.n316 B.n165 10.6151
R1022 B.n320 B.n165 10.6151
R1023 B.n321 B.n320 10.6151
R1024 B.n322 B.n321 10.6151
R1025 B.n322 B.n163 10.6151
R1026 B.n326 B.n163 10.6151
R1027 B.n327 B.n326 10.6151
R1028 B.n328 B.n327 10.6151
R1029 B.n328 B.n161 10.6151
R1030 B.n332 B.n161 10.6151
R1031 B.n333 B.n332 10.6151
R1032 B.n334 B.n333 10.6151
R1033 B.n334 B.n159 10.6151
R1034 B.n338 B.n159 10.6151
R1035 B.n341 B.n340 10.6151
R1036 B.n341 B.n155 10.6151
R1037 B.n345 B.n155 10.6151
R1038 B.n346 B.n345 10.6151
R1039 B.n347 B.n346 10.6151
R1040 B.n347 B.n153 10.6151
R1041 B.n351 B.n153 10.6151
R1042 B.n352 B.n351 10.6151
R1043 B.n353 B.n352 10.6151
R1044 B.n357 B.n356 10.6151
R1045 B.n358 B.n357 10.6151
R1046 B.n358 B.n147 10.6151
R1047 B.n362 B.n147 10.6151
R1048 B.n363 B.n362 10.6151
R1049 B.n364 B.n363 10.6151
R1050 B.n364 B.n145 10.6151
R1051 B.n368 B.n145 10.6151
R1052 B.n369 B.n368 10.6151
R1053 B.n370 B.n369 10.6151
R1054 B.n370 B.n143 10.6151
R1055 B.n374 B.n143 10.6151
R1056 B.n375 B.n374 10.6151
R1057 B.n376 B.n375 10.6151
R1058 B.n376 B.n141 10.6151
R1059 B.n380 B.n141 10.6151
R1060 B.n381 B.n380 10.6151
R1061 B.n382 B.n381 10.6151
R1062 B.n382 B.n139 10.6151
R1063 B.n386 B.n139 10.6151
R1064 B.n387 B.n386 10.6151
R1065 B.n388 B.n387 10.6151
R1066 B.n388 B.n137 10.6151
R1067 B.n392 B.n137 10.6151
R1068 B.n393 B.n392 10.6151
R1069 B.n394 B.n393 10.6151
R1070 B.n394 B.n135 10.6151
R1071 B.n398 B.n135 10.6151
R1072 B.n399 B.n398 10.6151
R1073 B.n400 B.n399 10.6151
R1074 B.n400 B.n133 10.6151
R1075 B.n404 B.n133 10.6151
R1076 B.n405 B.n404 10.6151
R1077 B.n406 B.n405 10.6151
R1078 B.n406 B.n131 10.6151
R1079 B.n410 B.n131 10.6151
R1080 B.n411 B.n410 10.6151
R1081 B.n412 B.n411 10.6151
R1082 B.n412 B.n129 10.6151
R1083 B.n416 B.n129 10.6151
R1084 B.n417 B.n416 10.6151
R1085 B.n418 B.n417 10.6151
R1086 B.n418 B.n127 10.6151
R1087 B.n422 B.n127 10.6151
R1088 B.n423 B.n422 10.6151
R1089 B.n424 B.n423 10.6151
R1090 B.n424 B.n125 10.6151
R1091 B.n428 B.n125 10.6151
R1092 B.n429 B.n428 10.6151
R1093 B.n262 B.n261 10.6151
R1094 B.n261 B.n260 10.6151
R1095 B.n260 B.n185 10.6151
R1096 B.n256 B.n185 10.6151
R1097 B.n256 B.n255 10.6151
R1098 B.n255 B.n254 10.6151
R1099 B.n254 B.n187 10.6151
R1100 B.n250 B.n187 10.6151
R1101 B.n250 B.n249 10.6151
R1102 B.n249 B.n248 10.6151
R1103 B.n248 B.n189 10.6151
R1104 B.n244 B.n189 10.6151
R1105 B.n244 B.n243 10.6151
R1106 B.n243 B.n242 10.6151
R1107 B.n242 B.n191 10.6151
R1108 B.n238 B.n191 10.6151
R1109 B.n238 B.n237 10.6151
R1110 B.n237 B.n236 10.6151
R1111 B.n236 B.n193 10.6151
R1112 B.n232 B.n193 10.6151
R1113 B.n232 B.n231 10.6151
R1114 B.n231 B.n230 10.6151
R1115 B.n230 B.n195 10.6151
R1116 B.n226 B.n195 10.6151
R1117 B.n226 B.n225 10.6151
R1118 B.n225 B.n224 10.6151
R1119 B.n224 B.n197 10.6151
R1120 B.n220 B.n197 10.6151
R1121 B.n220 B.n219 10.6151
R1122 B.n219 B.n218 10.6151
R1123 B.n218 B.n199 10.6151
R1124 B.n214 B.n199 10.6151
R1125 B.n214 B.n213 10.6151
R1126 B.n213 B.n212 10.6151
R1127 B.n212 B.n201 10.6151
R1128 B.n208 B.n201 10.6151
R1129 B.n208 B.n207 10.6151
R1130 B.n207 B.n206 10.6151
R1131 B.n206 B.n203 10.6151
R1132 B.n203 B.n0 10.6151
R1133 B.n779 B.n1 10.6151
R1134 B.n779 B.n778 10.6151
R1135 B.n778 B.n777 10.6151
R1136 B.n777 B.n4 10.6151
R1137 B.n773 B.n4 10.6151
R1138 B.n773 B.n772 10.6151
R1139 B.n772 B.n771 10.6151
R1140 B.n771 B.n6 10.6151
R1141 B.n767 B.n6 10.6151
R1142 B.n767 B.n766 10.6151
R1143 B.n766 B.n765 10.6151
R1144 B.n765 B.n8 10.6151
R1145 B.n761 B.n8 10.6151
R1146 B.n761 B.n760 10.6151
R1147 B.n760 B.n759 10.6151
R1148 B.n759 B.n10 10.6151
R1149 B.n755 B.n10 10.6151
R1150 B.n755 B.n754 10.6151
R1151 B.n754 B.n753 10.6151
R1152 B.n753 B.n12 10.6151
R1153 B.n749 B.n12 10.6151
R1154 B.n749 B.n748 10.6151
R1155 B.n748 B.n747 10.6151
R1156 B.n747 B.n14 10.6151
R1157 B.n743 B.n14 10.6151
R1158 B.n743 B.n742 10.6151
R1159 B.n742 B.n741 10.6151
R1160 B.n741 B.n16 10.6151
R1161 B.n737 B.n16 10.6151
R1162 B.n737 B.n736 10.6151
R1163 B.n736 B.n735 10.6151
R1164 B.n735 B.n18 10.6151
R1165 B.n731 B.n18 10.6151
R1166 B.n731 B.n730 10.6151
R1167 B.n730 B.n729 10.6151
R1168 B.n729 B.n20 10.6151
R1169 B.n725 B.n20 10.6151
R1170 B.n725 B.n724 10.6151
R1171 B.n724 B.n723 10.6151
R1172 B.n723 B.n22 10.6151
R1173 B.n646 B.n645 9.36635
R1174 B.n628 B.n58 9.36635
R1175 B.n339 B.n338 9.36635
R1176 B.n356 B.n151 9.36635
R1177 B.n783 B.n0 2.81026
R1178 B.n783 B.n1 2.81026
R1179 B.n645 B.n644 1.24928
R1180 B.n58 B.n54 1.24928
R1181 B.n340 B.n339 1.24928
R1182 B.n353 B.n151 1.24928
R1183 VN.n3 VN.t5 181.786
R1184 VN.n17 VN.t3 181.786
R1185 VN.n25 VN.n14 161.3
R1186 VN.n24 VN.n23 161.3
R1187 VN.n22 VN.n15 161.3
R1188 VN.n21 VN.n20 161.3
R1189 VN.n19 VN.n16 161.3
R1190 VN.n11 VN.n0 161.3
R1191 VN.n10 VN.n9 161.3
R1192 VN.n8 VN.n1 161.3
R1193 VN.n7 VN.n6 161.3
R1194 VN.n5 VN.n2 161.3
R1195 VN.n4 VN.t2 146.853
R1196 VN.n12 VN.t4 146.853
R1197 VN.n18 VN.t1 146.853
R1198 VN.n26 VN.t0 146.853
R1199 VN.n13 VN.n12 96.5656
R1200 VN.n27 VN.n26 96.5656
R1201 VN VN.n27 50.7216
R1202 VN.n6 VN.n1 50.6917
R1203 VN.n20 VN.n15 50.6917
R1204 VN.n4 VN.n3 48.0623
R1205 VN.n18 VN.n17 48.0623
R1206 VN.n10 VN.n1 30.2951
R1207 VN.n24 VN.n15 30.2951
R1208 VN.n5 VN.n4 24.4675
R1209 VN.n6 VN.n5 24.4675
R1210 VN.n11 VN.n10 24.4675
R1211 VN.n20 VN.n19 24.4675
R1212 VN.n19 VN.n18 24.4675
R1213 VN.n25 VN.n24 24.4675
R1214 VN.n12 VN.n11 14.1914
R1215 VN.n26 VN.n25 14.1914
R1216 VN.n17 VN.n16 6.56002
R1217 VN.n3 VN.n2 6.56002
R1218 VN.n27 VN.n14 0.278367
R1219 VN.n13 VN.n0 0.278367
R1220 VN.n23 VN.n14 0.189894
R1221 VN.n23 VN.n22 0.189894
R1222 VN.n22 VN.n21 0.189894
R1223 VN.n21 VN.n16 0.189894
R1224 VN.n7 VN.n2 0.189894
R1225 VN.n8 VN.n7 0.189894
R1226 VN.n9 VN.n8 0.189894
R1227 VN.n9 VN.n0 0.189894
R1228 VN VN.n13 0.153454
R1229 VTAIL.n7 VTAIL.t9 55.8009
R1230 VTAIL.n11 VTAIL.t10 55.8006
R1231 VTAIL.n2 VTAIL.t5 55.8006
R1232 VTAIL.n10 VTAIL.t3 55.8006
R1233 VTAIL.n9 VTAIL.n8 53.6324
R1234 VTAIL.n6 VTAIL.n5 53.6324
R1235 VTAIL.n1 VTAIL.n0 53.6322
R1236 VTAIL.n4 VTAIL.n3 53.6322
R1237 VTAIL.n6 VTAIL.n4 30.0996
R1238 VTAIL.n11 VTAIL.n10 27.6945
R1239 VTAIL.n7 VTAIL.n6 2.40567
R1240 VTAIL.n10 VTAIL.n9 2.40567
R1241 VTAIL.n4 VTAIL.n2 2.40567
R1242 VTAIL.n0 VTAIL.t11 2.16895
R1243 VTAIL.n0 VTAIL.t8 2.16895
R1244 VTAIL.n3 VTAIL.t1 2.16895
R1245 VTAIL.n3 VTAIL.t4 2.16895
R1246 VTAIL.n8 VTAIL.t2 2.16895
R1247 VTAIL.n8 VTAIL.t0 2.16895
R1248 VTAIL.n5 VTAIL.t6 2.16895
R1249 VTAIL.n5 VTAIL.t7 2.16895
R1250 VTAIL VTAIL.n11 1.74619
R1251 VTAIL.n9 VTAIL.n7 1.67291
R1252 VTAIL.n2 VTAIL.n1 1.67291
R1253 VTAIL VTAIL.n1 0.659983
R1254 VDD2.n1 VDD2.t0 74.2279
R1255 VDD2.n2 VDD2.t5 72.4797
R1256 VDD2.n1 VDD2.n0 70.8569
R1257 VDD2 VDD2.n3 70.8541
R1258 VDD2.n2 VDD2.n1 44.4545
R1259 VDD2.n3 VDD2.t4 2.16895
R1260 VDD2.n3 VDD2.t2 2.16895
R1261 VDD2.n0 VDD2.t3 2.16895
R1262 VDD2.n0 VDD2.t1 2.16895
R1263 VDD2 VDD2.n2 1.86257
R1264 VP.n9 VP.t2 181.786
R1265 VP.n11 VP.n8 161.3
R1266 VP.n13 VP.n12 161.3
R1267 VP.n14 VP.n7 161.3
R1268 VP.n16 VP.n15 161.3
R1269 VP.n17 VP.n6 161.3
R1270 VP.n37 VP.n0 161.3
R1271 VP.n36 VP.n35 161.3
R1272 VP.n34 VP.n1 161.3
R1273 VP.n33 VP.n32 161.3
R1274 VP.n31 VP.n2 161.3
R1275 VP.n30 VP.n29 161.3
R1276 VP.n28 VP.n3 161.3
R1277 VP.n27 VP.n26 161.3
R1278 VP.n25 VP.n4 161.3
R1279 VP.n24 VP.n23 161.3
R1280 VP.n22 VP.n5 161.3
R1281 VP.n30 VP.t1 146.853
R1282 VP.n20 VP.t4 146.853
R1283 VP.n38 VP.t0 146.853
R1284 VP.n10 VP.t5 146.853
R1285 VP.n18 VP.t3 146.853
R1286 VP.n21 VP.n20 96.5656
R1287 VP.n39 VP.n38 96.5656
R1288 VP.n19 VP.n18 96.5656
R1289 VP.n26 VP.n25 50.6917
R1290 VP.n32 VP.n1 50.6917
R1291 VP.n12 VP.n7 50.6917
R1292 VP.n21 VP.n19 50.4428
R1293 VP.n10 VP.n9 48.0623
R1294 VP.n25 VP.n24 30.2951
R1295 VP.n36 VP.n1 30.2951
R1296 VP.n16 VP.n7 30.2951
R1297 VP.n24 VP.n5 24.4675
R1298 VP.n26 VP.n3 24.4675
R1299 VP.n30 VP.n3 24.4675
R1300 VP.n31 VP.n30 24.4675
R1301 VP.n32 VP.n31 24.4675
R1302 VP.n37 VP.n36 24.4675
R1303 VP.n17 VP.n16 24.4675
R1304 VP.n11 VP.n10 24.4675
R1305 VP.n12 VP.n11 24.4675
R1306 VP.n20 VP.n5 14.1914
R1307 VP.n38 VP.n37 14.1914
R1308 VP.n18 VP.n17 14.1914
R1309 VP.n9 VP.n8 6.56002
R1310 VP.n19 VP.n6 0.278367
R1311 VP.n22 VP.n21 0.278367
R1312 VP.n39 VP.n0 0.278367
R1313 VP.n13 VP.n8 0.189894
R1314 VP.n14 VP.n13 0.189894
R1315 VP.n15 VP.n14 0.189894
R1316 VP.n15 VP.n6 0.189894
R1317 VP.n23 VP.n22 0.189894
R1318 VP.n23 VP.n4 0.189894
R1319 VP.n27 VP.n4 0.189894
R1320 VP.n28 VP.n27 0.189894
R1321 VP.n29 VP.n28 0.189894
R1322 VP.n29 VP.n2 0.189894
R1323 VP.n33 VP.n2 0.189894
R1324 VP.n34 VP.n33 0.189894
R1325 VP.n35 VP.n34 0.189894
R1326 VP.n35 VP.n0 0.189894
R1327 VP VP.n39 0.153454
R1328 VDD1 VDD1.t3 74.3417
R1329 VDD1.n1 VDD1.t1 74.2279
R1330 VDD1.n1 VDD1.n0 70.8569
R1331 VDD1.n3 VDD1.n2 70.311
R1332 VDD1.n3 VDD1.n1 46.2401
R1333 VDD1.n2 VDD1.t0 2.16895
R1334 VDD1.n2 VDD1.t2 2.16895
R1335 VDD1.n0 VDD1.t4 2.16895
R1336 VDD1.n0 VDD1.t5 2.16895
R1337 VDD1 VDD1.n3 0.543603
C0 VDD2 w_n3202_n3966# 2.54588f
C1 VDD2 VTAIL 8.867009f
C2 VDD2 VDD1 1.35258f
C3 VDD2 VN 8.21529f
C4 VDD2 VP 0.44667f
C5 VTAIL w_n3202_n3966# 3.38209f
C6 VDD1 w_n3202_n3966# 2.46528f
C7 VDD2 B 2.36174f
C8 VN w_n3202_n3966# 6.08323f
C9 VP w_n3202_n3966# 6.49682f
C10 VTAIL VDD1 8.818f
C11 VN VTAIL 8.207299f
C12 VTAIL VP 8.22164f
C13 VN VDD1 0.150512f
C14 VDD1 VP 8.507679f
C15 VN VP 7.34254f
C16 B w_n3202_n3966# 10.321f
C17 B VTAIL 4.29956f
C18 B VDD1 2.29101f
C19 B VN 1.17271f
C20 B VP 1.86253f
C21 VDD2 VSUBS 1.962347f
C22 VDD1 VSUBS 2.436224f
C23 VTAIL VSUBS 1.269354f
C24 VN VSUBS 5.8163f
C25 VP VSUBS 2.936023f
C26 B VSUBS 4.753628f
C27 w_n3202_n3966# VSUBS 0.155732p
C28 VDD1.t3 VSUBS 3.44483f
C29 VDD1.t1 VSUBS 3.4434f
C30 VDD1.t4 VSUBS 0.324899f
C31 VDD1.t5 VSUBS 0.324899f
C32 VDD1.n0 VSUBS 2.64051f
C33 VDD1.n1 VSUBS 4.0783f
C34 VDD1.t0 VSUBS 0.324899f
C35 VDD1.t2 VSUBS 0.324899f
C36 VDD1.n2 VSUBS 2.63434f
C37 VDD1.n3 VSUBS 3.56832f
C38 VP.n0 VSUBS 0.039872f
C39 VP.t0 VSUBS 3.05586f
C40 VP.n1 VSUBS 0.029022f
C41 VP.n2 VSUBS 0.030243f
C42 VP.t1 VSUBS 3.05586f
C43 VP.n3 VSUBS 0.056365f
C44 VP.n4 VSUBS 0.030243f
C45 VP.n5 VSUBS 0.044677f
C46 VP.n6 VSUBS 0.039872f
C47 VP.t3 VSUBS 3.05586f
C48 VP.n7 VSUBS 0.029022f
C49 VP.n8 VSUBS 0.287894f
C50 VP.t5 VSUBS 3.05586f
C51 VP.t2 VSUBS 3.29685f
C52 VP.n9 VSUBS 1.12307f
C53 VP.n10 VSUBS 1.17042f
C54 VP.n11 VSUBS 0.056365f
C55 VP.n12 VSUBS 0.055213f
C56 VP.n13 VSUBS 0.030243f
C57 VP.n14 VSUBS 0.030243f
C58 VP.n15 VSUBS 0.030243f
C59 VP.n16 VSUBS 0.060433f
C60 VP.n17 VSUBS 0.044677f
C61 VP.n18 VSUBS 1.17261f
C62 VP.n19 VSUBS 1.70033f
C63 VP.t4 VSUBS 3.05586f
C64 VP.n20 VSUBS 1.17261f
C65 VP.n21 VSUBS 1.72189f
C66 VP.n22 VSUBS 0.039872f
C67 VP.n23 VSUBS 0.030243f
C68 VP.n24 VSUBS 0.060433f
C69 VP.n25 VSUBS 0.029022f
C70 VP.n26 VSUBS 0.055213f
C71 VP.n27 VSUBS 0.030243f
C72 VP.n28 VSUBS 0.030243f
C73 VP.n29 VSUBS 0.030243f
C74 VP.n30 VSUBS 1.09815f
C75 VP.n31 VSUBS 0.056365f
C76 VP.n32 VSUBS 0.055213f
C77 VP.n33 VSUBS 0.030243f
C78 VP.n34 VSUBS 0.030243f
C79 VP.n35 VSUBS 0.030243f
C80 VP.n36 VSUBS 0.060433f
C81 VP.n37 VSUBS 0.044677f
C82 VP.n38 VSUBS 1.17261f
C83 VP.n39 VSUBS 0.04452f
C84 VDD2.t0 VSUBS 3.44361f
C85 VDD2.t3 VSUBS 0.324919f
C86 VDD2.t1 VSUBS 0.324919f
C87 VDD2.n0 VSUBS 2.64067f
C88 VDD2.n1 VSUBS 3.94408f
C89 VDD2.t5 VSUBS 3.42504f
C90 VDD2.n2 VSUBS 3.60128f
C91 VDD2.t4 VSUBS 0.324919f
C92 VDD2.t2 VSUBS 0.324919f
C93 VDD2.n3 VSUBS 2.64062f
C94 VTAIL.t11 VSUBS 0.33318f
C95 VTAIL.t8 VSUBS 0.33318f
C96 VTAIL.n0 VSUBS 2.53511f
C97 VTAIL.n1 VSUBS 0.879828f
C98 VTAIL.t5 VSUBS 3.32291f
C99 VTAIL.n2 VSUBS 1.15892f
C100 VTAIL.t1 VSUBS 0.33318f
C101 VTAIL.t4 VSUBS 0.33318f
C102 VTAIL.n3 VSUBS 2.53511f
C103 VTAIL.n4 VSUBS 2.87569f
C104 VTAIL.t6 VSUBS 0.33318f
C105 VTAIL.t7 VSUBS 0.33318f
C106 VTAIL.n5 VSUBS 2.53512f
C107 VTAIL.n6 VSUBS 2.87568f
C108 VTAIL.t9 VSUBS 3.32291f
C109 VTAIL.n7 VSUBS 1.15892f
C110 VTAIL.t2 VSUBS 0.33318f
C111 VTAIL.t0 VSUBS 0.33318f
C112 VTAIL.n8 VSUBS 2.53512f
C113 VTAIL.n9 VSUBS 1.03804f
C114 VTAIL.t3 VSUBS 3.32291f
C115 VTAIL.n10 VSUBS 2.77859f
C116 VTAIL.t10 VSUBS 3.32291f
C117 VTAIL.n11 VSUBS 2.71882f
C118 VN.n0 VSUBS 0.038903f
C119 VN.t4 VSUBS 2.98157f
C120 VN.n1 VSUBS 0.028317f
C121 VN.n2 VSUBS 0.280895f
C122 VN.t2 VSUBS 2.98157f
C123 VN.t5 VSUBS 3.2167f
C124 VN.n3 VSUBS 1.09577f
C125 VN.n4 VSUBS 1.14197f
C126 VN.n5 VSUBS 0.054995f
C127 VN.n6 VSUBS 0.053871f
C128 VN.n7 VSUBS 0.029508f
C129 VN.n8 VSUBS 0.029508f
C130 VN.n9 VSUBS 0.029508f
C131 VN.n10 VSUBS 0.058964f
C132 VN.n11 VSUBS 0.043591f
C133 VN.n12 VSUBS 1.1441f
C134 VN.n13 VSUBS 0.043438f
C135 VN.n14 VSUBS 0.038903f
C136 VN.t0 VSUBS 2.98157f
C137 VN.n15 VSUBS 0.028317f
C138 VN.n16 VSUBS 0.280895f
C139 VN.t1 VSUBS 2.98157f
C140 VN.t3 VSUBS 3.2167f
C141 VN.n17 VSUBS 1.09577f
C142 VN.n18 VSUBS 1.14197f
C143 VN.n19 VSUBS 0.054995f
C144 VN.n20 VSUBS 0.053871f
C145 VN.n21 VSUBS 0.029508f
C146 VN.n22 VSUBS 0.029508f
C147 VN.n23 VSUBS 0.029508f
C148 VN.n24 VSUBS 0.058964f
C149 VN.n25 VSUBS 0.043591f
C150 VN.n26 VSUBS 1.1441f
C151 VN.n27 VSUBS 1.67483f
C152 B.n0 VSUBS 0.004835f
C153 B.n1 VSUBS 0.004835f
C154 B.n2 VSUBS 0.007647f
C155 B.n3 VSUBS 0.007647f
C156 B.n4 VSUBS 0.007647f
C157 B.n5 VSUBS 0.007647f
C158 B.n6 VSUBS 0.007647f
C159 B.n7 VSUBS 0.007647f
C160 B.n8 VSUBS 0.007647f
C161 B.n9 VSUBS 0.007647f
C162 B.n10 VSUBS 0.007647f
C163 B.n11 VSUBS 0.007647f
C164 B.n12 VSUBS 0.007647f
C165 B.n13 VSUBS 0.007647f
C166 B.n14 VSUBS 0.007647f
C167 B.n15 VSUBS 0.007647f
C168 B.n16 VSUBS 0.007647f
C169 B.n17 VSUBS 0.007647f
C170 B.n18 VSUBS 0.007647f
C171 B.n19 VSUBS 0.007647f
C172 B.n20 VSUBS 0.007647f
C173 B.n21 VSUBS 0.007647f
C174 B.n22 VSUBS 0.018106f
C175 B.n23 VSUBS 0.007647f
C176 B.n24 VSUBS 0.007647f
C177 B.n25 VSUBS 0.007647f
C178 B.n26 VSUBS 0.007647f
C179 B.n27 VSUBS 0.007647f
C180 B.n28 VSUBS 0.007647f
C181 B.n29 VSUBS 0.007647f
C182 B.n30 VSUBS 0.007647f
C183 B.n31 VSUBS 0.007647f
C184 B.n32 VSUBS 0.007647f
C185 B.n33 VSUBS 0.007647f
C186 B.n34 VSUBS 0.007647f
C187 B.n35 VSUBS 0.007647f
C188 B.n36 VSUBS 0.007647f
C189 B.n37 VSUBS 0.007647f
C190 B.n38 VSUBS 0.007647f
C191 B.n39 VSUBS 0.007647f
C192 B.n40 VSUBS 0.007647f
C193 B.n41 VSUBS 0.007647f
C194 B.n42 VSUBS 0.007647f
C195 B.n43 VSUBS 0.007647f
C196 B.n44 VSUBS 0.007647f
C197 B.n45 VSUBS 0.007647f
C198 B.n46 VSUBS 0.007647f
C199 B.n47 VSUBS 0.007647f
C200 B.t11 VSUBS 0.545034f
C201 B.t10 VSUBS 0.567559f
C202 B.t9 VSUBS 1.80158f
C203 B.n48 VSUBS 0.296968f
C204 B.n49 VSUBS 0.078028f
C205 B.n50 VSUBS 0.007647f
C206 B.n51 VSUBS 0.007647f
C207 B.n52 VSUBS 0.007647f
C208 B.n53 VSUBS 0.007647f
C209 B.n54 VSUBS 0.004273f
C210 B.n55 VSUBS 0.007647f
C211 B.t5 VSUBS 0.545018f
C212 B.t4 VSUBS 0.567546f
C213 B.t3 VSUBS 1.80158f
C214 B.n56 VSUBS 0.296981f
C215 B.n57 VSUBS 0.078044f
C216 B.n58 VSUBS 0.017716f
C217 B.n59 VSUBS 0.007647f
C218 B.n60 VSUBS 0.007647f
C219 B.n61 VSUBS 0.007647f
C220 B.n62 VSUBS 0.007647f
C221 B.n63 VSUBS 0.007647f
C222 B.n64 VSUBS 0.007647f
C223 B.n65 VSUBS 0.007647f
C224 B.n66 VSUBS 0.007647f
C225 B.n67 VSUBS 0.007647f
C226 B.n68 VSUBS 0.007647f
C227 B.n69 VSUBS 0.007647f
C228 B.n70 VSUBS 0.007647f
C229 B.n71 VSUBS 0.007647f
C230 B.n72 VSUBS 0.007647f
C231 B.n73 VSUBS 0.007647f
C232 B.n74 VSUBS 0.007647f
C233 B.n75 VSUBS 0.007647f
C234 B.n76 VSUBS 0.007647f
C235 B.n77 VSUBS 0.007647f
C236 B.n78 VSUBS 0.007647f
C237 B.n79 VSUBS 0.007647f
C238 B.n80 VSUBS 0.007647f
C239 B.n81 VSUBS 0.007647f
C240 B.n82 VSUBS 0.018552f
C241 B.n83 VSUBS 0.007647f
C242 B.n84 VSUBS 0.007647f
C243 B.n85 VSUBS 0.007647f
C244 B.n86 VSUBS 0.007647f
C245 B.n87 VSUBS 0.007647f
C246 B.n88 VSUBS 0.007647f
C247 B.n89 VSUBS 0.007647f
C248 B.n90 VSUBS 0.007647f
C249 B.n91 VSUBS 0.007647f
C250 B.n92 VSUBS 0.007647f
C251 B.n93 VSUBS 0.007647f
C252 B.n94 VSUBS 0.007647f
C253 B.n95 VSUBS 0.007647f
C254 B.n96 VSUBS 0.007647f
C255 B.n97 VSUBS 0.007647f
C256 B.n98 VSUBS 0.007647f
C257 B.n99 VSUBS 0.007647f
C258 B.n100 VSUBS 0.007647f
C259 B.n101 VSUBS 0.007647f
C260 B.n102 VSUBS 0.007647f
C261 B.n103 VSUBS 0.007647f
C262 B.n104 VSUBS 0.007647f
C263 B.n105 VSUBS 0.007647f
C264 B.n106 VSUBS 0.007647f
C265 B.n107 VSUBS 0.007647f
C266 B.n108 VSUBS 0.007647f
C267 B.n109 VSUBS 0.007647f
C268 B.n110 VSUBS 0.007647f
C269 B.n111 VSUBS 0.007647f
C270 B.n112 VSUBS 0.007647f
C271 B.n113 VSUBS 0.007647f
C272 B.n114 VSUBS 0.007647f
C273 B.n115 VSUBS 0.007647f
C274 B.n116 VSUBS 0.007647f
C275 B.n117 VSUBS 0.007647f
C276 B.n118 VSUBS 0.007647f
C277 B.n119 VSUBS 0.007647f
C278 B.n120 VSUBS 0.007647f
C279 B.n121 VSUBS 0.007647f
C280 B.n122 VSUBS 0.007647f
C281 B.n123 VSUBS 0.007647f
C282 B.n124 VSUBS 0.018552f
C283 B.n125 VSUBS 0.007647f
C284 B.n126 VSUBS 0.007647f
C285 B.n127 VSUBS 0.007647f
C286 B.n128 VSUBS 0.007647f
C287 B.n129 VSUBS 0.007647f
C288 B.n130 VSUBS 0.007647f
C289 B.n131 VSUBS 0.007647f
C290 B.n132 VSUBS 0.007647f
C291 B.n133 VSUBS 0.007647f
C292 B.n134 VSUBS 0.007647f
C293 B.n135 VSUBS 0.007647f
C294 B.n136 VSUBS 0.007647f
C295 B.n137 VSUBS 0.007647f
C296 B.n138 VSUBS 0.007647f
C297 B.n139 VSUBS 0.007647f
C298 B.n140 VSUBS 0.007647f
C299 B.n141 VSUBS 0.007647f
C300 B.n142 VSUBS 0.007647f
C301 B.n143 VSUBS 0.007647f
C302 B.n144 VSUBS 0.007647f
C303 B.n145 VSUBS 0.007647f
C304 B.n146 VSUBS 0.007647f
C305 B.n147 VSUBS 0.007647f
C306 B.n148 VSUBS 0.007647f
C307 B.t1 VSUBS 0.545018f
C308 B.t2 VSUBS 0.567546f
C309 B.t0 VSUBS 1.80158f
C310 B.n149 VSUBS 0.296981f
C311 B.n150 VSUBS 0.078044f
C312 B.n151 VSUBS 0.017716f
C313 B.n152 VSUBS 0.007647f
C314 B.n153 VSUBS 0.007647f
C315 B.n154 VSUBS 0.007647f
C316 B.n155 VSUBS 0.007647f
C317 B.n156 VSUBS 0.007647f
C318 B.t7 VSUBS 0.545034f
C319 B.t8 VSUBS 0.567559f
C320 B.t6 VSUBS 1.80158f
C321 B.n157 VSUBS 0.296968f
C322 B.n158 VSUBS 0.078028f
C323 B.n159 VSUBS 0.007647f
C324 B.n160 VSUBS 0.007647f
C325 B.n161 VSUBS 0.007647f
C326 B.n162 VSUBS 0.007647f
C327 B.n163 VSUBS 0.007647f
C328 B.n164 VSUBS 0.007647f
C329 B.n165 VSUBS 0.007647f
C330 B.n166 VSUBS 0.007647f
C331 B.n167 VSUBS 0.007647f
C332 B.n168 VSUBS 0.007647f
C333 B.n169 VSUBS 0.007647f
C334 B.n170 VSUBS 0.007647f
C335 B.n171 VSUBS 0.007647f
C336 B.n172 VSUBS 0.007647f
C337 B.n173 VSUBS 0.007647f
C338 B.n174 VSUBS 0.007647f
C339 B.n175 VSUBS 0.007647f
C340 B.n176 VSUBS 0.007647f
C341 B.n177 VSUBS 0.007647f
C342 B.n178 VSUBS 0.007647f
C343 B.n179 VSUBS 0.007647f
C344 B.n180 VSUBS 0.007647f
C345 B.n181 VSUBS 0.007647f
C346 B.n182 VSUBS 0.007647f
C347 B.n183 VSUBS 0.018552f
C348 B.n184 VSUBS 0.007647f
C349 B.n185 VSUBS 0.007647f
C350 B.n186 VSUBS 0.007647f
C351 B.n187 VSUBS 0.007647f
C352 B.n188 VSUBS 0.007647f
C353 B.n189 VSUBS 0.007647f
C354 B.n190 VSUBS 0.007647f
C355 B.n191 VSUBS 0.007647f
C356 B.n192 VSUBS 0.007647f
C357 B.n193 VSUBS 0.007647f
C358 B.n194 VSUBS 0.007647f
C359 B.n195 VSUBS 0.007647f
C360 B.n196 VSUBS 0.007647f
C361 B.n197 VSUBS 0.007647f
C362 B.n198 VSUBS 0.007647f
C363 B.n199 VSUBS 0.007647f
C364 B.n200 VSUBS 0.007647f
C365 B.n201 VSUBS 0.007647f
C366 B.n202 VSUBS 0.007647f
C367 B.n203 VSUBS 0.007647f
C368 B.n204 VSUBS 0.007647f
C369 B.n205 VSUBS 0.007647f
C370 B.n206 VSUBS 0.007647f
C371 B.n207 VSUBS 0.007647f
C372 B.n208 VSUBS 0.007647f
C373 B.n209 VSUBS 0.007647f
C374 B.n210 VSUBS 0.007647f
C375 B.n211 VSUBS 0.007647f
C376 B.n212 VSUBS 0.007647f
C377 B.n213 VSUBS 0.007647f
C378 B.n214 VSUBS 0.007647f
C379 B.n215 VSUBS 0.007647f
C380 B.n216 VSUBS 0.007647f
C381 B.n217 VSUBS 0.007647f
C382 B.n218 VSUBS 0.007647f
C383 B.n219 VSUBS 0.007647f
C384 B.n220 VSUBS 0.007647f
C385 B.n221 VSUBS 0.007647f
C386 B.n222 VSUBS 0.007647f
C387 B.n223 VSUBS 0.007647f
C388 B.n224 VSUBS 0.007647f
C389 B.n225 VSUBS 0.007647f
C390 B.n226 VSUBS 0.007647f
C391 B.n227 VSUBS 0.007647f
C392 B.n228 VSUBS 0.007647f
C393 B.n229 VSUBS 0.007647f
C394 B.n230 VSUBS 0.007647f
C395 B.n231 VSUBS 0.007647f
C396 B.n232 VSUBS 0.007647f
C397 B.n233 VSUBS 0.007647f
C398 B.n234 VSUBS 0.007647f
C399 B.n235 VSUBS 0.007647f
C400 B.n236 VSUBS 0.007647f
C401 B.n237 VSUBS 0.007647f
C402 B.n238 VSUBS 0.007647f
C403 B.n239 VSUBS 0.007647f
C404 B.n240 VSUBS 0.007647f
C405 B.n241 VSUBS 0.007647f
C406 B.n242 VSUBS 0.007647f
C407 B.n243 VSUBS 0.007647f
C408 B.n244 VSUBS 0.007647f
C409 B.n245 VSUBS 0.007647f
C410 B.n246 VSUBS 0.007647f
C411 B.n247 VSUBS 0.007647f
C412 B.n248 VSUBS 0.007647f
C413 B.n249 VSUBS 0.007647f
C414 B.n250 VSUBS 0.007647f
C415 B.n251 VSUBS 0.007647f
C416 B.n252 VSUBS 0.007647f
C417 B.n253 VSUBS 0.007647f
C418 B.n254 VSUBS 0.007647f
C419 B.n255 VSUBS 0.007647f
C420 B.n256 VSUBS 0.007647f
C421 B.n257 VSUBS 0.007647f
C422 B.n258 VSUBS 0.007647f
C423 B.n259 VSUBS 0.007647f
C424 B.n260 VSUBS 0.007647f
C425 B.n261 VSUBS 0.007647f
C426 B.n262 VSUBS 0.018106f
C427 B.n263 VSUBS 0.018106f
C428 B.n264 VSUBS 0.018552f
C429 B.n265 VSUBS 0.007647f
C430 B.n266 VSUBS 0.007647f
C431 B.n267 VSUBS 0.007647f
C432 B.n268 VSUBS 0.007647f
C433 B.n269 VSUBS 0.007647f
C434 B.n270 VSUBS 0.007647f
C435 B.n271 VSUBS 0.007647f
C436 B.n272 VSUBS 0.007647f
C437 B.n273 VSUBS 0.007647f
C438 B.n274 VSUBS 0.007647f
C439 B.n275 VSUBS 0.007647f
C440 B.n276 VSUBS 0.007647f
C441 B.n277 VSUBS 0.007647f
C442 B.n278 VSUBS 0.007647f
C443 B.n279 VSUBS 0.007647f
C444 B.n280 VSUBS 0.007647f
C445 B.n281 VSUBS 0.007647f
C446 B.n282 VSUBS 0.007647f
C447 B.n283 VSUBS 0.007647f
C448 B.n284 VSUBS 0.007647f
C449 B.n285 VSUBS 0.007647f
C450 B.n286 VSUBS 0.007647f
C451 B.n287 VSUBS 0.007647f
C452 B.n288 VSUBS 0.007647f
C453 B.n289 VSUBS 0.007647f
C454 B.n290 VSUBS 0.007647f
C455 B.n291 VSUBS 0.007647f
C456 B.n292 VSUBS 0.007647f
C457 B.n293 VSUBS 0.007647f
C458 B.n294 VSUBS 0.007647f
C459 B.n295 VSUBS 0.007647f
C460 B.n296 VSUBS 0.007647f
C461 B.n297 VSUBS 0.007647f
C462 B.n298 VSUBS 0.007647f
C463 B.n299 VSUBS 0.007647f
C464 B.n300 VSUBS 0.007647f
C465 B.n301 VSUBS 0.007647f
C466 B.n302 VSUBS 0.007647f
C467 B.n303 VSUBS 0.007647f
C468 B.n304 VSUBS 0.007647f
C469 B.n305 VSUBS 0.007647f
C470 B.n306 VSUBS 0.007647f
C471 B.n307 VSUBS 0.007647f
C472 B.n308 VSUBS 0.007647f
C473 B.n309 VSUBS 0.007647f
C474 B.n310 VSUBS 0.007647f
C475 B.n311 VSUBS 0.007647f
C476 B.n312 VSUBS 0.007647f
C477 B.n313 VSUBS 0.007647f
C478 B.n314 VSUBS 0.007647f
C479 B.n315 VSUBS 0.007647f
C480 B.n316 VSUBS 0.007647f
C481 B.n317 VSUBS 0.007647f
C482 B.n318 VSUBS 0.007647f
C483 B.n319 VSUBS 0.007647f
C484 B.n320 VSUBS 0.007647f
C485 B.n321 VSUBS 0.007647f
C486 B.n322 VSUBS 0.007647f
C487 B.n323 VSUBS 0.007647f
C488 B.n324 VSUBS 0.007647f
C489 B.n325 VSUBS 0.007647f
C490 B.n326 VSUBS 0.007647f
C491 B.n327 VSUBS 0.007647f
C492 B.n328 VSUBS 0.007647f
C493 B.n329 VSUBS 0.007647f
C494 B.n330 VSUBS 0.007647f
C495 B.n331 VSUBS 0.007647f
C496 B.n332 VSUBS 0.007647f
C497 B.n333 VSUBS 0.007647f
C498 B.n334 VSUBS 0.007647f
C499 B.n335 VSUBS 0.007647f
C500 B.n336 VSUBS 0.007647f
C501 B.n337 VSUBS 0.007647f
C502 B.n338 VSUBS 0.007197f
C503 B.n339 VSUBS 0.017716f
C504 B.n340 VSUBS 0.004273f
C505 B.n341 VSUBS 0.007647f
C506 B.n342 VSUBS 0.007647f
C507 B.n343 VSUBS 0.007647f
C508 B.n344 VSUBS 0.007647f
C509 B.n345 VSUBS 0.007647f
C510 B.n346 VSUBS 0.007647f
C511 B.n347 VSUBS 0.007647f
C512 B.n348 VSUBS 0.007647f
C513 B.n349 VSUBS 0.007647f
C514 B.n350 VSUBS 0.007647f
C515 B.n351 VSUBS 0.007647f
C516 B.n352 VSUBS 0.007647f
C517 B.n353 VSUBS 0.004273f
C518 B.n354 VSUBS 0.007647f
C519 B.n355 VSUBS 0.007647f
C520 B.n356 VSUBS 0.007197f
C521 B.n357 VSUBS 0.007647f
C522 B.n358 VSUBS 0.007647f
C523 B.n359 VSUBS 0.007647f
C524 B.n360 VSUBS 0.007647f
C525 B.n361 VSUBS 0.007647f
C526 B.n362 VSUBS 0.007647f
C527 B.n363 VSUBS 0.007647f
C528 B.n364 VSUBS 0.007647f
C529 B.n365 VSUBS 0.007647f
C530 B.n366 VSUBS 0.007647f
C531 B.n367 VSUBS 0.007647f
C532 B.n368 VSUBS 0.007647f
C533 B.n369 VSUBS 0.007647f
C534 B.n370 VSUBS 0.007647f
C535 B.n371 VSUBS 0.007647f
C536 B.n372 VSUBS 0.007647f
C537 B.n373 VSUBS 0.007647f
C538 B.n374 VSUBS 0.007647f
C539 B.n375 VSUBS 0.007647f
C540 B.n376 VSUBS 0.007647f
C541 B.n377 VSUBS 0.007647f
C542 B.n378 VSUBS 0.007647f
C543 B.n379 VSUBS 0.007647f
C544 B.n380 VSUBS 0.007647f
C545 B.n381 VSUBS 0.007647f
C546 B.n382 VSUBS 0.007647f
C547 B.n383 VSUBS 0.007647f
C548 B.n384 VSUBS 0.007647f
C549 B.n385 VSUBS 0.007647f
C550 B.n386 VSUBS 0.007647f
C551 B.n387 VSUBS 0.007647f
C552 B.n388 VSUBS 0.007647f
C553 B.n389 VSUBS 0.007647f
C554 B.n390 VSUBS 0.007647f
C555 B.n391 VSUBS 0.007647f
C556 B.n392 VSUBS 0.007647f
C557 B.n393 VSUBS 0.007647f
C558 B.n394 VSUBS 0.007647f
C559 B.n395 VSUBS 0.007647f
C560 B.n396 VSUBS 0.007647f
C561 B.n397 VSUBS 0.007647f
C562 B.n398 VSUBS 0.007647f
C563 B.n399 VSUBS 0.007647f
C564 B.n400 VSUBS 0.007647f
C565 B.n401 VSUBS 0.007647f
C566 B.n402 VSUBS 0.007647f
C567 B.n403 VSUBS 0.007647f
C568 B.n404 VSUBS 0.007647f
C569 B.n405 VSUBS 0.007647f
C570 B.n406 VSUBS 0.007647f
C571 B.n407 VSUBS 0.007647f
C572 B.n408 VSUBS 0.007647f
C573 B.n409 VSUBS 0.007647f
C574 B.n410 VSUBS 0.007647f
C575 B.n411 VSUBS 0.007647f
C576 B.n412 VSUBS 0.007647f
C577 B.n413 VSUBS 0.007647f
C578 B.n414 VSUBS 0.007647f
C579 B.n415 VSUBS 0.007647f
C580 B.n416 VSUBS 0.007647f
C581 B.n417 VSUBS 0.007647f
C582 B.n418 VSUBS 0.007647f
C583 B.n419 VSUBS 0.007647f
C584 B.n420 VSUBS 0.007647f
C585 B.n421 VSUBS 0.007647f
C586 B.n422 VSUBS 0.007647f
C587 B.n423 VSUBS 0.007647f
C588 B.n424 VSUBS 0.007647f
C589 B.n425 VSUBS 0.007647f
C590 B.n426 VSUBS 0.007647f
C591 B.n427 VSUBS 0.007647f
C592 B.n428 VSUBS 0.007647f
C593 B.n429 VSUBS 0.018552f
C594 B.n430 VSUBS 0.018106f
C595 B.n431 VSUBS 0.018106f
C596 B.n432 VSUBS 0.007647f
C597 B.n433 VSUBS 0.007647f
C598 B.n434 VSUBS 0.007647f
C599 B.n435 VSUBS 0.007647f
C600 B.n436 VSUBS 0.007647f
C601 B.n437 VSUBS 0.007647f
C602 B.n438 VSUBS 0.007647f
C603 B.n439 VSUBS 0.007647f
C604 B.n440 VSUBS 0.007647f
C605 B.n441 VSUBS 0.007647f
C606 B.n442 VSUBS 0.007647f
C607 B.n443 VSUBS 0.007647f
C608 B.n444 VSUBS 0.007647f
C609 B.n445 VSUBS 0.007647f
C610 B.n446 VSUBS 0.007647f
C611 B.n447 VSUBS 0.007647f
C612 B.n448 VSUBS 0.007647f
C613 B.n449 VSUBS 0.007647f
C614 B.n450 VSUBS 0.007647f
C615 B.n451 VSUBS 0.007647f
C616 B.n452 VSUBS 0.007647f
C617 B.n453 VSUBS 0.007647f
C618 B.n454 VSUBS 0.007647f
C619 B.n455 VSUBS 0.007647f
C620 B.n456 VSUBS 0.007647f
C621 B.n457 VSUBS 0.007647f
C622 B.n458 VSUBS 0.007647f
C623 B.n459 VSUBS 0.007647f
C624 B.n460 VSUBS 0.007647f
C625 B.n461 VSUBS 0.007647f
C626 B.n462 VSUBS 0.007647f
C627 B.n463 VSUBS 0.007647f
C628 B.n464 VSUBS 0.007647f
C629 B.n465 VSUBS 0.007647f
C630 B.n466 VSUBS 0.007647f
C631 B.n467 VSUBS 0.007647f
C632 B.n468 VSUBS 0.007647f
C633 B.n469 VSUBS 0.007647f
C634 B.n470 VSUBS 0.007647f
C635 B.n471 VSUBS 0.007647f
C636 B.n472 VSUBS 0.007647f
C637 B.n473 VSUBS 0.007647f
C638 B.n474 VSUBS 0.007647f
C639 B.n475 VSUBS 0.007647f
C640 B.n476 VSUBS 0.007647f
C641 B.n477 VSUBS 0.007647f
C642 B.n478 VSUBS 0.007647f
C643 B.n479 VSUBS 0.007647f
C644 B.n480 VSUBS 0.007647f
C645 B.n481 VSUBS 0.007647f
C646 B.n482 VSUBS 0.007647f
C647 B.n483 VSUBS 0.007647f
C648 B.n484 VSUBS 0.007647f
C649 B.n485 VSUBS 0.007647f
C650 B.n486 VSUBS 0.007647f
C651 B.n487 VSUBS 0.007647f
C652 B.n488 VSUBS 0.007647f
C653 B.n489 VSUBS 0.007647f
C654 B.n490 VSUBS 0.007647f
C655 B.n491 VSUBS 0.007647f
C656 B.n492 VSUBS 0.007647f
C657 B.n493 VSUBS 0.007647f
C658 B.n494 VSUBS 0.007647f
C659 B.n495 VSUBS 0.007647f
C660 B.n496 VSUBS 0.007647f
C661 B.n497 VSUBS 0.007647f
C662 B.n498 VSUBS 0.007647f
C663 B.n499 VSUBS 0.007647f
C664 B.n500 VSUBS 0.007647f
C665 B.n501 VSUBS 0.007647f
C666 B.n502 VSUBS 0.007647f
C667 B.n503 VSUBS 0.007647f
C668 B.n504 VSUBS 0.007647f
C669 B.n505 VSUBS 0.007647f
C670 B.n506 VSUBS 0.007647f
C671 B.n507 VSUBS 0.007647f
C672 B.n508 VSUBS 0.007647f
C673 B.n509 VSUBS 0.007647f
C674 B.n510 VSUBS 0.007647f
C675 B.n511 VSUBS 0.007647f
C676 B.n512 VSUBS 0.007647f
C677 B.n513 VSUBS 0.007647f
C678 B.n514 VSUBS 0.007647f
C679 B.n515 VSUBS 0.007647f
C680 B.n516 VSUBS 0.007647f
C681 B.n517 VSUBS 0.007647f
C682 B.n518 VSUBS 0.007647f
C683 B.n519 VSUBS 0.007647f
C684 B.n520 VSUBS 0.007647f
C685 B.n521 VSUBS 0.007647f
C686 B.n522 VSUBS 0.007647f
C687 B.n523 VSUBS 0.007647f
C688 B.n524 VSUBS 0.007647f
C689 B.n525 VSUBS 0.007647f
C690 B.n526 VSUBS 0.007647f
C691 B.n527 VSUBS 0.007647f
C692 B.n528 VSUBS 0.007647f
C693 B.n529 VSUBS 0.007647f
C694 B.n530 VSUBS 0.007647f
C695 B.n531 VSUBS 0.007647f
C696 B.n532 VSUBS 0.007647f
C697 B.n533 VSUBS 0.007647f
C698 B.n534 VSUBS 0.007647f
C699 B.n535 VSUBS 0.007647f
C700 B.n536 VSUBS 0.007647f
C701 B.n537 VSUBS 0.007647f
C702 B.n538 VSUBS 0.007647f
C703 B.n539 VSUBS 0.007647f
C704 B.n540 VSUBS 0.007647f
C705 B.n541 VSUBS 0.007647f
C706 B.n542 VSUBS 0.007647f
C707 B.n543 VSUBS 0.007647f
C708 B.n544 VSUBS 0.007647f
C709 B.n545 VSUBS 0.007647f
C710 B.n546 VSUBS 0.007647f
C711 B.n547 VSUBS 0.007647f
C712 B.n548 VSUBS 0.007647f
C713 B.n549 VSUBS 0.007647f
C714 B.n550 VSUBS 0.007647f
C715 B.n551 VSUBS 0.007647f
C716 B.n552 VSUBS 0.007647f
C717 B.n553 VSUBS 0.018106f
C718 B.n554 VSUBS 0.018977f
C719 B.n555 VSUBS 0.017681f
C720 B.n556 VSUBS 0.007647f
C721 B.n557 VSUBS 0.007647f
C722 B.n558 VSUBS 0.007647f
C723 B.n559 VSUBS 0.007647f
C724 B.n560 VSUBS 0.007647f
C725 B.n561 VSUBS 0.007647f
C726 B.n562 VSUBS 0.007647f
C727 B.n563 VSUBS 0.007647f
C728 B.n564 VSUBS 0.007647f
C729 B.n565 VSUBS 0.007647f
C730 B.n566 VSUBS 0.007647f
C731 B.n567 VSUBS 0.007647f
C732 B.n568 VSUBS 0.007647f
C733 B.n569 VSUBS 0.007647f
C734 B.n570 VSUBS 0.007647f
C735 B.n571 VSUBS 0.007647f
C736 B.n572 VSUBS 0.007647f
C737 B.n573 VSUBS 0.007647f
C738 B.n574 VSUBS 0.007647f
C739 B.n575 VSUBS 0.007647f
C740 B.n576 VSUBS 0.007647f
C741 B.n577 VSUBS 0.007647f
C742 B.n578 VSUBS 0.007647f
C743 B.n579 VSUBS 0.007647f
C744 B.n580 VSUBS 0.007647f
C745 B.n581 VSUBS 0.007647f
C746 B.n582 VSUBS 0.007647f
C747 B.n583 VSUBS 0.007647f
C748 B.n584 VSUBS 0.007647f
C749 B.n585 VSUBS 0.007647f
C750 B.n586 VSUBS 0.007647f
C751 B.n587 VSUBS 0.007647f
C752 B.n588 VSUBS 0.007647f
C753 B.n589 VSUBS 0.007647f
C754 B.n590 VSUBS 0.007647f
C755 B.n591 VSUBS 0.007647f
C756 B.n592 VSUBS 0.007647f
C757 B.n593 VSUBS 0.007647f
C758 B.n594 VSUBS 0.007647f
C759 B.n595 VSUBS 0.007647f
C760 B.n596 VSUBS 0.007647f
C761 B.n597 VSUBS 0.007647f
C762 B.n598 VSUBS 0.007647f
C763 B.n599 VSUBS 0.007647f
C764 B.n600 VSUBS 0.007647f
C765 B.n601 VSUBS 0.007647f
C766 B.n602 VSUBS 0.007647f
C767 B.n603 VSUBS 0.007647f
C768 B.n604 VSUBS 0.007647f
C769 B.n605 VSUBS 0.007647f
C770 B.n606 VSUBS 0.007647f
C771 B.n607 VSUBS 0.007647f
C772 B.n608 VSUBS 0.007647f
C773 B.n609 VSUBS 0.007647f
C774 B.n610 VSUBS 0.007647f
C775 B.n611 VSUBS 0.007647f
C776 B.n612 VSUBS 0.007647f
C777 B.n613 VSUBS 0.007647f
C778 B.n614 VSUBS 0.007647f
C779 B.n615 VSUBS 0.007647f
C780 B.n616 VSUBS 0.007647f
C781 B.n617 VSUBS 0.007647f
C782 B.n618 VSUBS 0.007647f
C783 B.n619 VSUBS 0.007647f
C784 B.n620 VSUBS 0.007647f
C785 B.n621 VSUBS 0.007647f
C786 B.n622 VSUBS 0.007647f
C787 B.n623 VSUBS 0.007647f
C788 B.n624 VSUBS 0.007647f
C789 B.n625 VSUBS 0.007647f
C790 B.n626 VSUBS 0.007647f
C791 B.n627 VSUBS 0.007647f
C792 B.n628 VSUBS 0.007197f
C793 B.n629 VSUBS 0.007647f
C794 B.n630 VSUBS 0.007647f
C795 B.n631 VSUBS 0.007647f
C796 B.n632 VSUBS 0.007647f
C797 B.n633 VSUBS 0.007647f
C798 B.n634 VSUBS 0.007647f
C799 B.n635 VSUBS 0.007647f
C800 B.n636 VSUBS 0.007647f
C801 B.n637 VSUBS 0.007647f
C802 B.n638 VSUBS 0.007647f
C803 B.n639 VSUBS 0.007647f
C804 B.n640 VSUBS 0.007647f
C805 B.n641 VSUBS 0.007647f
C806 B.n642 VSUBS 0.007647f
C807 B.n643 VSUBS 0.007647f
C808 B.n644 VSUBS 0.004273f
C809 B.n645 VSUBS 0.017716f
C810 B.n646 VSUBS 0.007197f
C811 B.n647 VSUBS 0.007647f
C812 B.n648 VSUBS 0.007647f
C813 B.n649 VSUBS 0.007647f
C814 B.n650 VSUBS 0.007647f
C815 B.n651 VSUBS 0.007647f
C816 B.n652 VSUBS 0.007647f
C817 B.n653 VSUBS 0.007647f
C818 B.n654 VSUBS 0.007647f
C819 B.n655 VSUBS 0.007647f
C820 B.n656 VSUBS 0.007647f
C821 B.n657 VSUBS 0.007647f
C822 B.n658 VSUBS 0.007647f
C823 B.n659 VSUBS 0.007647f
C824 B.n660 VSUBS 0.007647f
C825 B.n661 VSUBS 0.007647f
C826 B.n662 VSUBS 0.007647f
C827 B.n663 VSUBS 0.007647f
C828 B.n664 VSUBS 0.007647f
C829 B.n665 VSUBS 0.007647f
C830 B.n666 VSUBS 0.007647f
C831 B.n667 VSUBS 0.007647f
C832 B.n668 VSUBS 0.007647f
C833 B.n669 VSUBS 0.007647f
C834 B.n670 VSUBS 0.007647f
C835 B.n671 VSUBS 0.007647f
C836 B.n672 VSUBS 0.007647f
C837 B.n673 VSUBS 0.007647f
C838 B.n674 VSUBS 0.007647f
C839 B.n675 VSUBS 0.007647f
C840 B.n676 VSUBS 0.007647f
C841 B.n677 VSUBS 0.007647f
C842 B.n678 VSUBS 0.007647f
C843 B.n679 VSUBS 0.007647f
C844 B.n680 VSUBS 0.007647f
C845 B.n681 VSUBS 0.007647f
C846 B.n682 VSUBS 0.007647f
C847 B.n683 VSUBS 0.007647f
C848 B.n684 VSUBS 0.007647f
C849 B.n685 VSUBS 0.007647f
C850 B.n686 VSUBS 0.007647f
C851 B.n687 VSUBS 0.007647f
C852 B.n688 VSUBS 0.007647f
C853 B.n689 VSUBS 0.007647f
C854 B.n690 VSUBS 0.007647f
C855 B.n691 VSUBS 0.007647f
C856 B.n692 VSUBS 0.007647f
C857 B.n693 VSUBS 0.007647f
C858 B.n694 VSUBS 0.007647f
C859 B.n695 VSUBS 0.007647f
C860 B.n696 VSUBS 0.007647f
C861 B.n697 VSUBS 0.007647f
C862 B.n698 VSUBS 0.007647f
C863 B.n699 VSUBS 0.007647f
C864 B.n700 VSUBS 0.007647f
C865 B.n701 VSUBS 0.007647f
C866 B.n702 VSUBS 0.007647f
C867 B.n703 VSUBS 0.007647f
C868 B.n704 VSUBS 0.007647f
C869 B.n705 VSUBS 0.007647f
C870 B.n706 VSUBS 0.007647f
C871 B.n707 VSUBS 0.007647f
C872 B.n708 VSUBS 0.007647f
C873 B.n709 VSUBS 0.007647f
C874 B.n710 VSUBS 0.007647f
C875 B.n711 VSUBS 0.007647f
C876 B.n712 VSUBS 0.007647f
C877 B.n713 VSUBS 0.007647f
C878 B.n714 VSUBS 0.007647f
C879 B.n715 VSUBS 0.007647f
C880 B.n716 VSUBS 0.007647f
C881 B.n717 VSUBS 0.007647f
C882 B.n718 VSUBS 0.007647f
C883 B.n719 VSUBS 0.018552f
C884 B.n720 VSUBS 0.018552f
C885 B.n721 VSUBS 0.018106f
C886 B.n722 VSUBS 0.007647f
C887 B.n723 VSUBS 0.007647f
C888 B.n724 VSUBS 0.007647f
C889 B.n725 VSUBS 0.007647f
C890 B.n726 VSUBS 0.007647f
C891 B.n727 VSUBS 0.007647f
C892 B.n728 VSUBS 0.007647f
C893 B.n729 VSUBS 0.007647f
C894 B.n730 VSUBS 0.007647f
C895 B.n731 VSUBS 0.007647f
C896 B.n732 VSUBS 0.007647f
C897 B.n733 VSUBS 0.007647f
C898 B.n734 VSUBS 0.007647f
C899 B.n735 VSUBS 0.007647f
C900 B.n736 VSUBS 0.007647f
C901 B.n737 VSUBS 0.007647f
C902 B.n738 VSUBS 0.007647f
C903 B.n739 VSUBS 0.007647f
C904 B.n740 VSUBS 0.007647f
C905 B.n741 VSUBS 0.007647f
C906 B.n742 VSUBS 0.007647f
C907 B.n743 VSUBS 0.007647f
C908 B.n744 VSUBS 0.007647f
C909 B.n745 VSUBS 0.007647f
C910 B.n746 VSUBS 0.007647f
C911 B.n747 VSUBS 0.007647f
C912 B.n748 VSUBS 0.007647f
C913 B.n749 VSUBS 0.007647f
C914 B.n750 VSUBS 0.007647f
C915 B.n751 VSUBS 0.007647f
C916 B.n752 VSUBS 0.007647f
C917 B.n753 VSUBS 0.007647f
C918 B.n754 VSUBS 0.007647f
C919 B.n755 VSUBS 0.007647f
C920 B.n756 VSUBS 0.007647f
C921 B.n757 VSUBS 0.007647f
C922 B.n758 VSUBS 0.007647f
C923 B.n759 VSUBS 0.007647f
C924 B.n760 VSUBS 0.007647f
C925 B.n761 VSUBS 0.007647f
C926 B.n762 VSUBS 0.007647f
C927 B.n763 VSUBS 0.007647f
C928 B.n764 VSUBS 0.007647f
C929 B.n765 VSUBS 0.007647f
C930 B.n766 VSUBS 0.007647f
C931 B.n767 VSUBS 0.007647f
C932 B.n768 VSUBS 0.007647f
C933 B.n769 VSUBS 0.007647f
C934 B.n770 VSUBS 0.007647f
C935 B.n771 VSUBS 0.007647f
C936 B.n772 VSUBS 0.007647f
C937 B.n773 VSUBS 0.007647f
C938 B.n774 VSUBS 0.007647f
C939 B.n775 VSUBS 0.007647f
C940 B.n776 VSUBS 0.007647f
C941 B.n777 VSUBS 0.007647f
C942 B.n778 VSUBS 0.007647f
C943 B.n779 VSUBS 0.007647f
C944 B.n780 VSUBS 0.007647f
C945 B.n781 VSUBS 0.007647f
C946 B.n782 VSUBS 0.007647f
C947 B.n783 VSUBS 0.017314f
.ends

