* NGSPICE file created from diff_pair_sample_0958.ext - technology: sky130A

.subckt diff_pair_sample_0958 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t7 VP.t0 VTAIL.t15 B.t2 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
X1 VTAIL.t1 VN.t0 VDD2.t7 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=1.49655 ps=9.4 w=9.07 l=0.28
X2 VDD1.t6 VP.t1 VTAIL.t14 B.t3 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=3.5373 ps=18.92 w=9.07 l=0.28
X3 VTAIL.t0 VN.t1 VDD2.t6 B.t0 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
X4 VDD2.t5 VN.t2 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
X5 VTAIL.t10 VP.t2 VDD1.t5 B.t1 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=1.49655 ps=9.4 w=9.07 l=0.28
X6 B.t21 B.t19 B.t20 B.t13 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=0 ps=0 w=9.07 l=0.28
X7 VDD1.t4 VP.t3 VTAIL.t9 B.t7 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
X8 B.t18 B.t16 B.t17 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=0 ps=0 w=9.07 l=0.28
X9 VTAIL.t4 VN.t3 VDD2.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=1.49655 ps=9.4 w=9.07 l=0.28
X10 VTAIL.t13 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
X11 B.t15 B.t12 B.t14 B.t13 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=0 ps=0 w=9.07 l=0.28
X12 VDD2.t3 VN.t4 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=3.5373 ps=18.92 w=9.07 l=0.28
X13 VTAIL.t12 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
X14 VTAIL.t8 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=1.49655 ps=9.4 w=9.07 l=0.28
X15 VDD2.t2 VN.t5 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=3.5373 ps=18.92 w=9.07 l=0.28
X16 VDD2.t1 VN.t6 VTAIL.t7 B.t7 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
X17 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=3.5373 pd=18.92 as=0 ps=0 w=9.07 l=0.28
X18 VDD1.t0 VP.t7 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=3.5373 ps=18.92 w=9.07 l=0.28
X19 VTAIL.t5 VN.t7 VDD2.t0 B.t5 sky130_fd_pr__nfet_01v8 ad=1.49655 pd=9.4 as=1.49655 ps=9.4 w=9.07 l=0.28
R0 VP.n17 VP.t7 917.521
R1 VP.n11 VP.t6 917.521
R2 VP.n4 VP.t2 917.521
R3 VP.n9 VP.t1 917.521
R4 VP.n16 VP.t5 893.422
R5 VP.n1 VP.t3 893.422
R6 VP.n3 VP.t0 893.422
R7 VP.n8 VP.t4 893.422
R8 VP.n5 VP.n4 161.489
R9 VP.n18 VP.n17 161.3
R10 VP.n6 VP.n5 161.3
R11 VP.n7 VP.n2 161.3
R12 VP.n10 VP.n9 161.3
R13 VP.n15 VP.n0 161.3
R14 VP.n14 VP.n13 161.3
R15 VP.n12 VP.n11 161.3
R16 VP.n15 VP.n14 73.0308
R17 VP.n7 VP.n6 73.0308
R18 VP.n11 VP.n1 64.9975
R19 VP.n17 VP.n16 64.9975
R20 VP.n4 VP.n3 64.9975
R21 VP.n9 VP.n8 64.9975
R22 VP.n12 VP.n10 37.796
R23 VP.n14 VP.n1 8.03383
R24 VP.n16 VP.n15 8.03383
R25 VP.n6 VP.n3 8.03383
R26 VP.n8 VP.n7 8.03383
R27 VP.n5 VP.n2 0.189894
R28 VP.n10 VP.n2 0.189894
R29 VP.n13 VP.n12 0.189894
R30 VP.n13 VP.n0 0.189894
R31 VP.n18 VP.n0 0.189894
R32 VP VP.n18 0.0516364
R33 VTAIL.n11 VTAIL.t10 52.3994
R34 VTAIL.n10 VTAIL.t6 52.3994
R35 VTAIL.n7 VTAIL.t4 52.3994
R36 VTAIL.n15 VTAIL.t3 52.3991
R37 VTAIL.n2 VTAIL.t1 52.3991
R38 VTAIL.n3 VTAIL.t11 52.3991
R39 VTAIL.n6 VTAIL.t8 52.3991
R40 VTAIL.n14 VTAIL.t14 52.3991
R41 VTAIL.n13 VTAIL.n12 50.2164
R42 VTAIL.n9 VTAIL.n8 50.2164
R43 VTAIL.n1 VTAIL.n0 50.2161
R44 VTAIL.n5 VTAIL.n4 50.2161
R45 VTAIL.n15 VTAIL.n14 20.7117
R46 VTAIL.n7 VTAIL.n6 20.7117
R47 VTAIL.n0 VTAIL.t2 2.18352
R48 VTAIL.n0 VTAIL.t5 2.18352
R49 VTAIL.n4 VTAIL.t9 2.18352
R50 VTAIL.n4 VTAIL.t12 2.18352
R51 VTAIL.n12 VTAIL.t15 2.18352
R52 VTAIL.n12 VTAIL.t13 2.18352
R53 VTAIL.n8 VTAIL.t7 2.18352
R54 VTAIL.n8 VTAIL.t0 2.18352
R55 VTAIL.n9 VTAIL.n7 0.526362
R56 VTAIL.n10 VTAIL.n9 0.526362
R57 VTAIL.n13 VTAIL.n11 0.526362
R58 VTAIL.n14 VTAIL.n13 0.526362
R59 VTAIL.n6 VTAIL.n5 0.526362
R60 VTAIL.n5 VTAIL.n3 0.526362
R61 VTAIL.n2 VTAIL.n1 0.526362
R62 VTAIL.n11 VTAIL.n10 0.470328
R63 VTAIL.n3 VTAIL.n2 0.470328
R64 VTAIL VTAIL.n15 0.468172
R65 VTAIL VTAIL.n1 0.0586897
R66 VDD1 VDD1.n0 67.2163
R67 VDD1.n3 VDD1.n2 67.1025
R68 VDD1.n3 VDD1.n1 67.1025
R69 VDD1.n5 VDD1.n4 66.895
R70 VDD1.n5 VDD1.n3 34.4837
R71 VDD1.n4 VDD1.t3 2.18352
R72 VDD1.n4 VDD1.t6 2.18352
R73 VDD1.n0 VDD1.t5 2.18352
R74 VDD1.n0 VDD1.t7 2.18352
R75 VDD1.n2 VDD1.t2 2.18352
R76 VDD1.n2 VDD1.t0 2.18352
R77 VDD1.n1 VDD1.t1 2.18352
R78 VDD1.n1 VDD1.t4 2.18352
R79 VDD1 VDD1.n5 0.205241
R80 B.n300 B.t19 999.804
R81 B.n297 B.t12 999.804
R82 B.n74 B.t16 999.804
R83 B.n72 B.t8 999.804
R84 B.n529 B.n528 585
R85 B.n226 B.n71 585
R86 B.n225 B.n224 585
R87 B.n223 B.n222 585
R88 B.n221 B.n220 585
R89 B.n219 B.n218 585
R90 B.n217 B.n216 585
R91 B.n215 B.n214 585
R92 B.n213 B.n212 585
R93 B.n211 B.n210 585
R94 B.n209 B.n208 585
R95 B.n207 B.n206 585
R96 B.n205 B.n204 585
R97 B.n203 B.n202 585
R98 B.n201 B.n200 585
R99 B.n199 B.n198 585
R100 B.n197 B.n196 585
R101 B.n195 B.n194 585
R102 B.n193 B.n192 585
R103 B.n191 B.n190 585
R104 B.n189 B.n188 585
R105 B.n187 B.n186 585
R106 B.n185 B.n184 585
R107 B.n183 B.n182 585
R108 B.n181 B.n180 585
R109 B.n179 B.n178 585
R110 B.n177 B.n176 585
R111 B.n175 B.n174 585
R112 B.n173 B.n172 585
R113 B.n171 B.n170 585
R114 B.n169 B.n168 585
R115 B.n167 B.n166 585
R116 B.n165 B.n164 585
R117 B.n162 B.n161 585
R118 B.n160 B.n159 585
R119 B.n158 B.n157 585
R120 B.n156 B.n155 585
R121 B.n154 B.n153 585
R122 B.n152 B.n151 585
R123 B.n150 B.n149 585
R124 B.n148 B.n147 585
R125 B.n146 B.n145 585
R126 B.n144 B.n143 585
R127 B.n141 B.n140 585
R128 B.n139 B.n138 585
R129 B.n137 B.n136 585
R130 B.n135 B.n134 585
R131 B.n133 B.n132 585
R132 B.n131 B.n130 585
R133 B.n129 B.n128 585
R134 B.n127 B.n126 585
R135 B.n125 B.n124 585
R136 B.n123 B.n122 585
R137 B.n121 B.n120 585
R138 B.n119 B.n118 585
R139 B.n117 B.n116 585
R140 B.n115 B.n114 585
R141 B.n113 B.n112 585
R142 B.n111 B.n110 585
R143 B.n109 B.n108 585
R144 B.n107 B.n106 585
R145 B.n105 B.n104 585
R146 B.n103 B.n102 585
R147 B.n101 B.n100 585
R148 B.n99 B.n98 585
R149 B.n97 B.n96 585
R150 B.n95 B.n94 585
R151 B.n93 B.n92 585
R152 B.n91 B.n90 585
R153 B.n89 B.n88 585
R154 B.n87 B.n86 585
R155 B.n85 B.n84 585
R156 B.n83 B.n82 585
R157 B.n81 B.n80 585
R158 B.n79 B.n78 585
R159 B.n77 B.n76 585
R160 B.n527 B.n33 585
R161 B.n532 B.n33 585
R162 B.n526 B.n32 585
R163 B.n533 B.n32 585
R164 B.n525 B.n524 585
R165 B.n524 B.n28 585
R166 B.n523 B.n27 585
R167 B.n539 B.n27 585
R168 B.n522 B.n26 585
R169 B.n540 B.n26 585
R170 B.n521 B.n25 585
R171 B.n541 B.n25 585
R172 B.n520 B.n519 585
R173 B.n519 B.n21 585
R174 B.n518 B.n20 585
R175 B.n547 B.n20 585
R176 B.n517 B.n19 585
R177 B.n548 B.n19 585
R178 B.n516 B.n18 585
R179 B.n549 B.n18 585
R180 B.n515 B.n514 585
R181 B.n514 B.n513 585
R182 B.n512 B.n14 585
R183 B.n555 B.n14 585
R184 B.n511 B.n13 585
R185 B.n556 B.n13 585
R186 B.n510 B.n12 585
R187 B.n557 B.n12 585
R188 B.n509 B.n508 585
R189 B.n508 B.n11 585
R190 B.n507 B.n7 585
R191 B.n563 B.n7 585
R192 B.n506 B.n6 585
R193 B.n564 B.n6 585
R194 B.n505 B.n5 585
R195 B.n565 B.n5 585
R196 B.n504 B.n503 585
R197 B.n503 B.n4 585
R198 B.n502 B.n227 585
R199 B.n502 B.n501 585
R200 B.n491 B.n228 585
R201 B.n494 B.n228 585
R202 B.n493 B.n492 585
R203 B.n495 B.n493 585
R204 B.n490 B.n232 585
R205 B.n235 B.n232 585
R206 B.n489 B.n488 585
R207 B.n488 B.n487 585
R208 B.n234 B.n233 585
R209 B.n480 B.n234 585
R210 B.n479 B.n478 585
R211 B.n481 B.n479 585
R212 B.n477 B.n240 585
R213 B.n240 B.n239 585
R214 B.n476 B.n475 585
R215 B.n475 B.n474 585
R216 B.n242 B.n241 585
R217 B.n243 B.n242 585
R218 B.n467 B.n466 585
R219 B.n468 B.n467 585
R220 B.n465 B.n247 585
R221 B.n251 B.n247 585
R222 B.n464 B.n463 585
R223 B.n463 B.n462 585
R224 B.n249 B.n248 585
R225 B.n250 B.n249 585
R226 B.n455 B.n454 585
R227 B.n456 B.n455 585
R228 B.n453 B.n256 585
R229 B.n256 B.n255 585
R230 B.n448 B.n447 585
R231 B.n446 B.n296 585
R232 B.n445 B.n295 585
R233 B.n450 B.n295 585
R234 B.n444 B.n443 585
R235 B.n442 B.n441 585
R236 B.n440 B.n439 585
R237 B.n438 B.n437 585
R238 B.n436 B.n435 585
R239 B.n434 B.n433 585
R240 B.n432 B.n431 585
R241 B.n430 B.n429 585
R242 B.n428 B.n427 585
R243 B.n426 B.n425 585
R244 B.n424 B.n423 585
R245 B.n422 B.n421 585
R246 B.n420 B.n419 585
R247 B.n418 B.n417 585
R248 B.n416 B.n415 585
R249 B.n414 B.n413 585
R250 B.n412 B.n411 585
R251 B.n410 B.n409 585
R252 B.n408 B.n407 585
R253 B.n406 B.n405 585
R254 B.n404 B.n403 585
R255 B.n402 B.n401 585
R256 B.n400 B.n399 585
R257 B.n398 B.n397 585
R258 B.n396 B.n395 585
R259 B.n394 B.n393 585
R260 B.n392 B.n391 585
R261 B.n390 B.n389 585
R262 B.n388 B.n387 585
R263 B.n386 B.n385 585
R264 B.n384 B.n383 585
R265 B.n382 B.n381 585
R266 B.n380 B.n379 585
R267 B.n378 B.n377 585
R268 B.n376 B.n375 585
R269 B.n374 B.n373 585
R270 B.n372 B.n371 585
R271 B.n370 B.n369 585
R272 B.n368 B.n367 585
R273 B.n366 B.n365 585
R274 B.n364 B.n363 585
R275 B.n362 B.n361 585
R276 B.n360 B.n359 585
R277 B.n358 B.n357 585
R278 B.n356 B.n355 585
R279 B.n354 B.n353 585
R280 B.n352 B.n351 585
R281 B.n350 B.n349 585
R282 B.n348 B.n347 585
R283 B.n346 B.n345 585
R284 B.n344 B.n343 585
R285 B.n342 B.n341 585
R286 B.n340 B.n339 585
R287 B.n338 B.n337 585
R288 B.n336 B.n335 585
R289 B.n334 B.n333 585
R290 B.n332 B.n331 585
R291 B.n330 B.n329 585
R292 B.n328 B.n327 585
R293 B.n326 B.n325 585
R294 B.n324 B.n323 585
R295 B.n322 B.n321 585
R296 B.n320 B.n319 585
R297 B.n318 B.n317 585
R298 B.n316 B.n315 585
R299 B.n314 B.n313 585
R300 B.n312 B.n311 585
R301 B.n310 B.n309 585
R302 B.n308 B.n307 585
R303 B.n306 B.n305 585
R304 B.n304 B.n303 585
R305 B.n258 B.n257 585
R306 B.n452 B.n451 585
R307 B.n451 B.n450 585
R308 B.n254 B.n253 585
R309 B.n255 B.n254 585
R310 B.n458 B.n457 585
R311 B.n457 B.n456 585
R312 B.n459 B.n252 585
R313 B.n252 B.n250 585
R314 B.n461 B.n460 585
R315 B.n462 B.n461 585
R316 B.n246 B.n245 585
R317 B.n251 B.n246 585
R318 B.n470 B.n469 585
R319 B.n469 B.n468 585
R320 B.n471 B.n244 585
R321 B.n244 B.n243 585
R322 B.n473 B.n472 585
R323 B.n474 B.n473 585
R324 B.n238 B.n237 585
R325 B.n239 B.n238 585
R326 B.n483 B.n482 585
R327 B.n482 B.n481 585
R328 B.n484 B.n236 585
R329 B.n480 B.n236 585
R330 B.n486 B.n485 585
R331 B.n487 B.n486 585
R332 B.n231 B.n230 585
R333 B.n235 B.n231 585
R334 B.n497 B.n496 585
R335 B.n496 B.n495 585
R336 B.n498 B.n229 585
R337 B.n494 B.n229 585
R338 B.n500 B.n499 585
R339 B.n501 B.n500 585
R340 B.n2 B.n0 585
R341 B.n4 B.n2 585
R342 B.n3 B.n1 585
R343 B.n564 B.n3 585
R344 B.n562 B.n561 585
R345 B.n563 B.n562 585
R346 B.n560 B.n8 585
R347 B.n11 B.n8 585
R348 B.n559 B.n558 585
R349 B.n558 B.n557 585
R350 B.n10 B.n9 585
R351 B.n556 B.n10 585
R352 B.n554 B.n553 585
R353 B.n555 B.n554 585
R354 B.n552 B.n15 585
R355 B.n513 B.n15 585
R356 B.n551 B.n550 585
R357 B.n550 B.n549 585
R358 B.n17 B.n16 585
R359 B.n548 B.n17 585
R360 B.n546 B.n545 585
R361 B.n547 B.n546 585
R362 B.n544 B.n22 585
R363 B.n22 B.n21 585
R364 B.n543 B.n542 585
R365 B.n542 B.n541 585
R366 B.n24 B.n23 585
R367 B.n540 B.n24 585
R368 B.n538 B.n537 585
R369 B.n539 B.n538 585
R370 B.n536 B.n29 585
R371 B.n29 B.n28 585
R372 B.n535 B.n534 585
R373 B.n534 B.n533 585
R374 B.n31 B.n30 585
R375 B.n532 B.n31 585
R376 B.n567 B.n566 585
R377 B.n566 B.n565 585
R378 B.n448 B.n254 478.086
R379 B.n76 B.n31 478.086
R380 B.n451 B.n256 478.086
R381 B.n529 B.n33 478.086
R382 B.n531 B.n530 256.663
R383 B.n531 B.n70 256.663
R384 B.n531 B.n69 256.663
R385 B.n531 B.n68 256.663
R386 B.n531 B.n67 256.663
R387 B.n531 B.n66 256.663
R388 B.n531 B.n65 256.663
R389 B.n531 B.n64 256.663
R390 B.n531 B.n63 256.663
R391 B.n531 B.n62 256.663
R392 B.n531 B.n61 256.663
R393 B.n531 B.n60 256.663
R394 B.n531 B.n59 256.663
R395 B.n531 B.n58 256.663
R396 B.n531 B.n57 256.663
R397 B.n531 B.n56 256.663
R398 B.n531 B.n55 256.663
R399 B.n531 B.n54 256.663
R400 B.n531 B.n53 256.663
R401 B.n531 B.n52 256.663
R402 B.n531 B.n51 256.663
R403 B.n531 B.n50 256.663
R404 B.n531 B.n49 256.663
R405 B.n531 B.n48 256.663
R406 B.n531 B.n47 256.663
R407 B.n531 B.n46 256.663
R408 B.n531 B.n45 256.663
R409 B.n531 B.n44 256.663
R410 B.n531 B.n43 256.663
R411 B.n531 B.n42 256.663
R412 B.n531 B.n41 256.663
R413 B.n531 B.n40 256.663
R414 B.n531 B.n39 256.663
R415 B.n531 B.n38 256.663
R416 B.n531 B.n37 256.663
R417 B.n531 B.n36 256.663
R418 B.n531 B.n35 256.663
R419 B.n531 B.n34 256.663
R420 B.n450 B.n449 256.663
R421 B.n450 B.n259 256.663
R422 B.n450 B.n260 256.663
R423 B.n450 B.n261 256.663
R424 B.n450 B.n262 256.663
R425 B.n450 B.n263 256.663
R426 B.n450 B.n264 256.663
R427 B.n450 B.n265 256.663
R428 B.n450 B.n266 256.663
R429 B.n450 B.n267 256.663
R430 B.n450 B.n268 256.663
R431 B.n450 B.n269 256.663
R432 B.n450 B.n270 256.663
R433 B.n450 B.n271 256.663
R434 B.n450 B.n272 256.663
R435 B.n450 B.n273 256.663
R436 B.n450 B.n274 256.663
R437 B.n450 B.n275 256.663
R438 B.n450 B.n276 256.663
R439 B.n450 B.n277 256.663
R440 B.n450 B.n278 256.663
R441 B.n450 B.n279 256.663
R442 B.n450 B.n280 256.663
R443 B.n450 B.n281 256.663
R444 B.n450 B.n282 256.663
R445 B.n450 B.n283 256.663
R446 B.n450 B.n284 256.663
R447 B.n450 B.n285 256.663
R448 B.n450 B.n286 256.663
R449 B.n450 B.n287 256.663
R450 B.n450 B.n288 256.663
R451 B.n450 B.n289 256.663
R452 B.n450 B.n290 256.663
R453 B.n450 B.n291 256.663
R454 B.n450 B.n292 256.663
R455 B.n450 B.n293 256.663
R456 B.n450 B.n294 256.663
R457 B.n457 B.n254 163.367
R458 B.n457 B.n252 163.367
R459 B.n461 B.n252 163.367
R460 B.n461 B.n246 163.367
R461 B.n469 B.n246 163.367
R462 B.n469 B.n244 163.367
R463 B.n473 B.n244 163.367
R464 B.n473 B.n238 163.367
R465 B.n482 B.n238 163.367
R466 B.n482 B.n236 163.367
R467 B.n486 B.n236 163.367
R468 B.n486 B.n231 163.367
R469 B.n496 B.n231 163.367
R470 B.n496 B.n229 163.367
R471 B.n500 B.n229 163.367
R472 B.n500 B.n2 163.367
R473 B.n566 B.n2 163.367
R474 B.n566 B.n3 163.367
R475 B.n562 B.n3 163.367
R476 B.n562 B.n8 163.367
R477 B.n558 B.n8 163.367
R478 B.n558 B.n10 163.367
R479 B.n554 B.n10 163.367
R480 B.n554 B.n15 163.367
R481 B.n550 B.n15 163.367
R482 B.n550 B.n17 163.367
R483 B.n546 B.n17 163.367
R484 B.n546 B.n22 163.367
R485 B.n542 B.n22 163.367
R486 B.n542 B.n24 163.367
R487 B.n538 B.n24 163.367
R488 B.n538 B.n29 163.367
R489 B.n534 B.n29 163.367
R490 B.n534 B.n31 163.367
R491 B.n296 B.n295 163.367
R492 B.n443 B.n295 163.367
R493 B.n441 B.n440 163.367
R494 B.n437 B.n436 163.367
R495 B.n433 B.n432 163.367
R496 B.n429 B.n428 163.367
R497 B.n425 B.n424 163.367
R498 B.n421 B.n420 163.367
R499 B.n417 B.n416 163.367
R500 B.n413 B.n412 163.367
R501 B.n409 B.n408 163.367
R502 B.n405 B.n404 163.367
R503 B.n401 B.n400 163.367
R504 B.n397 B.n396 163.367
R505 B.n393 B.n392 163.367
R506 B.n389 B.n388 163.367
R507 B.n385 B.n384 163.367
R508 B.n381 B.n380 163.367
R509 B.n377 B.n376 163.367
R510 B.n373 B.n372 163.367
R511 B.n369 B.n368 163.367
R512 B.n365 B.n364 163.367
R513 B.n361 B.n360 163.367
R514 B.n357 B.n356 163.367
R515 B.n353 B.n352 163.367
R516 B.n349 B.n348 163.367
R517 B.n345 B.n344 163.367
R518 B.n341 B.n340 163.367
R519 B.n337 B.n336 163.367
R520 B.n333 B.n332 163.367
R521 B.n329 B.n328 163.367
R522 B.n325 B.n324 163.367
R523 B.n321 B.n320 163.367
R524 B.n317 B.n316 163.367
R525 B.n313 B.n312 163.367
R526 B.n309 B.n308 163.367
R527 B.n305 B.n304 163.367
R528 B.n451 B.n258 163.367
R529 B.n455 B.n256 163.367
R530 B.n455 B.n249 163.367
R531 B.n463 B.n249 163.367
R532 B.n463 B.n247 163.367
R533 B.n467 B.n247 163.367
R534 B.n467 B.n242 163.367
R535 B.n475 B.n242 163.367
R536 B.n475 B.n240 163.367
R537 B.n479 B.n240 163.367
R538 B.n479 B.n234 163.367
R539 B.n488 B.n234 163.367
R540 B.n488 B.n232 163.367
R541 B.n493 B.n232 163.367
R542 B.n493 B.n228 163.367
R543 B.n502 B.n228 163.367
R544 B.n503 B.n502 163.367
R545 B.n503 B.n5 163.367
R546 B.n6 B.n5 163.367
R547 B.n7 B.n6 163.367
R548 B.n508 B.n7 163.367
R549 B.n508 B.n12 163.367
R550 B.n13 B.n12 163.367
R551 B.n14 B.n13 163.367
R552 B.n514 B.n14 163.367
R553 B.n514 B.n18 163.367
R554 B.n19 B.n18 163.367
R555 B.n20 B.n19 163.367
R556 B.n519 B.n20 163.367
R557 B.n519 B.n25 163.367
R558 B.n26 B.n25 163.367
R559 B.n27 B.n26 163.367
R560 B.n524 B.n27 163.367
R561 B.n524 B.n32 163.367
R562 B.n33 B.n32 163.367
R563 B.n80 B.n79 163.367
R564 B.n84 B.n83 163.367
R565 B.n88 B.n87 163.367
R566 B.n92 B.n91 163.367
R567 B.n96 B.n95 163.367
R568 B.n100 B.n99 163.367
R569 B.n104 B.n103 163.367
R570 B.n108 B.n107 163.367
R571 B.n112 B.n111 163.367
R572 B.n116 B.n115 163.367
R573 B.n120 B.n119 163.367
R574 B.n124 B.n123 163.367
R575 B.n128 B.n127 163.367
R576 B.n132 B.n131 163.367
R577 B.n136 B.n135 163.367
R578 B.n140 B.n139 163.367
R579 B.n145 B.n144 163.367
R580 B.n149 B.n148 163.367
R581 B.n153 B.n152 163.367
R582 B.n157 B.n156 163.367
R583 B.n161 B.n160 163.367
R584 B.n166 B.n165 163.367
R585 B.n170 B.n169 163.367
R586 B.n174 B.n173 163.367
R587 B.n178 B.n177 163.367
R588 B.n182 B.n181 163.367
R589 B.n186 B.n185 163.367
R590 B.n190 B.n189 163.367
R591 B.n194 B.n193 163.367
R592 B.n198 B.n197 163.367
R593 B.n202 B.n201 163.367
R594 B.n206 B.n205 163.367
R595 B.n210 B.n209 163.367
R596 B.n214 B.n213 163.367
R597 B.n218 B.n217 163.367
R598 B.n222 B.n221 163.367
R599 B.n224 B.n71 163.367
R600 B.n450 B.n255 98.92
R601 B.n532 B.n531 98.92
R602 B.n300 B.t21 84.6095
R603 B.n72 B.t10 84.6095
R604 B.n297 B.t15 84.5988
R605 B.n74 B.t17 84.5988
R606 B.n301 B.t20 72.7792
R607 B.n73 B.t11 72.7792
R608 B.n298 B.t14 72.7684
R609 B.n75 B.t18 72.7684
R610 B.n449 B.n448 71.676
R611 B.n443 B.n259 71.676
R612 B.n440 B.n260 71.676
R613 B.n436 B.n261 71.676
R614 B.n432 B.n262 71.676
R615 B.n428 B.n263 71.676
R616 B.n424 B.n264 71.676
R617 B.n420 B.n265 71.676
R618 B.n416 B.n266 71.676
R619 B.n412 B.n267 71.676
R620 B.n408 B.n268 71.676
R621 B.n404 B.n269 71.676
R622 B.n400 B.n270 71.676
R623 B.n396 B.n271 71.676
R624 B.n392 B.n272 71.676
R625 B.n388 B.n273 71.676
R626 B.n384 B.n274 71.676
R627 B.n380 B.n275 71.676
R628 B.n376 B.n276 71.676
R629 B.n372 B.n277 71.676
R630 B.n368 B.n278 71.676
R631 B.n364 B.n279 71.676
R632 B.n360 B.n280 71.676
R633 B.n356 B.n281 71.676
R634 B.n352 B.n282 71.676
R635 B.n348 B.n283 71.676
R636 B.n344 B.n284 71.676
R637 B.n340 B.n285 71.676
R638 B.n336 B.n286 71.676
R639 B.n332 B.n287 71.676
R640 B.n328 B.n288 71.676
R641 B.n324 B.n289 71.676
R642 B.n320 B.n290 71.676
R643 B.n316 B.n291 71.676
R644 B.n312 B.n292 71.676
R645 B.n308 B.n293 71.676
R646 B.n304 B.n294 71.676
R647 B.n76 B.n34 71.676
R648 B.n80 B.n35 71.676
R649 B.n84 B.n36 71.676
R650 B.n88 B.n37 71.676
R651 B.n92 B.n38 71.676
R652 B.n96 B.n39 71.676
R653 B.n100 B.n40 71.676
R654 B.n104 B.n41 71.676
R655 B.n108 B.n42 71.676
R656 B.n112 B.n43 71.676
R657 B.n116 B.n44 71.676
R658 B.n120 B.n45 71.676
R659 B.n124 B.n46 71.676
R660 B.n128 B.n47 71.676
R661 B.n132 B.n48 71.676
R662 B.n136 B.n49 71.676
R663 B.n140 B.n50 71.676
R664 B.n145 B.n51 71.676
R665 B.n149 B.n52 71.676
R666 B.n153 B.n53 71.676
R667 B.n157 B.n54 71.676
R668 B.n161 B.n55 71.676
R669 B.n166 B.n56 71.676
R670 B.n170 B.n57 71.676
R671 B.n174 B.n58 71.676
R672 B.n178 B.n59 71.676
R673 B.n182 B.n60 71.676
R674 B.n186 B.n61 71.676
R675 B.n190 B.n62 71.676
R676 B.n194 B.n63 71.676
R677 B.n198 B.n64 71.676
R678 B.n202 B.n65 71.676
R679 B.n206 B.n66 71.676
R680 B.n210 B.n67 71.676
R681 B.n214 B.n68 71.676
R682 B.n218 B.n69 71.676
R683 B.n222 B.n70 71.676
R684 B.n530 B.n71 71.676
R685 B.n530 B.n529 71.676
R686 B.n224 B.n70 71.676
R687 B.n221 B.n69 71.676
R688 B.n217 B.n68 71.676
R689 B.n213 B.n67 71.676
R690 B.n209 B.n66 71.676
R691 B.n205 B.n65 71.676
R692 B.n201 B.n64 71.676
R693 B.n197 B.n63 71.676
R694 B.n193 B.n62 71.676
R695 B.n189 B.n61 71.676
R696 B.n185 B.n60 71.676
R697 B.n181 B.n59 71.676
R698 B.n177 B.n58 71.676
R699 B.n173 B.n57 71.676
R700 B.n169 B.n56 71.676
R701 B.n165 B.n55 71.676
R702 B.n160 B.n54 71.676
R703 B.n156 B.n53 71.676
R704 B.n152 B.n52 71.676
R705 B.n148 B.n51 71.676
R706 B.n144 B.n50 71.676
R707 B.n139 B.n49 71.676
R708 B.n135 B.n48 71.676
R709 B.n131 B.n47 71.676
R710 B.n127 B.n46 71.676
R711 B.n123 B.n45 71.676
R712 B.n119 B.n44 71.676
R713 B.n115 B.n43 71.676
R714 B.n111 B.n42 71.676
R715 B.n107 B.n41 71.676
R716 B.n103 B.n40 71.676
R717 B.n99 B.n39 71.676
R718 B.n95 B.n38 71.676
R719 B.n91 B.n37 71.676
R720 B.n87 B.n36 71.676
R721 B.n83 B.n35 71.676
R722 B.n79 B.n34 71.676
R723 B.n449 B.n296 71.676
R724 B.n441 B.n259 71.676
R725 B.n437 B.n260 71.676
R726 B.n433 B.n261 71.676
R727 B.n429 B.n262 71.676
R728 B.n425 B.n263 71.676
R729 B.n421 B.n264 71.676
R730 B.n417 B.n265 71.676
R731 B.n413 B.n266 71.676
R732 B.n409 B.n267 71.676
R733 B.n405 B.n268 71.676
R734 B.n401 B.n269 71.676
R735 B.n397 B.n270 71.676
R736 B.n393 B.n271 71.676
R737 B.n389 B.n272 71.676
R738 B.n385 B.n273 71.676
R739 B.n381 B.n274 71.676
R740 B.n377 B.n275 71.676
R741 B.n373 B.n276 71.676
R742 B.n369 B.n277 71.676
R743 B.n365 B.n278 71.676
R744 B.n361 B.n279 71.676
R745 B.n357 B.n280 71.676
R746 B.n353 B.n281 71.676
R747 B.n349 B.n282 71.676
R748 B.n345 B.n283 71.676
R749 B.n341 B.n284 71.676
R750 B.n337 B.n285 71.676
R751 B.n333 B.n286 71.676
R752 B.n329 B.n287 71.676
R753 B.n325 B.n288 71.676
R754 B.n321 B.n289 71.676
R755 B.n317 B.n290 71.676
R756 B.n313 B.n291 71.676
R757 B.n309 B.n292 71.676
R758 B.n305 B.n293 71.676
R759 B.n294 B.n258 71.676
R760 B.n302 B.n301 59.5399
R761 B.n299 B.n298 59.5399
R762 B.n142 B.n75 59.5399
R763 B.n163 B.n73 59.5399
R764 B.n456 B.n255 52.1441
R765 B.n456 B.n250 52.1441
R766 B.n462 B.n250 52.1441
R767 B.n462 B.n251 52.1441
R768 B.n468 B.n243 52.1441
R769 B.n474 B.n243 52.1441
R770 B.n474 B.n239 52.1441
R771 B.n481 B.n239 52.1441
R772 B.n487 B.n235 52.1441
R773 B.n495 B.n494 52.1441
R774 B.n501 B.n4 52.1441
R775 B.n565 B.n4 52.1441
R776 B.n565 B.n564 52.1441
R777 B.n564 B.n563 52.1441
R778 B.n557 B.n11 52.1441
R779 B.n556 B.n555 52.1441
R780 B.n549 B.n548 52.1441
R781 B.n548 B.n547 52.1441
R782 B.n547 B.n21 52.1441
R783 B.n541 B.n21 52.1441
R784 B.n540 B.n539 52.1441
R785 B.n539 B.n28 52.1441
R786 B.n533 B.n28 52.1441
R787 B.n533 B.n532 52.1441
R788 B.n480 B.t7 47.5432
R789 B.n513 B.t5 47.5432
R790 B.n468 B.t13 46.0096
R791 B.t4 B.n480 46.0096
R792 B.n513 B.t3 46.0096
R793 B.n541 B.t9 46.0096
R794 B.n235 B.t0 36.8078
R795 B.t2 B.n556 36.8078
R796 B.n77 B.n30 31.0639
R797 B.n528 B.n527 31.0639
R798 B.n453 B.n452 31.0639
R799 B.n447 B.n253 31.0639
R800 B.n494 B.t6 26.0723
R801 B.n501 B.t6 26.0723
R802 B.n563 B.t1 26.0723
R803 B.n11 B.t1 26.0723
R804 B B.n567 18.0485
R805 B.n495 B.t0 15.3369
R806 B.n557 B.t2 15.3369
R807 B.n301 B.n300 11.8308
R808 B.n298 B.n297 11.8308
R809 B.n75 B.n74 11.8308
R810 B.n73 B.n72 11.8308
R811 B.n78 B.n77 10.6151
R812 B.n81 B.n78 10.6151
R813 B.n82 B.n81 10.6151
R814 B.n85 B.n82 10.6151
R815 B.n86 B.n85 10.6151
R816 B.n89 B.n86 10.6151
R817 B.n90 B.n89 10.6151
R818 B.n93 B.n90 10.6151
R819 B.n94 B.n93 10.6151
R820 B.n97 B.n94 10.6151
R821 B.n98 B.n97 10.6151
R822 B.n101 B.n98 10.6151
R823 B.n102 B.n101 10.6151
R824 B.n105 B.n102 10.6151
R825 B.n106 B.n105 10.6151
R826 B.n109 B.n106 10.6151
R827 B.n110 B.n109 10.6151
R828 B.n113 B.n110 10.6151
R829 B.n114 B.n113 10.6151
R830 B.n117 B.n114 10.6151
R831 B.n118 B.n117 10.6151
R832 B.n121 B.n118 10.6151
R833 B.n122 B.n121 10.6151
R834 B.n125 B.n122 10.6151
R835 B.n126 B.n125 10.6151
R836 B.n129 B.n126 10.6151
R837 B.n130 B.n129 10.6151
R838 B.n133 B.n130 10.6151
R839 B.n134 B.n133 10.6151
R840 B.n137 B.n134 10.6151
R841 B.n138 B.n137 10.6151
R842 B.n141 B.n138 10.6151
R843 B.n146 B.n143 10.6151
R844 B.n147 B.n146 10.6151
R845 B.n150 B.n147 10.6151
R846 B.n151 B.n150 10.6151
R847 B.n154 B.n151 10.6151
R848 B.n155 B.n154 10.6151
R849 B.n158 B.n155 10.6151
R850 B.n159 B.n158 10.6151
R851 B.n162 B.n159 10.6151
R852 B.n167 B.n164 10.6151
R853 B.n168 B.n167 10.6151
R854 B.n171 B.n168 10.6151
R855 B.n172 B.n171 10.6151
R856 B.n175 B.n172 10.6151
R857 B.n176 B.n175 10.6151
R858 B.n179 B.n176 10.6151
R859 B.n180 B.n179 10.6151
R860 B.n183 B.n180 10.6151
R861 B.n184 B.n183 10.6151
R862 B.n187 B.n184 10.6151
R863 B.n188 B.n187 10.6151
R864 B.n191 B.n188 10.6151
R865 B.n192 B.n191 10.6151
R866 B.n195 B.n192 10.6151
R867 B.n196 B.n195 10.6151
R868 B.n199 B.n196 10.6151
R869 B.n200 B.n199 10.6151
R870 B.n203 B.n200 10.6151
R871 B.n204 B.n203 10.6151
R872 B.n207 B.n204 10.6151
R873 B.n208 B.n207 10.6151
R874 B.n211 B.n208 10.6151
R875 B.n212 B.n211 10.6151
R876 B.n215 B.n212 10.6151
R877 B.n216 B.n215 10.6151
R878 B.n219 B.n216 10.6151
R879 B.n220 B.n219 10.6151
R880 B.n223 B.n220 10.6151
R881 B.n225 B.n223 10.6151
R882 B.n226 B.n225 10.6151
R883 B.n528 B.n226 10.6151
R884 B.n454 B.n453 10.6151
R885 B.n454 B.n248 10.6151
R886 B.n464 B.n248 10.6151
R887 B.n465 B.n464 10.6151
R888 B.n466 B.n465 10.6151
R889 B.n466 B.n241 10.6151
R890 B.n476 B.n241 10.6151
R891 B.n477 B.n476 10.6151
R892 B.n478 B.n477 10.6151
R893 B.n478 B.n233 10.6151
R894 B.n489 B.n233 10.6151
R895 B.n490 B.n489 10.6151
R896 B.n492 B.n490 10.6151
R897 B.n492 B.n491 10.6151
R898 B.n491 B.n227 10.6151
R899 B.n504 B.n227 10.6151
R900 B.n505 B.n504 10.6151
R901 B.n506 B.n505 10.6151
R902 B.n507 B.n506 10.6151
R903 B.n509 B.n507 10.6151
R904 B.n510 B.n509 10.6151
R905 B.n511 B.n510 10.6151
R906 B.n512 B.n511 10.6151
R907 B.n515 B.n512 10.6151
R908 B.n516 B.n515 10.6151
R909 B.n517 B.n516 10.6151
R910 B.n518 B.n517 10.6151
R911 B.n520 B.n518 10.6151
R912 B.n521 B.n520 10.6151
R913 B.n522 B.n521 10.6151
R914 B.n523 B.n522 10.6151
R915 B.n525 B.n523 10.6151
R916 B.n526 B.n525 10.6151
R917 B.n527 B.n526 10.6151
R918 B.n447 B.n446 10.6151
R919 B.n446 B.n445 10.6151
R920 B.n445 B.n444 10.6151
R921 B.n444 B.n442 10.6151
R922 B.n442 B.n439 10.6151
R923 B.n439 B.n438 10.6151
R924 B.n438 B.n435 10.6151
R925 B.n435 B.n434 10.6151
R926 B.n434 B.n431 10.6151
R927 B.n431 B.n430 10.6151
R928 B.n430 B.n427 10.6151
R929 B.n427 B.n426 10.6151
R930 B.n426 B.n423 10.6151
R931 B.n423 B.n422 10.6151
R932 B.n422 B.n419 10.6151
R933 B.n419 B.n418 10.6151
R934 B.n418 B.n415 10.6151
R935 B.n415 B.n414 10.6151
R936 B.n414 B.n411 10.6151
R937 B.n411 B.n410 10.6151
R938 B.n410 B.n407 10.6151
R939 B.n407 B.n406 10.6151
R940 B.n406 B.n403 10.6151
R941 B.n403 B.n402 10.6151
R942 B.n402 B.n399 10.6151
R943 B.n399 B.n398 10.6151
R944 B.n398 B.n395 10.6151
R945 B.n395 B.n394 10.6151
R946 B.n394 B.n391 10.6151
R947 B.n391 B.n390 10.6151
R948 B.n390 B.n387 10.6151
R949 B.n387 B.n386 10.6151
R950 B.n383 B.n382 10.6151
R951 B.n382 B.n379 10.6151
R952 B.n379 B.n378 10.6151
R953 B.n378 B.n375 10.6151
R954 B.n375 B.n374 10.6151
R955 B.n374 B.n371 10.6151
R956 B.n371 B.n370 10.6151
R957 B.n370 B.n367 10.6151
R958 B.n367 B.n366 10.6151
R959 B.n363 B.n362 10.6151
R960 B.n362 B.n359 10.6151
R961 B.n359 B.n358 10.6151
R962 B.n358 B.n355 10.6151
R963 B.n355 B.n354 10.6151
R964 B.n354 B.n351 10.6151
R965 B.n351 B.n350 10.6151
R966 B.n350 B.n347 10.6151
R967 B.n347 B.n346 10.6151
R968 B.n346 B.n343 10.6151
R969 B.n343 B.n342 10.6151
R970 B.n342 B.n339 10.6151
R971 B.n339 B.n338 10.6151
R972 B.n338 B.n335 10.6151
R973 B.n335 B.n334 10.6151
R974 B.n334 B.n331 10.6151
R975 B.n331 B.n330 10.6151
R976 B.n330 B.n327 10.6151
R977 B.n327 B.n326 10.6151
R978 B.n326 B.n323 10.6151
R979 B.n323 B.n322 10.6151
R980 B.n322 B.n319 10.6151
R981 B.n319 B.n318 10.6151
R982 B.n318 B.n315 10.6151
R983 B.n315 B.n314 10.6151
R984 B.n314 B.n311 10.6151
R985 B.n311 B.n310 10.6151
R986 B.n310 B.n307 10.6151
R987 B.n307 B.n306 10.6151
R988 B.n306 B.n303 10.6151
R989 B.n303 B.n257 10.6151
R990 B.n452 B.n257 10.6151
R991 B.n458 B.n253 10.6151
R992 B.n459 B.n458 10.6151
R993 B.n460 B.n459 10.6151
R994 B.n460 B.n245 10.6151
R995 B.n470 B.n245 10.6151
R996 B.n471 B.n470 10.6151
R997 B.n472 B.n471 10.6151
R998 B.n472 B.n237 10.6151
R999 B.n483 B.n237 10.6151
R1000 B.n484 B.n483 10.6151
R1001 B.n485 B.n484 10.6151
R1002 B.n485 B.n230 10.6151
R1003 B.n497 B.n230 10.6151
R1004 B.n498 B.n497 10.6151
R1005 B.n499 B.n498 10.6151
R1006 B.n499 B.n0 10.6151
R1007 B.n561 B.n1 10.6151
R1008 B.n561 B.n560 10.6151
R1009 B.n560 B.n559 10.6151
R1010 B.n559 B.n9 10.6151
R1011 B.n553 B.n9 10.6151
R1012 B.n553 B.n552 10.6151
R1013 B.n552 B.n551 10.6151
R1014 B.n551 B.n16 10.6151
R1015 B.n545 B.n16 10.6151
R1016 B.n545 B.n544 10.6151
R1017 B.n544 B.n543 10.6151
R1018 B.n543 B.n23 10.6151
R1019 B.n537 B.n23 10.6151
R1020 B.n537 B.n536 10.6151
R1021 B.n536 B.n535 10.6151
R1022 B.n535 B.n30 10.6151
R1023 B.n142 B.n141 9.36635
R1024 B.n164 B.n163 9.36635
R1025 B.n386 B.n299 9.36635
R1026 B.n363 B.n302 9.36635
R1027 B.n251 B.t13 6.13504
R1028 B.n481 B.t4 6.13504
R1029 B.n549 B.t3 6.13504
R1030 B.t9 B.n540 6.13504
R1031 B.n487 B.t7 4.60141
R1032 B.n555 B.t5 4.60141
R1033 B.n567 B.n0 2.81026
R1034 B.n567 B.n1 2.81026
R1035 B.n143 B.n142 1.24928
R1036 B.n163 B.n162 1.24928
R1037 B.n383 B.n299 1.24928
R1038 B.n366 B.n302 1.24928
R1039 VN.n7 VN.t5 917.521
R1040 VN.n2 VN.t0 917.521
R1041 VN.n16 VN.t3 917.521
R1042 VN.n11 VN.t4 917.521
R1043 VN.n6 VN.t7 893.422
R1044 VN.n1 VN.t2 893.422
R1045 VN.n15 VN.t6 893.422
R1046 VN.n10 VN.t1 893.422
R1047 VN.n12 VN.n11 161.489
R1048 VN.n3 VN.n2 161.489
R1049 VN.n8 VN.n7 161.3
R1050 VN.n17 VN.n16 161.3
R1051 VN.n14 VN.n9 161.3
R1052 VN.n13 VN.n12 161.3
R1053 VN.n5 VN.n0 161.3
R1054 VN.n4 VN.n3 161.3
R1055 VN.n5 VN.n4 73.0308
R1056 VN.n14 VN.n13 73.0308
R1057 VN.n2 VN.n1 64.9975
R1058 VN.n7 VN.n6 64.9975
R1059 VN.n16 VN.n15 64.9975
R1060 VN.n11 VN.n10 64.9975
R1061 VN VN.n17 38.1766
R1062 VN.n4 VN.n1 8.03383
R1063 VN.n6 VN.n5 8.03383
R1064 VN.n15 VN.n14 8.03383
R1065 VN.n13 VN.n10 8.03383
R1066 VN.n17 VN.n9 0.189894
R1067 VN.n12 VN.n9 0.189894
R1068 VN.n3 VN.n0 0.189894
R1069 VN.n8 VN.n0 0.189894
R1070 VN VN.n8 0.0516364
R1071 VDD2.n2 VDD2.n1 67.1025
R1072 VDD2.n2 VDD2.n0 67.1025
R1073 VDD2 VDD2.n5 67.0997
R1074 VDD2.n4 VDD2.n3 66.8952
R1075 VDD2.n4 VDD2.n2 33.9006
R1076 VDD2.n5 VDD2.t6 2.18352
R1077 VDD2.n5 VDD2.t3 2.18352
R1078 VDD2.n3 VDD2.t4 2.18352
R1079 VDD2.n3 VDD2.t1 2.18352
R1080 VDD2.n1 VDD2.t0 2.18352
R1081 VDD2.n1 VDD2.t2 2.18352
R1082 VDD2.n0 VDD2.t7 2.18352
R1083 VDD2.n0 VDD2.t5 2.18352
R1084 VDD2 VDD2.n4 0.321621
C0 VN VDD2 2.5011f
C1 VN VTAIL 2.18589f
C2 VDD2 VTAIL 13.2621f
C3 VN VDD1 0.147458f
C4 VDD1 VDD2 0.622516f
C5 VDD1 VTAIL 13.2233f
C6 VN VP 4.28643f
C7 VDD2 VP 0.272722f
C8 VTAIL VP 2.2f
C9 VDD1 VP 2.62615f
C10 VDD2 B 2.893951f
C11 VDD1 B 3.06781f
C12 VTAIL B 6.866367f
C13 VN B 6.83779f
C14 VP B 4.789098f
C15 VDD2.t7 B 0.242654f
C16 VDD2.t5 B 0.242654f
C17 VDD2.n0 B 2.12598f
C18 VDD2.t0 B 0.242654f
C19 VDD2.t2 B 0.242654f
C20 VDD2.n1 B 2.12598f
C21 VDD2.n2 B 2.35303f
C22 VDD2.t4 B 0.242654f
C23 VDD2.t1 B 0.242654f
C24 VDD2.n3 B 2.12485f
C25 VDD2.n4 B 2.58318f
C26 VDD2.t6 B 0.242654f
C27 VDD2.t3 B 0.242654f
C28 VDD2.n5 B 2.12595f
C29 VN.n0 B 0.055568f
C30 VN.t7 B 0.399994f
C31 VN.t2 B 0.399994f
C32 VN.n1 B 0.168f
C33 VN.t0 B 0.404357f
C34 VN.n2 B 0.184024f
C35 VN.n3 B 0.114836f
C36 VN.n4 B 0.020318f
C37 VN.n5 B 0.020318f
C38 VN.n6 B 0.168f
C39 VN.t5 B 0.404357f
C40 VN.n7 B 0.183955f
C41 VN.n8 B 0.043063f
C42 VN.n9 B 0.055568f
C43 VN.t3 B 0.404357f
C44 VN.t6 B 0.399994f
C45 VN.t1 B 0.399994f
C46 VN.n10 B 0.168f
C47 VN.t4 B 0.404357f
C48 VN.n11 B 0.184024f
C49 VN.n12 B 0.114836f
C50 VN.n13 B 0.020318f
C51 VN.n14 B 0.020318f
C52 VN.n15 B 0.168f
C53 VN.n16 B 0.183955f
C54 VN.n17 B 1.94753f
C55 VDD1.t5 B 0.240749f
C56 VDD1.t7 B 0.240749f
C57 VDD1.n0 B 2.10995f
C58 VDD1.t1 B 0.240749f
C59 VDD1.t4 B 0.240749f
C60 VDD1.n1 B 2.10929f
C61 VDD1.t2 B 0.240749f
C62 VDD1.t0 B 0.240749f
C63 VDD1.n2 B 2.10929f
C64 VDD1.n3 B 2.40691f
C65 VDD1.t3 B 0.240749f
C66 VDD1.t6 B 0.240749f
C67 VDD1.n4 B 2.10816f
C68 VDD1.n5 B 2.60202f
C69 VTAIL.t2 B 0.178407f
C70 VTAIL.t5 B 0.178407f
C71 VTAIL.n0 B 1.49785f
C72 VTAIL.n1 B 0.276074f
C73 VTAIL.t1 B 1.90917f
C74 VTAIL.n2 B 0.384332f
C75 VTAIL.t11 B 1.90917f
C76 VTAIL.n3 B 0.384332f
C77 VTAIL.t9 B 0.178407f
C78 VTAIL.t12 B 0.178407f
C79 VTAIL.n4 B 1.49785f
C80 VTAIL.n5 B 0.313585f
C81 VTAIL.t8 B 1.90917f
C82 VTAIL.n6 B 1.35408f
C83 VTAIL.t4 B 1.90918f
C84 VTAIL.n7 B 1.35407f
C85 VTAIL.t7 B 0.178407f
C86 VTAIL.t0 B 0.178407f
C87 VTAIL.n8 B 1.49785f
C88 VTAIL.n9 B 0.31358f
C89 VTAIL.t6 B 1.90918f
C90 VTAIL.n10 B 0.384327f
C91 VTAIL.t10 B 1.90918f
C92 VTAIL.n11 B 0.384327f
C93 VTAIL.t15 B 0.178407f
C94 VTAIL.t13 B 0.178407f
C95 VTAIL.n12 B 1.49785f
C96 VTAIL.n13 B 0.31358f
C97 VTAIL.t14 B 1.90917f
C98 VTAIL.n14 B 1.35408f
C99 VTAIL.t3 B 1.90917f
C100 VTAIL.n15 B 1.34941f
C101 VP.n0 B 0.056678f
C102 VP.t5 B 0.407979f
C103 VP.t3 B 0.407979f
C104 VP.n1 B 0.171354f
C105 VP.n2 B 0.056678f
C106 VP.t4 B 0.407979f
C107 VP.t0 B 0.407979f
C108 VP.n3 B 0.171354f
C109 VP.t2 B 0.412429f
C110 VP.n4 B 0.187698f
C111 VP.n5 B 0.117128f
C112 VP.n6 B 0.020724f
C113 VP.n7 B 0.020724f
C114 VP.n8 B 0.171354f
C115 VP.t1 B 0.412429f
C116 VP.n9 B 0.187627f
C117 VP.n10 B 1.94895f
C118 VP.t6 B 0.412429f
C119 VP.n11 B 0.187627f
C120 VP.n12 B 2.00285f
C121 VP.n13 B 0.056678f
C122 VP.n14 B 0.020724f
C123 VP.n15 B 0.020724f
C124 VP.n16 B 0.171354f
C125 VP.t7 B 0.412429f
C126 VP.n17 B 0.187627f
C127 VP.n18 B 0.043923f
.ends

