* NGSPICE file created from diff_pair_sample_0027.ext - technology: sky130A

.subckt diff_pair_sample_0027 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t14 VN.t0 VDD2.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=2.81325 ps=17.38 w=17.05 l=0.54
X1 VTAIL.t15 VP.t0 VDD1.t7 B.t21 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X2 VDD2.t5 VN.t1 VTAIL.t13 B.t1 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X3 VTAIL.t12 VN.t2 VDD2.t4 B.t21 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X4 VDD2.t7 VN.t3 VTAIL.t11 B.t6 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X5 B.t20 B.t18 B.t19 B.t12 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=0 ps=0 w=17.05 l=0.54
X6 VDD2.t6 VN.t4 VTAIL.t10 B.t3 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=6.6495 ps=34.88 w=17.05 l=0.54
X7 VDD1.t6 VP.t1 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=6.6495 ps=34.88 w=17.05 l=0.54
X8 VDD1.t5 VP.t2 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X9 VDD1.t4 VP.t3 VTAIL.t6 B.t6 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X10 B.t17 B.t15 B.t16 B.t8 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=0 ps=0 w=17.05 l=0.54
X11 VTAIL.t9 VN.t5 VDD2.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X12 B.t14 B.t11 B.t13 B.t12 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=0 ps=0 w=17.05 l=0.54
X13 VTAIL.t5 VP.t4 VDD1.t3 B.t5 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=2.81325 ps=17.38 w=17.05 l=0.54
X14 VDD2.t0 VN.t6 VTAIL.t8 B.t2 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=6.6495 ps=34.88 w=17.05 l=0.54
X15 VTAIL.t0 VP.t5 VDD1.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=2.81325 ps=17.38 w=17.05 l=0.54
X16 VTAIL.t4 VP.t6 VDD1.t1 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=2.81325 ps=17.38 w=17.05 l=0.54
X17 B.t10 B.t7 B.t9 B.t8 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=0 ps=0 w=17.05 l=0.54
X18 VDD1.t0 VP.t7 VTAIL.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=2.81325 pd=17.38 as=6.6495 ps=34.88 w=17.05 l=0.54
X19 VTAIL.t7 VN.t7 VDD2.t2 B.t4 sky130_fd_pr__nfet_01v8 ad=6.6495 pd=34.88 as=2.81325 ps=17.38 w=17.05 l=0.54
R0 VN.n2 VN.t0 859.521
R1 VN.n10 VN.t6 859.521
R2 VN.n1 VN.t3 834.129
R3 VN.n4 VN.t2 834.129
R4 VN.n6 VN.t4 834.129
R5 VN.n9 VN.t5 834.129
R6 VN.n12 VN.t1 834.129
R7 VN.n14 VN.t7 834.129
R8 VN.n7 VN.n6 161.3
R9 VN.n15 VN.n14 161.3
R10 VN.n13 VN.n8 161.3
R11 VN.n12 VN.n11 161.3
R12 VN.n5 VN.n0 161.3
R13 VN.n4 VN.n3 161.3
R14 VN.n4 VN.n1 48.2005
R15 VN.n12 VN.n9 48.2005
R16 VN VN.n15 45.4191
R17 VN.n11 VN.n10 45.0031
R18 VN.n3 VN.n2 45.0031
R19 VN.n6 VN.n5 41.6278
R20 VN.n14 VN.n13 41.6278
R21 VN.n2 VN.n1 15.6319
R22 VN.n10 VN.n9 15.6319
R23 VN.n5 VN.n4 6.57323
R24 VN.n13 VN.n12 6.57323
R25 VN.n15 VN.n8 0.189894
R26 VN.n11 VN.n8 0.189894
R27 VN.n3 VN.n0 0.189894
R28 VN.n7 VN.n0 0.189894
R29 VN VN.n7 0.0516364
R30 VDD2.n2 VDD2.n1 58.8881
R31 VDD2.n2 VDD2.n0 58.8881
R32 VDD2 VDD2.n5 58.8854
R33 VDD2.n4 VDD2.n3 58.5687
R34 VDD2.n4 VDD2.n2 41.7886
R35 VDD2.n5 VDD2.t1 1.16179
R36 VDD2.n5 VDD2.t0 1.16179
R37 VDD2.n3 VDD2.t2 1.16179
R38 VDD2.n3 VDD2.t5 1.16179
R39 VDD2.n1 VDD2.t4 1.16179
R40 VDD2.n1 VDD2.t6 1.16179
R41 VDD2.n0 VDD2.t3 1.16179
R42 VDD2.n0 VDD2.t7 1.16179
R43 VDD2 VDD2.n4 0.43369
R44 VTAIL.n11 VTAIL.t5 43.0512
R45 VTAIL.n10 VTAIL.t8 43.0512
R46 VTAIL.n7 VTAIL.t7 43.0512
R47 VTAIL.n15 VTAIL.t10 43.0511
R48 VTAIL.n2 VTAIL.t14 43.0511
R49 VTAIL.n3 VTAIL.t2 43.0511
R50 VTAIL.n6 VTAIL.t4 43.0511
R51 VTAIL.n14 VTAIL.t3 43.0511
R52 VTAIL.n13 VTAIL.n12 41.8899
R53 VTAIL.n9 VTAIL.n8 41.8899
R54 VTAIL.n1 VTAIL.n0 41.8897
R55 VTAIL.n5 VTAIL.n4 41.8897
R56 VTAIL.n15 VTAIL.n14 27.8152
R57 VTAIL.n7 VTAIL.n6 27.8152
R58 VTAIL.n0 VTAIL.t11 1.16179
R59 VTAIL.n0 VTAIL.t12 1.16179
R60 VTAIL.n4 VTAIL.t1 1.16179
R61 VTAIL.n4 VTAIL.t0 1.16179
R62 VTAIL.n12 VTAIL.t6 1.16179
R63 VTAIL.n12 VTAIL.t15 1.16179
R64 VTAIL.n8 VTAIL.t13 1.16179
R65 VTAIL.n8 VTAIL.t9 1.16179
R66 VTAIL.n9 VTAIL.n7 0.7505
R67 VTAIL.n10 VTAIL.n9 0.7505
R68 VTAIL.n13 VTAIL.n11 0.7505
R69 VTAIL.n14 VTAIL.n13 0.7505
R70 VTAIL.n6 VTAIL.n5 0.7505
R71 VTAIL.n5 VTAIL.n3 0.7505
R72 VTAIL.n2 VTAIL.n1 0.7505
R73 VTAIL VTAIL.n15 0.69231
R74 VTAIL.n11 VTAIL.n10 0.470328
R75 VTAIL.n3 VTAIL.n2 0.470328
R76 VTAIL VTAIL.n1 0.0586897
R77 B.n453 B.t7 966.451
R78 B.n451 B.t15 966.451
R79 B.n106 B.t18 966.451
R80 B.n103 B.t11 966.451
R81 B.n790 B.n789 585
R82 B.n349 B.n102 585
R83 B.n348 B.n347 585
R84 B.n346 B.n345 585
R85 B.n344 B.n343 585
R86 B.n342 B.n341 585
R87 B.n340 B.n339 585
R88 B.n338 B.n337 585
R89 B.n336 B.n335 585
R90 B.n334 B.n333 585
R91 B.n332 B.n331 585
R92 B.n330 B.n329 585
R93 B.n328 B.n327 585
R94 B.n326 B.n325 585
R95 B.n324 B.n323 585
R96 B.n322 B.n321 585
R97 B.n320 B.n319 585
R98 B.n318 B.n317 585
R99 B.n316 B.n315 585
R100 B.n314 B.n313 585
R101 B.n312 B.n311 585
R102 B.n310 B.n309 585
R103 B.n308 B.n307 585
R104 B.n306 B.n305 585
R105 B.n304 B.n303 585
R106 B.n302 B.n301 585
R107 B.n300 B.n299 585
R108 B.n298 B.n297 585
R109 B.n296 B.n295 585
R110 B.n294 B.n293 585
R111 B.n292 B.n291 585
R112 B.n290 B.n289 585
R113 B.n288 B.n287 585
R114 B.n286 B.n285 585
R115 B.n284 B.n283 585
R116 B.n282 B.n281 585
R117 B.n280 B.n279 585
R118 B.n278 B.n277 585
R119 B.n276 B.n275 585
R120 B.n274 B.n273 585
R121 B.n272 B.n271 585
R122 B.n270 B.n269 585
R123 B.n268 B.n267 585
R124 B.n266 B.n265 585
R125 B.n264 B.n263 585
R126 B.n262 B.n261 585
R127 B.n260 B.n259 585
R128 B.n258 B.n257 585
R129 B.n256 B.n255 585
R130 B.n254 B.n253 585
R131 B.n252 B.n251 585
R132 B.n250 B.n249 585
R133 B.n248 B.n247 585
R134 B.n246 B.n245 585
R135 B.n244 B.n243 585
R136 B.n242 B.n241 585
R137 B.n240 B.n239 585
R138 B.n238 B.n237 585
R139 B.n236 B.n235 585
R140 B.n234 B.n233 585
R141 B.n232 B.n231 585
R142 B.n230 B.n229 585
R143 B.n228 B.n227 585
R144 B.n226 B.n225 585
R145 B.n224 B.n223 585
R146 B.n222 B.n221 585
R147 B.n220 B.n219 585
R148 B.n218 B.n217 585
R149 B.n216 B.n215 585
R150 B.n214 B.n213 585
R151 B.n212 B.n211 585
R152 B.n210 B.n209 585
R153 B.n208 B.n207 585
R154 B.n206 B.n205 585
R155 B.n204 B.n203 585
R156 B.n202 B.n201 585
R157 B.n200 B.n199 585
R158 B.n198 B.n197 585
R159 B.n196 B.n195 585
R160 B.n194 B.n193 585
R161 B.n192 B.n191 585
R162 B.n190 B.n189 585
R163 B.n188 B.n187 585
R164 B.n186 B.n185 585
R165 B.n184 B.n183 585
R166 B.n182 B.n181 585
R167 B.n180 B.n179 585
R168 B.n178 B.n177 585
R169 B.n176 B.n175 585
R170 B.n174 B.n173 585
R171 B.n172 B.n171 585
R172 B.n170 B.n169 585
R173 B.n168 B.n167 585
R174 B.n166 B.n165 585
R175 B.n164 B.n163 585
R176 B.n162 B.n161 585
R177 B.n160 B.n159 585
R178 B.n158 B.n157 585
R179 B.n156 B.n155 585
R180 B.n154 B.n153 585
R181 B.n152 B.n151 585
R182 B.n150 B.n149 585
R183 B.n148 B.n147 585
R184 B.n146 B.n145 585
R185 B.n144 B.n143 585
R186 B.n142 B.n141 585
R187 B.n140 B.n139 585
R188 B.n138 B.n137 585
R189 B.n136 B.n135 585
R190 B.n134 B.n133 585
R191 B.n132 B.n131 585
R192 B.n130 B.n129 585
R193 B.n128 B.n127 585
R194 B.n126 B.n125 585
R195 B.n124 B.n123 585
R196 B.n122 B.n121 585
R197 B.n120 B.n119 585
R198 B.n118 B.n117 585
R199 B.n116 B.n115 585
R200 B.n114 B.n113 585
R201 B.n112 B.n111 585
R202 B.n110 B.n109 585
R203 B.n788 B.n41 585
R204 B.n793 B.n41 585
R205 B.n787 B.n40 585
R206 B.n794 B.n40 585
R207 B.n786 B.n785 585
R208 B.n785 B.n36 585
R209 B.n784 B.n35 585
R210 B.n800 B.n35 585
R211 B.n783 B.n34 585
R212 B.n801 B.n34 585
R213 B.n782 B.n33 585
R214 B.n802 B.n33 585
R215 B.n781 B.n780 585
R216 B.n780 B.n29 585
R217 B.n779 B.n28 585
R218 B.n808 B.n28 585
R219 B.n778 B.n27 585
R220 B.n809 B.n27 585
R221 B.n777 B.n26 585
R222 B.n810 B.n26 585
R223 B.n776 B.n775 585
R224 B.n775 B.n25 585
R225 B.n774 B.n21 585
R226 B.n816 B.n21 585
R227 B.n773 B.n20 585
R228 B.n817 B.n20 585
R229 B.n772 B.n19 585
R230 B.t21 B.n19 585
R231 B.n771 B.n770 585
R232 B.n770 B.n15 585
R233 B.n769 B.n14 585
R234 B.n823 B.n14 585
R235 B.n768 B.n13 585
R236 B.n824 B.n13 585
R237 B.n767 B.n12 585
R238 B.n825 B.n12 585
R239 B.n766 B.n765 585
R240 B.n765 B.n11 585
R241 B.n764 B.n7 585
R242 B.n831 B.n7 585
R243 B.n763 B.n6 585
R244 B.n832 B.n6 585
R245 B.n762 B.n5 585
R246 B.n833 B.n5 585
R247 B.n761 B.n760 585
R248 B.n760 B.n4 585
R249 B.n759 B.n350 585
R250 B.n759 B.n758 585
R251 B.n748 B.n351 585
R252 B.n751 B.n351 585
R253 B.n750 B.n749 585
R254 B.n752 B.n750 585
R255 B.n747 B.n356 585
R256 B.n356 B.n355 585
R257 B.n746 B.n745 585
R258 B.n745 B.n744 585
R259 B.n358 B.n357 585
R260 B.n359 B.n358 585
R261 B.n738 B.n737 585
R262 B.t1 B.n738 585
R263 B.n736 B.n364 585
R264 B.n364 B.n363 585
R265 B.n735 B.n734 585
R266 B.n734 B.n733 585
R267 B.n366 B.n365 585
R268 B.n726 B.n366 585
R269 B.n725 B.n724 585
R270 B.n727 B.n725 585
R271 B.n723 B.n371 585
R272 B.n371 B.n370 585
R273 B.n722 B.n721 585
R274 B.n721 B.n720 585
R275 B.n373 B.n372 585
R276 B.n374 B.n373 585
R277 B.n713 B.n712 585
R278 B.n714 B.n713 585
R279 B.n711 B.n378 585
R280 B.n382 B.n378 585
R281 B.n710 B.n709 585
R282 B.n709 B.n708 585
R283 B.n380 B.n379 585
R284 B.n381 B.n380 585
R285 B.n701 B.n700 585
R286 B.n702 B.n701 585
R287 B.n699 B.n387 585
R288 B.n387 B.n386 585
R289 B.n694 B.n693 585
R290 B.n692 B.n450 585
R291 B.n691 B.n449 585
R292 B.n696 B.n449 585
R293 B.n690 B.n689 585
R294 B.n688 B.n687 585
R295 B.n686 B.n685 585
R296 B.n684 B.n683 585
R297 B.n682 B.n681 585
R298 B.n680 B.n679 585
R299 B.n678 B.n677 585
R300 B.n676 B.n675 585
R301 B.n674 B.n673 585
R302 B.n672 B.n671 585
R303 B.n670 B.n669 585
R304 B.n668 B.n667 585
R305 B.n666 B.n665 585
R306 B.n664 B.n663 585
R307 B.n662 B.n661 585
R308 B.n660 B.n659 585
R309 B.n658 B.n657 585
R310 B.n656 B.n655 585
R311 B.n654 B.n653 585
R312 B.n652 B.n651 585
R313 B.n650 B.n649 585
R314 B.n648 B.n647 585
R315 B.n646 B.n645 585
R316 B.n644 B.n643 585
R317 B.n642 B.n641 585
R318 B.n640 B.n639 585
R319 B.n638 B.n637 585
R320 B.n636 B.n635 585
R321 B.n634 B.n633 585
R322 B.n632 B.n631 585
R323 B.n630 B.n629 585
R324 B.n628 B.n627 585
R325 B.n626 B.n625 585
R326 B.n624 B.n623 585
R327 B.n622 B.n621 585
R328 B.n620 B.n619 585
R329 B.n618 B.n617 585
R330 B.n616 B.n615 585
R331 B.n614 B.n613 585
R332 B.n612 B.n611 585
R333 B.n610 B.n609 585
R334 B.n608 B.n607 585
R335 B.n606 B.n605 585
R336 B.n604 B.n603 585
R337 B.n602 B.n601 585
R338 B.n600 B.n599 585
R339 B.n598 B.n597 585
R340 B.n596 B.n595 585
R341 B.n594 B.n593 585
R342 B.n592 B.n591 585
R343 B.n590 B.n589 585
R344 B.n588 B.n587 585
R345 B.n586 B.n585 585
R346 B.n583 B.n582 585
R347 B.n581 B.n580 585
R348 B.n579 B.n578 585
R349 B.n577 B.n576 585
R350 B.n575 B.n574 585
R351 B.n573 B.n572 585
R352 B.n571 B.n570 585
R353 B.n569 B.n568 585
R354 B.n567 B.n566 585
R355 B.n565 B.n564 585
R356 B.n562 B.n561 585
R357 B.n560 B.n559 585
R358 B.n558 B.n557 585
R359 B.n556 B.n555 585
R360 B.n554 B.n553 585
R361 B.n552 B.n551 585
R362 B.n550 B.n549 585
R363 B.n548 B.n547 585
R364 B.n546 B.n545 585
R365 B.n544 B.n543 585
R366 B.n542 B.n541 585
R367 B.n540 B.n539 585
R368 B.n538 B.n537 585
R369 B.n536 B.n535 585
R370 B.n534 B.n533 585
R371 B.n532 B.n531 585
R372 B.n530 B.n529 585
R373 B.n528 B.n527 585
R374 B.n526 B.n525 585
R375 B.n524 B.n523 585
R376 B.n522 B.n521 585
R377 B.n520 B.n519 585
R378 B.n518 B.n517 585
R379 B.n516 B.n515 585
R380 B.n514 B.n513 585
R381 B.n512 B.n511 585
R382 B.n510 B.n509 585
R383 B.n508 B.n507 585
R384 B.n506 B.n505 585
R385 B.n504 B.n503 585
R386 B.n502 B.n501 585
R387 B.n500 B.n499 585
R388 B.n498 B.n497 585
R389 B.n496 B.n495 585
R390 B.n494 B.n493 585
R391 B.n492 B.n491 585
R392 B.n490 B.n489 585
R393 B.n488 B.n487 585
R394 B.n486 B.n485 585
R395 B.n484 B.n483 585
R396 B.n482 B.n481 585
R397 B.n480 B.n479 585
R398 B.n478 B.n477 585
R399 B.n476 B.n475 585
R400 B.n474 B.n473 585
R401 B.n472 B.n471 585
R402 B.n470 B.n469 585
R403 B.n468 B.n467 585
R404 B.n466 B.n465 585
R405 B.n464 B.n463 585
R406 B.n462 B.n461 585
R407 B.n460 B.n459 585
R408 B.n458 B.n457 585
R409 B.n456 B.n455 585
R410 B.n389 B.n388 585
R411 B.n698 B.n697 585
R412 B.n697 B.n696 585
R413 B.n385 B.n384 585
R414 B.n386 B.n385 585
R415 B.n704 B.n703 585
R416 B.n703 B.n702 585
R417 B.n705 B.n383 585
R418 B.n383 B.n381 585
R419 B.n707 B.n706 585
R420 B.n708 B.n707 585
R421 B.n377 B.n376 585
R422 B.n382 B.n377 585
R423 B.n716 B.n715 585
R424 B.n715 B.n714 585
R425 B.n717 B.n375 585
R426 B.n375 B.n374 585
R427 B.n719 B.n718 585
R428 B.n720 B.n719 585
R429 B.n369 B.n368 585
R430 B.n370 B.n369 585
R431 B.n729 B.n728 585
R432 B.n728 B.n727 585
R433 B.n730 B.n367 585
R434 B.n726 B.n367 585
R435 B.n732 B.n731 585
R436 B.n733 B.n732 585
R437 B.n362 B.n361 585
R438 B.n363 B.n362 585
R439 B.n740 B.n739 585
R440 B.n739 B.t1 585
R441 B.n741 B.n360 585
R442 B.n360 B.n359 585
R443 B.n743 B.n742 585
R444 B.n744 B.n743 585
R445 B.n354 B.n353 585
R446 B.n355 B.n354 585
R447 B.n754 B.n753 585
R448 B.n753 B.n752 585
R449 B.n755 B.n352 585
R450 B.n751 B.n352 585
R451 B.n757 B.n756 585
R452 B.n758 B.n757 585
R453 B.n2 B.n0 585
R454 B.n4 B.n2 585
R455 B.n3 B.n1 585
R456 B.n832 B.n3 585
R457 B.n830 B.n829 585
R458 B.n831 B.n830 585
R459 B.n828 B.n8 585
R460 B.n11 B.n8 585
R461 B.n827 B.n826 585
R462 B.n826 B.n825 585
R463 B.n10 B.n9 585
R464 B.n824 B.n10 585
R465 B.n822 B.n821 585
R466 B.n823 B.n822 585
R467 B.n820 B.n16 585
R468 B.n16 B.n15 585
R469 B.n819 B.n818 585
R470 B.n818 B.t21 585
R471 B.n18 B.n17 585
R472 B.n817 B.n18 585
R473 B.n815 B.n814 585
R474 B.n816 B.n815 585
R475 B.n813 B.n22 585
R476 B.n25 B.n22 585
R477 B.n812 B.n811 585
R478 B.n811 B.n810 585
R479 B.n24 B.n23 585
R480 B.n809 B.n24 585
R481 B.n807 B.n806 585
R482 B.n808 B.n807 585
R483 B.n805 B.n30 585
R484 B.n30 B.n29 585
R485 B.n804 B.n803 585
R486 B.n803 B.n802 585
R487 B.n32 B.n31 585
R488 B.n801 B.n32 585
R489 B.n799 B.n798 585
R490 B.n800 B.n799 585
R491 B.n797 B.n37 585
R492 B.n37 B.n36 585
R493 B.n796 B.n795 585
R494 B.n795 B.n794 585
R495 B.n39 B.n38 585
R496 B.n793 B.n39 585
R497 B.n835 B.n834 585
R498 B.n834 B.n833 585
R499 B.n694 B.n385 526.135
R500 B.n109 B.n39 526.135
R501 B.n697 B.n387 526.135
R502 B.n790 B.n41 526.135
R503 B.n792 B.n791 256.663
R504 B.n792 B.n101 256.663
R505 B.n792 B.n100 256.663
R506 B.n792 B.n99 256.663
R507 B.n792 B.n98 256.663
R508 B.n792 B.n97 256.663
R509 B.n792 B.n96 256.663
R510 B.n792 B.n95 256.663
R511 B.n792 B.n94 256.663
R512 B.n792 B.n93 256.663
R513 B.n792 B.n92 256.663
R514 B.n792 B.n91 256.663
R515 B.n792 B.n90 256.663
R516 B.n792 B.n89 256.663
R517 B.n792 B.n88 256.663
R518 B.n792 B.n87 256.663
R519 B.n792 B.n86 256.663
R520 B.n792 B.n85 256.663
R521 B.n792 B.n84 256.663
R522 B.n792 B.n83 256.663
R523 B.n792 B.n82 256.663
R524 B.n792 B.n81 256.663
R525 B.n792 B.n80 256.663
R526 B.n792 B.n79 256.663
R527 B.n792 B.n78 256.663
R528 B.n792 B.n77 256.663
R529 B.n792 B.n76 256.663
R530 B.n792 B.n75 256.663
R531 B.n792 B.n74 256.663
R532 B.n792 B.n73 256.663
R533 B.n792 B.n72 256.663
R534 B.n792 B.n71 256.663
R535 B.n792 B.n70 256.663
R536 B.n792 B.n69 256.663
R537 B.n792 B.n68 256.663
R538 B.n792 B.n67 256.663
R539 B.n792 B.n66 256.663
R540 B.n792 B.n65 256.663
R541 B.n792 B.n64 256.663
R542 B.n792 B.n63 256.663
R543 B.n792 B.n62 256.663
R544 B.n792 B.n61 256.663
R545 B.n792 B.n60 256.663
R546 B.n792 B.n59 256.663
R547 B.n792 B.n58 256.663
R548 B.n792 B.n57 256.663
R549 B.n792 B.n56 256.663
R550 B.n792 B.n55 256.663
R551 B.n792 B.n54 256.663
R552 B.n792 B.n53 256.663
R553 B.n792 B.n52 256.663
R554 B.n792 B.n51 256.663
R555 B.n792 B.n50 256.663
R556 B.n792 B.n49 256.663
R557 B.n792 B.n48 256.663
R558 B.n792 B.n47 256.663
R559 B.n792 B.n46 256.663
R560 B.n792 B.n45 256.663
R561 B.n792 B.n44 256.663
R562 B.n792 B.n43 256.663
R563 B.n792 B.n42 256.663
R564 B.n696 B.n695 256.663
R565 B.n696 B.n390 256.663
R566 B.n696 B.n391 256.663
R567 B.n696 B.n392 256.663
R568 B.n696 B.n393 256.663
R569 B.n696 B.n394 256.663
R570 B.n696 B.n395 256.663
R571 B.n696 B.n396 256.663
R572 B.n696 B.n397 256.663
R573 B.n696 B.n398 256.663
R574 B.n696 B.n399 256.663
R575 B.n696 B.n400 256.663
R576 B.n696 B.n401 256.663
R577 B.n696 B.n402 256.663
R578 B.n696 B.n403 256.663
R579 B.n696 B.n404 256.663
R580 B.n696 B.n405 256.663
R581 B.n696 B.n406 256.663
R582 B.n696 B.n407 256.663
R583 B.n696 B.n408 256.663
R584 B.n696 B.n409 256.663
R585 B.n696 B.n410 256.663
R586 B.n696 B.n411 256.663
R587 B.n696 B.n412 256.663
R588 B.n696 B.n413 256.663
R589 B.n696 B.n414 256.663
R590 B.n696 B.n415 256.663
R591 B.n696 B.n416 256.663
R592 B.n696 B.n417 256.663
R593 B.n696 B.n418 256.663
R594 B.n696 B.n419 256.663
R595 B.n696 B.n420 256.663
R596 B.n696 B.n421 256.663
R597 B.n696 B.n422 256.663
R598 B.n696 B.n423 256.663
R599 B.n696 B.n424 256.663
R600 B.n696 B.n425 256.663
R601 B.n696 B.n426 256.663
R602 B.n696 B.n427 256.663
R603 B.n696 B.n428 256.663
R604 B.n696 B.n429 256.663
R605 B.n696 B.n430 256.663
R606 B.n696 B.n431 256.663
R607 B.n696 B.n432 256.663
R608 B.n696 B.n433 256.663
R609 B.n696 B.n434 256.663
R610 B.n696 B.n435 256.663
R611 B.n696 B.n436 256.663
R612 B.n696 B.n437 256.663
R613 B.n696 B.n438 256.663
R614 B.n696 B.n439 256.663
R615 B.n696 B.n440 256.663
R616 B.n696 B.n441 256.663
R617 B.n696 B.n442 256.663
R618 B.n696 B.n443 256.663
R619 B.n696 B.n444 256.663
R620 B.n696 B.n445 256.663
R621 B.n696 B.n446 256.663
R622 B.n696 B.n447 256.663
R623 B.n696 B.n448 256.663
R624 B.n703 B.n385 163.367
R625 B.n703 B.n383 163.367
R626 B.n707 B.n383 163.367
R627 B.n707 B.n377 163.367
R628 B.n715 B.n377 163.367
R629 B.n715 B.n375 163.367
R630 B.n719 B.n375 163.367
R631 B.n719 B.n369 163.367
R632 B.n728 B.n369 163.367
R633 B.n728 B.n367 163.367
R634 B.n732 B.n367 163.367
R635 B.n732 B.n362 163.367
R636 B.n739 B.n362 163.367
R637 B.n739 B.n360 163.367
R638 B.n743 B.n360 163.367
R639 B.n743 B.n354 163.367
R640 B.n753 B.n354 163.367
R641 B.n753 B.n352 163.367
R642 B.n757 B.n352 163.367
R643 B.n757 B.n2 163.367
R644 B.n834 B.n2 163.367
R645 B.n834 B.n3 163.367
R646 B.n830 B.n3 163.367
R647 B.n830 B.n8 163.367
R648 B.n826 B.n8 163.367
R649 B.n826 B.n10 163.367
R650 B.n822 B.n10 163.367
R651 B.n822 B.n16 163.367
R652 B.n818 B.n16 163.367
R653 B.n818 B.n18 163.367
R654 B.n815 B.n18 163.367
R655 B.n815 B.n22 163.367
R656 B.n811 B.n22 163.367
R657 B.n811 B.n24 163.367
R658 B.n807 B.n24 163.367
R659 B.n807 B.n30 163.367
R660 B.n803 B.n30 163.367
R661 B.n803 B.n32 163.367
R662 B.n799 B.n32 163.367
R663 B.n799 B.n37 163.367
R664 B.n795 B.n37 163.367
R665 B.n795 B.n39 163.367
R666 B.n450 B.n449 163.367
R667 B.n689 B.n449 163.367
R668 B.n687 B.n686 163.367
R669 B.n683 B.n682 163.367
R670 B.n679 B.n678 163.367
R671 B.n675 B.n674 163.367
R672 B.n671 B.n670 163.367
R673 B.n667 B.n666 163.367
R674 B.n663 B.n662 163.367
R675 B.n659 B.n658 163.367
R676 B.n655 B.n654 163.367
R677 B.n651 B.n650 163.367
R678 B.n647 B.n646 163.367
R679 B.n643 B.n642 163.367
R680 B.n639 B.n638 163.367
R681 B.n635 B.n634 163.367
R682 B.n631 B.n630 163.367
R683 B.n627 B.n626 163.367
R684 B.n623 B.n622 163.367
R685 B.n619 B.n618 163.367
R686 B.n615 B.n614 163.367
R687 B.n611 B.n610 163.367
R688 B.n607 B.n606 163.367
R689 B.n603 B.n602 163.367
R690 B.n599 B.n598 163.367
R691 B.n595 B.n594 163.367
R692 B.n591 B.n590 163.367
R693 B.n587 B.n586 163.367
R694 B.n582 B.n581 163.367
R695 B.n578 B.n577 163.367
R696 B.n574 B.n573 163.367
R697 B.n570 B.n569 163.367
R698 B.n566 B.n565 163.367
R699 B.n561 B.n560 163.367
R700 B.n557 B.n556 163.367
R701 B.n553 B.n552 163.367
R702 B.n549 B.n548 163.367
R703 B.n545 B.n544 163.367
R704 B.n541 B.n540 163.367
R705 B.n537 B.n536 163.367
R706 B.n533 B.n532 163.367
R707 B.n529 B.n528 163.367
R708 B.n525 B.n524 163.367
R709 B.n521 B.n520 163.367
R710 B.n517 B.n516 163.367
R711 B.n513 B.n512 163.367
R712 B.n509 B.n508 163.367
R713 B.n505 B.n504 163.367
R714 B.n501 B.n500 163.367
R715 B.n497 B.n496 163.367
R716 B.n493 B.n492 163.367
R717 B.n489 B.n488 163.367
R718 B.n485 B.n484 163.367
R719 B.n481 B.n480 163.367
R720 B.n477 B.n476 163.367
R721 B.n473 B.n472 163.367
R722 B.n469 B.n468 163.367
R723 B.n465 B.n464 163.367
R724 B.n461 B.n460 163.367
R725 B.n457 B.n456 163.367
R726 B.n697 B.n389 163.367
R727 B.n701 B.n387 163.367
R728 B.n701 B.n380 163.367
R729 B.n709 B.n380 163.367
R730 B.n709 B.n378 163.367
R731 B.n713 B.n378 163.367
R732 B.n713 B.n373 163.367
R733 B.n721 B.n373 163.367
R734 B.n721 B.n371 163.367
R735 B.n725 B.n371 163.367
R736 B.n725 B.n366 163.367
R737 B.n734 B.n366 163.367
R738 B.n734 B.n364 163.367
R739 B.n738 B.n364 163.367
R740 B.n738 B.n358 163.367
R741 B.n745 B.n358 163.367
R742 B.n745 B.n356 163.367
R743 B.n750 B.n356 163.367
R744 B.n750 B.n351 163.367
R745 B.n759 B.n351 163.367
R746 B.n760 B.n759 163.367
R747 B.n760 B.n5 163.367
R748 B.n6 B.n5 163.367
R749 B.n7 B.n6 163.367
R750 B.n765 B.n7 163.367
R751 B.n765 B.n12 163.367
R752 B.n13 B.n12 163.367
R753 B.n14 B.n13 163.367
R754 B.n770 B.n14 163.367
R755 B.n770 B.n19 163.367
R756 B.n20 B.n19 163.367
R757 B.n21 B.n20 163.367
R758 B.n775 B.n21 163.367
R759 B.n775 B.n26 163.367
R760 B.n27 B.n26 163.367
R761 B.n28 B.n27 163.367
R762 B.n780 B.n28 163.367
R763 B.n780 B.n33 163.367
R764 B.n34 B.n33 163.367
R765 B.n35 B.n34 163.367
R766 B.n785 B.n35 163.367
R767 B.n785 B.n40 163.367
R768 B.n41 B.n40 163.367
R769 B.n113 B.n112 163.367
R770 B.n117 B.n116 163.367
R771 B.n121 B.n120 163.367
R772 B.n125 B.n124 163.367
R773 B.n129 B.n128 163.367
R774 B.n133 B.n132 163.367
R775 B.n137 B.n136 163.367
R776 B.n141 B.n140 163.367
R777 B.n145 B.n144 163.367
R778 B.n149 B.n148 163.367
R779 B.n153 B.n152 163.367
R780 B.n157 B.n156 163.367
R781 B.n161 B.n160 163.367
R782 B.n165 B.n164 163.367
R783 B.n169 B.n168 163.367
R784 B.n173 B.n172 163.367
R785 B.n177 B.n176 163.367
R786 B.n181 B.n180 163.367
R787 B.n185 B.n184 163.367
R788 B.n189 B.n188 163.367
R789 B.n193 B.n192 163.367
R790 B.n197 B.n196 163.367
R791 B.n201 B.n200 163.367
R792 B.n205 B.n204 163.367
R793 B.n209 B.n208 163.367
R794 B.n213 B.n212 163.367
R795 B.n217 B.n216 163.367
R796 B.n221 B.n220 163.367
R797 B.n225 B.n224 163.367
R798 B.n229 B.n228 163.367
R799 B.n233 B.n232 163.367
R800 B.n237 B.n236 163.367
R801 B.n241 B.n240 163.367
R802 B.n245 B.n244 163.367
R803 B.n249 B.n248 163.367
R804 B.n253 B.n252 163.367
R805 B.n257 B.n256 163.367
R806 B.n261 B.n260 163.367
R807 B.n265 B.n264 163.367
R808 B.n269 B.n268 163.367
R809 B.n273 B.n272 163.367
R810 B.n277 B.n276 163.367
R811 B.n281 B.n280 163.367
R812 B.n285 B.n284 163.367
R813 B.n289 B.n288 163.367
R814 B.n293 B.n292 163.367
R815 B.n297 B.n296 163.367
R816 B.n301 B.n300 163.367
R817 B.n305 B.n304 163.367
R818 B.n309 B.n308 163.367
R819 B.n313 B.n312 163.367
R820 B.n317 B.n316 163.367
R821 B.n321 B.n320 163.367
R822 B.n325 B.n324 163.367
R823 B.n329 B.n328 163.367
R824 B.n333 B.n332 163.367
R825 B.n337 B.n336 163.367
R826 B.n341 B.n340 163.367
R827 B.n345 B.n344 163.367
R828 B.n347 B.n102 163.367
R829 B.n453 B.t10 85.1511
R830 B.n103 B.t13 85.1511
R831 B.n451 B.t17 85.1284
R832 B.n106 B.t19 85.1284
R833 B.n695 B.n694 71.676
R834 B.n689 B.n390 71.676
R835 B.n686 B.n391 71.676
R836 B.n682 B.n392 71.676
R837 B.n678 B.n393 71.676
R838 B.n674 B.n394 71.676
R839 B.n670 B.n395 71.676
R840 B.n666 B.n396 71.676
R841 B.n662 B.n397 71.676
R842 B.n658 B.n398 71.676
R843 B.n654 B.n399 71.676
R844 B.n650 B.n400 71.676
R845 B.n646 B.n401 71.676
R846 B.n642 B.n402 71.676
R847 B.n638 B.n403 71.676
R848 B.n634 B.n404 71.676
R849 B.n630 B.n405 71.676
R850 B.n626 B.n406 71.676
R851 B.n622 B.n407 71.676
R852 B.n618 B.n408 71.676
R853 B.n614 B.n409 71.676
R854 B.n610 B.n410 71.676
R855 B.n606 B.n411 71.676
R856 B.n602 B.n412 71.676
R857 B.n598 B.n413 71.676
R858 B.n594 B.n414 71.676
R859 B.n590 B.n415 71.676
R860 B.n586 B.n416 71.676
R861 B.n581 B.n417 71.676
R862 B.n577 B.n418 71.676
R863 B.n573 B.n419 71.676
R864 B.n569 B.n420 71.676
R865 B.n565 B.n421 71.676
R866 B.n560 B.n422 71.676
R867 B.n556 B.n423 71.676
R868 B.n552 B.n424 71.676
R869 B.n548 B.n425 71.676
R870 B.n544 B.n426 71.676
R871 B.n540 B.n427 71.676
R872 B.n536 B.n428 71.676
R873 B.n532 B.n429 71.676
R874 B.n528 B.n430 71.676
R875 B.n524 B.n431 71.676
R876 B.n520 B.n432 71.676
R877 B.n516 B.n433 71.676
R878 B.n512 B.n434 71.676
R879 B.n508 B.n435 71.676
R880 B.n504 B.n436 71.676
R881 B.n500 B.n437 71.676
R882 B.n496 B.n438 71.676
R883 B.n492 B.n439 71.676
R884 B.n488 B.n440 71.676
R885 B.n484 B.n441 71.676
R886 B.n480 B.n442 71.676
R887 B.n476 B.n443 71.676
R888 B.n472 B.n444 71.676
R889 B.n468 B.n445 71.676
R890 B.n464 B.n446 71.676
R891 B.n460 B.n447 71.676
R892 B.n456 B.n448 71.676
R893 B.n109 B.n42 71.676
R894 B.n113 B.n43 71.676
R895 B.n117 B.n44 71.676
R896 B.n121 B.n45 71.676
R897 B.n125 B.n46 71.676
R898 B.n129 B.n47 71.676
R899 B.n133 B.n48 71.676
R900 B.n137 B.n49 71.676
R901 B.n141 B.n50 71.676
R902 B.n145 B.n51 71.676
R903 B.n149 B.n52 71.676
R904 B.n153 B.n53 71.676
R905 B.n157 B.n54 71.676
R906 B.n161 B.n55 71.676
R907 B.n165 B.n56 71.676
R908 B.n169 B.n57 71.676
R909 B.n173 B.n58 71.676
R910 B.n177 B.n59 71.676
R911 B.n181 B.n60 71.676
R912 B.n185 B.n61 71.676
R913 B.n189 B.n62 71.676
R914 B.n193 B.n63 71.676
R915 B.n197 B.n64 71.676
R916 B.n201 B.n65 71.676
R917 B.n205 B.n66 71.676
R918 B.n209 B.n67 71.676
R919 B.n213 B.n68 71.676
R920 B.n217 B.n69 71.676
R921 B.n221 B.n70 71.676
R922 B.n225 B.n71 71.676
R923 B.n229 B.n72 71.676
R924 B.n233 B.n73 71.676
R925 B.n237 B.n74 71.676
R926 B.n241 B.n75 71.676
R927 B.n245 B.n76 71.676
R928 B.n249 B.n77 71.676
R929 B.n253 B.n78 71.676
R930 B.n257 B.n79 71.676
R931 B.n261 B.n80 71.676
R932 B.n265 B.n81 71.676
R933 B.n269 B.n82 71.676
R934 B.n273 B.n83 71.676
R935 B.n277 B.n84 71.676
R936 B.n281 B.n85 71.676
R937 B.n285 B.n86 71.676
R938 B.n289 B.n87 71.676
R939 B.n293 B.n88 71.676
R940 B.n297 B.n89 71.676
R941 B.n301 B.n90 71.676
R942 B.n305 B.n91 71.676
R943 B.n309 B.n92 71.676
R944 B.n313 B.n93 71.676
R945 B.n317 B.n94 71.676
R946 B.n321 B.n95 71.676
R947 B.n325 B.n96 71.676
R948 B.n329 B.n97 71.676
R949 B.n333 B.n98 71.676
R950 B.n337 B.n99 71.676
R951 B.n341 B.n100 71.676
R952 B.n345 B.n101 71.676
R953 B.n791 B.n102 71.676
R954 B.n791 B.n790 71.676
R955 B.n347 B.n101 71.676
R956 B.n344 B.n100 71.676
R957 B.n340 B.n99 71.676
R958 B.n336 B.n98 71.676
R959 B.n332 B.n97 71.676
R960 B.n328 B.n96 71.676
R961 B.n324 B.n95 71.676
R962 B.n320 B.n94 71.676
R963 B.n316 B.n93 71.676
R964 B.n312 B.n92 71.676
R965 B.n308 B.n91 71.676
R966 B.n304 B.n90 71.676
R967 B.n300 B.n89 71.676
R968 B.n296 B.n88 71.676
R969 B.n292 B.n87 71.676
R970 B.n288 B.n86 71.676
R971 B.n284 B.n85 71.676
R972 B.n280 B.n84 71.676
R973 B.n276 B.n83 71.676
R974 B.n272 B.n82 71.676
R975 B.n268 B.n81 71.676
R976 B.n264 B.n80 71.676
R977 B.n260 B.n79 71.676
R978 B.n256 B.n78 71.676
R979 B.n252 B.n77 71.676
R980 B.n248 B.n76 71.676
R981 B.n244 B.n75 71.676
R982 B.n240 B.n74 71.676
R983 B.n236 B.n73 71.676
R984 B.n232 B.n72 71.676
R985 B.n228 B.n71 71.676
R986 B.n224 B.n70 71.676
R987 B.n220 B.n69 71.676
R988 B.n216 B.n68 71.676
R989 B.n212 B.n67 71.676
R990 B.n208 B.n66 71.676
R991 B.n204 B.n65 71.676
R992 B.n200 B.n64 71.676
R993 B.n196 B.n63 71.676
R994 B.n192 B.n62 71.676
R995 B.n188 B.n61 71.676
R996 B.n184 B.n60 71.676
R997 B.n180 B.n59 71.676
R998 B.n176 B.n58 71.676
R999 B.n172 B.n57 71.676
R1000 B.n168 B.n56 71.676
R1001 B.n164 B.n55 71.676
R1002 B.n160 B.n54 71.676
R1003 B.n156 B.n53 71.676
R1004 B.n152 B.n52 71.676
R1005 B.n148 B.n51 71.676
R1006 B.n144 B.n50 71.676
R1007 B.n140 B.n49 71.676
R1008 B.n136 B.n48 71.676
R1009 B.n132 B.n47 71.676
R1010 B.n128 B.n46 71.676
R1011 B.n124 B.n45 71.676
R1012 B.n120 B.n44 71.676
R1013 B.n116 B.n43 71.676
R1014 B.n112 B.n42 71.676
R1015 B.n695 B.n450 71.676
R1016 B.n687 B.n390 71.676
R1017 B.n683 B.n391 71.676
R1018 B.n679 B.n392 71.676
R1019 B.n675 B.n393 71.676
R1020 B.n671 B.n394 71.676
R1021 B.n667 B.n395 71.676
R1022 B.n663 B.n396 71.676
R1023 B.n659 B.n397 71.676
R1024 B.n655 B.n398 71.676
R1025 B.n651 B.n399 71.676
R1026 B.n647 B.n400 71.676
R1027 B.n643 B.n401 71.676
R1028 B.n639 B.n402 71.676
R1029 B.n635 B.n403 71.676
R1030 B.n631 B.n404 71.676
R1031 B.n627 B.n405 71.676
R1032 B.n623 B.n406 71.676
R1033 B.n619 B.n407 71.676
R1034 B.n615 B.n408 71.676
R1035 B.n611 B.n409 71.676
R1036 B.n607 B.n410 71.676
R1037 B.n603 B.n411 71.676
R1038 B.n599 B.n412 71.676
R1039 B.n595 B.n413 71.676
R1040 B.n591 B.n414 71.676
R1041 B.n587 B.n415 71.676
R1042 B.n582 B.n416 71.676
R1043 B.n578 B.n417 71.676
R1044 B.n574 B.n418 71.676
R1045 B.n570 B.n419 71.676
R1046 B.n566 B.n420 71.676
R1047 B.n561 B.n421 71.676
R1048 B.n557 B.n422 71.676
R1049 B.n553 B.n423 71.676
R1050 B.n549 B.n424 71.676
R1051 B.n545 B.n425 71.676
R1052 B.n541 B.n426 71.676
R1053 B.n537 B.n427 71.676
R1054 B.n533 B.n428 71.676
R1055 B.n529 B.n429 71.676
R1056 B.n525 B.n430 71.676
R1057 B.n521 B.n431 71.676
R1058 B.n517 B.n432 71.676
R1059 B.n513 B.n433 71.676
R1060 B.n509 B.n434 71.676
R1061 B.n505 B.n435 71.676
R1062 B.n501 B.n436 71.676
R1063 B.n497 B.n437 71.676
R1064 B.n493 B.n438 71.676
R1065 B.n489 B.n439 71.676
R1066 B.n485 B.n440 71.676
R1067 B.n481 B.n441 71.676
R1068 B.n477 B.n442 71.676
R1069 B.n473 B.n443 71.676
R1070 B.n469 B.n444 71.676
R1071 B.n465 B.n445 71.676
R1072 B.n461 B.n446 71.676
R1073 B.n457 B.n447 71.676
R1074 B.n448 B.n389 71.676
R1075 B.n454 B.t9 68.2784
R1076 B.n104 B.t14 68.2784
R1077 B.n452 B.t16 68.2556
R1078 B.n107 B.t20 68.2556
R1079 B.n563 B.n454 59.5399
R1080 B.n584 B.n452 59.5399
R1081 B.n108 B.n107 59.5399
R1082 B.n105 B.n104 59.5399
R1083 B.n696 B.n386 57.6489
R1084 B.n793 B.n792 57.6489
R1085 B.n110 B.n38 34.1859
R1086 B.n789 B.n788 34.1859
R1087 B.n699 B.n698 34.1859
R1088 B.n693 B.n384 34.1859
R1089 B.n702 B.n386 33.5055
R1090 B.n702 B.n381 33.5055
R1091 B.n708 B.n381 33.5055
R1092 B.n708 B.n382 33.5055
R1093 B.n714 B.n374 33.5055
R1094 B.n720 B.n374 33.5055
R1095 B.n720 B.n370 33.5055
R1096 B.n727 B.n370 33.5055
R1097 B.n727 B.n726 33.5055
R1098 B.n733 B.n363 33.5055
R1099 B.t1 B.n363 33.5055
R1100 B.t1 B.n359 33.5055
R1101 B.n744 B.n359 33.5055
R1102 B.n752 B.n355 33.5055
R1103 B.n752 B.n751 33.5055
R1104 B.n758 B.n4 33.5055
R1105 B.n833 B.n4 33.5055
R1106 B.n833 B.n832 33.5055
R1107 B.n832 B.n831 33.5055
R1108 B.n825 B.n11 33.5055
R1109 B.n825 B.n824 33.5055
R1110 B.n823 B.n15 33.5055
R1111 B.t21 B.n15 33.5055
R1112 B.t21 B.n817 33.5055
R1113 B.n817 B.n816 33.5055
R1114 B.n810 B.n25 33.5055
R1115 B.n810 B.n809 33.5055
R1116 B.n809 B.n808 33.5055
R1117 B.n808 B.n29 33.5055
R1118 B.n802 B.n29 33.5055
R1119 B.n801 B.n800 33.5055
R1120 B.n800 B.n36 33.5055
R1121 B.n794 B.n36 33.5055
R1122 B.n794 B.n793 33.5055
R1123 B.n758 B.t2 29.5638
R1124 B.n831 B.t5 29.5638
R1125 B.n382 B.t8 22.6657
R1126 B.t12 B.n801 22.6657
R1127 B.n733 B.t4 18.7239
R1128 B.n744 B.t0 18.7239
R1129 B.t6 B.n823 18.7239
R1130 B.n816 B.t3 18.7239
R1131 B B.n835 18.0485
R1132 B.n454 B.n453 16.8732
R1133 B.n452 B.n451 16.8732
R1134 B.n107 B.n106 16.8732
R1135 B.n104 B.n103 16.8732
R1136 B.n726 B.t4 14.7821
R1137 B.t0 B.n355 14.7821
R1138 B.n824 B.t6 14.7821
R1139 B.n25 B.t3 14.7821
R1140 B.n714 B.t8 10.8404
R1141 B.n802 B.t12 10.8404
R1142 B.n111 B.n110 10.6151
R1143 B.n114 B.n111 10.6151
R1144 B.n115 B.n114 10.6151
R1145 B.n118 B.n115 10.6151
R1146 B.n119 B.n118 10.6151
R1147 B.n122 B.n119 10.6151
R1148 B.n123 B.n122 10.6151
R1149 B.n126 B.n123 10.6151
R1150 B.n127 B.n126 10.6151
R1151 B.n130 B.n127 10.6151
R1152 B.n131 B.n130 10.6151
R1153 B.n134 B.n131 10.6151
R1154 B.n135 B.n134 10.6151
R1155 B.n138 B.n135 10.6151
R1156 B.n139 B.n138 10.6151
R1157 B.n142 B.n139 10.6151
R1158 B.n143 B.n142 10.6151
R1159 B.n146 B.n143 10.6151
R1160 B.n147 B.n146 10.6151
R1161 B.n150 B.n147 10.6151
R1162 B.n151 B.n150 10.6151
R1163 B.n154 B.n151 10.6151
R1164 B.n155 B.n154 10.6151
R1165 B.n158 B.n155 10.6151
R1166 B.n159 B.n158 10.6151
R1167 B.n162 B.n159 10.6151
R1168 B.n163 B.n162 10.6151
R1169 B.n166 B.n163 10.6151
R1170 B.n167 B.n166 10.6151
R1171 B.n170 B.n167 10.6151
R1172 B.n171 B.n170 10.6151
R1173 B.n174 B.n171 10.6151
R1174 B.n175 B.n174 10.6151
R1175 B.n178 B.n175 10.6151
R1176 B.n179 B.n178 10.6151
R1177 B.n182 B.n179 10.6151
R1178 B.n183 B.n182 10.6151
R1179 B.n186 B.n183 10.6151
R1180 B.n187 B.n186 10.6151
R1181 B.n190 B.n187 10.6151
R1182 B.n191 B.n190 10.6151
R1183 B.n194 B.n191 10.6151
R1184 B.n195 B.n194 10.6151
R1185 B.n198 B.n195 10.6151
R1186 B.n199 B.n198 10.6151
R1187 B.n202 B.n199 10.6151
R1188 B.n203 B.n202 10.6151
R1189 B.n206 B.n203 10.6151
R1190 B.n207 B.n206 10.6151
R1191 B.n210 B.n207 10.6151
R1192 B.n211 B.n210 10.6151
R1193 B.n214 B.n211 10.6151
R1194 B.n215 B.n214 10.6151
R1195 B.n218 B.n215 10.6151
R1196 B.n219 B.n218 10.6151
R1197 B.n223 B.n222 10.6151
R1198 B.n226 B.n223 10.6151
R1199 B.n227 B.n226 10.6151
R1200 B.n230 B.n227 10.6151
R1201 B.n231 B.n230 10.6151
R1202 B.n234 B.n231 10.6151
R1203 B.n235 B.n234 10.6151
R1204 B.n238 B.n235 10.6151
R1205 B.n239 B.n238 10.6151
R1206 B.n243 B.n242 10.6151
R1207 B.n246 B.n243 10.6151
R1208 B.n247 B.n246 10.6151
R1209 B.n250 B.n247 10.6151
R1210 B.n251 B.n250 10.6151
R1211 B.n254 B.n251 10.6151
R1212 B.n255 B.n254 10.6151
R1213 B.n258 B.n255 10.6151
R1214 B.n259 B.n258 10.6151
R1215 B.n262 B.n259 10.6151
R1216 B.n263 B.n262 10.6151
R1217 B.n266 B.n263 10.6151
R1218 B.n267 B.n266 10.6151
R1219 B.n270 B.n267 10.6151
R1220 B.n271 B.n270 10.6151
R1221 B.n274 B.n271 10.6151
R1222 B.n275 B.n274 10.6151
R1223 B.n278 B.n275 10.6151
R1224 B.n279 B.n278 10.6151
R1225 B.n282 B.n279 10.6151
R1226 B.n283 B.n282 10.6151
R1227 B.n286 B.n283 10.6151
R1228 B.n287 B.n286 10.6151
R1229 B.n290 B.n287 10.6151
R1230 B.n291 B.n290 10.6151
R1231 B.n294 B.n291 10.6151
R1232 B.n295 B.n294 10.6151
R1233 B.n298 B.n295 10.6151
R1234 B.n299 B.n298 10.6151
R1235 B.n302 B.n299 10.6151
R1236 B.n303 B.n302 10.6151
R1237 B.n306 B.n303 10.6151
R1238 B.n307 B.n306 10.6151
R1239 B.n310 B.n307 10.6151
R1240 B.n311 B.n310 10.6151
R1241 B.n314 B.n311 10.6151
R1242 B.n315 B.n314 10.6151
R1243 B.n318 B.n315 10.6151
R1244 B.n319 B.n318 10.6151
R1245 B.n322 B.n319 10.6151
R1246 B.n323 B.n322 10.6151
R1247 B.n326 B.n323 10.6151
R1248 B.n327 B.n326 10.6151
R1249 B.n330 B.n327 10.6151
R1250 B.n331 B.n330 10.6151
R1251 B.n334 B.n331 10.6151
R1252 B.n335 B.n334 10.6151
R1253 B.n338 B.n335 10.6151
R1254 B.n339 B.n338 10.6151
R1255 B.n342 B.n339 10.6151
R1256 B.n343 B.n342 10.6151
R1257 B.n346 B.n343 10.6151
R1258 B.n348 B.n346 10.6151
R1259 B.n349 B.n348 10.6151
R1260 B.n789 B.n349 10.6151
R1261 B.n700 B.n699 10.6151
R1262 B.n700 B.n379 10.6151
R1263 B.n710 B.n379 10.6151
R1264 B.n711 B.n710 10.6151
R1265 B.n712 B.n711 10.6151
R1266 B.n712 B.n372 10.6151
R1267 B.n722 B.n372 10.6151
R1268 B.n723 B.n722 10.6151
R1269 B.n724 B.n723 10.6151
R1270 B.n724 B.n365 10.6151
R1271 B.n735 B.n365 10.6151
R1272 B.n736 B.n735 10.6151
R1273 B.n737 B.n736 10.6151
R1274 B.n737 B.n357 10.6151
R1275 B.n746 B.n357 10.6151
R1276 B.n747 B.n746 10.6151
R1277 B.n749 B.n747 10.6151
R1278 B.n749 B.n748 10.6151
R1279 B.n748 B.n350 10.6151
R1280 B.n761 B.n350 10.6151
R1281 B.n762 B.n761 10.6151
R1282 B.n763 B.n762 10.6151
R1283 B.n764 B.n763 10.6151
R1284 B.n766 B.n764 10.6151
R1285 B.n767 B.n766 10.6151
R1286 B.n768 B.n767 10.6151
R1287 B.n769 B.n768 10.6151
R1288 B.n771 B.n769 10.6151
R1289 B.n772 B.n771 10.6151
R1290 B.n773 B.n772 10.6151
R1291 B.n774 B.n773 10.6151
R1292 B.n776 B.n774 10.6151
R1293 B.n777 B.n776 10.6151
R1294 B.n778 B.n777 10.6151
R1295 B.n779 B.n778 10.6151
R1296 B.n781 B.n779 10.6151
R1297 B.n782 B.n781 10.6151
R1298 B.n783 B.n782 10.6151
R1299 B.n784 B.n783 10.6151
R1300 B.n786 B.n784 10.6151
R1301 B.n787 B.n786 10.6151
R1302 B.n788 B.n787 10.6151
R1303 B.n693 B.n692 10.6151
R1304 B.n692 B.n691 10.6151
R1305 B.n691 B.n690 10.6151
R1306 B.n690 B.n688 10.6151
R1307 B.n688 B.n685 10.6151
R1308 B.n685 B.n684 10.6151
R1309 B.n684 B.n681 10.6151
R1310 B.n681 B.n680 10.6151
R1311 B.n680 B.n677 10.6151
R1312 B.n677 B.n676 10.6151
R1313 B.n676 B.n673 10.6151
R1314 B.n673 B.n672 10.6151
R1315 B.n672 B.n669 10.6151
R1316 B.n669 B.n668 10.6151
R1317 B.n668 B.n665 10.6151
R1318 B.n665 B.n664 10.6151
R1319 B.n664 B.n661 10.6151
R1320 B.n661 B.n660 10.6151
R1321 B.n660 B.n657 10.6151
R1322 B.n657 B.n656 10.6151
R1323 B.n656 B.n653 10.6151
R1324 B.n653 B.n652 10.6151
R1325 B.n652 B.n649 10.6151
R1326 B.n649 B.n648 10.6151
R1327 B.n648 B.n645 10.6151
R1328 B.n645 B.n644 10.6151
R1329 B.n644 B.n641 10.6151
R1330 B.n641 B.n640 10.6151
R1331 B.n640 B.n637 10.6151
R1332 B.n637 B.n636 10.6151
R1333 B.n636 B.n633 10.6151
R1334 B.n633 B.n632 10.6151
R1335 B.n632 B.n629 10.6151
R1336 B.n629 B.n628 10.6151
R1337 B.n628 B.n625 10.6151
R1338 B.n625 B.n624 10.6151
R1339 B.n624 B.n621 10.6151
R1340 B.n621 B.n620 10.6151
R1341 B.n620 B.n617 10.6151
R1342 B.n617 B.n616 10.6151
R1343 B.n616 B.n613 10.6151
R1344 B.n613 B.n612 10.6151
R1345 B.n612 B.n609 10.6151
R1346 B.n609 B.n608 10.6151
R1347 B.n608 B.n605 10.6151
R1348 B.n605 B.n604 10.6151
R1349 B.n604 B.n601 10.6151
R1350 B.n601 B.n600 10.6151
R1351 B.n600 B.n597 10.6151
R1352 B.n597 B.n596 10.6151
R1353 B.n596 B.n593 10.6151
R1354 B.n593 B.n592 10.6151
R1355 B.n592 B.n589 10.6151
R1356 B.n589 B.n588 10.6151
R1357 B.n588 B.n585 10.6151
R1358 B.n583 B.n580 10.6151
R1359 B.n580 B.n579 10.6151
R1360 B.n579 B.n576 10.6151
R1361 B.n576 B.n575 10.6151
R1362 B.n575 B.n572 10.6151
R1363 B.n572 B.n571 10.6151
R1364 B.n571 B.n568 10.6151
R1365 B.n568 B.n567 10.6151
R1366 B.n567 B.n564 10.6151
R1367 B.n562 B.n559 10.6151
R1368 B.n559 B.n558 10.6151
R1369 B.n558 B.n555 10.6151
R1370 B.n555 B.n554 10.6151
R1371 B.n554 B.n551 10.6151
R1372 B.n551 B.n550 10.6151
R1373 B.n550 B.n547 10.6151
R1374 B.n547 B.n546 10.6151
R1375 B.n546 B.n543 10.6151
R1376 B.n543 B.n542 10.6151
R1377 B.n542 B.n539 10.6151
R1378 B.n539 B.n538 10.6151
R1379 B.n538 B.n535 10.6151
R1380 B.n535 B.n534 10.6151
R1381 B.n534 B.n531 10.6151
R1382 B.n531 B.n530 10.6151
R1383 B.n530 B.n527 10.6151
R1384 B.n527 B.n526 10.6151
R1385 B.n526 B.n523 10.6151
R1386 B.n523 B.n522 10.6151
R1387 B.n522 B.n519 10.6151
R1388 B.n519 B.n518 10.6151
R1389 B.n518 B.n515 10.6151
R1390 B.n515 B.n514 10.6151
R1391 B.n514 B.n511 10.6151
R1392 B.n511 B.n510 10.6151
R1393 B.n510 B.n507 10.6151
R1394 B.n507 B.n506 10.6151
R1395 B.n506 B.n503 10.6151
R1396 B.n503 B.n502 10.6151
R1397 B.n502 B.n499 10.6151
R1398 B.n499 B.n498 10.6151
R1399 B.n498 B.n495 10.6151
R1400 B.n495 B.n494 10.6151
R1401 B.n494 B.n491 10.6151
R1402 B.n491 B.n490 10.6151
R1403 B.n490 B.n487 10.6151
R1404 B.n487 B.n486 10.6151
R1405 B.n486 B.n483 10.6151
R1406 B.n483 B.n482 10.6151
R1407 B.n482 B.n479 10.6151
R1408 B.n479 B.n478 10.6151
R1409 B.n478 B.n475 10.6151
R1410 B.n475 B.n474 10.6151
R1411 B.n474 B.n471 10.6151
R1412 B.n471 B.n470 10.6151
R1413 B.n470 B.n467 10.6151
R1414 B.n467 B.n466 10.6151
R1415 B.n466 B.n463 10.6151
R1416 B.n463 B.n462 10.6151
R1417 B.n462 B.n459 10.6151
R1418 B.n459 B.n458 10.6151
R1419 B.n458 B.n455 10.6151
R1420 B.n455 B.n388 10.6151
R1421 B.n698 B.n388 10.6151
R1422 B.n704 B.n384 10.6151
R1423 B.n705 B.n704 10.6151
R1424 B.n706 B.n705 10.6151
R1425 B.n706 B.n376 10.6151
R1426 B.n716 B.n376 10.6151
R1427 B.n717 B.n716 10.6151
R1428 B.n718 B.n717 10.6151
R1429 B.n718 B.n368 10.6151
R1430 B.n729 B.n368 10.6151
R1431 B.n730 B.n729 10.6151
R1432 B.n731 B.n730 10.6151
R1433 B.n731 B.n361 10.6151
R1434 B.n740 B.n361 10.6151
R1435 B.n741 B.n740 10.6151
R1436 B.n742 B.n741 10.6151
R1437 B.n742 B.n353 10.6151
R1438 B.n754 B.n353 10.6151
R1439 B.n755 B.n754 10.6151
R1440 B.n756 B.n755 10.6151
R1441 B.n756 B.n0 10.6151
R1442 B.n829 B.n1 10.6151
R1443 B.n829 B.n828 10.6151
R1444 B.n828 B.n827 10.6151
R1445 B.n827 B.n9 10.6151
R1446 B.n821 B.n9 10.6151
R1447 B.n821 B.n820 10.6151
R1448 B.n820 B.n819 10.6151
R1449 B.n819 B.n17 10.6151
R1450 B.n814 B.n17 10.6151
R1451 B.n814 B.n813 10.6151
R1452 B.n813 B.n812 10.6151
R1453 B.n812 B.n23 10.6151
R1454 B.n806 B.n23 10.6151
R1455 B.n806 B.n805 10.6151
R1456 B.n805 B.n804 10.6151
R1457 B.n804 B.n31 10.6151
R1458 B.n798 B.n31 10.6151
R1459 B.n798 B.n797 10.6151
R1460 B.n797 B.n796 10.6151
R1461 B.n796 B.n38 10.6151
R1462 B.n219 B.n108 9.36635
R1463 B.n242 B.n105 9.36635
R1464 B.n585 B.n584 9.36635
R1465 B.n563 B.n562 9.36635
R1466 B.n751 B.t2 3.94227
R1467 B.n11 B.t5 3.94227
R1468 B.n835 B.n0 2.81026
R1469 B.n835 B.n1 2.81026
R1470 B.n222 B.n108 1.24928
R1471 B.n239 B.n105 1.24928
R1472 B.n584 B.n583 1.24928
R1473 B.n564 B.n563 1.24928
R1474 VP.n4 VP.t4 859.521
R1475 VP.n11 VP.t6 834.129
R1476 VP.n1 VP.t2 834.129
R1477 VP.n16 VP.t5 834.129
R1478 VP.n18 VP.t1 834.129
R1479 VP.n8 VP.t7 834.129
R1480 VP.n6 VP.t0 834.129
R1481 VP.n5 VP.t3 834.129
R1482 VP.n19 VP.n18 161.3
R1483 VP.n6 VP.n3 161.3
R1484 VP.n7 VP.n2 161.3
R1485 VP.n9 VP.n8 161.3
R1486 VP.n17 VP.n0 161.3
R1487 VP.n16 VP.n15 161.3
R1488 VP.n14 VP.n1 161.3
R1489 VP.n13 VP.n12 161.3
R1490 VP.n11 VP.n10 161.3
R1491 VP.n16 VP.n1 48.2005
R1492 VP.n6 VP.n5 48.2005
R1493 VP.n10 VP.n9 45.0384
R1494 VP.n4 VP.n3 45.0031
R1495 VP.n12 VP.n11 41.6278
R1496 VP.n18 VP.n17 41.6278
R1497 VP.n8 VP.n7 41.6278
R1498 VP.n5 VP.n4 15.6319
R1499 VP.n12 VP.n1 6.57323
R1500 VP.n17 VP.n16 6.57323
R1501 VP.n7 VP.n6 6.57323
R1502 VP.n3 VP.n2 0.189894
R1503 VP.n9 VP.n2 0.189894
R1504 VP.n13 VP.n10 0.189894
R1505 VP.n14 VP.n13 0.189894
R1506 VP.n15 VP.n14 0.189894
R1507 VP.n15 VP.n0 0.189894
R1508 VP.n19 VP.n0 0.189894
R1509 VP VP.n19 0.0516364
R1510 VDD1 VDD1.n0 59.0019
R1511 VDD1.n3 VDD1.n2 58.8881
R1512 VDD1.n3 VDD1.n1 58.8881
R1513 VDD1.n5 VDD1.n4 58.5686
R1514 VDD1.n5 VDD1.n3 42.3716
R1515 VDD1.n4 VDD1.t7 1.16179
R1516 VDD1.n4 VDD1.t0 1.16179
R1517 VDD1.n0 VDD1.t3 1.16179
R1518 VDD1.n0 VDD1.t4 1.16179
R1519 VDD1.n2 VDD1.t2 1.16179
R1520 VDD1.n2 VDD1.t6 1.16179
R1521 VDD1.n1 VDD1.t1 1.16179
R1522 VDD1.n1 VDD1.t5 1.16179
R1523 VDD1 VDD1.n5 0.31731
C0 VDD1 VDD2 0.746651f
C1 VDD2 VN 6.64184f
C2 VDD1 VP 6.79394f
C3 VDD2 VTAIL 16.9394f
C4 VP VN 6.08172f
C5 VDD1 VN 0.147865f
C6 VTAIL VP 6.14427f
C7 VDD1 VTAIL 16.8988f
C8 VTAIL VN 6.13016f
C9 VDD2 VP 0.300326f
C10 VDD2 B 3.740525f
C11 VDD1 B 3.960294f
C12 VTAIL B 11.575352f
C13 VN B 8.68567f
C14 VP B 6.349529f
C15 VDD1.t3 B 0.390972f
C16 VDD1.t4 B 0.390972f
C17 VDD1.n0 B 3.55302f
C18 VDD1.t1 B 0.390972f
C19 VDD1.t5 B 0.390972f
C20 VDD1.n1 B 3.55227f
C21 VDD1.t2 B 0.390972f
C22 VDD1.t6 B 0.390972f
C23 VDD1.n2 B 3.55227f
C24 VDD1.n3 B 2.84645f
C25 VDD1.t7 B 0.390972f
C26 VDD1.t0 B 0.390972f
C27 VDD1.n4 B 3.55032f
C28 VDD1.n5 B 3.08448f
C29 VP.n0 B 0.048309f
C30 VP.t2 B 1.26209f
C31 VP.n1 B 0.483851f
C32 VP.n2 B 0.048309f
C33 VP.t7 B 1.26209f
C34 VP.t0 B 1.26209f
C35 VP.n3 B 0.196749f
C36 VP.t3 B 1.26209f
C37 VP.t4 B 1.27633f
C38 VP.n4 B 0.470766f
C39 VP.n5 B 0.491931f
C40 VP.n6 B 0.483851f
C41 VP.n7 B 0.010962f
C42 VP.n8 B 0.48117f
C43 VP.n9 B 2.23437f
C44 VP.n10 B 2.27293f
C45 VP.t6 B 1.26209f
C46 VP.n11 B 0.48117f
C47 VP.n12 B 0.010962f
C48 VP.n13 B 0.048309f
C49 VP.n14 B 0.048309f
C50 VP.n15 B 0.048309f
C51 VP.t5 B 1.26209f
C52 VP.n16 B 0.483851f
C53 VP.n17 B 0.010962f
C54 VP.t1 B 1.26209f
C55 VP.n18 B 0.48117f
C56 VP.n19 B 0.037438f
C57 VTAIL.t11 B 0.275143f
C58 VTAIL.t12 B 0.275143f
C59 VTAIL.n0 B 2.43178f
C60 VTAIL.n1 B 0.263632f
C61 VTAIL.t14 B 3.10375f
C62 VTAIL.n2 B 0.369144f
C63 VTAIL.t2 B 3.10375f
C64 VTAIL.n3 B 0.369144f
C65 VTAIL.t1 B 0.275143f
C66 VTAIL.t0 B 0.275143f
C67 VTAIL.n4 B 2.43178f
C68 VTAIL.n5 B 0.309154f
C69 VTAIL.t4 B 3.10375f
C70 VTAIL.n6 B 1.63215f
C71 VTAIL.t7 B 3.10377f
C72 VTAIL.n7 B 1.63212f
C73 VTAIL.t13 B 0.275143f
C74 VTAIL.t9 B 0.275143f
C75 VTAIL.n8 B 2.43178f
C76 VTAIL.n9 B 0.30915f
C77 VTAIL.t8 B 3.10377f
C78 VTAIL.n10 B 0.369123f
C79 VTAIL.t5 B 3.10377f
C80 VTAIL.n11 B 0.369123f
C81 VTAIL.t6 B 0.275143f
C82 VTAIL.t15 B 0.275143f
C83 VTAIL.n12 B 2.43178f
C84 VTAIL.n13 B 0.30915f
C85 VTAIL.t3 B 3.10374f
C86 VTAIL.n14 B 1.63215f
C87 VTAIL.t10 B 3.10375f
C88 VTAIL.n15 B 1.62832f
C89 VDD2.t3 B 0.389434f
C90 VDD2.t7 B 0.389434f
C91 VDD2.n0 B 3.53829f
C92 VDD2.t4 B 0.389434f
C93 VDD2.t6 B 0.389434f
C94 VDD2.n1 B 3.53829f
C95 VDD2.n2 B 2.77378f
C96 VDD2.t2 B 0.389434f
C97 VDD2.t5 B 0.389434f
C98 VDD2.n3 B 3.53636f
C99 VDD2.n4 B 3.03789f
C100 VDD2.t1 B 0.389434f
C101 VDD2.t0 B 0.389434f
C102 VDD2.n5 B 3.53825f
C103 VN.n0 B 0.047631f
C104 VN.t3 B 1.24436f
C105 VN.n1 B 0.485019f
C106 VN.t0 B 1.2584f
C107 VN.n2 B 0.464152f
C108 VN.n3 B 0.193985f
C109 VN.t2 B 1.24436f
C110 VN.n4 B 0.477053f
C111 VN.n5 B 0.010808f
C112 VN.t4 B 1.24436f
C113 VN.n6 B 0.47441f
C114 VN.n7 B 0.036912f
C115 VN.n8 B 0.047631f
C116 VN.t5 B 1.24436f
C117 VN.n9 B 0.485019f
C118 VN.t1 B 1.24436f
C119 VN.t6 B 1.2584f
C120 VN.n10 B 0.464152f
C121 VN.n11 B 0.193985f
C122 VN.n12 B 0.477053f
C123 VN.n13 B 0.010808f
C124 VN.t7 B 1.24436f
C125 VN.n14 B 0.47441f
C126 VN.n15 B 2.23412f
.ends

