* NGSPICE file created from diff_pair_sample_1353.ext - technology: sky130A

.subckt diff_pair_sample_1353 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t3 VP.t0 VTAIL.t4 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9931 pd=18.47 as=7.0746 ps=37.06 w=18.14 l=0.52
X1 VTAIL.t3 VN.t0 VDD2.t3 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=2.9931 ps=18.47 w=18.14 l=0.52
X2 VDD1.t2 VP.t1 VTAIL.t7 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9931 pd=18.47 as=7.0746 ps=37.06 w=18.14 l=0.52
X3 B.t17 B.t15 B.t16 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=0 ps=0 w=18.14 l=0.52
X4 B.t14 B.t12 B.t13 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=0 ps=0 w=18.14 l=0.52
X5 B.t11 B.t8 B.t10 B.t9 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=0 ps=0 w=18.14 l=0.52
X6 VDD2.t2 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=2.9931 pd=18.47 as=7.0746 ps=37.06 w=18.14 l=0.52
X7 B.t7 B.t4 B.t6 B.t5 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=0 ps=0 w=18.14 l=0.52
X8 VTAIL.t2 VN.t2 VDD2.t1 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=2.9931 ps=18.47 w=18.14 l=0.52
X9 VTAIL.t6 VP.t2 VDD1.t1 B.t3 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=2.9931 ps=18.47 w=18.14 l=0.52
X10 VDD2.t0 VN.t3 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=2.9931 pd=18.47 as=7.0746 ps=37.06 w=18.14 l=0.52
X11 VTAIL.t5 VP.t3 VDD1.t0 B.t2 sky130_fd_pr__nfet_01v8 ad=7.0746 pd=37.06 as=2.9931 ps=18.47 w=18.14 l=0.52
R0 VP.n0 VP.t2 937.245
R1 VP.n0 VP.t0 937.221
R2 VP.n2 VP.t3 916.264
R3 VP.n3 VP.t1 916.264
R4 VP.n4 VP.n3 161.3
R5 VP.n2 VP.n1 161.3
R6 VP.n1 VP.n0 114.782
R7 VP.n3 VP.n2 48.2005
R8 VP.n4 VP.n1 0.189894
R9 VP VP.n4 0.0516364
R10 VTAIL.n810 VTAIL.n714 289.615
R11 VTAIL.n96 VTAIL.n0 289.615
R12 VTAIL.n198 VTAIL.n102 289.615
R13 VTAIL.n300 VTAIL.n204 289.615
R14 VTAIL.n708 VTAIL.n612 289.615
R15 VTAIL.n606 VTAIL.n510 289.615
R16 VTAIL.n504 VTAIL.n408 289.615
R17 VTAIL.n402 VTAIL.n306 289.615
R18 VTAIL.n746 VTAIL.n745 185
R19 VTAIL.n751 VTAIL.n750 185
R20 VTAIL.n753 VTAIL.n752 185
R21 VTAIL.n742 VTAIL.n741 185
R22 VTAIL.n759 VTAIL.n758 185
R23 VTAIL.n761 VTAIL.n760 185
R24 VTAIL.n738 VTAIL.n737 185
R25 VTAIL.n767 VTAIL.n766 185
R26 VTAIL.n769 VTAIL.n768 185
R27 VTAIL.n734 VTAIL.n733 185
R28 VTAIL.n775 VTAIL.n774 185
R29 VTAIL.n777 VTAIL.n776 185
R30 VTAIL.n730 VTAIL.n729 185
R31 VTAIL.n783 VTAIL.n782 185
R32 VTAIL.n785 VTAIL.n784 185
R33 VTAIL.n726 VTAIL.n725 185
R34 VTAIL.n792 VTAIL.n791 185
R35 VTAIL.n793 VTAIL.n724 185
R36 VTAIL.n795 VTAIL.n794 185
R37 VTAIL.n722 VTAIL.n721 185
R38 VTAIL.n801 VTAIL.n800 185
R39 VTAIL.n803 VTAIL.n802 185
R40 VTAIL.n718 VTAIL.n717 185
R41 VTAIL.n809 VTAIL.n808 185
R42 VTAIL.n811 VTAIL.n810 185
R43 VTAIL.n32 VTAIL.n31 185
R44 VTAIL.n37 VTAIL.n36 185
R45 VTAIL.n39 VTAIL.n38 185
R46 VTAIL.n28 VTAIL.n27 185
R47 VTAIL.n45 VTAIL.n44 185
R48 VTAIL.n47 VTAIL.n46 185
R49 VTAIL.n24 VTAIL.n23 185
R50 VTAIL.n53 VTAIL.n52 185
R51 VTAIL.n55 VTAIL.n54 185
R52 VTAIL.n20 VTAIL.n19 185
R53 VTAIL.n61 VTAIL.n60 185
R54 VTAIL.n63 VTAIL.n62 185
R55 VTAIL.n16 VTAIL.n15 185
R56 VTAIL.n69 VTAIL.n68 185
R57 VTAIL.n71 VTAIL.n70 185
R58 VTAIL.n12 VTAIL.n11 185
R59 VTAIL.n78 VTAIL.n77 185
R60 VTAIL.n79 VTAIL.n10 185
R61 VTAIL.n81 VTAIL.n80 185
R62 VTAIL.n8 VTAIL.n7 185
R63 VTAIL.n87 VTAIL.n86 185
R64 VTAIL.n89 VTAIL.n88 185
R65 VTAIL.n4 VTAIL.n3 185
R66 VTAIL.n95 VTAIL.n94 185
R67 VTAIL.n97 VTAIL.n96 185
R68 VTAIL.n134 VTAIL.n133 185
R69 VTAIL.n139 VTAIL.n138 185
R70 VTAIL.n141 VTAIL.n140 185
R71 VTAIL.n130 VTAIL.n129 185
R72 VTAIL.n147 VTAIL.n146 185
R73 VTAIL.n149 VTAIL.n148 185
R74 VTAIL.n126 VTAIL.n125 185
R75 VTAIL.n155 VTAIL.n154 185
R76 VTAIL.n157 VTAIL.n156 185
R77 VTAIL.n122 VTAIL.n121 185
R78 VTAIL.n163 VTAIL.n162 185
R79 VTAIL.n165 VTAIL.n164 185
R80 VTAIL.n118 VTAIL.n117 185
R81 VTAIL.n171 VTAIL.n170 185
R82 VTAIL.n173 VTAIL.n172 185
R83 VTAIL.n114 VTAIL.n113 185
R84 VTAIL.n180 VTAIL.n179 185
R85 VTAIL.n181 VTAIL.n112 185
R86 VTAIL.n183 VTAIL.n182 185
R87 VTAIL.n110 VTAIL.n109 185
R88 VTAIL.n189 VTAIL.n188 185
R89 VTAIL.n191 VTAIL.n190 185
R90 VTAIL.n106 VTAIL.n105 185
R91 VTAIL.n197 VTAIL.n196 185
R92 VTAIL.n199 VTAIL.n198 185
R93 VTAIL.n236 VTAIL.n235 185
R94 VTAIL.n241 VTAIL.n240 185
R95 VTAIL.n243 VTAIL.n242 185
R96 VTAIL.n232 VTAIL.n231 185
R97 VTAIL.n249 VTAIL.n248 185
R98 VTAIL.n251 VTAIL.n250 185
R99 VTAIL.n228 VTAIL.n227 185
R100 VTAIL.n257 VTAIL.n256 185
R101 VTAIL.n259 VTAIL.n258 185
R102 VTAIL.n224 VTAIL.n223 185
R103 VTAIL.n265 VTAIL.n264 185
R104 VTAIL.n267 VTAIL.n266 185
R105 VTAIL.n220 VTAIL.n219 185
R106 VTAIL.n273 VTAIL.n272 185
R107 VTAIL.n275 VTAIL.n274 185
R108 VTAIL.n216 VTAIL.n215 185
R109 VTAIL.n282 VTAIL.n281 185
R110 VTAIL.n283 VTAIL.n214 185
R111 VTAIL.n285 VTAIL.n284 185
R112 VTAIL.n212 VTAIL.n211 185
R113 VTAIL.n291 VTAIL.n290 185
R114 VTAIL.n293 VTAIL.n292 185
R115 VTAIL.n208 VTAIL.n207 185
R116 VTAIL.n299 VTAIL.n298 185
R117 VTAIL.n301 VTAIL.n300 185
R118 VTAIL.n709 VTAIL.n708 185
R119 VTAIL.n707 VTAIL.n706 185
R120 VTAIL.n616 VTAIL.n615 185
R121 VTAIL.n701 VTAIL.n700 185
R122 VTAIL.n699 VTAIL.n698 185
R123 VTAIL.n620 VTAIL.n619 185
R124 VTAIL.n693 VTAIL.n692 185
R125 VTAIL.n691 VTAIL.n622 185
R126 VTAIL.n690 VTAIL.n689 185
R127 VTAIL.n625 VTAIL.n623 185
R128 VTAIL.n684 VTAIL.n683 185
R129 VTAIL.n682 VTAIL.n681 185
R130 VTAIL.n629 VTAIL.n628 185
R131 VTAIL.n676 VTAIL.n675 185
R132 VTAIL.n674 VTAIL.n673 185
R133 VTAIL.n633 VTAIL.n632 185
R134 VTAIL.n668 VTAIL.n667 185
R135 VTAIL.n666 VTAIL.n665 185
R136 VTAIL.n637 VTAIL.n636 185
R137 VTAIL.n660 VTAIL.n659 185
R138 VTAIL.n658 VTAIL.n657 185
R139 VTAIL.n641 VTAIL.n640 185
R140 VTAIL.n652 VTAIL.n651 185
R141 VTAIL.n650 VTAIL.n649 185
R142 VTAIL.n645 VTAIL.n644 185
R143 VTAIL.n607 VTAIL.n606 185
R144 VTAIL.n605 VTAIL.n604 185
R145 VTAIL.n514 VTAIL.n513 185
R146 VTAIL.n599 VTAIL.n598 185
R147 VTAIL.n597 VTAIL.n596 185
R148 VTAIL.n518 VTAIL.n517 185
R149 VTAIL.n591 VTAIL.n590 185
R150 VTAIL.n589 VTAIL.n520 185
R151 VTAIL.n588 VTAIL.n587 185
R152 VTAIL.n523 VTAIL.n521 185
R153 VTAIL.n582 VTAIL.n581 185
R154 VTAIL.n580 VTAIL.n579 185
R155 VTAIL.n527 VTAIL.n526 185
R156 VTAIL.n574 VTAIL.n573 185
R157 VTAIL.n572 VTAIL.n571 185
R158 VTAIL.n531 VTAIL.n530 185
R159 VTAIL.n566 VTAIL.n565 185
R160 VTAIL.n564 VTAIL.n563 185
R161 VTAIL.n535 VTAIL.n534 185
R162 VTAIL.n558 VTAIL.n557 185
R163 VTAIL.n556 VTAIL.n555 185
R164 VTAIL.n539 VTAIL.n538 185
R165 VTAIL.n550 VTAIL.n549 185
R166 VTAIL.n548 VTAIL.n547 185
R167 VTAIL.n543 VTAIL.n542 185
R168 VTAIL.n505 VTAIL.n504 185
R169 VTAIL.n503 VTAIL.n502 185
R170 VTAIL.n412 VTAIL.n411 185
R171 VTAIL.n497 VTAIL.n496 185
R172 VTAIL.n495 VTAIL.n494 185
R173 VTAIL.n416 VTAIL.n415 185
R174 VTAIL.n489 VTAIL.n488 185
R175 VTAIL.n487 VTAIL.n418 185
R176 VTAIL.n486 VTAIL.n485 185
R177 VTAIL.n421 VTAIL.n419 185
R178 VTAIL.n480 VTAIL.n479 185
R179 VTAIL.n478 VTAIL.n477 185
R180 VTAIL.n425 VTAIL.n424 185
R181 VTAIL.n472 VTAIL.n471 185
R182 VTAIL.n470 VTAIL.n469 185
R183 VTAIL.n429 VTAIL.n428 185
R184 VTAIL.n464 VTAIL.n463 185
R185 VTAIL.n462 VTAIL.n461 185
R186 VTAIL.n433 VTAIL.n432 185
R187 VTAIL.n456 VTAIL.n455 185
R188 VTAIL.n454 VTAIL.n453 185
R189 VTAIL.n437 VTAIL.n436 185
R190 VTAIL.n448 VTAIL.n447 185
R191 VTAIL.n446 VTAIL.n445 185
R192 VTAIL.n441 VTAIL.n440 185
R193 VTAIL.n403 VTAIL.n402 185
R194 VTAIL.n401 VTAIL.n400 185
R195 VTAIL.n310 VTAIL.n309 185
R196 VTAIL.n395 VTAIL.n394 185
R197 VTAIL.n393 VTAIL.n392 185
R198 VTAIL.n314 VTAIL.n313 185
R199 VTAIL.n387 VTAIL.n386 185
R200 VTAIL.n385 VTAIL.n316 185
R201 VTAIL.n384 VTAIL.n383 185
R202 VTAIL.n319 VTAIL.n317 185
R203 VTAIL.n378 VTAIL.n377 185
R204 VTAIL.n376 VTAIL.n375 185
R205 VTAIL.n323 VTAIL.n322 185
R206 VTAIL.n370 VTAIL.n369 185
R207 VTAIL.n368 VTAIL.n367 185
R208 VTAIL.n327 VTAIL.n326 185
R209 VTAIL.n362 VTAIL.n361 185
R210 VTAIL.n360 VTAIL.n359 185
R211 VTAIL.n331 VTAIL.n330 185
R212 VTAIL.n354 VTAIL.n353 185
R213 VTAIL.n352 VTAIL.n351 185
R214 VTAIL.n335 VTAIL.n334 185
R215 VTAIL.n346 VTAIL.n345 185
R216 VTAIL.n344 VTAIL.n343 185
R217 VTAIL.n339 VTAIL.n338 185
R218 VTAIL.n747 VTAIL.t1 147.659
R219 VTAIL.n33 VTAIL.t3 147.659
R220 VTAIL.n135 VTAIL.t7 147.659
R221 VTAIL.n237 VTAIL.t5 147.659
R222 VTAIL.n646 VTAIL.t4 147.659
R223 VTAIL.n544 VTAIL.t6 147.659
R224 VTAIL.n442 VTAIL.t0 147.659
R225 VTAIL.n340 VTAIL.t2 147.659
R226 VTAIL.n751 VTAIL.n745 104.615
R227 VTAIL.n752 VTAIL.n751 104.615
R228 VTAIL.n752 VTAIL.n741 104.615
R229 VTAIL.n759 VTAIL.n741 104.615
R230 VTAIL.n760 VTAIL.n759 104.615
R231 VTAIL.n760 VTAIL.n737 104.615
R232 VTAIL.n767 VTAIL.n737 104.615
R233 VTAIL.n768 VTAIL.n767 104.615
R234 VTAIL.n768 VTAIL.n733 104.615
R235 VTAIL.n775 VTAIL.n733 104.615
R236 VTAIL.n776 VTAIL.n775 104.615
R237 VTAIL.n776 VTAIL.n729 104.615
R238 VTAIL.n783 VTAIL.n729 104.615
R239 VTAIL.n784 VTAIL.n783 104.615
R240 VTAIL.n784 VTAIL.n725 104.615
R241 VTAIL.n792 VTAIL.n725 104.615
R242 VTAIL.n793 VTAIL.n792 104.615
R243 VTAIL.n794 VTAIL.n793 104.615
R244 VTAIL.n794 VTAIL.n721 104.615
R245 VTAIL.n801 VTAIL.n721 104.615
R246 VTAIL.n802 VTAIL.n801 104.615
R247 VTAIL.n802 VTAIL.n717 104.615
R248 VTAIL.n809 VTAIL.n717 104.615
R249 VTAIL.n810 VTAIL.n809 104.615
R250 VTAIL.n37 VTAIL.n31 104.615
R251 VTAIL.n38 VTAIL.n37 104.615
R252 VTAIL.n38 VTAIL.n27 104.615
R253 VTAIL.n45 VTAIL.n27 104.615
R254 VTAIL.n46 VTAIL.n45 104.615
R255 VTAIL.n46 VTAIL.n23 104.615
R256 VTAIL.n53 VTAIL.n23 104.615
R257 VTAIL.n54 VTAIL.n53 104.615
R258 VTAIL.n54 VTAIL.n19 104.615
R259 VTAIL.n61 VTAIL.n19 104.615
R260 VTAIL.n62 VTAIL.n61 104.615
R261 VTAIL.n62 VTAIL.n15 104.615
R262 VTAIL.n69 VTAIL.n15 104.615
R263 VTAIL.n70 VTAIL.n69 104.615
R264 VTAIL.n70 VTAIL.n11 104.615
R265 VTAIL.n78 VTAIL.n11 104.615
R266 VTAIL.n79 VTAIL.n78 104.615
R267 VTAIL.n80 VTAIL.n79 104.615
R268 VTAIL.n80 VTAIL.n7 104.615
R269 VTAIL.n87 VTAIL.n7 104.615
R270 VTAIL.n88 VTAIL.n87 104.615
R271 VTAIL.n88 VTAIL.n3 104.615
R272 VTAIL.n95 VTAIL.n3 104.615
R273 VTAIL.n96 VTAIL.n95 104.615
R274 VTAIL.n139 VTAIL.n133 104.615
R275 VTAIL.n140 VTAIL.n139 104.615
R276 VTAIL.n140 VTAIL.n129 104.615
R277 VTAIL.n147 VTAIL.n129 104.615
R278 VTAIL.n148 VTAIL.n147 104.615
R279 VTAIL.n148 VTAIL.n125 104.615
R280 VTAIL.n155 VTAIL.n125 104.615
R281 VTAIL.n156 VTAIL.n155 104.615
R282 VTAIL.n156 VTAIL.n121 104.615
R283 VTAIL.n163 VTAIL.n121 104.615
R284 VTAIL.n164 VTAIL.n163 104.615
R285 VTAIL.n164 VTAIL.n117 104.615
R286 VTAIL.n171 VTAIL.n117 104.615
R287 VTAIL.n172 VTAIL.n171 104.615
R288 VTAIL.n172 VTAIL.n113 104.615
R289 VTAIL.n180 VTAIL.n113 104.615
R290 VTAIL.n181 VTAIL.n180 104.615
R291 VTAIL.n182 VTAIL.n181 104.615
R292 VTAIL.n182 VTAIL.n109 104.615
R293 VTAIL.n189 VTAIL.n109 104.615
R294 VTAIL.n190 VTAIL.n189 104.615
R295 VTAIL.n190 VTAIL.n105 104.615
R296 VTAIL.n197 VTAIL.n105 104.615
R297 VTAIL.n198 VTAIL.n197 104.615
R298 VTAIL.n241 VTAIL.n235 104.615
R299 VTAIL.n242 VTAIL.n241 104.615
R300 VTAIL.n242 VTAIL.n231 104.615
R301 VTAIL.n249 VTAIL.n231 104.615
R302 VTAIL.n250 VTAIL.n249 104.615
R303 VTAIL.n250 VTAIL.n227 104.615
R304 VTAIL.n257 VTAIL.n227 104.615
R305 VTAIL.n258 VTAIL.n257 104.615
R306 VTAIL.n258 VTAIL.n223 104.615
R307 VTAIL.n265 VTAIL.n223 104.615
R308 VTAIL.n266 VTAIL.n265 104.615
R309 VTAIL.n266 VTAIL.n219 104.615
R310 VTAIL.n273 VTAIL.n219 104.615
R311 VTAIL.n274 VTAIL.n273 104.615
R312 VTAIL.n274 VTAIL.n215 104.615
R313 VTAIL.n282 VTAIL.n215 104.615
R314 VTAIL.n283 VTAIL.n282 104.615
R315 VTAIL.n284 VTAIL.n283 104.615
R316 VTAIL.n284 VTAIL.n211 104.615
R317 VTAIL.n291 VTAIL.n211 104.615
R318 VTAIL.n292 VTAIL.n291 104.615
R319 VTAIL.n292 VTAIL.n207 104.615
R320 VTAIL.n299 VTAIL.n207 104.615
R321 VTAIL.n300 VTAIL.n299 104.615
R322 VTAIL.n708 VTAIL.n707 104.615
R323 VTAIL.n707 VTAIL.n615 104.615
R324 VTAIL.n700 VTAIL.n615 104.615
R325 VTAIL.n700 VTAIL.n699 104.615
R326 VTAIL.n699 VTAIL.n619 104.615
R327 VTAIL.n692 VTAIL.n619 104.615
R328 VTAIL.n692 VTAIL.n691 104.615
R329 VTAIL.n691 VTAIL.n690 104.615
R330 VTAIL.n690 VTAIL.n623 104.615
R331 VTAIL.n683 VTAIL.n623 104.615
R332 VTAIL.n683 VTAIL.n682 104.615
R333 VTAIL.n682 VTAIL.n628 104.615
R334 VTAIL.n675 VTAIL.n628 104.615
R335 VTAIL.n675 VTAIL.n674 104.615
R336 VTAIL.n674 VTAIL.n632 104.615
R337 VTAIL.n667 VTAIL.n632 104.615
R338 VTAIL.n667 VTAIL.n666 104.615
R339 VTAIL.n666 VTAIL.n636 104.615
R340 VTAIL.n659 VTAIL.n636 104.615
R341 VTAIL.n659 VTAIL.n658 104.615
R342 VTAIL.n658 VTAIL.n640 104.615
R343 VTAIL.n651 VTAIL.n640 104.615
R344 VTAIL.n651 VTAIL.n650 104.615
R345 VTAIL.n650 VTAIL.n644 104.615
R346 VTAIL.n606 VTAIL.n605 104.615
R347 VTAIL.n605 VTAIL.n513 104.615
R348 VTAIL.n598 VTAIL.n513 104.615
R349 VTAIL.n598 VTAIL.n597 104.615
R350 VTAIL.n597 VTAIL.n517 104.615
R351 VTAIL.n590 VTAIL.n517 104.615
R352 VTAIL.n590 VTAIL.n589 104.615
R353 VTAIL.n589 VTAIL.n588 104.615
R354 VTAIL.n588 VTAIL.n521 104.615
R355 VTAIL.n581 VTAIL.n521 104.615
R356 VTAIL.n581 VTAIL.n580 104.615
R357 VTAIL.n580 VTAIL.n526 104.615
R358 VTAIL.n573 VTAIL.n526 104.615
R359 VTAIL.n573 VTAIL.n572 104.615
R360 VTAIL.n572 VTAIL.n530 104.615
R361 VTAIL.n565 VTAIL.n530 104.615
R362 VTAIL.n565 VTAIL.n564 104.615
R363 VTAIL.n564 VTAIL.n534 104.615
R364 VTAIL.n557 VTAIL.n534 104.615
R365 VTAIL.n557 VTAIL.n556 104.615
R366 VTAIL.n556 VTAIL.n538 104.615
R367 VTAIL.n549 VTAIL.n538 104.615
R368 VTAIL.n549 VTAIL.n548 104.615
R369 VTAIL.n548 VTAIL.n542 104.615
R370 VTAIL.n504 VTAIL.n503 104.615
R371 VTAIL.n503 VTAIL.n411 104.615
R372 VTAIL.n496 VTAIL.n411 104.615
R373 VTAIL.n496 VTAIL.n495 104.615
R374 VTAIL.n495 VTAIL.n415 104.615
R375 VTAIL.n488 VTAIL.n415 104.615
R376 VTAIL.n488 VTAIL.n487 104.615
R377 VTAIL.n487 VTAIL.n486 104.615
R378 VTAIL.n486 VTAIL.n419 104.615
R379 VTAIL.n479 VTAIL.n419 104.615
R380 VTAIL.n479 VTAIL.n478 104.615
R381 VTAIL.n478 VTAIL.n424 104.615
R382 VTAIL.n471 VTAIL.n424 104.615
R383 VTAIL.n471 VTAIL.n470 104.615
R384 VTAIL.n470 VTAIL.n428 104.615
R385 VTAIL.n463 VTAIL.n428 104.615
R386 VTAIL.n463 VTAIL.n462 104.615
R387 VTAIL.n462 VTAIL.n432 104.615
R388 VTAIL.n455 VTAIL.n432 104.615
R389 VTAIL.n455 VTAIL.n454 104.615
R390 VTAIL.n454 VTAIL.n436 104.615
R391 VTAIL.n447 VTAIL.n436 104.615
R392 VTAIL.n447 VTAIL.n446 104.615
R393 VTAIL.n446 VTAIL.n440 104.615
R394 VTAIL.n402 VTAIL.n401 104.615
R395 VTAIL.n401 VTAIL.n309 104.615
R396 VTAIL.n394 VTAIL.n309 104.615
R397 VTAIL.n394 VTAIL.n393 104.615
R398 VTAIL.n393 VTAIL.n313 104.615
R399 VTAIL.n386 VTAIL.n313 104.615
R400 VTAIL.n386 VTAIL.n385 104.615
R401 VTAIL.n385 VTAIL.n384 104.615
R402 VTAIL.n384 VTAIL.n317 104.615
R403 VTAIL.n377 VTAIL.n317 104.615
R404 VTAIL.n377 VTAIL.n376 104.615
R405 VTAIL.n376 VTAIL.n322 104.615
R406 VTAIL.n369 VTAIL.n322 104.615
R407 VTAIL.n369 VTAIL.n368 104.615
R408 VTAIL.n368 VTAIL.n326 104.615
R409 VTAIL.n361 VTAIL.n326 104.615
R410 VTAIL.n361 VTAIL.n360 104.615
R411 VTAIL.n360 VTAIL.n330 104.615
R412 VTAIL.n353 VTAIL.n330 104.615
R413 VTAIL.n353 VTAIL.n352 104.615
R414 VTAIL.n352 VTAIL.n334 104.615
R415 VTAIL.n345 VTAIL.n334 104.615
R416 VTAIL.n345 VTAIL.n344 104.615
R417 VTAIL.n344 VTAIL.n338 104.615
R418 VTAIL.t1 VTAIL.n745 52.3082
R419 VTAIL.t3 VTAIL.n31 52.3082
R420 VTAIL.t7 VTAIL.n133 52.3082
R421 VTAIL.t5 VTAIL.n235 52.3082
R422 VTAIL.t4 VTAIL.n644 52.3082
R423 VTAIL.t6 VTAIL.n542 52.3082
R424 VTAIL.t0 VTAIL.n440 52.3082
R425 VTAIL.t2 VTAIL.n338 52.3082
R426 VTAIL.n815 VTAIL.n814 30.246
R427 VTAIL.n101 VTAIL.n100 30.246
R428 VTAIL.n203 VTAIL.n202 30.246
R429 VTAIL.n305 VTAIL.n304 30.246
R430 VTAIL.n713 VTAIL.n712 30.246
R431 VTAIL.n611 VTAIL.n610 30.246
R432 VTAIL.n509 VTAIL.n508 30.246
R433 VTAIL.n407 VTAIL.n406 30.246
R434 VTAIL.n815 VTAIL.n713 28.7376
R435 VTAIL.n407 VTAIL.n305 28.7376
R436 VTAIL.n747 VTAIL.n746 15.6677
R437 VTAIL.n33 VTAIL.n32 15.6677
R438 VTAIL.n135 VTAIL.n134 15.6677
R439 VTAIL.n237 VTAIL.n236 15.6677
R440 VTAIL.n646 VTAIL.n645 15.6677
R441 VTAIL.n544 VTAIL.n543 15.6677
R442 VTAIL.n442 VTAIL.n441 15.6677
R443 VTAIL.n340 VTAIL.n339 15.6677
R444 VTAIL.n795 VTAIL.n724 13.1884
R445 VTAIL.n81 VTAIL.n10 13.1884
R446 VTAIL.n183 VTAIL.n112 13.1884
R447 VTAIL.n285 VTAIL.n214 13.1884
R448 VTAIL.n693 VTAIL.n622 13.1884
R449 VTAIL.n591 VTAIL.n520 13.1884
R450 VTAIL.n489 VTAIL.n418 13.1884
R451 VTAIL.n387 VTAIL.n316 13.1884
R452 VTAIL.n750 VTAIL.n749 12.8005
R453 VTAIL.n791 VTAIL.n790 12.8005
R454 VTAIL.n796 VTAIL.n722 12.8005
R455 VTAIL.n36 VTAIL.n35 12.8005
R456 VTAIL.n77 VTAIL.n76 12.8005
R457 VTAIL.n82 VTAIL.n8 12.8005
R458 VTAIL.n138 VTAIL.n137 12.8005
R459 VTAIL.n179 VTAIL.n178 12.8005
R460 VTAIL.n184 VTAIL.n110 12.8005
R461 VTAIL.n240 VTAIL.n239 12.8005
R462 VTAIL.n281 VTAIL.n280 12.8005
R463 VTAIL.n286 VTAIL.n212 12.8005
R464 VTAIL.n694 VTAIL.n620 12.8005
R465 VTAIL.n689 VTAIL.n624 12.8005
R466 VTAIL.n649 VTAIL.n648 12.8005
R467 VTAIL.n592 VTAIL.n518 12.8005
R468 VTAIL.n587 VTAIL.n522 12.8005
R469 VTAIL.n547 VTAIL.n546 12.8005
R470 VTAIL.n490 VTAIL.n416 12.8005
R471 VTAIL.n485 VTAIL.n420 12.8005
R472 VTAIL.n445 VTAIL.n444 12.8005
R473 VTAIL.n388 VTAIL.n314 12.8005
R474 VTAIL.n383 VTAIL.n318 12.8005
R475 VTAIL.n343 VTAIL.n342 12.8005
R476 VTAIL.n753 VTAIL.n744 12.0247
R477 VTAIL.n789 VTAIL.n726 12.0247
R478 VTAIL.n800 VTAIL.n799 12.0247
R479 VTAIL.n39 VTAIL.n30 12.0247
R480 VTAIL.n75 VTAIL.n12 12.0247
R481 VTAIL.n86 VTAIL.n85 12.0247
R482 VTAIL.n141 VTAIL.n132 12.0247
R483 VTAIL.n177 VTAIL.n114 12.0247
R484 VTAIL.n188 VTAIL.n187 12.0247
R485 VTAIL.n243 VTAIL.n234 12.0247
R486 VTAIL.n279 VTAIL.n216 12.0247
R487 VTAIL.n290 VTAIL.n289 12.0247
R488 VTAIL.n698 VTAIL.n697 12.0247
R489 VTAIL.n688 VTAIL.n625 12.0247
R490 VTAIL.n652 VTAIL.n643 12.0247
R491 VTAIL.n596 VTAIL.n595 12.0247
R492 VTAIL.n586 VTAIL.n523 12.0247
R493 VTAIL.n550 VTAIL.n541 12.0247
R494 VTAIL.n494 VTAIL.n493 12.0247
R495 VTAIL.n484 VTAIL.n421 12.0247
R496 VTAIL.n448 VTAIL.n439 12.0247
R497 VTAIL.n392 VTAIL.n391 12.0247
R498 VTAIL.n382 VTAIL.n319 12.0247
R499 VTAIL.n346 VTAIL.n337 12.0247
R500 VTAIL.n754 VTAIL.n742 11.249
R501 VTAIL.n786 VTAIL.n785 11.249
R502 VTAIL.n803 VTAIL.n720 11.249
R503 VTAIL.n40 VTAIL.n28 11.249
R504 VTAIL.n72 VTAIL.n71 11.249
R505 VTAIL.n89 VTAIL.n6 11.249
R506 VTAIL.n142 VTAIL.n130 11.249
R507 VTAIL.n174 VTAIL.n173 11.249
R508 VTAIL.n191 VTAIL.n108 11.249
R509 VTAIL.n244 VTAIL.n232 11.249
R510 VTAIL.n276 VTAIL.n275 11.249
R511 VTAIL.n293 VTAIL.n210 11.249
R512 VTAIL.n701 VTAIL.n618 11.249
R513 VTAIL.n685 VTAIL.n684 11.249
R514 VTAIL.n653 VTAIL.n641 11.249
R515 VTAIL.n599 VTAIL.n516 11.249
R516 VTAIL.n583 VTAIL.n582 11.249
R517 VTAIL.n551 VTAIL.n539 11.249
R518 VTAIL.n497 VTAIL.n414 11.249
R519 VTAIL.n481 VTAIL.n480 11.249
R520 VTAIL.n449 VTAIL.n437 11.249
R521 VTAIL.n395 VTAIL.n312 11.249
R522 VTAIL.n379 VTAIL.n378 11.249
R523 VTAIL.n347 VTAIL.n335 11.249
R524 VTAIL.n758 VTAIL.n757 10.4732
R525 VTAIL.n782 VTAIL.n728 10.4732
R526 VTAIL.n804 VTAIL.n718 10.4732
R527 VTAIL.n44 VTAIL.n43 10.4732
R528 VTAIL.n68 VTAIL.n14 10.4732
R529 VTAIL.n90 VTAIL.n4 10.4732
R530 VTAIL.n146 VTAIL.n145 10.4732
R531 VTAIL.n170 VTAIL.n116 10.4732
R532 VTAIL.n192 VTAIL.n106 10.4732
R533 VTAIL.n248 VTAIL.n247 10.4732
R534 VTAIL.n272 VTAIL.n218 10.4732
R535 VTAIL.n294 VTAIL.n208 10.4732
R536 VTAIL.n702 VTAIL.n616 10.4732
R537 VTAIL.n681 VTAIL.n627 10.4732
R538 VTAIL.n657 VTAIL.n656 10.4732
R539 VTAIL.n600 VTAIL.n514 10.4732
R540 VTAIL.n579 VTAIL.n525 10.4732
R541 VTAIL.n555 VTAIL.n554 10.4732
R542 VTAIL.n498 VTAIL.n412 10.4732
R543 VTAIL.n477 VTAIL.n423 10.4732
R544 VTAIL.n453 VTAIL.n452 10.4732
R545 VTAIL.n396 VTAIL.n310 10.4732
R546 VTAIL.n375 VTAIL.n321 10.4732
R547 VTAIL.n351 VTAIL.n350 10.4732
R548 VTAIL.n761 VTAIL.n740 9.69747
R549 VTAIL.n781 VTAIL.n730 9.69747
R550 VTAIL.n808 VTAIL.n807 9.69747
R551 VTAIL.n47 VTAIL.n26 9.69747
R552 VTAIL.n67 VTAIL.n16 9.69747
R553 VTAIL.n94 VTAIL.n93 9.69747
R554 VTAIL.n149 VTAIL.n128 9.69747
R555 VTAIL.n169 VTAIL.n118 9.69747
R556 VTAIL.n196 VTAIL.n195 9.69747
R557 VTAIL.n251 VTAIL.n230 9.69747
R558 VTAIL.n271 VTAIL.n220 9.69747
R559 VTAIL.n298 VTAIL.n297 9.69747
R560 VTAIL.n706 VTAIL.n705 9.69747
R561 VTAIL.n680 VTAIL.n629 9.69747
R562 VTAIL.n660 VTAIL.n639 9.69747
R563 VTAIL.n604 VTAIL.n603 9.69747
R564 VTAIL.n578 VTAIL.n527 9.69747
R565 VTAIL.n558 VTAIL.n537 9.69747
R566 VTAIL.n502 VTAIL.n501 9.69747
R567 VTAIL.n476 VTAIL.n425 9.69747
R568 VTAIL.n456 VTAIL.n435 9.69747
R569 VTAIL.n400 VTAIL.n399 9.69747
R570 VTAIL.n374 VTAIL.n323 9.69747
R571 VTAIL.n354 VTAIL.n333 9.69747
R572 VTAIL.n814 VTAIL.n813 9.45567
R573 VTAIL.n100 VTAIL.n99 9.45567
R574 VTAIL.n202 VTAIL.n201 9.45567
R575 VTAIL.n304 VTAIL.n303 9.45567
R576 VTAIL.n712 VTAIL.n711 9.45567
R577 VTAIL.n610 VTAIL.n609 9.45567
R578 VTAIL.n508 VTAIL.n507 9.45567
R579 VTAIL.n406 VTAIL.n405 9.45567
R580 VTAIL.n813 VTAIL.n812 9.3005
R581 VTAIL.n716 VTAIL.n715 9.3005
R582 VTAIL.n807 VTAIL.n806 9.3005
R583 VTAIL.n805 VTAIL.n804 9.3005
R584 VTAIL.n720 VTAIL.n719 9.3005
R585 VTAIL.n799 VTAIL.n798 9.3005
R586 VTAIL.n797 VTAIL.n796 9.3005
R587 VTAIL.n736 VTAIL.n735 9.3005
R588 VTAIL.n765 VTAIL.n764 9.3005
R589 VTAIL.n763 VTAIL.n762 9.3005
R590 VTAIL.n740 VTAIL.n739 9.3005
R591 VTAIL.n757 VTAIL.n756 9.3005
R592 VTAIL.n755 VTAIL.n754 9.3005
R593 VTAIL.n744 VTAIL.n743 9.3005
R594 VTAIL.n749 VTAIL.n748 9.3005
R595 VTAIL.n771 VTAIL.n770 9.3005
R596 VTAIL.n773 VTAIL.n772 9.3005
R597 VTAIL.n732 VTAIL.n731 9.3005
R598 VTAIL.n779 VTAIL.n778 9.3005
R599 VTAIL.n781 VTAIL.n780 9.3005
R600 VTAIL.n728 VTAIL.n727 9.3005
R601 VTAIL.n787 VTAIL.n786 9.3005
R602 VTAIL.n789 VTAIL.n788 9.3005
R603 VTAIL.n790 VTAIL.n723 9.3005
R604 VTAIL.n99 VTAIL.n98 9.3005
R605 VTAIL.n2 VTAIL.n1 9.3005
R606 VTAIL.n93 VTAIL.n92 9.3005
R607 VTAIL.n91 VTAIL.n90 9.3005
R608 VTAIL.n6 VTAIL.n5 9.3005
R609 VTAIL.n85 VTAIL.n84 9.3005
R610 VTAIL.n83 VTAIL.n82 9.3005
R611 VTAIL.n22 VTAIL.n21 9.3005
R612 VTAIL.n51 VTAIL.n50 9.3005
R613 VTAIL.n49 VTAIL.n48 9.3005
R614 VTAIL.n26 VTAIL.n25 9.3005
R615 VTAIL.n43 VTAIL.n42 9.3005
R616 VTAIL.n41 VTAIL.n40 9.3005
R617 VTAIL.n30 VTAIL.n29 9.3005
R618 VTAIL.n35 VTAIL.n34 9.3005
R619 VTAIL.n57 VTAIL.n56 9.3005
R620 VTAIL.n59 VTAIL.n58 9.3005
R621 VTAIL.n18 VTAIL.n17 9.3005
R622 VTAIL.n65 VTAIL.n64 9.3005
R623 VTAIL.n67 VTAIL.n66 9.3005
R624 VTAIL.n14 VTAIL.n13 9.3005
R625 VTAIL.n73 VTAIL.n72 9.3005
R626 VTAIL.n75 VTAIL.n74 9.3005
R627 VTAIL.n76 VTAIL.n9 9.3005
R628 VTAIL.n201 VTAIL.n200 9.3005
R629 VTAIL.n104 VTAIL.n103 9.3005
R630 VTAIL.n195 VTAIL.n194 9.3005
R631 VTAIL.n193 VTAIL.n192 9.3005
R632 VTAIL.n108 VTAIL.n107 9.3005
R633 VTAIL.n187 VTAIL.n186 9.3005
R634 VTAIL.n185 VTAIL.n184 9.3005
R635 VTAIL.n124 VTAIL.n123 9.3005
R636 VTAIL.n153 VTAIL.n152 9.3005
R637 VTAIL.n151 VTAIL.n150 9.3005
R638 VTAIL.n128 VTAIL.n127 9.3005
R639 VTAIL.n145 VTAIL.n144 9.3005
R640 VTAIL.n143 VTAIL.n142 9.3005
R641 VTAIL.n132 VTAIL.n131 9.3005
R642 VTAIL.n137 VTAIL.n136 9.3005
R643 VTAIL.n159 VTAIL.n158 9.3005
R644 VTAIL.n161 VTAIL.n160 9.3005
R645 VTAIL.n120 VTAIL.n119 9.3005
R646 VTAIL.n167 VTAIL.n166 9.3005
R647 VTAIL.n169 VTAIL.n168 9.3005
R648 VTAIL.n116 VTAIL.n115 9.3005
R649 VTAIL.n175 VTAIL.n174 9.3005
R650 VTAIL.n177 VTAIL.n176 9.3005
R651 VTAIL.n178 VTAIL.n111 9.3005
R652 VTAIL.n303 VTAIL.n302 9.3005
R653 VTAIL.n206 VTAIL.n205 9.3005
R654 VTAIL.n297 VTAIL.n296 9.3005
R655 VTAIL.n295 VTAIL.n294 9.3005
R656 VTAIL.n210 VTAIL.n209 9.3005
R657 VTAIL.n289 VTAIL.n288 9.3005
R658 VTAIL.n287 VTAIL.n286 9.3005
R659 VTAIL.n226 VTAIL.n225 9.3005
R660 VTAIL.n255 VTAIL.n254 9.3005
R661 VTAIL.n253 VTAIL.n252 9.3005
R662 VTAIL.n230 VTAIL.n229 9.3005
R663 VTAIL.n247 VTAIL.n246 9.3005
R664 VTAIL.n245 VTAIL.n244 9.3005
R665 VTAIL.n234 VTAIL.n233 9.3005
R666 VTAIL.n239 VTAIL.n238 9.3005
R667 VTAIL.n261 VTAIL.n260 9.3005
R668 VTAIL.n263 VTAIL.n262 9.3005
R669 VTAIL.n222 VTAIL.n221 9.3005
R670 VTAIL.n269 VTAIL.n268 9.3005
R671 VTAIL.n271 VTAIL.n270 9.3005
R672 VTAIL.n218 VTAIL.n217 9.3005
R673 VTAIL.n277 VTAIL.n276 9.3005
R674 VTAIL.n279 VTAIL.n278 9.3005
R675 VTAIL.n280 VTAIL.n213 9.3005
R676 VTAIL.n672 VTAIL.n671 9.3005
R677 VTAIL.n631 VTAIL.n630 9.3005
R678 VTAIL.n678 VTAIL.n677 9.3005
R679 VTAIL.n680 VTAIL.n679 9.3005
R680 VTAIL.n627 VTAIL.n626 9.3005
R681 VTAIL.n686 VTAIL.n685 9.3005
R682 VTAIL.n688 VTAIL.n687 9.3005
R683 VTAIL.n624 VTAIL.n621 9.3005
R684 VTAIL.n711 VTAIL.n710 9.3005
R685 VTAIL.n614 VTAIL.n613 9.3005
R686 VTAIL.n705 VTAIL.n704 9.3005
R687 VTAIL.n703 VTAIL.n702 9.3005
R688 VTAIL.n618 VTAIL.n617 9.3005
R689 VTAIL.n697 VTAIL.n696 9.3005
R690 VTAIL.n695 VTAIL.n694 9.3005
R691 VTAIL.n670 VTAIL.n669 9.3005
R692 VTAIL.n635 VTAIL.n634 9.3005
R693 VTAIL.n664 VTAIL.n663 9.3005
R694 VTAIL.n662 VTAIL.n661 9.3005
R695 VTAIL.n639 VTAIL.n638 9.3005
R696 VTAIL.n656 VTAIL.n655 9.3005
R697 VTAIL.n654 VTAIL.n653 9.3005
R698 VTAIL.n643 VTAIL.n642 9.3005
R699 VTAIL.n648 VTAIL.n647 9.3005
R700 VTAIL.n570 VTAIL.n569 9.3005
R701 VTAIL.n529 VTAIL.n528 9.3005
R702 VTAIL.n576 VTAIL.n575 9.3005
R703 VTAIL.n578 VTAIL.n577 9.3005
R704 VTAIL.n525 VTAIL.n524 9.3005
R705 VTAIL.n584 VTAIL.n583 9.3005
R706 VTAIL.n586 VTAIL.n585 9.3005
R707 VTAIL.n522 VTAIL.n519 9.3005
R708 VTAIL.n609 VTAIL.n608 9.3005
R709 VTAIL.n512 VTAIL.n511 9.3005
R710 VTAIL.n603 VTAIL.n602 9.3005
R711 VTAIL.n601 VTAIL.n600 9.3005
R712 VTAIL.n516 VTAIL.n515 9.3005
R713 VTAIL.n595 VTAIL.n594 9.3005
R714 VTAIL.n593 VTAIL.n592 9.3005
R715 VTAIL.n568 VTAIL.n567 9.3005
R716 VTAIL.n533 VTAIL.n532 9.3005
R717 VTAIL.n562 VTAIL.n561 9.3005
R718 VTAIL.n560 VTAIL.n559 9.3005
R719 VTAIL.n537 VTAIL.n536 9.3005
R720 VTAIL.n554 VTAIL.n553 9.3005
R721 VTAIL.n552 VTAIL.n551 9.3005
R722 VTAIL.n541 VTAIL.n540 9.3005
R723 VTAIL.n546 VTAIL.n545 9.3005
R724 VTAIL.n468 VTAIL.n467 9.3005
R725 VTAIL.n427 VTAIL.n426 9.3005
R726 VTAIL.n474 VTAIL.n473 9.3005
R727 VTAIL.n476 VTAIL.n475 9.3005
R728 VTAIL.n423 VTAIL.n422 9.3005
R729 VTAIL.n482 VTAIL.n481 9.3005
R730 VTAIL.n484 VTAIL.n483 9.3005
R731 VTAIL.n420 VTAIL.n417 9.3005
R732 VTAIL.n507 VTAIL.n506 9.3005
R733 VTAIL.n410 VTAIL.n409 9.3005
R734 VTAIL.n501 VTAIL.n500 9.3005
R735 VTAIL.n499 VTAIL.n498 9.3005
R736 VTAIL.n414 VTAIL.n413 9.3005
R737 VTAIL.n493 VTAIL.n492 9.3005
R738 VTAIL.n491 VTAIL.n490 9.3005
R739 VTAIL.n466 VTAIL.n465 9.3005
R740 VTAIL.n431 VTAIL.n430 9.3005
R741 VTAIL.n460 VTAIL.n459 9.3005
R742 VTAIL.n458 VTAIL.n457 9.3005
R743 VTAIL.n435 VTAIL.n434 9.3005
R744 VTAIL.n452 VTAIL.n451 9.3005
R745 VTAIL.n450 VTAIL.n449 9.3005
R746 VTAIL.n439 VTAIL.n438 9.3005
R747 VTAIL.n444 VTAIL.n443 9.3005
R748 VTAIL.n366 VTAIL.n365 9.3005
R749 VTAIL.n325 VTAIL.n324 9.3005
R750 VTAIL.n372 VTAIL.n371 9.3005
R751 VTAIL.n374 VTAIL.n373 9.3005
R752 VTAIL.n321 VTAIL.n320 9.3005
R753 VTAIL.n380 VTAIL.n379 9.3005
R754 VTAIL.n382 VTAIL.n381 9.3005
R755 VTAIL.n318 VTAIL.n315 9.3005
R756 VTAIL.n405 VTAIL.n404 9.3005
R757 VTAIL.n308 VTAIL.n307 9.3005
R758 VTAIL.n399 VTAIL.n398 9.3005
R759 VTAIL.n397 VTAIL.n396 9.3005
R760 VTAIL.n312 VTAIL.n311 9.3005
R761 VTAIL.n391 VTAIL.n390 9.3005
R762 VTAIL.n389 VTAIL.n388 9.3005
R763 VTAIL.n364 VTAIL.n363 9.3005
R764 VTAIL.n329 VTAIL.n328 9.3005
R765 VTAIL.n358 VTAIL.n357 9.3005
R766 VTAIL.n356 VTAIL.n355 9.3005
R767 VTAIL.n333 VTAIL.n332 9.3005
R768 VTAIL.n350 VTAIL.n349 9.3005
R769 VTAIL.n348 VTAIL.n347 9.3005
R770 VTAIL.n337 VTAIL.n336 9.3005
R771 VTAIL.n342 VTAIL.n341 9.3005
R772 VTAIL.n762 VTAIL.n738 8.92171
R773 VTAIL.n778 VTAIL.n777 8.92171
R774 VTAIL.n811 VTAIL.n716 8.92171
R775 VTAIL.n48 VTAIL.n24 8.92171
R776 VTAIL.n64 VTAIL.n63 8.92171
R777 VTAIL.n97 VTAIL.n2 8.92171
R778 VTAIL.n150 VTAIL.n126 8.92171
R779 VTAIL.n166 VTAIL.n165 8.92171
R780 VTAIL.n199 VTAIL.n104 8.92171
R781 VTAIL.n252 VTAIL.n228 8.92171
R782 VTAIL.n268 VTAIL.n267 8.92171
R783 VTAIL.n301 VTAIL.n206 8.92171
R784 VTAIL.n709 VTAIL.n614 8.92171
R785 VTAIL.n677 VTAIL.n676 8.92171
R786 VTAIL.n661 VTAIL.n637 8.92171
R787 VTAIL.n607 VTAIL.n512 8.92171
R788 VTAIL.n575 VTAIL.n574 8.92171
R789 VTAIL.n559 VTAIL.n535 8.92171
R790 VTAIL.n505 VTAIL.n410 8.92171
R791 VTAIL.n473 VTAIL.n472 8.92171
R792 VTAIL.n457 VTAIL.n433 8.92171
R793 VTAIL.n403 VTAIL.n308 8.92171
R794 VTAIL.n371 VTAIL.n370 8.92171
R795 VTAIL.n355 VTAIL.n331 8.92171
R796 VTAIL.n766 VTAIL.n765 8.14595
R797 VTAIL.n774 VTAIL.n732 8.14595
R798 VTAIL.n812 VTAIL.n714 8.14595
R799 VTAIL.n52 VTAIL.n51 8.14595
R800 VTAIL.n60 VTAIL.n18 8.14595
R801 VTAIL.n98 VTAIL.n0 8.14595
R802 VTAIL.n154 VTAIL.n153 8.14595
R803 VTAIL.n162 VTAIL.n120 8.14595
R804 VTAIL.n200 VTAIL.n102 8.14595
R805 VTAIL.n256 VTAIL.n255 8.14595
R806 VTAIL.n264 VTAIL.n222 8.14595
R807 VTAIL.n302 VTAIL.n204 8.14595
R808 VTAIL.n710 VTAIL.n612 8.14595
R809 VTAIL.n673 VTAIL.n631 8.14595
R810 VTAIL.n665 VTAIL.n664 8.14595
R811 VTAIL.n608 VTAIL.n510 8.14595
R812 VTAIL.n571 VTAIL.n529 8.14595
R813 VTAIL.n563 VTAIL.n562 8.14595
R814 VTAIL.n506 VTAIL.n408 8.14595
R815 VTAIL.n469 VTAIL.n427 8.14595
R816 VTAIL.n461 VTAIL.n460 8.14595
R817 VTAIL.n404 VTAIL.n306 8.14595
R818 VTAIL.n367 VTAIL.n325 8.14595
R819 VTAIL.n359 VTAIL.n358 8.14595
R820 VTAIL.n769 VTAIL.n736 7.3702
R821 VTAIL.n773 VTAIL.n734 7.3702
R822 VTAIL.n55 VTAIL.n22 7.3702
R823 VTAIL.n59 VTAIL.n20 7.3702
R824 VTAIL.n157 VTAIL.n124 7.3702
R825 VTAIL.n161 VTAIL.n122 7.3702
R826 VTAIL.n259 VTAIL.n226 7.3702
R827 VTAIL.n263 VTAIL.n224 7.3702
R828 VTAIL.n672 VTAIL.n633 7.3702
R829 VTAIL.n668 VTAIL.n635 7.3702
R830 VTAIL.n570 VTAIL.n531 7.3702
R831 VTAIL.n566 VTAIL.n533 7.3702
R832 VTAIL.n468 VTAIL.n429 7.3702
R833 VTAIL.n464 VTAIL.n431 7.3702
R834 VTAIL.n366 VTAIL.n327 7.3702
R835 VTAIL.n362 VTAIL.n329 7.3702
R836 VTAIL.n770 VTAIL.n769 6.59444
R837 VTAIL.n770 VTAIL.n734 6.59444
R838 VTAIL.n56 VTAIL.n55 6.59444
R839 VTAIL.n56 VTAIL.n20 6.59444
R840 VTAIL.n158 VTAIL.n157 6.59444
R841 VTAIL.n158 VTAIL.n122 6.59444
R842 VTAIL.n260 VTAIL.n259 6.59444
R843 VTAIL.n260 VTAIL.n224 6.59444
R844 VTAIL.n669 VTAIL.n633 6.59444
R845 VTAIL.n669 VTAIL.n668 6.59444
R846 VTAIL.n567 VTAIL.n531 6.59444
R847 VTAIL.n567 VTAIL.n566 6.59444
R848 VTAIL.n465 VTAIL.n429 6.59444
R849 VTAIL.n465 VTAIL.n464 6.59444
R850 VTAIL.n363 VTAIL.n327 6.59444
R851 VTAIL.n363 VTAIL.n362 6.59444
R852 VTAIL.n766 VTAIL.n736 5.81868
R853 VTAIL.n774 VTAIL.n773 5.81868
R854 VTAIL.n814 VTAIL.n714 5.81868
R855 VTAIL.n52 VTAIL.n22 5.81868
R856 VTAIL.n60 VTAIL.n59 5.81868
R857 VTAIL.n100 VTAIL.n0 5.81868
R858 VTAIL.n154 VTAIL.n124 5.81868
R859 VTAIL.n162 VTAIL.n161 5.81868
R860 VTAIL.n202 VTAIL.n102 5.81868
R861 VTAIL.n256 VTAIL.n226 5.81868
R862 VTAIL.n264 VTAIL.n263 5.81868
R863 VTAIL.n304 VTAIL.n204 5.81868
R864 VTAIL.n712 VTAIL.n612 5.81868
R865 VTAIL.n673 VTAIL.n672 5.81868
R866 VTAIL.n665 VTAIL.n635 5.81868
R867 VTAIL.n610 VTAIL.n510 5.81868
R868 VTAIL.n571 VTAIL.n570 5.81868
R869 VTAIL.n563 VTAIL.n533 5.81868
R870 VTAIL.n508 VTAIL.n408 5.81868
R871 VTAIL.n469 VTAIL.n468 5.81868
R872 VTAIL.n461 VTAIL.n431 5.81868
R873 VTAIL.n406 VTAIL.n306 5.81868
R874 VTAIL.n367 VTAIL.n366 5.81868
R875 VTAIL.n359 VTAIL.n329 5.81868
R876 VTAIL.n765 VTAIL.n738 5.04292
R877 VTAIL.n777 VTAIL.n732 5.04292
R878 VTAIL.n812 VTAIL.n811 5.04292
R879 VTAIL.n51 VTAIL.n24 5.04292
R880 VTAIL.n63 VTAIL.n18 5.04292
R881 VTAIL.n98 VTAIL.n97 5.04292
R882 VTAIL.n153 VTAIL.n126 5.04292
R883 VTAIL.n165 VTAIL.n120 5.04292
R884 VTAIL.n200 VTAIL.n199 5.04292
R885 VTAIL.n255 VTAIL.n228 5.04292
R886 VTAIL.n267 VTAIL.n222 5.04292
R887 VTAIL.n302 VTAIL.n301 5.04292
R888 VTAIL.n710 VTAIL.n709 5.04292
R889 VTAIL.n676 VTAIL.n631 5.04292
R890 VTAIL.n664 VTAIL.n637 5.04292
R891 VTAIL.n608 VTAIL.n607 5.04292
R892 VTAIL.n574 VTAIL.n529 5.04292
R893 VTAIL.n562 VTAIL.n535 5.04292
R894 VTAIL.n506 VTAIL.n505 5.04292
R895 VTAIL.n472 VTAIL.n427 5.04292
R896 VTAIL.n460 VTAIL.n433 5.04292
R897 VTAIL.n404 VTAIL.n403 5.04292
R898 VTAIL.n370 VTAIL.n325 5.04292
R899 VTAIL.n358 VTAIL.n331 5.04292
R900 VTAIL.n748 VTAIL.n747 4.38563
R901 VTAIL.n34 VTAIL.n33 4.38563
R902 VTAIL.n136 VTAIL.n135 4.38563
R903 VTAIL.n238 VTAIL.n237 4.38563
R904 VTAIL.n647 VTAIL.n646 4.38563
R905 VTAIL.n545 VTAIL.n544 4.38563
R906 VTAIL.n443 VTAIL.n442 4.38563
R907 VTAIL.n341 VTAIL.n340 4.38563
R908 VTAIL.n762 VTAIL.n761 4.26717
R909 VTAIL.n778 VTAIL.n730 4.26717
R910 VTAIL.n808 VTAIL.n716 4.26717
R911 VTAIL.n48 VTAIL.n47 4.26717
R912 VTAIL.n64 VTAIL.n16 4.26717
R913 VTAIL.n94 VTAIL.n2 4.26717
R914 VTAIL.n150 VTAIL.n149 4.26717
R915 VTAIL.n166 VTAIL.n118 4.26717
R916 VTAIL.n196 VTAIL.n104 4.26717
R917 VTAIL.n252 VTAIL.n251 4.26717
R918 VTAIL.n268 VTAIL.n220 4.26717
R919 VTAIL.n298 VTAIL.n206 4.26717
R920 VTAIL.n706 VTAIL.n614 4.26717
R921 VTAIL.n677 VTAIL.n629 4.26717
R922 VTAIL.n661 VTAIL.n660 4.26717
R923 VTAIL.n604 VTAIL.n512 4.26717
R924 VTAIL.n575 VTAIL.n527 4.26717
R925 VTAIL.n559 VTAIL.n558 4.26717
R926 VTAIL.n502 VTAIL.n410 4.26717
R927 VTAIL.n473 VTAIL.n425 4.26717
R928 VTAIL.n457 VTAIL.n456 4.26717
R929 VTAIL.n400 VTAIL.n308 4.26717
R930 VTAIL.n371 VTAIL.n323 4.26717
R931 VTAIL.n355 VTAIL.n354 4.26717
R932 VTAIL.n758 VTAIL.n740 3.49141
R933 VTAIL.n782 VTAIL.n781 3.49141
R934 VTAIL.n807 VTAIL.n718 3.49141
R935 VTAIL.n44 VTAIL.n26 3.49141
R936 VTAIL.n68 VTAIL.n67 3.49141
R937 VTAIL.n93 VTAIL.n4 3.49141
R938 VTAIL.n146 VTAIL.n128 3.49141
R939 VTAIL.n170 VTAIL.n169 3.49141
R940 VTAIL.n195 VTAIL.n106 3.49141
R941 VTAIL.n248 VTAIL.n230 3.49141
R942 VTAIL.n272 VTAIL.n271 3.49141
R943 VTAIL.n297 VTAIL.n208 3.49141
R944 VTAIL.n705 VTAIL.n616 3.49141
R945 VTAIL.n681 VTAIL.n680 3.49141
R946 VTAIL.n657 VTAIL.n639 3.49141
R947 VTAIL.n603 VTAIL.n514 3.49141
R948 VTAIL.n579 VTAIL.n578 3.49141
R949 VTAIL.n555 VTAIL.n537 3.49141
R950 VTAIL.n501 VTAIL.n412 3.49141
R951 VTAIL.n477 VTAIL.n476 3.49141
R952 VTAIL.n453 VTAIL.n435 3.49141
R953 VTAIL.n399 VTAIL.n310 3.49141
R954 VTAIL.n375 VTAIL.n374 3.49141
R955 VTAIL.n351 VTAIL.n333 3.49141
R956 VTAIL.n757 VTAIL.n742 2.71565
R957 VTAIL.n785 VTAIL.n728 2.71565
R958 VTAIL.n804 VTAIL.n803 2.71565
R959 VTAIL.n43 VTAIL.n28 2.71565
R960 VTAIL.n71 VTAIL.n14 2.71565
R961 VTAIL.n90 VTAIL.n89 2.71565
R962 VTAIL.n145 VTAIL.n130 2.71565
R963 VTAIL.n173 VTAIL.n116 2.71565
R964 VTAIL.n192 VTAIL.n191 2.71565
R965 VTAIL.n247 VTAIL.n232 2.71565
R966 VTAIL.n275 VTAIL.n218 2.71565
R967 VTAIL.n294 VTAIL.n293 2.71565
R968 VTAIL.n702 VTAIL.n701 2.71565
R969 VTAIL.n684 VTAIL.n627 2.71565
R970 VTAIL.n656 VTAIL.n641 2.71565
R971 VTAIL.n600 VTAIL.n599 2.71565
R972 VTAIL.n582 VTAIL.n525 2.71565
R973 VTAIL.n554 VTAIL.n539 2.71565
R974 VTAIL.n498 VTAIL.n497 2.71565
R975 VTAIL.n480 VTAIL.n423 2.71565
R976 VTAIL.n452 VTAIL.n437 2.71565
R977 VTAIL.n396 VTAIL.n395 2.71565
R978 VTAIL.n378 VTAIL.n321 2.71565
R979 VTAIL.n350 VTAIL.n335 2.71565
R980 VTAIL.n754 VTAIL.n753 1.93989
R981 VTAIL.n786 VTAIL.n726 1.93989
R982 VTAIL.n800 VTAIL.n720 1.93989
R983 VTAIL.n40 VTAIL.n39 1.93989
R984 VTAIL.n72 VTAIL.n12 1.93989
R985 VTAIL.n86 VTAIL.n6 1.93989
R986 VTAIL.n142 VTAIL.n141 1.93989
R987 VTAIL.n174 VTAIL.n114 1.93989
R988 VTAIL.n188 VTAIL.n108 1.93989
R989 VTAIL.n244 VTAIL.n243 1.93989
R990 VTAIL.n276 VTAIL.n216 1.93989
R991 VTAIL.n290 VTAIL.n210 1.93989
R992 VTAIL.n698 VTAIL.n618 1.93989
R993 VTAIL.n685 VTAIL.n625 1.93989
R994 VTAIL.n653 VTAIL.n652 1.93989
R995 VTAIL.n596 VTAIL.n516 1.93989
R996 VTAIL.n583 VTAIL.n523 1.93989
R997 VTAIL.n551 VTAIL.n550 1.93989
R998 VTAIL.n494 VTAIL.n414 1.93989
R999 VTAIL.n481 VTAIL.n421 1.93989
R1000 VTAIL.n449 VTAIL.n448 1.93989
R1001 VTAIL.n392 VTAIL.n312 1.93989
R1002 VTAIL.n379 VTAIL.n319 1.93989
R1003 VTAIL.n347 VTAIL.n346 1.93989
R1004 VTAIL.n750 VTAIL.n744 1.16414
R1005 VTAIL.n791 VTAIL.n789 1.16414
R1006 VTAIL.n799 VTAIL.n722 1.16414
R1007 VTAIL.n36 VTAIL.n30 1.16414
R1008 VTAIL.n77 VTAIL.n75 1.16414
R1009 VTAIL.n85 VTAIL.n8 1.16414
R1010 VTAIL.n138 VTAIL.n132 1.16414
R1011 VTAIL.n179 VTAIL.n177 1.16414
R1012 VTAIL.n187 VTAIL.n110 1.16414
R1013 VTAIL.n240 VTAIL.n234 1.16414
R1014 VTAIL.n281 VTAIL.n279 1.16414
R1015 VTAIL.n289 VTAIL.n212 1.16414
R1016 VTAIL.n697 VTAIL.n620 1.16414
R1017 VTAIL.n689 VTAIL.n688 1.16414
R1018 VTAIL.n649 VTAIL.n643 1.16414
R1019 VTAIL.n595 VTAIL.n518 1.16414
R1020 VTAIL.n587 VTAIL.n586 1.16414
R1021 VTAIL.n547 VTAIL.n541 1.16414
R1022 VTAIL.n493 VTAIL.n416 1.16414
R1023 VTAIL.n485 VTAIL.n484 1.16414
R1024 VTAIL.n445 VTAIL.n439 1.16414
R1025 VTAIL.n391 VTAIL.n314 1.16414
R1026 VTAIL.n383 VTAIL.n382 1.16414
R1027 VTAIL.n343 VTAIL.n337 1.16414
R1028 VTAIL.n509 VTAIL.n407 0.733259
R1029 VTAIL.n713 VTAIL.n611 0.733259
R1030 VTAIL.n305 VTAIL.n203 0.733259
R1031 VTAIL.n611 VTAIL.n509 0.470328
R1032 VTAIL.n203 VTAIL.n101 0.470328
R1033 VTAIL VTAIL.n101 0.425069
R1034 VTAIL.n749 VTAIL.n746 0.388379
R1035 VTAIL.n790 VTAIL.n724 0.388379
R1036 VTAIL.n796 VTAIL.n795 0.388379
R1037 VTAIL.n35 VTAIL.n32 0.388379
R1038 VTAIL.n76 VTAIL.n10 0.388379
R1039 VTAIL.n82 VTAIL.n81 0.388379
R1040 VTAIL.n137 VTAIL.n134 0.388379
R1041 VTAIL.n178 VTAIL.n112 0.388379
R1042 VTAIL.n184 VTAIL.n183 0.388379
R1043 VTAIL.n239 VTAIL.n236 0.388379
R1044 VTAIL.n280 VTAIL.n214 0.388379
R1045 VTAIL.n286 VTAIL.n285 0.388379
R1046 VTAIL.n694 VTAIL.n693 0.388379
R1047 VTAIL.n624 VTAIL.n622 0.388379
R1048 VTAIL.n648 VTAIL.n645 0.388379
R1049 VTAIL.n592 VTAIL.n591 0.388379
R1050 VTAIL.n522 VTAIL.n520 0.388379
R1051 VTAIL.n546 VTAIL.n543 0.388379
R1052 VTAIL.n490 VTAIL.n489 0.388379
R1053 VTAIL.n420 VTAIL.n418 0.388379
R1054 VTAIL.n444 VTAIL.n441 0.388379
R1055 VTAIL.n388 VTAIL.n387 0.388379
R1056 VTAIL.n318 VTAIL.n316 0.388379
R1057 VTAIL.n342 VTAIL.n339 0.388379
R1058 VTAIL VTAIL.n815 0.30869
R1059 VTAIL.n748 VTAIL.n743 0.155672
R1060 VTAIL.n755 VTAIL.n743 0.155672
R1061 VTAIL.n756 VTAIL.n755 0.155672
R1062 VTAIL.n756 VTAIL.n739 0.155672
R1063 VTAIL.n763 VTAIL.n739 0.155672
R1064 VTAIL.n764 VTAIL.n763 0.155672
R1065 VTAIL.n764 VTAIL.n735 0.155672
R1066 VTAIL.n771 VTAIL.n735 0.155672
R1067 VTAIL.n772 VTAIL.n771 0.155672
R1068 VTAIL.n772 VTAIL.n731 0.155672
R1069 VTAIL.n779 VTAIL.n731 0.155672
R1070 VTAIL.n780 VTAIL.n779 0.155672
R1071 VTAIL.n780 VTAIL.n727 0.155672
R1072 VTAIL.n787 VTAIL.n727 0.155672
R1073 VTAIL.n788 VTAIL.n787 0.155672
R1074 VTAIL.n788 VTAIL.n723 0.155672
R1075 VTAIL.n797 VTAIL.n723 0.155672
R1076 VTAIL.n798 VTAIL.n797 0.155672
R1077 VTAIL.n798 VTAIL.n719 0.155672
R1078 VTAIL.n805 VTAIL.n719 0.155672
R1079 VTAIL.n806 VTAIL.n805 0.155672
R1080 VTAIL.n806 VTAIL.n715 0.155672
R1081 VTAIL.n813 VTAIL.n715 0.155672
R1082 VTAIL.n34 VTAIL.n29 0.155672
R1083 VTAIL.n41 VTAIL.n29 0.155672
R1084 VTAIL.n42 VTAIL.n41 0.155672
R1085 VTAIL.n42 VTAIL.n25 0.155672
R1086 VTAIL.n49 VTAIL.n25 0.155672
R1087 VTAIL.n50 VTAIL.n49 0.155672
R1088 VTAIL.n50 VTAIL.n21 0.155672
R1089 VTAIL.n57 VTAIL.n21 0.155672
R1090 VTAIL.n58 VTAIL.n57 0.155672
R1091 VTAIL.n58 VTAIL.n17 0.155672
R1092 VTAIL.n65 VTAIL.n17 0.155672
R1093 VTAIL.n66 VTAIL.n65 0.155672
R1094 VTAIL.n66 VTAIL.n13 0.155672
R1095 VTAIL.n73 VTAIL.n13 0.155672
R1096 VTAIL.n74 VTAIL.n73 0.155672
R1097 VTAIL.n74 VTAIL.n9 0.155672
R1098 VTAIL.n83 VTAIL.n9 0.155672
R1099 VTAIL.n84 VTAIL.n83 0.155672
R1100 VTAIL.n84 VTAIL.n5 0.155672
R1101 VTAIL.n91 VTAIL.n5 0.155672
R1102 VTAIL.n92 VTAIL.n91 0.155672
R1103 VTAIL.n92 VTAIL.n1 0.155672
R1104 VTAIL.n99 VTAIL.n1 0.155672
R1105 VTAIL.n136 VTAIL.n131 0.155672
R1106 VTAIL.n143 VTAIL.n131 0.155672
R1107 VTAIL.n144 VTAIL.n143 0.155672
R1108 VTAIL.n144 VTAIL.n127 0.155672
R1109 VTAIL.n151 VTAIL.n127 0.155672
R1110 VTAIL.n152 VTAIL.n151 0.155672
R1111 VTAIL.n152 VTAIL.n123 0.155672
R1112 VTAIL.n159 VTAIL.n123 0.155672
R1113 VTAIL.n160 VTAIL.n159 0.155672
R1114 VTAIL.n160 VTAIL.n119 0.155672
R1115 VTAIL.n167 VTAIL.n119 0.155672
R1116 VTAIL.n168 VTAIL.n167 0.155672
R1117 VTAIL.n168 VTAIL.n115 0.155672
R1118 VTAIL.n175 VTAIL.n115 0.155672
R1119 VTAIL.n176 VTAIL.n175 0.155672
R1120 VTAIL.n176 VTAIL.n111 0.155672
R1121 VTAIL.n185 VTAIL.n111 0.155672
R1122 VTAIL.n186 VTAIL.n185 0.155672
R1123 VTAIL.n186 VTAIL.n107 0.155672
R1124 VTAIL.n193 VTAIL.n107 0.155672
R1125 VTAIL.n194 VTAIL.n193 0.155672
R1126 VTAIL.n194 VTAIL.n103 0.155672
R1127 VTAIL.n201 VTAIL.n103 0.155672
R1128 VTAIL.n238 VTAIL.n233 0.155672
R1129 VTAIL.n245 VTAIL.n233 0.155672
R1130 VTAIL.n246 VTAIL.n245 0.155672
R1131 VTAIL.n246 VTAIL.n229 0.155672
R1132 VTAIL.n253 VTAIL.n229 0.155672
R1133 VTAIL.n254 VTAIL.n253 0.155672
R1134 VTAIL.n254 VTAIL.n225 0.155672
R1135 VTAIL.n261 VTAIL.n225 0.155672
R1136 VTAIL.n262 VTAIL.n261 0.155672
R1137 VTAIL.n262 VTAIL.n221 0.155672
R1138 VTAIL.n269 VTAIL.n221 0.155672
R1139 VTAIL.n270 VTAIL.n269 0.155672
R1140 VTAIL.n270 VTAIL.n217 0.155672
R1141 VTAIL.n277 VTAIL.n217 0.155672
R1142 VTAIL.n278 VTAIL.n277 0.155672
R1143 VTAIL.n278 VTAIL.n213 0.155672
R1144 VTAIL.n287 VTAIL.n213 0.155672
R1145 VTAIL.n288 VTAIL.n287 0.155672
R1146 VTAIL.n288 VTAIL.n209 0.155672
R1147 VTAIL.n295 VTAIL.n209 0.155672
R1148 VTAIL.n296 VTAIL.n295 0.155672
R1149 VTAIL.n296 VTAIL.n205 0.155672
R1150 VTAIL.n303 VTAIL.n205 0.155672
R1151 VTAIL.n711 VTAIL.n613 0.155672
R1152 VTAIL.n704 VTAIL.n613 0.155672
R1153 VTAIL.n704 VTAIL.n703 0.155672
R1154 VTAIL.n703 VTAIL.n617 0.155672
R1155 VTAIL.n696 VTAIL.n617 0.155672
R1156 VTAIL.n696 VTAIL.n695 0.155672
R1157 VTAIL.n695 VTAIL.n621 0.155672
R1158 VTAIL.n687 VTAIL.n621 0.155672
R1159 VTAIL.n687 VTAIL.n686 0.155672
R1160 VTAIL.n686 VTAIL.n626 0.155672
R1161 VTAIL.n679 VTAIL.n626 0.155672
R1162 VTAIL.n679 VTAIL.n678 0.155672
R1163 VTAIL.n678 VTAIL.n630 0.155672
R1164 VTAIL.n671 VTAIL.n630 0.155672
R1165 VTAIL.n671 VTAIL.n670 0.155672
R1166 VTAIL.n670 VTAIL.n634 0.155672
R1167 VTAIL.n663 VTAIL.n634 0.155672
R1168 VTAIL.n663 VTAIL.n662 0.155672
R1169 VTAIL.n662 VTAIL.n638 0.155672
R1170 VTAIL.n655 VTAIL.n638 0.155672
R1171 VTAIL.n655 VTAIL.n654 0.155672
R1172 VTAIL.n654 VTAIL.n642 0.155672
R1173 VTAIL.n647 VTAIL.n642 0.155672
R1174 VTAIL.n609 VTAIL.n511 0.155672
R1175 VTAIL.n602 VTAIL.n511 0.155672
R1176 VTAIL.n602 VTAIL.n601 0.155672
R1177 VTAIL.n601 VTAIL.n515 0.155672
R1178 VTAIL.n594 VTAIL.n515 0.155672
R1179 VTAIL.n594 VTAIL.n593 0.155672
R1180 VTAIL.n593 VTAIL.n519 0.155672
R1181 VTAIL.n585 VTAIL.n519 0.155672
R1182 VTAIL.n585 VTAIL.n584 0.155672
R1183 VTAIL.n584 VTAIL.n524 0.155672
R1184 VTAIL.n577 VTAIL.n524 0.155672
R1185 VTAIL.n577 VTAIL.n576 0.155672
R1186 VTAIL.n576 VTAIL.n528 0.155672
R1187 VTAIL.n569 VTAIL.n528 0.155672
R1188 VTAIL.n569 VTAIL.n568 0.155672
R1189 VTAIL.n568 VTAIL.n532 0.155672
R1190 VTAIL.n561 VTAIL.n532 0.155672
R1191 VTAIL.n561 VTAIL.n560 0.155672
R1192 VTAIL.n560 VTAIL.n536 0.155672
R1193 VTAIL.n553 VTAIL.n536 0.155672
R1194 VTAIL.n553 VTAIL.n552 0.155672
R1195 VTAIL.n552 VTAIL.n540 0.155672
R1196 VTAIL.n545 VTAIL.n540 0.155672
R1197 VTAIL.n507 VTAIL.n409 0.155672
R1198 VTAIL.n500 VTAIL.n409 0.155672
R1199 VTAIL.n500 VTAIL.n499 0.155672
R1200 VTAIL.n499 VTAIL.n413 0.155672
R1201 VTAIL.n492 VTAIL.n413 0.155672
R1202 VTAIL.n492 VTAIL.n491 0.155672
R1203 VTAIL.n491 VTAIL.n417 0.155672
R1204 VTAIL.n483 VTAIL.n417 0.155672
R1205 VTAIL.n483 VTAIL.n482 0.155672
R1206 VTAIL.n482 VTAIL.n422 0.155672
R1207 VTAIL.n475 VTAIL.n422 0.155672
R1208 VTAIL.n475 VTAIL.n474 0.155672
R1209 VTAIL.n474 VTAIL.n426 0.155672
R1210 VTAIL.n467 VTAIL.n426 0.155672
R1211 VTAIL.n467 VTAIL.n466 0.155672
R1212 VTAIL.n466 VTAIL.n430 0.155672
R1213 VTAIL.n459 VTAIL.n430 0.155672
R1214 VTAIL.n459 VTAIL.n458 0.155672
R1215 VTAIL.n458 VTAIL.n434 0.155672
R1216 VTAIL.n451 VTAIL.n434 0.155672
R1217 VTAIL.n451 VTAIL.n450 0.155672
R1218 VTAIL.n450 VTAIL.n438 0.155672
R1219 VTAIL.n443 VTAIL.n438 0.155672
R1220 VTAIL.n405 VTAIL.n307 0.155672
R1221 VTAIL.n398 VTAIL.n307 0.155672
R1222 VTAIL.n398 VTAIL.n397 0.155672
R1223 VTAIL.n397 VTAIL.n311 0.155672
R1224 VTAIL.n390 VTAIL.n311 0.155672
R1225 VTAIL.n390 VTAIL.n389 0.155672
R1226 VTAIL.n389 VTAIL.n315 0.155672
R1227 VTAIL.n381 VTAIL.n315 0.155672
R1228 VTAIL.n381 VTAIL.n380 0.155672
R1229 VTAIL.n380 VTAIL.n320 0.155672
R1230 VTAIL.n373 VTAIL.n320 0.155672
R1231 VTAIL.n373 VTAIL.n372 0.155672
R1232 VTAIL.n372 VTAIL.n324 0.155672
R1233 VTAIL.n365 VTAIL.n324 0.155672
R1234 VTAIL.n365 VTAIL.n364 0.155672
R1235 VTAIL.n364 VTAIL.n328 0.155672
R1236 VTAIL.n357 VTAIL.n328 0.155672
R1237 VTAIL.n357 VTAIL.n356 0.155672
R1238 VTAIL.n356 VTAIL.n332 0.155672
R1239 VTAIL.n349 VTAIL.n332 0.155672
R1240 VTAIL.n349 VTAIL.n348 0.155672
R1241 VTAIL.n348 VTAIL.n336 0.155672
R1242 VTAIL.n341 VTAIL.n336 0.155672
R1243 VDD1 VDD1.n1 100.784
R1244 VDD1 VDD1.n0 58.7669
R1245 VDD1.n0 VDD1.t1 1.09201
R1246 VDD1.n0 VDD1.t3 1.09201
R1247 VDD1.n1 VDD1.t0 1.09201
R1248 VDD1.n1 VDD1.t2 1.09201
R1249 B.n101 B.t4 1046.66
R1250 B.n99 B.t15 1046.66
R1251 B.n450 B.t12 1046.66
R1252 B.n448 B.t8 1046.66
R1253 B.n779 B.n778 585
R1254 B.n780 B.n779 585
R1255 B.n355 B.n97 585
R1256 B.n354 B.n353 585
R1257 B.n352 B.n351 585
R1258 B.n350 B.n349 585
R1259 B.n348 B.n347 585
R1260 B.n346 B.n345 585
R1261 B.n344 B.n343 585
R1262 B.n342 B.n341 585
R1263 B.n340 B.n339 585
R1264 B.n338 B.n337 585
R1265 B.n336 B.n335 585
R1266 B.n334 B.n333 585
R1267 B.n332 B.n331 585
R1268 B.n330 B.n329 585
R1269 B.n328 B.n327 585
R1270 B.n326 B.n325 585
R1271 B.n324 B.n323 585
R1272 B.n322 B.n321 585
R1273 B.n320 B.n319 585
R1274 B.n318 B.n317 585
R1275 B.n316 B.n315 585
R1276 B.n314 B.n313 585
R1277 B.n312 B.n311 585
R1278 B.n310 B.n309 585
R1279 B.n308 B.n307 585
R1280 B.n306 B.n305 585
R1281 B.n304 B.n303 585
R1282 B.n302 B.n301 585
R1283 B.n300 B.n299 585
R1284 B.n298 B.n297 585
R1285 B.n296 B.n295 585
R1286 B.n294 B.n293 585
R1287 B.n292 B.n291 585
R1288 B.n290 B.n289 585
R1289 B.n288 B.n287 585
R1290 B.n286 B.n285 585
R1291 B.n284 B.n283 585
R1292 B.n282 B.n281 585
R1293 B.n280 B.n279 585
R1294 B.n278 B.n277 585
R1295 B.n276 B.n275 585
R1296 B.n274 B.n273 585
R1297 B.n272 B.n271 585
R1298 B.n270 B.n269 585
R1299 B.n268 B.n267 585
R1300 B.n266 B.n265 585
R1301 B.n264 B.n263 585
R1302 B.n262 B.n261 585
R1303 B.n260 B.n259 585
R1304 B.n258 B.n257 585
R1305 B.n256 B.n255 585
R1306 B.n254 B.n253 585
R1307 B.n252 B.n251 585
R1308 B.n250 B.n249 585
R1309 B.n248 B.n247 585
R1310 B.n246 B.n245 585
R1311 B.n244 B.n243 585
R1312 B.n242 B.n241 585
R1313 B.n240 B.n239 585
R1314 B.n237 B.n236 585
R1315 B.n235 B.n234 585
R1316 B.n233 B.n232 585
R1317 B.n231 B.n230 585
R1318 B.n229 B.n228 585
R1319 B.n227 B.n226 585
R1320 B.n225 B.n224 585
R1321 B.n223 B.n222 585
R1322 B.n221 B.n220 585
R1323 B.n219 B.n218 585
R1324 B.n217 B.n216 585
R1325 B.n215 B.n214 585
R1326 B.n213 B.n212 585
R1327 B.n211 B.n210 585
R1328 B.n209 B.n208 585
R1329 B.n207 B.n206 585
R1330 B.n205 B.n204 585
R1331 B.n203 B.n202 585
R1332 B.n201 B.n200 585
R1333 B.n199 B.n198 585
R1334 B.n197 B.n196 585
R1335 B.n195 B.n194 585
R1336 B.n193 B.n192 585
R1337 B.n191 B.n190 585
R1338 B.n189 B.n188 585
R1339 B.n187 B.n186 585
R1340 B.n185 B.n184 585
R1341 B.n183 B.n182 585
R1342 B.n181 B.n180 585
R1343 B.n179 B.n178 585
R1344 B.n177 B.n176 585
R1345 B.n175 B.n174 585
R1346 B.n173 B.n172 585
R1347 B.n171 B.n170 585
R1348 B.n169 B.n168 585
R1349 B.n167 B.n166 585
R1350 B.n165 B.n164 585
R1351 B.n163 B.n162 585
R1352 B.n161 B.n160 585
R1353 B.n159 B.n158 585
R1354 B.n157 B.n156 585
R1355 B.n155 B.n154 585
R1356 B.n153 B.n152 585
R1357 B.n151 B.n150 585
R1358 B.n149 B.n148 585
R1359 B.n147 B.n146 585
R1360 B.n145 B.n144 585
R1361 B.n143 B.n142 585
R1362 B.n141 B.n140 585
R1363 B.n139 B.n138 585
R1364 B.n137 B.n136 585
R1365 B.n135 B.n134 585
R1366 B.n133 B.n132 585
R1367 B.n131 B.n130 585
R1368 B.n129 B.n128 585
R1369 B.n127 B.n126 585
R1370 B.n125 B.n124 585
R1371 B.n123 B.n122 585
R1372 B.n121 B.n120 585
R1373 B.n119 B.n118 585
R1374 B.n117 B.n116 585
R1375 B.n115 B.n114 585
R1376 B.n113 B.n112 585
R1377 B.n111 B.n110 585
R1378 B.n109 B.n108 585
R1379 B.n107 B.n106 585
R1380 B.n105 B.n104 585
R1381 B.n33 B.n32 585
R1382 B.n783 B.n782 585
R1383 B.n777 B.n98 585
R1384 B.n98 B.n30 585
R1385 B.n776 B.n29 585
R1386 B.n787 B.n29 585
R1387 B.n775 B.n28 585
R1388 B.n788 B.n28 585
R1389 B.n774 B.n27 585
R1390 B.n789 B.n27 585
R1391 B.n773 B.n772 585
R1392 B.n772 B.n26 585
R1393 B.n771 B.n22 585
R1394 B.n795 B.n22 585
R1395 B.n770 B.n21 585
R1396 B.n796 B.n21 585
R1397 B.n769 B.n20 585
R1398 B.n797 B.n20 585
R1399 B.n768 B.n767 585
R1400 B.n767 B.n16 585
R1401 B.n766 B.n15 585
R1402 B.n803 B.n15 585
R1403 B.n765 B.n14 585
R1404 B.n804 B.n14 585
R1405 B.n764 B.n13 585
R1406 B.n805 B.n13 585
R1407 B.n763 B.n762 585
R1408 B.n762 B.n12 585
R1409 B.n761 B.n760 585
R1410 B.n761 B.n8 585
R1411 B.n759 B.n7 585
R1412 B.n812 B.n7 585
R1413 B.n758 B.n6 585
R1414 B.n813 B.n6 585
R1415 B.n757 B.n5 585
R1416 B.n814 B.n5 585
R1417 B.n756 B.n755 585
R1418 B.n755 B.n4 585
R1419 B.n754 B.n356 585
R1420 B.n754 B.n753 585
R1421 B.n743 B.n357 585
R1422 B.n746 B.n357 585
R1423 B.n745 B.n744 585
R1424 B.n747 B.n745 585
R1425 B.n742 B.n361 585
R1426 B.n365 B.n361 585
R1427 B.n741 B.n740 585
R1428 B.n740 B.n739 585
R1429 B.n363 B.n362 585
R1430 B.n364 B.n363 585
R1431 B.n732 B.n731 585
R1432 B.n733 B.n732 585
R1433 B.n730 B.n370 585
R1434 B.n370 B.n369 585
R1435 B.n729 B.n728 585
R1436 B.n728 B.n727 585
R1437 B.n372 B.n371 585
R1438 B.n720 B.n372 585
R1439 B.n719 B.n718 585
R1440 B.n721 B.n719 585
R1441 B.n717 B.n377 585
R1442 B.n377 B.n376 585
R1443 B.n716 B.n715 585
R1444 B.n715 B.n714 585
R1445 B.n379 B.n378 585
R1446 B.n380 B.n379 585
R1447 B.n710 B.n709 585
R1448 B.n383 B.n382 585
R1449 B.n706 B.n705 585
R1450 B.n707 B.n706 585
R1451 B.n704 B.n447 585
R1452 B.n703 B.n702 585
R1453 B.n701 B.n700 585
R1454 B.n699 B.n698 585
R1455 B.n697 B.n696 585
R1456 B.n695 B.n694 585
R1457 B.n693 B.n692 585
R1458 B.n691 B.n690 585
R1459 B.n689 B.n688 585
R1460 B.n687 B.n686 585
R1461 B.n685 B.n684 585
R1462 B.n683 B.n682 585
R1463 B.n681 B.n680 585
R1464 B.n679 B.n678 585
R1465 B.n677 B.n676 585
R1466 B.n675 B.n674 585
R1467 B.n673 B.n672 585
R1468 B.n671 B.n670 585
R1469 B.n669 B.n668 585
R1470 B.n667 B.n666 585
R1471 B.n665 B.n664 585
R1472 B.n663 B.n662 585
R1473 B.n661 B.n660 585
R1474 B.n659 B.n658 585
R1475 B.n657 B.n656 585
R1476 B.n655 B.n654 585
R1477 B.n653 B.n652 585
R1478 B.n651 B.n650 585
R1479 B.n649 B.n648 585
R1480 B.n647 B.n646 585
R1481 B.n645 B.n644 585
R1482 B.n643 B.n642 585
R1483 B.n641 B.n640 585
R1484 B.n639 B.n638 585
R1485 B.n637 B.n636 585
R1486 B.n635 B.n634 585
R1487 B.n633 B.n632 585
R1488 B.n631 B.n630 585
R1489 B.n629 B.n628 585
R1490 B.n627 B.n626 585
R1491 B.n625 B.n624 585
R1492 B.n623 B.n622 585
R1493 B.n621 B.n620 585
R1494 B.n619 B.n618 585
R1495 B.n617 B.n616 585
R1496 B.n615 B.n614 585
R1497 B.n613 B.n612 585
R1498 B.n611 B.n610 585
R1499 B.n609 B.n608 585
R1500 B.n607 B.n606 585
R1501 B.n605 B.n604 585
R1502 B.n603 B.n602 585
R1503 B.n601 B.n600 585
R1504 B.n599 B.n598 585
R1505 B.n597 B.n596 585
R1506 B.n595 B.n594 585
R1507 B.n593 B.n592 585
R1508 B.n590 B.n589 585
R1509 B.n588 B.n587 585
R1510 B.n586 B.n585 585
R1511 B.n584 B.n583 585
R1512 B.n582 B.n581 585
R1513 B.n580 B.n579 585
R1514 B.n578 B.n577 585
R1515 B.n576 B.n575 585
R1516 B.n574 B.n573 585
R1517 B.n572 B.n571 585
R1518 B.n570 B.n569 585
R1519 B.n568 B.n567 585
R1520 B.n566 B.n565 585
R1521 B.n564 B.n563 585
R1522 B.n562 B.n561 585
R1523 B.n560 B.n559 585
R1524 B.n558 B.n557 585
R1525 B.n556 B.n555 585
R1526 B.n554 B.n553 585
R1527 B.n552 B.n551 585
R1528 B.n550 B.n549 585
R1529 B.n548 B.n547 585
R1530 B.n546 B.n545 585
R1531 B.n544 B.n543 585
R1532 B.n542 B.n541 585
R1533 B.n540 B.n539 585
R1534 B.n538 B.n537 585
R1535 B.n536 B.n535 585
R1536 B.n534 B.n533 585
R1537 B.n532 B.n531 585
R1538 B.n530 B.n529 585
R1539 B.n528 B.n527 585
R1540 B.n526 B.n525 585
R1541 B.n524 B.n523 585
R1542 B.n522 B.n521 585
R1543 B.n520 B.n519 585
R1544 B.n518 B.n517 585
R1545 B.n516 B.n515 585
R1546 B.n514 B.n513 585
R1547 B.n512 B.n511 585
R1548 B.n510 B.n509 585
R1549 B.n508 B.n507 585
R1550 B.n506 B.n505 585
R1551 B.n504 B.n503 585
R1552 B.n502 B.n501 585
R1553 B.n500 B.n499 585
R1554 B.n498 B.n497 585
R1555 B.n496 B.n495 585
R1556 B.n494 B.n493 585
R1557 B.n492 B.n491 585
R1558 B.n490 B.n489 585
R1559 B.n488 B.n487 585
R1560 B.n486 B.n485 585
R1561 B.n484 B.n483 585
R1562 B.n482 B.n481 585
R1563 B.n480 B.n479 585
R1564 B.n478 B.n477 585
R1565 B.n476 B.n475 585
R1566 B.n474 B.n473 585
R1567 B.n472 B.n471 585
R1568 B.n470 B.n469 585
R1569 B.n468 B.n467 585
R1570 B.n466 B.n465 585
R1571 B.n464 B.n463 585
R1572 B.n462 B.n461 585
R1573 B.n460 B.n459 585
R1574 B.n458 B.n457 585
R1575 B.n456 B.n455 585
R1576 B.n454 B.n453 585
R1577 B.n711 B.n381 585
R1578 B.n381 B.n380 585
R1579 B.n713 B.n712 585
R1580 B.n714 B.n713 585
R1581 B.n375 B.n374 585
R1582 B.n376 B.n375 585
R1583 B.n723 B.n722 585
R1584 B.n722 B.n721 585
R1585 B.n724 B.n373 585
R1586 B.n720 B.n373 585
R1587 B.n726 B.n725 585
R1588 B.n727 B.n726 585
R1589 B.n368 B.n367 585
R1590 B.n369 B.n368 585
R1591 B.n735 B.n734 585
R1592 B.n734 B.n733 585
R1593 B.n736 B.n366 585
R1594 B.n366 B.n364 585
R1595 B.n738 B.n737 585
R1596 B.n739 B.n738 585
R1597 B.n360 B.n359 585
R1598 B.n365 B.n360 585
R1599 B.n749 B.n748 585
R1600 B.n748 B.n747 585
R1601 B.n750 B.n358 585
R1602 B.n746 B.n358 585
R1603 B.n752 B.n751 585
R1604 B.n753 B.n752 585
R1605 B.n3 B.n0 585
R1606 B.n4 B.n3 585
R1607 B.n811 B.n1 585
R1608 B.n812 B.n811 585
R1609 B.n810 B.n809 585
R1610 B.n810 B.n8 585
R1611 B.n808 B.n9 585
R1612 B.n12 B.n9 585
R1613 B.n807 B.n806 585
R1614 B.n806 B.n805 585
R1615 B.n11 B.n10 585
R1616 B.n804 B.n11 585
R1617 B.n802 B.n801 585
R1618 B.n803 B.n802 585
R1619 B.n800 B.n17 585
R1620 B.n17 B.n16 585
R1621 B.n799 B.n798 585
R1622 B.n798 B.n797 585
R1623 B.n19 B.n18 585
R1624 B.n796 B.n19 585
R1625 B.n794 B.n793 585
R1626 B.n795 B.n794 585
R1627 B.n792 B.n23 585
R1628 B.n26 B.n23 585
R1629 B.n791 B.n790 585
R1630 B.n790 B.n789 585
R1631 B.n25 B.n24 585
R1632 B.n788 B.n25 585
R1633 B.n786 B.n785 585
R1634 B.n787 B.n786 585
R1635 B.n784 B.n31 585
R1636 B.n31 B.n30 585
R1637 B.n815 B.n814 585
R1638 B.n813 B.n2 585
R1639 B.n782 B.n31 511.721
R1640 B.n779 B.n98 511.721
R1641 B.n453 B.n379 511.721
R1642 B.n709 B.n381 511.721
R1643 B.n99 B.t16 404.293
R1644 B.n450 B.t14 404.293
R1645 B.n101 B.t6 404.293
R1646 B.n448 B.t11 404.293
R1647 B.n100 B.t17 387.808
R1648 B.n451 B.t13 387.808
R1649 B.n102 B.t7 387.808
R1650 B.n449 B.t10 387.808
R1651 B.n780 B.n96 256.663
R1652 B.n780 B.n95 256.663
R1653 B.n780 B.n94 256.663
R1654 B.n780 B.n93 256.663
R1655 B.n780 B.n92 256.663
R1656 B.n780 B.n91 256.663
R1657 B.n780 B.n90 256.663
R1658 B.n780 B.n89 256.663
R1659 B.n780 B.n88 256.663
R1660 B.n780 B.n87 256.663
R1661 B.n780 B.n86 256.663
R1662 B.n780 B.n85 256.663
R1663 B.n780 B.n84 256.663
R1664 B.n780 B.n83 256.663
R1665 B.n780 B.n82 256.663
R1666 B.n780 B.n81 256.663
R1667 B.n780 B.n80 256.663
R1668 B.n780 B.n79 256.663
R1669 B.n780 B.n78 256.663
R1670 B.n780 B.n77 256.663
R1671 B.n780 B.n76 256.663
R1672 B.n780 B.n75 256.663
R1673 B.n780 B.n74 256.663
R1674 B.n780 B.n73 256.663
R1675 B.n780 B.n72 256.663
R1676 B.n780 B.n71 256.663
R1677 B.n780 B.n70 256.663
R1678 B.n780 B.n69 256.663
R1679 B.n780 B.n68 256.663
R1680 B.n780 B.n67 256.663
R1681 B.n780 B.n66 256.663
R1682 B.n780 B.n65 256.663
R1683 B.n780 B.n64 256.663
R1684 B.n780 B.n63 256.663
R1685 B.n780 B.n62 256.663
R1686 B.n780 B.n61 256.663
R1687 B.n780 B.n60 256.663
R1688 B.n780 B.n59 256.663
R1689 B.n780 B.n58 256.663
R1690 B.n780 B.n57 256.663
R1691 B.n780 B.n56 256.663
R1692 B.n780 B.n55 256.663
R1693 B.n780 B.n54 256.663
R1694 B.n780 B.n53 256.663
R1695 B.n780 B.n52 256.663
R1696 B.n780 B.n51 256.663
R1697 B.n780 B.n50 256.663
R1698 B.n780 B.n49 256.663
R1699 B.n780 B.n48 256.663
R1700 B.n780 B.n47 256.663
R1701 B.n780 B.n46 256.663
R1702 B.n780 B.n45 256.663
R1703 B.n780 B.n44 256.663
R1704 B.n780 B.n43 256.663
R1705 B.n780 B.n42 256.663
R1706 B.n780 B.n41 256.663
R1707 B.n780 B.n40 256.663
R1708 B.n780 B.n39 256.663
R1709 B.n780 B.n38 256.663
R1710 B.n780 B.n37 256.663
R1711 B.n780 B.n36 256.663
R1712 B.n780 B.n35 256.663
R1713 B.n780 B.n34 256.663
R1714 B.n781 B.n780 256.663
R1715 B.n708 B.n707 256.663
R1716 B.n707 B.n384 256.663
R1717 B.n707 B.n385 256.663
R1718 B.n707 B.n386 256.663
R1719 B.n707 B.n387 256.663
R1720 B.n707 B.n388 256.663
R1721 B.n707 B.n389 256.663
R1722 B.n707 B.n390 256.663
R1723 B.n707 B.n391 256.663
R1724 B.n707 B.n392 256.663
R1725 B.n707 B.n393 256.663
R1726 B.n707 B.n394 256.663
R1727 B.n707 B.n395 256.663
R1728 B.n707 B.n396 256.663
R1729 B.n707 B.n397 256.663
R1730 B.n707 B.n398 256.663
R1731 B.n707 B.n399 256.663
R1732 B.n707 B.n400 256.663
R1733 B.n707 B.n401 256.663
R1734 B.n707 B.n402 256.663
R1735 B.n707 B.n403 256.663
R1736 B.n707 B.n404 256.663
R1737 B.n707 B.n405 256.663
R1738 B.n707 B.n406 256.663
R1739 B.n707 B.n407 256.663
R1740 B.n707 B.n408 256.663
R1741 B.n707 B.n409 256.663
R1742 B.n707 B.n410 256.663
R1743 B.n707 B.n411 256.663
R1744 B.n707 B.n412 256.663
R1745 B.n707 B.n413 256.663
R1746 B.n707 B.n414 256.663
R1747 B.n707 B.n415 256.663
R1748 B.n707 B.n416 256.663
R1749 B.n707 B.n417 256.663
R1750 B.n707 B.n418 256.663
R1751 B.n707 B.n419 256.663
R1752 B.n707 B.n420 256.663
R1753 B.n707 B.n421 256.663
R1754 B.n707 B.n422 256.663
R1755 B.n707 B.n423 256.663
R1756 B.n707 B.n424 256.663
R1757 B.n707 B.n425 256.663
R1758 B.n707 B.n426 256.663
R1759 B.n707 B.n427 256.663
R1760 B.n707 B.n428 256.663
R1761 B.n707 B.n429 256.663
R1762 B.n707 B.n430 256.663
R1763 B.n707 B.n431 256.663
R1764 B.n707 B.n432 256.663
R1765 B.n707 B.n433 256.663
R1766 B.n707 B.n434 256.663
R1767 B.n707 B.n435 256.663
R1768 B.n707 B.n436 256.663
R1769 B.n707 B.n437 256.663
R1770 B.n707 B.n438 256.663
R1771 B.n707 B.n439 256.663
R1772 B.n707 B.n440 256.663
R1773 B.n707 B.n441 256.663
R1774 B.n707 B.n442 256.663
R1775 B.n707 B.n443 256.663
R1776 B.n707 B.n444 256.663
R1777 B.n707 B.n445 256.663
R1778 B.n707 B.n446 256.663
R1779 B.n817 B.n816 256.663
R1780 B.n104 B.n33 163.367
R1781 B.n108 B.n107 163.367
R1782 B.n112 B.n111 163.367
R1783 B.n116 B.n115 163.367
R1784 B.n120 B.n119 163.367
R1785 B.n124 B.n123 163.367
R1786 B.n128 B.n127 163.367
R1787 B.n132 B.n131 163.367
R1788 B.n136 B.n135 163.367
R1789 B.n140 B.n139 163.367
R1790 B.n144 B.n143 163.367
R1791 B.n148 B.n147 163.367
R1792 B.n152 B.n151 163.367
R1793 B.n156 B.n155 163.367
R1794 B.n160 B.n159 163.367
R1795 B.n164 B.n163 163.367
R1796 B.n168 B.n167 163.367
R1797 B.n172 B.n171 163.367
R1798 B.n176 B.n175 163.367
R1799 B.n180 B.n179 163.367
R1800 B.n184 B.n183 163.367
R1801 B.n188 B.n187 163.367
R1802 B.n192 B.n191 163.367
R1803 B.n196 B.n195 163.367
R1804 B.n200 B.n199 163.367
R1805 B.n204 B.n203 163.367
R1806 B.n208 B.n207 163.367
R1807 B.n212 B.n211 163.367
R1808 B.n216 B.n215 163.367
R1809 B.n220 B.n219 163.367
R1810 B.n224 B.n223 163.367
R1811 B.n228 B.n227 163.367
R1812 B.n232 B.n231 163.367
R1813 B.n236 B.n235 163.367
R1814 B.n241 B.n240 163.367
R1815 B.n245 B.n244 163.367
R1816 B.n249 B.n248 163.367
R1817 B.n253 B.n252 163.367
R1818 B.n257 B.n256 163.367
R1819 B.n261 B.n260 163.367
R1820 B.n265 B.n264 163.367
R1821 B.n269 B.n268 163.367
R1822 B.n273 B.n272 163.367
R1823 B.n277 B.n276 163.367
R1824 B.n281 B.n280 163.367
R1825 B.n285 B.n284 163.367
R1826 B.n289 B.n288 163.367
R1827 B.n293 B.n292 163.367
R1828 B.n297 B.n296 163.367
R1829 B.n301 B.n300 163.367
R1830 B.n305 B.n304 163.367
R1831 B.n309 B.n308 163.367
R1832 B.n313 B.n312 163.367
R1833 B.n317 B.n316 163.367
R1834 B.n321 B.n320 163.367
R1835 B.n325 B.n324 163.367
R1836 B.n329 B.n328 163.367
R1837 B.n333 B.n332 163.367
R1838 B.n337 B.n336 163.367
R1839 B.n341 B.n340 163.367
R1840 B.n345 B.n344 163.367
R1841 B.n349 B.n348 163.367
R1842 B.n353 B.n352 163.367
R1843 B.n779 B.n97 163.367
R1844 B.n715 B.n379 163.367
R1845 B.n715 B.n377 163.367
R1846 B.n719 B.n377 163.367
R1847 B.n719 B.n372 163.367
R1848 B.n728 B.n372 163.367
R1849 B.n728 B.n370 163.367
R1850 B.n732 B.n370 163.367
R1851 B.n732 B.n363 163.367
R1852 B.n740 B.n363 163.367
R1853 B.n740 B.n361 163.367
R1854 B.n745 B.n361 163.367
R1855 B.n745 B.n357 163.367
R1856 B.n754 B.n357 163.367
R1857 B.n755 B.n754 163.367
R1858 B.n755 B.n5 163.367
R1859 B.n6 B.n5 163.367
R1860 B.n7 B.n6 163.367
R1861 B.n761 B.n7 163.367
R1862 B.n762 B.n761 163.367
R1863 B.n762 B.n13 163.367
R1864 B.n14 B.n13 163.367
R1865 B.n15 B.n14 163.367
R1866 B.n767 B.n15 163.367
R1867 B.n767 B.n20 163.367
R1868 B.n21 B.n20 163.367
R1869 B.n22 B.n21 163.367
R1870 B.n772 B.n22 163.367
R1871 B.n772 B.n27 163.367
R1872 B.n28 B.n27 163.367
R1873 B.n29 B.n28 163.367
R1874 B.n98 B.n29 163.367
R1875 B.n706 B.n383 163.367
R1876 B.n706 B.n447 163.367
R1877 B.n702 B.n701 163.367
R1878 B.n698 B.n697 163.367
R1879 B.n694 B.n693 163.367
R1880 B.n690 B.n689 163.367
R1881 B.n686 B.n685 163.367
R1882 B.n682 B.n681 163.367
R1883 B.n678 B.n677 163.367
R1884 B.n674 B.n673 163.367
R1885 B.n670 B.n669 163.367
R1886 B.n666 B.n665 163.367
R1887 B.n662 B.n661 163.367
R1888 B.n658 B.n657 163.367
R1889 B.n654 B.n653 163.367
R1890 B.n650 B.n649 163.367
R1891 B.n646 B.n645 163.367
R1892 B.n642 B.n641 163.367
R1893 B.n638 B.n637 163.367
R1894 B.n634 B.n633 163.367
R1895 B.n630 B.n629 163.367
R1896 B.n626 B.n625 163.367
R1897 B.n622 B.n621 163.367
R1898 B.n618 B.n617 163.367
R1899 B.n614 B.n613 163.367
R1900 B.n610 B.n609 163.367
R1901 B.n606 B.n605 163.367
R1902 B.n602 B.n601 163.367
R1903 B.n598 B.n597 163.367
R1904 B.n594 B.n593 163.367
R1905 B.n589 B.n588 163.367
R1906 B.n585 B.n584 163.367
R1907 B.n581 B.n580 163.367
R1908 B.n577 B.n576 163.367
R1909 B.n573 B.n572 163.367
R1910 B.n569 B.n568 163.367
R1911 B.n565 B.n564 163.367
R1912 B.n561 B.n560 163.367
R1913 B.n557 B.n556 163.367
R1914 B.n553 B.n552 163.367
R1915 B.n549 B.n548 163.367
R1916 B.n545 B.n544 163.367
R1917 B.n541 B.n540 163.367
R1918 B.n537 B.n536 163.367
R1919 B.n533 B.n532 163.367
R1920 B.n529 B.n528 163.367
R1921 B.n525 B.n524 163.367
R1922 B.n521 B.n520 163.367
R1923 B.n517 B.n516 163.367
R1924 B.n513 B.n512 163.367
R1925 B.n509 B.n508 163.367
R1926 B.n505 B.n504 163.367
R1927 B.n501 B.n500 163.367
R1928 B.n497 B.n496 163.367
R1929 B.n493 B.n492 163.367
R1930 B.n489 B.n488 163.367
R1931 B.n485 B.n484 163.367
R1932 B.n481 B.n480 163.367
R1933 B.n477 B.n476 163.367
R1934 B.n473 B.n472 163.367
R1935 B.n469 B.n468 163.367
R1936 B.n465 B.n464 163.367
R1937 B.n461 B.n460 163.367
R1938 B.n457 B.n456 163.367
R1939 B.n713 B.n381 163.367
R1940 B.n713 B.n375 163.367
R1941 B.n722 B.n375 163.367
R1942 B.n722 B.n373 163.367
R1943 B.n726 B.n373 163.367
R1944 B.n726 B.n368 163.367
R1945 B.n734 B.n368 163.367
R1946 B.n734 B.n366 163.367
R1947 B.n738 B.n366 163.367
R1948 B.n738 B.n360 163.367
R1949 B.n748 B.n360 163.367
R1950 B.n748 B.n358 163.367
R1951 B.n752 B.n358 163.367
R1952 B.n752 B.n3 163.367
R1953 B.n815 B.n3 163.367
R1954 B.n811 B.n2 163.367
R1955 B.n811 B.n810 163.367
R1956 B.n810 B.n9 163.367
R1957 B.n806 B.n9 163.367
R1958 B.n806 B.n11 163.367
R1959 B.n802 B.n11 163.367
R1960 B.n802 B.n17 163.367
R1961 B.n798 B.n17 163.367
R1962 B.n798 B.n19 163.367
R1963 B.n794 B.n19 163.367
R1964 B.n794 B.n23 163.367
R1965 B.n790 B.n23 163.367
R1966 B.n790 B.n25 163.367
R1967 B.n786 B.n25 163.367
R1968 B.n786 B.n31 163.367
R1969 B.n782 B.n781 71.676
R1970 B.n104 B.n34 71.676
R1971 B.n108 B.n35 71.676
R1972 B.n112 B.n36 71.676
R1973 B.n116 B.n37 71.676
R1974 B.n120 B.n38 71.676
R1975 B.n124 B.n39 71.676
R1976 B.n128 B.n40 71.676
R1977 B.n132 B.n41 71.676
R1978 B.n136 B.n42 71.676
R1979 B.n140 B.n43 71.676
R1980 B.n144 B.n44 71.676
R1981 B.n148 B.n45 71.676
R1982 B.n152 B.n46 71.676
R1983 B.n156 B.n47 71.676
R1984 B.n160 B.n48 71.676
R1985 B.n164 B.n49 71.676
R1986 B.n168 B.n50 71.676
R1987 B.n172 B.n51 71.676
R1988 B.n176 B.n52 71.676
R1989 B.n180 B.n53 71.676
R1990 B.n184 B.n54 71.676
R1991 B.n188 B.n55 71.676
R1992 B.n192 B.n56 71.676
R1993 B.n196 B.n57 71.676
R1994 B.n200 B.n58 71.676
R1995 B.n204 B.n59 71.676
R1996 B.n208 B.n60 71.676
R1997 B.n212 B.n61 71.676
R1998 B.n216 B.n62 71.676
R1999 B.n220 B.n63 71.676
R2000 B.n224 B.n64 71.676
R2001 B.n228 B.n65 71.676
R2002 B.n232 B.n66 71.676
R2003 B.n236 B.n67 71.676
R2004 B.n241 B.n68 71.676
R2005 B.n245 B.n69 71.676
R2006 B.n249 B.n70 71.676
R2007 B.n253 B.n71 71.676
R2008 B.n257 B.n72 71.676
R2009 B.n261 B.n73 71.676
R2010 B.n265 B.n74 71.676
R2011 B.n269 B.n75 71.676
R2012 B.n273 B.n76 71.676
R2013 B.n277 B.n77 71.676
R2014 B.n281 B.n78 71.676
R2015 B.n285 B.n79 71.676
R2016 B.n289 B.n80 71.676
R2017 B.n293 B.n81 71.676
R2018 B.n297 B.n82 71.676
R2019 B.n301 B.n83 71.676
R2020 B.n305 B.n84 71.676
R2021 B.n309 B.n85 71.676
R2022 B.n313 B.n86 71.676
R2023 B.n317 B.n87 71.676
R2024 B.n321 B.n88 71.676
R2025 B.n325 B.n89 71.676
R2026 B.n329 B.n90 71.676
R2027 B.n333 B.n91 71.676
R2028 B.n337 B.n92 71.676
R2029 B.n341 B.n93 71.676
R2030 B.n345 B.n94 71.676
R2031 B.n349 B.n95 71.676
R2032 B.n353 B.n96 71.676
R2033 B.n97 B.n96 71.676
R2034 B.n352 B.n95 71.676
R2035 B.n348 B.n94 71.676
R2036 B.n344 B.n93 71.676
R2037 B.n340 B.n92 71.676
R2038 B.n336 B.n91 71.676
R2039 B.n332 B.n90 71.676
R2040 B.n328 B.n89 71.676
R2041 B.n324 B.n88 71.676
R2042 B.n320 B.n87 71.676
R2043 B.n316 B.n86 71.676
R2044 B.n312 B.n85 71.676
R2045 B.n308 B.n84 71.676
R2046 B.n304 B.n83 71.676
R2047 B.n300 B.n82 71.676
R2048 B.n296 B.n81 71.676
R2049 B.n292 B.n80 71.676
R2050 B.n288 B.n79 71.676
R2051 B.n284 B.n78 71.676
R2052 B.n280 B.n77 71.676
R2053 B.n276 B.n76 71.676
R2054 B.n272 B.n75 71.676
R2055 B.n268 B.n74 71.676
R2056 B.n264 B.n73 71.676
R2057 B.n260 B.n72 71.676
R2058 B.n256 B.n71 71.676
R2059 B.n252 B.n70 71.676
R2060 B.n248 B.n69 71.676
R2061 B.n244 B.n68 71.676
R2062 B.n240 B.n67 71.676
R2063 B.n235 B.n66 71.676
R2064 B.n231 B.n65 71.676
R2065 B.n227 B.n64 71.676
R2066 B.n223 B.n63 71.676
R2067 B.n219 B.n62 71.676
R2068 B.n215 B.n61 71.676
R2069 B.n211 B.n60 71.676
R2070 B.n207 B.n59 71.676
R2071 B.n203 B.n58 71.676
R2072 B.n199 B.n57 71.676
R2073 B.n195 B.n56 71.676
R2074 B.n191 B.n55 71.676
R2075 B.n187 B.n54 71.676
R2076 B.n183 B.n53 71.676
R2077 B.n179 B.n52 71.676
R2078 B.n175 B.n51 71.676
R2079 B.n171 B.n50 71.676
R2080 B.n167 B.n49 71.676
R2081 B.n163 B.n48 71.676
R2082 B.n159 B.n47 71.676
R2083 B.n155 B.n46 71.676
R2084 B.n151 B.n45 71.676
R2085 B.n147 B.n44 71.676
R2086 B.n143 B.n43 71.676
R2087 B.n139 B.n42 71.676
R2088 B.n135 B.n41 71.676
R2089 B.n131 B.n40 71.676
R2090 B.n127 B.n39 71.676
R2091 B.n123 B.n38 71.676
R2092 B.n119 B.n37 71.676
R2093 B.n115 B.n36 71.676
R2094 B.n111 B.n35 71.676
R2095 B.n107 B.n34 71.676
R2096 B.n781 B.n33 71.676
R2097 B.n709 B.n708 71.676
R2098 B.n447 B.n384 71.676
R2099 B.n701 B.n385 71.676
R2100 B.n697 B.n386 71.676
R2101 B.n693 B.n387 71.676
R2102 B.n689 B.n388 71.676
R2103 B.n685 B.n389 71.676
R2104 B.n681 B.n390 71.676
R2105 B.n677 B.n391 71.676
R2106 B.n673 B.n392 71.676
R2107 B.n669 B.n393 71.676
R2108 B.n665 B.n394 71.676
R2109 B.n661 B.n395 71.676
R2110 B.n657 B.n396 71.676
R2111 B.n653 B.n397 71.676
R2112 B.n649 B.n398 71.676
R2113 B.n645 B.n399 71.676
R2114 B.n641 B.n400 71.676
R2115 B.n637 B.n401 71.676
R2116 B.n633 B.n402 71.676
R2117 B.n629 B.n403 71.676
R2118 B.n625 B.n404 71.676
R2119 B.n621 B.n405 71.676
R2120 B.n617 B.n406 71.676
R2121 B.n613 B.n407 71.676
R2122 B.n609 B.n408 71.676
R2123 B.n605 B.n409 71.676
R2124 B.n601 B.n410 71.676
R2125 B.n597 B.n411 71.676
R2126 B.n593 B.n412 71.676
R2127 B.n588 B.n413 71.676
R2128 B.n584 B.n414 71.676
R2129 B.n580 B.n415 71.676
R2130 B.n576 B.n416 71.676
R2131 B.n572 B.n417 71.676
R2132 B.n568 B.n418 71.676
R2133 B.n564 B.n419 71.676
R2134 B.n560 B.n420 71.676
R2135 B.n556 B.n421 71.676
R2136 B.n552 B.n422 71.676
R2137 B.n548 B.n423 71.676
R2138 B.n544 B.n424 71.676
R2139 B.n540 B.n425 71.676
R2140 B.n536 B.n426 71.676
R2141 B.n532 B.n427 71.676
R2142 B.n528 B.n428 71.676
R2143 B.n524 B.n429 71.676
R2144 B.n520 B.n430 71.676
R2145 B.n516 B.n431 71.676
R2146 B.n512 B.n432 71.676
R2147 B.n508 B.n433 71.676
R2148 B.n504 B.n434 71.676
R2149 B.n500 B.n435 71.676
R2150 B.n496 B.n436 71.676
R2151 B.n492 B.n437 71.676
R2152 B.n488 B.n438 71.676
R2153 B.n484 B.n439 71.676
R2154 B.n480 B.n440 71.676
R2155 B.n476 B.n441 71.676
R2156 B.n472 B.n442 71.676
R2157 B.n468 B.n443 71.676
R2158 B.n464 B.n444 71.676
R2159 B.n460 B.n445 71.676
R2160 B.n456 B.n446 71.676
R2161 B.n708 B.n383 71.676
R2162 B.n702 B.n384 71.676
R2163 B.n698 B.n385 71.676
R2164 B.n694 B.n386 71.676
R2165 B.n690 B.n387 71.676
R2166 B.n686 B.n388 71.676
R2167 B.n682 B.n389 71.676
R2168 B.n678 B.n390 71.676
R2169 B.n674 B.n391 71.676
R2170 B.n670 B.n392 71.676
R2171 B.n666 B.n393 71.676
R2172 B.n662 B.n394 71.676
R2173 B.n658 B.n395 71.676
R2174 B.n654 B.n396 71.676
R2175 B.n650 B.n397 71.676
R2176 B.n646 B.n398 71.676
R2177 B.n642 B.n399 71.676
R2178 B.n638 B.n400 71.676
R2179 B.n634 B.n401 71.676
R2180 B.n630 B.n402 71.676
R2181 B.n626 B.n403 71.676
R2182 B.n622 B.n404 71.676
R2183 B.n618 B.n405 71.676
R2184 B.n614 B.n406 71.676
R2185 B.n610 B.n407 71.676
R2186 B.n606 B.n408 71.676
R2187 B.n602 B.n409 71.676
R2188 B.n598 B.n410 71.676
R2189 B.n594 B.n411 71.676
R2190 B.n589 B.n412 71.676
R2191 B.n585 B.n413 71.676
R2192 B.n581 B.n414 71.676
R2193 B.n577 B.n415 71.676
R2194 B.n573 B.n416 71.676
R2195 B.n569 B.n417 71.676
R2196 B.n565 B.n418 71.676
R2197 B.n561 B.n419 71.676
R2198 B.n557 B.n420 71.676
R2199 B.n553 B.n421 71.676
R2200 B.n549 B.n422 71.676
R2201 B.n545 B.n423 71.676
R2202 B.n541 B.n424 71.676
R2203 B.n537 B.n425 71.676
R2204 B.n533 B.n426 71.676
R2205 B.n529 B.n427 71.676
R2206 B.n525 B.n428 71.676
R2207 B.n521 B.n429 71.676
R2208 B.n517 B.n430 71.676
R2209 B.n513 B.n431 71.676
R2210 B.n509 B.n432 71.676
R2211 B.n505 B.n433 71.676
R2212 B.n501 B.n434 71.676
R2213 B.n497 B.n435 71.676
R2214 B.n493 B.n436 71.676
R2215 B.n489 B.n437 71.676
R2216 B.n485 B.n438 71.676
R2217 B.n481 B.n439 71.676
R2218 B.n477 B.n440 71.676
R2219 B.n473 B.n441 71.676
R2220 B.n469 B.n442 71.676
R2221 B.n465 B.n443 71.676
R2222 B.n461 B.n444 71.676
R2223 B.n457 B.n445 71.676
R2224 B.n453 B.n446 71.676
R2225 B.n816 B.n815 71.676
R2226 B.n816 B.n2 71.676
R2227 B.n707 B.n380 61.5422
R2228 B.n780 B.n30 61.5422
R2229 B.n103 B.n102 59.5399
R2230 B.n238 B.n100 59.5399
R2231 B.n452 B.n451 59.5399
R2232 B.n591 B.n449 59.5399
R2233 B.n711 B.n710 33.2493
R2234 B.n454 B.n378 33.2493
R2235 B.n778 B.n777 33.2493
R2236 B.n784 B.n783 33.2493
R2237 B.n714 B.n380 31.9458
R2238 B.n714 B.n376 31.9458
R2239 B.n721 B.n376 31.9458
R2240 B.n721 B.n720 31.9458
R2241 B.n727 B.n369 31.9458
R2242 B.n733 B.n369 31.9458
R2243 B.n733 B.n364 31.9458
R2244 B.n739 B.n364 31.9458
R2245 B.n739 B.n365 31.9458
R2246 B.n747 B.n746 31.9458
R2247 B.n753 B.n4 31.9458
R2248 B.n814 B.n4 31.9458
R2249 B.n814 B.n813 31.9458
R2250 B.n813 B.n812 31.9458
R2251 B.n812 B.n8 31.9458
R2252 B.n805 B.n12 31.9458
R2253 B.n804 B.n803 31.9458
R2254 B.n803 B.n16 31.9458
R2255 B.n797 B.n16 31.9458
R2256 B.n797 B.n796 31.9458
R2257 B.n796 B.n795 31.9458
R2258 B.n789 B.n26 31.9458
R2259 B.n789 B.n788 31.9458
R2260 B.n788 B.n787 31.9458
R2261 B.n787 B.n30 31.9458
R2262 B.n747 B.t2 27.248
R2263 B.n805 B.t1 27.248
R2264 B.n746 B.t0 20.671
R2265 B.n12 B.t3 20.671
R2266 B B.n817 18.0485
R2267 B.n727 B.t9 17.8523
R2268 B.n795 B.t5 17.8523
R2269 B.n102 B.n101 16.4853
R2270 B.n100 B.n99 16.4853
R2271 B.n451 B.n450 16.4853
R2272 B.n449 B.n448 16.4853
R2273 B.n720 B.t9 14.094
R2274 B.n26 B.t5 14.094
R2275 B.n753 B.t0 11.2753
R2276 B.t3 B.n8 11.2753
R2277 B.n712 B.n711 10.6151
R2278 B.n712 B.n374 10.6151
R2279 B.n723 B.n374 10.6151
R2280 B.n724 B.n723 10.6151
R2281 B.n725 B.n724 10.6151
R2282 B.n725 B.n367 10.6151
R2283 B.n735 B.n367 10.6151
R2284 B.n736 B.n735 10.6151
R2285 B.n737 B.n736 10.6151
R2286 B.n737 B.n359 10.6151
R2287 B.n749 B.n359 10.6151
R2288 B.n750 B.n749 10.6151
R2289 B.n751 B.n750 10.6151
R2290 B.n751 B.n0 10.6151
R2291 B.n710 B.n382 10.6151
R2292 B.n705 B.n382 10.6151
R2293 B.n705 B.n704 10.6151
R2294 B.n704 B.n703 10.6151
R2295 B.n703 B.n700 10.6151
R2296 B.n700 B.n699 10.6151
R2297 B.n699 B.n696 10.6151
R2298 B.n696 B.n695 10.6151
R2299 B.n695 B.n692 10.6151
R2300 B.n692 B.n691 10.6151
R2301 B.n691 B.n688 10.6151
R2302 B.n688 B.n687 10.6151
R2303 B.n687 B.n684 10.6151
R2304 B.n684 B.n683 10.6151
R2305 B.n683 B.n680 10.6151
R2306 B.n680 B.n679 10.6151
R2307 B.n679 B.n676 10.6151
R2308 B.n676 B.n675 10.6151
R2309 B.n675 B.n672 10.6151
R2310 B.n672 B.n671 10.6151
R2311 B.n671 B.n668 10.6151
R2312 B.n668 B.n667 10.6151
R2313 B.n667 B.n664 10.6151
R2314 B.n664 B.n663 10.6151
R2315 B.n663 B.n660 10.6151
R2316 B.n660 B.n659 10.6151
R2317 B.n659 B.n656 10.6151
R2318 B.n656 B.n655 10.6151
R2319 B.n655 B.n652 10.6151
R2320 B.n652 B.n651 10.6151
R2321 B.n651 B.n648 10.6151
R2322 B.n648 B.n647 10.6151
R2323 B.n647 B.n644 10.6151
R2324 B.n644 B.n643 10.6151
R2325 B.n643 B.n640 10.6151
R2326 B.n640 B.n639 10.6151
R2327 B.n639 B.n636 10.6151
R2328 B.n636 B.n635 10.6151
R2329 B.n635 B.n632 10.6151
R2330 B.n632 B.n631 10.6151
R2331 B.n631 B.n628 10.6151
R2332 B.n628 B.n627 10.6151
R2333 B.n627 B.n624 10.6151
R2334 B.n624 B.n623 10.6151
R2335 B.n623 B.n620 10.6151
R2336 B.n620 B.n619 10.6151
R2337 B.n619 B.n616 10.6151
R2338 B.n616 B.n615 10.6151
R2339 B.n615 B.n612 10.6151
R2340 B.n612 B.n611 10.6151
R2341 B.n611 B.n608 10.6151
R2342 B.n608 B.n607 10.6151
R2343 B.n607 B.n604 10.6151
R2344 B.n604 B.n603 10.6151
R2345 B.n603 B.n600 10.6151
R2346 B.n600 B.n599 10.6151
R2347 B.n599 B.n596 10.6151
R2348 B.n596 B.n595 10.6151
R2349 B.n595 B.n592 10.6151
R2350 B.n590 B.n587 10.6151
R2351 B.n587 B.n586 10.6151
R2352 B.n586 B.n583 10.6151
R2353 B.n583 B.n582 10.6151
R2354 B.n582 B.n579 10.6151
R2355 B.n579 B.n578 10.6151
R2356 B.n578 B.n575 10.6151
R2357 B.n575 B.n574 10.6151
R2358 B.n571 B.n570 10.6151
R2359 B.n570 B.n567 10.6151
R2360 B.n567 B.n566 10.6151
R2361 B.n566 B.n563 10.6151
R2362 B.n563 B.n562 10.6151
R2363 B.n562 B.n559 10.6151
R2364 B.n559 B.n558 10.6151
R2365 B.n558 B.n555 10.6151
R2366 B.n555 B.n554 10.6151
R2367 B.n554 B.n551 10.6151
R2368 B.n551 B.n550 10.6151
R2369 B.n550 B.n547 10.6151
R2370 B.n547 B.n546 10.6151
R2371 B.n546 B.n543 10.6151
R2372 B.n543 B.n542 10.6151
R2373 B.n542 B.n539 10.6151
R2374 B.n539 B.n538 10.6151
R2375 B.n538 B.n535 10.6151
R2376 B.n535 B.n534 10.6151
R2377 B.n534 B.n531 10.6151
R2378 B.n531 B.n530 10.6151
R2379 B.n530 B.n527 10.6151
R2380 B.n527 B.n526 10.6151
R2381 B.n526 B.n523 10.6151
R2382 B.n523 B.n522 10.6151
R2383 B.n522 B.n519 10.6151
R2384 B.n519 B.n518 10.6151
R2385 B.n518 B.n515 10.6151
R2386 B.n515 B.n514 10.6151
R2387 B.n514 B.n511 10.6151
R2388 B.n511 B.n510 10.6151
R2389 B.n510 B.n507 10.6151
R2390 B.n507 B.n506 10.6151
R2391 B.n506 B.n503 10.6151
R2392 B.n503 B.n502 10.6151
R2393 B.n502 B.n499 10.6151
R2394 B.n499 B.n498 10.6151
R2395 B.n498 B.n495 10.6151
R2396 B.n495 B.n494 10.6151
R2397 B.n494 B.n491 10.6151
R2398 B.n491 B.n490 10.6151
R2399 B.n490 B.n487 10.6151
R2400 B.n487 B.n486 10.6151
R2401 B.n486 B.n483 10.6151
R2402 B.n483 B.n482 10.6151
R2403 B.n482 B.n479 10.6151
R2404 B.n479 B.n478 10.6151
R2405 B.n478 B.n475 10.6151
R2406 B.n475 B.n474 10.6151
R2407 B.n474 B.n471 10.6151
R2408 B.n471 B.n470 10.6151
R2409 B.n470 B.n467 10.6151
R2410 B.n467 B.n466 10.6151
R2411 B.n466 B.n463 10.6151
R2412 B.n463 B.n462 10.6151
R2413 B.n462 B.n459 10.6151
R2414 B.n459 B.n458 10.6151
R2415 B.n458 B.n455 10.6151
R2416 B.n455 B.n454 10.6151
R2417 B.n716 B.n378 10.6151
R2418 B.n717 B.n716 10.6151
R2419 B.n718 B.n717 10.6151
R2420 B.n718 B.n371 10.6151
R2421 B.n729 B.n371 10.6151
R2422 B.n730 B.n729 10.6151
R2423 B.n731 B.n730 10.6151
R2424 B.n731 B.n362 10.6151
R2425 B.n741 B.n362 10.6151
R2426 B.n742 B.n741 10.6151
R2427 B.n744 B.n742 10.6151
R2428 B.n744 B.n743 10.6151
R2429 B.n743 B.n356 10.6151
R2430 B.n756 B.n356 10.6151
R2431 B.n757 B.n756 10.6151
R2432 B.n758 B.n757 10.6151
R2433 B.n759 B.n758 10.6151
R2434 B.n760 B.n759 10.6151
R2435 B.n763 B.n760 10.6151
R2436 B.n764 B.n763 10.6151
R2437 B.n765 B.n764 10.6151
R2438 B.n766 B.n765 10.6151
R2439 B.n768 B.n766 10.6151
R2440 B.n769 B.n768 10.6151
R2441 B.n770 B.n769 10.6151
R2442 B.n771 B.n770 10.6151
R2443 B.n773 B.n771 10.6151
R2444 B.n774 B.n773 10.6151
R2445 B.n775 B.n774 10.6151
R2446 B.n776 B.n775 10.6151
R2447 B.n777 B.n776 10.6151
R2448 B.n809 B.n1 10.6151
R2449 B.n809 B.n808 10.6151
R2450 B.n808 B.n807 10.6151
R2451 B.n807 B.n10 10.6151
R2452 B.n801 B.n10 10.6151
R2453 B.n801 B.n800 10.6151
R2454 B.n800 B.n799 10.6151
R2455 B.n799 B.n18 10.6151
R2456 B.n793 B.n18 10.6151
R2457 B.n793 B.n792 10.6151
R2458 B.n792 B.n791 10.6151
R2459 B.n791 B.n24 10.6151
R2460 B.n785 B.n24 10.6151
R2461 B.n785 B.n784 10.6151
R2462 B.n783 B.n32 10.6151
R2463 B.n105 B.n32 10.6151
R2464 B.n106 B.n105 10.6151
R2465 B.n109 B.n106 10.6151
R2466 B.n110 B.n109 10.6151
R2467 B.n113 B.n110 10.6151
R2468 B.n114 B.n113 10.6151
R2469 B.n117 B.n114 10.6151
R2470 B.n118 B.n117 10.6151
R2471 B.n121 B.n118 10.6151
R2472 B.n122 B.n121 10.6151
R2473 B.n125 B.n122 10.6151
R2474 B.n126 B.n125 10.6151
R2475 B.n129 B.n126 10.6151
R2476 B.n130 B.n129 10.6151
R2477 B.n133 B.n130 10.6151
R2478 B.n134 B.n133 10.6151
R2479 B.n137 B.n134 10.6151
R2480 B.n138 B.n137 10.6151
R2481 B.n141 B.n138 10.6151
R2482 B.n142 B.n141 10.6151
R2483 B.n145 B.n142 10.6151
R2484 B.n146 B.n145 10.6151
R2485 B.n149 B.n146 10.6151
R2486 B.n150 B.n149 10.6151
R2487 B.n153 B.n150 10.6151
R2488 B.n154 B.n153 10.6151
R2489 B.n157 B.n154 10.6151
R2490 B.n158 B.n157 10.6151
R2491 B.n161 B.n158 10.6151
R2492 B.n162 B.n161 10.6151
R2493 B.n165 B.n162 10.6151
R2494 B.n166 B.n165 10.6151
R2495 B.n169 B.n166 10.6151
R2496 B.n170 B.n169 10.6151
R2497 B.n173 B.n170 10.6151
R2498 B.n174 B.n173 10.6151
R2499 B.n177 B.n174 10.6151
R2500 B.n178 B.n177 10.6151
R2501 B.n181 B.n178 10.6151
R2502 B.n182 B.n181 10.6151
R2503 B.n185 B.n182 10.6151
R2504 B.n186 B.n185 10.6151
R2505 B.n189 B.n186 10.6151
R2506 B.n190 B.n189 10.6151
R2507 B.n193 B.n190 10.6151
R2508 B.n194 B.n193 10.6151
R2509 B.n197 B.n194 10.6151
R2510 B.n198 B.n197 10.6151
R2511 B.n201 B.n198 10.6151
R2512 B.n202 B.n201 10.6151
R2513 B.n205 B.n202 10.6151
R2514 B.n206 B.n205 10.6151
R2515 B.n209 B.n206 10.6151
R2516 B.n210 B.n209 10.6151
R2517 B.n213 B.n210 10.6151
R2518 B.n214 B.n213 10.6151
R2519 B.n217 B.n214 10.6151
R2520 B.n218 B.n217 10.6151
R2521 B.n222 B.n221 10.6151
R2522 B.n225 B.n222 10.6151
R2523 B.n226 B.n225 10.6151
R2524 B.n229 B.n226 10.6151
R2525 B.n230 B.n229 10.6151
R2526 B.n233 B.n230 10.6151
R2527 B.n234 B.n233 10.6151
R2528 B.n237 B.n234 10.6151
R2529 B.n242 B.n239 10.6151
R2530 B.n243 B.n242 10.6151
R2531 B.n246 B.n243 10.6151
R2532 B.n247 B.n246 10.6151
R2533 B.n250 B.n247 10.6151
R2534 B.n251 B.n250 10.6151
R2535 B.n254 B.n251 10.6151
R2536 B.n255 B.n254 10.6151
R2537 B.n258 B.n255 10.6151
R2538 B.n259 B.n258 10.6151
R2539 B.n262 B.n259 10.6151
R2540 B.n263 B.n262 10.6151
R2541 B.n266 B.n263 10.6151
R2542 B.n267 B.n266 10.6151
R2543 B.n270 B.n267 10.6151
R2544 B.n271 B.n270 10.6151
R2545 B.n274 B.n271 10.6151
R2546 B.n275 B.n274 10.6151
R2547 B.n278 B.n275 10.6151
R2548 B.n279 B.n278 10.6151
R2549 B.n282 B.n279 10.6151
R2550 B.n283 B.n282 10.6151
R2551 B.n286 B.n283 10.6151
R2552 B.n287 B.n286 10.6151
R2553 B.n290 B.n287 10.6151
R2554 B.n291 B.n290 10.6151
R2555 B.n294 B.n291 10.6151
R2556 B.n295 B.n294 10.6151
R2557 B.n298 B.n295 10.6151
R2558 B.n299 B.n298 10.6151
R2559 B.n302 B.n299 10.6151
R2560 B.n303 B.n302 10.6151
R2561 B.n306 B.n303 10.6151
R2562 B.n307 B.n306 10.6151
R2563 B.n310 B.n307 10.6151
R2564 B.n311 B.n310 10.6151
R2565 B.n314 B.n311 10.6151
R2566 B.n315 B.n314 10.6151
R2567 B.n318 B.n315 10.6151
R2568 B.n319 B.n318 10.6151
R2569 B.n322 B.n319 10.6151
R2570 B.n323 B.n322 10.6151
R2571 B.n326 B.n323 10.6151
R2572 B.n327 B.n326 10.6151
R2573 B.n330 B.n327 10.6151
R2574 B.n331 B.n330 10.6151
R2575 B.n334 B.n331 10.6151
R2576 B.n335 B.n334 10.6151
R2577 B.n338 B.n335 10.6151
R2578 B.n339 B.n338 10.6151
R2579 B.n342 B.n339 10.6151
R2580 B.n343 B.n342 10.6151
R2581 B.n346 B.n343 10.6151
R2582 B.n347 B.n346 10.6151
R2583 B.n350 B.n347 10.6151
R2584 B.n351 B.n350 10.6151
R2585 B.n354 B.n351 10.6151
R2586 B.n355 B.n354 10.6151
R2587 B.n778 B.n355 10.6151
R2588 B.n817 B.n0 8.11757
R2589 B.n817 B.n1 8.11757
R2590 B.n591 B.n590 6.5566
R2591 B.n574 B.n452 6.5566
R2592 B.n221 B.n103 6.5566
R2593 B.n238 B.n237 6.5566
R2594 B.n365 B.t2 4.69834
R2595 B.t1 B.n804 4.69834
R2596 B.n592 B.n591 4.05904
R2597 B.n571 B.n452 4.05904
R2598 B.n218 B.n103 4.05904
R2599 B.n239 B.n238 4.05904
R2600 VN.n0 VN.t0 937.245
R2601 VN.n1 VN.t1 937.245
R2602 VN.n0 VN.t3 937.221
R2603 VN.n1 VN.t2 937.221
R2604 VN VN.n1 115.162
R2605 VN VN.n0 70.265
R2606 VDD2.n2 VDD2.n0 100.26
R2607 VDD2.n2 VDD2.n1 58.7087
R2608 VDD2.n1 VDD2.t1 1.09201
R2609 VDD2.n1 VDD2.t2 1.09201
R2610 VDD2.n0 VDD2.t3 1.09201
R2611 VDD2.n0 VDD2.t0 1.09201
R2612 VDD2 VDD2.n2 0.0586897
C0 VDD1 VP 4.11947f
C1 VP VTAIL 3.32114f
C2 VDD2 VP 0.262389f
C3 VDD1 VTAIL 10.77f
C4 VDD1 VDD2 0.527935f
C5 VP VN 5.82666f
C6 VDD2 VTAIL 10.8103f
C7 VDD1 VN 0.147558f
C8 VN VTAIL 3.30703f
C9 VDD2 VN 4.00485f
C10 VDD2 B 3.08326f
C11 VDD1 B 7.661f
C12 VTAIL B 12.104782f
C13 VN B 9.1596f
C14 VP B 4.928979f
C15 VDD2.t3 B 0.426473f
C16 VDD2.t0 B 0.426473f
C17 VDD2.n0 B 4.77933f
C18 VDD2.t1 B 0.426473f
C19 VDD2.t2 B 0.426473f
C20 VDD2.n1 B 3.88275f
C21 VDD2.n2 B 4.35538f
C22 VN.t0 B 1.45264f
C23 VN.t3 B 1.45263f
C24 VN.n0 B 1.06925f
C25 VN.t1 B 1.45264f
C26 VN.t2 B 1.45263f
C27 VN.n1 B 2.06491f
C28 VDD1.t1 B 0.42619f
C29 VDD1.t3 B 0.42619f
C30 VDD1.n0 B 3.88051f
C31 VDD1.t0 B 0.42619f
C32 VDD1.t2 B 0.42619f
C33 VDD1.n1 B 4.80763f
C34 VTAIL.n0 B 0.022149f
C35 VTAIL.n1 B 0.016552f
C36 VTAIL.n2 B 0.008894f
C37 VTAIL.n3 B 0.021023f
C38 VTAIL.n4 B 0.009418f
C39 VTAIL.n5 B 0.016552f
C40 VTAIL.n6 B 0.008894f
C41 VTAIL.n7 B 0.021023f
C42 VTAIL.n8 B 0.009418f
C43 VTAIL.n9 B 0.016552f
C44 VTAIL.n10 B 0.009156f
C45 VTAIL.n11 B 0.021023f
C46 VTAIL.n12 B 0.009418f
C47 VTAIL.n13 B 0.016552f
C48 VTAIL.n14 B 0.008894f
C49 VTAIL.n15 B 0.021023f
C50 VTAIL.n16 B 0.009418f
C51 VTAIL.n17 B 0.016552f
C52 VTAIL.n18 B 0.008894f
C53 VTAIL.n19 B 0.021023f
C54 VTAIL.n20 B 0.009418f
C55 VTAIL.n21 B 0.016552f
C56 VTAIL.n22 B 0.008894f
C57 VTAIL.n23 B 0.021023f
C58 VTAIL.n24 B 0.009418f
C59 VTAIL.n25 B 0.016552f
C60 VTAIL.n26 B 0.008894f
C61 VTAIL.n27 B 0.021023f
C62 VTAIL.n28 B 0.009418f
C63 VTAIL.n29 B 0.016552f
C64 VTAIL.n30 B 0.008894f
C65 VTAIL.n31 B 0.015767f
C66 VTAIL.n32 B 0.012419f
C67 VTAIL.t3 B 0.034843f
C68 VTAIL.n33 B 0.120988f
C69 VTAIL.n34 B 1.31511f
C70 VTAIL.n35 B 0.008894f
C71 VTAIL.n36 B 0.009418f
C72 VTAIL.n37 B 0.021023f
C73 VTAIL.n38 B 0.021023f
C74 VTAIL.n39 B 0.009418f
C75 VTAIL.n40 B 0.008894f
C76 VTAIL.n41 B 0.016552f
C77 VTAIL.n42 B 0.016552f
C78 VTAIL.n43 B 0.008894f
C79 VTAIL.n44 B 0.009418f
C80 VTAIL.n45 B 0.021023f
C81 VTAIL.n46 B 0.021023f
C82 VTAIL.n47 B 0.009418f
C83 VTAIL.n48 B 0.008894f
C84 VTAIL.n49 B 0.016552f
C85 VTAIL.n50 B 0.016552f
C86 VTAIL.n51 B 0.008894f
C87 VTAIL.n52 B 0.009418f
C88 VTAIL.n53 B 0.021023f
C89 VTAIL.n54 B 0.021023f
C90 VTAIL.n55 B 0.009418f
C91 VTAIL.n56 B 0.008894f
C92 VTAIL.n57 B 0.016552f
C93 VTAIL.n58 B 0.016552f
C94 VTAIL.n59 B 0.008894f
C95 VTAIL.n60 B 0.009418f
C96 VTAIL.n61 B 0.021023f
C97 VTAIL.n62 B 0.021023f
C98 VTAIL.n63 B 0.009418f
C99 VTAIL.n64 B 0.008894f
C100 VTAIL.n65 B 0.016552f
C101 VTAIL.n66 B 0.016552f
C102 VTAIL.n67 B 0.008894f
C103 VTAIL.n68 B 0.009418f
C104 VTAIL.n69 B 0.021023f
C105 VTAIL.n70 B 0.021023f
C106 VTAIL.n71 B 0.009418f
C107 VTAIL.n72 B 0.008894f
C108 VTAIL.n73 B 0.016552f
C109 VTAIL.n74 B 0.016552f
C110 VTAIL.n75 B 0.008894f
C111 VTAIL.n76 B 0.008894f
C112 VTAIL.n77 B 0.009418f
C113 VTAIL.n78 B 0.021023f
C114 VTAIL.n79 B 0.021023f
C115 VTAIL.n80 B 0.021023f
C116 VTAIL.n81 B 0.009156f
C117 VTAIL.n82 B 0.008894f
C118 VTAIL.n83 B 0.016552f
C119 VTAIL.n84 B 0.016552f
C120 VTAIL.n85 B 0.008894f
C121 VTAIL.n86 B 0.009418f
C122 VTAIL.n87 B 0.021023f
C123 VTAIL.n88 B 0.021023f
C124 VTAIL.n89 B 0.009418f
C125 VTAIL.n90 B 0.008894f
C126 VTAIL.n91 B 0.016552f
C127 VTAIL.n92 B 0.016552f
C128 VTAIL.n93 B 0.008894f
C129 VTAIL.n94 B 0.009418f
C130 VTAIL.n95 B 0.021023f
C131 VTAIL.n96 B 0.043537f
C132 VTAIL.n97 B 0.009418f
C133 VTAIL.n98 B 0.008894f
C134 VTAIL.n99 B 0.035998f
C135 VTAIL.n100 B 0.024086f
C136 VTAIL.n101 B 0.060565f
C137 VTAIL.n102 B 0.022149f
C138 VTAIL.n103 B 0.016552f
C139 VTAIL.n104 B 0.008894f
C140 VTAIL.n105 B 0.021023f
C141 VTAIL.n106 B 0.009418f
C142 VTAIL.n107 B 0.016552f
C143 VTAIL.n108 B 0.008894f
C144 VTAIL.n109 B 0.021023f
C145 VTAIL.n110 B 0.009418f
C146 VTAIL.n111 B 0.016552f
C147 VTAIL.n112 B 0.009156f
C148 VTAIL.n113 B 0.021023f
C149 VTAIL.n114 B 0.009418f
C150 VTAIL.n115 B 0.016552f
C151 VTAIL.n116 B 0.008894f
C152 VTAIL.n117 B 0.021023f
C153 VTAIL.n118 B 0.009418f
C154 VTAIL.n119 B 0.016552f
C155 VTAIL.n120 B 0.008894f
C156 VTAIL.n121 B 0.021023f
C157 VTAIL.n122 B 0.009418f
C158 VTAIL.n123 B 0.016552f
C159 VTAIL.n124 B 0.008894f
C160 VTAIL.n125 B 0.021023f
C161 VTAIL.n126 B 0.009418f
C162 VTAIL.n127 B 0.016552f
C163 VTAIL.n128 B 0.008894f
C164 VTAIL.n129 B 0.021023f
C165 VTAIL.n130 B 0.009418f
C166 VTAIL.n131 B 0.016552f
C167 VTAIL.n132 B 0.008894f
C168 VTAIL.n133 B 0.015767f
C169 VTAIL.n134 B 0.012419f
C170 VTAIL.t7 B 0.034843f
C171 VTAIL.n135 B 0.120988f
C172 VTAIL.n136 B 1.31511f
C173 VTAIL.n137 B 0.008894f
C174 VTAIL.n138 B 0.009418f
C175 VTAIL.n139 B 0.021023f
C176 VTAIL.n140 B 0.021023f
C177 VTAIL.n141 B 0.009418f
C178 VTAIL.n142 B 0.008894f
C179 VTAIL.n143 B 0.016552f
C180 VTAIL.n144 B 0.016552f
C181 VTAIL.n145 B 0.008894f
C182 VTAIL.n146 B 0.009418f
C183 VTAIL.n147 B 0.021023f
C184 VTAIL.n148 B 0.021023f
C185 VTAIL.n149 B 0.009418f
C186 VTAIL.n150 B 0.008894f
C187 VTAIL.n151 B 0.016552f
C188 VTAIL.n152 B 0.016552f
C189 VTAIL.n153 B 0.008894f
C190 VTAIL.n154 B 0.009418f
C191 VTAIL.n155 B 0.021023f
C192 VTAIL.n156 B 0.021023f
C193 VTAIL.n157 B 0.009418f
C194 VTAIL.n158 B 0.008894f
C195 VTAIL.n159 B 0.016552f
C196 VTAIL.n160 B 0.016552f
C197 VTAIL.n161 B 0.008894f
C198 VTAIL.n162 B 0.009418f
C199 VTAIL.n163 B 0.021023f
C200 VTAIL.n164 B 0.021023f
C201 VTAIL.n165 B 0.009418f
C202 VTAIL.n166 B 0.008894f
C203 VTAIL.n167 B 0.016552f
C204 VTAIL.n168 B 0.016552f
C205 VTAIL.n169 B 0.008894f
C206 VTAIL.n170 B 0.009418f
C207 VTAIL.n171 B 0.021023f
C208 VTAIL.n172 B 0.021023f
C209 VTAIL.n173 B 0.009418f
C210 VTAIL.n174 B 0.008894f
C211 VTAIL.n175 B 0.016552f
C212 VTAIL.n176 B 0.016552f
C213 VTAIL.n177 B 0.008894f
C214 VTAIL.n178 B 0.008894f
C215 VTAIL.n179 B 0.009418f
C216 VTAIL.n180 B 0.021023f
C217 VTAIL.n181 B 0.021023f
C218 VTAIL.n182 B 0.021023f
C219 VTAIL.n183 B 0.009156f
C220 VTAIL.n184 B 0.008894f
C221 VTAIL.n185 B 0.016552f
C222 VTAIL.n186 B 0.016552f
C223 VTAIL.n187 B 0.008894f
C224 VTAIL.n188 B 0.009418f
C225 VTAIL.n189 B 0.021023f
C226 VTAIL.n190 B 0.021023f
C227 VTAIL.n191 B 0.009418f
C228 VTAIL.n192 B 0.008894f
C229 VTAIL.n193 B 0.016552f
C230 VTAIL.n194 B 0.016552f
C231 VTAIL.n195 B 0.008894f
C232 VTAIL.n196 B 0.009418f
C233 VTAIL.n197 B 0.021023f
C234 VTAIL.n198 B 0.043537f
C235 VTAIL.n199 B 0.009418f
C236 VTAIL.n200 B 0.008894f
C237 VTAIL.n201 B 0.035998f
C238 VTAIL.n202 B 0.024086f
C239 VTAIL.n203 B 0.077002f
C240 VTAIL.n204 B 0.022149f
C241 VTAIL.n205 B 0.016552f
C242 VTAIL.n206 B 0.008894f
C243 VTAIL.n207 B 0.021023f
C244 VTAIL.n208 B 0.009418f
C245 VTAIL.n209 B 0.016552f
C246 VTAIL.n210 B 0.008894f
C247 VTAIL.n211 B 0.021023f
C248 VTAIL.n212 B 0.009418f
C249 VTAIL.n213 B 0.016552f
C250 VTAIL.n214 B 0.009156f
C251 VTAIL.n215 B 0.021023f
C252 VTAIL.n216 B 0.009418f
C253 VTAIL.n217 B 0.016552f
C254 VTAIL.n218 B 0.008894f
C255 VTAIL.n219 B 0.021023f
C256 VTAIL.n220 B 0.009418f
C257 VTAIL.n221 B 0.016552f
C258 VTAIL.n222 B 0.008894f
C259 VTAIL.n223 B 0.021023f
C260 VTAIL.n224 B 0.009418f
C261 VTAIL.n225 B 0.016552f
C262 VTAIL.n226 B 0.008894f
C263 VTAIL.n227 B 0.021023f
C264 VTAIL.n228 B 0.009418f
C265 VTAIL.n229 B 0.016552f
C266 VTAIL.n230 B 0.008894f
C267 VTAIL.n231 B 0.021023f
C268 VTAIL.n232 B 0.009418f
C269 VTAIL.n233 B 0.016552f
C270 VTAIL.n234 B 0.008894f
C271 VTAIL.n235 B 0.015767f
C272 VTAIL.n236 B 0.012419f
C273 VTAIL.t5 B 0.034843f
C274 VTAIL.n237 B 0.120988f
C275 VTAIL.n238 B 1.31511f
C276 VTAIL.n239 B 0.008894f
C277 VTAIL.n240 B 0.009418f
C278 VTAIL.n241 B 0.021023f
C279 VTAIL.n242 B 0.021023f
C280 VTAIL.n243 B 0.009418f
C281 VTAIL.n244 B 0.008894f
C282 VTAIL.n245 B 0.016552f
C283 VTAIL.n246 B 0.016552f
C284 VTAIL.n247 B 0.008894f
C285 VTAIL.n248 B 0.009418f
C286 VTAIL.n249 B 0.021023f
C287 VTAIL.n250 B 0.021023f
C288 VTAIL.n251 B 0.009418f
C289 VTAIL.n252 B 0.008894f
C290 VTAIL.n253 B 0.016552f
C291 VTAIL.n254 B 0.016552f
C292 VTAIL.n255 B 0.008894f
C293 VTAIL.n256 B 0.009418f
C294 VTAIL.n257 B 0.021023f
C295 VTAIL.n258 B 0.021023f
C296 VTAIL.n259 B 0.009418f
C297 VTAIL.n260 B 0.008894f
C298 VTAIL.n261 B 0.016552f
C299 VTAIL.n262 B 0.016552f
C300 VTAIL.n263 B 0.008894f
C301 VTAIL.n264 B 0.009418f
C302 VTAIL.n265 B 0.021023f
C303 VTAIL.n266 B 0.021023f
C304 VTAIL.n267 B 0.009418f
C305 VTAIL.n268 B 0.008894f
C306 VTAIL.n269 B 0.016552f
C307 VTAIL.n270 B 0.016552f
C308 VTAIL.n271 B 0.008894f
C309 VTAIL.n272 B 0.009418f
C310 VTAIL.n273 B 0.021023f
C311 VTAIL.n274 B 0.021023f
C312 VTAIL.n275 B 0.009418f
C313 VTAIL.n276 B 0.008894f
C314 VTAIL.n277 B 0.016552f
C315 VTAIL.n278 B 0.016552f
C316 VTAIL.n279 B 0.008894f
C317 VTAIL.n280 B 0.008894f
C318 VTAIL.n281 B 0.009418f
C319 VTAIL.n282 B 0.021023f
C320 VTAIL.n283 B 0.021023f
C321 VTAIL.n284 B 0.021023f
C322 VTAIL.n285 B 0.009156f
C323 VTAIL.n286 B 0.008894f
C324 VTAIL.n287 B 0.016552f
C325 VTAIL.n288 B 0.016552f
C326 VTAIL.n289 B 0.008894f
C327 VTAIL.n290 B 0.009418f
C328 VTAIL.n291 B 0.021023f
C329 VTAIL.n292 B 0.021023f
C330 VTAIL.n293 B 0.009418f
C331 VTAIL.n294 B 0.008894f
C332 VTAIL.n295 B 0.016552f
C333 VTAIL.n296 B 0.016552f
C334 VTAIL.n297 B 0.008894f
C335 VTAIL.n298 B 0.009418f
C336 VTAIL.n299 B 0.021023f
C337 VTAIL.n300 B 0.043537f
C338 VTAIL.n301 B 0.009418f
C339 VTAIL.n302 B 0.008894f
C340 VTAIL.n303 B 0.035998f
C341 VTAIL.n304 B 0.024086f
C342 VTAIL.n305 B 1.14991f
C343 VTAIL.n306 B 0.022149f
C344 VTAIL.n307 B 0.016552f
C345 VTAIL.n308 B 0.008894f
C346 VTAIL.n309 B 0.021023f
C347 VTAIL.n310 B 0.009418f
C348 VTAIL.n311 B 0.016552f
C349 VTAIL.n312 B 0.008894f
C350 VTAIL.n313 B 0.021023f
C351 VTAIL.n314 B 0.009418f
C352 VTAIL.n315 B 0.016552f
C353 VTAIL.n316 B 0.009156f
C354 VTAIL.n317 B 0.021023f
C355 VTAIL.n318 B 0.008894f
C356 VTAIL.n319 B 0.009418f
C357 VTAIL.n320 B 0.016552f
C358 VTAIL.n321 B 0.008894f
C359 VTAIL.n322 B 0.021023f
C360 VTAIL.n323 B 0.009418f
C361 VTAIL.n324 B 0.016552f
C362 VTAIL.n325 B 0.008894f
C363 VTAIL.n326 B 0.021023f
C364 VTAIL.n327 B 0.009418f
C365 VTAIL.n328 B 0.016552f
C366 VTAIL.n329 B 0.008894f
C367 VTAIL.n330 B 0.021023f
C368 VTAIL.n331 B 0.009418f
C369 VTAIL.n332 B 0.016552f
C370 VTAIL.n333 B 0.008894f
C371 VTAIL.n334 B 0.021023f
C372 VTAIL.n335 B 0.009418f
C373 VTAIL.n336 B 0.016552f
C374 VTAIL.n337 B 0.008894f
C375 VTAIL.n338 B 0.015767f
C376 VTAIL.n339 B 0.012419f
C377 VTAIL.t2 B 0.034843f
C378 VTAIL.n340 B 0.120988f
C379 VTAIL.n341 B 1.31511f
C380 VTAIL.n342 B 0.008894f
C381 VTAIL.n343 B 0.009418f
C382 VTAIL.n344 B 0.021023f
C383 VTAIL.n345 B 0.021023f
C384 VTAIL.n346 B 0.009418f
C385 VTAIL.n347 B 0.008894f
C386 VTAIL.n348 B 0.016552f
C387 VTAIL.n349 B 0.016552f
C388 VTAIL.n350 B 0.008894f
C389 VTAIL.n351 B 0.009418f
C390 VTAIL.n352 B 0.021023f
C391 VTAIL.n353 B 0.021023f
C392 VTAIL.n354 B 0.009418f
C393 VTAIL.n355 B 0.008894f
C394 VTAIL.n356 B 0.016552f
C395 VTAIL.n357 B 0.016552f
C396 VTAIL.n358 B 0.008894f
C397 VTAIL.n359 B 0.009418f
C398 VTAIL.n360 B 0.021023f
C399 VTAIL.n361 B 0.021023f
C400 VTAIL.n362 B 0.009418f
C401 VTAIL.n363 B 0.008894f
C402 VTAIL.n364 B 0.016552f
C403 VTAIL.n365 B 0.016552f
C404 VTAIL.n366 B 0.008894f
C405 VTAIL.n367 B 0.009418f
C406 VTAIL.n368 B 0.021023f
C407 VTAIL.n369 B 0.021023f
C408 VTAIL.n370 B 0.009418f
C409 VTAIL.n371 B 0.008894f
C410 VTAIL.n372 B 0.016552f
C411 VTAIL.n373 B 0.016552f
C412 VTAIL.n374 B 0.008894f
C413 VTAIL.n375 B 0.009418f
C414 VTAIL.n376 B 0.021023f
C415 VTAIL.n377 B 0.021023f
C416 VTAIL.n378 B 0.009418f
C417 VTAIL.n379 B 0.008894f
C418 VTAIL.n380 B 0.016552f
C419 VTAIL.n381 B 0.016552f
C420 VTAIL.n382 B 0.008894f
C421 VTAIL.n383 B 0.009418f
C422 VTAIL.n384 B 0.021023f
C423 VTAIL.n385 B 0.021023f
C424 VTAIL.n386 B 0.021023f
C425 VTAIL.n387 B 0.009156f
C426 VTAIL.n388 B 0.008894f
C427 VTAIL.n389 B 0.016552f
C428 VTAIL.n390 B 0.016552f
C429 VTAIL.n391 B 0.008894f
C430 VTAIL.n392 B 0.009418f
C431 VTAIL.n393 B 0.021023f
C432 VTAIL.n394 B 0.021023f
C433 VTAIL.n395 B 0.009418f
C434 VTAIL.n396 B 0.008894f
C435 VTAIL.n397 B 0.016552f
C436 VTAIL.n398 B 0.016552f
C437 VTAIL.n399 B 0.008894f
C438 VTAIL.n400 B 0.009418f
C439 VTAIL.n401 B 0.021023f
C440 VTAIL.n402 B 0.043537f
C441 VTAIL.n403 B 0.009418f
C442 VTAIL.n404 B 0.008894f
C443 VTAIL.n405 B 0.035998f
C444 VTAIL.n406 B 0.024086f
C445 VTAIL.n407 B 1.14991f
C446 VTAIL.n408 B 0.022149f
C447 VTAIL.n409 B 0.016552f
C448 VTAIL.n410 B 0.008894f
C449 VTAIL.n411 B 0.021023f
C450 VTAIL.n412 B 0.009418f
C451 VTAIL.n413 B 0.016552f
C452 VTAIL.n414 B 0.008894f
C453 VTAIL.n415 B 0.021023f
C454 VTAIL.n416 B 0.009418f
C455 VTAIL.n417 B 0.016552f
C456 VTAIL.n418 B 0.009156f
C457 VTAIL.n419 B 0.021023f
C458 VTAIL.n420 B 0.008894f
C459 VTAIL.n421 B 0.009418f
C460 VTAIL.n422 B 0.016552f
C461 VTAIL.n423 B 0.008894f
C462 VTAIL.n424 B 0.021023f
C463 VTAIL.n425 B 0.009418f
C464 VTAIL.n426 B 0.016552f
C465 VTAIL.n427 B 0.008894f
C466 VTAIL.n428 B 0.021023f
C467 VTAIL.n429 B 0.009418f
C468 VTAIL.n430 B 0.016552f
C469 VTAIL.n431 B 0.008894f
C470 VTAIL.n432 B 0.021023f
C471 VTAIL.n433 B 0.009418f
C472 VTAIL.n434 B 0.016552f
C473 VTAIL.n435 B 0.008894f
C474 VTAIL.n436 B 0.021023f
C475 VTAIL.n437 B 0.009418f
C476 VTAIL.n438 B 0.016552f
C477 VTAIL.n439 B 0.008894f
C478 VTAIL.n440 B 0.015767f
C479 VTAIL.n441 B 0.012419f
C480 VTAIL.t0 B 0.034843f
C481 VTAIL.n442 B 0.120988f
C482 VTAIL.n443 B 1.31511f
C483 VTAIL.n444 B 0.008894f
C484 VTAIL.n445 B 0.009418f
C485 VTAIL.n446 B 0.021023f
C486 VTAIL.n447 B 0.021023f
C487 VTAIL.n448 B 0.009418f
C488 VTAIL.n449 B 0.008894f
C489 VTAIL.n450 B 0.016552f
C490 VTAIL.n451 B 0.016552f
C491 VTAIL.n452 B 0.008894f
C492 VTAIL.n453 B 0.009418f
C493 VTAIL.n454 B 0.021023f
C494 VTAIL.n455 B 0.021023f
C495 VTAIL.n456 B 0.009418f
C496 VTAIL.n457 B 0.008894f
C497 VTAIL.n458 B 0.016552f
C498 VTAIL.n459 B 0.016552f
C499 VTAIL.n460 B 0.008894f
C500 VTAIL.n461 B 0.009418f
C501 VTAIL.n462 B 0.021023f
C502 VTAIL.n463 B 0.021023f
C503 VTAIL.n464 B 0.009418f
C504 VTAIL.n465 B 0.008894f
C505 VTAIL.n466 B 0.016552f
C506 VTAIL.n467 B 0.016552f
C507 VTAIL.n468 B 0.008894f
C508 VTAIL.n469 B 0.009418f
C509 VTAIL.n470 B 0.021023f
C510 VTAIL.n471 B 0.021023f
C511 VTAIL.n472 B 0.009418f
C512 VTAIL.n473 B 0.008894f
C513 VTAIL.n474 B 0.016552f
C514 VTAIL.n475 B 0.016552f
C515 VTAIL.n476 B 0.008894f
C516 VTAIL.n477 B 0.009418f
C517 VTAIL.n478 B 0.021023f
C518 VTAIL.n479 B 0.021023f
C519 VTAIL.n480 B 0.009418f
C520 VTAIL.n481 B 0.008894f
C521 VTAIL.n482 B 0.016552f
C522 VTAIL.n483 B 0.016552f
C523 VTAIL.n484 B 0.008894f
C524 VTAIL.n485 B 0.009418f
C525 VTAIL.n486 B 0.021023f
C526 VTAIL.n487 B 0.021023f
C527 VTAIL.n488 B 0.021023f
C528 VTAIL.n489 B 0.009156f
C529 VTAIL.n490 B 0.008894f
C530 VTAIL.n491 B 0.016552f
C531 VTAIL.n492 B 0.016552f
C532 VTAIL.n493 B 0.008894f
C533 VTAIL.n494 B 0.009418f
C534 VTAIL.n495 B 0.021023f
C535 VTAIL.n496 B 0.021023f
C536 VTAIL.n497 B 0.009418f
C537 VTAIL.n498 B 0.008894f
C538 VTAIL.n499 B 0.016552f
C539 VTAIL.n500 B 0.016552f
C540 VTAIL.n501 B 0.008894f
C541 VTAIL.n502 B 0.009418f
C542 VTAIL.n503 B 0.021023f
C543 VTAIL.n504 B 0.043537f
C544 VTAIL.n505 B 0.009418f
C545 VTAIL.n506 B 0.008894f
C546 VTAIL.n507 B 0.035998f
C547 VTAIL.n508 B 0.024086f
C548 VTAIL.n509 B 0.077002f
C549 VTAIL.n510 B 0.022149f
C550 VTAIL.n511 B 0.016552f
C551 VTAIL.n512 B 0.008894f
C552 VTAIL.n513 B 0.021023f
C553 VTAIL.n514 B 0.009418f
C554 VTAIL.n515 B 0.016552f
C555 VTAIL.n516 B 0.008894f
C556 VTAIL.n517 B 0.021023f
C557 VTAIL.n518 B 0.009418f
C558 VTAIL.n519 B 0.016552f
C559 VTAIL.n520 B 0.009156f
C560 VTAIL.n521 B 0.021023f
C561 VTAIL.n522 B 0.008894f
C562 VTAIL.n523 B 0.009418f
C563 VTAIL.n524 B 0.016552f
C564 VTAIL.n525 B 0.008894f
C565 VTAIL.n526 B 0.021023f
C566 VTAIL.n527 B 0.009418f
C567 VTAIL.n528 B 0.016552f
C568 VTAIL.n529 B 0.008894f
C569 VTAIL.n530 B 0.021023f
C570 VTAIL.n531 B 0.009418f
C571 VTAIL.n532 B 0.016552f
C572 VTAIL.n533 B 0.008894f
C573 VTAIL.n534 B 0.021023f
C574 VTAIL.n535 B 0.009418f
C575 VTAIL.n536 B 0.016552f
C576 VTAIL.n537 B 0.008894f
C577 VTAIL.n538 B 0.021023f
C578 VTAIL.n539 B 0.009418f
C579 VTAIL.n540 B 0.016552f
C580 VTAIL.n541 B 0.008894f
C581 VTAIL.n542 B 0.015767f
C582 VTAIL.n543 B 0.012419f
C583 VTAIL.t6 B 0.034843f
C584 VTAIL.n544 B 0.120988f
C585 VTAIL.n545 B 1.31511f
C586 VTAIL.n546 B 0.008894f
C587 VTAIL.n547 B 0.009418f
C588 VTAIL.n548 B 0.021023f
C589 VTAIL.n549 B 0.021023f
C590 VTAIL.n550 B 0.009418f
C591 VTAIL.n551 B 0.008894f
C592 VTAIL.n552 B 0.016552f
C593 VTAIL.n553 B 0.016552f
C594 VTAIL.n554 B 0.008894f
C595 VTAIL.n555 B 0.009418f
C596 VTAIL.n556 B 0.021023f
C597 VTAIL.n557 B 0.021023f
C598 VTAIL.n558 B 0.009418f
C599 VTAIL.n559 B 0.008894f
C600 VTAIL.n560 B 0.016552f
C601 VTAIL.n561 B 0.016552f
C602 VTAIL.n562 B 0.008894f
C603 VTAIL.n563 B 0.009418f
C604 VTAIL.n564 B 0.021023f
C605 VTAIL.n565 B 0.021023f
C606 VTAIL.n566 B 0.009418f
C607 VTAIL.n567 B 0.008894f
C608 VTAIL.n568 B 0.016552f
C609 VTAIL.n569 B 0.016552f
C610 VTAIL.n570 B 0.008894f
C611 VTAIL.n571 B 0.009418f
C612 VTAIL.n572 B 0.021023f
C613 VTAIL.n573 B 0.021023f
C614 VTAIL.n574 B 0.009418f
C615 VTAIL.n575 B 0.008894f
C616 VTAIL.n576 B 0.016552f
C617 VTAIL.n577 B 0.016552f
C618 VTAIL.n578 B 0.008894f
C619 VTAIL.n579 B 0.009418f
C620 VTAIL.n580 B 0.021023f
C621 VTAIL.n581 B 0.021023f
C622 VTAIL.n582 B 0.009418f
C623 VTAIL.n583 B 0.008894f
C624 VTAIL.n584 B 0.016552f
C625 VTAIL.n585 B 0.016552f
C626 VTAIL.n586 B 0.008894f
C627 VTAIL.n587 B 0.009418f
C628 VTAIL.n588 B 0.021023f
C629 VTAIL.n589 B 0.021023f
C630 VTAIL.n590 B 0.021023f
C631 VTAIL.n591 B 0.009156f
C632 VTAIL.n592 B 0.008894f
C633 VTAIL.n593 B 0.016552f
C634 VTAIL.n594 B 0.016552f
C635 VTAIL.n595 B 0.008894f
C636 VTAIL.n596 B 0.009418f
C637 VTAIL.n597 B 0.021023f
C638 VTAIL.n598 B 0.021023f
C639 VTAIL.n599 B 0.009418f
C640 VTAIL.n600 B 0.008894f
C641 VTAIL.n601 B 0.016552f
C642 VTAIL.n602 B 0.016552f
C643 VTAIL.n603 B 0.008894f
C644 VTAIL.n604 B 0.009418f
C645 VTAIL.n605 B 0.021023f
C646 VTAIL.n606 B 0.043537f
C647 VTAIL.n607 B 0.009418f
C648 VTAIL.n608 B 0.008894f
C649 VTAIL.n609 B 0.035998f
C650 VTAIL.n610 B 0.024086f
C651 VTAIL.n611 B 0.077002f
C652 VTAIL.n612 B 0.022149f
C653 VTAIL.n613 B 0.016552f
C654 VTAIL.n614 B 0.008894f
C655 VTAIL.n615 B 0.021023f
C656 VTAIL.n616 B 0.009418f
C657 VTAIL.n617 B 0.016552f
C658 VTAIL.n618 B 0.008894f
C659 VTAIL.n619 B 0.021023f
C660 VTAIL.n620 B 0.009418f
C661 VTAIL.n621 B 0.016552f
C662 VTAIL.n622 B 0.009156f
C663 VTAIL.n623 B 0.021023f
C664 VTAIL.n624 B 0.008894f
C665 VTAIL.n625 B 0.009418f
C666 VTAIL.n626 B 0.016552f
C667 VTAIL.n627 B 0.008894f
C668 VTAIL.n628 B 0.021023f
C669 VTAIL.n629 B 0.009418f
C670 VTAIL.n630 B 0.016552f
C671 VTAIL.n631 B 0.008894f
C672 VTAIL.n632 B 0.021023f
C673 VTAIL.n633 B 0.009418f
C674 VTAIL.n634 B 0.016552f
C675 VTAIL.n635 B 0.008894f
C676 VTAIL.n636 B 0.021023f
C677 VTAIL.n637 B 0.009418f
C678 VTAIL.n638 B 0.016552f
C679 VTAIL.n639 B 0.008894f
C680 VTAIL.n640 B 0.021023f
C681 VTAIL.n641 B 0.009418f
C682 VTAIL.n642 B 0.016552f
C683 VTAIL.n643 B 0.008894f
C684 VTAIL.n644 B 0.015767f
C685 VTAIL.n645 B 0.012419f
C686 VTAIL.t4 B 0.034843f
C687 VTAIL.n646 B 0.120988f
C688 VTAIL.n647 B 1.31511f
C689 VTAIL.n648 B 0.008894f
C690 VTAIL.n649 B 0.009418f
C691 VTAIL.n650 B 0.021023f
C692 VTAIL.n651 B 0.021023f
C693 VTAIL.n652 B 0.009418f
C694 VTAIL.n653 B 0.008894f
C695 VTAIL.n654 B 0.016552f
C696 VTAIL.n655 B 0.016552f
C697 VTAIL.n656 B 0.008894f
C698 VTAIL.n657 B 0.009418f
C699 VTAIL.n658 B 0.021023f
C700 VTAIL.n659 B 0.021023f
C701 VTAIL.n660 B 0.009418f
C702 VTAIL.n661 B 0.008894f
C703 VTAIL.n662 B 0.016552f
C704 VTAIL.n663 B 0.016552f
C705 VTAIL.n664 B 0.008894f
C706 VTAIL.n665 B 0.009418f
C707 VTAIL.n666 B 0.021023f
C708 VTAIL.n667 B 0.021023f
C709 VTAIL.n668 B 0.009418f
C710 VTAIL.n669 B 0.008894f
C711 VTAIL.n670 B 0.016552f
C712 VTAIL.n671 B 0.016552f
C713 VTAIL.n672 B 0.008894f
C714 VTAIL.n673 B 0.009418f
C715 VTAIL.n674 B 0.021023f
C716 VTAIL.n675 B 0.021023f
C717 VTAIL.n676 B 0.009418f
C718 VTAIL.n677 B 0.008894f
C719 VTAIL.n678 B 0.016552f
C720 VTAIL.n679 B 0.016552f
C721 VTAIL.n680 B 0.008894f
C722 VTAIL.n681 B 0.009418f
C723 VTAIL.n682 B 0.021023f
C724 VTAIL.n683 B 0.021023f
C725 VTAIL.n684 B 0.009418f
C726 VTAIL.n685 B 0.008894f
C727 VTAIL.n686 B 0.016552f
C728 VTAIL.n687 B 0.016552f
C729 VTAIL.n688 B 0.008894f
C730 VTAIL.n689 B 0.009418f
C731 VTAIL.n690 B 0.021023f
C732 VTAIL.n691 B 0.021023f
C733 VTAIL.n692 B 0.021023f
C734 VTAIL.n693 B 0.009156f
C735 VTAIL.n694 B 0.008894f
C736 VTAIL.n695 B 0.016552f
C737 VTAIL.n696 B 0.016552f
C738 VTAIL.n697 B 0.008894f
C739 VTAIL.n698 B 0.009418f
C740 VTAIL.n699 B 0.021023f
C741 VTAIL.n700 B 0.021023f
C742 VTAIL.n701 B 0.009418f
C743 VTAIL.n702 B 0.008894f
C744 VTAIL.n703 B 0.016552f
C745 VTAIL.n704 B 0.016552f
C746 VTAIL.n705 B 0.008894f
C747 VTAIL.n706 B 0.009418f
C748 VTAIL.n707 B 0.021023f
C749 VTAIL.n708 B 0.043537f
C750 VTAIL.n709 B 0.009418f
C751 VTAIL.n710 B 0.008894f
C752 VTAIL.n711 B 0.035998f
C753 VTAIL.n712 B 0.024086f
C754 VTAIL.n713 B 1.14991f
C755 VTAIL.n714 B 0.022149f
C756 VTAIL.n715 B 0.016552f
C757 VTAIL.n716 B 0.008894f
C758 VTAIL.n717 B 0.021023f
C759 VTAIL.n718 B 0.009418f
C760 VTAIL.n719 B 0.016552f
C761 VTAIL.n720 B 0.008894f
C762 VTAIL.n721 B 0.021023f
C763 VTAIL.n722 B 0.009418f
C764 VTAIL.n723 B 0.016552f
C765 VTAIL.n724 B 0.009156f
C766 VTAIL.n725 B 0.021023f
C767 VTAIL.n726 B 0.009418f
C768 VTAIL.n727 B 0.016552f
C769 VTAIL.n728 B 0.008894f
C770 VTAIL.n729 B 0.021023f
C771 VTAIL.n730 B 0.009418f
C772 VTAIL.n731 B 0.016552f
C773 VTAIL.n732 B 0.008894f
C774 VTAIL.n733 B 0.021023f
C775 VTAIL.n734 B 0.009418f
C776 VTAIL.n735 B 0.016552f
C777 VTAIL.n736 B 0.008894f
C778 VTAIL.n737 B 0.021023f
C779 VTAIL.n738 B 0.009418f
C780 VTAIL.n739 B 0.016552f
C781 VTAIL.n740 B 0.008894f
C782 VTAIL.n741 B 0.021023f
C783 VTAIL.n742 B 0.009418f
C784 VTAIL.n743 B 0.016552f
C785 VTAIL.n744 B 0.008894f
C786 VTAIL.n745 B 0.015767f
C787 VTAIL.n746 B 0.012419f
C788 VTAIL.t1 B 0.034843f
C789 VTAIL.n747 B 0.120988f
C790 VTAIL.n748 B 1.31511f
C791 VTAIL.n749 B 0.008894f
C792 VTAIL.n750 B 0.009418f
C793 VTAIL.n751 B 0.021023f
C794 VTAIL.n752 B 0.021023f
C795 VTAIL.n753 B 0.009418f
C796 VTAIL.n754 B 0.008894f
C797 VTAIL.n755 B 0.016552f
C798 VTAIL.n756 B 0.016552f
C799 VTAIL.n757 B 0.008894f
C800 VTAIL.n758 B 0.009418f
C801 VTAIL.n759 B 0.021023f
C802 VTAIL.n760 B 0.021023f
C803 VTAIL.n761 B 0.009418f
C804 VTAIL.n762 B 0.008894f
C805 VTAIL.n763 B 0.016552f
C806 VTAIL.n764 B 0.016552f
C807 VTAIL.n765 B 0.008894f
C808 VTAIL.n766 B 0.009418f
C809 VTAIL.n767 B 0.021023f
C810 VTAIL.n768 B 0.021023f
C811 VTAIL.n769 B 0.009418f
C812 VTAIL.n770 B 0.008894f
C813 VTAIL.n771 B 0.016552f
C814 VTAIL.n772 B 0.016552f
C815 VTAIL.n773 B 0.008894f
C816 VTAIL.n774 B 0.009418f
C817 VTAIL.n775 B 0.021023f
C818 VTAIL.n776 B 0.021023f
C819 VTAIL.n777 B 0.009418f
C820 VTAIL.n778 B 0.008894f
C821 VTAIL.n779 B 0.016552f
C822 VTAIL.n780 B 0.016552f
C823 VTAIL.n781 B 0.008894f
C824 VTAIL.n782 B 0.009418f
C825 VTAIL.n783 B 0.021023f
C826 VTAIL.n784 B 0.021023f
C827 VTAIL.n785 B 0.009418f
C828 VTAIL.n786 B 0.008894f
C829 VTAIL.n787 B 0.016552f
C830 VTAIL.n788 B 0.016552f
C831 VTAIL.n789 B 0.008894f
C832 VTAIL.n790 B 0.008894f
C833 VTAIL.n791 B 0.009418f
C834 VTAIL.n792 B 0.021023f
C835 VTAIL.n793 B 0.021023f
C836 VTAIL.n794 B 0.021023f
C837 VTAIL.n795 B 0.009156f
C838 VTAIL.n796 B 0.008894f
C839 VTAIL.n797 B 0.016552f
C840 VTAIL.n798 B 0.016552f
C841 VTAIL.n799 B 0.008894f
C842 VTAIL.n800 B 0.009418f
C843 VTAIL.n801 B 0.021023f
C844 VTAIL.n802 B 0.021023f
C845 VTAIL.n803 B 0.009418f
C846 VTAIL.n804 B 0.008894f
C847 VTAIL.n805 B 0.016552f
C848 VTAIL.n806 B 0.016552f
C849 VTAIL.n807 B 0.008894f
C850 VTAIL.n808 B 0.009418f
C851 VTAIL.n809 B 0.021023f
C852 VTAIL.n810 B 0.043537f
C853 VTAIL.n811 B 0.009418f
C854 VTAIL.n812 B 0.008894f
C855 VTAIL.n813 B 0.035998f
C856 VTAIL.n814 B 0.024086f
C857 VTAIL.n815 B 1.12727f
C858 VP.t0 B 1.47223f
C859 VP.t2 B 1.47224f
C860 VP.n0 B 2.07367f
C861 VP.n1 B 4.08683f
C862 VP.t3 B 1.45984f
C863 VP.n2 B 0.554158f
C864 VP.t1 B 1.45984f
C865 VP.n3 B 0.554158f
C866 VP.n4 B 0.042306f
.ends

