* NGSPICE file created from diff_pair_sample_0040.ext - technology: sky130A

.subckt diff_pair_sample_0040 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t1 VP.t0 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0.7449 ps=4.6 w=1.91 l=2.29
X1 VDD1.t0 VP.t1 VTAIL.t2 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0.7449 ps=4.6 w=1.91 l=2.29
X2 B.t15 B.t13 B.t14 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0 ps=0 w=1.91 l=2.29
X3 VDD2.t1 VN.t0 VTAIL.t3 B.t1 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0.7449 ps=4.6 w=1.91 l=2.29
X4 B.t12 B.t10 B.t11 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0 ps=0 w=1.91 l=2.29
X5 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0 ps=0 w=1.91 l=2.29
X6 B.t5 B.t2 B.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0 ps=0 w=1.91 l=2.29
X7 VDD2.t0 VN.t1 VTAIL.t0 B.t0 sky130_fd_pr__nfet_01v8 ad=0.7449 pd=4.6 as=0.7449 ps=4.6 w=1.91 l=2.29
R0 VP.n0 VP.t1 105.463
R1 VP.n0 VP.t0 69.2717
R2 VP VP.n0 0.336784
R3 VTAIL.n26 VTAIL.n24 289.615
R4 VTAIL.n2 VTAIL.n0 289.615
R5 VTAIL.n18 VTAIL.n16 289.615
R6 VTAIL.n10 VTAIL.n8 289.615
R7 VTAIL.n27 VTAIL.n26 185
R8 VTAIL.n3 VTAIL.n2 185
R9 VTAIL.n19 VTAIL.n18 185
R10 VTAIL.n11 VTAIL.n10 185
R11 VTAIL.t0 VTAIL.n25 164.876
R12 VTAIL.t1 VTAIL.n1 164.876
R13 VTAIL.t2 VTAIL.n17 164.876
R14 VTAIL.t3 VTAIL.n9 164.876
R15 VTAIL.n26 VTAIL.t0 52.3082
R16 VTAIL.n2 VTAIL.t1 52.3082
R17 VTAIL.n18 VTAIL.t2 52.3082
R18 VTAIL.n10 VTAIL.t3 52.3082
R19 VTAIL.n31 VTAIL.n30 36.646
R20 VTAIL.n7 VTAIL.n6 36.646
R21 VTAIL.n23 VTAIL.n22 36.646
R22 VTAIL.n15 VTAIL.n14 36.646
R23 VTAIL.n15 VTAIL.n7 18.5307
R24 VTAIL.n31 VTAIL.n23 16.2721
R25 VTAIL.n27 VTAIL.n25 14.7318
R26 VTAIL.n3 VTAIL.n1 14.7318
R27 VTAIL.n19 VTAIL.n17 14.7318
R28 VTAIL.n11 VTAIL.n9 14.7318
R29 VTAIL.n28 VTAIL.n24 12.8005
R30 VTAIL.n4 VTAIL.n0 12.8005
R31 VTAIL.n20 VTAIL.n16 12.8005
R32 VTAIL.n12 VTAIL.n8 12.8005
R33 VTAIL.n30 VTAIL.n29 9.45567
R34 VTAIL.n6 VTAIL.n5 9.45567
R35 VTAIL.n22 VTAIL.n21 9.45567
R36 VTAIL.n14 VTAIL.n13 9.45567
R37 VTAIL.n29 VTAIL.n28 9.3005
R38 VTAIL.n5 VTAIL.n4 9.3005
R39 VTAIL.n21 VTAIL.n20 9.3005
R40 VTAIL.n13 VTAIL.n12 9.3005
R41 VTAIL.n29 VTAIL.n25 5.62509
R42 VTAIL.n5 VTAIL.n1 5.62509
R43 VTAIL.n21 VTAIL.n17 5.62509
R44 VTAIL.n13 VTAIL.n9 5.62509
R45 VTAIL.n23 VTAIL.n15 1.59964
R46 VTAIL.n30 VTAIL.n24 1.16414
R47 VTAIL.n6 VTAIL.n0 1.16414
R48 VTAIL.n22 VTAIL.n16 1.16414
R49 VTAIL.n14 VTAIL.n8 1.16414
R50 VTAIL VTAIL.n7 1.09317
R51 VTAIL VTAIL.n31 0.506965
R52 VTAIL.n28 VTAIL.n27 0.388379
R53 VTAIL.n4 VTAIL.n3 0.388379
R54 VTAIL.n20 VTAIL.n19 0.388379
R55 VTAIL.n12 VTAIL.n11 0.388379
R56 VDD1.n2 VDD1.n0 289.615
R57 VDD1.n9 VDD1.n7 289.615
R58 VDD1.n3 VDD1.n2 185
R59 VDD1.n10 VDD1.n9 185
R60 VDD1.t0 VDD1.n1 164.876
R61 VDD1.t1 VDD1.n8 164.876
R62 VDD1 VDD1.n13 84.2375
R63 VDD1 VDD1.n6 53.9476
R64 VDD1.n2 VDD1.t0 52.3082
R65 VDD1.n9 VDD1.t1 52.3082
R66 VDD1.n3 VDD1.n1 14.7318
R67 VDD1.n10 VDD1.n8 14.7318
R68 VDD1.n4 VDD1.n0 12.8005
R69 VDD1.n11 VDD1.n7 12.8005
R70 VDD1.n6 VDD1.n5 9.45567
R71 VDD1.n13 VDD1.n12 9.45567
R72 VDD1.n5 VDD1.n4 9.3005
R73 VDD1.n12 VDD1.n11 9.3005
R74 VDD1.n5 VDD1.n1 5.62509
R75 VDD1.n12 VDD1.n8 5.62509
R76 VDD1.n6 VDD1.n0 1.16414
R77 VDD1.n13 VDD1.n7 1.16414
R78 VDD1.n4 VDD1.n3 0.388379
R79 VDD1.n11 VDD1.n10 0.388379
R80 B.n363 B.n362 585
R81 B.n364 B.n363 585
R82 B.n129 B.n63 585
R83 B.n128 B.n127 585
R84 B.n126 B.n125 585
R85 B.n124 B.n123 585
R86 B.n122 B.n121 585
R87 B.n120 B.n119 585
R88 B.n118 B.n117 585
R89 B.n116 B.n115 585
R90 B.n114 B.n113 585
R91 B.n112 B.n111 585
R92 B.n110 B.n109 585
R93 B.n107 B.n106 585
R94 B.n105 B.n104 585
R95 B.n103 B.n102 585
R96 B.n101 B.n100 585
R97 B.n99 B.n98 585
R98 B.n97 B.n96 585
R99 B.n95 B.n94 585
R100 B.n93 B.n92 585
R101 B.n91 B.n90 585
R102 B.n89 B.n88 585
R103 B.n87 B.n86 585
R104 B.n85 B.n84 585
R105 B.n83 B.n82 585
R106 B.n81 B.n80 585
R107 B.n79 B.n78 585
R108 B.n77 B.n76 585
R109 B.n75 B.n74 585
R110 B.n73 B.n72 585
R111 B.n71 B.n70 585
R112 B.n47 B.n46 585
R113 B.n367 B.n366 585
R114 B.n361 B.n64 585
R115 B.n64 B.n44 585
R116 B.n360 B.n43 585
R117 B.n371 B.n43 585
R118 B.n359 B.n42 585
R119 B.n372 B.n42 585
R120 B.n358 B.n41 585
R121 B.n373 B.n41 585
R122 B.n357 B.n356 585
R123 B.n356 B.n37 585
R124 B.n355 B.n36 585
R125 B.n379 B.n36 585
R126 B.n354 B.n35 585
R127 B.n380 B.n35 585
R128 B.n353 B.n34 585
R129 B.n381 B.n34 585
R130 B.n352 B.n351 585
R131 B.n351 B.n30 585
R132 B.n350 B.n29 585
R133 B.n387 B.n29 585
R134 B.n349 B.n28 585
R135 B.n388 B.n28 585
R136 B.n348 B.n27 585
R137 B.n389 B.n27 585
R138 B.n347 B.n346 585
R139 B.n346 B.n23 585
R140 B.n345 B.n22 585
R141 B.n395 B.n22 585
R142 B.n344 B.n21 585
R143 B.n396 B.n21 585
R144 B.n343 B.n20 585
R145 B.n397 B.n20 585
R146 B.n342 B.n341 585
R147 B.n341 B.n16 585
R148 B.n340 B.n15 585
R149 B.n403 B.n15 585
R150 B.n339 B.n14 585
R151 B.n404 B.n14 585
R152 B.n338 B.n13 585
R153 B.n405 B.n13 585
R154 B.n337 B.n336 585
R155 B.n336 B.n12 585
R156 B.n335 B.n334 585
R157 B.n335 B.n8 585
R158 B.n333 B.n7 585
R159 B.n412 B.n7 585
R160 B.n332 B.n6 585
R161 B.n413 B.n6 585
R162 B.n331 B.n5 585
R163 B.n414 B.n5 585
R164 B.n330 B.n329 585
R165 B.n329 B.n4 585
R166 B.n328 B.n130 585
R167 B.n328 B.n327 585
R168 B.n318 B.n131 585
R169 B.n132 B.n131 585
R170 B.n320 B.n319 585
R171 B.n321 B.n320 585
R172 B.n317 B.n136 585
R173 B.n140 B.n136 585
R174 B.n316 B.n315 585
R175 B.n315 B.n314 585
R176 B.n138 B.n137 585
R177 B.n139 B.n138 585
R178 B.n307 B.n306 585
R179 B.n308 B.n307 585
R180 B.n305 B.n145 585
R181 B.n145 B.n144 585
R182 B.n304 B.n303 585
R183 B.n303 B.n302 585
R184 B.n147 B.n146 585
R185 B.n148 B.n147 585
R186 B.n295 B.n294 585
R187 B.n296 B.n295 585
R188 B.n293 B.n153 585
R189 B.n153 B.n152 585
R190 B.n292 B.n291 585
R191 B.n291 B.n290 585
R192 B.n155 B.n154 585
R193 B.n156 B.n155 585
R194 B.n283 B.n282 585
R195 B.n284 B.n283 585
R196 B.n281 B.n161 585
R197 B.n161 B.n160 585
R198 B.n280 B.n279 585
R199 B.n279 B.n278 585
R200 B.n163 B.n162 585
R201 B.n164 B.n163 585
R202 B.n271 B.n270 585
R203 B.n272 B.n271 585
R204 B.n269 B.n169 585
R205 B.n169 B.n168 585
R206 B.n268 B.n267 585
R207 B.n267 B.n266 585
R208 B.n171 B.n170 585
R209 B.n172 B.n171 585
R210 B.n262 B.n261 585
R211 B.n175 B.n174 585
R212 B.n258 B.n257 585
R213 B.n259 B.n258 585
R214 B.n256 B.n191 585
R215 B.n255 B.n254 585
R216 B.n253 B.n252 585
R217 B.n251 B.n250 585
R218 B.n249 B.n248 585
R219 B.n247 B.n246 585
R220 B.n245 B.n244 585
R221 B.n243 B.n242 585
R222 B.n241 B.n240 585
R223 B.n238 B.n237 585
R224 B.n236 B.n235 585
R225 B.n234 B.n233 585
R226 B.n232 B.n231 585
R227 B.n230 B.n229 585
R228 B.n228 B.n227 585
R229 B.n226 B.n225 585
R230 B.n224 B.n223 585
R231 B.n222 B.n221 585
R232 B.n220 B.n219 585
R233 B.n218 B.n217 585
R234 B.n216 B.n215 585
R235 B.n214 B.n213 585
R236 B.n212 B.n211 585
R237 B.n210 B.n209 585
R238 B.n208 B.n207 585
R239 B.n206 B.n205 585
R240 B.n204 B.n203 585
R241 B.n202 B.n201 585
R242 B.n200 B.n199 585
R243 B.n198 B.n197 585
R244 B.n263 B.n173 585
R245 B.n173 B.n172 585
R246 B.n265 B.n264 585
R247 B.n266 B.n265 585
R248 B.n167 B.n166 585
R249 B.n168 B.n167 585
R250 B.n274 B.n273 585
R251 B.n273 B.n272 585
R252 B.n275 B.n165 585
R253 B.n165 B.n164 585
R254 B.n277 B.n276 585
R255 B.n278 B.n277 585
R256 B.n159 B.n158 585
R257 B.n160 B.n159 585
R258 B.n286 B.n285 585
R259 B.n285 B.n284 585
R260 B.n287 B.n157 585
R261 B.n157 B.n156 585
R262 B.n289 B.n288 585
R263 B.n290 B.n289 585
R264 B.n151 B.n150 585
R265 B.n152 B.n151 585
R266 B.n298 B.n297 585
R267 B.n297 B.n296 585
R268 B.n299 B.n149 585
R269 B.n149 B.n148 585
R270 B.n301 B.n300 585
R271 B.n302 B.n301 585
R272 B.n143 B.n142 585
R273 B.n144 B.n143 585
R274 B.n310 B.n309 585
R275 B.n309 B.n308 585
R276 B.n311 B.n141 585
R277 B.n141 B.n139 585
R278 B.n313 B.n312 585
R279 B.n314 B.n313 585
R280 B.n135 B.n134 585
R281 B.n140 B.n135 585
R282 B.n323 B.n322 585
R283 B.n322 B.n321 585
R284 B.n324 B.n133 585
R285 B.n133 B.n132 585
R286 B.n326 B.n325 585
R287 B.n327 B.n326 585
R288 B.n3 B.n0 585
R289 B.n4 B.n3 585
R290 B.n411 B.n1 585
R291 B.n412 B.n411 585
R292 B.n410 B.n409 585
R293 B.n410 B.n8 585
R294 B.n408 B.n9 585
R295 B.n12 B.n9 585
R296 B.n407 B.n406 585
R297 B.n406 B.n405 585
R298 B.n11 B.n10 585
R299 B.n404 B.n11 585
R300 B.n402 B.n401 585
R301 B.n403 B.n402 585
R302 B.n400 B.n17 585
R303 B.n17 B.n16 585
R304 B.n399 B.n398 585
R305 B.n398 B.n397 585
R306 B.n19 B.n18 585
R307 B.n396 B.n19 585
R308 B.n394 B.n393 585
R309 B.n395 B.n394 585
R310 B.n392 B.n24 585
R311 B.n24 B.n23 585
R312 B.n391 B.n390 585
R313 B.n390 B.n389 585
R314 B.n26 B.n25 585
R315 B.n388 B.n26 585
R316 B.n386 B.n385 585
R317 B.n387 B.n386 585
R318 B.n384 B.n31 585
R319 B.n31 B.n30 585
R320 B.n383 B.n382 585
R321 B.n382 B.n381 585
R322 B.n33 B.n32 585
R323 B.n380 B.n33 585
R324 B.n378 B.n377 585
R325 B.n379 B.n378 585
R326 B.n376 B.n38 585
R327 B.n38 B.n37 585
R328 B.n375 B.n374 585
R329 B.n374 B.n373 585
R330 B.n40 B.n39 585
R331 B.n372 B.n40 585
R332 B.n370 B.n369 585
R333 B.n371 B.n370 585
R334 B.n368 B.n45 585
R335 B.n45 B.n44 585
R336 B.n415 B.n414 585
R337 B.n413 B.n2 585
R338 B.n366 B.n45 540.549
R339 B.n363 B.n64 540.549
R340 B.n197 B.n171 540.549
R341 B.n261 B.n173 540.549
R342 B.n364 B.n62 256.663
R343 B.n364 B.n61 256.663
R344 B.n364 B.n60 256.663
R345 B.n364 B.n59 256.663
R346 B.n364 B.n58 256.663
R347 B.n364 B.n57 256.663
R348 B.n364 B.n56 256.663
R349 B.n364 B.n55 256.663
R350 B.n364 B.n54 256.663
R351 B.n364 B.n53 256.663
R352 B.n364 B.n52 256.663
R353 B.n364 B.n51 256.663
R354 B.n364 B.n50 256.663
R355 B.n364 B.n49 256.663
R356 B.n364 B.n48 256.663
R357 B.n365 B.n364 256.663
R358 B.n260 B.n259 256.663
R359 B.n259 B.n176 256.663
R360 B.n259 B.n177 256.663
R361 B.n259 B.n178 256.663
R362 B.n259 B.n179 256.663
R363 B.n259 B.n180 256.663
R364 B.n259 B.n181 256.663
R365 B.n259 B.n182 256.663
R366 B.n259 B.n183 256.663
R367 B.n259 B.n184 256.663
R368 B.n259 B.n185 256.663
R369 B.n259 B.n186 256.663
R370 B.n259 B.n187 256.663
R371 B.n259 B.n188 256.663
R372 B.n259 B.n189 256.663
R373 B.n259 B.n190 256.663
R374 B.n417 B.n416 256.663
R375 B.n67 B.t6 227.626
R376 B.n65 B.t13 227.626
R377 B.n194 B.t10 227.626
R378 B.n192 B.t2 227.626
R379 B.n259 B.n172 191.371
R380 B.n364 B.n44 191.371
R381 B.n65 B.t14 172.085
R382 B.n194 B.t12 172.085
R383 B.n67 B.t8 172.084
R384 B.n192 B.t5 172.084
R385 B.n70 B.n47 163.367
R386 B.n74 B.n73 163.367
R387 B.n78 B.n77 163.367
R388 B.n82 B.n81 163.367
R389 B.n86 B.n85 163.367
R390 B.n90 B.n89 163.367
R391 B.n94 B.n93 163.367
R392 B.n98 B.n97 163.367
R393 B.n102 B.n101 163.367
R394 B.n106 B.n105 163.367
R395 B.n111 B.n110 163.367
R396 B.n115 B.n114 163.367
R397 B.n119 B.n118 163.367
R398 B.n123 B.n122 163.367
R399 B.n127 B.n126 163.367
R400 B.n363 B.n63 163.367
R401 B.n267 B.n171 163.367
R402 B.n267 B.n169 163.367
R403 B.n271 B.n169 163.367
R404 B.n271 B.n163 163.367
R405 B.n279 B.n163 163.367
R406 B.n279 B.n161 163.367
R407 B.n283 B.n161 163.367
R408 B.n283 B.n155 163.367
R409 B.n291 B.n155 163.367
R410 B.n291 B.n153 163.367
R411 B.n295 B.n153 163.367
R412 B.n295 B.n147 163.367
R413 B.n303 B.n147 163.367
R414 B.n303 B.n145 163.367
R415 B.n307 B.n145 163.367
R416 B.n307 B.n138 163.367
R417 B.n315 B.n138 163.367
R418 B.n315 B.n136 163.367
R419 B.n320 B.n136 163.367
R420 B.n320 B.n131 163.367
R421 B.n328 B.n131 163.367
R422 B.n329 B.n328 163.367
R423 B.n329 B.n5 163.367
R424 B.n6 B.n5 163.367
R425 B.n7 B.n6 163.367
R426 B.n335 B.n7 163.367
R427 B.n336 B.n335 163.367
R428 B.n336 B.n13 163.367
R429 B.n14 B.n13 163.367
R430 B.n15 B.n14 163.367
R431 B.n341 B.n15 163.367
R432 B.n341 B.n20 163.367
R433 B.n21 B.n20 163.367
R434 B.n22 B.n21 163.367
R435 B.n346 B.n22 163.367
R436 B.n346 B.n27 163.367
R437 B.n28 B.n27 163.367
R438 B.n29 B.n28 163.367
R439 B.n351 B.n29 163.367
R440 B.n351 B.n34 163.367
R441 B.n35 B.n34 163.367
R442 B.n36 B.n35 163.367
R443 B.n356 B.n36 163.367
R444 B.n356 B.n41 163.367
R445 B.n42 B.n41 163.367
R446 B.n43 B.n42 163.367
R447 B.n64 B.n43 163.367
R448 B.n258 B.n175 163.367
R449 B.n258 B.n191 163.367
R450 B.n254 B.n253 163.367
R451 B.n250 B.n249 163.367
R452 B.n246 B.n245 163.367
R453 B.n242 B.n241 163.367
R454 B.n237 B.n236 163.367
R455 B.n233 B.n232 163.367
R456 B.n229 B.n228 163.367
R457 B.n225 B.n224 163.367
R458 B.n221 B.n220 163.367
R459 B.n217 B.n216 163.367
R460 B.n213 B.n212 163.367
R461 B.n209 B.n208 163.367
R462 B.n205 B.n204 163.367
R463 B.n201 B.n200 163.367
R464 B.n265 B.n173 163.367
R465 B.n265 B.n167 163.367
R466 B.n273 B.n167 163.367
R467 B.n273 B.n165 163.367
R468 B.n277 B.n165 163.367
R469 B.n277 B.n159 163.367
R470 B.n285 B.n159 163.367
R471 B.n285 B.n157 163.367
R472 B.n289 B.n157 163.367
R473 B.n289 B.n151 163.367
R474 B.n297 B.n151 163.367
R475 B.n297 B.n149 163.367
R476 B.n301 B.n149 163.367
R477 B.n301 B.n143 163.367
R478 B.n309 B.n143 163.367
R479 B.n309 B.n141 163.367
R480 B.n313 B.n141 163.367
R481 B.n313 B.n135 163.367
R482 B.n322 B.n135 163.367
R483 B.n322 B.n133 163.367
R484 B.n326 B.n133 163.367
R485 B.n326 B.n3 163.367
R486 B.n415 B.n3 163.367
R487 B.n411 B.n2 163.367
R488 B.n411 B.n410 163.367
R489 B.n410 B.n9 163.367
R490 B.n406 B.n9 163.367
R491 B.n406 B.n11 163.367
R492 B.n402 B.n11 163.367
R493 B.n402 B.n17 163.367
R494 B.n398 B.n17 163.367
R495 B.n398 B.n19 163.367
R496 B.n394 B.n19 163.367
R497 B.n394 B.n24 163.367
R498 B.n390 B.n24 163.367
R499 B.n390 B.n26 163.367
R500 B.n386 B.n26 163.367
R501 B.n386 B.n31 163.367
R502 B.n382 B.n31 163.367
R503 B.n382 B.n33 163.367
R504 B.n378 B.n33 163.367
R505 B.n378 B.n38 163.367
R506 B.n374 B.n38 163.367
R507 B.n374 B.n40 163.367
R508 B.n370 B.n40 163.367
R509 B.n370 B.n45 163.367
R510 B.n66 B.t15 121.272
R511 B.n195 B.t11 121.272
R512 B.n68 B.t9 121.272
R513 B.n193 B.t4 121.272
R514 B.n266 B.n172 104.106
R515 B.n266 B.n168 104.106
R516 B.n272 B.n168 104.106
R517 B.n272 B.n164 104.106
R518 B.n278 B.n164 104.106
R519 B.n278 B.n160 104.106
R520 B.n284 B.n160 104.106
R521 B.n290 B.n156 104.106
R522 B.n290 B.n152 104.106
R523 B.n296 B.n152 104.106
R524 B.n296 B.n148 104.106
R525 B.n302 B.n148 104.106
R526 B.n302 B.n144 104.106
R527 B.n308 B.n144 104.106
R528 B.n308 B.n139 104.106
R529 B.n314 B.n139 104.106
R530 B.n314 B.n140 104.106
R531 B.n321 B.n132 104.106
R532 B.n327 B.n132 104.106
R533 B.n327 B.n4 104.106
R534 B.n414 B.n4 104.106
R535 B.n414 B.n413 104.106
R536 B.n413 B.n412 104.106
R537 B.n412 B.n8 104.106
R538 B.n12 B.n8 104.106
R539 B.n405 B.n12 104.106
R540 B.n404 B.n403 104.106
R541 B.n403 B.n16 104.106
R542 B.n397 B.n16 104.106
R543 B.n397 B.n396 104.106
R544 B.n396 B.n395 104.106
R545 B.n395 B.n23 104.106
R546 B.n389 B.n23 104.106
R547 B.n389 B.n388 104.106
R548 B.n388 B.n387 104.106
R549 B.n387 B.n30 104.106
R550 B.n381 B.n380 104.106
R551 B.n380 B.n379 104.106
R552 B.n379 B.n37 104.106
R553 B.n373 B.n37 104.106
R554 B.n373 B.n372 104.106
R555 B.n372 B.n371 104.106
R556 B.n371 B.n44 104.106
R557 B.n321 B.t1 99.5134
R558 B.n405 B.t0 99.5134
R559 B.t3 B.n156 90.3276
R560 B.t7 B.n30 90.3276
R561 B.n366 B.n365 71.676
R562 B.n70 B.n48 71.676
R563 B.n74 B.n49 71.676
R564 B.n78 B.n50 71.676
R565 B.n82 B.n51 71.676
R566 B.n86 B.n52 71.676
R567 B.n90 B.n53 71.676
R568 B.n94 B.n54 71.676
R569 B.n98 B.n55 71.676
R570 B.n102 B.n56 71.676
R571 B.n106 B.n57 71.676
R572 B.n111 B.n58 71.676
R573 B.n115 B.n59 71.676
R574 B.n119 B.n60 71.676
R575 B.n123 B.n61 71.676
R576 B.n127 B.n62 71.676
R577 B.n63 B.n62 71.676
R578 B.n126 B.n61 71.676
R579 B.n122 B.n60 71.676
R580 B.n118 B.n59 71.676
R581 B.n114 B.n58 71.676
R582 B.n110 B.n57 71.676
R583 B.n105 B.n56 71.676
R584 B.n101 B.n55 71.676
R585 B.n97 B.n54 71.676
R586 B.n93 B.n53 71.676
R587 B.n89 B.n52 71.676
R588 B.n85 B.n51 71.676
R589 B.n81 B.n50 71.676
R590 B.n77 B.n49 71.676
R591 B.n73 B.n48 71.676
R592 B.n365 B.n47 71.676
R593 B.n261 B.n260 71.676
R594 B.n191 B.n176 71.676
R595 B.n253 B.n177 71.676
R596 B.n249 B.n178 71.676
R597 B.n245 B.n179 71.676
R598 B.n241 B.n180 71.676
R599 B.n236 B.n181 71.676
R600 B.n232 B.n182 71.676
R601 B.n228 B.n183 71.676
R602 B.n224 B.n184 71.676
R603 B.n220 B.n185 71.676
R604 B.n216 B.n186 71.676
R605 B.n212 B.n187 71.676
R606 B.n208 B.n188 71.676
R607 B.n204 B.n189 71.676
R608 B.n200 B.n190 71.676
R609 B.n260 B.n175 71.676
R610 B.n254 B.n176 71.676
R611 B.n250 B.n177 71.676
R612 B.n246 B.n178 71.676
R613 B.n242 B.n179 71.676
R614 B.n237 B.n180 71.676
R615 B.n233 B.n181 71.676
R616 B.n229 B.n182 71.676
R617 B.n225 B.n183 71.676
R618 B.n221 B.n184 71.676
R619 B.n217 B.n185 71.676
R620 B.n213 B.n186 71.676
R621 B.n209 B.n187 71.676
R622 B.n205 B.n188 71.676
R623 B.n201 B.n189 71.676
R624 B.n197 B.n190 71.676
R625 B.n416 B.n415 71.676
R626 B.n416 B.n2 71.676
R627 B.n69 B.n68 59.5399
R628 B.n108 B.n66 59.5399
R629 B.n196 B.n195 59.5399
R630 B.n239 B.n193 59.5399
R631 B.n68 B.n67 50.8126
R632 B.n66 B.n65 50.8126
R633 B.n195 B.n194 50.8126
R634 B.n193 B.n192 50.8126
R635 B.n263 B.n262 35.1225
R636 B.n198 B.n170 35.1225
R637 B.n362 B.n361 35.1225
R638 B.n368 B.n367 35.1225
R639 B B.n417 18.0485
R640 B.n284 B.t3 13.7792
R641 B.n381 B.t7 13.7792
R642 B.n264 B.n263 10.6151
R643 B.n264 B.n166 10.6151
R644 B.n274 B.n166 10.6151
R645 B.n275 B.n274 10.6151
R646 B.n276 B.n275 10.6151
R647 B.n276 B.n158 10.6151
R648 B.n286 B.n158 10.6151
R649 B.n287 B.n286 10.6151
R650 B.n288 B.n287 10.6151
R651 B.n288 B.n150 10.6151
R652 B.n298 B.n150 10.6151
R653 B.n299 B.n298 10.6151
R654 B.n300 B.n299 10.6151
R655 B.n300 B.n142 10.6151
R656 B.n310 B.n142 10.6151
R657 B.n311 B.n310 10.6151
R658 B.n312 B.n311 10.6151
R659 B.n312 B.n134 10.6151
R660 B.n323 B.n134 10.6151
R661 B.n324 B.n323 10.6151
R662 B.n325 B.n324 10.6151
R663 B.n325 B.n0 10.6151
R664 B.n262 B.n174 10.6151
R665 B.n257 B.n174 10.6151
R666 B.n257 B.n256 10.6151
R667 B.n256 B.n255 10.6151
R668 B.n255 B.n252 10.6151
R669 B.n252 B.n251 10.6151
R670 B.n251 B.n248 10.6151
R671 B.n248 B.n247 10.6151
R672 B.n247 B.n244 10.6151
R673 B.n244 B.n243 10.6151
R674 B.n243 B.n240 10.6151
R675 B.n238 B.n235 10.6151
R676 B.n235 B.n234 10.6151
R677 B.n234 B.n231 10.6151
R678 B.n231 B.n230 10.6151
R679 B.n230 B.n227 10.6151
R680 B.n227 B.n226 10.6151
R681 B.n226 B.n223 10.6151
R682 B.n223 B.n222 10.6151
R683 B.n219 B.n218 10.6151
R684 B.n218 B.n215 10.6151
R685 B.n215 B.n214 10.6151
R686 B.n214 B.n211 10.6151
R687 B.n211 B.n210 10.6151
R688 B.n210 B.n207 10.6151
R689 B.n207 B.n206 10.6151
R690 B.n206 B.n203 10.6151
R691 B.n203 B.n202 10.6151
R692 B.n202 B.n199 10.6151
R693 B.n199 B.n198 10.6151
R694 B.n268 B.n170 10.6151
R695 B.n269 B.n268 10.6151
R696 B.n270 B.n269 10.6151
R697 B.n270 B.n162 10.6151
R698 B.n280 B.n162 10.6151
R699 B.n281 B.n280 10.6151
R700 B.n282 B.n281 10.6151
R701 B.n282 B.n154 10.6151
R702 B.n292 B.n154 10.6151
R703 B.n293 B.n292 10.6151
R704 B.n294 B.n293 10.6151
R705 B.n294 B.n146 10.6151
R706 B.n304 B.n146 10.6151
R707 B.n305 B.n304 10.6151
R708 B.n306 B.n305 10.6151
R709 B.n306 B.n137 10.6151
R710 B.n316 B.n137 10.6151
R711 B.n317 B.n316 10.6151
R712 B.n319 B.n317 10.6151
R713 B.n319 B.n318 10.6151
R714 B.n318 B.n130 10.6151
R715 B.n330 B.n130 10.6151
R716 B.n331 B.n330 10.6151
R717 B.n332 B.n331 10.6151
R718 B.n333 B.n332 10.6151
R719 B.n334 B.n333 10.6151
R720 B.n337 B.n334 10.6151
R721 B.n338 B.n337 10.6151
R722 B.n339 B.n338 10.6151
R723 B.n340 B.n339 10.6151
R724 B.n342 B.n340 10.6151
R725 B.n343 B.n342 10.6151
R726 B.n344 B.n343 10.6151
R727 B.n345 B.n344 10.6151
R728 B.n347 B.n345 10.6151
R729 B.n348 B.n347 10.6151
R730 B.n349 B.n348 10.6151
R731 B.n350 B.n349 10.6151
R732 B.n352 B.n350 10.6151
R733 B.n353 B.n352 10.6151
R734 B.n354 B.n353 10.6151
R735 B.n355 B.n354 10.6151
R736 B.n357 B.n355 10.6151
R737 B.n358 B.n357 10.6151
R738 B.n359 B.n358 10.6151
R739 B.n360 B.n359 10.6151
R740 B.n361 B.n360 10.6151
R741 B.n409 B.n1 10.6151
R742 B.n409 B.n408 10.6151
R743 B.n408 B.n407 10.6151
R744 B.n407 B.n10 10.6151
R745 B.n401 B.n10 10.6151
R746 B.n401 B.n400 10.6151
R747 B.n400 B.n399 10.6151
R748 B.n399 B.n18 10.6151
R749 B.n393 B.n18 10.6151
R750 B.n393 B.n392 10.6151
R751 B.n392 B.n391 10.6151
R752 B.n391 B.n25 10.6151
R753 B.n385 B.n25 10.6151
R754 B.n385 B.n384 10.6151
R755 B.n384 B.n383 10.6151
R756 B.n383 B.n32 10.6151
R757 B.n377 B.n32 10.6151
R758 B.n377 B.n376 10.6151
R759 B.n376 B.n375 10.6151
R760 B.n375 B.n39 10.6151
R761 B.n369 B.n39 10.6151
R762 B.n369 B.n368 10.6151
R763 B.n367 B.n46 10.6151
R764 B.n71 B.n46 10.6151
R765 B.n72 B.n71 10.6151
R766 B.n75 B.n72 10.6151
R767 B.n76 B.n75 10.6151
R768 B.n79 B.n76 10.6151
R769 B.n80 B.n79 10.6151
R770 B.n83 B.n80 10.6151
R771 B.n84 B.n83 10.6151
R772 B.n87 B.n84 10.6151
R773 B.n88 B.n87 10.6151
R774 B.n92 B.n91 10.6151
R775 B.n95 B.n92 10.6151
R776 B.n96 B.n95 10.6151
R777 B.n99 B.n96 10.6151
R778 B.n100 B.n99 10.6151
R779 B.n103 B.n100 10.6151
R780 B.n104 B.n103 10.6151
R781 B.n107 B.n104 10.6151
R782 B.n112 B.n109 10.6151
R783 B.n113 B.n112 10.6151
R784 B.n116 B.n113 10.6151
R785 B.n117 B.n116 10.6151
R786 B.n120 B.n117 10.6151
R787 B.n121 B.n120 10.6151
R788 B.n124 B.n121 10.6151
R789 B.n125 B.n124 10.6151
R790 B.n128 B.n125 10.6151
R791 B.n129 B.n128 10.6151
R792 B.n362 B.n129 10.6151
R793 B.n417 B.n0 8.11757
R794 B.n417 B.n1 8.11757
R795 B.n239 B.n238 6.5566
R796 B.n222 B.n196 6.5566
R797 B.n91 B.n69 6.5566
R798 B.n108 B.n107 6.5566
R799 B.n140 B.t1 4.5934
R800 B.t0 B.n404 4.5934
R801 B.n240 B.n239 4.05904
R802 B.n219 B.n196 4.05904
R803 B.n88 B.n69 4.05904
R804 B.n109 B.n108 4.05904
R805 VN VN.t0 105.558
R806 VN VN.t1 69.608
R807 VDD2.n9 VDD2.n7 289.615
R808 VDD2.n2 VDD2.n0 289.615
R809 VDD2.n10 VDD2.n9 185
R810 VDD2.n3 VDD2.n2 185
R811 VDD2.t1 VDD2.n8 164.876
R812 VDD2.t0 VDD2.n1 164.876
R813 VDD2.n14 VDD2.n6 83.148
R814 VDD2.n14 VDD2.n13 53.3247
R815 VDD2.n9 VDD2.t1 52.3082
R816 VDD2.n2 VDD2.t0 52.3082
R817 VDD2.n10 VDD2.n8 14.7318
R818 VDD2.n3 VDD2.n1 14.7318
R819 VDD2.n11 VDD2.n7 12.8005
R820 VDD2.n4 VDD2.n0 12.8005
R821 VDD2.n13 VDD2.n12 9.45567
R822 VDD2.n6 VDD2.n5 9.45567
R823 VDD2.n12 VDD2.n11 9.3005
R824 VDD2.n5 VDD2.n4 9.3005
R825 VDD2.n12 VDD2.n8 5.62509
R826 VDD2.n5 VDD2.n1 5.62509
R827 VDD2.n13 VDD2.n7 1.16414
R828 VDD2.n6 VDD2.n0 1.16414
R829 VDD2 VDD2.n14 0.623345
R830 VDD2.n11 VDD2.n10 0.388379
R831 VDD2.n4 VDD2.n3 0.388379
C0 VTAIL VP 0.914816f
C1 VTAIL VDD1 2.30113f
C2 VP VDD1 0.817206f
C3 VN VDD2 0.646842f
C4 VTAIL VN 0.900676f
C5 VTAIL VDD2 2.35194f
C6 VN VP 3.45063f
C7 VDD2 VP 0.326373f
C8 VN VDD1 0.154407f
C9 VDD2 VDD1 0.636242f
C10 VDD2 B 2.476978f
C11 VDD1 B 3.98724f
C12 VTAIL B 2.849394f
C13 VN B 7.21534f
C14 VP B 5.131906f
C15 VDD2.n0 B 0.024928f
C16 VDD2.n1 B 0.058457f
C17 VDD2.t0 B 0.041216f
C18 VDD2.n2 B 0.043129f
C19 VDD2.n3 B 0.011797f
C20 VDD2.n4 B 0.009576f
C21 VDD2.n5 B 0.115483f
C22 VDD2.n6 B 0.272194f
C23 VDD2.n7 B 0.024928f
C24 VDD2.n8 B 0.058457f
C25 VDD2.t1 B 0.041216f
C26 VDD2.n9 B 0.043129f
C27 VDD2.n10 B 0.011797f
C28 VDD2.n11 B 0.009576f
C29 VDD2.n12 B 0.115483f
C30 VDD2.n13 B 0.039706f
C31 VDD2.n14 B 1.37782f
C32 VN.t1 B 0.544928f
C33 VN.t0 B 0.950205f
C34 VDD1.n0 B 0.023252f
C35 VDD1.n1 B 0.054526f
C36 VDD1.t0 B 0.038444f
C37 VDD1.n2 B 0.040228f
C38 VDD1.n3 B 0.011004f
C39 VDD1.n4 B 0.008932f
C40 VDD1.n5 B 0.107717f
C41 VDD1.n6 B 0.037825f
C42 VDD1.n7 B 0.023252f
C43 VDD1.n8 B 0.054526f
C44 VDD1.t1 B 0.038444f
C45 VDD1.n9 B 0.040228f
C46 VDD1.n10 B 0.011004f
C47 VDD1.n11 B 0.008932f
C48 VDD1.n12 B 0.107717f
C49 VDD1.n13 B 0.27722f
C50 VTAIL.n0 B 0.030091f
C51 VTAIL.n1 B 0.070564f
C52 VTAIL.t1 B 0.049752f
C53 VTAIL.n2 B 0.05206f
C54 VTAIL.n3 B 0.01424f
C55 VTAIL.n4 B 0.011559f
C56 VTAIL.n5 B 0.139399f
C57 VTAIL.n6 B 0.033122f
C58 VTAIL.n7 B 0.817385f
C59 VTAIL.n8 B 0.030091f
C60 VTAIL.n9 B 0.070564f
C61 VTAIL.t3 B 0.049752f
C62 VTAIL.n10 B 0.05206f
C63 VTAIL.n11 B 0.01424f
C64 VTAIL.n12 B 0.011559f
C65 VTAIL.n13 B 0.139399f
C66 VTAIL.n14 B 0.033122f
C67 VTAIL.n15 B 0.85249f
C68 VTAIL.n16 B 0.030091f
C69 VTAIL.n17 B 0.070564f
C70 VTAIL.t2 B 0.049752f
C71 VTAIL.n18 B 0.05206f
C72 VTAIL.n19 B 0.01424f
C73 VTAIL.n20 B 0.011559f
C74 VTAIL.n21 B 0.139399f
C75 VTAIL.n22 B 0.033122f
C76 VTAIL.n23 B 0.695935f
C77 VTAIL.n24 B 0.030091f
C78 VTAIL.n25 B 0.070564f
C79 VTAIL.t0 B 0.049752f
C80 VTAIL.n26 B 0.05206f
C81 VTAIL.n27 B 0.01424f
C82 VTAIL.n28 B 0.011559f
C83 VTAIL.n29 B 0.139399f
C84 VTAIL.n30 B 0.033122f
C85 VTAIL.n31 B 0.620197f
C86 VP.t1 B 0.956982f
C87 VP.t0 B 0.550591f
C88 VP.n0 B 1.92791f
.ends

