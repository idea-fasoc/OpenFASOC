* NGSPICE file created from diff_pair_sample_1249.ext - technology: sky130A

.subckt diff_pair_sample_1249 VTAIL VN VP B VDD2 VDD1
X0 VDD1.t5 VP.t0 VTAIL.t10 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=1.2144 ps=7.69 w=7.36 l=1.4
X1 VDD2.t5 VN.t0 VTAIL.t2 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=1.2144 ps=7.69 w=7.36 l=1.4
X2 VTAIL.t8 VP.t1 VDD1.t4 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=1.2144 ps=7.69 w=7.36 l=1.4
X3 VDD1.t3 VP.t2 VTAIL.t11 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=2.8704 ps=15.5 w=7.36 l=1.4
X4 VDD1.t2 VP.t3 VTAIL.t6 B.t2 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=1.2144 ps=7.69 w=7.36 l=1.4
X5 B.t19 B.t17 B.t18 B.t14 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=0 ps=0 w=7.36 l=1.4
X6 VTAIL.t9 VP.t4 VDD1.t1 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=1.2144 ps=7.69 w=7.36 l=1.4
X7 VDD1.t0 VP.t5 VTAIL.t7 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=2.8704 ps=15.5 w=7.36 l=1.4
X8 B.t16 B.t13 B.t15 B.t14 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=0 ps=0 w=7.36 l=1.4
X9 VDD2.t4 VN.t1 VTAIL.t1 B.t1 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=2.8704 ps=15.5 w=7.36 l=1.4
X10 VTAIL.t0 VN.t2 VDD2.t3 B.t0 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=1.2144 ps=7.69 w=7.36 l=1.4
X11 VDD2.t2 VN.t3 VTAIL.t4 B.t4 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=2.8704 ps=15.5 w=7.36 l=1.4
X12 VDD2.t1 VN.t4 VTAIL.t5 B.t5 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=1.2144 ps=7.69 w=7.36 l=1.4
X13 VTAIL.t3 VN.t5 VDD2.t0 B.t3 sky130_fd_pr__nfet_01v8 ad=1.2144 pd=7.69 as=1.2144 ps=7.69 w=7.36 l=1.4
X14 B.t12 B.t10 B.t11 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=0 ps=0 w=7.36 l=1.4
X15 B.t9 B.t6 B.t8 B.t7 sky130_fd_pr__nfet_01v8 ad=2.8704 pd=15.5 as=0 ps=0 w=7.36 l=1.4
R0 VP.n15 VP.n14 174.581
R1 VP.n27 VP.n26 174.581
R2 VP.n13 VP.n12 174.581
R3 VP.n7 VP.t0 161.577
R4 VP.n8 VP.n5 161.3
R5 VP.n10 VP.n9 161.3
R6 VP.n11 VP.n4 161.3
R7 VP.n25 VP.n0 161.3
R8 VP.n24 VP.n23 161.3
R9 VP.n22 VP.n1 161.3
R10 VP.n21 VP.n20 161.3
R11 VP.n19 VP.n2 161.3
R12 VP.n18 VP.n17 161.3
R13 VP.n16 VP.n3 161.3
R14 VP.n20 VP.t1 126.698
R15 VP.n14 VP.t3 126.698
R16 VP.n26 VP.t2 126.698
R17 VP.n6 VP.t4 126.698
R18 VP.n12 VP.t5 126.698
R19 VP.n19 VP.n18 53.6554
R20 VP.n24 VP.n1 53.6554
R21 VP.n10 VP.n5 53.6554
R22 VP.n7 VP.n6 41.8949
R23 VP.n15 VP.n13 40.3755
R24 VP.n18 VP.n3 27.4986
R25 VP.n25 VP.n24 27.4986
R26 VP.n11 VP.n10 27.4986
R27 VP.n20 VP.n19 24.5923
R28 VP.n20 VP.n1 24.5923
R29 VP.n6 VP.n5 24.5923
R30 VP.n8 VP.n7 17.6108
R31 VP.n14 VP.n3 11.3127
R32 VP.n26 VP.n25 11.3127
R33 VP.n12 VP.n11 11.3127
R34 VP.n9 VP.n8 0.189894
R35 VP.n9 VP.n4 0.189894
R36 VP.n13 VP.n4 0.189894
R37 VP.n16 VP.n15 0.189894
R38 VP.n17 VP.n16 0.189894
R39 VP.n17 VP.n2 0.189894
R40 VP.n21 VP.n2 0.189894
R41 VP.n22 VP.n21 0.189894
R42 VP.n23 VP.n22 0.189894
R43 VP.n23 VP.n0 0.189894
R44 VP.n27 VP.n0 0.189894
R45 VP VP.n27 0.0516364
R46 VTAIL.n162 VTAIL.n128 289.615
R47 VTAIL.n36 VTAIL.n2 289.615
R48 VTAIL.n122 VTAIL.n88 289.615
R49 VTAIL.n80 VTAIL.n46 289.615
R50 VTAIL.n140 VTAIL.n139 185
R51 VTAIL.n145 VTAIL.n144 185
R52 VTAIL.n147 VTAIL.n146 185
R53 VTAIL.n136 VTAIL.n135 185
R54 VTAIL.n153 VTAIL.n152 185
R55 VTAIL.n155 VTAIL.n154 185
R56 VTAIL.n132 VTAIL.n131 185
R57 VTAIL.n161 VTAIL.n160 185
R58 VTAIL.n163 VTAIL.n162 185
R59 VTAIL.n14 VTAIL.n13 185
R60 VTAIL.n19 VTAIL.n18 185
R61 VTAIL.n21 VTAIL.n20 185
R62 VTAIL.n10 VTAIL.n9 185
R63 VTAIL.n27 VTAIL.n26 185
R64 VTAIL.n29 VTAIL.n28 185
R65 VTAIL.n6 VTAIL.n5 185
R66 VTAIL.n35 VTAIL.n34 185
R67 VTAIL.n37 VTAIL.n36 185
R68 VTAIL.n123 VTAIL.n122 185
R69 VTAIL.n121 VTAIL.n120 185
R70 VTAIL.n92 VTAIL.n91 185
R71 VTAIL.n115 VTAIL.n114 185
R72 VTAIL.n113 VTAIL.n112 185
R73 VTAIL.n96 VTAIL.n95 185
R74 VTAIL.n107 VTAIL.n106 185
R75 VTAIL.n105 VTAIL.n104 185
R76 VTAIL.n100 VTAIL.n99 185
R77 VTAIL.n81 VTAIL.n80 185
R78 VTAIL.n79 VTAIL.n78 185
R79 VTAIL.n50 VTAIL.n49 185
R80 VTAIL.n73 VTAIL.n72 185
R81 VTAIL.n71 VTAIL.n70 185
R82 VTAIL.n54 VTAIL.n53 185
R83 VTAIL.n65 VTAIL.n64 185
R84 VTAIL.n63 VTAIL.n62 185
R85 VTAIL.n58 VTAIL.n57 185
R86 VTAIL.n141 VTAIL.t4 147.659
R87 VTAIL.n15 VTAIL.t11 147.659
R88 VTAIL.n101 VTAIL.t7 147.659
R89 VTAIL.n59 VTAIL.t1 147.659
R90 VTAIL.n145 VTAIL.n139 104.615
R91 VTAIL.n146 VTAIL.n145 104.615
R92 VTAIL.n146 VTAIL.n135 104.615
R93 VTAIL.n153 VTAIL.n135 104.615
R94 VTAIL.n154 VTAIL.n153 104.615
R95 VTAIL.n154 VTAIL.n131 104.615
R96 VTAIL.n161 VTAIL.n131 104.615
R97 VTAIL.n162 VTAIL.n161 104.615
R98 VTAIL.n19 VTAIL.n13 104.615
R99 VTAIL.n20 VTAIL.n19 104.615
R100 VTAIL.n20 VTAIL.n9 104.615
R101 VTAIL.n27 VTAIL.n9 104.615
R102 VTAIL.n28 VTAIL.n27 104.615
R103 VTAIL.n28 VTAIL.n5 104.615
R104 VTAIL.n35 VTAIL.n5 104.615
R105 VTAIL.n36 VTAIL.n35 104.615
R106 VTAIL.n122 VTAIL.n121 104.615
R107 VTAIL.n121 VTAIL.n91 104.615
R108 VTAIL.n114 VTAIL.n91 104.615
R109 VTAIL.n114 VTAIL.n113 104.615
R110 VTAIL.n113 VTAIL.n95 104.615
R111 VTAIL.n106 VTAIL.n95 104.615
R112 VTAIL.n106 VTAIL.n105 104.615
R113 VTAIL.n105 VTAIL.n99 104.615
R114 VTAIL.n80 VTAIL.n79 104.615
R115 VTAIL.n79 VTAIL.n49 104.615
R116 VTAIL.n72 VTAIL.n49 104.615
R117 VTAIL.n72 VTAIL.n71 104.615
R118 VTAIL.n71 VTAIL.n53 104.615
R119 VTAIL.n64 VTAIL.n53 104.615
R120 VTAIL.n64 VTAIL.n63 104.615
R121 VTAIL.n63 VTAIL.n57 104.615
R122 VTAIL.t4 VTAIL.n139 52.3082
R123 VTAIL.t11 VTAIL.n13 52.3082
R124 VTAIL.t7 VTAIL.n99 52.3082
R125 VTAIL.t1 VTAIL.n57 52.3082
R126 VTAIL.n87 VTAIL.n86 46.9702
R127 VTAIL.n45 VTAIL.n44 46.9702
R128 VTAIL.n1 VTAIL.n0 46.97
R129 VTAIL.n43 VTAIL.n42 46.97
R130 VTAIL.n167 VTAIL.n166 30.6338
R131 VTAIL.n41 VTAIL.n40 30.6338
R132 VTAIL.n127 VTAIL.n126 30.6338
R133 VTAIL.n85 VTAIL.n84 30.6338
R134 VTAIL.n45 VTAIL.n43 21.6945
R135 VTAIL.n167 VTAIL.n127 20.2031
R136 VTAIL.n141 VTAIL.n140 15.6677
R137 VTAIL.n15 VTAIL.n14 15.6677
R138 VTAIL.n101 VTAIL.n100 15.6677
R139 VTAIL.n59 VTAIL.n58 15.6677
R140 VTAIL.n144 VTAIL.n143 12.8005
R141 VTAIL.n18 VTAIL.n17 12.8005
R142 VTAIL.n104 VTAIL.n103 12.8005
R143 VTAIL.n62 VTAIL.n61 12.8005
R144 VTAIL.n147 VTAIL.n138 12.0247
R145 VTAIL.n21 VTAIL.n12 12.0247
R146 VTAIL.n107 VTAIL.n98 12.0247
R147 VTAIL.n65 VTAIL.n56 12.0247
R148 VTAIL.n148 VTAIL.n136 11.249
R149 VTAIL.n22 VTAIL.n10 11.249
R150 VTAIL.n108 VTAIL.n96 11.249
R151 VTAIL.n66 VTAIL.n54 11.249
R152 VTAIL.n152 VTAIL.n151 10.4732
R153 VTAIL.n26 VTAIL.n25 10.4732
R154 VTAIL.n112 VTAIL.n111 10.4732
R155 VTAIL.n70 VTAIL.n69 10.4732
R156 VTAIL.n155 VTAIL.n134 9.69747
R157 VTAIL.n29 VTAIL.n8 9.69747
R158 VTAIL.n115 VTAIL.n94 9.69747
R159 VTAIL.n73 VTAIL.n52 9.69747
R160 VTAIL.n166 VTAIL.n165 9.45567
R161 VTAIL.n40 VTAIL.n39 9.45567
R162 VTAIL.n126 VTAIL.n125 9.45567
R163 VTAIL.n84 VTAIL.n83 9.45567
R164 VTAIL.n165 VTAIL.n164 9.3005
R165 VTAIL.n159 VTAIL.n158 9.3005
R166 VTAIL.n157 VTAIL.n156 9.3005
R167 VTAIL.n134 VTAIL.n133 9.3005
R168 VTAIL.n151 VTAIL.n150 9.3005
R169 VTAIL.n149 VTAIL.n148 9.3005
R170 VTAIL.n138 VTAIL.n137 9.3005
R171 VTAIL.n143 VTAIL.n142 9.3005
R172 VTAIL.n130 VTAIL.n129 9.3005
R173 VTAIL.n39 VTAIL.n38 9.3005
R174 VTAIL.n33 VTAIL.n32 9.3005
R175 VTAIL.n31 VTAIL.n30 9.3005
R176 VTAIL.n8 VTAIL.n7 9.3005
R177 VTAIL.n25 VTAIL.n24 9.3005
R178 VTAIL.n23 VTAIL.n22 9.3005
R179 VTAIL.n12 VTAIL.n11 9.3005
R180 VTAIL.n17 VTAIL.n16 9.3005
R181 VTAIL.n4 VTAIL.n3 9.3005
R182 VTAIL.n125 VTAIL.n124 9.3005
R183 VTAIL.n90 VTAIL.n89 9.3005
R184 VTAIL.n119 VTAIL.n118 9.3005
R185 VTAIL.n117 VTAIL.n116 9.3005
R186 VTAIL.n94 VTAIL.n93 9.3005
R187 VTAIL.n111 VTAIL.n110 9.3005
R188 VTAIL.n109 VTAIL.n108 9.3005
R189 VTAIL.n98 VTAIL.n97 9.3005
R190 VTAIL.n103 VTAIL.n102 9.3005
R191 VTAIL.n83 VTAIL.n82 9.3005
R192 VTAIL.n48 VTAIL.n47 9.3005
R193 VTAIL.n77 VTAIL.n76 9.3005
R194 VTAIL.n75 VTAIL.n74 9.3005
R195 VTAIL.n52 VTAIL.n51 9.3005
R196 VTAIL.n69 VTAIL.n68 9.3005
R197 VTAIL.n67 VTAIL.n66 9.3005
R198 VTAIL.n56 VTAIL.n55 9.3005
R199 VTAIL.n61 VTAIL.n60 9.3005
R200 VTAIL.n156 VTAIL.n132 8.92171
R201 VTAIL.n30 VTAIL.n6 8.92171
R202 VTAIL.n116 VTAIL.n92 8.92171
R203 VTAIL.n74 VTAIL.n50 8.92171
R204 VTAIL.n160 VTAIL.n159 8.14595
R205 VTAIL.n34 VTAIL.n33 8.14595
R206 VTAIL.n120 VTAIL.n119 8.14595
R207 VTAIL.n78 VTAIL.n77 8.14595
R208 VTAIL.n163 VTAIL.n130 7.3702
R209 VTAIL.n166 VTAIL.n128 7.3702
R210 VTAIL.n37 VTAIL.n4 7.3702
R211 VTAIL.n40 VTAIL.n2 7.3702
R212 VTAIL.n126 VTAIL.n88 7.3702
R213 VTAIL.n123 VTAIL.n90 7.3702
R214 VTAIL.n84 VTAIL.n46 7.3702
R215 VTAIL.n81 VTAIL.n48 7.3702
R216 VTAIL.n164 VTAIL.n163 6.59444
R217 VTAIL.n164 VTAIL.n128 6.59444
R218 VTAIL.n38 VTAIL.n37 6.59444
R219 VTAIL.n38 VTAIL.n2 6.59444
R220 VTAIL.n124 VTAIL.n88 6.59444
R221 VTAIL.n124 VTAIL.n123 6.59444
R222 VTAIL.n82 VTAIL.n46 6.59444
R223 VTAIL.n82 VTAIL.n81 6.59444
R224 VTAIL.n160 VTAIL.n130 5.81868
R225 VTAIL.n34 VTAIL.n4 5.81868
R226 VTAIL.n120 VTAIL.n90 5.81868
R227 VTAIL.n78 VTAIL.n48 5.81868
R228 VTAIL.n159 VTAIL.n132 5.04292
R229 VTAIL.n33 VTAIL.n6 5.04292
R230 VTAIL.n119 VTAIL.n92 5.04292
R231 VTAIL.n77 VTAIL.n50 5.04292
R232 VTAIL.n102 VTAIL.n101 4.38565
R233 VTAIL.n60 VTAIL.n59 4.38565
R234 VTAIL.n142 VTAIL.n141 4.38565
R235 VTAIL.n16 VTAIL.n15 4.38565
R236 VTAIL.n156 VTAIL.n155 4.26717
R237 VTAIL.n30 VTAIL.n29 4.26717
R238 VTAIL.n116 VTAIL.n115 4.26717
R239 VTAIL.n74 VTAIL.n73 4.26717
R240 VTAIL.n152 VTAIL.n134 3.49141
R241 VTAIL.n26 VTAIL.n8 3.49141
R242 VTAIL.n112 VTAIL.n94 3.49141
R243 VTAIL.n70 VTAIL.n52 3.49141
R244 VTAIL.n151 VTAIL.n136 2.71565
R245 VTAIL.n25 VTAIL.n10 2.71565
R246 VTAIL.n111 VTAIL.n96 2.71565
R247 VTAIL.n69 VTAIL.n54 2.71565
R248 VTAIL.n0 VTAIL.t5 2.69072
R249 VTAIL.n0 VTAIL.t0 2.69072
R250 VTAIL.n42 VTAIL.t6 2.69072
R251 VTAIL.n42 VTAIL.t8 2.69072
R252 VTAIL.n86 VTAIL.t10 2.69072
R253 VTAIL.n86 VTAIL.t9 2.69072
R254 VTAIL.n44 VTAIL.t2 2.69072
R255 VTAIL.n44 VTAIL.t3 2.69072
R256 VTAIL.n148 VTAIL.n147 1.93989
R257 VTAIL.n22 VTAIL.n21 1.93989
R258 VTAIL.n108 VTAIL.n107 1.93989
R259 VTAIL.n66 VTAIL.n65 1.93989
R260 VTAIL.n85 VTAIL.n45 1.49188
R261 VTAIL.n127 VTAIL.n87 1.49188
R262 VTAIL.n43 VTAIL.n41 1.49188
R263 VTAIL.n87 VTAIL.n85 1.21602
R264 VTAIL.n41 VTAIL.n1 1.21602
R265 VTAIL.n144 VTAIL.n138 1.16414
R266 VTAIL.n18 VTAIL.n12 1.16414
R267 VTAIL.n104 VTAIL.n98 1.16414
R268 VTAIL.n62 VTAIL.n56 1.16414
R269 VTAIL VTAIL.n167 1.06084
R270 VTAIL VTAIL.n1 0.431534
R271 VTAIL.n143 VTAIL.n140 0.388379
R272 VTAIL.n17 VTAIL.n14 0.388379
R273 VTAIL.n103 VTAIL.n100 0.388379
R274 VTAIL.n61 VTAIL.n58 0.388379
R275 VTAIL.n142 VTAIL.n137 0.155672
R276 VTAIL.n149 VTAIL.n137 0.155672
R277 VTAIL.n150 VTAIL.n149 0.155672
R278 VTAIL.n150 VTAIL.n133 0.155672
R279 VTAIL.n157 VTAIL.n133 0.155672
R280 VTAIL.n158 VTAIL.n157 0.155672
R281 VTAIL.n158 VTAIL.n129 0.155672
R282 VTAIL.n165 VTAIL.n129 0.155672
R283 VTAIL.n16 VTAIL.n11 0.155672
R284 VTAIL.n23 VTAIL.n11 0.155672
R285 VTAIL.n24 VTAIL.n23 0.155672
R286 VTAIL.n24 VTAIL.n7 0.155672
R287 VTAIL.n31 VTAIL.n7 0.155672
R288 VTAIL.n32 VTAIL.n31 0.155672
R289 VTAIL.n32 VTAIL.n3 0.155672
R290 VTAIL.n39 VTAIL.n3 0.155672
R291 VTAIL.n125 VTAIL.n89 0.155672
R292 VTAIL.n118 VTAIL.n89 0.155672
R293 VTAIL.n118 VTAIL.n117 0.155672
R294 VTAIL.n117 VTAIL.n93 0.155672
R295 VTAIL.n110 VTAIL.n93 0.155672
R296 VTAIL.n110 VTAIL.n109 0.155672
R297 VTAIL.n109 VTAIL.n97 0.155672
R298 VTAIL.n102 VTAIL.n97 0.155672
R299 VTAIL.n83 VTAIL.n47 0.155672
R300 VTAIL.n76 VTAIL.n47 0.155672
R301 VTAIL.n76 VTAIL.n75 0.155672
R302 VTAIL.n75 VTAIL.n51 0.155672
R303 VTAIL.n68 VTAIL.n51 0.155672
R304 VTAIL.n68 VTAIL.n67 0.155672
R305 VTAIL.n67 VTAIL.n55 0.155672
R306 VTAIL.n60 VTAIL.n55 0.155672
R307 VDD1.n34 VDD1.n0 289.615
R308 VDD1.n73 VDD1.n39 289.615
R309 VDD1.n35 VDD1.n34 185
R310 VDD1.n33 VDD1.n32 185
R311 VDD1.n4 VDD1.n3 185
R312 VDD1.n27 VDD1.n26 185
R313 VDD1.n25 VDD1.n24 185
R314 VDD1.n8 VDD1.n7 185
R315 VDD1.n19 VDD1.n18 185
R316 VDD1.n17 VDD1.n16 185
R317 VDD1.n12 VDD1.n11 185
R318 VDD1.n51 VDD1.n50 185
R319 VDD1.n56 VDD1.n55 185
R320 VDD1.n58 VDD1.n57 185
R321 VDD1.n47 VDD1.n46 185
R322 VDD1.n64 VDD1.n63 185
R323 VDD1.n66 VDD1.n65 185
R324 VDD1.n43 VDD1.n42 185
R325 VDD1.n72 VDD1.n71 185
R326 VDD1.n74 VDD1.n73 185
R327 VDD1.n13 VDD1.t5 147.659
R328 VDD1.n52 VDD1.t2 147.659
R329 VDD1.n34 VDD1.n33 104.615
R330 VDD1.n33 VDD1.n3 104.615
R331 VDD1.n26 VDD1.n3 104.615
R332 VDD1.n26 VDD1.n25 104.615
R333 VDD1.n25 VDD1.n7 104.615
R334 VDD1.n18 VDD1.n7 104.615
R335 VDD1.n18 VDD1.n17 104.615
R336 VDD1.n17 VDD1.n11 104.615
R337 VDD1.n56 VDD1.n50 104.615
R338 VDD1.n57 VDD1.n56 104.615
R339 VDD1.n57 VDD1.n46 104.615
R340 VDD1.n64 VDD1.n46 104.615
R341 VDD1.n65 VDD1.n64 104.615
R342 VDD1.n65 VDD1.n42 104.615
R343 VDD1.n72 VDD1.n42 104.615
R344 VDD1.n73 VDD1.n72 104.615
R345 VDD1.n79 VDD1.n78 63.9663
R346 VDD1.n81 VDD1.n80 63.6488
R347 VDD1.t5 VDD1.n11 52.3082
R348 VDD1.t2 VDD1.n50 52.3082
R349 VDD1 VDD1.n38 48.4893
R350 VDD1.n79 VDD1.n77 48.3758
R351 VDD1.n81 VDD1.n79 36.2358
R352 VDD1.n13 VDD1.n12 15.6677
R353 VDD1.n52 VDD1.n51 15.6677
R354 VDD1.n16 VDD1.n15 12.8005
R355 VDD1.n55 VDD1.n54 12.8005
R356 VDD1.n19 VDD1.n10 12.0247
R357 VDD1.n58 VDD1.n49 12.0247
R358 VDD1.n20 VDD1.n8 11.249
R359 VDD1.n59 VDD1.n47 11.249
R360 VDD1.n24 VDD1.n23 10.4732
R361 VDD1.n63 VDD1.n62 10.4732
R362 VDD1.n27 VDD1.n6 9.69747
R363 VDD1.n66 VDD1.n45 9.69747
R364 VDD1.n38 VDD1.n37 9.45567
R365 VDD1.n77 VDD1.n76 9.45567
R366 VDD1.n37 VDD1.n36 9.3005
R367 VDD1.n2 VDD1.n1 9.3005
R368 VDD1.n31 VDD1.n30 9.3005
R369 VDD1.n29 VDD1.n28 9.3005
R370 VDD1.n6 VDD1.n5 9.3005
R371 VDD1.n23 VDD1.n22 9.3005
R372 VDD1.n21 VDD1.n20 9.3005
R373 VDD1.n10 VDD1.n9 9.3005
R374 VDD1.n15 VDD1.n14 9.3005
R375 VDD1.n76 VDD1.n75 9.3005
R376 VDD1.n70 VDD1.n69 9.3005
R377 VDD1.n68 VDD1.n67 9.3005
R378 VDD1.n45 VDD1.n44 9.3005
R379 VDD1.n62 VDD1.n61 9.3005
R380 VDD1.n60 VDD1.n59 9.3005
R381 VDD1.n49 VDD1.n48 9.3005
R382 VDD1.n54 VDD1.n53 9.3005
R383 VDD1.n41 VDD1.n40 9.3005
R384 VDD1.n28 VDD1.n4 8.92171
R385 VDD1.n67 VDD1.n43 8.92171
R386 VDD1.n32 VDD1.n31 8.14595
R387 VDD1.n71 VDD1.n70 8.14595
R388 VDD1.n38 VDD1.n0 7.3702
R389 VDD1.n35 VDD1.n2 7.3702
R390 VDD1.n74 VDD1.n41 7.3702
R391 VDD1.n77 VDD1.n39 7.3702
R392 VDD1.n36 VDD1.n0 6.59444
R393 VDD1.n36 VDD1.n35 6.59444
R394 VDD1.n75 VDD1.n74 6.59444
R395 VDD1.n75 VDD1.n39 6.59444
R396 VDD1.n32 VDD1.n2 5.81868
R397 VDD1.n71 VDD1.n41 5.81868
R398 VDD1.n31 VDD1.n4 5.04292
R399 VDD1.n70 VDD1.n43 5.04292
R400 VDD1.n14 VDD1.n13 4.38565
R401 VDD1.n53 VDD1.n52 4.38565
R402 VDD1.n28 VDD1.n27 4.26717
R403 VDD1.n67 VDD1.n66 4.26717
R404 VDD1.n24 VDD1.n6 3.49141
R405 VDD1.n63 VDD1.n45 3.49141
R406 VDD1.n23 VDD1.n8 2.71565
R407 VDD1.n62 VDD1.n47 2.71565
R408 VDD1.n80 VDD1.t1 2.69072
R409 VDD1.n80 VDD1.t0 2.69072
R410 VDD1.n78 VDD1.t4 2.69072
R411 VDD1.n78 VDD1.t3 2.69072
R412 VDD1.n20 VDD1.n19 1.93989
R413 VDD1.n59 VDD1.n58 1.93989
R414 VDD1.n16 VDD1.n10 1.16414
R415 VDD1.n55 VDD1.n49 1.16414
R416 VDD1.n15 VDD1.n12 0.388379
R417 VDD1.n54 VDD1.n51 0.388379
R418 VDD1 VDD1.n81 0.315155
R419 VDD1.n37 VDD1.n1 0.155672
R420 VDD1.n30 VDD1.n1 0.155672
R421 VDD1.n30 VDD1.n29 0.155672
R422 VDD1.n29 VDD1.n5 0.155672
R423 VDD1.n22 VDD1.n5 0.155672
R424 VDD1.n22 VDD1.n21 0.155672
R425 VDD1.n21 VDD1.n9 0.155672
R426 VDD1.n14 VDD1.n9 0.155672
R427 VDD1.n53 VDD1.n48 0.155672
R428 VDD1.n60 VDD1.n48 0.155672
R429 VDD1.n61 VDD1.n60 0.155672
R430 VDD1.n61 VDD1.n44 0.155672
R431 VDD1.n68 VDD1.n44 0.155672
R432 VDD1.n69 VDD1.n68 0.155672
R433 VDD1.n69 VDD1.n40 0.155672
R434 VDD1.n76 VDD1.n40 0.155672
R435 B.n569 B.n568 585
R436 B.n220 B.n87 585
R437 B.n219 B.n218 585
R438 B.n217 B.n216 585
R439 B.n215 B.n214 585
R440 B.n213 B.n212 585
R441 B.n211 B.n210 585
R442 B.n209 B.n208 585
R443 B.n207 B.n206 585
R444 B.n205 B.n204 585
R445 B.n203 B.n202 585
R446 B.n201 B.n200 585
R447 B.n199 B.n198 585
R448 B.n197 B.n196 585
R449 B.n195 B.n194 585
R450 B.n193 B.n192 585
R451 B.n191 B.n190 585
R452 B.n189 B.n188 585
R453 B.n187 B.n186 585
R454 B.n185 B.n184 585
R455 B.n183 B.n182 585
R456 B.n181 B.n180 585
R457 B.n179 B.n178 585
R458 B.n177 B.n176 585
R459 B.n175 B.n174 585
R460 B.n173 B.n172 585
R461 B.n171 B.n170 585
R462 B.n169 B.n168 585
R463 B.n167 B.n166 585
R464 B.n165 B.n164 585
R465 B.n163 B.n162 585
R466 B.n161 B.n160 585
R467 B.n159 B.n158 585
R468 B.n157 B.n156 585
R469 B.n155 B.n154 585
R470 B.n153 B.n152 585
R471 B.n151 B.n150 585
R472 B.n149 B.n148 585
R473 B.n147 B.n146 585
R474 B.n145 B.n144 585
R475 B.n143 B.n142 585
R476 B.n141 B.n140 585
R477 B.n139 B.n138 585
R478 B.n137 B.n136 585
R479 B.n135 B.n134 585
R480 B.n133 B.n132 585
R481 B.n131 B.n130 585
R482 B.n129 B.n128 585
R483 B.n127 B.n126 585
R484 B.n125 B.n124 585
R485 B.n123 B.n122 585
R486 B.n121 B.n120 585
R487 B.n119 B.n118 585
R488 B.n117 B.n116 585
R489 B.n115 B.n114 585
R490 B.n113 B.n112 585
R491 B.n111 B.n110 585
R492 B.n109 B.n108 585
R493 B.n107 B.n106 585
R494 B.n105 B.n104 585
R495 B.n103 B.n102 585
R496 B.n101 B.n100 585
R497 B.n99 B.n98 585
R498 B.n97 B.n96 585
R499 B.n95 B.n94 585
R500 B.n53 B.n52 585
R501 B.n567 B.n54 585
R502 B.n572 B.n54 585
R503 B.n566 B.n565 585
R504 B.n565 B.n50 585
R505 B.n564 B.n49 585
R506 B.n578 B.n49 585
R507 B.n563 B.n48 585
R508 B.n579 B.n48 585
R509 B.n562 B.n47 585
R510 B.n580 B.n47 585
R511 B.n561 B.n560 585
R512 B.n560 B.n46 585
R513 B.n559 B.n42 585
R514 B.n586 B.n42 585
R515 B.n558 B.n41 585
R516 B.n587 B.n41 585
R517 B.n557 B.n40 585
R518 B.n588 B.n40 585
R519 B.n556 B.n555 585
R520 B.n555 B.n36 585
R521 B.n554 B.n35 585
R522 B.n594 B.n35 585
R523 B.n553 B.n34 585
R524 B.n595 B.n34 585
R525 B.n552 B.n33 585
R526 B.n596 B.n33 585
R527 B.n551 B.n550 585
R528 B.n550 B.n29 585
R529 B.n549 B.n28 585
R530 B.n602 B.n28 585
R531 B.n548 B.n27 585
R532 B.n603 B.n27 585
R533 B.n547 B.n26 585
R534 B.n604 B.n26 585
R535 B.n546 B.n545 585
R536 B.n545 B.n22 585
R537 B.n544 B.n21 585
R538 B.n610 B.n21 585
R539 B.n543 B.n20 585
R540 B.n611 B.n20 585
R541 B.n542 B.n19 585
R542 B.n612 B.n19 585
R543 B.n541 B.n540 585
R544 B.n540 B.n15 585
R545 B.n539 B.n14 585
R546 B.n618 B.n14 585
R547 B.n538 B.n13 585
R548 B.n619 B.n13 585
R549 B.n537 B.n12 585
R550 B.n620 B.n12 585
R551 B.n536 B.n535 585
R552 B.n535 B.n534 585
R553 B.n533 B.n532 585
R554 B.n533 B.n8 585
R555 B.n531 B.n7 585
R556 B.n627 B.n7 585
R557 B.n530 B.n6 585
R558 B.n628 B.n6 585
R559 B.n529 B.n5 585
R560 B.n629 B.n5 585
R561 B.n528 B.n527 585
R562 B.n527 B.n4 585
R563 B.n526 B.n221 585
R564 B.n526 B.n525 585
R565 B.n516 B.n222 585
R566 B.n223 B.n222 585
R567 B.n518 B.n517 585
R568 B.n519 B.n518 585
R569 B.n515 B.n228 585
R570 B.n228 B.n227 585
R571 B.n514 B.n513 585
R572 B.n513 B.n512 585
R573 B.n230 B.n229 585
R574 B.n231 B.n230 585
R575 B.n505 B.n504 585
R576 B.n506 B.n505 585
R577 B.n503 B.n235 585
R578 B.n239 B.n235 585
R579 B.n502 B.n501 585
R580 B.n501 B.n500 585
R581 B.n237 B.n236 585
R582 B.n238 B.n237 585
R583 B.n493 B.n492 585
R584 B.n494 B.n493 585
R585 B.n491 B.n244 585
R586 B.n244 B.n243 585
R587 B.n490 B.n489 585
R588 B.n489 B.n488 585
R589 B.n246 B.n245 585
R590 B.n247 B.n246 585
R591 B.n481 B.n480 585
R592 B.n482 B.n481 585
R593 B.n479 B.n252 585
R594 B.n252 B.n251 585
R595 B.n478 B.n477 585
R596 B.n477 B.n476 585
R597 B.n254 B.n253 585
R598 B.n255 B.n254 585
R599 B.n469 B.n468 585
R600 B.n470 B.n469 585
R601 B.n467 B.n260 585
R602 B.n260 B.n259 585
R603 B.n466 B.n465 585
R604 B.n465 B.n464 585
R605 B.n262 B.n261 585
R606 B.n457 B.n262 585
R607 B.n456 B.n455 585
R608 B.n458 B.n456 585
R609 B.n454 B.n267 585
R610 B.n267 B.n266 585
R611 B.n453 B.n452 585
R612 B.n452 B.n451 585
R613 B.n269 B.n268 585
R614 B.n270 B.n269 585
R615 B.n444 B.n443 585
R616 B.n445 B.n444 585
R617 B.n273 B.n272 585
R618 B.n312 B.n310 585
R619 B.n313 B.n309 585
R620 B.n313 B.n274 585
R621 B.n316 B.n315 585
R622 B.n317 B.n308 585
R623 B.n319 B.n318 585
R624 B.n321 B.n307 585
R625 B.n324 B.n323 585
R626 B.n325 B.n306 585
R627 B.n327 B.n326 585
R628 B.n329 B.n305 585
R629 B.n332 B.n331 585
R630 B.n333 B.n304 585
R631 B.n335 B.n334 585
R632 B.n337 B.n303 585
R633 B.n340 B.n339 585
R634 B.n341 B.n302 585
R635 B.n343 B.n342 585
R636 B.n345 B.n301 585
R637 B.n348 B.n347 585
R638 B.n349 B.n300 585
R639 B.n351 B.n350 585
R640 B.n353 B.n299 585
R641 B.n356 B.n355 585
R642 B.n357 B.n298 585
R643 B.n359 B.n358 585
R644 B.n361 B.n297 585
R645 B.n364 B.n363 585
R646 B.n366 B.n294 585
R647 B.n368 B.n367 585
R648 B.n370 B.n293 585
R649 B.n373 B.n372 585
R650 B.n374 B.n292 585
R651 B.n376 B.n375 585
R652 B.n378 B.n291 585
R653 B.n381 B.n380 585
R654 B.n382 B.n290 585
R655 B.n387 B.n386 585
R656 B.n389 B.n289 585
R657 B.n392 B.n391 585
R658 B.n393 B.n288 585
R659 B.n395 B.n394 585
R660 B.n397 B.n287 585
R661 B.n400 B.n399 585
R662 B.n401 B.n286 585
R663 B.n403 B.n402 585
R664 B.n405 B.n285 585
R665 B.n408 B.n407 585
R666 B.n409 B.n284 585
R667 B.n411 B.n410 585
R668 B.n413 B.n283 585
R669 B.n416 B.n415 585
R670 B.n417 B.n282 585
R671 B.n419 B.n418 585
R672 B.n421 B.n281 585
R673 B.n424 B.n423 585
R674 B.n425 B.n280 585
R675 B.n427 B.n426 585
R676 B.n429 B.n279 585
R677 B.n432 B.n431 585
R678 B.n433 B.n278 585
R679 B.n435 B.n434 585
R680 B.n437 B.n277 585
R681 B.n438 B.n276 585
R682 B.n441 B.n440 585
R683 B.n442 B.n275 585
R684 B.n275 B.n274 585
R685 B.n447 B.n446 585
R686 B.n446 B.n445 585
R687 B.n448 B.n271 585
R688 B.n271 B.n270 585
R689 B.n450 B.n449 585
R690 B.n451 B.n450 585
R691 B.n265 B.n264 585
R692 B.n266 B.n265 585
R693 B.n460 B.n459 585
R694 B.n459 B.n458 585
R695 B.n461 B.n263 585
R696 B.n457 B.n263 585
R697 B.n463 B.n462 585
R698 B.n464 B.n463 585
R699 B.n258 B.n257 585
R700 B.n259 B.n258 585
R701 B.n472 B.n471 585
R702 B.n471 B.n470 585
R703 B.n473 B.n256 585
R704 B.n256 B.n255 585
R705 B.n475 B.n474 585
R706 B.n476 B.n475 585
R707 B.n250 B.n249 585
R708 B.n251 B.n250 585
R709 B.n484 B.n483 585
R710 B.n483 B.n482 585
R711 B.n485 B.n248 585
R712 B.n248 B.n247 585
R713 B.n487 B.n486 585
R714 B.n488 B.n487 585
R715 B.n242 B.n241 585
R716 B.n243 B.n242 585
R717 B.n496 B.n495 585
R718 B.n495 B.n494 585
R719 B.n497 B.n240 585
R720 B.n240 B.n238 585
R721 B.n499 B.n498 585
R722 B.n500 B.n499 585
R723 B.n234 B.n233 585
R724 B.n239 B.n234 585
R725 B.n508 B.n507 585
R726 B.n507 B.n506 585
R727 B.n509 B.n232 585
R728 B.n232 B.n231 585
R729 B.n511 B.n510 585
R730 B.n512 B.n511 585
R731 B.n226 B.n225 585
R732 B.n227 B.n226 585
R733 B.n521 B.n520 585
R734 B.n520 B.n519 585
R735 B.n522 B.n224 585
R736 B.n224 B.n223 585
R737 B.n524 B.n523 585
R738 B.n525 B.n524 585
R739 B.n3 B.n0 585
R740 B.n4 B.n3 585
R741 B.n626 B.n1 585
R742 B.n627 B.n626 585
R743 B.n625 B.n624 585
R744 B.n625 B.n8 585
R745 B.n623 B.n9 585
R746 B.n534 B.n9 585
R747 B.n622 B.n621 585
R748 B.n621 B.n620 585
R749 B.n11 B.n10 585
R750 B.n619 B.n11 585
R751 B.n617 B.n616 585
R752 B.n618 B.n617 585
R753 B.n615 B.n16 585
R754 B.n16 B.n15 585
R755 B.n614 B.n613 585
R756 B.n613 B.n612 585
R757 B.n18 B.n17 585
R758 B.n611 B.n18 585
R759 B.n609 B.n608 585
R760 B.n610 B.n609 585
R761 B.n607 B.n23 585
R762 B.n23 B.n22 585
R763 B.n606 B.n605 585
R764 B.n605 B.n604 585
R765 B.n25 B.n24 585
R766 B.n603 B.n25 585
R767 B.n601 B.n600 585
R768 B.n602 B.n601 585
R769 B.n599 B.n30 585
R770 B.n30 B.n29 585
R771 B.n598 B.n597 585
R772 B.n597 B.n596 585
R773 B.n32 B.n31 585
R774 B.n595 B.n32 585
R775 B.n593 B.n592 585
R776 B.n594 B.n593 585
R777 B.n591 B.n37 585
R778 B.n37 B.n36 585
R779 B.n590 B.n589 585
R780 B.n589 B.n588 585
R781 B.n39 B.n38 585
R782 B.n587 B.n39 585
R783 B.n585 B.n584 585
R784 B.n586 B.n585 585
R785 B.n583 B.n43 585
R786 B.n46 B.n43 585
R787 B.n582 B.n581 585
R788 B.n581 B.n580 585
R789 B.n45 B.n44 585
R790 B.n579 B.n45 585
R791 B.n577 B.n576 585
R792 B.n578 B.n577 585
R793 B.n575 B.n51 585
R794 B.n51 B.n50 585
R795 B.n574 B.n573 585
R796 B.n573 B.n572 585
R797 B.n630 B.n629 585
R798 B.n628 B.n2 585
R799 B.n573 B.n53 454.062
R800 B.n569 B.n54 454.062
R801 B.n444 B.n275 454.062
R802 B.n446 B.n273 454.062
R803 B.n91 B.t17 331.745
R804 B.n88 B.t13 331.745
R805 B.n383 B.t10 331.745
R806 B.n295 B.t6 331.745
R807 B.n571 B.n570 256.663
R808 B.n571 B.n86 256.663
R809 B.n571 B.n85 256.663
R810 B.n571 B.n84 256.663
R811 B.n571 B.n83 256.663
R812 B.n571 B.n82 256.663
R813 B.n571 B.n81 256.663
R814 B.n571 B.n80 256.663
R815 B.n571 B.n79 256.663
R816 B.n571 B.n78 256.663
R817 B.n571 B.n77 256.663
R818 B.n571 B.n76 256.663
R819 B.n571 B.n75 256.663
R820 B.n571 B.n74 256.663
R821 B.n571 B.n73 256.663
R822 B.n571 B.n72 256.663
R823 B.n571 B.n71 256.663
R824 B.n571 B.n70 256.663
R825 B.n571 B.n69 256.663
R826 B.n571 B.n68 256.663
R827 B.n571 B.n67 256.663
R828 B.n571 B.n66 256.663
R829 B.n571 B.n65 256.663
R830 B.n571 B.n64 256.663
R831 B.n571 B.n63 256.663
R832 B.n571 B.n62 256.663
R833 B.n571 B.n61 256.663
R834 B.n571 B.n60 256.663
R835 B.n571 B.n59 256.663
R836 B.n571 B.n58 256.663
R837 B.n571 B.n57 256.663
R838 B.n571 B.n56 256.663
R839 B.n571 B.n55 256.663
R840 B.n311 B.n274 256.663
R841 B.n314 B.n274 256.663
R842 B.n320 B.n274 256.663
R843 B.n322 B.n274 256.663
R844 B.n328 B.n274 256.663
R845 B.n330 B.n274 256.663
R846 B.n336 B.n274 256.663
R847 B.n338 B.n274 256.663
R848 B.n344 B.n274 256.663
R849 B.n346 B.n274 256.663
R850 B.n352 B.n274 256.663
R851 B.n354 B.n274 256.663
R852 B.n360 B.n274 256.663
R853 B.n362 B.n274 256.663
R854 B.n369 B.n274 256.663
R855 B.n371 B.n274 256.663
R856 B.n377 B.n274 256.663
R857 B.n379 B.n274 256.663
R858 B.n388 B.n274 256.663
R859 B.n390 B.n274 256.663
R860 B.n396 B.n274 256.663
R861 B.n398 B.n274 256.663
R862 B.n404 B.n274 256.663
R863 B.n406 B.n274 256.663
R864 B.n412 B.n274 256.663
R865 B.n414 B.n274 256.663
R866 B.n420 B.n274 256.663
R867 B.n422 B.n274 256.663
R868 B.n428 B.n274 256.663
R869 B.n430 B.n274 256.663
R870 B.n436 B.n274 256.663
R871 B.n439 B.n274 256.663
R872 B.n632 B.n631 256.663
R873 B.n88 B.t15 235.913
R874 B.n383 B.t12 235.913
R875 B.n91 B.t18 235.913
R876 B.n295 B.t9 235.913
R877 B.n89 B.t16 202.362
R878 B.n384 B.t11 202.362
R879 B.n92 B.t19 202.362
R880 B.n296 B.t8 202.362
R881 B.n96 B.n95 163.367
R882 B.n100 B.n99 163.367
R883 B.n104 B.n103 163.367
R884 B.n108 B.n107 163.367
R885 B.n112 B.n111 163.367
R886 B.n116 B.n115 163.367
R887 B.n120 B.n119 163.367
R888 B.n124 B.n123 163.367
R889 B.n128 B.n127 163.367
R890 B.n132 B.n131 163.367
R891 B.n136 B.n135 163.367
R892 B.n140 B.n139 163.367
R893 B.n144 B.n143 163.367
R894 B.n148 B.n147 163.367
R895 B.n152 B.n151 163.367
R896 B.n156 B.n155 163.367
R897 B.n160 B.n159 163.367
R898 B.n164 B.n163 163.367
R899 B.n168 B.n167 163.367
R900 B.n172 B.n171 163.367
R901 B.n176 B.n175 163.367
R902 B.n180 B.n179 163.367
R903 B.n184 B.n183 163.367
R904 B.n188 B.n187 163.367
R905 B.n192 B.n191 163.367
R906 B.n196 B.n195 163.367
R907 B.n200 B.n199 163.367
R908 B.n204 B.n203 163.367
R909 B.n208 B.n207 163.367
R910 B.n212 B.n211 163.367
R911 B.n216 B.n215 163.367
R912 B.n218 B.n87 163.367
R913 B.n444 B.n269 163.367
R914 B.n452 B.n269 163.367
R915 B.n452 B.n267 163.367
R916 B.n456 B.n267 163.367
R917 B.n456 B.n262 163.367
R918 B.n465 B.n262 163.367
R919 B.n465 B.n260 163.367
R920 B.n469 B.n260 163.367
R921 B.n469 B.n254 163.367
R922 B.n477 B.n254 163.367
R923 B.n477 B.n252 163.367
R924 B.n481 B.n252 163.367
R925 B.n481 B.n246 163.367
R926 B.n489 B.n246 163.367
R927 B.n489 B.n244 163.367
R928 B.n493 B.n244 163.367
R929 B.n493 B.n237 163.367
R930 B.n501 B.n237 163.367
R931 B.n501 B.n235 163.367
R932 B.n505 B.n235 163.367
R933 B.n505 B.n230 163.367
R934 B.n513 B.n230 163.367
R935 B.n513 B.n228 163.367
R936 B.n518 B.n228 163.367
R937 B.n518 B.n222 163.367
R938 B.n526 B.n222 163.367
R939 B.n527 B.n526 163.367
R940 B.n527 B.n5 163.367
R941 B.n6 B.n5 163.367
R942 B.n7 B.n6 163.367
R943 B.n533 B.n7 163.367
R944 B.n535 B.n533 163.367
R945 B.n535 B.n12 163.367
R946 B.n13 B.n12 163.367
R947 B.n14 B.n13 163.367
R948 B.n540 B.n14 163.367
R949 B.n540 B.n19 163.367
R950 B.n20 B.n19 163.367
R951 B.n21 B.n20 163.367
R952 B.n545 B.n21 163.367
R953 B.n545 B.n26 163.367
R954 B.n27 B.n26 163.367
R955 B.n28 B.n27 163.367
R956 B.n550 B.n28 163.367
R957 B.n550 B.n33 163.367
R958 B.n34 B.n33 163.367
R959 B.n35 B.n34 163.367
R960 B.n555 B.n35 163.367
R961 B.n555 B.n40 163.367
R962 B.n41 B.n40 163.367
R963 B.n42 B.n41 163.367
R964 B.n560 B.n42 163.367
R965 B.n560 B.n47 163.367
R966 B.n48 B.n47 163.367
R967 B.n49 B.n48 163.367
R968 B.n565 B.n49 163.367
R969 B.n565 B.n54 163.367
R970 B.n313 B.n312 163.367
R971 B.n315 B.n313 163.367
R972 B.n319 B.n308 163.367
R973 B.n323 B.n321 163.367
R974 B.n327 B.n306 163.367
R975 B.n331 B.n329 163.367
R976 B.n335 B.n304 163.367
R977 B.n339 B.n337 163.367
R978 B.n343 B.n302 163.367
R979 B.n347 B.n345 163.367
R980 B.n351 B.n300 163.367
R981 B.n355 B.n353 163.367
R982 B.n359 B.n298 163.367
R983 B.n363 B.n361 163.367
R984 B.n368 B.n294 163.367
R985 B.n372 B.n370 163.367
R986 B.n376 B.n292 163.367
R987 B.n380 B.n378 163.367
R988 B.n387 B.n290 163.367
R989 B.n391 B.n389 163.367
R990 B.n395 B.n288 163.367
R991 B.n399 B.n397 163.367
R992 B.n403 B.n286 163.367
R993 B.n407 B.n405 163.367
R994 B.n411 B.n284 163.367
R995 B.n415 B.n413 163.367
R996 B.n419 B.n282 163.367
R997 B.n423 B.n421 163.367
R998 B.n427 B.n280 163.367
R999 B.n431 B.n429 163.367
R1000 B.n435 B.n278 163.367
R1001 B.n438 B.n437 163.367
R1002 B.n440 B.n275 163.367
R1003 B.n446 B.n271 163.367
R1004 B.n450 B.n271 163.367
R1005 B.n450 B.n265 163.367
R1006 B.n459 B.n265 163.367
R1007 B.n459 B.n263 163.367
R1008 B.n463 B.n263 163.367
R1009 B.n463 B.n258 163.367
R1010 B.n471 B.n258 163.367
R1011 B.n471 B.n256 163.367
R1012 B.n475 B.n256 163.367
R1013 B.n475 B.n250 163.367
R1014 B.n483 B.n250 163.367
R1015 B.n483 B.n248 163.367
R1016 B.n487 B.n248 163.367
R1017 B.n487 B.n242 163.367
R1018 B.n495 B.n242 163.367
R1019 B.n495 B.n240 163.367
R1020 B.n499 B.n240 163.367
R1021 B.n499 B.n234 163.367
R1022 B.n507 B.n234 163.367
R1023 B.n507 B.n232 163.367
R1024 B.n511 B.n232 163.367
R1025 B.n511 B.n226 163.367
R1026 B.n520 B.n226 163.367
R1027 B.n520 B.n224 163.367
R1028 B.n524 B.n224 163.367
R1029 B.n524 B.n3 163.367
R1030 B.n630 B.n3 163.367
R1031 B.n626 B.n2 163.367
R1032 B.n626 B.n625 163.367
R1033 B.n625 B.n9 163.367
R1034 B.n621 B.n9 163.367
R1035 B.n621 B.n11 163.367
R1036 B.n617 B.n11 163.367
R1037 B.n617 B.n16 163.367
R1038 B.n613 B.n16 163.367
R1039 B.n613 B.n18 163.367
R1040 B.n609 B.n18 163.367
R1041 B.n609 B.n23 163.367
R1042 B.n605 B.n23 163.367
R1043 B.n605 B.n25 163.367
R1044 B.n601 B.n25 163.367
R1045 B.n601 B.n30 163.367
R1046 B.n597 B.n30 163.367
R1047 B.n597 B.n32 163.367
R1048 B.n593 B.n32 163.367
R1049 B.n593 B.n37 163.367
R1050 B.n589 B.n37 163.367
R1051 B.n589 B.n39 163.367
R1052 B.n585 B.n39 163.367
R1053 B.n585 B.n43 163.367
R1054 B.n581 B.n43 163.367
R1055 B.n581 B.n45 163.367
R1056 B.n577 B.n45 163.367
R1057 B.n577 B.n51 163.367
R1058 B.n573 B.n51 163.367
R1059 B.n445 B.n274 105.343
R1060 B.n572 B.n571 105.343
R1061 B.n55 B.n53 71.676
R1062 B.n96 B.n56 71.676
R1063 B.n100 B.n57 71.676
R1064 B.n104 B.n58 71.676
R1065 B.n108 B.n59 71.676
R1066 B.n112 B.n60 71.676
R1067 B.n116 B.n61 71.676
R1068 B.n120 B.n62 71.676
R1069 B.n124 B.n63 71.676
R1070 B.n128 B.n64 71.676
R1071 B.n132 B.n65 71.676
R1072 B.n136 B.n66 71.676
R1073 B.n140 B.n67 71.676
R1074 B.n144 B.n68 71.676
R1075 B.n148 B.n69 71.676
R1076 B.n152 B.n70 71.676
R1077 B.n156 B.n71 71.676
R1078 B.n160 B.n72 71.676
R1079 B.n164 B.n73 71.676
R1080 B.n168 B.n74 71.676
R1081 B.n172 B.n75 71.676
R1082 B.n176 B.n76 71.676
R1083 B.n180 B.n77 71.676
R1084 B.n184 B.n78 71.676
R1085 B.n188 B.n79 71.676
R1086 B.n192 B.n80 71.676
R1087 B.n196 B.n81 71.676
R1088 B.n200 B.n82 71.676
R1089 B.n204 B.n83 71.676
R1090 B.n208 B.n84 71.676
R1091 B.n212 B.n85 71.676
R1092 B.n216 B.n86 71.676
R1093 B.n570 B.n87 71.676
R1094 B.n570 B.n569 71.676
R1095 B.n218 B.n86 71.676
R1096 B.n215 B.n85 71.676
R1097 B.n211 B.n84 71.676
R1098 B.n207 B.n83 71.676
R1099 B.n203 B.n82 71.676
R1100 B.n199 B.n81 71.676
R1101 B.n195 B.n80 71.676
R1102 B.n191 B.n79 71.676
R1103 B.n187 B.n78 71.676
R1104 B.n183 B.n77 71.676
R1105 B.n179 B.n76 71.676
R1106 B.n175 B.n75 71.676
R1107 B.n171 B.n74 71.676
R1108 B.n167 B.n73 71.676
R1109 B.n163 B.n72 71.676
R1110 B.n159 B.n71 71.676
R1111 B.n155 B.n70 71.676
R1112 B.n151 B.n69 71.676
R1113 B.n147 B.n68 71.676
R1114 B.n143 B.n67 71.676
R1115 B.n139 B.n66 71.676
R1116 B.n135 B.n65 71.676
R1117 B.n131 B.n64 71.676
R1118 B.n127 B.n63 71.676
R1119 B.n123 B.n62 71.676
R1120 B.n119 B.n61 71.676
R1121 B.n115 B.n60 71.676
R1122 B.n111 B.n59 71.676
R1123 B.n107 B.n58 71.676
R1124 B.n103 B.n57 71.676
R1125 B.n99 B.n56 71.676
R1126 B.n95 B.n55 71.676
R1127 B.n311 B.n273 71.676
R1128 B.n315 B.n314 71.676
R1129 B.n320 B.n319 71.676
R1130 B.n323 B.n322 71.676
R1131 B.n328 B.n327 71.676
R1132 B.n331 B.n330 71.676
R1133 B.n336 B.n335 71.676
R1134 B.n339 B.n338 71.676
R1135 B.n344 B.n343 71.676
R1136 B.n347 B.n346 71.676
R1137 B.n352 B.n351 71.676
R1138 B.n355 B.n354 71.676
R1139 B.n360 B.n359 71.676
R1140 B.n363 B.n362 71.676
R1141 B.n369 B.n368 71.676
R1142 B.n372 B.n371 71.676
R1143 B.n377 B.n376 71.676
R1144 B.n380 B.n379 71.676
R1145 B.n388 B.n387 71.676
R1146 B.n391 B.n390 71.676
R1147 B.n396 B.n395 71.676
R1148 B.n399 B.n398 71.676
R1149 B.n404 B.n403 71.676
R1150 B.n407 B.n406 71.676
R1151 B.n412 B.n411 71.676
R1152 B.n415 B.n414 71.676
R1153 B.n420 B.n419 71.676
R1154 B.n423 B.n422 71.676
R1155 B.n428 B.n427 71.676
R1156 B.n431 B.n430 71.676
R1157 B.n436 B.n435 71.676
R1158 B.n439 B.n438 71.676
R1159 B.n312 B.n311 71.676
R1160 B.n314 B.n308 71.676
R1161 B.n321 B.n320 71.676
R1162 B.n322 B.n306 71.676
R1163 B.n329 B.n328 71.676
R1164 B.n330 B.n304 71.676
R1165 B.n337 B.n336 71.676
R1166 B.n338 B.n302 71.676
R1167 B.n345 B.n344 71.676
R1168 B.n346 B.n300 71.676
R1169 B.n353 B.n352 71.676
R1170 B.n354 B.n298 71.676
R1171 B.n361 B.n360 71.676
R1172 B.n362 B.n294 71.676
R1173 B.n370 B.n369 71.676
R1174 B.n371 B.n292 71.676
R1175 B.n378 B.n377 71.676
R1176 B.n379 B.n290 71.676
R1177 B.n389 B.n388 71.676
R1178 B.n390 B.n288 71.676
R1179 B.n397 B.n396 71.676
R1180 B.n398 B.n286 71.676
R1181 B.n405 B.n404 71.676
R1182 B.n406 B.n284 71.676
R1183 B.n413 B.n412 71.676
R1184 B.n414 B.n282 71.676
R1185 B.n421 B.n420 71.676
R1186 B.n422 B.n280 71.676
R1187 B.n429 B.n428 71.676
R1188 B.n430 B.n278 71.676
R1189 B.n437 B.n436 71.676
R1190 B.n440 B.n439 71.676
R1191 B.n631 B.n630 71.676
R1192 B.n631 B.n2 71.676
R1193 B.n93 B.n92 59.5399
R1194 B.n90 B.n89 59.5399
R1195 B.n385 B.n384 59.5399
R1196 B.n365 B.n296 59.5399
R1197 B.n445 B.n270 59.2011
R1198 B.n451 B.n270 59.2011
R1199 B.n451 B.n266 59.2011
R1200 B.n458 B.n266 59.2011
R1201 B.n458 B.n457 59.2011
R1202 B.n464 B.n259 59.2011
R1203 B.n470 B.n259 59.2011
R1204 B.n470 B.n255 59.2011
R1205 B.n476 B.n255 59.2011
R1206 B.n476 B.n251 59.2011
R1207 B.n482 B.n251 59.2011
R1208 B.n482 B.n247 59.2011
R1209 B.n488 B.n247 59.2011
R1210 B.n494 B.n243 59.2011
R1211 B.n494 B.n238 59.2011
R1212 B.n500 B.n238 59.2011
R1213 B.n500 B.n239 59.2011
R1214 B.n506 B.n231 59.2011
R1215 B.n512 B.n231 59.2011
R1216 B.n512 B.n227 59.2011
R1217 B.n519 B.n227 59.2011
R1218 B.n525 B.n223 59.2011
R1219 B.n525 B.n4 59.2011
R1220 B.n629 B.n4 59.2011
R1221 B.n629 B.n628 59.2011
R1222 B.n628 B.n627 59.2011
R1223 B.n627 B.n8 59.2011
R1224 B.n534 B.n8 59.2011
R1225 B.n620 B.n619 59.2011
R1226 B.n619 B.n618 59.2011
R1227 B.n618 B.n15 59.2011
R1228 B.n612 B.n15 59.2011
R1229 B.n611 B.n610 59.2011
R1230 B.n610 B.n22 59.2011
R1231 B.n604 B.n22 59.2011
R1232 B.n604 B.n603 59.2011
R1233 B.n602 B.n29 59.2011
R1234 B.n596 B.n29 59.2011
R1235 B.n596 B.n595 59.2011
R1236 B.n595 B.n594 59.2011
R1237 B.n594 B.n36 59.2011
R1238 B.n588 B.n36 59.2011
R1239 B.n588 B.n587 59.2011
R1240 B.n587 B.n586 59.2011
R1241 B.n580 B.n46 59.2011
R1242 B.n580 B.n579 59.2011
R1243 B.n579 B.n578 59.2011
R1244 B.n578 B.n50 59.2011
R1245 B.n572 B.n50 59.2011
R1246 B.n457 B.t7 52.2364
R1247 B.n46 B.t14 52.2364
R1248 B.t2 B.n243 48.754
R1249 B.n603 B.t4 48.754
R1250 B.n506 B.t3 43.5304
R1251 B.n612 B.t0 43.5304
R1252 B.t1 B.n223 38.3068
R1253 B.n534 B.t5 38.3068
R1254 B.n92 B.n91 33.552
R1255 B.n89 B.n88 33.552
R1256 B.n384 B.n383 33.552
R1257 B.n296 B.n295 33.552
R1258 B.n568 B.n567 29.5029
R1259 B.n447 B.n272 29.5029
R1260 B.n443 B.n442 29.5029
R1261 B.n574 B.n52 29.5029
R1262 B.n519 B.t1 20.8948
R1263 B.n620 B.t5 20.8948
R1264 B B.n632 18.0485
R1265 B.n239 B.t3 15.6713
R1266 B.t0 B.n611 15.6713
R1267 B.n448 B.n447 10.6151
R1268 B.n449 B.n448 10.6151
R1269 B.n449 B.n264 10.6151
R1270 B.n460 B.n264 10.6151
R1271 B.n461 B.n460 10.6151
R1272 B.n462 B.n461 10.6151
R1273 B.n462 B.n257 10.6151
R1274 B.n472 B.n257 10.6151
R1275 B.n473 B.n472 10.6151
R1276 B.n474 B.n473 10.6151
R1277 B.n474 B.n249 10.6151
R1278 B.n484 B.n249 10.6151
R1279 B.n485 B.n484 10.6151
R1280 B.n486 B.n485 10.6151
R1281 B.n486 B.n241 10.6151
R1282 B.n496 B.n241 10.6151
R1283 B.n497 B.n496 10.6151
R1284 B.n498 B.n497 10.6151
R1285 B.n498 B.n233 10.6151
R1286 B.n508 B.n233 10.6151
R1287 B.n509 B.n508 10.6151
R1288 B.n510 B.n509 10.6151
R1289 B.n510 B.n225 10.6151
R1290 B.n521 B.n225 10.6151
R1291 B.n522 B.n521 10.6151
R1292 B.n523 B.n522 10.6151
R1293 B.n523 B.n0 10.6151
R1294 B.n310 B.n272 10.6151
R1295 B.n310 B.n309 10.6151
R1296 B.n316 B.n309 10.6151
R1297 B.n317 B.n316 10.6151
R1298 B.n318 B.n317 10.6151
R1299 B.n318 B.n307 10.6151
R1300 B.n324 B.n307 10.6151
R1301 B.n325 B.n324 10.6151
R1302 B.n326 B.n325 10.6151
R1303 B.n326 B.n305 10.6151
R1304 B.n332 B.n305 10.6151
R1305 B.n333 B.n332 10.6151
R1306 B.n334 B.n333 10.6151
R1307 B.n334 B.n303 10.6151
R1308 B.n340 B.n303 10.6151
R1309 B.n341 B.n340 10.6151
R1310 B.n342 B.n341 10.6151
R1311 B.n342 B.n301 10.6151
R1312 B.n348 B.n301 10.6151
R1313 B.n349 B.n348 10.6151
R1314 B.n350 B.n349 10.6151
R1315 B.n350 B.n299 10.6151
R1316 B.n356 B.n299 10.6151
R1317 B.n357 B.n356 10.6151
R1318 B.n358 B.n357 10.6151
R1319 B.n358 B.n297 10.6151
R1320 B.n364 B.n297 10.6151
R1321 B.n367 B.n366 10.6151
R1322 B.n367 B.n293 10.6151
R1323 B.n373 B.n293 10.6151
R1324 B.n374 B.n373 10.6151
R1325 B.n375 B.n374 10.6151
R1326 B.n375 B.n291 10.6151
R1327 B.n381 B.n291 10.6151
R1328 B.n382 B.n381 10.6151
R1329 B.n386 B.n382 10.6151
R1330 B.n392 B.n289 10.6151
R1331 B.n393 B.n392 10.6151
R1332 B.n394 B.n393 10.6151
R1333 B.n394 B.n287 10.6151
R1334 B.n400 B.n287 10.6151
R1335 B.n401 B.n400 10.6151
R1336 B.n402 B.n401 10.6151
R1337 B.n402 B.n285 10.6151
R1338 B.n408 B.n285 10.6151
R1339 B.n409 B.n408 10.6151
R1340 B.n410 B.n409 10.6151
R1341 B.n410 B.n283 10.6151
R1342 B.n416 B.n283 10.6151
R1343 B.n417 B.n416 10.6151
R1344 B.n418 B.n417 10.6151
R1345 B.n418 B.n281 10.6151
R1346 B.n424 B.n281 10.6151
R1347 B.n425 B.n424 10.6151
R1348 B.n426 B.n425 10.6151
R1349 B.n426 B.n279 10.6151
R1350 B.n432 B.n279 10.6151
R1351 B.n433 B.n432 10.6151
R1352 B.n434 B.n433 10.6151
R1353 B.n434 B.n277 10.6151
R1354 B.n277 B.n276 10.6151
R1355 B.n441 B.n276 10.6151
R1356 B.n442 B.n441 10.6151
R1357 B.n443 B.n268 10.6151
R1358 B.n453 B.n268 10.6151
R1359 B.n454 B.n453 10.6151
R1360 B.n455 B.n454 10.6151
R1361 B.n455 B.n261 10.6151
R1362 B.n466 B.n261 10.6151
R1363 B.n467 B.n466 10.6151
R1364 B.n468 B.n467 10.6151
R1365 B.n468 B.n253 10.6151
R1366 B.n478 B.n253 10.6151
R1367 B.n479 B.n478 10.6151
R1368 B.n480 B.n479 10.6151
R1369 B.n480 B.n245 10.6151
R1370 B.n490 B.n245 10.6151
R1371 B.n491 B.n490 10.6151
R1372 B.n492 B.n491 10.6151
R1373 B.n492 B.n236 10.6151
R1374 B.n502 B.n236 10.6151
R1375 B.n503 B.n502 10.6151
R1376 B.n504 B.n503 10.6151
R1377 B.n504 B.n229 10.6151
R1378 B.n514 B.n229 10.6151
R1379 B.n515 B.n514 10.6151
R1380 B.n517 B.n515 10.6151
R1381 B.n517 B.n516 10.6151
R1382 B.n516 B.n221 10.6151
R1383 B.n528 B.n221 10.6151
R1384 B.n529 B.n528 10.6151
R1385 B.n530 B.n529 10.6151
R1386 B.n531 B.n530 10.6151
R1387 B.n532 B.n531 10.6151
R1388 B.n536 B.n532 10.6151
R1389 B.n537 B.n536 10.6151
R1390 B.n538 B.n537 10.6151
R1391 B.n539 B.n538 10.6151
R1392 B.n541 B.n539 10.6151
R1393 B.n542 B.n541 10.6151
R1394 B.n543 B.n542 10.6151
R1395 B.n544 B.n543 10.6151
R1396 B.n546 B.n544 10.6151
R1397 B.n547 B.n546 10.6151
R1398 B.n548 B.n547 10.6151
R1399 B.n549 B.n548 10.6151
R1400 B.n551 B.n549 10.6151
R1401 B.n552 B.n551 10.6151
R1402 B.n553 B.n552 10.6151
R1403 B.n554 B.n553 10.6151
R1404 B.n556 B.n554 10.6151
R1405 B.n557 B.n556 10.6151
R1406 B.n558 B.n557 10.6151
R1407 B.n559 B.n558 10.6151
R1408 B.n561 B.n559 10.6151
R1409 B.n562 B.n561 10.6151
R1410 B.n563 B.n562 10.6151
R1411 B.n564 B.n563 10.6151
R1412 B.n566 B.n564 10.6151
R1413 B.n567 B.n566 10.6151
R1414 B.n624 B.n1 10.6151
R1415 B.n624 B.n623 10.6151
R1416 B.n623 B.n622 10.6151
R1417 B.n622 B.n10 10.6151
R1418 B.n616 B.n10 10.6151
R1419 B.n616 B.n615 10.6151
R1420 B.n615 B.n614 10.6151
R1421 B.n614 B.n17 10.6151
R1422 B.n608 B.n17 10.6151
R1423 B.n608 B.n607 10.6151
R1424 B.n607 B.n606 10.6151
R1425 B.n606 B.n24 10.6151
R1426 B.n600 B.n24 10.6151
R1427 B.n600 B.n599 10.6151
R1428 B.n599 B.n598 10.6151
R1429 B.n598 B.n31 10.6151
R1430 B.n592 B.n31 10.6151
R1431 B.n592 B.n591 10.6151
R1432 B.n591 B.n590 10.6151
R1433 B.n590 B.n38 10.6151
R1434 B.n584 B.n38 10.6151
R1435 B.n584 B.n583 10.6151
R1436 B.n583 B.n582 10.6151
R1437 B.n582 B.n44 10.6151
R1438 B.n576 B.n44 10.6151
R1439 B.n576 B.n575 10.6151
R1440 B.n575 B.n574 10.6151
R1441 B.n94 B.n52 10.6151
R1442 B.n97 B.n94 10.6151
R1443 B.n98 B.n97 10.6151
R1444 B.n101 B.n98 10.6151
R1445 B.n102 B.n101 10.6151
R1446 B.n105 B.n102 10.6151
R1447 B.n106 B.n105 10.6151
R1448 B.n109 B.n106 10.6151
R1449 B.n110 B.n109 10.6151
R1450 B.n113 B.n110 10.6151
R1451 B.n114 B.n113 10.6151
R1452 B.n117 B.n114 10.6151
R1453 B.n118 B.n117 10.6151
R1454 B.n121 B.n118 10.6151
R1455 B.n122 B.n121 10.6151
R1456 B.n125 B.n122 10.6151
R1457 B.n126 B.n125 10.6151
R1458 B.n129 B.n126 10.6151
R1459 B.n130 B.n129 10.6151
R1460 B.n133 B.n130 10.6151
R1461 B.n134 B.n133 10.6151
R1462 B.n137 B.n134 10.6151
R1463 B.n138 B.n137 10.6151
R1464 B.n141 B.n138 10.6151
R1465 B.n142 B.n141 10.6151
R1466 B.n145 B.n142 10.6151
R1467 B.n146 B.n145 10.6151
R1468 B.n150 B.n149 10.6151
R1469 B.n153 B.n150 10.6151
R1470 B.n154 B.n153 10.6151
R1471 B.n157 B.n154 10.6151
R1472 B.n158 B.n157 10.6151
R1473 B.n161 B.n158 10.6151
R1474 B.n162 B.n161 10.6151
R1475 B.n165 B.n162 10.6151
R1476 B.n166 B.n165 10.6151
R1477 B.n170 B.n169 10.6151
R1478 B.n173 B.n170 10.6151
R1479 B.n174 B.n173 10.6151
R1480 B.n177 B.n174 10.6151
R1481 B.n178 B.n177 10.6151
R1482 B.n181 B.n178 10.6151
R1483 B.n182 B.n181 10.6151
R1484 B.n185 B.n182 10.6151
R1485 B.n186 B.n185 10.6151
R1486 B.n189 B.n186 10.6151
R1487 B.n190 B.n189 10.6151
R1488 B.n193 B.n190 10.6151
R1489 B.n194 B.n193 10.6151
R1490 B.n197 B.n194 10.6151
R1491 B.n198 B.n197 10.6151
R1492 B.n201 B.n198 10.6151
R1493 B.n202 B.n201 10.6151
R1494 B.n205 B.n202 10.6151
R1495 B.n206 B.n205 10.6151
R1496 B.n209 B.n206 10.6151
R1497 B.n210 B.n209 10.6151
R1498 B.n213 B.n210 10.6151
R1499 B.n214 B.n213 10.6151
R1500 B.n217 B.n214 10.6151
R1501 B.n219 B.n217 10.6151
R1502 B.n220 B.n219 10.6151
R1503 B.n568 B.n220 10.6151
R1504 B.n488 B.t2 10.4477
R1505 B.t4 B.n602 10.4477
R1506 B.n365 B.n364 9.36635
R1507 B.n385 B.n289 9.36635
R1508 B.n146 B.n93 9.36635
R1509 B.n169 B.n90 9.36635
R1510 B.n632 B.n0 8.11757
R1511 B.n632 B.n1 8.11757
R1512 B.n464 B.t7 6.96528
R1513 B.n586 B.t14 6.96528
R1514 B.n366 B.n365 1.24928
R1515 B.n386 B.n385 1.24928
R1516 B.n149 B.n93 1.24928
R1517 B.n166 B.n90 1.24928
R1518 VN.n9 VN.n8 174.581
R1519 VN.n19 VN.n18 174.581
R1520 VN.n3 VN.t4 161.577
R1521 VN.n13 VN.t1 161.577
R1522 VN.n17 VN.n10 161.3
R1523 VN.n16 VN.n15 161.3
R1524 VN.n14 VN.n11 161.3
R1525 VN.n7 VN.n0 161.3
R1526 VN.n6 VN.n5 161.3
R1527 VN.n4 VN.n1 161.3
R1528 VN.n2 VN.t2 126.698
R1529 VN.n8 VN.t3 126.698
R1530 VN.n12 VN.t5 126.698
R1531 VN.n18 VN.t0 126.698
R1532 VN.n6 VN.n1 53.6554
R1533 VN.n16 VN.n11 53.6554
R1534 VN.n3 VN.n2 41.8949
R1535 VN.n13 VN.n12 41.8949
R1536 VN VN.n19 40.7562
R1537 VN.n7 VN.n6 27.4986
R1538 VN.n17 VN.n16 27.4986
R1539 VN.n2 VN.n1 24.5923
R1540 VN.n12 VN.n11 24.5923
R1541 VN.n14 VN.n13 17.6108
R1542 VN.n4 VN.n3 17.6108
R1543 VN.n8 VN.n7 11.3127
R1544 VN.n18 VN.n17 11.3127
R1545 VN.n19 VN.n10 0.189894
R1546 VN.n15 VN.n10 0.189894
R1547 VN.n15 VN.n14 0.189894
R1548 VN.n5 VN.n4 0.189894
R1549 VN.n5 VN.n0 0.189894
R1550 VN.n9 VN.n0 0.189894
R1551 VN VN.n9 0.0516364
R1552 VDD2.n75 VDD2.n41 289.615
R1553 VDD2.n34 VDD2.n0 289.615
R1554 VDD2.n76 VDD2.n75 185
R1555 VDD2.n74 VDD2.n73 185
R1556 VDD2.n45 VDD2.n44 185
R1557 VDD2.n68 VDD2.n67 185
R1558 VDD2.n66 VDD2.n65 185
R1559 VDD2.n49 VDD2.n48 185
R1560 VDD2.n60 VDD2.n59 185
R1561 VDD2.n58 VDD2.n57 185
R1562 VDD2.n53 VDD2.n52 185
R1563 VDD2.n12 VDD2.n11 185
R1564 VDD2.n17 VDD2.n16 185
R1565 VDD2.n19 VDD2.n18 185
R1566 VDD2.n8 VDD2.n7 185
R1567 VDD2.n25 VDD2.n24 185
R1568 VDD2.n27 VDD2.n26 185
R1569 VDD2.n4 VDD2.n3 185
R1570 VDD2.n33 VDD2.n32 185
R1571 VDD2.n35 VDD2.n34 185
R1572 VDD2.n54 VDD2.t5 147.659
R1573 VDD2.n13 VDD2.t1 147.659
R1574 VDD2.n75 VDD2.n74 104.615
R1575 VDD2.n74 VDD2.n44 104.615
R1576 VDD2.n67 VDD2.n44 104.615
R1577 VDD2.n67 VDD2.n66 104.615
R1578 VDD2.n66 VDD2.n48 104.615
R1579 VDD2.n59 VDD2.n48 104.615
R1580 VDD2.n59 VDD2.n58 104.615
R1581 VDD2.n58 VDD2.n52 104.615
R1582 VDD2.n17 VDD2.n11 104.615
R1583 VDD2.n18 VDD2.n17 104.615
R1584 VDD2.n18 VDD2.n7 104.615
R1585 VDD2.n25 VDD2.n7 104.615
R1586 VDD2.n26 VDD2.n25 104.615
R1587 VDD2.n26 VDD2.n3 104.615
R1588 VDD2.n33 VDD2.n3 104.615
R1589 VDD2.n34 VDD2.n33 104.615
R1590 VDD2.n40 VDD2.n39 63.9663
R1591 VDD2 VDD2.n81 63.9635
R1592 VDD2.t5 VDD2.n52 52.3082
R1593 VDD2.t1 VDD2.n11 52.3082
R1594 VDD2.n40 VDD2.n38 48.3758
R1595 VDD2.n80 VDD2.n79 47.3126
R1596 VDD2.n80 VDD2.n40 34.9071
R1597 VDD2.n54 VDD2.n53 15.6677
R1598 VDD2.n13 VDD2.n12 15.6677
R1599 VDD2.n57 VDD2.n56 12.8005
R1600 VDD2.n16 VDD2.n15 12.8005
R1601 VDD2.n60 VDD2.n51 12.0247
R1602 VDD2.n19 VDD2.n10 12.0247
R1603 VDD2.n61 VDD2.n49 11.249
R1604 VDD2.n20 VDD2.n8 11.249
R1605 VDD2.n65 VDD2.n64 10.4732
R1606 VDD2.n24 VDD2.n23 10.4732
R1607 VDD2.n68 VDD2.n47 9.69747
R1608 VDD2.n27 VDD2.n6 9.69747
R1609 VDD2.n79 VDD2.n78 9.45567
R1610 VDD2.n38 VDD2.n37 9.45567
R1611 VDD2.n78 VDD2.n77 9.3005
R1612 VDD2.n43 VDD2.n42 9.3005
R1613 VDD2.n72 VDD2.n71 9.3005
R1614 VDD2.n70 VDD2.n69 9.3005
R1615 VDD2.n47 VDD2.n46 9.3005
R1616 VDD2.n64 VDD2.n63 9.3005
R1617 VDD2.n62 VDD2.n61 9.3005
R1618 VDD2.n51 VDD2.n50 9.3005
R1619 VDD2.n56 VDD2.n55 9.3005
R1620 VDD2.n37 VDD2.n36 9.3005
R1621 VDD2.n31 VDD2.n30 9.3005
R1622 VDD2.n29 VDD2.n28 9.3005
R1623 VDD2.n6 VDD2.n5 9.3005
R1624 VDD2.n23 VDD2.n22 9.3005
R1625 VDD2.n21 VDD2.n20 9.3005
R1626 VDD2.n10 VDD2.n9 9.3005
R1627 VDD2.n15 VDD2.n14 9.3005
R1628 VDD2.n2 VDD2.n1 9.3005
R1629 VDD2.n69 VDD2.n45 8.92171
R1630 VDD2.n28 VDD2.n4 8.92171
R1631 VDD2.n73 VDD2.n72 8.14595
R1632 VDD2.n32 VDD2.n31 8.14595
R1633 VDD2.n79 VDD2.n41 7.3702
R1634 VDD2.n76 VDD2.n43 7.3702
R1635 VDD2.n35 VDD2.n2 7.3702
R1636 VDD2.n38 VDD2.n0 7.3702
R1637 VDD2.n77 VDD2.n41 6.59444
R1638 VDD2.n77 VDD2.n76 6.59444
R1639 VDD2.n36 VDD2.n35 6.59444
R1640 VDD2.n36 VDD2.n0 6.59444
R1641 VDD2.n73 VDD2.n43 5.81868
R1642 VDD2.n32 VDD2.n2 5.81868
R1643 VDD2.n72 VDD2.n45 5.04292
R1644 VDD2.n31 VDD2.n4 5.04292
R1645 VDD2.n55 VDD2.n54 4.38565
R1646 VDD2.n14 VDD2.n13 4.38565
R1647 VDD2.n69 VDD2.n68 4.26717
R1648 VDD2.n28 VDD2.n27 4.26717
R1649 VDD2.n65 VDD2.n47 3.49141
R1650 VDD2.n24 VDD2.n6 3.49141
R1651 VDD2.n64 VDD2.n49 2.71565
R1652 VDD2.n23 VDD2.n8 2.71565
R1653 VDD2.n81 VDD2.t0 2.69072
R1654 VDD2.n81 VDD2.t4 2.69072
R1655 VDD2.n39 VDD2.t3 2.69072
R1656 VDD2.n39 VDD2.t2 2.69072
R1657 VDD2.n61 VDD2.n60 1.93989
R1658 VDD2.n20 VDD2.n19 1.93989
R1659 VDD2 VDD2.n80 1.17722
R1660 VDD2.n57 VDD2.n51 1.16414
R1661 VDD2.n16 VDD2.n10 1.16414
R1662 VDD2.n56 VDD2.n53 0.388379
R1663 VDD2.n15 VDD2.n12 0.388379
R1664 VDD2.n78 VDD2.n42 0.155672
R1665 VDD2.n71 VDD2.n42 0.155672
R1666 VDD2.n71 VDD2.n70 0.155672
R1667 VDD2.n70 VDD2.n46 0.155672
R1668 VDD2.n63 VDD2.n46 0.155672
R1669 VDD2.n63 VDD2.n62 0.155672
R1670 VDD2.n62 VDD2.n50 0.155672
R1671 VDD2.n55 VDD2.n50 0.155672
R1672 VDD2.n14 VDD2.n9 0.155672
R1673 VDD2.n21 VDD2.n9 0.155672
R1674 VDD2.n22 VDD2.n21 0.155672
R1675 VDD2.n22 VDD2.n5 0.155672
R1676 VDD2.n29 VDD2.n5 0.155672
R1677 VDD2.n30 VDD2.n29 0.155672
R1678 VDD2.n30 VDD2.n1 0.155672
R1679 VDD2.n37 VDD2.n1 0.155672
C0 VN VP 4.89822f
C1 VTAIL VP 3.74582f
C2 VTAIL VN 3.73151f
C3 VDD1 VP 3.86859f
C4 VDD2 VP 0.356522f
C5 VDD1 VN 0.149435f
C6 VDD2 VN 3.66407f
C7 VDD1 VTAIL 5.90021f
C8 VDD2 VTAIL 5.94289f
C9 VDD2 VDD1 0.968635f
C10 VDD2 B 4.211111f
C11 VDD1 B 4.27143f
C12 VTAIL B 5.185142f
C13 VN B 9.04932f
C14 VP B 7.55766f
C15 VDD2.n0 B 0.030923f
C16 VDD2.n1 B 0.022f
C17 VDD2.n2 B 0.011822f
C18 VDD2.n3 B 0.027942f
C19 VDD2.n4 B 0.012517f
C20 VDD2.n5 B 0.022f
C21 VDD2.n6 B 0.011822f
C22 VDD2.n7 B 0.027942f
C23 VDD2.n8 B 0.012517f
C24 VDD2.n9 B 0.022f
C25 VDD2.n10 B 0.011822f
C26 VDD2.n11 B 0.020957f
C27 VDD2.n12 B 0.016506f
C28 VDD2.t1 B 0.045533f
C29 VDD2.n13 B 0.101421f
C30 VDD2.n14 B 0.66092f
C31 VDD2.n15 B 0.011822f
C32 VDD2.n16 B 0.012517f
C33 VDD2.n17 B 0.027942f
C34 VDD2.n18 B 0.027942f
C35 VDD2.n19 B 0.012517f
C36 VDD2.n20 B 0.011822f
C37 VDD2.n21 B 0.022f
C38 VDD2.n22 B 0.022f
C39 VDD2.n23 B 0.011822f
C40 VDD2.n24 B 0.012517f
C41 VDD2.n25 B 0.027942f
C42 VDD2.n26 B 0.027942f
C43 VDD2.n27 B 0.012517f
C44 VDD2.n28 B 0.011822f
C45 VDD2.n29 B 0.022f
C46 VDD2.n30 B 0.022f
C47 VDD2.n31 B 0.011822f
C48 VDD2.n32 B 0.012517f
C49 VDD2.n33 B 0.027942f
C50 VDD2.n34 B 0.06049f
C51 VDD2.n35 B 0.012517f
C52 VDD2.n36 B 0.011822f
C53 VDD2.n37 B 0.048447f
C54 VDD2.n38 B 0.051549f
C55 VDD2.t3 B 0.127953f
C56 VDD2.t2 B 0.127953f
C57 VDD2.n39 B 1.09229f
C58 VDD2.n40 B 1.65334f
C59 VDD2.n41 B 0.030923f
C60 VDD2.n42 B 0.022f
C61 VDD2.n43 B 0.011822f
C62 VDD2.n44 B 0.027942f
C63 VDD2.n45 B 0.012517f
C64 VDD2.n46 B 0.022f
C65 VDD2.n47 B 0.011822f
C66 VDD2.n48 B 0.027942f
C67 VDD2.n49 B 0.012517f
C68 VDD2.n50 B 0.022f
C69 VDD2.n51 B 0.011822f
C70 VDD2.n52 B 0.020957f
C71 VDD2.n53 B 0.016506f
C72 VDD2.t5 B 0.045533f
C73 VDD2.n54 B 0.101421f
C74 VDD2.n55 B 0.66092f
C75 VDD2.n56 B 0.011822f
C76 VDD2.n57 B 0.012517f
C77 VDD2.n58 B 0.027942f
C78 VDD2.n59 B 0.027942f
C79 VDD2.n60 B 0.012517f
C80 VDD2.n61 B 0.011822f
C81 VDD2.n62 B 0.022f
C82 VDD2.n63 B 0.022f
C83 VDD2.n64 B 0.011822f
C84 VDD2.n65 B 0.012517f
C85 VDD2.n66 B 0.027942f
C86 VDD2.n67 B 0.027942f
C87 VDD2.n68 B 0.012517f
C88 VDD2.n69 B 0.011822f
C89 VDD2.n70 B 0.022f
C90 VDD2.n71 B 0.022f
C91 VDD2.n72 B 0.011822f
C92 VDD2.n73 B 0.012517f
C93 VDD2.n74 B 0.027942f
C94 VDD2.n75 B 0.06049f
C95 VDD2.n76 B 0.012517f
C96 VDD2.n77 B 0.011822f
C97 VDD2.n78 B 0.048447f
C98 VDD2.n79 B 0.048982f
C99 VDD2.n80 B 1.64331f
C100 VDD2.t0 B 0.127953f
C101 VDD2.t4 B 0.127953f
C102 VDD2.n81 B 1.09227f
C103 VN.n0 B 0.034948f
C104 VN.t3 B 0.963487f
C105 VN.n1 B 0.061343f
C106 VN.t4 B 1.07065f
C107 VN.t2 B 0.963487f
C108 VN.n2 B 0.447299f
C109 VN.n3 B 0.435606f
C110 VN.n4 B 0.219246f
C111 VN.n5 B 0.034948f
C112 VN.n6 B 0.037288f
C113 VN.n7 B 0.050507f
C114 VN.n8 B 0.435957f
C115 VN.n9 B 0.032646f
C116 VN.n10 B 0.034948f
C117 VN.t0 B 0.963487f
C118 VN.n11 B 0.061343f
C119 VN.t1 B 1.07065f
C120 VN.t5 B 0.963487f
C121 VN.n12 B 0.447299f
C122 VN.n13 B 0.435606f
C123 VN.n14 B 0.219246f
C124 VN.n15 B 0.034948f
C125 VN.n16 B 0.037288f
C126 VN.n17 B 0.050507f
C127 VN.n18 B 0.435957f
C128 VN.n19 B 1.37807f
C129 VDD1.n0 B 0.031302f
C130 VDD1.n1 B 0.02227f
C131 VDD1.n2 B 0.011967f
C132 VDD1.n3 B 0.028285f
C133 VDD1.n4 B 0.012671f
C134 VDD1.n5 B 0.02227f
C135 VDD1.n6 B 0.011967f
C136 VDD1.n7 B 0.028285f
C137 VDD1.n8 B 0.012671f
C138 VDD1.n9 B 0.02227f
C139 VDD1.n10 B 0.011967f
C140 VDD1.n11 B 0.021214f
C141 VDD1.n12 B 0.016709f
C142 VDD1.t5 B 0.046092f
C143 VDD1.n13 B 0.102665f
C144 VDD1.n14 B 0.669026f
C145 VDD1.n15 B 0.011967f
C146 VDD1.n16 B 0.012671f
C147 VDD1.n17 B 0.028285f
C148 VDD1.n18 B 0.028285f
C149 VDD1.n19 B 0.012671f
C150 VDD1.n20 B 0.011967f
C151 VDD1.n21 B 0.02227f
C152 VDD1.n22 B 0.02227f
C153 VDD1.n23 B 0.011967f
C154 VDD1.n24 B 0.012671f
C155 VDD1.n25 B 0.028285f
C156 VDD1.n26 B 0.028285f
C157 VDD1.n27 B 0.012671f
C158 VDD1.n28 B 0.011967f
C159 VDD1.n29 B 0.02227f
C160 VDD1.n30 B 0.02227f
C161 VDD1.n31 B 0.011967f
C162 VDD1.n32 B 0.012671f
C163 VDD1.n33 B 0.028285f
C164 VDD1.n34 B 0.061232f
C165 VDD1.n35 B 0.012671f
C166 VDD1.n36 B 0.011967f
C167 VDD1.n37 B 0.049041f
C168 VDD1.n38 B 0.052638f
C169 VDD1.n39 B 0.031302f
C170 VDD1.n40 B 0.02227f
C171 VDD1.n41 B 0.011967f
C172 VDD1.n42 B 0.028285f
C173 VDD1.n43 B 0.012671f
C174 VDD1.n44 B 0.02227f
C175 VDD1.n45 B 0.011967f
C176 VDD1.n46 B 0.028285f
C177 VDD1.n47 B 0.012671f
C178 VDD1.n48 B 0.02227f
C179 VDD1.n49 B 0.011967f
C180 VDD1.n50 B 0.021214f
C181 VDD1.n51 B 0.016709f
C182 VDD1.t2 B 0.046092f
C183 VDD1.n52 B 0.102665f
C184 VDD1.n53 B 0.669026f
C185 VDD1.n54 B 0.011967f
C186 VDD1.n55 B 0.012671f
C187 VDD1.n56 B 0.028285f
C188 VDD1.n57 B 0.028285f
C189 VDD1.n58 B 0.012671f
C190 VDD1.n59 B 0.011967f
C191 VDD1.n60 B 0.02227f
C192 VDD1.n61 B 0.02227f
C193 VDD1.n62 B 0.011967f
C194 VDD1.n63 B 0.012671f
C195 VDD1.n64 B 0.028285f
C196 VDD1.n65 B 0.028285f
C197 VDD1.n66 B 0.012671f
C198 VDD1.n67 B 0.011967f
C199 VDD1.n68 B 0.02227f
C200 VDD1.n69 B 0.02227f
C201 VDD1.n70 B 0.011967f
C202 VDD1.n71 B 0.012671f
C203 VDD1.n72 B 0.028285f
C204 VDD1.n73 B 0.061232f
C205 VDD1.n74 B 0.012671f
C206 VDD1.n75 B 0.011967f
C207 VDD1.n76 B 0.049041f
C208 VDD1.n77 B 0.052182f
C209 VDD1.t4 B 0.129522f
C210 VDD1.t3 B 0.129522f
C211 VDD1.n78 B 1.10569f
C212 VDD1.n79 B 1.75462f
C213 VDD1.t1 B 0.129522f
C214 VDD1.t0 B 0.129522f
C215 VDD1.n80 B 1.10407f
C216 VDD1.n81 B 1.86237f
C217 VTAIL.t5 B 0.142937f
C218 VTAIL.t0 B 0.142937f
C219 VTAIL.n0 B 1.14758f
C220 VTAIL.n1 B 0.372009f
C221 VTAIL.n2 B 0.034544f
C222 VTAIL.n3 B 0.024576f
C223 VTAIL.n4 B 0.013206f
C224 VTAIL.n5 B 0.031215f
C225 VTAIL.n6 B 0.013983f
C226 VTAIL.n7 B 0.024576f
C227 VTAIL.n8 B 0.013206f
C228 VTAIL.n9 B 0.031215f
C229 VTAIL.n10 B 0.013983f
C230 VTAIL.n11 B 0.024576f
C231 VTAIL.n12 B 0.013206f
C232 VTAIL.n13 B 0.023411f
C233 VTAIL.n14 B 0.018439f
C234 VTAIL.t11 B 0.050865f
C235 VTAIL.n15 B 0.113299f
C236 VTAIL.n16 B 0.73832f
C237 VTAIL.n17 B 0.013206f
C238 VTAIL.n18 B 0.013983f
C239 VTAIL.n19 B 0.031215f
C240 VTAIL.n20 B 0.031215f
C241 VTAIL.n21 B 0.013983f
C242 VTAIL.n22 B 0.013206f
C243 VTAIL.n23 B 0.024576f
C244 VTAIL.n24 B 0.024576f
C245 VTAIL.n25 B 0.013206f
C246 VTAIL.n26 B 0.013983f
C247 VTAIL.n27 B 0.031215f
C248 VTAIL.n28 B 0.031215f
C249 VTAIL.n29 B 0.013983f
C250 VTAIL.n30 B 0.013206f
C251 VTAIL.n31 B 0.024576f
C252 VTAIL.n32 B 0.024576f
C253 VTAIL.n33 B 0.013206f
C254 VTAIL.n34 B 0.013983f
C255 VTAIL.n35 B 0.031215f
C256 VTAIL.n36 B 0.067574f
C257 VTAIL.n37 B 0.013983f
C258 VTAIL.n38 B 0.013206f
C259 VTAIL.n39 B 0.054121f
C260 VTAIL.n40 B 0.037726f
C261 VTAIL.n41 B 0.233834f
C262 VTAIL.t6 B 0.142937f
C263 VTAIL.t8 B 0.142937f
C264 VTAIL.n42 B 1.14758f
C265 VTAIL.n43 B 1.43221f
C266 VTAIL.t2 B 0.142937f
C267 VTAIL.t3 B 0.142937f
C268 VTAIL.n44 B 1.14759f
C269 VTAIL.n45 B 1.4322f
C270 VTAIL.n46 B 0.034544f
C271 VTAIL.n47 B 0.024576f
C272 VTAIL.n48 B 0.013206f
C273 VTAIL.n49 B 0.031215f
C274 VTAIL.n50 B 0.013983f
C275 VTAIL.n51 B 0.024576f
C276 VTAIL.n52 B 0.013206f
C277 VTAIL.n53 B 0.031215f
C278 VTAIL.n54 B 0.013983f
C279 VTAIL.n55 B 0.024576f
C280 VTAIL.n56 B 0.013206f
C281 VTAIL.n57 B 0.023411f
C282 VTAIL.n58 B 0.018439f
C283 VTAIL.t1 B 0.050865f
C284 VTAIL.n59 B 0.113299f
C285 VTAIL.n60 B 0.73832f
C286 VTAIL.n61 B 0.013206f
C287 VTAIL.n62 B 0.013983f
C288 VTAIL.n63 B 0.031215f
C289 VTAIL.n64 B 0.031215f
C290 VTAIL.n65 B 0.013983f
C291 VTAIL.n66 B 0.013206f
C292 VTAIL.n67 B 0.024576f
C293 VTAIL.n68 B 0.024576f
C294 VTAIL.n69 B 0.013206f
C295 VTAIL.n70 B 0.013983f
C296 VTAIL.n71 B 0.031215f
C297 VTAIL.n72 B 0.031215f
C298 VTAIL.n73 B 0.013983f
C299 VTAIL.n74 B 0.013206f
C300 VTAIL.n75 B 0.024576f
C301 VTAIL.n76 B 0.024576f
C302 VTAIL.n77 B 0.013206f
C303 VTAIL.n78 B 0.013983f
C304 VTAIL.n79 B 0.031215f
C305 VTAIL.n80 B 0.067574f
C306 VTAIL.n81 B 0.013983f
C307 VTAIL.n82 B 0.013206f
C308 VTAIL.n83 B 0.054121f
C309 VTAIL.n84 B 0.037726f
C310 VTAIL.n85 B 0.233834f
C311 VTAIL.t10 B 0.142937f
C312 VTAIL.t9 B 0.142937f
C313 VTAIL.n86 B 1.14759f
C314 VTAIL.n87 B 0.455969f
C315 VTAIL.n88 B 0.034544f
C316 VTAIL.n89 B 0.024576f
C317 VTAIL.n90 B 0.013206f
C318 VTAIL.n91 B 0.031215f
C319 VTAIL.n92 B 0.013983f
C320 VTAIL.n93 B 0.024576f
C321 VTAIL.n94 B 0.013206f
C322 VTAIL.n95 B 0.031215f
C323 VTAIL.n96 B 0.013983f
C324 VTAIL.n97 B 0.024576f
C325 VTAIL.n98 B 0.013206f
C326 VTAIL.n99 B 0.023411f
C327 VTAIL.n100 B 0.018439f
C328 VTAIL.t7 B 0.050865f
C329 VTAIL.n101 B 0.113299f
C330 VTAIL.n102 B 0.73832f
C331 VTAIL.n103 B 0.013206f
C332 VTAIL.n104 B 0.013983f
C333 VTAIL.n105 B 0.031215f
C334 VTAIL.n106 B 0.031215f
C335 VTAIL.n107 B 0.013983f
C336 VTAIL.n108 B 0.013206f
C337 VTAIL.n109 B 0.024576f
C338 VTAIL.n110 B 0.024576f
C339 VTAIL.n111 B 0.013206f
C340 VTAIL.n112 B 0.013983f
C341 VTAIL.n113 B 0.031215f
C342 VTAIL.n114 B 0.031215f
C343 VTAIL.n115 B 0.013983f
C344 VTAIL.n116 B 0.013206f
C345 VTAIL.n117 B 0.024576f
C346 VTAIL.n118 B 0.024576f
C347 VTAIL.n119 B 0.013206f
C348 VTAIL.n120 B 0.013983f
C349 VTAIL.n121 B 0.031215f
C350 VTAIL.n122 B 0.067574f
C351 VTAIL.n123 B 0.013983f
C352 VTAIL.n124 B 0.013206f
C353 VTAIL.n125 B 0.054121f
C354 VTAIL.n126 B 0.037726f
C355 VTAIL.n127 B 1.09196f
C356 VTAIL.n128 B 0.034544f
C357 VTAIL.n129 B 0.024576f
C358 VTAIL.n130 B 0.013206f
C359 VTAIL.n131 B 0.031215f
C360 VTAIL.n132 B 0.013983f
C361 VTAIL.n133 B 0.024576f
C362 VTAIL.n134 B 0.013206f
C363 VTAIL.n135 B 0.031215f
C364 VTAIL.n136 B 0.013983f
C365 VTAIL.n137 B 0.024576f
C366 VTAIL.n138 B 0.013206f
C367 VTAIL.n139 B 0.023411f
C368 VTAIL.n140 B 0.018439f
C369 VTAIL.t4 B 0.050865f
C370 VTAIL.n141 B 0.113299f
C371 VTAIL.n142 B 0.73832f
C372 VTAIL.n143 B 0.013206f
C373 VTAIL.n144 B 0.013983f
C374 VTAIL.n145 B 0.031215f
C375 VTAIL.n146 B 0.031215f
C376 VTAIL.n147 B 0.013983f
C377 VTAIL.n148 B 0.013206f
C378 VTAIL.n149 B 0.024576f
C379 VTAIL.n150 B 0.024576f
C380 VTAIL.n151 B 0.013206f
C381 VTAIL.n152 B 0.013983f
C382 VTAIL.n153 B 0.031215f
C383 VTAIL.n154 B 0.031215f
C384 VTAIL.n155 B 0.013983f
C385 VTAIL.n156 B 0.013206f
C386 VTAIL.n157 B 0.024576f
C387 VTAIL.n158 B 0.024576f
C388 VTAIL.n159 B 0.013206f
C389 VTAIL.n160 B 0.013983f
C390 VTAIL.n161 B 0.031215f
C391 VTAIL.n162 B 0.067574f
C392 VTAIL.n163 B 0.013983f
C393 VTAIL.n164 B 0.013206f
C394 VTAIL.n165 B 0.054121f
C395 VTAIL.n166 B 0.037726f
C396 VTAIL.n167 B 1.05783f
C397 VP.n0 B 0.035659f
C398 VP.t2 B 0.98308f
C399 VP.n1 B 0.06259f
C400 VP.n2 B 0.035659f
C401 VP.t1 B 0.98308f
C402 VP.n3 B 0.051534f
C403 VP.n4 B 0.035659f
C404 VP.t5 B 0.98308f
C405 VP.n5 B 0.06259f
C406 VP.t0 B 1.09242f
C407 VP.t4 B 0.98308f
C408 VP.n6 B 0.456395f
C409 VP.n7 B 0.444464f
C410 VP.n8 B 0.223705f
C411 VP.n9 B 0.035659f
C412 VP.n10 B 0.038046f
C413 VP.n11 B 0.051534f
C414 VP.n12 B 0.444822f
C415 VP.n13 B 1.38263f
C416 VP.t3 B 0.98308f
C417 VP.n14 B 0.444822f
C418 VP.n15 B 1.41447f
C419 VP.n16 B 0.035659f
C420 VP.n17 B 0.035659f
C421 VP.n18 B 0.038046f
C422 VP.n19 B 0.06259f
C423 VP.n20 B 0.409365f
C424 VP.n21 B 0.035659f
C425 VP.n22 B 0.035659f
C426 VP.n23 B 0.035659f
C427 VP.n24 B 0.038046f
C428 VP.n25 B 0.051534f
C429 VP.n26 B 0.444822f
C430 VP.n27 B 0.03331f
.ends

