* NGSPICE file created from diff_pair_sample_1145.ext - technology: sky130A

.subckt diff_pair_sample_1145 VTAIL VN VP B VDD2 VDD1
X0 VTAIL.t15 VP.t0 VDD1.t7 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=1.67805 ps=10.5 w=10.17 l=0.98
X1 B.t11 B.t9 B.t10 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=0 ps=0 w=10.17 l=0.98
X2 VDD1.t4 VP.t1 VTAIL.t14 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=3.9663 ps=21.12 w=10.17 l=0.98
X3 VDD2.t7 VN.t0 VTAIL.t0 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X4 B.t8 B.t6 B.t7 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=0 ps=0 w=10.17 l=0.98
X5 VDD1.t5 VP.t2 VTAIL.t13 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X6 VDD1.t1 VP.t3 VTAIL.t12 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X7 VTAIL.t11 VP.t4 VDD1.t2 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=1.67805 ps=10.5 w=10.17 l=0.98
X8 VDD1.t0 VP.t5 VTAIL.t10 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=3.9663 ps=21.12 w=10.17 l=0.98
X9 VDD2.t6 VN.t1 VTAIL.t5 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=3.9663 ps=21.12 w=10.17 l=0.98
X10 VTAIL.t9 VP.t6 VDD1.t6 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X11 VTAIL.t4 VN.t2 VDD2.t5 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X12 VTAIL.t3 VN.t3 VDD2.t4 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=1.67805 ps=10.5 w=10.17 l=0.98
X13 VDD2.t3 VN.t4 VTAIL.t1 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=3.9663 ps=21.12 w=10.17 l=0.98
X14 B.t5 B.t3 B.t4 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=0 ps=0 w=10.17 l=0.98
X15 VTAIL.t8 VP.t7 VDD1.t3 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X16 B.t2 B.t0 B.t1 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=0 ps=0 w=10.17 l=0.98
X17 VDD2.t2 VN.t5 VTAIL.t7 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X18 VTAIL.t2 VN.t6 VDD2.t1 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=1.67805 pd=10.5 as=1.67805 ps=10.5 w=10.17 l=0.98
X19 VTAIL.t6 VN.t7 VDD2.t0 w_n2280_n3002# sky130_fd_pr__pfet_01v8 ad=3.9663 pd=21.12 as=1.67805 ps=10.5 w=10.17 l=0.98
R0 VP.n5 VP.t0 305.466
R1 VP.n17 VP.t4 290.43
R2 VP.n27 VP.t5 290.43
R3 VP.n14 VP.t1 290.43
R4 VP.n19 VP.t3 250.1
R5 VP.n25 VP.t6 250.1
R6 VP.n12 VP.t7 250.1
R7 VP.n6 VP.t2 250.1
R8 VP.n8 VP.n7 161.3
R9 VP.n9 VP.n4 161.3
R10 VP.n11 VP.n10 161.3
R11 VP.n13 VP.n3 161.3
R12 VP.n26 VP.n0 161.3
R13 VP.n24 VP.n23 161.3
R14 VP.n22 VP.n1 161.3
R15 VP.n21 VP.n20 161.3
R16 VP.n18 VP.n2 161.3
R17 VP.n15 VP.n14 80.6037
R18 VP.n28 VP.n27 80.6037
R19 VP.n17 VP.n16 80.6037
R20 VP.n18 VP.n17 55.2959
R21 VP.n27 VP.n26 55.2959
R22 VP.n14 VP.n13 55.2959
R23 VP.n6 VP.n5 46.8653
R24 VP.n8 VP.n5 44.049
R25 VP.n16 VP.n15 42.115
R26 VP.n20 VP.n1 40.4934
R27 VP.n24 VP.n1 40.4934
R28 VP.n11 VP.n4 40.4934
R29 VP.n7 VP.n4 40.4934
R30 VP.n19 VP.n18 16.8827
R31 VP.n26 VP.n25 16.8827
R32 VP.n13 VP.n12 16.8827
R33 VP.n20 VP.n19 7.58527
R34 VP.n25 VP.n24 7.58527
R35 VP.n12 VP.n11 7.58527
R36 VP.n7 VP.n6 7.58527
R37 VP.n15 VP.n3 0.285035
R38 VP.n16 VP.n2 0.285035
R39 VP.n28 VP.n0 0.285035
R40 VP.n9 VP.n8 0.189894
R41 VP.n10 VP.n9 0.189894
R42 VP.n10 VP.n3 0.189894
R43 VP.n21 VP.n2 0.189894
R44 VP.n22 VP.n21 0.189894
R45 VP.n23 VP.n22 0.189894
R46 VP.n23 VP.n0 0.189894
R47 VP VP.n28 0.146778
R48 VDD1 VDD1.n0 81.8145
R49 VDD1.n3 VDD1.n2 81.7008
R50 VDD1.n3 VDD1.n1 81.7008
R51 VDD1.n5 VDD1.n4 81.1915
R52 VDD1.n5 VDD1.n3 38.1474
R53 VDD1.n4 VDD1.t3 3.19667
R54 VDD1.n4 VDD1.t4 3.19667
R55 VDD1.n0 VDD1.t7 3.19667
R56 VDD1.n0 VDD1.t5 3.19667
R57 VDD1.n2 VDD1.t6 3.19667
R58 VDD1.n2 VDD1.t0 3.19667
R59 VDD1.n1 VDD1.t2 3.19667
R60 VDD1.n1 VDD1.t1 3.19667
R61 VDD1 VDD1.n5 0.506965
R62 VTAIL.n434 VTAIL.n386 756.745
R63 VTAIL.n50 VTAIL.n2 756.745
R64 VTAIL.n104 VTAIL.n56 756.745
R65 VTAIL.n160 VTAIL.n112 756.745
R66 VTAIL.n380 VTAIL.n332 756.745
R67 VTAIL.n324 VTAIL.n276 756.745
R68 VTAIL.n270 VTAIL.n222 756.745
R69 VTAIL.n214 VTAIL.n166 756.745
R70 VTAIL.n402 VTAIL.n401 585
R71 VTAIL.n407 VTAIL.n406 585
R72 VTAIL.n409 VTAIL.n408 585
R73 VTAIL.n398 VTAIL.n397 585
R74 VTAIL.n415 VTAIL.n414 585
R75 VTAIL.n417 VTAIL.n416 585
R76 VTAIL.n394 VTAIL.n393 585
R77 VTAIL.n424 VTAIL.n423 585
R78 VTAIL.n425 VTAIL.n392 585
R79 VTAIL.n427 VTAIL.n426 585
R80 VTAIL.n390 VTAIL.n389 585
R81 VTAIL.n433 VTAIL.n432 585
R82 VTAIL.n435 VTAIL.n434 585
R83 VTAIL.n18 VTAIL.n17 585
R84 VTAIL.n23 VTAIL.n22 585
R85 VTAIL.n25 VTAIL.n24 585
R86 VTAIL.n14 VTAIL.n13 585
R87 VTAIL.n31 VTAIL.n30 585
R88 VTAIL.n33 VTAIL.n32 585
R89 VTAIL.n10 VTAIL.n9 585
R90 VTAIL.n40 VTAIL.n39 585
R91 VTAIL.n41 VTAIL.n8 585
R92 VTAIL.n43 VTAIL.n42 585
R93 VTAIL.n6 VTAIL.n5 585
R94 VTAIL.n49 VTAIL.n48 585
R95 VTAIL.n51 VTAIL.n50 585
R96 VTAIL.n72 VTAIL.n71 585
R97 VTAIL.n77 VTAIL.n76 585
R98 VTAIL.n79 VTAIL.n78 585
R99 VTAIL.n68 VTAIL.n67 585
R100 VTAIL.n85 VTAIL.n84 585
R101 VTAIL.n87 VTAIL.n86 585
R102 VTAIL.n64 VTAIL.n63 585
R103 VTAIL.n94 VTAIL.n93 585
R104 VTAIL.n95 VTAIL.n62 585
R105 VTAIL.n97 VTAIL.n96 585
R106 VTAIL.n60 VTAIL.n59 585
R107 VTAIL.n103 VTAIL.n102 585
R108 VTAIL.n105 VTAIL.n104 585
R109 VTAIL.n128 VTAIL.n127 585
R110 VTAIL.n133 VTAIL.n132 585
R111 VTAIL.n135 VTAIL.n134 585
R112 VTAIL.n124 VTAIL.n123 585
R113 VTAIL.n141 VTAIL.n140 585
R114 VTAIL.n143 VTAIL.n142 585
R115 VTAIL.n120 VTAIL.n119 585
R116 VTAIL.n150 VTAIL.n149 585
R117 VTAIL.n151 VTAIL.n118 585
R118 VTAIL.n153 VTAIL.n152 585
R119 VTAIL.n116 VTAIL.n115 585
R120 VTAIL.n159 VTAIL.n158 585
R121 VTAIL.n161 VTAIL.n160 585
R122 VTAIL.n381 VTAIL.n380 585
R123 VTAIL.n379 VTAIL.n378 585
R124 VTAIL.n336 VTAIL.n335 585
R125 VTAIL.n373 VTAIL.n372 585
R126 VTAIL.n371 VTAIL.n338 585
R127 VTAIL.n370 VTAIL.n369 585
R128 VTAIL.n341 VTAIL.n339 585
R129 VTAIL.n364 VTAIL.n363 585
R130 VTAIL.n362 VTAIL.n361 585
R131 VTAIL.n345 VTAIL.n344 585
R132 VTAIL.n356 VTAIL.n355 585
R133 VTAIL.n354 VTAIL.n353 585
R134 VTAIL.n349 VTAIL.n348 585
R135 VTAIL.n325 VTAIL.n324 585
R136 VTAIL.n323 VTAIL.n322 585
R137 VTAIL.n280 VTAIL.n279 585
R138 VTAIL.n317 VTAIL.n316 585
R139 VTAIL.n315 VTAIL.n282 585
R140 VTAIL.n314 VTAIL.n313 585
R141 VTAIL.n285 VTAIL.n283 585
R142 VTAIL.n308 VTAIL.n307 585
R143 VTAIL.n306 VTAIL.n305 585
R144 VTAIL.n289 VTAIL.n288 585
R145 VTAIL.n300 VTAIL.n299 585
R146 VTAIL.n298 VTAIL.n297 585
R147 VTAIL.n293 VTAIL.n292 585
R148 VTAIL.n271 VTAIL.n270 585
R149 VTAIL.n269 VTAIL.n268 585
R150 VTAIL.n226 VTAIL.n225 585
R151 VTAIL.n263 VTAIL.n262 585
R152 VTAIL.n261 VTAIL.n228 585
R153 VTAIL.n260 VTAIL.n259 585
R154 VTAIL.n231 VTAIL.n229 585
R155 VTAIL.n254 VTAIL.n253 585
R156 VTAIL.n252 VTAIL.n251 585
R157 VTAIL.n235 VTAIL.n234 585
R158 VTAIL.n246 VTAIL.n245 585
R159 VTAIL.n244 VTAIL.n243 585
R160 VTAIL.n239 VTAIL.n238 585
R161 VTAIL.n215 VTAIL.n214 585
R162 VTAIL.n213 VTAIL.n212 585
R163 VTAIL.n170 VTAIL.n169 585
R164 VTAIL.n207 VTAIL.n206 585
R165 VTAIL.n205 VTAIL.n172 585
R166 VTAIL.n204 VTAIL.n203 585
R167 VTAIL.n175 VTAIL.n173 585
R168 VTAIL.n198 VTAIL.n197 585
R169 VTAIL.n196 VTAIL.n195 585
R170 VTAIL.n179 VTAIL.n178 585
R171 VTAIL.n190 VTAIL.n189 585
R172 VTAIL.n188 VTAIL.n187 585
R173 VTAIL.n183 VTAIL.n182 585
R174 VTAIL.n403 VTAIL.t1 329.038
R175 VTAIL.n19 VTAIL.t6 329.038
R176 VTAIL.n73 VTAIL.t10 329.038
R177 VTAIL.n129 VTAIL.t11 329.038
R178 VTAIL.n350 VTAIL.t14 329.038
R179 VTAIL.n294 VTAIL.t15 329.038
R180 VTAIL.n240 VTAIL.t5 329.038
R181 VTAIL.n184 VTAIL.t3 329.038
R182 VTAIL.n407 VTAIL.n401 171.744
R183 VTAIL.n408 VTAIL.n407 171.744
R184 VTAIL.n408 VTAIL.n397 171.744
R185 VTAIL.n415 VTAIL.n397 171.744
R186 VTAIL.n416 VTAIL.n415 171.744
R187 VTAIL.n416 VTAIL.n393 171.744
R188 VTAIL.n424 VTAIL.n393 171.744
R189 VTAIL.n425 VTAIL.n424 171.744
R190 VTAIL.n426 VTAIL.n425 171.744
R191 VTAIL.n426 VTAIL.n389 171.744
R192 VTAIL.n433 VTAIL.n389 171.744
R193 VTAIL.n434 VTAIL.n433 171.744
R194 VTAIL.n23 VTAIL.n17 171.744
R195 VTAIL.n24 VTAIL.n23 171.744
R196 VTAIL.n24 VTAIL.n13 171.744
R197 VTAIL.n31 VTAIL.n13 171.744
R198 VTAIL.n32 VTAIL.n31 171.744
R199 VTAIL.n32 VTAIL.n9 171.744
R200 VTAIL.n40 VTAIL.n9 171.744
R201 VTAIL.n41 VTAIL.n40 171.744
R202 VTAIL.n42 VTAIL.n41 171.744
R203 VTAIL.n42 VTAIL.n5 171.744
R204 VTAIL.n49 VTAIL.n5 171.744
R205 VTAIL.n50 VTAIL.n49 171.744
R206 VTAIL.n77 VTAIL.n71 171.744
R207 VTAIL.n78 VTAIL.n77 171.744
R208 VTAIL.n78 VTAIL.n67 171.744
R209 VTAIL.n85 VTAIL.n67 171.744
R210 VTAIL.n86 VTAIL.n85 171.744
R211 VTAIL.n86 VTAIL.n63 171.744
R212 VTAIL.n94 VTAIL.n63 171.744
R213 VTAIL.n95 VTAIL.n94 171.744
R214 VTAIL.n96 VTAIL.n95 171.744
R215 VTAIL.n96 VTAIL.n59 171.744
R216 VTAIL.n103 VTAIL.n59 171.744
R217 VTAIL.n104 VTAIL.n103 171.744
R218 VTAIL.n133 VTAIL.n127 171.744
R219 VTAIL.n134 VTAIL.n133 171.744
R220 VTAIL.n134 VTAIL.n123 171.744
R221 VTAIL.n141 VTAIL.n123 171.744
R222 VTAIL.n142 VTAIL.n141 171.744
R223 VTAIL.n142 VTAIL.n119 171.744
R224 VTAIL.n150 VTAIL.n119 171.744
R225 VTAIL.n151 VTAIL.n150 171.744
R226 VTAIL.n152 VTAIL.n151 171.744
R227 VTAIL.n152 VTAIL.n115 171.744
R228 VTAIL.n159 VTAIL.n115 171.744
R229 VTAIL.n160 VTAIL.n159 171.744
R230 VTAIL.n380 VTAIL.n379 171.744
R231 VTAIL.n379 VTAIL.n335 171.744
R232 VTAIL.n372 VTAIL.n335 171.744
R233 VTAIL.n372 VTAIL.n371 171.744
R234 VTAIL.n371 VTAIL.n370 171.744
R235 VTAIL.n370 VTAIL.n339 171.744
R236 VTAIL.n363 VTAIL.n339 171.744
R237 VTAIL.n363 VTAIL.n362 171.744
R238 VTAIL.n362 VTAIL.n344 171.744
R239 VTAIL.n355 VTAIL.n344 171.744
R240 VTAIL.n355 VTAIL.n354 171.744
R241 VTAIL.n354 VTAIL.n348 171.744
R242 VTAIL.n324 VTAIL.n323 171.744
R243 VTAIL.n323 VTAIL.n279 171.744
R244 VTAIL.n316 VTAIL.n279 171.744
R245 VTAIL.n316 VTAIL.n315 171.744
R246 VTAIL.n315 VTAIL.n314 171.744
R247 VTAIL.n314 VTAIL.n283 171.744
R248 VTAIL.n307 VTAIL.n283 171.744
R249 VTAIL.n307 VTAIL.n306 171.744
R250 VTAIL.n306 VTAIL.n288 171.744
R251 VTAIL.n299 VTAIL.n288 171.744
R252 VTAIL.n299 VTAIL.n298 171.744
R253 VTAIL.n298 VTAIL.n292 171.744
R254 VTAIL.n270 VTAIL.n269 171.744
R255 VTAIL.n269 VTAIL.n225 171.744
R256 VTAIL.n262 VTAIL.n225 171.744
R257 VTAIL.n262 VTAIL.n261 171.744
R258 VTAIL.n261 VTAIL.n260 171.744
R259 VTAIL.n260 VTAIL.n229 171.744
R260 VTAIL.n253 VTAIL.n229 171.744
R261 VTAIL.n253 VTAIL.n252 171.744
R262 VTAIL.n252 VTAIL.n234 171.744
R263 VTAIL.n245 VTAIL.n234 171.744
R264 VTAIL.n245 VTAIL.n244 171.744
R265 VTAIL.n244 VTAIL.n238 171.744
R266 VTAIL.n214 VTAIL.n213 171.744
R267 VTAIL.n213 VTAIL.n169 171.744
R268 VTAIL.n206 VTAIL.n169 171.744
R269 VTAIL.n206 VTAIL.n205 171.744
R270 VTAIL.n205 VTAIL.n204 171.744
R271 VTAIL.n204 VTAIL.n173 171.744
R272 VTAIL.n197 VTAIL.n173 171.744
R273 VTAIL.n197 VTAIL.n196 171.744
R274 VTAIL.n196 VTAIL.n178 171.744
R275 VTAIL.n189 VTAIL.n178 171.744
R276 VTAIL.n189 VTAIL.n188 171.744
R277 VTAIL.n188 VTAIL.n182 171.744
R278 VTAIL.t1 VTAIL.n401 85.8723
R279 VTAIL.t6 VTAIL.n17 85.8723
R280 VTAIL.t10 VTAIL.n71 85.8723
R281 VTAIL.t11 VTAIL.n127 85.8723
R282 VTAIL.t14 VTAIL.n348 85.8723
R283 VTAIL.t15 VTAIL.n292 85.8723
R284 VTAIL.t5 VTAIL.n238 85.8723
R285 VTAIL.t3 VTAIL.n182 85.8723
R286 VTAIL.n331 VTAIL.n330 64.5129
R287 VTAIL.n221 VTAIL.n220 64.5129
R288 VTAIL.n1 VTAIL.n0 64.5127
R289 VTAIL.n111 VTAIL.n110 64.5127
R290 VTAIL.n439 VTAIL.n438 36.2581
R291 VTAIL.n55 VTAIL.n54 36.2581
R292 VTAIL.n109 VTAIL.n108 36.2581
R293 VTAIL.n165 VTAIL.n164 36.2581
R294 VTAIL.n385 VTAIL.n384 36.2581
R295 VTAIL.n329 VTAIL.n328 36.2581
R296 VTAIL.n275 VTAIL.n274 36.2581
R297 VTAIL.n219 VTAIL.n218 36.2581
R298 VTAIL.n439 VTAIL.n385 22.2634
R299 VTAIL.n219 VTAIL.n165 22.2634
R300 VTAIL.n427 VTAIL.n392 13.1884
R301 VTAIL.n43 VTAIL.n8 13.1884
R302 VTAIL.n97 VTAIL.n62 13.1884
R303 VTAIL.n153 VTAIL.n118 13.1884
R304 VTAIL.n373 VTAIL.n338 13.1884
R305 VTAIL.n317 VTAIL.n282 13.1884
R306 VTAIL.n263 VTAIL.n228 13.1884
R307 VTAIL.n207 VTAIL.n172 13.1884
R308 VTAIL.n423 VTAIL.n422 12.8005
R309 VTAIL.n428 VTAIL.n390 12.8005
R310 VTAIL.n39 VTAIL.n38 12.8005
R311 VTAIL.n44 VTAIL.n6 12.8005
R312 VTAIL.n93 VTAIL.n92 12.8005
R313 VTAIL.n98 VTAIL.n60 12.8005
R314 VTAIL.n149 VTAIL.n148 12.8005
R315 VTAIL.n154 VTAIL.n116 12.8005
R316 VTAIL.n374 VTAIL.n336 12.8005
R317 VTAIL.n369 VTAIL.n340 12.8005
R318 VTAIL.n318 VTAIL.n280 12.8005
R319 VTAIL.n313 VTAIL.n284 12.8005
R320 VTAIL.n264 VTAIL.n226 12.8005
R321 VTAIL.n259 VTAIL.n230 12.8005
R322 VTAIL.n208 VTAIL.n170 12.8005
R323 VTAIL.n203 VTAIL.n174 12.8005
R324 VTAIL.n421 VTAIL.n394 12.0247
R325 VTAIL.n432 VTAIL.n431 12.0247
R326 VTAIL.n37 VTAIL.n10 12.0247
R327 VTAIL.n48 VTAIL.n47 12.0247
R328 VTAIL.n91 VTAIL.n64 12.0247
R329 VTAIL.n102 VTAIL.n101 12.0247
R330 VTAIL.n147 VTAIL.n120 12.0247
R331 VTAIL.n158 VTAIL.n157 12.0247
R332 VTAIL.n378 VTAIL.n377 12.0247
R333 VTAIL.n368 VTAIL.n341 12.0247
R334 VTAIL.n322 VTAIL.n321 12.0247
R335 VTAIL.n312 VTAIL.n285 12.0247
R336 VTAIL.n268 VTAIL.n267 12.0247
R337 VTAIL.n258 VTAIL.n231 12.0247
R338 VTAIL.n212 VTAIL.n211 12.0247
R339 VTAIL.n202 VTAIL.n175 12.0247
R340 VTAIL.n418 VTAIL.n417 11.249
R341 VTAIL.n435 VTAIL.n388 11.249
R342 VTAIL.n34 VTAIL.n33 11.249
R343 VTAIL.n51 VTAIL.n4 11.249
R344 VTAIL.n88 VTAIL.n87 11.249
R345 VTAIL.n105 VTAIL.n58 11.249
R346 VTAIL.n144 VTAIL.n143 11.249
R347 VTAIL.n161 VTAIL.n114 11.249
R348 VTAIL.n381 VTAIL.n334 11.249
R349 VTAIL.n365 VTAIL.n364 11.249
R350 VTAIL.n325 VTAIL.n278 11.249
R351 VTAIL.n309 VTAIL.n308 11.249
R352 VTAIL.n271 VTAIL.n224 11.249
R353 VTAIL.n255 VTAIL.n254 11.249
R354 VTAIL.n215 VTAIL.n168 11.249
R355 VTAIL.n199 VTAIL.n198 11.249
R356 VTAIL.n403 VTAIL.n402 10.7239
R357 VTAIL.n19 VTAIL.n18 10.7239
R358 VTAIL.n73 VTAIL.n72 10.7239
R359 VTAIL.n129 VTAIL.n128 10.7239
R360 VTAIL.n350 VTAIL.n349 10.7239
R361 VTAIL.n294 VTAIL.n293 10.7239
R362 VTAIL.n240 VTAIL.n239 10.7239
R363 VTAIL.n184 VTAIL.n183 10.7239
R364 VTAIL.n414 VTAIL.n396 10.4732
R365 VTAIL.n436 VTAIL.n386 10.4732
R366 VTAIL.n30 VTAIL.n12 10.4732
R367 VTAIL.n52 VTAIL.n2 10.4732
R368 VTAIL.n84 VTAIL.n66 10.4732
R369 VTAIL.n106 VTAIL.n56 10.4732
R370 VTAIL.n140 VTAIL.n122 10.4732
R371 VTAIL.n162 VTAIL.n112 10.4732
R372 VTAIL.n382 VTAIL.n332 10.4732
R373 VTAIL.n361 VTAIL.n343 10.4732
R374 VTAIL.n326 VTAIL.n276 10.4732
R375 VTAIL.n305 VTAIL.n287 10.4732
R376 VTAIL.n272 VTAIL.n222 10.4732
R377 VTAIL.n251 VTAIL.n233 10.4732
R378 VTAIL.n216 VTAIL.n166 10.4732
R379 VTAIL.n195 VTAIL.n177 10.4732
R380 VTAIL.n413 VTAIL.n398 9.69747
R381 VTAIL.n29 VTAIL.n14 9.69747
R382 VTAIL.n83 VTAIL.n68 9.69747
R383 VTAIL.n139 VTAIL.n124 9.69747
R384 VTAIL.n360 VTAIL.n345 9.69747
R385 VTAIL.n304 VTAIL.n289 9.69747
R386 VTAIL.n250 VTAIL.n235 9.69747
R387 VTAIL.n194 VTAIL.n179 9.69747
R388 VTAIL.n438 VTAIL.n437 9.45567
R389 VTAIL.n54 VTAIL.n53 9.45567
R390 VTAIL.n108 VTAIL.n107 9.45567
R391 VTAIL.n164 VTAIL.n163 9.45567
R392 VTAIL.n384 VTAIL.n383 9.45567
R393 VTAIL.n328 VTAIL.n327 9.45567
R394 VTAIL.n274 VTAIL.n273 9.45567
R395 VTAIL.n218 VTAIL.n217 9.45567
R396 VTAIL.n437 VTAIL.n436 9.3005
R397 VTAIL.n388 VTAIL.n387 9.3005
R398 VTAIL.n431 VTAIL.n430 9.3005
R399 VTAIL.n429 VTAIL.n428 9.3005
R400 VTAIL.n405 VTAIL.n404 9.3005
R401 VTAIL.n400 VTAIL.n399 9.3005
R402 VTAIL.n411 VTAIL.n410 9.3005
R403 VTAIL.n413 VTAIL.n412 9.3005
R404 VTAIL.n396 VTAIL.n395 9.3005
R405 VTAIL.n419 VTAIL.n418 9.3005
R406 VTAIL.n421 VTAIL.n420 9.3005
R407 VTAIL.n422 VTAIL.n391 9.3005
R408 VTAIL.n53 VTAIL.n52 9.3005
R409 VTAIL.n4 VTAIL.n3 9.3005
R410 VTAIL.n47 VTAIL.n46 9.3005
R411 VTAIL.n45 VTAIL.n44 9.3005
R412 VTAIL.n21 VTAIL.n20 9.3005
R413 VTAIL.n16 VTAIL.n15 9.3005
R414 VTAIL.n27 VTAIL.n26 9.3005
R415 VTAIL.n29 VTAIL.n28 9.3005
R416 VTAIL.n12 VTAIL.n11 9.3005
R417 VTAIL.n35 VTAIL.n34 9.3005
R418 VTAIL.n37 VTAIL.n36 9.3005
R419 VTAIL.n38 VTAIL.n7 9.3005
R420 VTAIL.n107 VTAIL.n106 9.3005
R421 VTAIL.n58 VTAIL.n57 9.3005
R422 VTAIL.n101 VTAIL.n100 9.3005
R423 VTAIL.n99 VTAIL.n98 9.3005
R424 VTAIL.n75 VTAIL.n74 9.3005
R425 VTAIL.n70 VTAIL.n69 9.3005
R426 VTAIL.n81 VTAIL.n80 9.3005
R427 VTAIL.n83 VTAIL.n82 9.3005
R428 VTAIL.n66 VTAIL.n65 9.3005
R429 VTAIL.n89 VTAIL.n88 9.3005
R430 VTAIL.n91 VTAIL.n90 9.3005
R431 VTAIL.n92 VTAIL.n61 9.3005
R432 VTAIL.n163 VTAIL.n162 9.3005
R433 VTAIL.n114 VTAIL.n113 9.3005
R434 VTAIL.n157 VTAIL.n156 9.3005
R435 VTAIL.n155 VTAIL.n154 9.3005
R436 VTAIL.n131 VTAIL.n130 9.3005
R437 VTAIL.n126 VTAIL.n125 9.3005
R438 VTAIL.n137 VTAIL.n136 9.3005
R439 VTAIL.n139 VTAIL.n138 9.3005
R440 VTAIL.n122 VTAIL.n121 9.3005
R441 VTAIL.n145 VTAIL.n144 9.3005
R442 VTAIL.n147 VTAIL.n146 9.3005
R443 VTAIL.n148 VTAIL.n117 9.3005
R444 VTAIL.n352 VTAIL.n351 9.3005
R445 VTAIL.n347 VTAIL.n346 9.3005
R446 VTAIL.n358 VTAIL.n357 9.3005
R447 VTAIL.n360 VTAIL.n359 9.3005
R448 VTAIL.n343 VTAIL.n342 9.3005
R449 VTAIL.n366 VTAIL.n365 9.3005
R450 VTAIL.n368 VTAIL.n367 9.3005
R451 VTAIL.n340 VTAIL.n337 9.3005
R452 VTAIL.n383 VTAIL.n382 9.3005
R453 VTAIL.n334 VTAIL.n333 9.3005
R454 VTAIL.n377 VTAIL.n376 9.3005
R455 VTAIL.n375 VTAIL.n374 9.3005
R456 VTAIL.n296 VTAIL.n295 9.3005
R457 VTAIL.n291 VTAIL.n290 9.3005
R458 VTAIL.n302 VTAIL.n301 9.3005
R459 VTAIL.n304 VTAIL.n303 9.3005
R460 VTAIL.n287 VTAIL.n286 9.3005
R461 VTAIL.n310 VTAIL.n309 9.3005
R462 VTAIL.n312 VTAIL.n311 9.3005
R463 VTAIL.n284 VTAIL.n281 9.3005
R464 VTAIL.n327 VTAIL.n326 9.3005
R465 VTAIL.n278 VTAIL.n277 9.3005
R466 VTAIL.n321 VTAIL.n320 9.3005
R467 VTAIL.n319 VTAIL.n318 9.3005
R468 VTAIL.n242 VTAIL.n241 9.3005
R469 VTAIL.n237 VTAIL.n236 9.3005
R470 VTAIL.n248 VTAIL.n247 9.3005
R471 VTAIL.n250 VTAIL.n249 9.3005
R472 VTAIL.n233 VTAIL.n232 9.3005
R473 VTAIL.n256 VTAIL.n255 9.3005
R474 VTAIL.n258 VTAIL.n257 9.3005
R475 VTAIL.n230 VTAIL.n227 9.3005
R476 VTAIL.n273 VTAIL.n272 9.3005
R477 VTAIL.n224 VTAIL.n223 9.3005
R478 VTAIL.n267 VTAIL.n266 9.3005
R479 VTAIL.n265 VTAIL.n264 9.3005
R480 VTAIL.n186 VTAIL.n185 9.3005
R481 VTAIL.n181 VTAIL.n180 9.3005
R482 VTAIL.n192 VTAIL.n191 9.3005
R483 VTAIL.n194 VTAIL.n193 9.3005
R484 VTAIL.n177 VTAIL.n176 9.3005
R485 VTAIL.n200 VTAIL.n199 9.3005
R486 VTAIL.n202 VTAIL.n201 9.3005
R487 VTAIL.n174 VTAIL.n171 9.3005
R488 VTAIL.n217 VTAIL.n216 9.3005
R489 VTAIL.n168 VTAIL.n167 9.3005
R490 VTAIL.n211 VTAIL.n210 9.3005
R491 VTAIL.n209 VTAIL.n208 9.3005
R492 VTAIL.n410 VTAIL.n409 8.92171
R493 VTAIL.n26 VTAIL.n25 8.92171
R494 VTAIL.n80 VTAIL.n79 8.92171
R495 VTAIL.n136 VTAIL.n135 8.92171
R496 VTAIL.n357 VTAIL.n356 8.92171
R497 VTAIL.n301 VTAIL.n300 8.92171
R498 VTAIL.n247 VTAIL.n246 8.92171
R499 VTAIL.n191 VTAIL.n190 8.92171
R500 VTAIL.n406 VTAIL.n400 8.14595
R501 VTAIL.n22 VTAIL.n16 8.14595
R502 VTAIL.n76 VTAIL.n70 8.14595
R503 VTAIL.n132 VTAIL.n126 8.14595
R504 VTAIL.n353 VTAIL.n347 8.14595
R505 VTAIL.n297 VTAIL.n291 8.14595
R506 VTAIL.n243 VTAIL.n237 8.14595
R507 VTAIL.n187 VTAIL.n181 8.14595
R508 VTAIL.n405 VTAIL.n402 7.3702
R509 VTAIL.n21 VTAIL.n18 7.3702
R510 VTAIL.n75 VTAIL.n72 7.3702
R511 VTAIL.n131 VTAIL.n128 7.3702
R512 VTAIL.n352 VTAIL.n349 7.3702
R513 VTAIL.n296 VTAIL.n293 7.3702
R514 VTAIL.n242 VTAIL.n239 7.3702
R515 VTAIL.n186 VTAIL.n183 7.3702
R516 VTAIL.n406 VTAIL.n405 5.81868
R517 VTAIL.n22 VTAIL.n21 5.81868
R518 VTAIL.n76 VTAIL.n75 5.81868
R519 VTAIL.n132 VTAIL.n131 5.81868
R520 VTAIL.n353 VTAIL.n352 5.81868
R521 VTAIL.n297 VTAIL.n296 5.81868
R522 VTAIL.n243 VTAIL.n242 5.81868
R523 VTAIL.n187 VTAIL.n186 5.81868
R524 VTAIL.n409 VTAIL.n400 5.04292
R525 VTAIL.n25 VTAIL.n16 5.04292
R526 VTAIL.n79 VTAIL.n70 5.04292
R527 VTAIL.n135 VTAIL.n126 5.04292
R528 VTAIL.n356 VTAIL.n347 5.04292
R529 VTAIL.n300 VTAIL.n291 5.04292
R530 VTAIL.n246 VTAIL.n237 5.04292
R531 VTAIL.n190 VTAIL.n181 5.04292
R532 VTAIL.n410 VTAIL.n398 4.26717
R533 VTAIL.n26 VTAIL.n14 4.26717
R534 VTAIL.n80 VTAIL.n68 4.26717
R535 VTAIL.n136 VTAIL.n124 4.26717
R536 VTAIL.n357 VTAIL.n345 4.26717
R537 VTAIL.n301 VTAIL.n289 4.26717
R538 VTAIL.n247 VTAIL.n235 4.26717
R539 VTAIL.n191 VTAIL.n179 4.26717
R540 VTAIL.n414 VTAIL.n413 3.49141
R541 VTAIL.n438 VTAIL.n386 3.49141
R542 VTAIL.n30 VTAIL.n29 3.49141
R543 VTAIL.n54 VTAIL.n2 3.49141
R544 VTAIL.n84 VTAIL.n83 3.49141
R545 VTAIL.n108 VTAIL.n56 3.49141
R546 VTAIL.n140 VTAIL.n139 3.49141
R547 VTAIL.n164 VTAIL.n112 3.49141
R548 VTAIL.n384 VTAIL.n332 3.49141
R549 VTAIL.n361 VTAIL.n360 3.49141
R550 VTAIL.n328 VTAIL.n276 3.49141
R551 VTAIL.n305 VTAIL.n304 3.49141
R552 VTAIL.n274 VTAIL.n222 3.49141
R553 VTAIL.n251 VTAIL.n250 3.49141
R554 VTAIL.n218 VTAIL.n166 3.49141
R555 VTAIL.n195 VTAIL.n194 3.49141
R556 VTAIL.n0 VTAIL.t7 3.19667
R557 VTAIL.n0 VTAIL.t4 3.19667
R558 VTAIL.n110 VTAIL.t12 3.19667
R559 VTAIL.n110 VTAIL.t9 3.19667
R560 VTAIL.n330 VTAIL.t13 3.19667
R561 VTAIL.n330 VTAIL.t8 3.19667
R562 VTAIL.n220 VTAIL.t0 3.19667
R563 VTAIL.n220 VTAIL.t2 3.19667
R564 VTAIL.n417 VTAIL.n396 2.71565
R565 VTAIL.n436 VTAIL.n435 2.71565
R566 VTAIL.n33 VTAIL.n12 2.71565
R567 VTAIL.n52 VTAIL.n51 2.71565
R568 VTAIL.n87 VTAIL.n66 2.71565
R569 VTAIL.n106 VTAIL.n105 2.71565
R570 VTAIL.n143 VTAIL.n122 2.71565
R571 VTAIL.n162 VTAIL.n161 2.71565
R572 VTAIL.n382 VTAIL.n381 2.71565
R573 VTAIL.n364 VTAIL.n343 2.71565
R574 VTAIL.n326 VTAIL.n325 2.71565
R575 VTAIL.n308 VTAIL.n287 2.71565
R576 VTAIL.n272 VTAIL.n271 2.71565
R577 VTAIL.n254 VTAIL.n233 2.71565
R578 VTAIL.n216 VTAIL.n215 2.71565
R579 VTAIL.n198 VTAIL.n177 2.71565
R580 VTAIL.n404 VTAIL.n403 2.41283
R581 VTAIL.n20 VTAIL.n19 2.41283
R582 VTAIL.n74 VTAIL.n73 2.41283
R583 VTAIL.n130 VTAIL.n129 2.41283
R584 VTAIL.n351 VTAIL.n350 2.41283
R585 VTAIL.n295 VTAIL.n294 2.41283
R586 VTAIL.n241 VTAIL.n240 2.41283
R587 VTAIL.n185 VTAIL.n184 2.41283
R588 VTAIL.n418 VTAIL.n394 1.93989
R589 VTAIL.n432 VTAIL.n388 1.93989
R590 VTAIL.n34 VTAIL.n10 1.93989
R591 VTAIL.n48 VTAIL.n4 1.93989
R592 VTAIL.n88 VTAIL.n64 1.93989
R593 VTAIL.n102 VTAIL.n58 1.93989
R594 VTAIL.n144 VTAIL.n120 1.93989
R595 VTAIL.n158 VTAIL.n114 1.93989
R596 VTAIL.n378 VTAIL.n334 1.93989
R597 VTAIL.n365 VTAIL.n341 1.93989
R598 VTAIL.n322 VTAIL.n278 1.93989
R599 VTAIL.n309 VTAIL.n285 1.93989
R600 VTAIL.n268 VTAIL.n224 1.93989
R601 VTAIL.n255 VTAIL.n231 1.93989
R602 VTAIL.n212 VTAIL.n168 1.93989
R603 VTAIL.n199 VTAIL.n175 1.93989
R604 VTAIL.n423 VTAIL.n421 1.16414
R605 VTAIL.n431 VTAIL.n390 1.16414
R606 VTAIL.n39 VTAIL.n37 1.16414
R607 VTAIL.n47 VTAIL.n6 1.16414
R608 VTAIL.n93 VTAIL.n91 1.16414
R609 VTAIL.n101 VTAIL.n60 1.16414
R610 VTAIL.n149 VTAIL.n147 1.16414
R611 VTAIL.n157 VTAIL.n116 1.16414
R612 VTAIL.n377 VTAIL.n336 1.16414
R613 VTAIL.n369 VTAIL.n368 1.16414
R614 VTAIL.n321 VTAIL.n280 1.16414
R615 VTAIL.n313 VTAIL.n312 1.16414
R616 VTAIL.n267 VTAIL.n226 1.16414
R617 VTAIL.n259 VTAIL.n258 1.16414
R618 VTAIL.n211 VTAIL.n170 1.16414
R619 VTAIL.n203 VTAIL.n202 1.16414
R620 VTAIL.n221 VTAIL.n219 1.12981
R621 VTAIL.n275 VTAIL.n221 1.12981
R622 VTAIL.n331 VTAIL.n329 1.12981
R623 VTAIL.n385 VTAIL.n331 1.12981
R624 VTAIL.n165 VTAIL.n111 1.12981
R625 VTAIL.n111 VTAIL.n109 1.12981
R626 VTAIL.n55 VTAIL.n1 1.12981
R627 VTAIL VTAIL.n439 1.07162
R628 VTAIL.n329 VTAIL.n275 0.470328
R629 VTAIL.n109 VTAIL.n55 0.470328
R630 VTAIL.n422 VTAIL.n392 0.388379
R631 VTAIL.n428 VTAIL.n427 0.388379
R632 VTAIL.n38 VTAIL.n8 0.388379
R633 VTAIL.n44 VTAIL.n43 0.388379
R634 VTAIL.n92 VTAIL.n62 0.388379
R635 VTAIL.n98 VTAIL.n97 0.388379
R636 VTAIL.n148 VTAIL.n118 0.388379
R637 VTAIL.n154 VTAIL.n153 0.388379
R638 VTAIL.n374 VTAIL.n373 0.388379
R639 VTAIL.n340 VTAIL.n338 0.388379
R640 VTAIL.n318 VTAIL.n317 0.388379
R641 VTAIL.n284 VTAIL.n282 0.388379
R642 VTAIL.n264 VTAIL.n263 0.388379
R643 VTAIL.n230 VTAIL.n228 0.388379
R644 VTAIL.n208 VTAIL.n207 0.388379
R645 VTAIL.n174 VTAIL.n172 0.388379
R646 VTAIL.n404 VTAIL.n399 0.155672
R647 VTAIL.n411 VTAIL.n399 0.155672
R648 VTAIL.n412 VTAIL.n411 0.155672
R649 VTAIL.n412 VTAIL.n395 0.155672
R650 VTAIL.n419 VTAIL.n395 0.155672
R651 VTAIL.n420 VTAIL.n419 0.155672
R652 VTAIL.n420 VTAIL.n391 0.155672
R653 VTAIL.n429 VTAIL.n391 0.155672
R654 VTAIL.n430 VTAIL.n429 0.155672
R655 VTAIL.n430 VTAIL.n387 0.155672
R656 VTAIL.n437 VTAIL.n387 0.155672
R657 VTAIL.n20 VTAIL.n15 0.155672
R658 VTAIL.n27 VTAIL.n15 0.155672
R659 VTAIL.n28 VTAIL.n27 0.155672
R660 VTAIL.n28 VTAIL.n11 0.155672
R661 VTAIL.n35 VTAIL.n11 0.155672
R662 VTAIL.n36 VTAIL.n35 0.155672
R663 VTAIL.n36 VTAIL.n7 0.155672
R664 VTAIL.n45 VTAIL.n7 0.155672
R665 VTAIL.n46 VTAIL.n45 0.155672
R666 VTAIL.n46 VTAIL.n3 0.155672
R667 VTAIL.n53 VTAIL.n3 0.155672
R668 VTAIL.n74 VTAIL.n69 0.155672
R669 VTAIL.n81 VTAIL.n69 0.155672
R670 VTAIL.n82 VTAIL.n81 0.155672
R671 VTAIL.n82 VTAIL.n65 0.155672
R672 VTAIL.n89 VTAIL.n65 0.155672
R673 VTAIL.n90 VTAIL.n89 0.155672
R674 VTAIL.n90 VTAIL.n61 0.155672
R675 VTAIL.n99 VTAIL.n61 0.155672
R676 VTAIL.n100 VTAIL.n99 0.155672
R677 VTAIL.n100 VTAIL.n57 0.155672
R678 VTAIL.n107 VTAIL.n57 0.155672
R679 VTAIL.n130 VTAIL.n125 0.155672
R680 VTAIL.n137 VTAIL.n125 0.155672
R681 VTAIL.n138 VTAIL.n137 0.155672
R682 VTAIL.n138 VTAIL.n121 0.155672
R683 VTAIL.n145 VTAIL.n121 0.155672
R684 VTAIL.n146 VTAIL.n145 0.155672
R685 VTAIL.n146 VTAIL.n117 0.155672
R686 VTAIL.n155 VTAIL.n117 0.155672
R687 VTAIL.n156 VTAIL.n155 0.155672
R688 VTAIL.n156 VTAIL.n113 0.155672
R689 VTAIL.n163 VTAIL.n113 0.155672
R690 VTAIL.n383 VTAIL.n333 0.155672
R691 VTAIL.n376 VTAIL.n333 0.155672
R692 VTAIL.n376 VTAIL.n375 0.155672
R693 VTAIL.n375 VTAIL.n337 0.155672
R694 VTAIL.n367 VTAIL.n337 0.155672
R695 VTAIL.n367 VTAIL.n366 0.155672
R696 VTAIL.n366 VTAIL.n342 0.155672
R697 VTAIL.n359 VTAIL.n342 0.155672
R698 VTAIL.n359 VTAIL.n358 0.155672
R699 VTAIL.n358 VTAIL.n346 0.155672
R700 VTAIL.n351 VTAIL.n346 0.155672
R701 VTAIL.n327 VTAIL.n277 0.155672
R702 VTAIL.n320 VTAIL.n277 0.155672
R703 VTAIL.n320 VTAIL.n319 0.155672
R704 VTAIL.n319 VTAIL.n281 0.155672
R705 VTAIL.n311 VTAIL.n281 0.155672
R706 VTAIL.n311 VTAIL.n310 0.155672
R707 VTAIL.n310 VTAIL.n286 0.155672
R708 VTAIL.n303 VTAIL.n286 0.155672
R709 VTAIL.n303 VTAIL.n302 0.155672
R710 VTAIL.n302 VTAIL.n290 0.155672
R711 VTAIL.n295 VTAIL.n290 0.155672
R712 VTAIL.n273 VTAIL.n223 0.155672
R713 VTAIL.n266 VTAIL.n223 0.155672
R714 VTAIL.n266 VTAIL.n265 0.155672
R715 VTAIL.n265 VTAIL.n227 0.155672
R716 VTAIL.n257 VTAIL.n227 0.155672
R717 VTAIL.n257 VTAIL.n256 0.155672
R718 VTAIL.n256 VTAIL.n232 0.155672
R719 VTAIL.n249 VTAIL.n232 0.155672
R720 VTAIL.n249 VTAIL.n248 0.155672
R721 VTAIL.n248 VTAIL.n236 0.155672
R722 VTAIL.n241 VTAIL.n236 0.155672
R723 VTAIL.n217 VTAIL.n167 0.155672
R724 VTAIL.n210 VTAIL.n167 0.155672
R725 VTAIL.n210 VTAIL.n209 0.155672
R726 VTAIL.n209 VTAIL.n171 0.155672
R727 VTAIL.n201 VTAIL.n171 0.155672
R728 VTAIL.n201 VTAIL.n200 0.155672
R729 VTAIL.n200 VTAIL.n176 0.155672
R730 VTAIL.n193 VTAIL.n176 0.155672
R731 VTAIL.n193 VTAIL.n192 0.155672
R732 VTAIL.n192 VTAIL.n180 0.155672
R733 VTAIL.n185 VTAIL.n180 0.155672
R734 VTAIL VTAIL.n1 0.0586897
R735 B.n311 B.n310 585
R736 B.n309 B.n90 585
R737 B.n308 B.n307 585
R738 B.n306 B.n91 585
R739 B.n305 B.n304 585
R740 B.n303 B.n92 585
R741 B.n302 B.n301 585
R742 B.n300 B.n93 585
R743 B.n299 B.n298 585
R744 B.n297 B.n94 585
R745 B.n296 B.n295 585
R746 B.n294 B.n95 585
R747 B.n293 B.n292 585
R748 B.n291 B.n96 585
R749 B.n290 B.n289 585
R750 B.n288 B.n97 585
R751 B.n287 B.n286 585
R752 B.n285 B.n98 585
R753 B.n284 B.n283 585
R754 B.n282 B.n99 585
R755 B.n281 B.n280 585
R756 B.n279 B.n100 585
R757 B.n278 B.n277 585
R758 B.n276 B.n101 585
R759 B.n275 B.n274 585
R760 B.n273 B.n102 585
R761 B.n272 B.n271 585
R762 B.n270 B.n103 585
R763 B.n269 B.n268 585
R764 B.n267 B.n104 585
R765 B.n266 B.n265 585
R766 B.n264 B.n105 585
R767 B.n263 B.n262 585
R768 B.n261 B.n106 585
R769 B.n260 B.n259 585
R770 B.n258 B.n107 585
R771 B.n257 B.n256 585
R772 B.n252 B.n108 585
R773 B.n251 B.n250 585
R774 B.n249 B.n109 585
R775 B.n248 B.n247 585
R776 B.n246 B.n110 585
R777 B.n245 B.n244 585
R778 B.n243 B.n111 585
R779 B.n242 B.n241 585
R780 B.n240 B.n112 585
R781 B.n238 B.n237 585
R782 B.n236 B.n115 585
R783 B.n235 B.n234 585
R784 B.n233 B.n116 585
R785 B.n232 B.n231 585
R786 B.n230 B.n117 585
R787 B.n229 B.n228 585
R788 B.n227 B.n118 585
R789 B.n226 B.n225 585
R790 B.n224 B.n119 585
R791 B.n223 B.n222 585
R792 B.n221 B.n120 585
R793 B.n220 B.n219 585
R794 B.n218 B.n121 585
R795 B.n217 B.n216 585
R796 B.n215 B.n122 585
R797 B.n214 B.n213 585
R798 B.n212 B.n123 585
R799 B.n211 B.n210 585
R800 B.n209 B.n124 585
R801 B.n208 B.n207 585
R802 B.n206 B.n125 585
R803 B.n205 B.n204 585
R804 B.n203 B.n126 585
R805 B.n202 B.n201 585
R806 B.n200 B.n127 585
R807 B.n199 B.n198 585
R808 B.n197 B.n128 585
R809 B.n196 B.n195 585
R810 B.n194 B.n129 585
R811 B.n193 B.n192 585
R812 B.n191 B.n130 585
R813 B.n190 B.n189 585
R814 B.n188 B.n131 585
R815 B.n187 B.n186 585
R816 B.n185 B.n132 585
R817 B.n312 B.n89 585
R818 B.n314 B.n313 585
R819 B.n315 B.n88 585
R820 B.n317 B.n316 585
R821 B.n318 B.n87 585
R822 B.n320 B.n319 585
R823 B.n321 B.n86 585
R824 B.n323 B.n322 585
R825 B.n324 B.n85 585
R826 B.n326 B.n325 585
R827 B.n327 B.n84 585
R828 B.n329 B.n328 585
R829 B.n330 B.n83 585
R830 B.n332 B.n331 585
R831 B.n333 B.n82 585
R832 B.n335 B.n334 585
R833 B.n336 B.n81 585
R834 B.n338 B.n337 585
R835 B.n339 B.n80 585
R836 B.n341 B.n340 585
R837 B.n342 B.n79 585
R838 B.n344 B.n343 585
R839 B.n345 B.n78 585
R840 B.n347 B.n346 585
R841 B.n348 B.n77 585
R842 B.n350 B.n349 585
R843 B.n351 B.n76 585
R844 B.n353 B.n352 585
R845 B.n354 B.n75 585
R846 B.n356 B.n355 585
R847 B.n357 B.n74 585
R848 B.n359 B.n358 585
R849 B.n360 B.n73 585
R850 B.n362 B.n361 585
R851 B.n363 B.n72 585
R852 B.n365 B.n364 585
R853 B.n366 B.n71 585
R854 B.n368 B.n367 585
R855 B.n369 B.n70 585
R856 B.n371 B.n370 585
R857 B.n372 B.n69 585
R858 B.n374 B.n373 585
R859 B.n375 B.n68 585
R860 B.n377 B.n376 585
R861 B.n378 B.n67 585
R862 B.n380 B.n379 585
R863 B.n381 B.n66 585
R864 B.n383 B.n382 585
R865 B.n384 B.n65 585
R866 B.n386 B.n385 585
R867 B.n387 B.n64 585
R868 B.n389 B.n388 585
R869 B.n390 B.n63 585
R870 B.n392 B.n391 585
R871 B.n393 B.n62 585
R872 B.n395 B.n394 585
R873 B.n519 B.n518 585
R874 B.n517 B.n16 585
R875 B.n516 B.n515 585
R876 B.n514 B.n17 585
R877 B.n513 B.n512 585
R878 B.n511 B.n18 585
R879 B.n510 B.n509 585
R880 B.n508 B.n19 585
R881 B.n507 B.n506 585
R882 B.n505 B.n20 585
R883 B.n504 B.n503 585
R884 B.n502 B.n21 585
R885 B.n501 B.n500 585
R886 B.n499 B.n22 585
R887 B.n498 B.n497 585
R888 B.n496 B.n23 585
R889 B.n495 B.n494 585
R890 B.n493 B.n24 585
R891 B.n492 B.n491 585
R892 B.n490 B.n25 585
R893 B.n489 B.n488 585
R894 B.n487 B.n26 585
R895 B.n486 B.n485 585
R896 B.n484 B.n27 585
R897 B.n483 B.n482 585
R898 B.n481 B.n28 585
R899 B.n480 B.n479 585
R900 B.n478 B.n29 585
R901 B.n477 B.n476 585
R902 B.n475 B.n30 585
R903 B.n474 B.n473 585
R904 B.n472 B.n31 585
R905 B.n471 B.n470 585
R906 B.n469 B.n32 585
R907 B.n468 B.n467 585
R908 B.n466 B.n33 585
R909 B.n464 B.n463 585
R910 B.n462 B.n36 585
R911 B.n461 B.n460 585
R912 B.n459 B.n37 585
R913 B.n458 B.n457 585
R914 B.n456 B.n38 585
R915 B.n455 B.n454 585
R916 B.n453 B.n39 585
R917 B.n452 B.n451 585
R918 B.n450 B.n40 585
R919 B.n449 B.n448 585
R920 B.n447 B.n41 585
R921 B.n446 B.n445 585
R922 B.n444 B.n45 585
R923 B.n443 B.n442 585
R924 B.n441 B.n46 585
R925 B.n440 B.n439 585
R926 B.n438 B.n47 585
R927 B.n437 B.n436 585
R928 B.n435 B.n48 585
R929 B.n434 B.n433 585
R930 B.n432 B.n49 585
R931 B.n431 B.n430 585
R932 B.n429 B.n50 585
R933 B.n428 B.n427 585
R934 B.n426 B.n51 585
R935 B.n425 B.n424 585
R936 B.n423 B.n52 585
R937 B.n422 B.n421 585
R938 B.n420 B.n53 585
R939 B.n419 B.n418 585
R940 B.n417 B.n54 585
R941 B.n416 B.n415 585
R942 B.n414 B.n55 585
R943 B.n413 B.n412 585
R944 B.n411 B.n56 585
R945 B.n410 B.n409 585
R946 B.n408 B.n57 585
R947 B.n407 B.n406 585
R948 B.n405 B.n58 585
R949 B.n404 B.n403 585
R950 B.n402 B.n59 585
R951 B.n401 B.n400 585
R952 B.n399 B.n60 585
R953 B.n398 B.n397 585
R954 B.n396 B.n61 585
R955 B.n520 B.n15 585
R956 B.n522 B.n521 585
R957 B.n523 B.n14 585
R958 B.n525 B.n524 585
R959 B.n526 B.n13 585
R960 B.n528 B.n527 585
R961 B.n529 B.n12 585
R962 B.n531 B.n530 585
R963 B.n532 B.n11 585
R964 B.n534 B.n533 585
R965 B.n535 B.n10 585
R966 B.n537 B.n536 585
R967 B.n538 B.n9 585
R968 B.n540 B.n539 585
R969 B.n541 B.n8 585
R970 B.n543 B.n542 585
R971 B.n544 B.n7 585
R972 B.n546 B.n545 585
R973 B.n547 B.n6 585
R974 B.n549 B.n548 585
R975 B.n550 B.n5 585
R976 B.n552 B.n551 585
R977 B.n553 B.n4 585
R978 B.n555 B.n554 585
R979 B.n556 B.n3 585
R980 B.n558 B.n557 585
R981 B.n559 B.n0 585
R982 B.n2 B.n1 585
R983 B.n146 B.n145 585
R984 B.n148 B.n147 585
R985 B.n149 B.n144 585
R986 B.n151 B.n150 585
R987 B.n152 B.n143 585
R988 B.n154 B.n153 585
R989 B.n155 B.n142 585
R990 B.n157 B.n156 585
R991 B.n158 B.n141 585
R992 B.n160 B.n159 585
R993 B.n161 B.n140 585
R994 B.n163 B.n162 585
R995 B.n164 B.n139 585
R996 B.n166 B.n165 585
R997 B.n167 B.n138 585
R998 B.n169 B.n168 585
R999 B.n170 B.n137 585
R1000 B.n172 B.n171 585
R1001 B.n173 B.n136 585
R1002 B.n175 B.n174 585
R1003 B.n176 B.n135 585
R1004 B.n178 B.n177 585
R1005 B.n179 B.n134 585
R1006 B.n181 B.n180 585
R1007 B.n182 B.n133 585
R1008 B.n184 B.n183 585
R1009 B.n183 B.n132 482.89
R1010 B.n312 B.n311 482.89
R1011 B.n396 B.n395 482.89
R1012 B.n518 B.n15 482.89
R1013 B.n113 B.t9 452.887
R1014 B.n253 B.t3 452.887
R1015 B.n42 B.t6 452.887
R1016 B.n34 B.t0 452.887
R1017 B.n253 B.t4 368.279
R1018 B.n42 B.t8 368.279
R1019 B.n113 B.t10 368.279
R1020 B.n34 B.t2 368.279
R1021 B.n254 B.t5 342.873
R1022 B.n43 B.t7 342.873
R1023 B.n114 B.t11 342.873
R1024 B.n35 B.t1 342.873
R1025 B.n561 B.n560 256.663
R1026 B.n560 B.n559 235.042
R1027 B.n560 B.n2 235.042
R1028 B.n187 B.n132 163.367
R1029 B.n188 B.n187 163.367
R1030 B.n189 B.n188 163.367
R1031 B.n189 B.n130 163.367
R1032 B.n193 B.n130 163.367
R1033 B.n194 B.n193 163.367
R1034 B.n195 B.n194 163.367
R1035 B.n195 B.n128 163.367
R1036 B.n199 B.n128 163.367
R1037 B.n200 B.n199 163.367
R1038 B.n201 B.n200 163.367
R1039 B.n201 B.n126 163.367
R1040 B.n205 B.n126 163.367
R1041 B.n206 B.n205 163.367
R1042 B.n207 B.n206 163.367
R1043 B.n207 B.n124 163.367
R1044 B.n211 B.n124 163.367
R1045 B.n212 B.n211 163.367
R1046 B.n213 B.n212 163.367
R1047 B.n213 B.n122 163.367
R1048 B.n217 B.n122 163.367
R1049 B.n218 B.n217 163.367
R1050 B.n219 B.n218 163.367
R1051 B.n219 B.n120 163.367
R1052 B.n223 B.n120 163.367
R1053 B.n224 B.n223 163.367
R1054 B.n225 B.n224 163.367
R1055 B.n225 B.n118 163.367
R1056 B.n229 B.n118 163.367
R1057 B.n230 B.n229 163.367
R1058 B.n231 B.n230 163.367
R1059 B.n231 B.n116 163.367
R1060 B.n235 B.n116 163.367
R1061 B.n236 B.n235 163.367
R1062 B.n237 B.n236 163.367
R1063 B.n237 B.n112 163.367
R1064 B.n242 B.n112 163.367
R1065 B.n243 B.n242 163.367
R1066 B.n244 B.n243 163.367
R1067 B.n244 B.n110 163.367
R1068 B.n248 B.n110 163.367
R1069 B.n249 B.n248 163.367
R1070 B.n250 B.n249 163.367
R1071 B.n250 B.n108 163.367
R1072 B.n257 B.n108 163.367
R1073 B.n258 B.n257 163.367
R1074 B.n259 B.n258 163.367
R1075 B.n259 B.n106 163.367
R1076 B.n263 B.n106 163.367
R1077 B.n264 B.n263 163.367
R1078 B.n265 B.n264 163.367
R1079 B.n265 B.n104 163.367
R1080 B.n269 B.n104 163.367
R1081 B.n270 B.n269 163.367
R1082 B.n271 B.n270 163.367
R1083 B.n271 B.n102 163.367
R1084 B.n275 B.n102 163.367
R1085 B.n276 B.n275 163.367
R1086 B.n277 B.n276 163.367
R1087 B.n277 B.n100 163.367
R1088 B.n281 B.n100 163.367
R1089 B.n282 B.n281 163.367
R1090 B.n283 B.n282 163.367
R1091 B.n283 B.n98 163.367
R1092 B.n287 B.n98 163.367
R1093 B.n288 B.n287 163.367
R1094 B.n289 B.n288 163.367
R1095 B.n289 B.n96 163.367
R1096 B.n293 B.n96 163.367
R1097 B.n294 B.n293 163.367
R1098 B.n295 B.n294 163.367
R1099 B.n295 B.n94 163.367
R1100 B.n299 B.n94 163.367
R1101 B.n300 B.n299 163.367
R1102 B.n301 B.n300 163.367
R1103 B.n301 B.n92 163.367
R1104 B.n305 B.n92 163.367
R1105 B.n306 B.n305 163.367
R1106 B.n307 B.n306 163.367
R1107 B.n307 B.n90 163.367
R1108 B.n311 B.n90 163.367
R1109 B.n395 B.n62 163.367
R1110 B.n391 B.n62 163.367
R1111 B.n391 B.n390 163.367
R1112 B.n390 B.n389 163.367
R1113 B.n389 B.n64 163.367
R1114 B.n385 B.n64 163.367
R1115 B.n385 B.n384 163.367
R1116 B.n384 B.n383 163.367
R1117 B.n383 B.n66 163.367
R1118 B.n379 B.n66 163.367
R1119 B.n379 B.n378 163.367
R1120 B.n378 B.n377 163.367
R1121 B.n377 B.n68 163.367
R1122 B.n373 B.n68 163.367
R1123 B.n373 B.n372 163.367
R1124 B.n372 B.n371 163.367
R1125 B.n371 B.n70 163.367
R1126 B.n367 B.n70 163.367
R1127 B.n367 B.n366 163.367
R1128 B.n366 B.n365 163.367
R1129 B.n365 B.n72 163.367
R1130 B.n361 B.n72 163.367
R1131 B.n361 B.n360 163.367
R1132 B.n360 B.n359 163.367
R1133 B.n359 B.n74 163.367
R1134 B.n355 B.n74 163.367
R1135 B.n355 B.n354 163.367
R1136 B.n354 B.n353 163.367
R1137 B.n353 B.n76 163.367
R1138 B.n349 B.n76 163.367
R1139 B.n349 B.n348 163.367
R1140 B.n348 B.n347 163.367
R1141 B.n347 B.n78 163.367
R1142 B.n343 B.n78 163.367
R1143 B.n343 B.n342 163.367
R1144 B.n342 B.n341 163.367
R1145 B.n341 B.n80 163.367
R1146 B.n337 B.n80 163.367
R1147 B.n337 B.n336 163.367
R1148 B.n336 B.n335 163.367
R1149 B.n335 B.n82 163.367
R1150 B.n331 B.n82 163.367
R1151 B.n331 B.n330 163.367
R1152 B.n330 B.n329 163.367
R1153 B.n329 B.n84 163.367
R1154 B.n325 B.n84 163.367
R1155 B.n325 B.n324 163.367
R1156 B.n324 B.n323 163.367
R1157 B.n323 B.n86 163.367
R1158 B.n319 B.n86 163.367
R1159 B.n319 B.n318 163.367
R1160 B.n318 B.n317 163.367
R1161 B.n317 B.n88 163.367
R1162 B.n313 B.n88 163.367
R1163 B.n313 B.n312 163.367
R1164 B.n518 B.n517 163.367
R1165 B.n517 B.n516 163.367
R1166 B.n516 B.n17 163.367
R1167 B.n512 B.n17 163.367
R1168 B.n512 B.n511 163.367
R1169 B.n511 B.n510 163.367
R1170 B.n510 B.n19 163.367
R1171 B.n506 B.n19 163.367
R1172 B.n506 B.n505 163.367
R1173 B.n505 B.n504 163.367
R1174 B.n504 B.n21 163.367
R1175 B.n500 B.n21 163.367
R1176 B.n500 B.n499 163.367
R1177 B.n499 B.n498 163.367
R1178 B.n498 B.n23 163.367
R1179 B.n494 B.n23 163.367
R1180 B.n494 B.n493 163.367
R1181 B.n493 B.n492 163.367
R1182 B.n492 B.n25 163.367
R1183 B.n488 B.n25 163.367
R1184 B.n488 B.n487 163.367
R1185 B.n487 B.n486 163.367
R1186 B.n486 B.n27 163.367
R1187 B.n482 B.n27 163.367
R1188 B.n482 B.n481 163.367
R1189 B.n481 B.n480 163.367
R1190 B.n480 B.n29 163.367
R1191 B.n476 B.n29 163.367
R1192 B.n476 B.n475 163.367
R1193 B.n475 B.n474 163.367
R1194 B.n474 B.n31 163.367
R1195 B.n470 B.n31 163.367
R1196 B.n470 B.n469 163.367
R1197 B.n469 B.n468 163.367
R1198 B.n468 B.n33 163.367
R1199 B.n463 B.n33 163.367
R1200 B.n463 B.n462 163.367
R1201 B.n462 B.n461 163.367
R1202 B.n461 B.n37 163.367
R1203 B.n457 B.n37 163.367
R1204 B.n457 B.n456 163.367
R1205 B.n456 B.n455 163.367
R1206 B.n455 B.n39 163.367
R1207 B.n451 B.n39 163.367
R1208 B.n451 B.n450 163.367
R1209 B.n450 B.n449 163.367
R1210 B.n449 B.n41 163.367
R1211 B.n445 B.n41 163.367
R1212 B.n445 B.n444 163.367
R1213 B.n444 B.n443 163.367
R1214 B.n443 B.n46 163.367
R1215 B.n439 B.n46 163.367
R1216 B.n439 B.n438 163.367
R1217 B.n438 B.n437 163.367
R1218 B.n437 B.n48 163.367
R1219 B.n433 B.n48 163.367
R1220 B.n433 B.n432 163.367
R1221 B.n432 B.n431 163.367
R1222 B.n431 B.n50 163.367
R1223 B.n427 B.n50 163.367
R1224 B.n427 B.n426 163.367
R1225 B.n426 B.n425 163.367
R1226 B.n425 B.n52 163.367
R1227 B.n421 B.n52 163.367
R1228 B.n421 B.n420 163.367
R1229 B.n420 B.n419 163.367
R1230 B.n419 B.n54 163.367
R1231 B.n415 B.n54 163.367
R1232 B.n415 B.n414 163.367
R1233 B.n414 B.n413 163.367
R1234 B.n413 B.n56 163.367
R1235 B.n409 B.n56 163.367
R1236 B.n409 B.n408 163.367
R1237 B.n408 B.n407 163.367
R1238 B.n407 B.n58 163.367
R1239 B.n403 B.n58 163.367
R1240 B.n403 B.n402 163.367
R1241 B.n402 B.n401 163.367
R1242 B.n401 B.n60 163.367
R1243 B.n397 B.n60 163.367
R1244 B.n397 B.n396 163.367
R1245 B.n522 B.n15 163.367
R1246 B.n523 B.n522 163.367
R1247 B.n524 B.n523 163.367
R1248 B.n524 B.n13 163.367
R1249 B.n528 B.n13 163.367
R1250 B.n529 B.n528 163.367
R1251 B.n530 B.n529 163.367
R1252 B.n530 B.n11 163.367
R1253 B.n534 B.n11 163.367
R1254 B.n535 B.n534 163.367
R1255 B.n536 B.n535 163.367
R1256 B.n536 B.n9 163.367
R1257 B.n540 B.n9 163.367
R1258 B.n541 B.n540 163.367
R1259 B.n542 B.n541 163.367
R1260 B.n542 B.n7 163.367
R1261 B.n546 B.n7 163.367
R1262 B.n547 B.n546 163.367
R1263 B.n548 B.n547 163.367
R1264 B.n548 B.n5 163.367
R1265 B.n552 B.n5 163.367
R1266 B.n553 B.n552 163.367
R1267 B.n554 B.n553 163.367
R1268 B.n554 B.n3 163.367
R1269 B.n558 B.n3 163.367
R1270 B.n559 B.n558 163.367
R1271 B.n146 B.n2 163.367
R1272 B.n147 B.n146 163.367
R1273 B.n147 B.n144 163.367
R1274 B.n151 B.n144 163.367
R1275 B.n152 B.n151 163.367
R1276 B.n153 B.n152 163.367
R1277 B.n153 B.n142 163.367
R1278 B.n157 B.n142 163.367
R1279 B.n158 B.n157 163.367
R1280 B.n159 B.n158 163.367
R1281 B.n159 B.n140 163.367
R1282 B.n163 B.n140 163.367
R1283 B.n164 B.n163 163.367
R1284 B.n165 B.n164 163.367
R1285 B.n165 B.n138 163.367
R1286 B.n169 B.n138 163.367
R1287 B.n170 B.n169 163.367
R1288 B.n171 B.n170 163.367
R1289 B.n171 B.n136 163.367
R1290 B.n175 B.n136 163.367
R1291 B.n176 B.n175 163.367
R1292 B.n177 B.n176 163.367
R1293 B.n177 B.n134 163.367
R1294 B.n181 B.n134 163.367
R1295 B.n182 B.n181 163.367
R1296 B.n183 B.n182 163.367
R1297 B.n239 B.n114 59.5399
R1298 B.n255 B.n254 59.5399
R1299 B.n44 B.n43 59.5399
R1300 B.n465 B.n35 59.5399
R1301 B.n520 B.n519 31.3761
R1302 B.n394 B.n61 31.3761
R1303 B.n310 B.n89 31.3761
R1304 B.n185 B.n184 31.3761
R1305 B.n114 B.n113 25.4066
R1306 B.n254 B.n253 25.4066
R1307 B.n43 B.n42 25.4066
R1308 B.n35 B.n34 25.4066
R1309 B B.n561 18.0485
R1310 B.n521 B.n520 10.6151
R1311 B.n521 B.n14 10.6151
R1312 B.n525 B.n14 10.6151
R1313 B.n526 B.n525 10.6151
R1314 B.n527 B.n526 10.6151
R1315 B.n527 B.n12 10.6151
R1316 B.n531 B.n12 10.6151
R1317 B.n532 B.n531 10.6151
R1318 B.n533 B.n532 10.6151
R1319 B.n533 B.n10 10.6151
R1320 B.n537 B.n10 10.6151
R1321 B.n538 B.n537 10.6151
R1322 B.n539 B.n538 10.6151
R1323 B.n539 B.n8 10.6151
R1324 B.n543 B.n8 10.6151
R1325 B.n544 B.n543 10.6151
R1326 B.n545 B.n544 10.6151
R1327 B.n545 B.n6 10.6151
R1328 B.n549 B.n6 10.6151
R1329 B.n550 B.n549 10.6151
R1330 B.n551 B.n550 10.6151
R1331 B.n551 B.n4 10.6151
R1332 B.n555 B.n4 10.6151
R1333 B.n556 B.n555 10.6151
R1334 B.n557 B.n556 10.6151
R1335 B.n557 B.n0 10.6151
R1336 B.n519 B.n16 10.6151
R1337 B.n515 B.n16 10.6151
R1338 B.n515 B.n514 10.6151
R1339 B.n514 B.n513 10.6151
R1340 B.n513 B.n18 10.6151
R1341 B.n509 B.n18 10.6151
R1342 B.n509 B.n508 10.6151
R1343 B.n508 B.n507 10.6151
R1344 B.n507 B.n20 10.6151
R1345 B.n503 B.n20 10.6151
R1346 B.n503 B.n502 10.6151
R1347 B.n502 B.n501 10.6151
R1348 B.n501 B.n22 10.6151
R1349 B.n497 B.n22 10.6151
R1350 B.n497 B.n496 10.6151
R1351 B.n496 B.n495 10.6151
R1352 B.n495 B.n24 10.6151
R1353 B.n491 B.n24 10.6151
R1354 B.n491 B.n490 10.6151
R1355 B.n490 B.n489 10.6151
R1356 B.n489 B.n26 10.6151
R1357 B.n485 B.n26 10.6151
R1358 B.n485 B.n484 10.6151
R1359 B.n484 B.n483 10.6151
R1360 B.n483 B.n28 10.6151
R1361 B.n479 B.n28 10.6151
R1362 B.n479 B.n478 10.6151
R1363 B.n478 B.n477 10.6151
R1364 B.n477 B.n30 10.6151
R1365 B.n473 B.n30 10.6151
R1366 B.n473 B.n472 10.6151
R1367 B.n472 B.n471 10.6151
R1368 B.n471 B.n32 10.6151
R1369 B.n467 B.n32 10.6151
R1370 B.n467 B.n466 10.6151
R1371 B.n464 B.n36 10.6151
R1372 B.n460 B.n36 10.6151
R1373 B.n460 B.n459 10.6151
R1374 B.n459 B.n458 10.6151
R1375 B.n458 B.n38 10.6151
R1376 B.n454 B.n38 10.6151
R1377 B.n454 B.n453 10.6151
R1378 B.n453 B.n452 10.6151
R1379 B.n452 B.n40 10.6151
R1380 B.n448 B.n447 10.6151
R1381 B.n447 B.n446 10.6151
R1382 B.n446 B.n45 10.6151
R1383 B.n442 B.n45 10.6151
R1384 B.n442 B.n441 10.6151
R1385 B.n441 B.n440 10.6151
R1386 B.n440 B.n47 10.6151
R1387 B.n436 B.n47 10.6151
R1388 B.n436 B.n435 10.6151
R1389 B.n435 B.n434 10.6151
R1390 B.n434 B.n49 10.6151
R1391 B.n430 B.n49 10.6151
R1392 B.n430 B.n429 10.6151
R1393 B.n429 B.n428 10.6151
R1394 B.n428 B.n51 10.6151
R1395 B.n424 B.n51 10.6151
R1396 B.n424 B.n423 10.6151
R1397 B.n423 B.n422 10.6151
R1398 B.n422 B.n53 10.6151
R1399 B.n418 B.n53 10.6151
R1400 B.n418 B.n417 10.6151
R1401 B.n417 B.n416 10.6151
R1402 B.n416 B.n55 10.6151
R1403 B.n412 B.n55 10.6151
R1404 B.n412 B.n411 10.6151
R1405 B.n411 B.n410 10.6151
R1406 B.n410 B.n57 10.6151
R1407 B.n406 B.n57 10.6151
R1408 B.n406 B.n405 10.6151
R1409 B.n405 B.n404 10.6151
R1410 B.n404 B.n59 10.6151
R1411 B.n400 B.n59 10.6151
R1412 B.n400 B.n399 10.6151
R1413 B.n399 B.n398 10.6151
R1414 B.n398 B.n61 10.6151
R1415 B.n394 B.n393 10.6151
R1416 B.n393 B.n392 10.6151
R1417 B.n392 B.n63 10.6151
R1418 B.n388 B.n63 10.6151
R1419 B.n388 B.n387 10.6151
R1420 B.n387 B.n386 10.6151
R1421 B.n386 B.n65 10.6151
R1422 B.n382 B.n65 10.6151
R1423 B.n382 B.n381 10.6151
R1424 B.n381 B.n380 10.6151
R1425 B.n380 B.n67 10.6151
R1426 B.n376 B.n67 10.6151
R1427 B.n376 B.n375 10.6151
R1428 B.n375 B.n374 10.6151
R1429 B.n374 B.n69 10.6151
R1430 B.n370 B.n69 10.6151
R1431 B.n370 B.n369 10.6151
R1432 B.n369 B.n368 10.6151
R1433 B.n368 B.n71 10.6151
R1434 B.n364 B.n71 10.6151
R1435 B.n364 B.n363 10.6151
R1436 B.n363 B.n362 10.6151
R1437 B.n362 B.n73 10.6151
R1438 B.n358 B.n73 10.6151
R1439 B.n358 B.n357 10.6151
R1440 B.n357 B.n356 10.6151
R1441 B.n356 B.n75 10.6151
R1442 B.n352 B.n75 10.6151
R1443 B.n352 B.n351 10.6151
R1444 B.n351 B.n350 10.6151
R1445 B.n350 B.n77 10.6151
R1446 B.n346 B.n77 10.6151
R1447 B.n346 B.n345 10.6151
R1448 B.n345 B.n344 10.6151
R1449 B.n344 B.n79 10.6151
R1450 B.n340 B.n79 10.6151
R1451 B.n340 B.n339 10.6151
R1452 B.n339 B.n338 10.6151
R1453 B.n338 B.n81 10.6151
R1454 B.n334 B.n81 10.6151
R1455 B.n334 B.n333 10.6151
R1456 B.n333 B.n332 10.6151
R1457 B.n332 B.n83 10.6151
R1458 B.n328 B.n83 10.6151
R1459 B.n328 B.n327 10.6151
R1460 B.n327 B.n326 10.6151
R1461 B.n326 B.n85 10.6151
R1462 B.n322 B.n85 10.6151
R1463 B.n322 B.n321 10.6151
R1464 B.n321 B.n320 10.6151
R1465 B.n320 B.n87 10.6151
R1466 B.n316 B.n87 10.6151
R1467 B.n316 B.n315 10.6151
R1468 B.n315 B.n314 10.6151
R1469 B.n314 B.n89 10.6151
R1470 B.n145 B.n1 10.6151
R1471 B.n148 B.n145 10.6151
R1472 B.n149 B.n148 10.6151
R1473 B.n150 B.n149 10.6151
R1474 B.n150 B.n143 10.6151
R1475 B.n154 B.n143 10.6151
R1476 B.n155 B.n154 10.6151
R1477 B.n156 B.n155 10.6151
R1478 B.n156 B.n141 10.6151
R1479 B.n160 B.n141 10.6151
R1480 B.n161 B.n160 10.6151
R1481 B.n162 B.n161 10.6151
R1482 B.n162 B.n139 10.6151
R1483 B.n166 B.n139 10.6151
R1484 B.n167 B.n166 10.6151
R1485 B.n168 B.n167 10.6151
R1486 B.n168 B.n137 10.6151
R1487 B.n172 B.n137 10.6151
R1488 B.n173 B.n172 10.6151
R1489 B.n174 B.n173 10.6151
R1490 B.n174 B.n135 10.6151
R1491 B.n178 B.n135 10.6151
R1492 B.n179 B.n178 10.6151
R1493 B.n180 B.n179 10.6151
R1494 B.n180 B.n133 10.6151
R1495 B.n184 B.n133 10.6151
R1496 B.n186 B.n185 10.6151
R1497 B.n186 B.n131 10.6151
R1498 B.n190 B.n131 10.6151
R1499 B.n191 B.n190 10.6151
R1500 B.n192 B.n191 10.6151
R1501 B.n192 B.n129 10.6151
R1502 B.n196 B.n129 10.6151
R1503 B.n197 B.n196 10.6151
R1504 B.n198 B.n197 10.6151
R1505 B.n198 B.n127 10.6151
R1506 B.n202 B.n127 10.6151
R1507 B.n203 B.n202 10.6151
R1508 B.n204 B.n203 10.6151
R1509 B.n204 B.n125 10.6151
R1510 B.n208 B.n125 10.6151
R1511 B.n209 B.n208 10.6151
R1512 B.n210 B.n209 10.6151
R1513 B.n210 B.n123 10.6151
R1514 B.n214 B.n123 10.6151
R1515 B.n215 B.n214 10.6151
R1516 B.n216 B.n215 10.6151
R1517 B.n216 B.n121 10.6151
R1518 B.n220 B.n121 10.6151
R1519 B.n221 B.n220 10.6151
R1520 B.n222 B.n221 10.6151
R1521 B.n222 B.n119 10.6151
R1522 B.n226 B.n119 10.6151
R1523 B.n227 B.n226 10.6151
R1524 B.n228 B.n227 10.6151
R1525 B.n228 B.n117 10.6151
R1526 B.n232 B.n117 10.6151
R1527 B.n233 B.n232 10.6151
R1528 B.n234 B.n233 10.6151
R1529 B.n234 B.n115 10.6151
R1530 B.n238 B.n115 10.6151
R1531 B.n241 B.n240 10.6151
R1532 B.n241 B.n111 10.6151
R1533 B.n245 B.n111 10.6151
R1534 B.n246 B.n245 10.6151
R1535 B.n247 B.n246 10.6151
R1536 B.n247 B.n109 10.6151
R1537 B.n251 B.n109 10.6151
R1538 B.n252 B.n251 10.6151
R1539 B.n256 B.n252 10.6151
R1540 B.n260 B.n107 10.6151
R1541 B.n261 B.n260 10.6151
R1542 B.n262 B.n261 10.6151
R1543 B.n262 B.n105 10.6151
R1544 B.n266 B.n105 10.6151
R1545 B.n267 B.n266 10.6151
R1546 B.n268 B.n267 10.6151
R1547 B.n268 B.n103 10.6151
R1548 B.n272 B.n103 10.6151
R1549 B.n273 B.n272 10.6151
R1550 B.n274 B.n273 10.6151
R1551 B.n274 B.n101 10.6151
R1552 B.n278 B.n101 10.6151
R1553 B.n279 B.n278 10.6151
R1554 B.n280 B.n279 10.6151
R1555 B.n280 B.n99 10.6151
R1556 B.n284 B.n99 10.6151
R1557 B.n285 B.n284 10.6151
R1558 B.n286 B.n285 10.6151
R1559 B.n286 B.n97 10.6151
R1560 B.n290 B.n97 10.6151
R1561 B.n291 B.n290 10.6151
R1562 B.n292 B.n291 10.6151
R1563 B.n292 B.n95 10.6151
R1564 B.n296 B.n95 10.6151
R1565 B.n297 B.n296 10.6151
R1566 B.n298 B.n297 10.6151
R1567 B.n298 B.n93 10.6151
R1568 B.n302 B.n93 10.6151
R1569 B.n303 B.n302 10.6151
R1570 B.n304 B.n303 10.6151
R1571 B.n304 B.n91 10.6151
R1572 B.n308 B.n91 10.6151
R1573 B.n309 B.n308 10.6151
R1574 B.n310 B.n309 10.6151
R1575 B.n466 B.n465 9.36635
R1576 B.n448 B.n44 9.36635
R1577 B.n239 B.n238 9.36635
R1578 B.n255 B.n107 9.36635
R1579 B.n561 B.n0 8.11757
R1580 B.n561 B.n1 8.11757
R1581 B.n465 B.n464 1.24928
R1582 B.n44 B.n40 1.24928
R1583 B.n240 B.n239 1.24928
R1584 B.n256 B.n255 1.24928
R1585 VN.n2 VN.t7 305.466
R1586 VN.n15 VN.t1 305.466
R1587 VN.n11 VN.t4 290.43
R1588 VN.n24 VN.t3 290.43
R1589 VN.n3 VN.t5 250.1
R1590 VN.n9 VN.t2 250.1
R1591 VN.n16 VN.t6 250.1
R1592 VN.n22 VN.t0 250.1
R1593 VN.n23 VN.n13 161.3
R1594 VN.n21 VN.n20 161.3
R1595 VN.n19 VN.n14 161.3
R1596 VN.n18 VN.n17 161.3
R1597 VN.n10 VN.n0 161.3
R1598 VN.n8 VN.n7 161.3
R1599 VN.n6 VN.n1 161.3
R1600 VN.n5 VN.n4 161.3
R1601 VN.n25 VN.n24 80.6037
R1602 VN.n12 VN.n11 80.6037
R1603 VN.n11 VN.n10 55.2959
R1604 VN.n24 VN.n23 55.2959
R1605 VN.n3 VN.n2 46.8653
R1606 VN.n16 VN.n15 46.8653
R1607 VN.n18 VN.n15 44.049
R1608 VN.n5 VN.n2 44.049
R1609 VN VN.n25 42.4006
R1610 VN.n4 VN.n1 40.4934
R1611 VN.n8 VN.n1 40.4934
R1612 VN.n17 VN.n14 40.4934
R1613 VN.n21 VN.n14 40.4934
R1614 VN.n10 VN.n9 16.8827
R1615 VN.n23 VN.n22 16.8827
R1616 VN.n4 VN.n3 7.58527
R1617 VN.n9 VN.n8 7.58527
R1618 VN.n17 VN.n16 7.58527
R1619 VN.n22 VN.n21 7.58527
R1620 VN.n25 VN.n13 0.285035
R1621 VN.n12 VN.n0 0.285035
R1622 VN.n20 VN.n13 0.189894
R1623 VN.n20 VN.n19 0.189894
R1624 VN.n19 VN.n18 0.189894
R1625 VN.n6 VN.n5 0.189894
R1626 VN.n7 VN.n6 0.189894
R1627 VN.n7 VN.n0 0.189894
R1628 VN VN.n12 0.146778
R1629 VDD2.n2 VDD2.n1 81.7008
R1630 VDD2.n2 VDD2.n0 81.7008
R1631 VDD2 VDD2.n5 81.698
R1632 VDD2.n4 VDD2.n3 81.1917
R1633 VDD2.n4 VDD2.n2 37.5644
R1634 VDD2.n5 VDD2.t1 3.19667
R1635 VDD2.n5 VDD2.t6 3.19667
R1636 VDD2.n3 VDD2.t4 3.19667
R1637 VDD2.n3 VDD2.t7 3.19667
R1638 VDD2.n1 VDD2.t5 3.19667
R1639 VDD2.n1 VDD2.t3 3.19667
R1640 VDD2.n0 VDD2.t0 3.19667
R1641 VDD2.n0 VDD2.t2 3.19667
R1642 VDD2 VDD2.n4 0.623345
C0 VDD1 VTAIL 8.53727f
C1 VP VTAIL 5.49425f
C2 VDD2 w_n2280_n3002# 1.40527f
C3 VN w_n2280_n3002# 4.15182f
C4 B w_n2280_n3002# 7.12275f
C5 VDD1 w_n2280_n3002# 1.35878f
C6 VP w_n2280_n3002# 4.443029f
C7 VN VDD2 5.52784f
C8 B VDD2 1.15159f
C9 VN B 0.825802f
C10 VTAIL w_n2280_n3002# 3.70841f
C11 VDD1 VDD2 0.966157f
C12 VDD1 VN 0.148851f
C13 VDD1 B 1.10627f
C14 VP VDD2 0.347337f
C15 VN VP 5.3418f
C16 VP B 1.30534f
C17 VDD1 VP 5.72575f
C18 VTAIL VDD2 8.580821f
C19 VN VTAIL 5.48014f
C20 B VTAIL 3.53895f
C21 VDD2 VSUBS 1.307353f
C22 VDD1 VSUBS 1.661378f
C23 VTAIL VSUBS 0.927299f
C24 VN VSUBS 4.79363f
C25 VP VSUBS 1.884199f
C26 B VSUBS 3.043378f
C27 w_n2280_n3002# VSUBS 84.515f
C28 VDD2.t0 VSUBS 0.208321f
C29 VDD2.t2 VSUBS 0.208321f
C30 VDD2.n0 VSUBS 1.59341f
C31 VDD2.t5 VSUBS 0.208321f
C32 VDD2.t3 VSUBS 0.208321f
C33 VDD2.n1 VSUBS 1.59341f
C34 VDD2.n2 VSUBS 2.79441f
C35 VDD2.t4 VSUBS 0.208321f
C36 VDD2.t7 VSUBS 0.208321f
C37 VDD2.n3 VSUBS 1.58964f
C38 VDD2.n4 VSUBS 2.573f
C39 VDD2.t1 VSUBS 0.208321f
C40 VDD2.t6 VSUBS 0.208321f
C41 VDD2.n5 VSUBS 1.59338f
C42 VN.n0 VSUBS 0.064607f
C43 VN.t2 VSUBS 1.30802f
C44 VN.n1 VSUBS 0.039141f
C45 VN.t7 VSUBS 1.40868f
C46 VN.n2 VSUBS 0.564099f
C47 VN.t5 VSUBS 1.30802f
C48 VN.n3 VSUBS 0.536683f
C49 VN.n4 VSUBS 0.065487f
C50 VN.n5 VSUBS 0.204906f
C51 VN.n6 VSUBS 0.048417f
C52 VN.n7 VSUBS 0.048417f
C53 VN.n8 VSUBS 0.065487f
C54 VN.n9 VSUBS 0.49533f
C55 VN.n10 VSUBS 0.064638f
C56 VN.t4 VSUBS 1.38072f
C57 VN.n11 VSUBS 0.567775f
C58 VN.n12 VSUBS 0.045345f
C59 VN.n13 VSUBS 0.064607f
C60 VN.t0 VSUBS 1.30802f
C61 VN.n14 VSUBS 0.039141f
C62 VN.t1 VSUBS 1.40868f
C63 VN.n15 VSUBS 0.564099f
C64 VN.t6 VSUBS 1.30802f
C65 VN.n16 VSUBS 0.536683f
C66 VN.n17 VSUBS 0.065487f
C67 VN.n18 VSUBS 0.204906f
C68 VN.n19 VSUBS 0.048417f
C69 VN.n20 VSUBS 0.048417f
C70 VN.n21 VSUBS 0.065487f
C71 VN.n22 VSUBS 0.49533f
C72 VN.n23 VSUBS 0.064638f
C73 VN.t3 VSUBS 1.38072f
C74 VN.n24 VSUBS 0.567775f
C75 VN.n25 VSUBS 2.05202f
C76 B.n0 VSUBS 0.007103f
C77 B.n1 VSUBS 0.007103f
C78 B.n2 VSUBS 0.010504f
C79 B.n3 VSUBS 0.00805f
C80 B.n4 VSUBS 0.00805f
C81 B.n5 VSUBS 0.00805f
C82 B.n6 VSUBS 0.00805f
C83 B.n7 VSUBS 0.00805f
C84 B.n8 VSUBS 0.00805f
C85 B.n9 VSUBS 0.00805f
C86 B.n10 VSUBS 0.00805f
C87 B.n11 VSUBS 0.00805f
C88 B.n12 VSUBS 0.00805f
C89 B.n13 VSUBS 0.00805f
C90 B.n14 VSUBS 0.00805f
C91 B.n15 VSUBS 0.017998f
C92 B.n16 VSUBS 0.00805f
C93 B.n17 VSUBS 0.00805f
C94 B.n18 VSUBS 0.00805f
C95 B.n19 VSUBS 0.00805f
C96 B.n20 VSUBS 0.00805f
C97 B.n21 VSUBS 0.00805f
C98 B.n22 VSUBS 0.00805f
C99 B.n23 VSUBS 0.00805f
C100 B.n24 VSUBS 0.00805f
C101 B.n25 VSUBS 0.00805f
C102 B.n26 VSUBS 0.00805f
C103 B.n27 VSUBS 0.00805f
C104 B.n28 VSUBS 0.00805f
C105 B.n29 VSUBS 0.00805f
C106 B.n30 VSUBS 0.00805f
C107 B.n31 VSUBS 0.00805f
C108 B.n32 VSUBS 0.00805f
C109 B.n33 VSUBS 0.00805f
C110 B.t1 VSUBS 0.197077f
C111 B.t2 VSUBS 0.213627f
C112 B.t0 VSUBS 0.490286f
C113 B.n34 VSUBS 0.327353f
C114 B.n35 VSUBS 0.251382f
C115 B.n36 VSUBS 0.00805f
C116 B.n37 VSUBS 0.00805f
C117 B.n38 VSUBS 0.00805f
C118 B.n39 VSUBS 0.00805f
C119 B.n40 VSUBS 0.004498f
C120 B.n41 VSUBS 0.00805f
C121 B.t7 VSUBS 0.197081f
C122 B.t8 VSUBS 0.21363f
C123 B.t6 VSUBS 0.490286f
C124 B.n42 VSUBS 0.32735f
C125 B.n43 VSUBS 0.251379f
C126 B.n44 VSUBS 0.01865f
C127 B.n45 VSUBS 0.00805f
C128 B.n46 VSUBS 0.00805f
C129 B.n47 VSUBS 0.00805f
C130 B.n48 VSUBS 0.00805f
C131 B.n49 VSUBS 0.00805f
C132 B.n50 VSUBS 0.00805f
C133 B.n51 VSUBS 0.00805f
C134 B.n52 VSUBS 0.00805f
C135 B.n53 VSUBS 0.00805f
C136 B.n54 VSUBS 0.00805f
C137 B.n55 VSUBS 0.00805f
C138 B.n56 VSUBS 0.00805f
C139 B.n57 VSUBS 0.00805f
C140 B.n58 VSUBS 0.00805f
C141 B.n59 VSUBS 0.00805f
C142 B.n60 VSUBS 0.00805f
C143 B.n61 VSUBS 0.018699f
C144 B.n62 VSUBS 0.00805f
C145 B.n63 VSUBS 0.00805f
C146 B.n64 VSUBS 0.00805f
C147 B.n65 VSUBS 0.00805f
C148 B.n66 VSUBS 0.00805f
C149 B.n67 VSUBS 0.00805f
C150 B.n68 VSUBS 0.00805f
C151 B.n69 VSUBS 0.00805f
C152 B.n70 VSUBS 0.00805f
C153 B.n71 VSUBS 0.00805f
C154 B.n72 VSUBS 0.00805f
C155 B.n73 VSUBS 0.00805f
C156 B.n74 VSUBS 0.00805f
C157 B.n75 VSUBS 0.00805f
C158 B.n76 VSUBS 0.00805f
C159 B.n77 VSUBS 0.00805f
C160 B.n78 VSUBS 0.00805f
C161 B.n79 VSUBS 0.00805f
C162 B.n80 VSUBS 0.00805f
C163 B.n81 VSUBS 0.00805f
C164 B.n82 VSUBS 0.00805f
C165 B.n83 VSUBS 0.00805f
C166 B.n84 VSUBS 0.00805f
C167 B.n85 VSUBS 0.00805f
C168 B.n86 VSUBS 0.00805f
C169 B.n87 VSUBS 0.00805f
C170 B.n88 VSUBS 0.00805f
C171 B.n89 VSUBS 0.018988f
C172 B.n90 VSUBS 0.00805f
C173 B.n91 VSUBS 0.00805f
C174 B.n92 VSUBS 0.00805f
C175 B.n93 VSUBS 0.00805f
C176 B.n94 VSUBS 0.00805f
C177 B.n95 VSUBS 0.00805f
C178 B.n96 VSUBS 0.00805f
C179 B.n97 VSUBS 0.00805f
C180 B.n98 VSUBS 0.00805f
C181 B.n99 VSUBS 0.00805f
C182 B.n100 VSUBS 0.00805f
C183 B.n101 VSUBS 0.00805f
C184 B.n102 VSUBS 0.00805f
C185 B.n103 VSUBS 0.00805f
C186 B.n104 VSUBS 0.00805f
C187 B.n105 VSUBS 0.00805f
C188 B.n106 VSUBS 0.00805f
C189 B.n107 VSUBS 0.007576f
C190 B.n108 VSUBS 0.00805f
C191 B.n109 VSUBS 0.00805f
C192 B.n110 VSUBS 0.00805f
C193 B.n111 VSUBS 0.00805f
C194 B.n112 VSUBS 0.00805f
C195 B.t11 VSUBS 0.197077f
C196 B.t10 VSUBS 0.213627f
C197 B.t9 VSUBS 0.490286f
C198 B.n113 VSUBS 0.327353f
C199 B.n114 VSUBS 0.251382f
C200 B.n115 VSUBS 0.00805f
C201 B.n116 VSUBS 0.00805f
C202 B.n117 VSUBS 0.00805f
C203 B.n118 VSUBS 0.00805f
C204 B.n119 VSUBS 0.00805f
C205 B.n120 VSUBS 0.00805f
C206 B.n121 VSUBS 0.00805f
C207 B.n122 VSUBS 0.00805f
C208 B.n123 VSUBS 0.00805f
C209 B.n124 VSUBS 0.00805f
C210 B.n125 VSUBS 0.00805f
C211 B.n126 VSUBS 0.00805f
C212 B.n127 VSUBS 0.00805f
C213 B.n128 VSUBS 0.00805f
C214 B.n129 VSUBS 0.00805f
C215 B.n130 VSUBS 0.00805f
C216 B.n131 VSUBS 0.00805f
C217 B.n132 VSUBS 0.018699f
C218 B.n133 VSUBS 0.00805f
C219 B.n134 VSUBS 0.00805f
C220 B.n135 VSUBS 0.00805f
C221 B.n136 VSUBS 0.00805f
C222 B.n137 VSUBS 0.00805f
C223 B.n138 VSUBS 0.00805f
C224 B.n139 VSUBS 0.00805f
C225 B.n140 VSUBS 0.00805f
C226 B.n141 VSUBS 0.00805f
C227 B.n142 VSUBS 0.00805f
C228 B.n143 VSUBS 0.00805f
C229 B.n144 VSUBS 0.00805f
C230 B.n145 VSUBS 0.00805f
C231 B.n146 VSUBS 0.00805f
C232 B.n147 VSUBS 0.00805f
C233 B.n148 VSUBS 0.00805f
C234 B.n149 VSUBS 0.00805f
C235 B.n150 VSUBS 0.00805f
C236 B.n151 VSUBS 0.00805f
C237 B.n152 VSUBS 0.00805f
C238 B.n153 VSUBS 0.00805f
C239 B.n154 VSUBS 0.00805f
C240 B.n155 VSUBS 0.00805f
C241 B.n156 VSUBS 0.00805f
C242 B.n157 VSUBS 0.00805f
C243 B.n158 VSUBS 0.00805f
C244 B.n159 VSUBS 0.00805f
C245 B.n160 VSUBS 0.00805f
C246 B.n161 VSUBS 0.00805f
C247 B.n162 VSUBS 0.00805f
C248 B.n163 VSUBS 0.00805f
C249 B.n164 VSUBS 0.00805f
C250 B.n165 VSUBS 0.00805f
C251 B.n166 VSUBS 0.00805f
C252 B.n167 VSUBS 0.00805f
C253 B.n168 VSUBS 0.00805f
C254 B.n169 VSUBS 0.00805f
C255 B.n170 VSUBS 0.00805f
C256 B.n171 VSUBS 0.00805f
C257 B.n172 VSUBS 0.00805f
C258 B.n173 VSUBS 0.00805f
C259 B.n174 VSUBS 0.00805f
C260 B.n175 VSUBS 0.00805f
C261 B.n176 VSUBS 0.00805f
C262 B.n177 VSUBS 0.00805f
C263 B.n178 VSUBS 0.00805f
C264 B.n179 VSUBS 0.00805f
C265 B.n180 VSUBS 0.00805f
C266 B.n181 VSUBS 0.00805f
C267 B.n182 VSUBS 0.00805f
C268 B.n183 VSUBS 0.017998f
C269 B.n184 VSUBS 0.017998f
C270 B.n185 VSUBS 0.018699f
C271 B.n186 VSUBS 0.00805f
C272 B.n187 VSUBS 0.00805f
C273 B.n188 VSUBS 0.00805f
C274 B.n189 VSUBS 0.00805f
C275 B.n190 VSUBS 0.00805f
C276 B.n191 VSUBS 0.00805f
C277 B.n192 VSUBS 0.00805f
C278 B.n193 VSUBS 0.00805f
C279 B.n194 VSUBS 0.00805f
C280 B.n195 VSUBS 0.00805f
C281 B.n196 VSUBS 0.00805f
C282 B.n197 VSUBS 0.00805f
C283 B.n198 VSUBS 0.00805f
C284 B.n199 VSUBS 0.00805f
C285 B.n200 VSUBS 0.00805f
C286 B.n201 VSUBS 0.00805f
C287 B.n202 VSUBS 0.00805f
C288 B.n203 VSUBS 0.00805f
C289 B.n204 VSUBS 0.00805f
C290 B.n205 VSUBS 0.00805f
C291 B.n206 VSUBS 0.00805f
C292 B.n207 VSUBS 0.00805f
C293 B.n208 VSUBS 0.00805f
C294 B.n209 VSUBS 0.00805f
C295 B.n210 VSUBS 0.00805f
C296 B.n211 VSUBS 0.00805f
C297 B.n212 VSUBS 0.00805f
C298 B.n213 VSUBS 0.00805f
C299 B.n214 VSUBS 0.00805f
C300 B.n215 VSUBS 0.00805f
C301 B.n216 VSUBS 0.00805f
C302 B.n217 VSUBS 0.00805f
C303 B.n218 VSUBS 0.00805f
C304 B.n219 VSUBS 0.00805f
C305 B.n220 VSUBS 0.00805f
C306 B.n221 VSUBS 0.00805f
C307 B.n222 VSUBS 0.00805f
C308 B.n223 VSUBS 0.00805f
C309 B.n224 VSUBS 0.00805f
C310 B.n225 VSUBS 0.00805f
C311 B.n226 VSUBS 0.00805f
C312 B.n227 VSUBS 0.00805f
C313 B.n228 VSUBS 0.00805f
C314 B.n229 VSUBS 0.00805f
C315 B.n230 VSUBS 0.00805f
C316 B.n231 VSUBS 0.00805f
C317 B.n232 VSUBS 0.00805f
C318 B.n233 VSUBS 0.00805f
C319 B.n234 VSUBS 0.00805f
C320 B.n235 VSUBS 0.00805f
C321 B.n236 VSUBS 0.00805f
C322 B.n237 VSUBS 0.00805f
C323 B.n238 VSUBS 0.007576f
C324 B.n239 VSUBS 0.01865f
C325 B.n240 VSUBS 0.004498f
C326 B.n241 VSUBS 0.00805f
C327 B.n242 VSUBS 0.00805f
C328 B.n243 VSUBS 0.00805f
C329 B.n244 VSUBS 0.00805f
C330 B.n245 VSUBS 0.00805f
C331 B.n246 VSUBS 0.00805f
C332 B.n247 VSUBS 0.00805f
C333 B.n248 VSUBS 0.00805f
C334 B.n249 VSUBS 0.00805f
C335 B.n250 VSUBS 0.00805f
C336 B.n251 VSUBS 0.00805f
C337 B.n252 VSUBS 0.00805f
C338 B.t5 VSUBS 0.197081f
C339 B.t4 VSUBS 0.21363f
C340 B.t3 VSUBS 0.490286f
C341 B.n253 VSUBS 0.32735f
C342 B.n254 VSUBS 0.251379f
C343 B.n255 VSUBS 0.01865f
C344 B.n256 VSUBS 0.004498f
C345 B.n257 VSUBS 0.00805f
C346 B.n258 VSUBS 0.00805f
C347 B.n259 VSUBS 0.00805f
C348 B.n260 VSUBS 0.00805f
C349 B.n261 VSUBS 0.00805f
C350 B.n262 VSUBS 0.00805f
C351 B.n263 VSUBS 0.00805f
C352 B.n264 VSUBS 0.00805f
C353 B.n265 VSUBS 0.00805f
C354 B.n266 VSUBS 0.00805f
C355 B.n267 VSUBS 0.00805f
C356 B.n268 VSUBS 0.00805f
C357 B.n269 VSUBS 0.00805f
C358 B.n270 VSUBS 0.00805f
C359 B.n271 VSUBS 0.00805f
C360 B.n272 VSUBS 0.00805f
C361 B.n273 VSUBS 0.00805f
C362 B.n274 VSUBS 0.00805f
C363 B.n275 VSUBS 0.00805f
C364 B.n276 VSUBS 0.00805f
C365 B.n277 VSUBS 0.00805f
C366 B.n278 VSUBS 0.00805f
C367 B.n279 VSUBS 0.00805f
C368 B.n280 VSUBS 0.00805f
C369 B.n281 VSUBS 0.00805f
C370 B.n282 VSUBS 0.00805f
C371 B.n283 VSUBS 0.00805f
C372 B.n284 VSUBS 0.00805f
C373 B.n285 VSUBS 0.00805f
C374 B.n286 VSUBS 0.00805f
C375 B.n287 VSUBS 0.00805f
C376 B.n288 VSUBS 0.00805f
C377 B.n289 VSUBS 0.00805f
C378 B.n290 VSUBS 0.00805f
C379 B.n291 VSUBS 0.00805f
C380 B.n292 VSUBS 0.00805f
C381 B.n293 VSUBS 0.00805f
C382 B.n294 VSUBS 0.00805f
C383 B.n295 VSUBS 0.00805f
C384 B.n296 VSUBS 0.00805f
C385 B.n297 VSUBS 0.00805f
C386 B.n298 VSUBS 0.00805f
C387 B.n299 VSUBS 0.00805f
C388 B.n300 VSUBS 0.00805f
C389 B.n301 VSUBS 0.00805f
C390 B.n302 VSUBS 0.00805f
C391 B.n303 VSUBS 0.00805f
C392 B.n304 VSUBS 0.00805f
C393 B.n305 VSUBS 0.00805f
C394 B.n306 VSUBS 0.00805f
C395 B.n307 VSUBS 0.00805f
C396 B.n308 VSUBS 0.00805f
C397 B.n309 VSUBS 0.00805f
C398 B.n310 VSUBS 0.017708f
C399 B.n311 VSUBS 0.018699f
C400 B.n312 VSUBS 0.017998f
C401 B.n313 VSUBS 0.00805f
C402 B.n314 VSUBS 0.00805f
C403 B.n315 VSUBS 0.00805f
C404 B.n316 VSUBS 0.00805f
C405 B.n317 VSUBS 0.00805f
C406 B.n318 VSUBS 0.00805f
C407 B.n319 VSUBS 0.00805f
C408 B.n320 VSUBS 0.00805f
C409 B.n321 VSUBS 0.00805f
C410 B.n322 VSUBS 0.00805f
C411 B.n323 VSUBS 0.00805f
C412 B.n324 VSUBS 0.00805f
C413 B.n325 VSUBS 0.00805f
C414 B.n326 VSUBS 0.00805f
C415 B.n327 VSUBS 0.00805f
C416 B.n328 VSUBS 0.00805f
C417 B.n329 VSUBS 0.00805f
C418 B.n330 VSUBS 0.00805f
C419 B.n331 VSUBS 0.00805f
C420 B.n332 VSUBS 0.00805f
C421 B.n333 VSUBS 0.00805f
C422 B.n334 VSUBS 0.00805f
C423 B.n335 VSUBS 0.00805f
C424 B.n336 VSUBS 0.00805f
C425 B.n337 VSUBS 0.00805f
C426 B.n338 VSUBS 0.00805f
C427 B.n339 VSUBS 0.00805f
C428 B.n340 VSUBS 0.00805f
C429 B.n341 VSUBS 0.00805f
C430 B.n342 VSUBS 0.00805f
C431 B.n343 VSUBS 0.00805f
C432 B.n344 VSUBS 0.00805f
C433 B.n345 VSUBS 0.00805f
C434 B.n346 VSUBS 0.00805f
C435 B.n347 VSUBS 0.00805f
C436 B.n348 VSUBS 0.00805f
C437 B.n349 VSUBS 0.00805f
C438 B.n350 VSUBS 0.00805f
C439 B.n351 VSUBS 0.00805f
C440 B.n352 VSUBS 0.00805f
C441 B.n353 VSUBS 0.00805f
C442 B.n354 VSUBS 0.00805f
C443 B.n355 VSUBS 0.00805f
C444 B.n356 VSUBS 0.00805f
C445 B.n357 VSUBS 0.00805f
C446 B.n358 VSUBS 0.00805f
C447 B.n359 VSUBS 0.00805f
C448 B.n360 VSUBS 0.00805f
C449 B.n361 VSUBS 0.00805f
C450 B.n362 VSUBS 0.00805f
C451 B.n363 VSUBS 0.00805f
C452 B.n364 VSUBS 0.00805f
C453 B.n365 VSUBS 0.00805f
C454 B.n366 VSUBS 0.00805f
C455 B.n367 VSUBS 0.00805f
C456 B.n368 VSUBS 0.00805f
C457 B.n369 VSUBS 0.00805f
C458 B.n370 VSUBS 0.00805f
C459 B.n371 VSUBS 0.00805f
C460 B.n372 VSUBS 0.00805f
C461 B.n373 VSUBS 0.00805f
C462 B.n374 VSUBS 0.00805f
C463 B.n375 VSUBS 0.00805f
C464 B.n376 VSUBS 0.00805f
C465 B.n377 VSUBS 0.00805f
C466 B.n378 VSUBS 0.00805f
C467 B.n379 VSUBS 0.00805f
C468 B.n380 VSUBS 0.00805f
C469 B.n381 VSUBS 0.00805f
C470 B.n382 VSUBS 0.00805f
C471 B.n383 VSUBS 0.00805f
C472 B.n384 VSUBS 0.00805f
C473 B.n385 VSUBS 0.00805f
C474 B.n386 VSUBS 0.00805f
C475 B.n387 VSUBS 0.00805f
C476 B.n388 VSUBS 0.00805f
C477 B.n389 VSUBS 0.00805f
C478 B.n390 VSUBS 0.00805f
C479 B.n391 VSUBS 0.00805f
C480 B.n392 VSUBS 0.00805f
C481 B.n393 VSUBS 0.00805f
C482 B.n394 VSUBS 0.017998f
C483 B.n395 VSUBS 0.017998f
C484 B.n396 VSUBS 0.018699f
C485 B.n397 VSUBS 0.00805f
C486 B.n398 VSUBS 0.00805f
C487 B.n399 VSUBS 0.00805f
C488 B.n400 VSUBS 0.00805f
C489 B.n401 VSUBS 0.00805f
C490 B.n402 VSUBS 0.00805f
C491 B.n403 VSUBS 0.00805f
C492 B.n404 VSUBS 0.00805f
C493 B.n405 VSUBS 0.00805f
C494 B.n406 VSUBS 0.00805f
C495 B.n407 VSUBS 0.00805f
C496 B.n408 VSUBS 0.00805f
C497 B.n409 VSUBS 0.00805f
C498 B.n410 VSUBS 0.00805f
C499 B.n411 VSUBS 0.00805f
C500 B.n412 VSUBS 0.00805f
C501 B.n413 VSUBS 0.00805f
C502 B.n414 VSUBS 0.00805f
C503 B.n415 VSUBS 0.00805f
C504 B.n416 VSUBS 0.00805f
C505 B.n417 VSUBS 0.00805f
C506 B.n418 VSUBS 0.00805f
C507 B.n419 VSUBS 0.00805f
C508 B.n420 VSUBS 0.00805f
C509 B.n421 VSUBS 0.00805f
C510 B.n422 VSUBS 0.00805f
C511 B.n423 VSUBS 0.00805f
C512 B.n424 VSUBS 0.00805f
C513 B.n425 VSUBS 0.00805f
C514 B.n426 VSUBS 0.00805f
C515 B.n427 VSUBS 0.00805f
C516 B.n428 VSUBS 0.00805f
C517 B.n429 VSUBS 0.00805f
C518 B.n430 VSUBS 0.00805f
C519 B.n431 VSUBS 0.00805f
C520 B.n432 VSUBS 0.00805f
C521 B.n433 VSUBS 0.00805f
C522 B.n434 VSUBS 0.00805f
C523 B.n435 VSUBS 0.00805f
C524 B.n436 VSUBS 0.00805f
C525 B.n437 VSUBS 0.00805f
C526 B.n438 VSUBS 0.00805f
C527 B.n439 VSUBS 0.00805f
C528 B.n440 VSUBS 0.00805f
C529 B.n441 VSUBS 0.00805f
C530 B.n442 VSUBS 0.00805f
C531 B.n443 VSUBS 0.00805f
C532 B.n444 VSUBS 0.00805f
C533 B.n445 VSUBS 0.00805f
C534 B.n446 VSUBS 0.00805f
C535 B.n447 VSUBS 0.00805f
C536 B.n448 VSUBS 0.007576f
C537 B.n449 VSUBS 0.00805f
C538 B.n450 VSUBS 0.00805f
C539 B.n451 VSUBS 0.00805f
C540 B.n452 VSUBS 0.00805f
C541 B.n453 VSUBS 0.00805f
C542 B.n454 VSUBS 0.00805f
C543 B.n455 VSUBS 0.00805f
C544 B.n456 VSUBS 0.00805f
C545 B.n457 VSUBS 0.00805f
C546 B.n458 VSUBS 0.00805f
C547 B.n459 VSUBS 0.00805f
C548 B.n460 VSUBS 0.00805f
C549 B.n461 VSUBS 0.00805f
C550 B.n462 VSUBS 0.00805f
C551 B.n463 VSUBS 0.00805f
C552 B.n464 VSUBS 0.004498f
C553 B.n465 VSUBS 0.01865f
C554 B.n466 VSUBS 0.007576f
C555 B.n467 VSUBS 0.00805f
C556 B.n468 VSUBS 0.00805f
C557 B.n469 VSUBS 0.00805f
C558 B.n470 VSUBS 0.00805f
C559 B.n471 VSUBS 0.00805f
C560 B.n472 VSUBS 0.00805f
C561 B.n473 VSUBS 0.00805f
C562 B.n474 VSUBS 0.00805f
C563 B.n475 VSUBS 0.00805f
C564 B.n476 VSUBS 0.00805f
C565 B.n477 VSUBS 0.00805f
C566 B.n478 VSUBS 0.00805f
C567 B.n479 VSUBS 0.00805f
C568 B.n480 VSUBS 0.00805f
C569 B.n481 VSUBS 0.00805f
C570 B.n482 VSUBS 0.00805f
C571 B.n483 VSUBS 0.00805f
C572 B.n484 VSUBS 0.00805f
C573 B.n485 VSUBS 0.00805f
C574 B.n486 VSUBS 0.00805f
C575 B.n487 VSUBS 0.00805f
C576 B.n488 VSUBS 0.00805f
C577 B.n489 VSUBS 0.00805f
C578 B.n490 VSUBS 0.00805f
C579 B.n491 VSUBS 0.00805f
C580 B.n492 VSUBS 0.00805f
C581 B.n493 VSUBS 0.00805f
C582 B.n494 VSUBS 0.00805f
C583 B.n495 VSUBS 0.00805f
C584 B.n496 VSUBS 0.00805f
C585 B.n497 VSUBS 0.00805f
C586 B.n498 VSUBS 0.00805f
C587 B.n499 VSUBS 0.00805f
C588 B.n500 VSUBS 0.00805f
C589 B.n501 VSUBS 0.00805f
C590 B.n502 VSUBS 0.00805f
C591 B.n503 VSUBS 0.00805f
C592 B.n504 VSUBS 0.00805f
C593 B.n505 VSUBS 0.00805f
C594 B.n506 VSUBS 0.00805f
C595 B.n507 VSUBS 0.00805f
C596 B.n508 VSUBS 0.00805f
C597 B.n509 VSUBS 0.00805f
C598 B.n510 VSUBS 0.00805f
C599 B.n511 VSUBS 0.00805f
C600 B.n512 VSUBS 0.00805f
C601 B.n513 VSUBS 0.00805f
C602 B.n514 VSUBS 0.00805f
C603 B.n515 VSUBS 0.00805f
C604 B.n516 VSUBS 0.00805f
C605 B.n517 VSUBS 0.00805f
C606 B.n518 VSUBS 0.018699f
C607 B.n519 VSUBS 0.018699f
C608 B.n520 VSUBS 0.017998f
C609 B.n521 VSUBS 0.00805f
C610 B.n522 VSUBS 0.00805f
C611 B.n523 VSUBS 0.00805f
C612 B.n524 VSUBS 0.00805f
C613 B.n525 VSUBS 0.00805f
C614 B.n526 VSUBS 0.00805f
C615 B.n527 VSUBS 0.00805f
C616 B.n528 VSUBS 0.00805f
C617 B.n529 VSUBS 0.00805f
C618 B.n530 VSUBS 0.00805f
C619 B.n531 VSUBS 0.00805f
C620 B.n532 VSUBS 0.00805f
C621 B.n533 VSUBS 0.00805f
C622 B.n534 VSUBS 0.00805f
C623 B.n535 VSUBS 0.00805f
C624 B.n536 VSUBS 0.00805f
C625 B.n537 VSUBS 0.00805f
C626 B.n538 VSUBS 0.00805f
C627 B.n539 VSUBS 0.00805f
C628 B.n540 VSUBS 0.00805f
C629 B.n541 VSUBS 0.00805f
C630 B.n542 VSUBS 0.00805f
C631 B.n543 VSUBS 0.00805f
C632 B.n544 VSUBS 0.00805f
C633 B.n545 VSUBS 0.00805f
C634 B.n546 VSUBS 0.00805f
C635 B.n547 VSUBS 0.00805f
C636 B.n548 VSUBS 0.00805f
C637 B.n549 VSUBS 0.00805f
C638 B.n550 VSUBS 0.00805f
C639 B.n551 VSUBS 0.00805f
C640 B.n552 VSUBS 0.00805f
C641 B.n553 VSUBS 0.00805f
C642 B.n554 VSUBS 0.00805f
C643 B.n555 VSUBS 0.00805f
C644 B.n556 VSUBS 0.00805f
C645 B.n557 VSUBS 0.00805f
C646 B.n558 VSUBS 0.00805f
C647 B.n559 VSUBS 0.010504f
C648 B.n560 VSUBS 0.01119f
C649 B.n561 VSUBS 0.022252f
C650 VTAIL.t7 VSUBS 0.200113f
C651 VTAIL.t4 VSUBS 0.200113f
C652 VTAIL.n0 VSUBS 1.41434f
C653 VTAIL.n1 VSUBS 0.61455f
C654 VTAIL.n2 VSUBS 0.028206f
C655 VTAIL.n3 VSUBS 0.0249f
C656 VTAIL.n4 VSUBS 0.01338f
C657 VTAIL.n5 VSUBS 0.031626f
C658 VTAIL.n6 VSUBS 0.014167f
C659 VTAIL.n7 VSUBS 0.0249f
C660 VTAIL.n8 VSUBS 0.013774f
C661 VTAIL.n9 VSUBS 0.031626f
C662 VTAIL.n10 VSUBS 0.014167f
C663 VTAIL.n11 VSUBS 0.0249f
C664 VTAIL.n12 VSUBS 0.01338f
C665 VTAIL.n13 VSUBS 0.031626f
C666 VTAIL.n14 VSUBS 0.014167f
C667 VTAIL.n15 VSUBS 0.0249f
C668 VTAIL.n16 VSUBS 0.01338f
C669 VTAIL.n17 VSUBS 0.023719f
C670 VTAIL.n18 VSUBS 0.023791f
C671 VTAIL.t6 VSUBS 0.068025f
C672 VTAIL.n19 VSUBS 0.175523f
C673 VTAIL.n20 VSUBS 1.02371f
C674 VTAIL.n21 VSUBS 0.01338f
C675 VTAIL.n22 VSUBS 0.014167f
C676 VTAIL.n23 VSUBS 0.031626f
C677 VTAIL.n24 VSUBS 0.031626f
C678 VTAIL.n25 VSUBS 0.014167f
C679 VTAIL.n26 VSUBS 0.01338f
C680 VTAIL.n27 VSUBS 0.0249f
C681 VTAIL.n28 VSUBS 0.0249f
C682 VTAIL.n29 VSUBS 0.01338f
C683 VTAIL.n30 VSUBS 0.014167f
C684 VTAIL.n31 VSUBS 0.031626f
C685 VTAIL.n32 VSUBS 0.031626f
C686 VTAIL.n33 VSUBS 0.014167f
C687 VTAIL.n34 VSUBS 0.01338f
C688 VTAIL.n35 VSUBS 0.0249f
C689 VTAIL.n36 VSUBS 0.0249f
C690 VTAIL.n37 VSUBS 0.01338f
C691 VTAIL.n38 VSUBS 0.01338f
C692 VTAIL.n39 VSUBS 0.014167f
C693 VTAIL.n40 VSUBS 0.031626f
C694 VTAIL.n41 VSUBS 0.031626f
C695 VTAIL.n42 VSUBS 0.031626f
C696 VTAIL.n43 VSUBS 0.013774f
C697 VTAIL.n44 VSUBS 0.01338f
C698 VTAIL.n45 VSUBS 0.0249f
C699 VTAIL.n46 VSUBS 0.0249f
C700 VTAIL.n47 VSUBS 0.01338f
C701 VTAIL.n48 VSUBS 0.014167f
C702 VTAIL.n49 VSUBS 0.031626f
C703 VTAIL.n50 VSUBS 0.079444f
C704 VTAIL.n51 VSUBS 0.014167f
C705 VTAIL.n52 VSUBS 0.01338f
C706 VTAIL.n53 VSUBS 0.064699f
C707 VTAIL.n54 VSUBS 0.040288f
C708 VTAIL.n55 VSUBS 0.153614f
C709 VTAIL.n56 VSUBS 0.028206f
C710 VTAIL.n57 VSUBS 0.0249f
C711 VTAIL.n58 VSUBS 0.01338f
C712 VTAIL.n59 VSUBS 0.031626f
C713 VTAIL.n60 VSUBS 0.014167f
C714 VTAIL.n61 VSUBS 0.0249f
C715 VTAIL.n62 VSUBS 0.013774f
C716 VTAIL.n63 VSUBS 0.031626f
C717 VTAIL.n64 VSUBS 0.014167f
C718 VTAIL.n65 VSUBS 0.0249f
C719 VTAIL.n66 VSUBS 0.01338f
C720 VTAIL.n67 VSUBS 0.031626f
C721 VTAIL.n68 VSUBS 0.014167f
C722 VTAIL.n69 VSUBS 0.0249f
C723 VTAIL.n70 VSUBS 0.01338f
C724 VTAIL.n71 VSUBS 0.023719f
C725 VTAIL.n72 VSUBS 0.023791f
C726 VTAIL.t10 VSUBS 0.068025f
C727 VTAIL.n73 VSUBS 0.175523f
C728 VTAIL.n74 VSUBS 1.02371f
C729 VTAIL.n75 VSUBS 0.01338f
C730 VTAIL.n76 VSUBS 0.014167f
C731 VTAIL.n77 VSUBS 0.031626f
C732 VTAIL.n78 VSUBS 0.031626f
C733 VTAIL.n79 VSUBS 0.014167f
C734 VTAIL.n80 VSUBS 0.01338f
C735 VTAIL.n81 VSUBS 0.0249f
C736 VTAIL.n82 VSUBS 0.0249f
C737 VTAIL.n83 VSUBS 0.01338f
C738 VTAIL.n84 VSUBS 0.014167f
C739 VTAIL.n85 VSUBS 0.031626f
C740 VTAIL.n86 VSUBS 0.031626f
C741 VTAIL.n87 VSUBS 0.014167f
C742 VTAIL.n88 VSUBS 0.01338f
C743 VTAIL.n89 VSUBS 0.0249f
C744 VTAIL.n90 VSUBS 0.0249f
C745 VTAIL.n91 VSUBS 0.01338f
C746 VTAIL.n92 VSUBS 0.01338f
C747 VTAIL.n93 VSUBS 0.014167f
C748 VTAIL.n94 VSUBS 0.031626f
C749 VTAIL.n95 VSUBS 0.031626f
C750 VTAIL.n96 VSUBS 0.031626f
C751 VTAIL.n97 VSUBS 0.013774f
C752 VTAIL.n98 VSUBS 0.01338f
C753 VTAIL.n99 VSUBS 0.0249f
C754 VTAIL.n100 VSUBS 0.0249f
C755 VTAIL.n101 VSUBS 0.01338f
C756 VTAIL.n102 VSUBS 0.014167f
C757 VTAIL.n103 VSUBS 0.031626f
C758 VTAIL.n104 VSUBS 0.079444f
C759 VTAIL.n105 VSUBS 0.014167f
C760 VTAIL.n106 VSUBS 0.01338f
C761 VTAIL.n107 VSUBS 0.064699f
C762 VTAIL.n108 VSUBS 0.040288f
C763 VTAIL.n109 VSUBS 0.153614f
C764 VTAIL.t12 VSUBS 0.200113f
C765 VTAIL.t9 VSUBS 0.200113f
C766 VTAIL.n110 VSUBS 1.41434f
C767 VTAIL.n111 VSUBS 0.70049f
C768 VTAIL.n112 VSUBS 0.028206f
C769 VTAIL.n113 VSUBS 0.0249f
C770 VTAIL.n114 VSUBS 0.01338f
C771 VTAIL.n115 VSUBS 0.031626f
C772 VTAIL.n116 VSUBS 0.014167f
C773 VTAIL.n117 VSUBS 0.0249f
C774 VTAIL.n118 VSUBS 0.013774f
C775 VTAIL.n119 VSUBS 0.031626f
C776 VTAIL.n120 VSUBS 0.014167f
C777 VTAIL.n121 VSUBS 0.0249f
C778 VTAIL.n122 VSUBS 0.01338f
C779 VTAIL.n123 VSUBS 0.031626f
C780 VTAIL.n124 VSUBS 0.014167f
C781 VTAIL.n125 VSUBS 0.0249f
C782 VTAIL.n126 VSUBS 0.01338f
C783 VTAIL.n127 VSUBS 0.023719f
C784 VTAIL.n128 VSUBS 0.023791f
C785 VTAIL.t11 VSUBS 0.068025f
C786 VTAIL.n129 VSUBS 0.175523f
C787 VTAIL.n130 VSUBS 1.02371f
C788 VTAIL.n131 VSUBS 0.01338f
C789 VTAIL.n132 VSUBS 0.014167f
C790 VTAIL.n133 VSUBS 0.031626f
C791 VTAIL.n134 VSUBS 0.031626f
C792 VTAIL.n135 VSUBS 0.014167f
C793 VTAIL.n136 VSUBS 0.01338f
C794 VTAIL.n137 VSUBS 0.0249f
C795 VTAIL.n138 VSUBS 0.0249f
C796 VTAIL.n139 VSUBS 0.01338f
C797 VTAIL.n140 VSUBS 0.014167f
C798 VTAIL.n141 VSUBS 0.031626f
C799 VTAIL.n142 VSUBS 0.031626f
C800 VTAIL.n143 VSUBS 0.014167f
C801 VTAIL.n144 VSUBS 0.01338f
C802 VTAIL.n145 VSUBS 0.0249f
C803 VTAIL.n146 VSUBS 0.0249f
C804 VTAIL.n147 VSUBS 0.01338f
C805 VTAIL.n148 VSUBS 0.01338f
C806 VTAIL.n149 VSUBS 0.014167f
C807 VTAIL.n150 VSUBS 0.031626f
C808 VTAIL.n151 VSUBS 0.031626f
C809 VTAIL.n152 VSUBS 0.031626f
C810 VTAIL.n153 VSUBS 0.013774f
C811 VTAIL.n154 VSUBS 0.01338f
C812 VTAIL.n155 VSUBS 0.0249f
C813 VTAIL.n156 VSUBS 0.0249f
C814 VTAIL.n157 VSUBS 0.01338f
C815 VTAIL.n158 VSUBS 0.014167f
C816 VTAIL.n159 VSUBS 0.031626f
C817 VTAIL.n160 VSUBS 0.079444f
C818 VTAIL.n161 VSUBS 0.014167f
C819 VTAIL.n162 VSUBS 0.01338f
C820 VTAIL.n163 VSUBS 0.064699f
C821 VTAIL.n164 VSUBS 0.040288f
C822 VTAIL.n165 VSUBS 1.24819f
C823 VTAIL.n166 VSUBS 0.028206f
C824 VTAIL.n167 VSUBS 0.0249f
C825 VTAIL.n168 VSUBS 0.01338f
C826 VTAIL.n169 VSUBS 0.031626f
C827 VTAIL.n170 VSUBS 0.014167f
C828 VTAIL.n171 VSUBS 0.0249f
C829 VTAIL.n172 VSUBS 0.013774f
C830 VTAIL.n173 VSUBS 0.031626f
C831 VTAIL.n174 VSUBS 0.01338f
C832 VTAIL.n175 VSUBS 0.014167f
C833 VTAIL.n176 VSUBS 0.0249f
C834 VTAIL.n177 VSUBS 0.01338f
C835 VTAIL.n178 VSUBS 0.031626f
C836 VTAIL.n179 VSUBS 0.014167f
C837 VTAIL.n180 VSUBS 0.0249f
C838 VTAIL.n181 VSUBS 0.01338f
C839 VTAIL.n182 VSUBS 0.023719f
C840 VTAIL.n183 VSUBS 0.023791f
C841 VTAIL.t3 VSUBS 0.068025f
C842 VTAIL.n184 VSUBS 0.175523f
C843 VTAIL.n185 VSUBS 1.02371f
C844 VTAIL.n186 VSUBS 0.01338f
C845 VTAIL.n187 VSUBS 0.014167f
C846 VTAIL.n188 VSUBS 0.031626f
C847 VTAIL.n189 VSUBS 0.031626f
C848 VTAIL.n190 VSUBS 0.014167f
C849 VTAIL.n191 VSUBS 0.01338f
C850 VTAIL.n192 VSUBS 0.0249f
C851 VTAIL.n193 VSUBS 0.0249f
C852 VTAIL.n194 VSUBS 0.01338f
C853 VTAIL.n195 VSUBS 0.014167f
C854 VTAIL.n196 VSUBS 0.031626f
C855 VTAIL.n197 VSUBS 0.031626f
C856 VTAIL.n198 VSUBS 0.014167f
C857 VTAIL.n199 VSUBS 0.01338f
C858 VTAIL.n200 VSUBS 0.0249f
C859 VTAIL.n201 VSUBS 0.0249f
C860 VTAIL.n202 VSUBS 0.01338f
C861 VTAIL.n203 VSUBS 0.014167f
C862 VTAIL.n204 VSUBS 0.031626f
C863 VTAIL.n205 VSUBS 0.031626f
C864 VTAIL.n206 VSUBS 0.031626f
C865 VTAIL.n207 VSUBS 0.013774f
C866 VTAIL.n208 VSUBS 0.01338f
C867 VTAIL.n209 VSUBS 0.0249f
C868 VTAIL.n210 VSUBS 0.0249f
C869 VTAIL.n211 VSUBS 0.01338f
C870 VTAIL.n212 VSUBS 0.014167f
C871 VTAIL.n213 VSUBS 0.031626f
C872 VTAIL.n214 VSUBS 0.079444f
C873 VTAIL.n215 VSUBS 0.014167f
C874 VTAIL.n216 VSUBS 0.01338f
C875 VTAIL.n217 VSUBS 0.064699f
C876 VTAIL.n218 VSUBS 0.040288f
C877 VTAIL.n219 VSUBS 1.24819f
C878 VTAIL.t0 VSUBS 0.200113f
C879 VTAIL.t2 VSUBS 0.200113f
C880 VTAIL.n220 VSUBS 1.41435f
C881 VTAIL.n221 VSUBS 0.700481f
C882 VTAIL.n222 VSUBS 0.028206f
C883 VTAIL.n223 VSUBS 0.0249f
C884 VTAIL.n224 VSUBS 0.01338f
C885 VTAIL.n225 VSUBS 0.031626f
C886 VTAIL.n226 VSUBS 0.014167f
C887 VTAIL.n227 VSUBS 0.0249f
C888 VTAIL.n228 VSUBS 0.013774f
C889 VTAIL.n229 VSUBS 0.031626f
C890 VTAIL.n230 VSUBS 0.01338f
C891 VTAIL.n231 VSUBS 0.014167f
C892 VTAIL.n232 VSUBS 0.0249f
C893 VTAIL.n233 VSUBS 0.01338f
C894 VTAIL.n234 VSUBS 0.031626f
C895 VTAIL.n235 VSUBS 0.014167f
C896 VTAIL.n236 VSUBS 0.0249f
C897 VTAIL.n237 VSUBS 0.01338f
C898 VTAIL.n238 VSUBS 0.023719f
C899 VTAIL.n239 VSUBS 0.023791f
C900 VTAIL.t5 VSUBS 0.068025f
C901 VTAIL.n240 VSUBS 0.175523f
C902 VTAIL.n241 VSUBS 1.02371f
C903 VTAIL.n242 VSUBS 0.01338f
C904 VTAIL.n243 VSUBS 0.014167f
C905 VTAIL.n244 VSUBS 0.031626f
C906 VTAIL.n245 VSUBS 0.031626f
C907 VTAIL.n246 VSUBS 0.014167f
C908 VTAIL.n247 VSUBS 0.01338f
C909 VTAIL.n248 VSUBS 0.0249f
C910 VTAIL.n249 VSUBS 0.0249f
C911 VTAIL.n250 VSUBS 0.01338f
C912 VTAIL.n251 VSUBS 0.014167f
C913 VTAIL.n252 VSUBS 0.031626f
C914 VTAIL.n253 VSUBS 0.031626f
C915 VTAIL.n254 VSUBS 0.014167f
C916 VTAIL.n255 VSUBS 0.01338f
C917 VTAIL.n256 VSUBS 0.0249f
C918 VTAIL.n257 VSUBS 0.0249f
C919 VTAIL.n258 VSUBS 0.01338f
C920 VTAIL.n259 VSUBS 0.014167f
C921 VTAIL.n260 VSUBS 0.031626f
C922 VTAIL.n261 VSUBS 0.031626f
C923 VTAIL.n262 VSUBS 0.031626f
C924 VTAIL.n263 VSUBS 0.013774f
C925 VTAIL.n264 VSUBS 0.01338f
C926 VTAIL.n265 VSUBS 0.0249f
C927 VTAIL.n266 VSUBS 0.0249f
C928 VTAIL.n267 VSUBS 0.01338f
C929 VTAIL.n268 VSUBS 0.014167f
C930 VTAIL.n269 VSUBS 0.031626f
C931 VTAIL.n270 VSUBS 0.079444f
C932 VTAIL.n271 VSUBS 0.014167f
C933 VTAIL.n272 VSUBS 0.01338f
C934 VTAIL.n273 VSUBS 0.064699f
C935 VTAIL.n274 VSUBS 0.040288f
C936 VTAIL.n275 VSUBS 0.153614f
C937 VTAIL.n276 VSUBS 0.028206f
C938 VTAIL.n277 VSUBS 0.0249f
C939 VTAIL.n278 VSUBS 0.01338f
C940 VTAIL.n279 VSUBS 0.031626f
C941 VTAIL.n280 VSUBS 0.014167f
C942 VTAIL.n281 VSUBS 0.0249f
C943 VTAIL.n282 VSUBS 0.013774f
C944 VTAIL.n283 VSUBS 0.031626f
C945 VTAIL.n284 VSUBS 0.01338f
C946 VTAIL.n285 VSUBS 0.014167f
C947 VTAIL.n286 VSUBS 0.0249f
C948 VTAIL.n287 VSUBS 0.01338f
C949 VTAIL.n288 VSUBS 0.031626f
C950 VTAIL.n289 VSUBS 0.014167f
C951 VTAIL.n290 VSUBS 0.0249f
C952 VTAIL.n291 VSUBS 0.01338f
C953 VTAIL.n292 VSUBS 0.023719f
C954 VTAIL.n293 VSUBS 0.023791f
C955 VTAIL.t15 VSUBS 0.068025f
C956 VTAIL.n294 VSUBS 0.175523f
C957 VTAIL.n295 VSUBS 1.02371f
C958 VTAIL.n296 VSUBS 0.01338f
C959 VTAIL.n297 VSUBS 0.014167f
C960 VTAIL.n298 VSUBS 0.031626f
C961 VTAIL.n299 VSUBS 0.031626f
C962 VTAIL.n300 VSUBS 0.014167f
C963 VTAIL.n301 VSUBS 0.01338f
C964 VTAIL.n302 VSUBS 0.0249f
C965 VTAIL.n303 VSUBS 0.0249f
C966 VTAIL.n304 VSUBS 0.01338f
C967 VTAIL.n305 VSUBS 0.014167f
C968 VTAIL.n306 VSUBS 0.031626f
C969 VTAIL.n307 VSUBS 0.031626f
C970 VTAIL.n308 VSUBS 0.014167f
C971 VTAIL.n309 VSUBS 0.01338f
C972 VTAIL.n310 VSUBS 0.0249f
C973 VTAIL.n311 VSUBS 0.0249f
C974 VTAIL.n312 VSUBS 0.01338f
C975 VTAIL.n313 VSUBS 0.014167f
C976 VTAIL.n314 VSUBS 0.031626f
C977 VTAIL.n315 VSUBS 0.031626f
C978 VTAIL.n316 VSUBS 0.031626f
C979 VTAIL.n317 VSUBS 0.013774f
C980 VTAIL.n318 VSUBS 0.01338f
C981 VTAIL.n319 VSUBS 0.0249f
C982 VTAIL.n320 VSUBS 0.0249f
C983 VTAIL.n321 VSUBS 0.01338f
C984 VTAIL.n322 VSUBS 0.014167f
C985 VTAIL.n323 VSUBS 0.031626f
C986 VTAIL.n324 VSUBS 0.079444f
C987 VTAIL.n325 VSUBS 0.014167f
C988 VTAIL.n326 VSUBS 0.01338f
C989 VTAIL.n327 VSUBS 0.064699f
C990 VTAIL.n328 VSUBS 0.040288f
C991 VTAIL.n329 VSUBS 0.153614f
C992 VTAIL.t13 VSUBS 0.200113f
C993 VTAIL.t8 VSUBS 0.200113f
C994 VTAIL.n330 VSUBS 1.41435f
C995 VTAIL.n331 VSUBS 0.700481f
C996 VTAIL.n332 VSUBS 0.028206f
C997 VTAIL.n333 VSUBS 0.0249f
C998 VTAIL.n334 VSUBS 0.01338f
C999 VTAIL.n335 VSUBS 0.031626f
C1000 VTAIL.n336 VSUBS 0.014167f
C1001 VTAIL.n337 VSUBS 0.0249f
C1002 VTAIL.n338 VSUBS 0.013774f
C1003 VTAIL.n339 VSUBS 0.031626f
C1004 VTAIL.n340 VSUBS 0.01338f
C1005 VTAIL.n341 VSUBS 0.014167f
C1006 VTAIL.n342 VSUBS 0.0249f
C1007 VTAIL.n343 VSUBS 0.01338f
C1008 VTAIL.n344 VSUBS 0.031626f
C1009 VTAIL.n345 VSUBS 0.014167f
C1010 VTAIL.n346 VSUBS 0.0249f
C1011 VTAIL.n347 VSUBS 0.01338f
C1012 VTAIL.n348 VSUBS 0.023719f
C1013 VTAIL.n349 VSUBS 0.023791f
C1014 VTAIL.t14 VSUBS 0.068025f
C1015 VTAIL.n350 VSUBS 0.175523f
C1016 VTAIL.n351 VSUBS 1.02371f
C1017 VTAIL.n352 VSUBS 0.01338f
C1018 VTAIL.n353 VSUBS 0.014167f
C1019 VTAIL.n354 VSUBS 0.031626f
C1020 VTAIL.n355 VSUBS 0.031626f
C1021 VTAIL.n356 VSUBS 0.014167f
C1022 VTAIL.n357 VSUBS 0.01338f
C1023 VTAIL.n358 VSUBS 0.0249f
C1024 VTAIL.n359 VSUBS 0.0249f
C1025 VTAIL.n360 VSUBS 0.01338f
C1026 VTAIL.n361 VSUBS 0.014167f
C1027 VTAIL.n362 VSUBS 0.031626f
C1028 VTAIL.n363 VSUBS 0.031626f
C1029 VTAIL.n364 VSUBS 0.014167f
C1030 VTAIL.n365 VSUBS 0.01338f
C1031 VTAIL.n366 VSUBS 0.0249f
C1032 VTAIL.n367 VSUBS 0.0249f
C1033 VTAIL.n368 VSUBS 0.01338f
C1034 VTAIL.n369 VSUBS 0.014167f
C1035 VTAIL.n370 VSUBS 0.031626f
C1036 VTAIL.n371 VSUBS 0.031626f
C1037 VTAIL.n372 VSUBS 0.031626f
C1038 VTAIL.n373 VSUBS 0.013774f
C1039 VTAIL.n374 VSUBS 0.01338f
C1040 VTAIL.n375 VSUBS 0.0249f
C1041 VTAIL.n376 VSUBS 0.0249f
C1042 VTAIL.n377 VSUBS 0.01338f
C1043 VTAIL.n378 VSUBS 0.014167f
C1044 VTAIL.n379 VSUBS 0.031626f
C1045 VTAIL.n380 VSUBS 0.079444f
C1046 VTAIL.n381 VSUBS 0.014167f
C1047 VTAIL.n382 VSUBS 0.01338f
C1048 VTAIL.n383 VSUBS 0.064699f
C1049 VTAIL.n384 VSUBS 0.040288f
C1050 VTAIL.n385 VSUBS 1.24819f
C1051 VTAIL.n386 VSUBS 0.028206f
C1052 VTAIL.n387 VSUBS 0.0249f
C1053 VTAIL.n388 VSUBS 0.01338f
C1054 VTAIL.n389 VSUBS 0.031626f
C1055 VTAIL.n390 VSUBS 0.014167f
C1056 VTAIL.n391 VSUBS 0.0249f
C1057 VTAIL.n392 VSUBS 0.013774f
C1058 VTAIL.n393 VSUBS 0.031626f
C1059 VTAIL.n394 VSUBS 0.014167f
C1060 VTAIL.n395 VSUBS 0.0249f
C1061 VTAIL.n396 VSUBS 0.01338f
C1062 VTAIL.n397 VSUBS 0.031626f
C1063 VTAIL.n398 VSUBS 0.014167f
C1064 VTAIL.n399 VSUBS 0.0249f
C1065 VTAIL.n400 VSUBS 0.01338f
C1066 VTAIL.n401 VSUBS 0.023719f
C1067 VTAIL.n402 VSUBS 0.023791f
C1068 VTAIL.t1 VSUBS 0.068025f
C1069 VTAIL.n403 VSUBS 0.175523f
C1070 VTAIL.n404 VSUBS 1.02371f
C1071 VTAIL.n405 VSUBS 0.01338f
C1072 VTAIL.n406 VSUBS 0.014167f
C1073 VTAIL.n407 VSUBS 0.031626f
C1074 VTAIL.n408 VSUBS 0.031626f
C1075 VTAIL.n409 VSUBS 0.014167f
C1076 VTAIL.n410 VSUBS 0.01338f
C1077 VTAIL.n411 VSUBS 0.0249f
C1078 VTAIL.n412 VSUBS 0.0249f
C1079 VTAIL.n413 VSUBS 0.01338f
C1080 VTAIL.n414 VSUBS 0.014167f
C1081 VTAIL.n415 VSUBS 0.031626f
C1082 VTAIL.n416 VSUBS 0.031626f
C1083 VTAIL.n417 VSUBS 0.014167f
C1084 VTAIL.n418 VSUBS 0.01338f
C1085 VTAIL.n419 VSUBS 0.0249f
C1086 VTAIL.n420 VSUBS 0.0249f
C1087 VTAIL.n421 VSUBS 0.01338f
C1088 VTAIL.n422 VSUBS 0.01338f
C1089 VTAIL.n423 VSUBS 0.014167f
C1090 VTAIL.n424 VSUBS 0.031626f
C1091 VTAIL.n425 VSUBS 0.031626f
C1092 VTAIL.n426 VSUBS 0.031626f
C1093 VTAIL.n427 VSUBS 0.013774f
C1094 VTAIL.n428 VSUBS 0.01338f
C1095 VTAIL.n429 VSUBS 0.0249f
C1096 VTAIL.n430 VSUBS 0.0249f
C1097 VTAIL.n431 VSUBS 0.01338f
C1098 VTAIL.n432 VSUBS 0.014167f
C1099 VTAIL.n433 VSUBS 0.031626f
C1100 VTAIL.n434 VSUBS 0.079444f
C1101 VTAIL.n435 VSUBS 0.014167f
C1102 VTAIL.n436 VSUBS 0.01338f
C1103 VTAIL.n437 VSUBS 0.064699f
C1104 VTAIL.n438 VSUBS 0.040288f
C1105 VTAIL.n439 VSUBS 1.24352f
C1106 VDD1.t7 VSUBS 0.208383f
C1107 VDD1.t5 VSUBS 0.208383f
C1108 VDD1.n0 VSUBS 1.5948f
C1109 VDD1.t2 VSUBS 0.208383f
C1110 VDD1.t1 VSUBS 0.208383f
C1111 VDD1.n1 VSUBS 1.59389f
C1112 VDD1.t6 VSUBS 0.208383f
C1113 VDD1.t0 VSUBS 0.208383f
C1114 VDD1.n2 VSUBS 1.59389f
C1115 VDD1.n3 VSUBS 2.85044f
C1116 VDD1.t3 VSUBS 0.208383f
C1117 VDD1.t4 VSUBS 0.208383f
C1118 VDD1.n4 VSUBS 1.59011f
C1119 VDD1.n5 VSUBS 2.60463f
C1120 VP.n0 VSUBS 0.066087f
C1121 VP.t6 VSUBS 1.33799f
C1122 VP.n1 VSUBS 0.040038f
C1123 VP.n2 VSUBS 0.066087f
C1124 VP.t3 VSUBS 1.33799f
C1125 VP.n3 VSUBS 0.066087f
C1126 VP.t1 VSUBS 1.41235f
C1127 VP.t7 VSUBS 1.33799f
C1128 VP.n4 VSUBS 0.040038f
C1129 VP.t0 VSUBS 1.44095f
C1130 VP.n5 VSUBS 0.577021f
C1131 VP.t2 VSUBS 1.33799f
C1132 VP.n6 VSUBS 0.548978f
C1133 VP.n7 VSUBS 0.066987f
C1134 VP.n8 VSUBS 0.2096f
C1135 VP.n9 VSUBS 0.049526f
C1136 VP.n10 VSUBS 0.049526f
C1137 VP.n11 VSUBS 0.066987f
C1138 VP.n12 VSUBS 0.506677f
C1139 VP.n13 VSUBS 0.066119f
C1140 VP.n14 VSUBS 0.580781f
C1141 VP.n15 VSUBS 2.07126f
C1142 VP.n16 VSUBS 2.11353f
C1143 VP.t4 VSUBS 1.41235f
C1144 VP.n17 VSUBS 0.580781f
C1145 VP.n18 VSUBS 0.066119f
C1146 VP.n19 VSUBS 0.506677f
C1147 VP.n20 VSUBS 0.066987f
C1148 VP.n21 VSUBS 0.049526f
C1149 VP.n22 VSUBS 0.049526f
C1150 VP.n23 VSUBS 0.049526f
C1151 VP.n24 VSUBS 0.066987f
C1152 VP.n25 VSUBS 0.506677f
C1153 VP.n26 VSUBS 0.066119f
C1154 VP.t5 VSUBS 1.41235f
C1155 VP.n27 VSUBS 0.580781f
C1156 VP.n28 VSUBS 0.046384f
.ends

